module basic_750_5000_1000_5_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_582,In_145);
or U1 (N_1,In_15,In_82);
and U2 (N_2,In_556,In_429);
nand U3 (N_3,In_632,In_127);
nand U4 (N_4,In_741,In_560);
or U5 (N_5,In_409,In_45);
or U6 (N_6,In_514,In_184);
nor U7 (N_7,In_364,In_72);
and U8 (N_8,In_618,In_320);
and U9 (N_9,In_506,In_368);
and U10 (N_10,In_236,In_118);
nor U11 (N_11,In_695,In_14);
nand U12 (N_12,In_32,In_74);
or U13 (N_13,In_546,In_119);
nand U14 (N_14,In_259,In_331);
nor U15 (N_15,In_473,In_54);
and U16 (N_16,In_636,In_410);
xor U17 (N_17,In_722,In_126);
xnor U18 (N_18,In_624,In_716);
or U19 (N_19,In_438,In_165);
or U20 (N_20,In_372,In_69);
nand U21 (N_21,In_691,In_466);
and U22 (N_22,In_218,In_665);
nor U23 (N_23,In_278,In_534);
xnor U24 (N_24,In_73,In_591);
nor U25 (N_25,In_8,In_196);
nand U26 (N_26,In_672,In_204);
and U27 (N_27,In_106,In_551);
and U28 (N_28,In_22,In_192);
or U29 (N_29,In_562,In_412);
xnor U30 (N_30,In_290,In_205);
xor U31 (N_31,In_676,In_497);
nand U32 (N_32,In_443,In_326);
xor U33 (N_33,In_345,In_155);
nand U34 (N_34,In_311,In_219);
or U35 (N_35,In_46,In_356);
nor U36 (N_36,In_605,In_511);
nor U37 (N_37,In_365,In_85);
xnor U38 (N_38,In_325,In_697);
and U39 (N_39,In_130,In_708);
xnor U40 (N_40,In_474,In_226);
or U41 (N_41,In_629,In_689);
xor U42 (N_42,In_44,In_59);
nand U43 (N_43,In_210,In_554);
nor U44 (N_44,In_314,In_682);
nor U45 (N_45,In_454,In_743);
and U46 (N_46,In_688,In_673);
nand U47 (N_47,In_488,In_481);
xor U48 (N_48,In_84,In_542);
or U49 (N_49,In_283,In_735);
and U50 (N_50,In_467,In_492);
and U51 (N_51,In_586,In_262);
xor U52 (N_52,In_243,In_104);
or U53 (N_53,In_726,In_515);
and U54 (N_54,In_424,In_107);
nor U55 (N_55,In_384,In_723);
nor U56 (N_56,In_423,In_298);
or U57 (N_57,In_241,In_164);
nor U58 (N_58,In_745,In_569);
nor U59 (N_59,In_646,In_92);
nand U60 (N_60,In_707,In_96);
and U61 (N_61,In_389,In_416);
xnor U62 (N_62,In_195,In_437);
and U63 (N_63,In_614,In_472);
nand U64 (N_64,In_299,In_304);
xnor U65 (N_65,In_110,In_491);
or U66 (N_66,In_150,In_622);
and U67 (N_67,In_198,In_575);
nand U68 (N_68,In_124,In_264);
or U69 (N_69,In_432,In_200);
nor U70 (N_70,In_538,In_272);
nor U71 (N_71,In_584,In_293);
nor U72 (N_72,In_201,In_17);
and U73 (N_73,In_237,In_539);
nand U74 (N_74,In_394,In_163);
nand U75 (N_75,In_238,In_690);
or U76 (N_76,In_434,In_611);
nand U77 (N_77,In_3,In_616);
nand U78 (N_78,In_38,In_683);
nand U79 (N_79,In_520,In_197);
and U80 (N_80,In_49,In_21);
nor U81 (N_81,In_144,In_700);
or U82 (N_82,In_220,In_711);
xor U83 (N_83,In_216,In_271);
nand U84 (N_84,In_313,In_292);
or U85 (N_85,In_308,In_40);
nor U86 (N_86,In_6,In_340);
xnor U87 (N_87,In_567,In_570);
and U88 (N_88,In_390,In_425);
nor U89 (N_89,In_373,In_275);
and U90 (N_90,In_9,In_536);
xor U91 (N_91,In_53,In_407);
nor U92 (N_92,In_746,In_213);
and U93 (N_93,In_561,In_628);
xor U94 (N_94,In_666,In_337);
and U95 (N_95,In_300,In_451);
xnor U96 (N_96,In_18,In_194);
or U97 (N_97,In_51,In_79);
nor U98 (N_98,In_181,In_43);
xnor U99 (N_99,In_258,In_422);
or U100 (N_100,In_86,In_612);
or U101 (N_101,In_552,In_510);
or U102 (N_102,In_327,In_146);
or U103 (N_103,In_129,In_81);
xnor U104 (N_104,In_744,In_495);
and U105 (N_105,In_95,In_670);
xor U106 (N_106,In_535,In_55);
and U107 (N_107,In_202,In_214);
and U108 (N_108,In_75,In_475);
nand U109 (N_109,In_553,In_532);
xnor U110 (N_110,In_228,In_247);
or U111 (N_111,In_504,In_633);
nand U112 (N_112,In_693,In_329);
xnor U113 (N_113,In_459,In_748);
nand U114 (N_114,In_349,In_717);
or U115 (N_115,In_668,In_125);
or U116 (N_116,In_548,In_608);
nor U117 (N_117,In_169,In_244);
and U118 (N_118,In_317,In_427);
nand U119 (N_119,In_193,In_659);
and U120 (N_120,In_12,In_421);
nand U121 (N_121,In_479,In_25);
xnor U122 (N_122,In_477,In_48);
or U123 (N_123,In_112,In_348);
or U124 (N_124,In_580,In_732);
xor U125 (N_125,In_530,In_179);
and U126 (N_126,In_378,In_211);
or U127 (N_127,In_650,In_186);
or U128 (N_128,In_11,In_286);
xnor U129 (N_129,In_660,In_159);
or U130 (N_130,In_120,In_638);
and U131 (N_131,In_5,In_602);
or U132 (N_132,In_157,In_573);
nor U133 (N_133,In_328,In_235);
or U134 (N_134,In_692,In_625);
nand U135 (N_135,In_122,In_566);
or U136 (N_136,In_486,In_720);
xor U137 (N_137,In_585,In_440);
and U138 (N_138,In_139,In_623);
or U139 (N_139,In_724,In_170);
nor U140 (N_140,In_102,In_590);
nor U141 (N_141,In_382,In_305);
nor U142 (N_142,In_65,In_607);
nor U143 (N_143,In_10,In_600);
xnor U144 (N_144,In_154,In_281);
nor U145 (N_145,In_316,In_199);
nor U146 (N_146,In_563,In_249);
xnor U147 (N_147,In_674,In_503);
or U148 (N_148,In_583,In_370);
xor U149 (N_149,In_469,In_100);
nor U150 (N_150,In_62,In_435);
or U151 (N_151,In_675,In_89);
nor U152 (N_152,In_288,In_606);
nand U153 (N_153,In_94,In_557);
or U154 (N_154,In_136,In_285);
or U155 (N_155,In_547,In_703);
nor U156 (N_156,In_667,In_677);
xor U157 (N_157,In_452,In_725);
and U158 (N_158,In_315,In_684);
nor U159 (N_159,In_284,In_77);
xor U160 (N_160,In_191,In_734);
nor U161 (N_161,In_489,In_704);
and U162 (N_162,In_428,In_696);
nor U163 (N_163,In_635,In_577);
and U164 (N_164,In_270,In_453);
and U165 (N_165,In_521,In_90);
nor U166 (N_166,In_685,In_56);
or U167 (N_167,In_496,In_307);
nor U168 (N_168,In_217,In_559);
xor U169 (N_169,In_721,In_261);
xor U170 (N_170,In_401,In_571);
or U171 (N_171,In_587,In_621);
nor U172 (N_172,In_652,In_265);
xnor U173 (N_173,In_468,In_168);
or U174 (N_174,In_76,In_442);
nor U175 (N_175,In_52,In_729);
nor U176 (N_176,In_63,In_543);
nand U177 (N_177,In_318,In_594);
xnor U178 (N_178,In_341,In_111);
or U179 (N_179,In_456,In_309);
nand U180 (N_180,In_680,In_206);
xor U181 (N_181,In_291,In_246);
nor U182 (N_182,In_524,In_487);
or U183 (N_183,In_742,In_29);
nor U184 (N_184,In_297,In_253);
and U185 (N_185,In_493,In_256);
or U186 (N_186,In_36,In_531);
and U187 (N_187,In_257,In_678);
xor U188 (N_188,In_446,In_572);
nor U189 (N_189,In_537,In_502);
or U190 (N_190,In_333,In_395);
nand U191 (N_191,In_108,In_215);
xor U192 (N_192,In_183,In_354);
and U193 (N_193,In_248,In_371);
nor U194 (N_194,In_60,In_457);
nor U195 (N_195,In_706,In_67);
or U196 (N_196,In_355,In_174);
nor U197 (N_197,In_224,In_545);
and U198 (N_198,In_91,In_519);
or U199 (N_199,In_156,In_718);
nand U200 (N_200,In_361,In_233);
nor U201 (N_201,In_705,In_109);
xnor U202 (N_202,In_282,In_458);
nor U203 (N_203,In_448,In_417);
and U204 (N_204,In_363,In_701);
xnor U205 (N_205,In_588,In_604);
and U206 (N_206,In_113,In_737);
nand U207 (N_207,In_686,In_230);
and U208 (N_208,In_358,In_509);
nand U209 (N_209,In_399,In_431);
xnor U210 (N_210,In_66,In_330);
and U211 (N_211,In_544,In_287);
nand U212 (N_212,In_596,In_630);
and U213 (N_213,In_523,In_252);
nand U214 (N_214,In_242,In_518);
nor U215 (N_215,In_657,In_388);
and U216 (N_216,In_460,In_739);
and U217 (N_217,In_478,In_221);
or U218 (N_218,In_500,In_450);
and U219 (N_219,In_362,In_263);
nand U220 (N_220,In_517,In_494);
and U221 (N_221,In_637,In_80);
nand U222 (N_222,In_47,In_749);
nor U223 (N_223,In_88,In_490);
xnor U224 (N_224,In_411,In_426);
xor U225 (N_225,In_610,In_171);
nand U226 (N_226,In_369,In_232);
xor U227 (N_227,In_393,In_461);
and U228 (N_228,In_603,In_240);
nand U229 (N_229,In_574,In_462);
and U230 (N_230,In_87,In_656);
nor U231 (N_231,In_267,In_375);
and U232 (N_232,In_335,In_351);
or U233 (N_233,In_643,In_26);
and U234 (N_234,In_280,In_30);
nand U235 (N_235,In_34,In_499);
or U236 (N_236,In_182,In_642);
nor U237 (N_237,In_589,In_508);
nand U238 (N_238,In_255,In_507);
nor U239 (N_239,In_415,In_408);
or U240 (N_240,In_463,In_114);
or U241 (N_241,In_640,In_480);
xnor U242 (N_242,In_344,In_27);
nor U243 (N_243,In_250,In_631);
nor U244 (N_244,In_302,In_301);
xnor U245 (N_245,In_387,In_28);
and U246 (N_246,In_296,In_702);
and U247 (N_247,In_208,In_445);
nor U248 (N_248,In_550,In_135);
nor U249 (N_249,In_592,In_151);
and U250 (N_250,In_42,In_68);
xor U251 (N_251,In_449,In_484);
or U252 (N_252,In_687,In_529);
and U253 (N_253,In_649,In_276);
or U254 (N_254,In_339,In_143);
xnor U255 (N_255,In_279,In_360);
or U256 (N_256,In_324,In_190);
nand U257 (N_257,In_441,In_541);
or U258 (N_258,In_180,In_57);
or U259 (N_259,In_597,In_414);
nor U260 (N_260,In_347,In_471);
xnor U261 (N_261,In_392,In_715);
xnor U262 (N_262,In_679,In_343);
nand U263 (N_263,In_698,In_131);
nor U264 (N_264,In_430,In_483);
nor U265 (N_265,In_533,In_303);
nor U266 (N_266,In_403,In_598);
or U267 (N_267,In_385,In_20);
xor U268 (N_268,In_465,In_172);
nand U269 (N_269,In_319,In_227);
and U270 (N_270,In_641,In_138);
xor U271 (N_271,In_476,In_386);
nor U272 (N_272,In_234,In_615);
and U273 (N_273,In_260,In_16);
and U274 (N_274,In_418,In_485);
nand U275 (N_275,In_555,In_397);
xnor U276 (N_276,In_223,In_207);
or U277 (N_277,In_398,In_439);
nand U278 (N_278,In_322,In_39);
or U279 (N_279,In_274,In_142);
nand U280 (N_280,In_176,In_37);
and U281 (N_281,In_133,In_661);
nand U282 (N_282,In_160,In_400);
nor U283 (N_283,In_404,In_99);
and U284 (N_284,In_728,In_1);
xor U285 (N_285,In_647,In_336);
and U286 (N_286,In_70,In_455);
nor U287 (N_287,In_105,In_187);
or U288 (N_288,In_312,In_644);
nor U289 (N_289,In_482,In_527);
nand U290 (N_290,In_357,In_153);
xor U291 (N_291,In_501,In_645);
xnor U292 (N_292,In_595,In_498);
or U293 (N_293,In_391,In_712);
nor U294 (N_294,In_576,In_374);
and U295 (N_295,In_103,In_681);
nor U296 (N_296,In_323,In_13);
xor U297 (N_297,In_19,In_413);
or U298 (N_298,In_350,In_101);
nand U299 (N_299,In_188,In_352);
nand U300 (N_300,In_121,In_377);
or U301 (N_301,In_83,In_627);
xnor U302 (N_302,In_134,In_671);
nor U303 (N_303,In_332,In_558);
xor U304 (N_304,In_620,In_225);
xor U305 (N_305,In_212,In_117);
or U306 (N_306,In_626,In_599);
or U307 (N_307,In_710,In_166);
nand U308 (N_308,In_733,In_222);
and U309 (N_309,In_366,In_376);
nand U310 (N_310,In_123,In_526);
or U311 (N_311,In_185,In_116);
nand U312 (N_312,In_653,In_41);
or U313 (N_313,In_229,In_50);
or U314 (N_314,In_310,In_346);
nor U315 (N_315,In_564,In_420);
xor U316 (N_316,In_231,In_173);
or U317 (N_317,In_7,In_512);
nor U318 (N_318,In_464,In_669);
xnor U319 (N_319,In_406,In_664);
xor U320 (N_320,In_266,In_731);
nor U321 (N_321,In_0,In_209);
nor U322 (N_322,In_175,In_64);
nand U323 (N_323,In_565,In_152);
or U324 (N_324,In_662,In_31);
nor U325 (N_325,In_730,In_23);
xor U326 (N_326,In_132,In_540);
nor U327 (N_327,In_699,In_289);
xor U328 (N_328,In_203,In_161);
xor U329 (N_329,In_522,In_433);
nand U330 (N_330,In_342,In_71);
nor U331 (N_331,In_334,In_359);
nand U332 (N_332,In_613,In_609);
nand U333 (N_333,In_601,In_239);
nand U334 (N_334,In_58,In_367);
or U335 (N_335,In_747,In_713);
xor U336 (N_336,In_269,In_516);
xnor U337 (N_337,In_137,In_141);
nor U338 (N_338,In_245,In_578);
or U339 (N_339,In_189,In_98);
and U340 (N_340,In_419,In_727);
nor U341 (N_341,In_177,In_97);
nor U342 (N_342,In_648,In_405);
xor U343 (N_343,In_380,In_651);
nand U344 (N_344,In_617,In_549);
nor U345 (N_345,In_738,In_306);
xnor U346 (N_346,In_93,In_149);
nor U347 (N_347,In_436,In_148);
nand U348 (N_348,In_277,In_634);
xnor U349 (N_349,In_402,In_295);
and U350 (N_350,In_251,In_78);
and U351 (N_351,In_528,In_694);
xnor U352 (N_352,In_663,In_709);
nand U353 (N_353,In_654,In_568);
and U354 (N_354,In_353,In_35);
nand U355 (N_355,In_61,In_24);
nor U356 (N_356,In_655,In_4);
nor U357 (N_357,In_470,In_639);
nand U358 (N_358,In_167,In_2);
xnor U359 (N_359,In_740,In_513);
xnor U360 (N_360,In_714,In_719);
or U361 (N_361,In_140,In_147);
xnor U362 (N_362,In_658,In_505);
or U363 (N_363,In_383,In_447);
and U364 (N_364,In_736,In_593);
nand U365 (N_365,In_444,In_525);
nor U366 (N_366,In_619,In_115);
nand U367 (N_367,In_294,In_158);
nor U368 (N_368,In_379,In_254);
xor U369 (N_369,In_128,In_381);
nor U370 (N_370,In_581,In_273);
xnor U371 (N_371,In_579,In_33);
or U372 (N_372,In_321,In_162);
xnor U373 (N_373,In_338,In_268);
nand U374 (N_374,In_396,In_178);
nand U375 (N_375,In_227,In_344);
xor U376 (N_376,In_72,In_547);
or U377 (N_377,In_485,In_237);
nand U378 (N_378,In_724,In_250);
or U379 (N_379,In_180,In_390);
and U380 (N_380,In_382,In_516);
nor U381 (N_381,In_124,In_157);
nor U382 (N_382,In_553,In_147);
nor U383 (N_383,In_667,In_197);
xnor U384 (N_384,In_711,In_84);
or U385 (N_385,In_467,In_169);
nor U386 (N_386,In_275,In_197);
and U387 (N_387,In_561,In_670);
or U388 (N_388,In_244,In_606);
nand U389 (N_389,In_674,In_161);
or U390 (N_390,In_415,In_466);
nor U391 (N_391,In_81,In_396);
or U392 (N_392,In_348,In_415);
nor U393 (N_393,In_743,In_519);
nor U394 (N_394,In_509,In_712);
xor U395 (N_395,In_199,In_484);
and U396 (N_396,In_262,In_297);
nor U397 (N_397,In_347,In_212);
nor U398 (N_398,In_537,In_550);
nand U399 (N_399,In_97,In_700);
and U400 (N_400,In_10,In_68);
nand U401 (N_401,In_288,In_643);
or U402 (N_402,In_631,In_493);
nand U403 (N_403,In_373,In_7);
and U404 (N_404,In_319,In_138);
nand U405 (N_405,In_655,In_571);
nand U406 (N_406,In_355,In_562);
xnor U407 (N_407,In_662,In_79);
or U408 (N_408,In_566,In_291);
xor U409 (N_409,In_604,In_748);
or U410 (N_410,In_235,In_384);
and U411 (N_411,In_338,In_684);
or U412 (N_412,In_480,In_719);
nand U413 (N_413,In_154,In_425);
nor U414 (N_414,In_538,In_89);
xor U415 (N_415,In_679,In_380);
or U416 (N_416,In_152,In_134);
nor U417 (N_417,In_495,In_400);
or U418 (N_418,In_453,In_642);
nand U419 (N_419,In_664,In_119);
xnor U420 (N_420,In_740,In_454);
nand U421 (N_421,In_193,In_96);
or U422 (N_422,In_656,In_109);
or U423 (N_423,In_681,In_227);
or U424 (N_424,In_136,In_29);
nor U425 (N_425,In_564,In_321);
nand U426 (N_426,In_282,In_157);
and U427 (N_427,In_372,In_386);
and U428 (N_428,In_643,In_227);
and U429 (N_429,In_610,In_434);
or U430 (N_430,In_203,In_200);
and U431 (N_431,In_483,In_63);
nand U432 (N_432,In_386,In_430);
nor U433 (N_433,In_354,In_639);
nand U434 (N_434,In_391,In_398);
or U435 (N_435,In_418,In_742);
or U436 (N_436,In_697,In_297);
nand U437 (N_437,In_126,In_324);
nor U438 (N_438,In_88,In_57);
nor U439 (N_439,In_163,In_413);
and U440 (N_440,In_143,In_458);
nand U441 (N_441,In_74,In_42);
or U442 (N_442,In_705,In_222);
or U443 (N_443,In_276,In_464);
or U444 (N_444,In_146,In_294);
xnor U445 (N_445,In_504,In_636);
xor U446 (N_446,In_271,In_125);
nor U447 (N_447,In_437,In_516);
nand U448 (N_448,In_318,In_611);
nor U449 (N_449,In_410,In_454);
nand U450 (N_450,In_138,In_654);
nand U451 (N_451,In_264,In_302);
and U452 (N_452,In_252,In_377);
and U453 (N_453,In_609,In_125);
and U454 (N_454,In_301,In_528);
nand U455 (N_455,In_599,In_187);
or U456 (N_456,In_316,In_723);
nand U457 (N_457,In_727,In_586);
xor U458 (N_458,In_437,In_537);
nor U459 (N_459,In_437,In_193);
and U460 (N_460,In_6,In_253);
and U461 (N_461,In_528,In_462);
or U462 (N_462,In_346,In_344);
and U463 (N_463,In_21,In_326);
and U464 (N_464,In_256,In_421);
and U465 (N_465,In_227,In_339);
xnor U466 (N_466,In_614,In_664);
xor U467 (N_467,In_716,In_268);
and U468 (N_468,In_426,In_242);
nor U469 (N_469,In_749,In_86);
or U470 (N_470,In_62,In_294);
and U471 (N_471,In_671,In_199);
xor U472 (N_472,In_167,In_463);
nor U473 (N_473,In_661,In_42);
or U474 (N_474,In_404,In_218);
xnor U475 (N_475,In_480,In_34);
or U476 (N_476,In_534,In_568);
and U477 (N_477,In_208,In_166);
and U478 (N_478,In_45,In_27);
nand U479 (N_479,In_596,In_504);
nand U480 (N_480,In_484,In_350);
nor U481 (N_481,In_497,In_345);
nor U482 (N_482,In_29,In_330);
or U483 (N_483,In_557,In_263);
and U484 (N_484,In_743,In_172);
nand U485 (N_485,In_96,In_491);
xnor U486 (N_486,In_592,In_51);
nor U487 (N_487,In_270,In_210);
nor U488 (N_488,In_453,In_160);
or U489 (N_489,In_226,In_342);
nand U490 (N_490,In_192,In_182);
nand U491 (N_491,In_92,In_33);
nor U492 (N_492,In_112,In_2);
or U493 (N_493,In_133,In_716);
or U494 (N_494,In_35,In_663);
and U495 (N_495,In_44,In_310);
and U496 (N_496,In_657,In_584);
or U497 (N_497,In_300,In_229);
xnor U498 (N_498,In_55,In_160);
xnor U499 (N_499,In_201,In_244);
nor U500 (N_500,In_165,In_627);
nor U501 (N_501,In_320,In_732);
nor U502 (N_502,In_112,In_192);
or U503 (N_503,In_305,In_631);
nand U504 (N_504,In_720,In_662);
or U505 (N_505,In_23,In_10);
nand U506 (N_506,In_97,In_688);
nor U507 (N_507,In_491,In_222);
xor U508 (N_508,In_716,In_176);
nor U509 (N_509,In_532,In_392);
or U510 (N_510,In_675,In_115);
or U511 (N_511,In_126,In_690);
xor U512 (N_512,In_717,In_632);
nand U513 (N_513,In_407,In_654);
or U514 (N_514,In_602,In_435);
nor U515 (N_515,In_169,In_441);
nor U516 (N_516,In_416,In_340);
nand U517 (N_517,In_430,In_315);
nand U518 (N_518,In_383,In_549);
nor U519 (N_519,In_140,In_607);
nor U520 (N_520,In_537,In_518);
and U521 (N_521,In_717,In_76);
or U522 (N_522,In_552,In_611);
and U523 (N_523,In_207,In_642);
or U524 (N_524,In_459,In_352);
nand U525 (N_525,In_588,In_720);
nand U526 (N_526,In_697,In_8);
or U527 (N_527,In_30,In_658);
xor U528 (N_528,In_598,In_168);
and U529 (N_529,In_468,In_145);
xnor U530 (N_530,In_470,In_325);
xnor U531 (N_531,In_120,In_714);
nor U532 (N_532,In_25,In_653);
nand U533 (N_533,In_139,In_711);
xor U534 (N_534,In_308,In_294);
xor U535 (N_535,In_478,In_557);
and U536 (N_536,In_275,In_613);
and U537 (N_537,In_68,In_210);
xnor U538 (N_538,In_335,In_611);
xor U539 (N_539,In_345,In_628);
nand U540 (N_540,In_706,In_232);
nand U541 (N_541,In_434,In_101);
or U542 (N_542,In_415,In_707);
nor U543 (N_543,In_142,In_437);
or U544 (N_544,In_256,In_659);
nand U545 (N_545,In_26,In_447);
or U546 (N_546,In_735,In_56);
and U547 (N_547,In_123,In_601);
xor U548 (N_548,In_508,In_748);
and U549 (N_549,In_49,In_689);
and U550 (N_550,In_359,In_66);
nand U551 (N_551,In_629,In_239);
and U552 (N_552,In_63,In_220);
nand U553 (N_553,In_472,In_424);
and U554 (N_554,In_528,In_655);
nor U555 (N_555,In_722,In_171);
and U556 (N_556,In_428,In_137);
or U557 (N_557,In_36,In_42);
nor U558 (N_558,In_482,In_706);
nand U559 (N_559,In_613,In_540);
nand U560 (N_560,In_408,In_16);
and U561 (N_561,In_530,In_155);
or U562 (N_562,In_722,In_402);
xor U563 (N_563,In_463,In_581);
and U564 (N_564,In_586,In_188);
nor U565 (N_565,In_664,In_23);
nor U566 (N_566,In_162,In_452);
or U567 (N_567,In_637,In_356);
or U568 (N_568,In_661,In_348);
xor U569 (N_569,In_543,In_77);
or U570 (N_570,In_506,In_133);
and U571 (N_571,In_721,In_623);
and U572 (N_572,In_356,In_7);
or U573 (N_573,In_563,In_620);
or U574 (N_574,In_495,In_425);
xor U575 (N_575,In_1,In_241);
nor U576 (N_576,In_0,In_60);
xnor U577 (N_577,In_57,In_430);
nor U578 (N_578,In_28,In_20);
and U579 (N_579,In_497,In_530);
xor U580 (N_580,In_205,In_719);
and U581 (N_581,In_645,In_653);
or U582 (N_582,In_320,In_354);
or U583 (N_583,In_694,In_302);
and U584 (N_584,In_122,In_725);
nand U585 (N_585,In_732,In_323);
or U586 (N_586,In_313,In_239);
nand U587 (N_587,In_398,In_670);
nand U588 (N_588,In_111,In_332);
nor U589 (N_589,In_3,In_539);
nor U590 (N_590,In_409,In_64);
or U591 (N_591,In_51,In_688);
and U592 (N_592,In_728,In_111);
and U593 (N_593,In_241,In_17);
nand U594 (N_594,In_744,In_91);
nor U595 (N_595,In_733,In_415);
nand U596 (N_596,In_98,In_266);
or U597 (N_597,In_480,In_471);
xor U598 (N_598,In_687,In_172);
xnor U599 (N_599,In_665,In_705);
or U600 (N_600,In_51,In_485);
xor U601 (N_601,In_714,In_404);
nor U602 (N_602,In_440,In_430);
or U603 (N_603,In_253,In_103);
xor U604 (N_604,In_331,In_478);
and U605 (N_605,In_121,In_562);
and U606 (N_606,In_111,In_197);
nor U607 (N_607,In_52,In_333);
nand U608 (N_608,In_388,In_602);
or U609 (N_609,In_711,In_366);
nor U610 (N_610,In_74,In_87);
or U611 (N_611,In_430,In_405);
and U612 (N_612,In_747,In_607);
nand U613 (N_613,In_58,In_288);
nor U614 (N_614,In_238,In_260);
nor U615 (N_615,In_214,In_377);
xnor U616 (N_616,In_370,In_186);
nand U617 (N_617,In_714,In_492);
xor U618 (N_618,In_477,In_412);
nand U619 (N_619,In_135,In_636);
xor U620 (N_620,In_498,In_319);
nand U621 (N_621,In_43,In_50);
xor U622 (N_622,In_336,In_525);
nor U623 (N_623,In_482,In_246);
nor U624 (N_624,In_402,In_563);
xnor U625 (N_625,In_177,In_136);
or U626 (N_626,In_48,In_517);
nor U627 (N_627,In_653,In_705);
xnor U628 (N_628,In_637,In_453);
xnor U629 (N_629,In_708,In_606);
xnor U630 (N_630,In_671,In_295);
nand U631 (N_631,In_37,In_537);
and U632 (N_632,In_132,In_16);
nand U633 (N_633,In_555,In_120);
or U634 (N_634,In_746,In_21);
and U635 (N_635,In_629,In_56);
and U636 (N_636,In_19,In_300);
nor U637 (N_637,In_217,In_392);
nor U638 (N_638,In_538,In_256);
nor U639 (N_639,In_684,In_668);
or U640 (N_640,In_146,In_55);
nor U641 (N_641,In_477,In_717);
nand U642 (N_642,In_547,In_332);
and U643 (N_643,In_355,In_322);
nand U644 (N_644,In_77,In_325);
or U645 (N_645,In_253,In_354);
xnor U646 (N_646,In_211,In_288);
or U647 (N_647,In_226,In_257);
nand U648 (N_648,In_168,In_720);
xnor U649 (N_649,In_184,In_465);
nand U650 (N_650,In_174,In_319);
nand U651 (N_651,In_511,In_68);
xor U652 (N_652,In_739,In_160);
nand U653 (N_653,In_623,In_241);
xnor U654 (N_654,In_501,In_319);
xnor U655 (N_655,In_191,In_114);
or U656 (N_656,In_523,In_392);
nand U657 (N_657,In_123,In_327);
and U658 (N_658,In_252,In_147);
nand U659 (N_659,In_395,In_94);
xnor U660 (N_660,In_131,In_382);
nor U661 (N_661,In_83,In_227);
nand U662 (N_662,In_140,In_544);
nor U663 (N_663,In_534,In_75);
xor U664 (N_664,In_438,In_330);
and U665 (N_665,In_156,In_607);
or U666 (N_666,In_379,In_12);
xnor U667 (N_667,In_626,In_256);
or U668 (N_668,In_434,In_222);
nand U669 (N_669,In_561,In_515);
xnor U670 (N_670,In_34,In_666);
nand U671 (N_671,In_572,In_503);
and U672 (N_672,In_533,In_138);
and U673 (N_673,In_61,In_23);
and U674 (N_674,In_343,In_712);
xnor U675 (N_675,In_366,In_566);
and U676 (N_676,In_697,In_596);
xor U677 (N_677,In_150,In_296);
nand U678 (N_678,In_631,In_330);
xnor U679 (N_679,In_660,In_141);
xnor U680 (N_680,In_565,In_581);
or U681 (N_681,In_87,In_4);
nand U682 (N_682,In_321,In_587);
or U683 (N_683,In_629,In_378);
and U684 (N_684,In_247,In_545);
nor U685 (N_685,In_342,In_57);
xor U686 (N_686,In_69,In_241);
and U687 (N_687,In_71,In_243);
or U688 (N_688,In_241,In_402);
nand U689 (N_689,In_47,In_240);
nor U690 (N_690,In_284,In_730);
nand U691 (N_691,In_59,In_376);
nor U692 (N_692,In_504,In_585);
xor U693 (N_693,In_152,In_340);
nand U694 (N_694,In_491,In_236);
nor U695 (N_695,In_518,In_231);
nor U696 (N_696,In_378,In_208);
nand U697 (N_697,In_302,In_303);
or U698 (N_698,In_596,In_403);
xnor U699 (N_699,In_271,In_714);
or U700 (N_700,In_155,In_34);
xor U701 (N_701,In_242,In_22);
nor U702 (N_702,In_694,In_232);
and U703 (N_703,In_441,In_411);
and U704 (N_704,In_144,In_453);
nand U705 (N_705,In_403,In_536);
or U706 (N_706,In_471,In_399);
or U707 (N_707,In_88,In_282);
or U708 (N_708,In_357,In_23);
nor U709 (N_709,In_237,In_694);
nor U710 (N_710,In_434,In_408);
or U711 (N_711,In_603,In_446);
xor U712 (N_712,In_461,In_447);
or U713 (N_713,In_146,In_28);
and U714 (N_714,In_609,In_224);
and U715 (N_715,In_166,In_158);
and U716 (N_716,In_78,In_247);
nor U717 (N_717,In_295,In_31);
nor U718 (N_718,In_721,In_205);
and U719 (N_719,In_53,In_600);
xnor U720 (N_720,In_46,In_720);
or U721 (N_721,In_525,In_372);
xor U722 (N_722,In_301,In_9);
xnor U723 (N_723,In_319,In_106);
or U724 (N_724,In_459,In_609);
or U725 (N_725,In_599,In_186);
or U726 (N_726,In_457,In_479);
or U727 (N_727,In_2,In_581);
xor U728 (N_728,In_354,In_192);
nand U729 (N_729,In_316,In_517);
or U730 (N_730,In_720,In_684);
or U731 (N_731,In_402,In_711);
nor U732 (N_732,In_71,In_497);
and U733 (N_733,In_712,In_490);
xnor U734 (N_734,In_120,In_669);
xor U735 (N_735,In_201,In_496);
and U736 (N_736,In_184,In_717);
nor U737 (N_737,In_426,In_347);
nand U738 (N_738,In_528,In_288);
nand U739 (N_739,In_310,In_442);
xor U740 (N_740,In_640,In_388);
xnor U741 (N_741,In_110,In_458);
or U742 (N_742,In_517,In_585);
or U743 (N_743,In_366,In_243);
and U744 (N_744,In_734,In_103);
or U745 (N_745,In_275,In_124);
xnor U746 (N_746,In_543,In_599);
or U747 (N_747,In_339,In_637);
xnor U748 (N_748,In_353,In_480);
or U749 (N_749,In_424,In_500);
xnor U750 (N_750,In_121,In_520);
or U751 (N_751,In_564,In_142);
nor U752 (N_752,In_728,In_590);
xnor U753 (N_753,In_694,In_712);
xor U754 (N_754,In_292,In_308);
xor U755 (N_755,In_47,In_547);
nand U756 (N_756,In_65,In_449);
xnor U757 (N_757,In_653,In_386);
and U758 (N_758,In_436,In_586);
xnor U759 (N_759,In_98,In_421);
xnor U760 (N_760,In_80,In_266);
nand U761 (N_761,In_156,In_340);
nor U762 (N_762,In_723,In_265);
nor U763 (N_763,In_292,In_184);
xnor U764 (N_764,In_580,In_296);
or U765 (N_765,In_464,In_506);
xor U766 (N_766,In_221,In_249);
xor U767 (N_767,In_109,In_419);
xor U768 (N_768,In_307,In_321);
nand U769 (N_769,In_250,In_597);
and U770 (N_770,In_666,In_212);
and U771 (N_771,In_26,In_681);
and U772 (N_772,In_129,In_121);
nand U773 (N_773,In_19,In_172);
nor U774 (N_774,In_221,In_180);
and U775 (N_775,In_62,In_155);
nor U776 (N_776,In_391,In_466);
or U777 (N_777,In_21,In_540);
nand U778 (N_778,In_46,In_296);
nand U779 (N_779,In_721,In_631);
nand U780 (N_780,In_30,In_117);
xor U781 (N_781,In_567,In_632);
nand U782 (N_782,In_65,In_589);
nor U783 (N_783,In_588,In_543);
nor U784 (N_784,In_351,In_484);
nor U785 (N_785,In_196,In_383);
and U786 (N_786,In_512,In_525);
xor U787 (N_787,In_215,In_748);
and U788 (N_788,In_688,In_651);
or U789 (N_789,In_351,In_517);
and U790 (N_790,In_346,In_583);
and U791 (N_791,In_709,In_73);
and U792 (N_792,In_331,In_173);
xnor U793 (N_793,In_351,In_680);
nor U794 (N_794,In_232,In_508);
xnor U795 (N_795,In_1,In_19);
nand U796 (N_796,In_731,In_322);
or U797 (N_797,In_168,In_626);
or U798 (N_798,In_568,In_60);
nor U799 (N_799,In_602,In_59);
and U800 (N_800,In_161,In_123);
nor U801 (N_801,In_194,In_624);
xor U802 (N_802,In_601,In_709);
and U803 (N_803,In_61,In_204);
nand U804 (N_804,In_135,In_472);
nor U805 (N_805,In_75,In_10);
xor U806 (N_806,In_649,In_439);
and U807 (N_807,In_369,In_650);
xor U808 (N_808,In_376,In_164);
nand U809 (N_809,In_646,In_37);
and U810 (N_810,In_677,In_540);
xnor U811 (N_811,In_334,In_307);
and U812 (N_812,In_39,In_534);
or U813 (N_813,In_134,In_120);
nand U814 (N_814,In_443,In_142);
nor U815 (N_815,In_314,In_337);
nand U816 (N_816,In_656,In_36);
nand U817 (N_817,In_48,In_449);
and U818 (N_818,In_441,In_747);
and U819 (N_819,In_97,In_363);
xnor U820 (N_820,In_455,In_218);
nor U821 (N_821,In_123,In_580);
nand U822 (N_822,In_188,In_206);
xnor U823 (N_823,In_694,In_386);
and U824 (N_824,In_472,In_171);
or U825 (N_825,In_10,In_725);
and U826 (N_826,In_481,In_590);
or U827 (N_827,In_307,In_441);
and U828 (N_828,In_528,In_227);
nand U829 (N_829,In_321,In_632);
nand U830 (N_830,In_445,In_737);
nand U831 (N_831,In_394,In_195);
nor U832 (N_832,In_675,In_140);
and U833 (N_833,In_482,In_80);
nor U834 (N_834,In_567,In_519);
nor U835 (N_835,In_116,In_366);
or U836 (N_836,In_365,In_132);
nand U837 (N_837,In_300,In_682);
nand U838 (N_838,In_634,In_371);
and U839 (N_839,In_480,In_432);
or U840 (N_840,In_701,In_473);
and U841 (N_841,In_185,In_37);
nand U842 (N_842,In_544,In_275);
and U843 (N_843,In_231,In_20);
and U844 (N_844,In_285,In_526);
xor U845 (N_845,In_569,In_743);
or U846 (N_846,In_308,In_22);
nor U847 (N_847,In_294,In_3);
nand U848 (N_848,In_570,In_598);
nor U849 (N_849,In_13,In_366);
or U850 (N_850,In_584,In_362);
xnor U851 (N_851,In_197,In_210);
nor U852 (N_852,In_378,In_84);
nand U853 (N_853,In_171,In_179);
or U854 (N_854,In_42,In_144);
nor U855 (N_855,In_233,In_18);
or U856 (N_856,In_265,In_406);
nand U857 (N_857,In_595,In_385);
or U858 (N_858,In_684,In_395);
xnor U859 (N_859,In_2,In_425);
nor U860 (N_860,In_630,In_309);
nand U861 (N_861,In_573,In_635);
nor U862 (N_862,In_192,In_73);
xor U863 (N_863,In_5,In_144);
xnor U864 (N_864,In_588,In_600);
nor U865 (N_865,In_143,In_687);
xnor U866 (N_866,In_314,In_128);
or U867 (N_867,In_88,In_381);
nor U868 (N_868,In_480,In_239);
or U869 (N_869,In_516,In_634);
or U870 (N_870,In_186,In_707);
nand U871 (N_871,In_381,In_182);
nor U872 (N_872,In_318,In_251);
xor U873 (N_873,In_572,In_681);
or U874 (N_874,In_226,In_512);
and U875 (N_875,In_214,In_363);
nor U876 (N_876,In_539,In_706);
nand U877 (N_877,In_80,In_232);
nor U878 (N_878,In_350,In_50);
or U879 (N_879,In_693,In_362);
nand U880 (N_880,In_415,In_42);
xnor U881 (N_881,In_713,In_201);
nor U882 (N_882,In_218,In_251);
xnor U883 (N_883,In_668,In_266);
nand U884 (N_884,In_171,In_256);
nor U885 (N_885,In_56,In_258);
and U886 (N_886,In_331,In_82);
or U887 (N_887,In_496,In_550);
or U888 (N_888,In_502,In_446);
xor U889 (N_889,In_56,In_472);
or U890 (N_890,In_334,In_82);
or U891 (N_891,In_268,In_718);
xnor U892 (N_892,In_603,In_249);
nand U893 (N_893,In_565,In_244);
nand U894 (N_894,In_652,In_369);
or U895 (N_895,In_423,In_46);
xor U896 (N_896,In_723,In_134);
nand U897 (N_897,In_366,In_143);
or U898 (N_898,In_76,In_87);
and U899 (N_899,In_589,In_571);
or U900 (N_900,In_473,In_298);
nand U901 (N_901,In_135,In_222);
or U902 (N_902,In_249,In_98);
or U903 (N_903,In_255,In_686);
nand U904 (N_904,In_41,In_588);
xnor U905 (N_905,In_455,In_461);
or U906 (N_906,In_111,In_504);
and U907 (N_907,In_303,In_155);
nor U908 (N_908,In_161,In_373);
or U909 (N_909,In_633,In_744);
or U910 (N_910,In_411,In_703);
nor U911 (N_911,In_437,In_206);
or U912 (N_912,In_417,In_320);
or U913 (N_913,In_77,In_322);
and U914 (N_914,In_320,In_576);
and U915 (N_915,In_10,In_286);
nand U916 (N_916,In_128,In_511);
or U917 (N_917,In_238,In_193);
and U918 (N_918,In_609,In_417);
nor U919 (N_919,In_268,In_354);
nor U920 (N_920,In_386,In_377);
or U921 (N_921,In_585,In_70);
xor U922 (N_922,In_214,In_551);
and U923 (N_923,In_215,In_389);
xor U924 (N_924,In_566,In_585);
xnor U925 (N_925,In_416,In_450);
nor U926 (N_926,In_275,In_92);
nand U927 (N_927,In_202,In_123);
or U928 (N_928,In_466,In_706);
nor U929 (N_929,In_691,In_177);
and U930 (N_930,In_399,In_195);
nand U931 (N_931,In_331,In_40);
xor U932 (N_932,In_67,In_317);
nor U933 (N_933,In_391,In_414);
nand U934 (N_934,In_132,In_560);
nor U935 (N_935,In_18,In_172);
or U936 (N_936,In_334,In_444);
or U937 (N_937,In_440,In_639);
nand U938 (N_938,In_659,In_106);
nor U939 (N_939,In_538,In_635);
nand U940 (N_940,In_112,In_57);
nor U941 (N_941,In_670,In_599);
nor U942 (N_942,In_65,In_613);
or U943 (N_943,In_355,In_483);
xnor U944 (N_944,In_84,In_551);
nand U945 (N_945,In_518,In_192);
xnor U946 (N_946,In_163,In_634);
nor U947 (N_947,In_459,In_435);
or U948 (N_948,In_180,In_502);
xnor U949 (N_949,In_548,In_169);
xnor U950 (N_950,In_651,In_466);
nor U951 (N_951,In_545,In_400);
and U952 (N_952,In_273,In_616);
nor U953 (N_953,In_32,In_609);
or U954 (N_954,In_472,In_406);
and U955 (N_955,In_116,In_125);
xnor U956 (N_956,In_249,In_639);
xnor U957 (N_957,In_498,In_712);
nand U958 (N_958,In_156,In_747);
nor U959 (N_959,In_98,In_50);
xnor U960 (N_960,In_571,In_131);
and U961 (N_961,In_46,In_654);
nor U962 (N_962,In_512,In_319);
nor U963 (N_963,In_710,In_726);
xnor U964 (N_964,In_334,In_592);
nor U965 (N_965,In_43,In_448);
nor U966 (N_966,In_150,In_326);
or U967 (N_967,In_32,In_622);
nor U968 (N_968,In_127,In_565);
nand U969 (N_969,In_436,In_615);
nand U970 (N_970,In_465,In_266);
or U971 (N_971,In_429,In_255);
nor U972 (N_972,In_723,In_6);
or U973 (N_973,In_353,In_291);
or U974 (N_974,In_76,In_133);
nand U975 (N_975,In_415,In_673);
xor U976 (N_976,In_479,In_53);
xnor U977 (N_977,In_348,In_359);
or U978 (N_978,In_710,In_251);
xnor U979 (N_979,In_690,In_618);
nor U980 (N_980,In_26,In_361);
and U981 (N_981,In_520,In_1);
nor U982 (N_982,In_335,In_566);
nand U983 (N_983,In_173,In_409);
or U984 (N_984,In_695,In_620);
nor U985 (N_985,In_717,In_106);
nand U986 (N_986,In_135,In_28);
nand U987 (N_987,In_295,In_577);
or U988 (N_988,In_50,In_49);
xor U989 (N_989,In_563,In_166);
nor U990 (N_990,In_142,In_72);
or U991 (N_991,In_141,In_726);
and U992 (N_992,In_687,In_314);
and U993 (N_993,In_130,In_229);
xor U994 (N_994,In_408,In_141);
or U995 (N_995,In_187,In_269);
or U996 (N_996,In_255,In_379);
nand U997 (N_997,In_583,In_547);
or U998 (N_998,In_57,In_246);
nor U999 (N_999,In_337,In_244);
xor U1000 (N_1000,N_118,N_610);
and U1001 (N_1001,N_218,N_614);
nand U1002 (N_1002,N_102,N_660);
nor U1003 (N_1003,N_127,N_580);
and U1004 (N_1004,N_898,N_282);
nor U1005 (N_1005,N_55,N_223);
xor U1006 (N_1006,N_843,N_917);
xor U1007 (N_1007,N_592,N_452);
nor U1008 (N_1008,N_44,N_585);
and U1009 (N_1009,N_725,N_745);
nand U1010 (N_1010,N_908,N_24);
nand U1011 (N_1011,N_357,N_685);
xnor U1012 (N_1012,N_20,N_695);
and U1013 (N_1013,N_265,N_663);
nor U1014 (N_1014,N_617,N_151);
nor U1015 (N_1015,N_573,N_18);
nand U1016 (N_1016,N_906,N_674);
xnor U1017 (N_1017,N_266,N_719);
xnor U1018 (N_1018,N_647,N_801);
and U1019 (N_1019,N_973,N_176);
nor U1020 (N_1020,N_974,N_53);
and U1021 (N_1021,N_572,N_181);
nor U1022 (N_1022,N_857,N_528);
nand U1023 (N_1023,N_839,N_829);
nor U1024 (N_1024,N_943,N_816);
nand U1025 (N_1025,N_72,N_246);
nor U1026 (N_1026,N_915,N_778);
nor U1027 (N_1027,N_620,N_830);
and U1028 (N_1028,N_810,N_712);
and U1029 (N_1029,N_208,N_64);
nor U1030 (N_1030,N_85,N_893);
xor U1031 (N_1031,N_413,N_992);
or U1032 (N_1032,N_30,N_26);
or U1033 (N_1033,N_379,N_133);
nand U1034 (N_1034,N_588,N_329);
xnor U1035 (N_1035,N_502,N_467);
or U1036 (N_1036,N_365,N_213);
nor U1037 (N_1037,N_203,N_478);
nand U1038 (N_1038,N_336,N_288);
and U1039 (N_1039,N_22,N_99);
nor U1040 (N_1040,N_986,N_684);
xor U1041 (N_1041,N_602,N_408);
nand U1042 (N_1042,N_308,N_871);
nor U1043 (N_1043,N_404,N_277);
and U1044 (N_1044,N_979,N_319);
xor U1045 (N_1045,N_561,N_993);
xor U1046 (N_1046,N_146,N_971);
xnor U1047 (N_1047,N_394,N_383);
or U1048 (N_1048,N_390,N_96);
or U1049 (N_1049,N_761,N_527);
and U1050 (N_1050,N_862,N_946);
and U1051 (N_1051,N_501,N_3);
or U1052 (N_1052,N_791,N_814);
nor U1053 (N_1053,N_370,N_782);
or U1054 (N_1054,N_513,N_727);
xnor U1055 (N_1055,N_728,N_866);
and U1056 (N_1056,N_518,N_395);
and U1057 (N_1057,N_207,N_444);
nor U1058 (N_1058,N_587,N_454);
xor U1059 (N_1059,N_988,N_364);
nor U1060 (N_1060,N_362,N_556);
nor U1061 (N_1061,N_476,N_98);
and U1062 (N_1062,N_8,N_382);
or U1063 (N_1063,N_461,N_380);
xor U1064 (N_1064,N_419,N_922);
or U1065 (N_1065,N_978,N_516);
or U1066 (N_1066,N_576,N_432);
or U1067 (N_1067,N_892,N_4);
or U1068 (N_1068,N_239,N_604);
or U1069 (N_1069,N_568,N_81);
nand U1070 (N_1070,N_631,N_51);
and U1071 (N_1071,N_124,N_799);
xor U1072 (N_1072,N_780,N_594);
or U1073 (N_1073,N_564,N_86);
and U1074 (N_1074,N_31,N_255);
xor U1075 (N_1075,N_312,N_437);
nand U1076 (N_1076,N_253,N_537);
nand U1077 (N_1077,N_515,N_637);
nand U1078 (N_1078,N_804,N_338);
xor U1079 (N_1079,N_733,N_903);
or U1080 (N_1080,N_640,N_865);
xor U1081 (N_1081,N_271,N_701);
and U1082 (N_1082,N_784,N_540);
nor U1083 (N_1083,N_194,N_872);
and U1084 (N_1084,N_536,N_738);
or U1085 (N_1085,N_835,N_403);
nor U1086 (N_1086,N_916,N_658);
and U1087 (N_1087,N_422,N_205);
nor U1088 (N_1088,N_311,N_760);
nor U1089 (N_1089,N_555,N_14);
nor U1090 (N_1090,N_32,N_430);
nor U1091 (N_1091,N_7,N_578);
or U1092 (N_1092,N_339,N_655);
xor U1093 (N_1093,N_41,N_486);
xnor U1094 (N_1094,N_928,N_877);
nand U1095 (N_1095,N_995,N_68);
and U1096 (N_1096,N_62,N_171);
or U1097 (N_1097,N_976,N_888);
nor U1098 (N_1098,N_508,N_850);
xor U1099 (N_1099,N_797,N_393);
xnor U1100 (N_1100,N_763,N_170);
and U1101 (N_1101,N_165,N_87);
nand U1102 (N_1102,N_268,N_899);
xnor U1103 (N_1103,N_115,N_284);
or U1104 (N_1104,N_441,N_927);
and U1105 (N_1105,N_608,N_938);
or U1106 (N_1106,N_914,N_37);
nor U1107 (N_1107,N_214,N_683);
xnor U1108 (N_1108,N_128,N_689);
nor U1109 (N_1109,N_818,N_129);
nand U1110 (N_1110,N_199,N_227);
nor U1111 (N_1111,N_896,N_547);
and U1112 (N_1112,N_652,N_356);
xor U1113 (N_1113,N_638,N_158);
xor U1114 (N_1114,N_786,N_964);
xnor U1115 (N_1115,N_942,N_249);
and U1116 (N_1116,N_889,N_581);
or U1117 (N_1117,N_632,N_273);
and U1118 (N_1118,N_653,N_27);
xnor U1119 (N_1119,N_807,N_226);
nor U1120 (N_1120,N_93,N_939);
xor U1121 (N_1121,N_177,N_112);
or U1122 (N_1122,N_316,N_79);
xnor U1123 (N_1123,N_793,N_700);
and U1124 (N_1124,N_464,N_425);
nor U1125 (N_1125,N_345,N_285);
and U1126 (N_1126,N_377,N_428);
xor U1127 (N_1127,N_317,N_178);
nand U1128 (N_1128,N_824,N_856);
xnor U1129 (N_1129,N_245,N_673);
or U1130 (N_1130,N_539,N_509);
or U1131 (N_1131,N_325,N_254);
nor U1132 (N_1132,N_813,N_426);
xor U1133 (N_1133,N_16,N_307);
xor U1134 (N_1134,N_56,N_634);
nor U1135 (N_1135,N_770,N_15);
xnor U1136 (N_1136,N_193,N_827);
or U1137 (N_1137,N_635,N_174);
xor U1138 (N_1138,N_867,N_676);
or U1139 (N_1139,N_766,N_78);
nand U1140 (N_1140,N_969,N_94);
and U1141 (N_1141,N_474,N_876);
nand U1142 (N_1142,N_551,N_812);
or U1143 (N_1143,N_233,N_263);
xnor U1144 (N_1144,N_142,N_76);
nand U1145 (N_1145,N_645,N_729);
xor U1146 (N_1146,N_229,N_546);
nand U1147 (N_1147,N_232,N_526);
and U1148 (N_1148,N_870,N_303);
and U1149 (N_1149,N_163,N_458);
or U1150 (N_1150,N_961,N_344);
and U1151 (N_1151,N_295,N_815);
nand U1152 (N_1152,N_584,N_720);
nand U1153 (N_1153,N_490,N_941);
nor U1154 (N_1154,N_929,N_145);
and U1155 (N_1155,N_967,N_292);
and U1156 (N_1156,N_672,N_741);
nor U1157 (N_1157,N_597,N_332);
or U1158 (N_1158,N_694,N_407);
nor U1159 (N_1159,N_999,N_260);
nand U1160 (N_1160,N_755,N_693);
nand U1161 (N_1161,N_438,N_542);
or U1162 (N_1162,N_429,N_500);
nand U1163 (N_1163,N_601,N_228);
xor U1164 (N_1164,N_730,N_443);
nor U1165 (N_1165,N_117,N_711);
or U1166 (N_1166,N_140,N_465);
xor U1167 (N_1167,N_703,N_936);
nand U1168 (N_1168,N_753,N_483);
nand U1169 (N_1169,N_590,N_71);
or U1170 (N_1170,N_415,N_103);
nor U1171 (N_1171,N_744,N_38);
xor U1172 (N_1172,N_952,N_781);
and U1173 (N_1173,N_657,N_854);
nand U1174 (N_1174,N_708,N_34);
or U1175 (N_1175,N_912,N_543);
or U1176 (N_1176,N_368,N_958);
nand U1177 (N_1177,N_525,N_777);
nor U1178 (N_1178,N_678,N_805);
nor U1179 (N_1179,N_299,N_350);
nor U1180 (N_1180,N_475,N_863);
nand U1181 (N_1181,N_479,N_636);
nor U1182 (N_1182,N_180,N_963);
xnor U1183 (N_1183,N_553,N_251);
or U1184 (N_1184,N_541,N_667);
xnor U1185 (N_1185,N_433,N_977);
or U1186 (N_1186,N_951,N_82);
xor U1187 (N_1187,N_398,N_788);
and U1188 (N_1188,N_164,N_692);
or U1189 (N_1189,N_983,N_1);
and U1190 (N_1190,N_73,N_715);
nor U1191 (N_1191,N_837,N_574);
or U1192 (N_1192,N_794,N_758);
and U1193 (N_1193,N_722,N_982);
xnor U1194 (N_1194,N_264,N_363);
nand U1195 (N_1195,N_449,N_405);
or U1196 (N_1196,N_58,N_886);
and U1197 (N_1197,N_742,N_931);
or U1198 (N_1198,N_846,N_157);
or U1199 (N_1199,N_358,N_477);
nand U1200 (N_1200,N_234,N_460);
and U1201 (N_1201,N_890,N_447);
nand U1202 (N_1202,N_654,N_902);
and U1203 (N_1203,N_644,N_291);
or U1204 (N_1204,N_323,N_834);
nor U1205 (N_1205,N_346,N_217);
or U1206 (N_1206,N_534,N_947);
xor U1207 (N_1207,N_281,N_114);
nor U1208 (N_1208,N_523,N_153);
and U1209 (N_1209,N_107,N_101);
nor U1210 (N_1210,N_399,N_354);
or U1211 (N_1211,N_57,N_385);
or U1212 (N_1212,N_119,N_949);
and U1213 (N_1213,N_396,N_498);
or U1214 (N_1214,N_446,N_397);
nor U1215 (N_1215,N_792,N_192);
nand U1216 (N_1216,N_195,N_175);
nand U1217 (N_1217,N_29,N_11);
nor U1218 (N_1218,N_67,N_686);
nand U1219 (N_1219,N_125,N_707);
and U1220 (N_1220,N_661,N_326);
nor U1221 (N_1221,N_371,N_409);
nand U1222 (N_1222,N_940,N_548);
nand U1223 (N_1223,N_185,N_734);
and U1224 (N_1224,N_267,N_488);
or U1225 (N_1225,N_283,N_337);
xor U1226 (N_1226,N_416,N_340);
nor U1227 (N_1227,N_562,N_844);
nand U1228 (N_1228,N_216,N_533);
nor U1229 (N_1229,N_910,N_819);
and U1230 (N_1230,N_154,N_343);
nand U1231 (N_1231,N_648,N_159);
nand U1232 (N_1232,N_802,N_66);
nand U1233 (N_1233,N_414,N_297);
or U1234 (N_1234,N_45,N_321);
and U1235 (N_1235,N_705,N_296);
xor U1236 (N_1236,N_959,N_275);
nor U1237 (N_1237,N_932,N_49);
xnor U1238 (N_1238,N_47,N_361);
nor U1239 (N_1239,N_987,N_531);
or U1240 (N_1240,N_769,N_933);
nor U1241 (N_1241,N_417,N_197);
nor U1242 (N_1242,N_909,N_565);
nand U1243 (N_1243,N_463,N_421);
and U1244 (N_1244,N_450,N_52);
nor U1245 (N_1245,N_111,N_400);
and U1246 (N_1246,N_298,N_209);
xnor U1247 (N_1247,N_764,N_605);
xnor U1248 (N_1248,N_504,N_897);
nor U1249 (N_1249,N_981,N_148);
xnor U1250 (N_1250,N_420,N_322);
nor U1251 (N_1251,N_747,N_726);
or U1252 (N_1252,N_554,N_716);
xor U1253 (N_1253,N_833,N_823);
and U1254 (N_1254,N_828,N_168);
nor U1255 (N_1255,N_762,N_704);
nor U1256 (N_1256,N_43,N_318);
and U1257 (N_1257,N_519,N_732);
nand U1258 (N_1258,N_682,N_427);
nand U1259 (N_1259,N_348,N_497);
and U1260 (N_1260,N_334,N_161);
or U1261 (N_1261,N_373,N_962);
or U1262 (N_1262,N_424,N_46);
and U1263 (N_1263,N_878,N_10);
xnor U1264 (N_1264,N_293,N_538);
nand U1265 (N_1265,N_595,N_996);
xor U1266 (N_1266,N_873,N_706);
xnor U1267 (N_1267,N_775,N_110);
nor U1268 (N_1268,N_520,N_184);
xor U1269 (N_1269,N_615,N_126);
or U1270 (N_1270,N_545,N_607);
nor U1271 (N_1271,N_493,N_972);
xor U1272 (N_1272,N_25,N_410);
nand U1273 (N_1273,N_290,N_681);
nor U1274 (N_1274,N_659,N_261);
xor U1275 (N_1275,N_859,N_328);
xor U1276 (N_1276,N_800,N_221);
nand U1277 (N_1277,N_852,N_558);
xnor U1278 (N_1278,N_975,N_524);
and U1279 (N_1279,N_5,N_529);
nor U1280 (N_1280,N_690,N_492);
nor U1281 (N_1281,N_309,N_120);
nor U1282 (N_1282,N_42,N_924);
xnor U1283 (N_1283,N_522,N_579);
nand U1284 (N_1284,N_306,N_74);
or U1285 (N_1285,N_984,N_147);
xnor U1286 (N_1286,N_629,N_649);
nand U1287 (N_1287,N_6,N_905);
xor U1288 (N_1288,N_847,N_990);
and U1289 (N_1289,N_259,N_998);
and U1290 (N_1290,N_262,N_521);
nor U1291 (N_1291,N_935,N_869);
nand U1292 (N_1292,N_108,N_855);
nor U1293 (N_1293,N_470,N_287);
and U1294 (N_1294,N_469,N_589);
xnor U1295 (N_1295,N_70,N_968);
nand U1296 (N_1296,N_826,N_269);
xnor U1297 (N_1297,N_480,N_880);
xnor U1298 (N_1298,N_149,N_434);
or U1299 (N_1299,N_330,N_225);
nor U1300 (N_1300,N_305,N_367);
nand U1301 (N_1301,N_646,N_445);
and U1302 (N_1302,N_808,N_603);
or U1303 (N_1303,N_774,N_59);
or U1304 (N_1304,N_628,N_511);
and U1305 (N_1305,N_13,N_392);
nand U1306 (N_1306,N_820,N_625);
nor U1307 (N_1307,N_756,N_335);
xnor U1308 (N_1308,N_378,N_560);
xnor U1309 (N_1309,N_662,N_131);
nor U1310 (N_1310,N_771,N_435);
or U1311 (N_1311,N_289,N_593);
and U1312 (N_1312,N_459,N_768);
and U1313 (N_1313,N_384,N_506);
and U1314 (N_1314,N_359,N_577);
nand U1315 (N_1315,N_806,N_247);
or U1316 (N_1316,N_202,N_466);
xnor U1317 (N_1317,N_624,N_136);
and U1318 (N_1318,N_853,N_630);
nand U1319 (N_1319,N_122,N_173);
nand U1320 (N_1320,N_215,N_187);
or U1321 (N_1321,N_135,N_50);
xnor U1322 (N_1322,N_116,N_945);
and U1323 (N_1323,N_505,N_842);
or U1324 (N_1324,N_256,N_104);
or U1325 (N_1325,N_822,N_473);
and U1326 (N_1326,N_402,N_456);
nand U1327 (N_1327,N_63,N_535);
or U1328 (N_1328,N_751,N_95);
or U1329 (N_1329,N_439,N_132);
and U1330 (N_1330,N_36,N_713);
and U1331 (N_1331,N_406,N_582);
xnor U1332 (N_1332,N_864,N_746);
nor U1333 (N_1333,N_575,N_765);
xor U1334 (N_1334,N_622,N_65);
xor U1335 (N_1335,N_918,N_201);
xnor U1336 (N_1336,N_489,N_472);
nor U1337 (N_1337,N_33,N_436);
nor U1338 (N_1338,N_210,N_200);
nor U1339 (N_1339,N_586,N_376);
nor U1340 (N_1340,N_731,N_710);
or U1341 (N_1341,N_567,N_381);
nand U1342 (N_1342,N_374,N_883);
nand U1343 (N_1343,N_491,N_28);
and U1344 (N_1344,N_9,N_301);
xor U1345 (N_1345,N_613,N_569);
and U1346 (N_1346,N_858,N_276);
nand U1347 (N_1347,N_391,N_736);
or U1348 (N_1348,N_349,N_485);
nand U1349 (N_1349,N_144,N_162);
nand U1350 (N_1350,N_724,N_671);
nor U1351 (N_1351,N_907,N_327);
xor U1352 (N_1352,N_570,N_167);
xnor U1353 (N_1353,N_809,N_698);
or U1354 (N_1354,N_484,N_143);
nor U1355 (N_1355,N_514,N_887);
nand U1356 (N_1356,N_235,N_219);
or U1357 (N_1357,N_457,N_411);
nor U1358 (N_1358,N_583,N_294);
nand U1359 (N_1359,N_669,N_507);
nor U1360 (N_1360,N_709,N_596);
nand U1361 (N_1361,N_286,N_956);
xor U1362 (N_1362,N_718,N_641);
nor U1363 (N_1363,N_137,N_369);
xnor U1364 (N_1364,N_244,N_313);
and U1365 (N_1365,N_189,N_776);
and U1366 (N_1366,N_848,N_832);
nor U1367 (N_1367,N_714,N_944);
or U1368 (N_1368,N_591,N_190);
and U1369 (N_1369,N_243,N_900);
xnor U1370 (N_1370,N_222,N_891);
xor U1371 (N_1371,N_304,N_191);
or U1372 (N_1372,N_677,N_186);
and U1373 (N_1373,N_453,N_544);
nor U1374 (N_1374,N_687,N_656);
nor U1375 (N_1375,N_650,N_759);
nor U1376 (N_1376,N_994,N_302);
xor U1377 (N_1377,N_894,N_90);
nor U1378 (N_1378,N_389,N_626);
nand U1379 (N_1379,N_623,N_743);
xnor U1380 (N_1380,N_23,N_599);
xnor U1381 (N_1381,N_183,N_113);
or U1382 (N_1382,N_803,N_904);
nand U1383 (N_1383,N_783,N_836);
and U1384 (N_1384,N_875,N_559);
nand U1385 (N_1385,N_767,N_600);
or U1386 (N_1386,N_851,N_451);
nand U1387 (N_1387,N_885,N_966);
nor U1388 (N_1388,N_423,N_923);
and U1389 (N_1389,N_749,N_75);
or U1390 (N_1390,N_487,N_83);
nor U1391 (N_1391,N_372,N_980);
nor U1392 (N_1392,N_238,N_412);
and U1393 (N_1393,N_258,N_611);
nand U1394 (N_1394,N_80,N_911);
and U1395 (N_1395,N_152,N_550);
and U1396 (N_1396,N_355,N_196);
nand U1397 (N_1397,N_735,N_665);
nand U1398 (N_1398,N_106,N_670);
and U1399 (N_1399,N_960,N_785);
xor U1400 (N_1400,N_401,N_532);
nand U1401 (N_1401,N_950,N_621);
nor U1402 (N_1402,N_757,N_787);
and U1403 (N_1403,N_206,N_39);
nor U1404 (N_1404,N_557,N_320);
and U1405 (N_1405,N_212,N_881);
and U1406 (N_1406,N_69,N_48);
and U1407 (N_1407,N_351,N_77);
and U1408 (N_1408,N_619,N_825);
nor U1409 (N_1409,N_552,N_643);
or U1410 (N_1410,N_274,N_440);
xor U1411 (N_1411,N_699,N_0);
nand U1412 (N_1412,N_347,N_606);
and U1413 (N_1413,N_779,N_182);
nor U1414 (N_1414,N_954,N_879);
or U1415 (N_1415,N_211,N_737);
nor U1416 (N_1416,N_431,N_130);
xor U1417 (N_1417,N_324,N_2);
and U1418 (N_1418,N_895,N_821);
or U1419 (N_1419,N_868,N_495);
nand U1420 (N_1420,N_970,N_188);
nand U1421 (N_1421,N_353,N_861);
xnor U1422 (N_1422,N_811,N_97);
nand U1423 (N_1423,N_270,N_252);
xnor U1424 (N_1424,N_789,N_333);
xnor U1425 (N_1425,N_169,N_697);
and U1426 (N_1426,N_691,N_642);
nor U1427 (N_1427,N_985,N_499);
xnor U1428 (N_1428,N_138,N_198);
nor U1429 (N_1429,N_21,N_633);
nand U1430 (N_1430,N_503,N_530);
nand U1431 (N_1431,N_386,N_874);
and U1432 (N_1432,N_242,N_752);
or U1433 (N_1433,N_717,N_748);
nor U1434 (N_1434,N_310,N_612);
and U1435 (N_1435,N_919,N_240);
or U1436 (N_1436,N_230,N_627);
and U1437 (N_1437,N_224,N_937);
xnor U1438 (N_1438,N_989,N_123);
xnor U1439 (N_1439,N_618,N_639);
or U1440 (N_1440,N_12,N_315);
and U1441 (N_1441,N_442,N_237);
xnor U1442 (N_1442,N_278,N_664);
xor U1443 (N_1443,N_17,N_882);
nand U1444 (N_1444,N_675,N_61);
nand U1445 (N_1445,N_352,N_481);
nor U1446 (N_1446,N_668,N_166);
xor U1447 (N_1447,N_598,N_121);
and U1448 (N_1448,N_566,N_84);
or U1449 (N_1449,N_248,N_884);
xnor U1450 (N_1450,N_40,N_930);
or U1451 (N_1451,N_666,N_849);
or U1452 (N_1452,N_817,N_510);
xnor U1453 (N_1453,N_772,N_236);
xnor U1454 (N_1454,N_798,N_616);
xor U1455 (N_1455,N_341,N_455);
or U1456 (N_1456,N_279,N_272);
and U1457 (N_1457,N_257,N_549);
nand U1458 (N_1458,N_19,N_141);
and U1459 (N_1459,N_680,N_957);
or U1460 (N_1460,N_723,N_721);
nor U1461 (N_1461,N_241,N_841);
or U1462 (N_1462,N_92,N_54);
xor U1463 (N_1463,N_925,N_300);
or U1464 (N_1464,N_179,N_139);
nand U1465 (N_1465,N_342,N_831);
nor U1466 (N_1466,N_60,N_991);
and U1467 (N_1467,N_468,N_679);
nor U1468 (N_1468,N_156,N_388);
xnor U1469 (N_1469,N_471,N_934);
xnor U1470 (N_1470,N_462,N_109);
or U1471 (N_1471,N_840,N_696);
nand U1472 (N_1472,N_860,N_997);
nand U1473 (N_1473,N_496,N_688);
or U1474 (N_1474,N_160,N_91);
xor U1475 (N_1475,N_89,N_651);
and U1476 (N_1476,N_387,N_920);
nor U1477 (N_1477,N_754,N_773);
xnor U1478 (N_1478,N_795,N_375);
nor U1479 (N_1479,N_134,N_204);
nor U1480 (N_1480,N_845,N_482);
nand U1481 (N_1481,N_512,N_702);
nand U1482 (N_1482,N_448,N_948);
nand U1483 (N_1483,N_901,N_926);
nor U1484 (N_1484,N_35,N_517);
nor U1485 (N_1485,N_494,N_913);
and U1486 (N_1486,N_155,N_740);
nor U1487 (N_1487,N_921,N_750);
and U1488 (N_1488,N_366,N_150);
or U1489 (N_1489,N_360,N_965);
nand U1490 (N_1490,N_280,N_955);
and U1491 (N_1491,N_838,N_331);
or U1492 (N_1492,N_100,N_105);
or U1493 (N_1493,N_563,N_88);
xor U1494 (N_1494,N_220,N_418);
and U1495 (N_1495,N_250,N_172);
or U1496 (N_1496,N_790,N_796);
nor U1497 (N_1497,N_314,N_739);
and U1498 (N_1498,N_571,N_953);
nand U1499 (N_1499,N_231,N_609);
or U1500 (N_1500,N_753,N_969);
and U1501 (N_1501,N_795,N_565);
nand U1502 (N_1502,N_563,N_778);
and U1503 (N_1503,N_853,N_394);
nor U1504 (N_1504,N_37,N_166);
nand U1505 (N_1505,N_755,N_119);
nor U1506 (N_1506,N_966,N_768);
xnor U1507 (N_1507,N_740,N_618);
nand U1508 (N_1508,N_586,N_653);
xnor U1509 (N_1509,N_173,N_537);
or U1510 (N_1510,N_44,N_490);
or U1511 (N_1511,N_714,N_953);
nor U1512 (N_1512,N_192,N_518);
nand U1513 (N_1513,N_385,N_161);
or U1514 (N_1514,N_14,N_263);
xnor U1515 (N_1515,N_350,N_271);
nand U1516 (N_1516,N_601,N_467);
and U1517 (N_1517,N_580,N_234);
and U1518 (N_1518,N_47,N_22);
nand U1519 (N_1519,N_523,N_867);
or U1520 (N_1520,N_819,N_769);
or U1521 (N_1521,N_130,N_749);
nor U1522 (N_1522,N_234,N_253);
and U1523 (N_1523,N_665,N_620);
xor U1524 (N_1524,N_737,N_926);
xor U1525 (N_1525,N_692,N_382);
xnor U1526 (N_1526,N_224,N_659);
or U1527 (N_1527,N_580,N_106);
xor U1528 (N_1528,N_839,N_506);
xnor U1529 (N_1529,N_385,N_721);
nand U1530 (N_1530,N_543,N_740);
or U1531 (N_1531,N_521,N_936);
nor U1532 (N_1532,N_373,N_448);
nand U1533 (N_1533,N_736,N_967);
nor U1534 (N_1534,N_632,N_397);
nor U1535 (N_1535,N_92,N_953);
nor U1536 (N_1536,N_903,N_831);
nand U1537 (N_1537,N_805,N_88);
and U1538 (N_1538,N_597,N_635);
and U1539 (N_1539,N_731,N_576);
or U1540 (N_1540,N_463,N_729);
nor U1541 (N_1541,N_220,N_725);
nor U1542 (N_1542,N_506,N_195);
nor U1543 (N_1543,N_244,N_848);
or U1544 (N_1544,N_485,N_127);
nand U1545 (N_1545,N_873,N_629);
nor U1546 (N_1546,N_927,N_873);
nand U1547 (N_1547,N_241,N_412);
nor U1548 (N_1548,N_956,N_52);
nand U1549 (N_1549,N_671,N_932);
nand U1550 (N_1550,N_432,N_825);
xnor U1551 (N_1551,N_79,N_870);
and U1552 (N_1552,N_563,N_887);
xnor U1553 (N_1553,N_668,N_752);
xor U1554 (N_1554,N_726,N_92);
nor U1555 (N_1555,N_750,N_440);
and U1556 (N_1556,N_741,N_386);
nand U1557 (N_1557,N_715,N_912);
or U1558 (N_1558,N_324,N_350);
nor U1559 (N_1559,N_906,N_569);
xor U1560 (N_1560,N_33,N_933);
and U1561 (N_1561,N_476,N_623);
nor U1562 (N_1562,N_747,N_911);
nand U1563 (N_1563,N_223,N_280);
and U1564 (N_1564,N_17,N_274);
xnor U1565 (N_1565,N_813,N_2);
nor U1566 (N_1566,N_827,N_965);
nor U1567 (N_1567,N_167,N_528);
nor U1568 (N_1568,N_901,N_191);
nand U1569 (N_1569,N_629,N_743);
or U1570 (N_1570,N_440,N_455);
or U1571 (N_1571,N_533,N_697);
nor U1572 (N_1572,N_948,N_263);
or U1573 (N_1573,N_903,N_271);
xor U1574 (N_1574,N_544,N_751);
xnor U1575 (N_1575,N_717,N_538);
and U1576 (N_1576,N_707,N_835);
xnor U1577 (N_1577,N_459,N_33);
xnor U1578 (N_1578,N_497,N_188);
or U1579 (N_1579,N_702,N_350);
or U1580 (N_1580,N_972,N_800);
xnor U1581 (N_1581,N_315,N_73);
nand U1582 (N_1582,N_249,N_540);
nor U1583 (N_1583,N_331,N_307);
and U1584 (N_1584,N_343,N_900);
nand U1585 (N_1585,N_810,N_43);
and U1586 (N_1586,N_263,N_84);
nor U1587 (N_1587,N_366,N_400);
or U1588 (N_1588,N_347,N_319);
and U1589 (N_1589,N_590,N_52);
xnor U1590 (N_1590,N_112,N_975);
xor U1591 (N_1591,N_748,N_628);
xor U1592 (N_1592,N_773,N_913);
xnor U1593 (N_1593,N_748,N_55);
or U1594 (N_1594,N_295,N_663);
and U1595 (N_1595,N_962,N_312);
xor U1596 (N_1596,N_197,N_845);
nor U1597 (N_1597,N_936,N_433);
and U1598 (N_1598,N_245,N_584);
or U1599 (N_1599,N_174,N_807);
xnor U1600 (N_1600,N_597,N_47);
xor U1601 (N_1601,N_330,N_251);
nor U1602 (N_1602,N_728,N_413);
nor U1603 (N_1603,N_958,N_907);
xor U1604 (N_1604,N_302,N_589);
nor U1605 (N_1605,N_12,N_907);
xnor U1606 (N_1606,N_203,N_275);
or U1607 (N_1607,N_72,N_675);
nand U1608 (N_1608,N_932,N_888);
and U1609 (N_1609,N_921,N_205);
nor U1610 (N_1610,N_362,N_435);
xnor U1611 (N_1611,N_136,N_876);
and U1612 (N_1612,N_286,N_452);
xor U1613 (N_1613,N_739,N_802);
and U1614 (N_1614,N_840,N_471);
nor U1615 (N_1615,N_504,N_165);
or U1616 (N_1616,N_155,N_686);
and U1617 (N_1617,N_196,N_401);
xnor U1618 (N_1618,N_512,N_934);
xnor U1619 (N_1619,N_80,N_430);
nand U1620 (N_1620,N_89,N_307);
nor U1621 (N_1621,N_641,N_914);
nand U1622 (N_1622,N_997,N_237);
and U1623 (N_1623,N_918,N_956);
nor U1624 (N_1624,N_478,N_700);
xnor U1625 (N_1625,N_616,N_607);
nor U1626 (N_1626,N_392,N_366);
nor U1627 (N_1627,N_175,N_924);
nor U1628 (N_1628,N_12,N_807);
or U1629 (N_1629,N_703,N_415);
or U1630 (N_1630,N_4,N_253);
nor U1631 (N_1631,N_514,N_874);
nand U1632 (N_1632,N_215,N_747);
xnor U1633 (N_1633,N_876,N_824);
nor U1634 (N_1634,N_108,N_383);
and U1635 (N_1635,N_496,N_55);
and U1636 (N_1636,N_299,N_464);
xor U1637 (N_1637,N_364,N_866);
nand U1638 (N_1638,N_609,N_762);
xor U1639 (N_1639,N_356,N_184);
nor U1640 (N_1640,N_748,N_994);
and U1641 (N_1641,N_540,N_908);
and U1642 (N_1642,N_291,N_151);
nand U1643 (N_1643,N_49,N_89);
and U1644 (N_1644,N_801,N_968);
nor U1645 (N_1645,N_439,N_286);
nor U1646 (N_1646,N_979,N_284);
and U1647 (N_1647,N_269,N_536);
and U1648 (N_1648,N_533,N_263);
or U1649 (N_1649,N_404,N_11);
xor U1650 (N_1650,N_448,N_901);
xnor U1651 (N_1651,N_743,N_194);
nand U1652 (N_1652,N_997,N_454);
nor U1653 (N_1653,N_815,N_732);
nand U1654 (N_1654,N_227,N_622);
or U1655 (N_1655,N_554,N_420);
xnor U1656 (N_1656,N_378,N_832);
xor U1657 (N_1657,N_788,N_851);
and U1658 (N_1658,N_393,N_435);
or U1659 (N_1659,N_76,N_622);
and U1660 (N_1660,N_857,N_710);
nand U1661 (N_1661,N_897,N_808);
nor U1662 (N_1662,N_418,N_692);
nand U1663 (N_1663,N_266,N_843);
and U1664 (N_1664,N_582,N_910);
nor U1665 (N_1665,N_689,N_408);
nor U1666 (N_1666,N_898,N_460);
or U1667 (N_1667,N_695,N_963);
or U1668 (N_1668,N_160,N_261);
and U1669 (N_1669,N_260,N_423);
xnor U1670 (N_1670,N_879,N_117);
nor U1671 (N_1671,N_878,N_317);
or U1672 (N_1672,N_561,N_845);
nand U1673 (N_1673,N_391,N_828);
xor U1674 (N_1674,N_778,N_314);
nor U1675 (N_1675,N_138,N_521);
nand U1676 (N_1676,N_293,N_544);
xnor U1677 (N_1677,N_337,N_853);
and U1678 (N_1678,N_510,N_177);
or U1679 (N_1679,N_475,N_882);
nor U1680 (N_1680,N_884,N_701);
and U1681 (N_1681,N_558,N_983);
and U1682 (N_1682,N_654,N_446);
or U1683 (N_1683,N_842,N_402);
and U1684 (N_1684,N_262,N_861);
nand U1685 (N_1685,N_336,N_679);
nor U1686 (N_1686,N_611,N_679);
xnor U1687 (N_1687,N_517,N_7);
xnor U1688 (N_1688,N_926,N_860);
and U1689 (N_1689,N_730,N_839);
nand U1690 (N_1690,N_776,N_812);
xor U1691 (N_1691,N_14,N_205);
nor U1692 (N_1692,N_823,N_995);
or U1693 (N_1693,N_404,N_224);
or U1694 (N_1694,N_989,N_606);
xnor U1695 (N_1695,N_550,N_509);
nand U1696 (N_1696,N_507,N_603);
or U1697 (N_1697,N_374,N_284);
xor U1698 (N_1698,N_346,N_45);
nand U1699 (N_1699,N_787,N_3);
and U1700 (N_1700,N_239,N_561);
xor U1701 (N_1701,N_243,N_435);
xor U1702 (N_1702,N_62,N_511);
or U1703 (N_1703,N_864,N_872);
nor U1704 (N_1704,N_667,N_10);
nor U1705 (N_1705,N_972,N_931);
and U1706 (N_1706,N_832,N_901);
xnor U1707 (N_1707,N_153,N_103);
and U1708 (N_1708,N_109,N_562);
and U1709 (N_1709,N_566,N_41);
and U1710 (N_1710,N_708,N_924);
or U1711 (N_1711,N_492,N_120);
or U1712 (N_1712,N_734,N_340);
or U1713 (N_1713,N_880,N_73);
or U1714 (N_1714,N_394,N_95);
nor U1715 (N_1715,N_476,N_491);
nand U1716 (N_1716,N_128,N_449);
nand U1717 (N_1717,N_581,N_365);
nand U1718 (N_1718,N_426,N_769);
nor U1719 (N_1719,N_974,N_399);
or U1720 (N_1720,N_734,N_557);
nor U1721 (N_1721,N_539,N_828);
or U1722 (N_1722,N_880,N_64);
xor U1723 (N_1723,N_394,N_423);
xor U1724 (N_1724,N_999,N_409);
or U1725 (N_1725,N_356,N_444);
and U1726 (N_1726,N_928,N_452);
or U1727 (N_1727,N_9,N_874);
or U1728 (N_1728,N_610,N_386);
nor U1729 (N_1729,N_242,N_888);
nand U1730 (N_1730,N_918,N_457);
nand U1731 (N_1731,N_504,N_836);
or U1732 (N_1732,N_93,N_625);
or U1733 (N_1733,N_340,N_276);
or U1734 (N_1734,N_129,N_515);
or U1735 (N_1735,N_567,N_73);
nand U1736 (N_1736,N_546,N_803);
or U1737 (N_1737,N_956,N_701);
or U1738 (N_1738,N_454,N_936);
and U1739 (N_1739,N_715,N_401);
nand U1740 (N_1740,N_708,N_473);
nand U1741 (N_1741,N_72,N_232);
or U1742 (N_1742,N_32,N_68);
or U1743 (N_1743,N_60,N_162);
nand U1744 (N_1744,N_812,N_719);
nand U1745 (N_1745,N_644,N_804);
nand U1746 (N_1746,N_5,N_611);
and U1747 (N_1747,N_878,N_362);
nor U1748 (N_1748,N_978,N_340);
nand U1749 (N_1749,N_580,N_156);
or U1750 (N_1750,N_836,N_123);
and U1751 (N_1751,N_293,N_914);
and U1752 (N_1752,N_259,N_936);
or U1753 (N_1753,N_341,N_21);
nand U1754 (N_1754,N_48,N_335);
nand U1755 (N_1755,N_305,N_782);
nand U1756 (N_1756,N_345,N_399);
or U1757 (N_1757,N_506,N_783);
and U1758 (N_1758,N_624,N_42);
nand U1759 (N_1759,N_793,N_971);
nand U1760 (N_1760,N_133,N_110);
nor U1761 (N_1761,N_809,N_420);
nand U1762 (N_1762,N_947,N_567);
or U1763 (N_1763,N_421,N_966);
xor U1764 (N_1764,N_942,N_139);
and U1765 (N_1765,N_498,N_69);
or U1766 (N_1766,N_200,N_142);
nand U1767 (N_1767,N_579,N_955);
or U1768 (N_1768,N_172,N_395);
nand U1769 (N_1769,N_947,N_741);
nor U1770 (N_1770,N_80,N_401);
nor U1771 (N_1771,N_140,N_131);
nor U1772 (N_1772,N_906,N_137);
and U1773 (N_1773,N_935,N_809);
or U1774 (N_1774,N_371,N_769);
or U1775 (N_1775,N_301,N_423);
nor U1776 (N_1776,N_291,N_912);
or U1777 (N_1777,N_379,N_163);
and U1778 (N_1778,N_722,N_209);
xnor U1779 (N_1779,N_837,N_461);
or U1780 (N_1780,N_622,N_229);
nand U1781 (N_1781,N_80,N_165);
and U1782 (N_1782,N_106,N_934);
nand U1783 (N_1783,N_686,N_330);
or U1784 (N_1784,N_836,N_468);
nand U1785 (N_1785,N_372,N_423);
nand U1786 (N_1786,N_860,N_545);
nand U1787 (N_1787,N_339,N_539);
nand U1788 (N_1788,N_237,N_18);
nand U1789 (N_1789,N_863,N_623);
nand U1790 (N_1790,N_213,N_101);
or U1791 (N_1791,N_664,N_74);
nor U1792 (N_1792,N_936,N_782);
and U1793 (N_1793,N_761,N_995);
xnor U1794 (N_1794,N_503,N_534);
and U1795 (N_1795,N_424,N_237);
nor U1796 (N_1796,N_653,N_885);
and U1797 (N_1797,N_275,N_354);
nand U1798 (N_1798,N_948,N_904);
and U1799 (N_1799,N_213,N_382);
or U1800 (N_1800,N_478,N_818);
or U1801 (N_1801,N_711,N_157);
and U1802 (N_1802,N_649,N_979);
nand U1803 (N_1803,N_298,N_409);
and U1804 (N_1804,N_682,N_612);
or U1805 (N_1805,N_864,N_584);
nor U1806 (N_1806,N_302,N_598);
and U1807 (N_1807,N_444,N_935);
xor U1808 (N_1808,N_436,N_280);
and U1809 (N_1809,N_635,N_674);
nand U1810 (N_1810,N_256,N_334);
nor U1811 (N_1811,N_334,N_889);
or U1812 (N_1812,N_539,N_307);
xor U1813 (N_1813,N_336,N_493);
nor U1814 (N_1814,N_946,N_338);
nor U1815 (N_1815,N_101,N_443);
or U1816 (N_1816,N_920,N_125);
nor U1817 (N_1817,N_958,N_836);
nor U1818 (N_1818,N_584,N_556);
or U1819 (N_1819,N_144,N_207);
nand U1820 (N_1820,N_692,N_511);
nand U1821 (N_1821,N_641,N_453);
or U1822 (N_1822,N_44,N_900);
nand U1823 (N_1823,N_721,N_991);
or U1824 (N_1824,N_6,N_612);
or U1825 (N_1825,N_827,N_660);
nor U1826 (N_1826,N_7,N_389);
nor U1827 (N_1827,N_285,N_237);
nor U1828 (N_1828,N_616,N_199);
nand U1829 (N_1829,N_451,N_553);
xor U1830 (N_1830,N_878,N_805);
and U1831 (N_1831,N_988,N_872);
or U1832 (N_1832,N_149,N_440);
xnor U1833 (N_1833,N_366,N_826);
and U1834 (N_1834,N_96,N_209);
or U1835 (N_1835,N_684,N_424);
nand U1836 (N_1836,N_863,N_430);
and U1837 (N_1837,N_491,N_388);
xor U1838 (N_1838,N_991,N_833);
nand U1839 (N_1839,N_663,N_924);
and U1840 (N_1840,N_106,N_549);
nor U1841 (N_1841,N_689,N_518);
or U1842 (N_1842,N_460,N_968);
nor U1843 (N_1843,N_910,N_75);
or U1844 (N_1844,N_594,N_240);
nand U1845 (N_1845,N_662,N_56);
nand U1846 (N_1846,N_129,N_430);
nand U1847 (N_1847,N_416,N_335);
nor U1848 (N_1848,N_760,N_2);
or U1849 (N_1849,N_866,N_403);
nand U1850 (N_1850,N_449,N_678);
and U1851 (N_1851,N_293,N_660);
xor U1852 (N_1852,N_225,N_306);
nor U1853 (N_1853,N_851,N_420);
or U1854 (N_1854,N_515,N_465);
and U1855 (N_1855,N_23,N_621);
nand U1856 (N_1856,N_601,N_181);
xnor U1857 (N_1857,N_167,N_917);
nand U1858 (N_1858,N_99,N_544);
xor U1859 (N_1859,N_551,N_290);
xnor U1860 (N_1860,N_866,N_541);
nor U1861 (N_1861,N_201,N_257);
or U1862 (N_1862,N_307,N_555);
nand U1863 (N_1863,N_592,N_48);
xnor U1864 (N_1864,N_522,N_774);
nor U1865 (N_1865,N_483,N_902);
nand U1866 (N_1866,N_738,N_528);
nand U1867 (N_1867,N_741,N_944);
xor U1868 (N_1868,N_776,N_777);
xnor U1869 (N_1869,N_907,N_423);
nor U1870 (N_1870,N_744,N_348);
and U1871 (N_1871,N_186,N_486);
nor U1872 (N_1872,N_564,N_603);
and U1873 (N_1873,N_692,N_472);
or U1874 (N_1874,N_655,N_67);
or U1875 (N_1875,N_473,N_429);
and U1876 (N_1876,N_312,N_583);
xor U1877 (N_1877,N_772,N_324);
nand U1878 (N_1878,N_713,N_708);
or U1879 (N_1879,N_551,N_662);
xnor U1880 (N_1880,N_628,N_829);
nand U1881 (N_1881,N_475,N_895);
nand U1882 (N_1882,N_392,N_466);
nand U1883 (N_1883,N_663,N_302);
xor U1884 (N_1884,N_77,N_395);
nand U1885 (N_1885,N_961,N_78);
and U1886 (N_1886,N_36,N_208);
and U1887 (N_1887,N_402,N_785);
nand U1888 (N_1888,N_708,N_786);
or U1889 (N_1889,N_915,N_303);
or U1890 (N_1890,N_719,N_885);
xnor U1891 (N_1891,N_197,N_941);
or U1892 (N_1892,N_322,N_208);
or U1893 (N_1893,N_294,N_287);
or U1894 (N_1894,N_432,N_677);
and U1895 (N_1895,N_564,N_695);
xor U1896 (N_1896,N_406,N_752);
nand U1897 (N_1897,N_860,N_460);
xor U1898 (N_1898,N_808,N_994);
xor U1899 (N_1899,N_995,N_323);
or U1900 (N_1900,N_565,N_781);
or U1901 (N_1901,N_853,N_176);
or U1902 (N_1902,N_223,N_286);
xor U1903 (N_1903,N_206,N_473);
or U1904 (N_1904,N_211,N_514);
nand U1905 (N_1905,N_171,N_568);
or U1906 (N_1906,N_151,N_126);
nor U1907 (N_1907,N_778,N_411);
and U1908 (N_1908,N_227,N_168);
xnor U1909 (N_1909,N_79,N_760);
and U1910 (N_1910,N_721,N_786);
xnor U1911 (N_1911,N_366,N_0);
nor U1912 (N_1912,N_592,N_35);
or U1913 (N_1913,N_334,N_427);
nand U1914 (N_1914,N_654,N_677);
or U1915 (N_1915,N_366,N_919);
or U1916 (N_1916,N_897,N_317);
and U1917 (N_1917,N_87,N_140);
and U1918 (N_1918,N_494,N_515);
nor U1919 (N_1919,N_560,N_200);
nand U1920 (N_1920,N_861,N_351);
nor U1921 (N_1921,N_310,N_343);
or U1922 (N_1922,N_593,N_656);
or U1923 (N_1923,N_126,N_197);
nand U1924 (N_1924,N_798,N_254);
and U1925 (N_1925,N_664,N_325);
and U1926 (N_1926,N_399,N_385);
nand U1927 (N_1927,N_735,N_579);
xnor U1928 (N_1928,N_128,N_237);
nand U1929 (N_1929,N_368,N_939);
and U1930 (N_1930,N_722,N_181);
nor U1931 (N_1931,N_535,N_875);
and U1932 (N_1932,N_195,N_676);
nand U1933 (N_1933,N_972,N_476);
nand U1934 (N_1934,N_827,N_396);
or U1935 (N_1935,N_561,N_675);
or U1936 (N_1936,N_754,N_609);
and U1937 (N_1937,N_586,N_54);
nand U1938 (N_1938,N_41,N_299);
and U1939 (N_1939,N_915,N_686);
nand U1940 (N_1940,N_550,N_699);
and U1941 (N_1941,N_502,N_591);
or U1942 (N_1942,N_248,N_680);
nand U1943 (N_1943,N_582,N_880);
and U1944 (N_1944,N_158,N_198);
nor U1945 (N_1945,N_455,N_38);
xnor U1946 (N_1946,N_173,N_138);
xor U1947 (N_1947,N_150,N_609);
and U1948 (N_1948,N_348,N_430);
or U1949 (N_1949,N_155,N_465);
nor U1950 (N_1950,N_508,N_538);
nand U1951 (N_1951,N_809,N_501);
xnor U1952 (N_1952,N_985,N_212);
nand U1953 (N_1953,N_722,N_551);
or U1954 (N_1954,N_305,N_668);
and U1955 (N_1955,N_21,N_12);
xor U1956 (N_1956,N_642,N_4);
xnor U1957 (N_1957,N_618,N_120);
nor U1958 (N_1958,N_641,N_77);
xnor U1959 (N_1959,N_294,N_26);
nor U1960 (N_1960,N_440,N_624);
or U1961 (N_1961,N_181,N_799);
nand U1962 (N_1962,N_694,N_944);
and U1963 (N_1963,N_144,N_798);
xnor U1964 (N_1964,N_73,N_886);
and U1965 (N_1965,N_219,N_852);
nand U1966 (N_1966,N_439,N_515);
xor U1967 (N_1967,N_680,N_955);
nor U1968 (N_1968,N_542,N_8);
or U1969 (N_1969,N_593,N_603);
nand U1970 (N_1970,N_273,N_924);
or U1971 (N_1971,N_37,N_327);
and U1972 (N_1972,N_411,N_441);
or U1973 (N_1973,N_86,N_227);
nor U1974 (N_1974,N_400,N_708);
or U1975 (N_1975,N_492,N_617);
nand U1976 (N_1976,N_718,N_359);
nand U1977 (N_1977,N_881,N_440);
nand U1978 (N_1978,N_835,N_866);
and U1979 (N_1979,N_885,N_529);
or U1980 (N_1980,N_380,N_411);
nand U1981 (N_1981,N_55,N_747);
xor U1982 (N_1982,N_155,N_93);
xnor U1983 (N_1983,N_302,N_639);
or U1984 (N_1984,N_870,N_686);
nand U1985 (N_1985,N_255,N_624);
nor U1986 (N_1986,N_988,N_267);
nand U1987 (N_1987,N_498,N_169);
nand U1988 (N_1988,N_268,N_768);
xnor U1989 (N_1989,N_143,N_483);
and U1990 (N_1990,N_173,N_668);
xor U1991 (N_1991,N_67,N_847);
nor U1992 (N_1992,N_681,N_456);
or U1993 (N_1993,N_358,N_116);
and U1994 (N_1994,N_13,N_262);
or U1995 (N_1995,N_174,N_52);
nor U1996 (N_1996,N_416,N_689);
xor U1997 (N_1997,N_414,N_703);
nand U1998 (N_1998,N_334,N_559);
nand U1999 (N_1999,N_219,N_672);
xnor U2000 (N_2000,N_1261,N_1539);
and U2001 (N_2001,N_1784,N_1637);
nand U2002 (N_2002,N_1945,N_1478);
nor U2003 (N_2003,N_1781,N_1812);
and U2004 (N_2004,N_1880,N_1447);
or U2005 (N_2005,N_1832,N_1062);
or U2006 (N_2006,N_1077,N_1896);
and U2007 (N_2007,N_1234,N_1434);
or U2008 (N_2008,N_1382,N_1170);
and U2009 (N_2009,N_1425,N_1676);
and U2010 (N_2010,N_1758,N_1599);
and U2011 (N_2011,N_1641,N_1767);
nor U2012 (N_2012,N_1191,N_1356);
and U2013 (N_2013,N_1439,N_1757);
nand U2014 (N_2014,N_1888,N_1215);
or U2015 (N_2015,N_1472,N_1798);
nor U2016 (N_2016,N_1760,N_1881);
and U2017 (N_2017,N_1253,N_1890);
xor U2018 (N_2018,N_1803,N_1155);
xor U2019 (N_2019,N_1931,N_1403);
xor U2020 (N_2020,N_1932,N_1492);
and U2021 (N_2021,N_1840,N_1267);
nand U2022 (N_2022,N_1994,N_1202);
nor U2023 (N_2023,N_1393,N_1631);
xor U2024 (N_2024,N_1795,N_1033);
and U2025 (N_2025,N_1604,N_1870);
and U2026 (N_2026,N_1441,N_1058);
xnor U2027 (N_2027,N_1534,N_1216);
nand U2028 (N_2028,N_1969,N_1011);
and U2029 (N_2029,N_1728,N_1893);
and U2030 (N_2030,N_1823,N_1834);
and U2031 (N_2031,N_1943,N_1491);
nand U2032 (N_2032,N_1620,N_1293);
nor U2033 (N_2033,N_1549,N_1868);
and U2034 (N_2034,N_1410,N_1626);
or U2035 (N_2035,N_1362,N_1379);
nand U2036 (N_2036,N_1486,N_1642);
or U2037 (N_2037,N_1804,N_1210);
and U2038 (N_2038,N_1591,N_1465);
nor U2039 (N_2039,N_1424,N_1181);
and U2040 (N_2040,N_1041,N_1948);
nor U2041 (N_2041,N_1968,N_1493);
nor U2042 (N_2042,N_1302,N_1712);
or U2043 (N_2043,N_1962,N_1485);
and U2044 (N_2044,N_1756,N_1245);
or U2045 (N_2045,N_1652,N_1929);
and U2046 (N_2046,N_1583,N_1866);
and U2047 (N_2047,N_1231,N_1954);
and U2048 (N_2048,N_1100,N_1937);
nand U2049 (N_2049,N_1841,N_1061);
and U2050 (N_2050,N_1076,N_1350);
and U2051 (N_2051,N_1214,N_1071);
and U2052 (N_2052,N_1108,N_1902);
nor U2053 (N_2053,N_1819,N_1649);
or U2054 (N_2054,N_1917,N_1698);
nor U2055 (N_2055,N_1960,N_1279);
nor U2056 (N_2056,N_1653,N_1249);
nand U2057 (N_2057,N_1675,N_1255);
and U2058 (N_2058,N_1411,N_1312);
nor U2059 (N_2059,N_1254,N_1034);
xor U2060 (N_2060,N_1974,N_1188);
or U2061 (N_2061,N_1487,N_1734);
xor U2062 (N_2062,N_1276,N_1999);
xor U2063 (N_2063,N_1218,N_1225);
or U2064 (N_2064,N_1783,N_1855);
or U2065 (N_2065,N_1949,N_1295);
or U2066 (N_2066,N_1050,N_1311);
nor U2067 (N_2067,N_1891,N_1294);
nand U2068 (N_2068,N_1520,N_1369);
nand U2069 (N_2069,N_1262,N_1420);
or U2070 (N_2070,N_1754,N_1205);
nand U2071 (N_2071,N_1574,N_1019);
nor U2072 (N_2072,N_1512,N_1814);
nor U2073 (N_2073,N_1538,N_1887);
nor U2074 (N_2074,N_1407,N_1501);
xnor U2075 (N_2075,N_1739,N_1703);
or U2076 (N_2076,N_1115,N_1044);
nor U2077 (N_2077,N_1381,N_1087);
nor U2078 (N_2078,N_1506,N_1094);
or U2079 (N_2079,N_1685,N_1828);
or U2080 (N_2080,N_1633,N_1707);
nand U2081 (N_2081,N_1730,N_1180);
nor U2082 (N_2082,N_1149,N_1313);
xor U2083 (N_2083,N_1632,N_1030);
xor U2084 (N_2084,N_1553,N_1341);
and U2085 (N_2085,N_1608,N_1263);
nand U2086 (N_2086,N_1530,N_1093);
nand U2087 (N_2087,N_1628,N_1102);
or U2088 (N_2088,N_1724,N_1809);
xor U2089 (N_2089,N_1152,N_1151);
and U2090 (N_2090,N_1168,N_1482);
and U2091 (N_2091,N_1014,N_1377);
and U2092 (N_2092,N_1413,N_1397);
nor U2093 (N_2093,N_1127,N_1933);
and U2094 (N_2094,N_1959,N_1680);
nand U2095 (N_2095,N_1119,N_1727);
xnor U2096 (N_2096,N_1004,N_1694);
nor U2097 (N_2097,N_1989,N_1519);
or U2098 (N_2098,N_1836,N_1372);
xnor U2099 (N_2099,N_1113,N_1390);
nand U2100 (N_2100,N_1750,N_1616);
or U2101 (N_2101,N_1634,N_1444);
and U2102 (N_2102,N_1722,N_1572);
nor U2103 (N_2103,N_1164,N_1726);
and U2104 (N_2104,N_1250,N_1349);
nor U2105 (N_2105,N_1097,N_1230);
xnor U2106 (N_2106,N_1961,N_1330);
nand U2107 (N_2107,N_1045,N_1473);
xnor U2108 (N_2108,N_1299,N_1923);
nand U2109 (N_2109,N_1301,N_1072);
or U2110 (N_2110,N_1701,N_1822);
or U2111 (N_2111,N_1592,N_1010);
nand U2112 (N_2112,N_1587,N_1236);
xnor U2113 (N_2113,N_1308,N_1412);
xnor U2114 (N_2114,N_1281,N_1913);
xor U2115 (N_2115,N_1359,N_1342);
nand U2116 (N_2116,N_1008,N_1209);
or U2117 (N_2117,N_1057,N_1875);
or U2118 (N_2118,N_1507,N_1017);
nor U2119 (N_2119,N_1638,N_1082);
and U2120 (N_2120,N_1557,N_1455);
or U2121 (N_2121,N_1612,N_1398);
and U2122 (N_2122,N_1112,N_1762);
xnor U2123 (N_2123,N_1116,N_1047);
or U2124 (N_2124,N_1842,N_1785);
and U2125 (N_2125,N_1233,N_1623);
or U2126 (N_2126,N_1856,N_1835);
and U2127 (N_2127,N_1496,N_1720);
nand U2128 (N_2128,N_1273,N_1851);
nand U2129 (N_2129,N_1521,N_1993);
xnor U2130 (N_2130,N_1597,N_1857);
xnor U2131 (N_2131,N_1192,N_1195);
xor U2132 (N_2132,N_1600,N_1338);
nor U2133 (N_2133,N_1667,N_1663);
or U2134 (N_2134,N_1918,N_1714);
or U2135 (N_2135,N_1665,N_1981);
nand U2136 (N_2136,N_1055,N_1169);
or U2137 (N_2137,N_1298,N_1443);
or U2138 (N_2138,N_1158,N_1001);
and U2139 (N_2139,N_1049,N_1518);
nand U2140 (N_2140,N_1440,N_1345);
nor U2141 (N_2141,N_1309,N_1458);
xnor U2142 (N_2142,N_1753,N_1573);
or U2143 (N_2143,N_1366,N_1992);
nor U2144 (N_2144,N_1167,N_1297);
or U2145 (N_2145,N_1884,N_1522);
nor U2146 (N_2146,N_1334,N_1636);
nand U2147 (N_2147,N_1246,N_1548);
nor U2148 (N_2148,N_1787,N_1498);
nor U2149 (N_2149,N_1159,N_1860);
or U2150 (N_2150,N_1833,N_1421);
nand U2151 (N_2151,N_1740,N_1752);
nand U2152 (N_2152,N_1380,N_1029);
nand U2153 (N_2153,N_1952,N_1805);
xor U2154 (N_2154,N_1602,N_1024);
nor U2155 (N_2155,N_1679,N_1640);
xnor U2156 (N_2156,N_1817,N_1831);
and U2157 (N_2157,N_1474,N_1850);
nor U2158 (N_2158,N_1448,N_1596);
and U2159 (N_2159,N_1509,N_1776);
or U2160 (N_2160,N_1562,N_1985);
nor U2161 (N_2161,N_1537,N_1373);
xnor U2162 (N_2162,N_1419,N_1328);
nor U2163 (N_2163,N_1260,N_1069);
nand U2164 (N_2164,N_1723,N_1639);
xor U2165 (N_2165,N_1745,N_1394);
or U2166 (N_2166,N_1532,N_1696);
or U2167 (N_2167,N_1399,N_1074);
nor U2168 (N_2168,N_1609,N_1508);
xnor U2169 (N_2169,N_1437,N_1543);
xnor U2170 (N_2170,N_1593,N_1105);
and U2171 (N_2171,N_1089,N_1883);
xnor U2172 (N_2172,N_1688,N_1830);
or U2173 (N_2173,N_1934,N_1719);
nand U2174 (N_2174,N_1775,N_1683);
or U2175 (N_2175,N_1416,N_1898);
nand U2176 (N_2176,N_1285,N_1436);
nor U2177 (N_2177,N_1237,N_1497);
and U2178 (N_2178,N_1951,N_1171);
or U2179 (N_2179,N_1315,N_1141);
xor U2180 (N_2180,N_1031,N_1438);
and U2181 (N_2181,N_1577,N_1348);
xor U2182 (N_2182,N_1361,N_1614);
xnor U2183 (N_2183,N_1384,N_1963);
nor U2184 (N_2184,N_1729,N_1671);
xnor U2185 (N_2185,N_1147,N_1204);
and U2186 (N_2186,N_1207,N_1721);
and U2187 (N_2187,N_1343,N_1489);
nor U2188 (N_2188,N_1930,N_1846);
and U2189 (N_2189,N_1125,N_1241);
xor U2190 (N_2190,N_1938,N_1504);
and U2191 (N_2191,N_1669,N_1920);
xnor U2192 (N_2192,N_1161,N_1409);
or U2193 (N_2193,N_1575,N_1725);
nor U2194 (N_2194,N_1759,N_1408);
or U2195 (N_2195,N_1924,N_1184);
or U2196 (N_2196,N_1582,N_1718);
and U2197 (N_2197,N_1477,N_1621);
and U2198 (N_2198,N_1461,N_1792);
xor U2199 (N_2199,N_1091,N_1217);
or U2200 (N_2200,N_1405,N_1429);
xnor U2201 (N_2201,N_1568,N_1259);
xor U2202 (N_2202,N_1432,N_1526);
or U2203 (N_2203,N_1736,N_1551);
nor U2204 (N_2204,N_1956,N_1874);
nor U2205 (N_2205,N_1743,N_1148);
nand U2206 (N_2206,N_1107,N_1535);
or U2207 (N_2207,N_1678,N_1660);
or U2208 (N_2208,N_1916,N_1370);
nor U2209 (N_2209,N_1821,N_1702);
xor U2210 (N_2210,N_1475,N_1305);
nand U2211 (N_2211,N_1120,N_1677);
xor U2212 (N_2212,N_1670,N_1879);
nor U2213 (N_2213,N_1153,N_1764);
nor U2214 (N_2214,N_1877,N_1513);
xnor U2215 (N_2215,N_1777,N_1386);
nor U2216 (N_2216,N_1732,N_1337);
xnor U2217 (N_2217,N_1456,N_1808);
nand U2218 (N_2218,N_1054,N_1894);
xor U2219 (N_2219,N_1163,N_1627);
nor U2220 (N_2220,N_1690,N_1901);
and U2221 (N_2221,N_1065,N_1570);
nand U2222 (N_2222,N_1975,N_1865);
or U2223 (N_2223,N_1912,N_1709);
nor U2224 (N_2224,N_1053,N_1326);
xor U2225 (N_2225,N_1738,N_1121);
nand U2226 (N_2226,N_1385,N_1598);
nor U2227 (N_2227,N_1027,N_1650);
xnor U2228 (N_2228,N_1389,N_1092);
or U2229 (N_2229,N_1189,N_1873);
nor U2230 (N_2230,N_1067,N_1561);
nor U2231 (N_2231,N_1942,N_1300);
or U2232 (N_2232,N_1275,N_1569);
and U2233 (N_2233,N_1283,N_1778);
and U2234 (N_2234,N_1023,N_1769);
xor U2235 (N_2235,N_1186,N_1987);
nor U2236 (N_2236,N_1606,N_1950);
nor U2237 (N_2237,N_1200,N_1944);
or U2238 (N_2238,N_1242,N_1862);
xnor U2239 (N_2239,N_1051,N_1318);
and U2240 (N_2240,N_1415,N_1026);
or U2241 (N_2241,N_1247,N_1829);
nand U2242 (N_2242,N_1414,N_1287);
or U2243 (N_2243,N_1863,N_1317);
and U2244 (N_2244,N_1861,N_1172);
nor U2245 (N_2245,N_1220,N_1126);
and U2246 (N_2246,N_1693,N_1580);
nand U2247 (N_2247,N_1355,N_1815);
xnor U2248 (N_2248,N_1387,N_1375);
nor U2249 (N_2249,N_1935,N_1321);
nor U2250 (N_2250,N_1006,N_1015);
nand U2251 (N_2251,N_1248,N_1132);
and U2252 (N_2252,N_1523,N_1586);
xnor U2253 (N_2253,N_1555,N_1040);
or U2254 (N_2254,N_1201,N_1183);
xnor U2255 (N_2255,N_1463,N_1766);
or U2256 (N_2256,N_1936,N_1354);
and U2257 (N_2257,N_1666,N_1325);
nand U2258 (N_2258,N_1129,N_1578);
or U2259 (N_2259,N_1590,N_1635);
or U2260 (N_2260,N_1176,N_1048);
and U2261 (N_2261,N_1657,N_1266);
nor U2262 (N_2262,N_1229,N_1998);
or U2263 (N_2263,N_1700,N_1824);
nor U2264 (N_2264,N_1774,N_1142);
and U2265 (N_2265,N_1624,N_1540);
nand U2266 (N_2266,N_1779,N_1388);
nor U2267 (N_2267,N_1547,N_1018);
xnor U2268 (N_2268,N_1905,N_1022);
and U2269 (N_2269,N_1615,N_1630);
or U2270 (N_2270,N_1307,N_1643);
or U2271 (N_2271,N_1079,N_1344);
and U2272 (N_2272,N_1859,N_1768);
or U2273 (N_2273,N_1052,N_1571);
xnor U2274 (N_2274,N_1222,N_1140);
and U2275 (N_2275,N_1088,N_1695);
and U2276 (N_2276,N_1117,N_1291);
nand U2277 (N_2277,N_1005,N_1849);
nor U2278 (N_2278,N_1658,N_1122);
or U2279 (N_2279,N_1710,N_1687);
or U2280 (N_2280,N_1984,N_1617);
xor U2281 (N_2281,N_1716,N_1043);
xor U2282 (N_2282,N_1763,N_1320);
or U2283 (N_2283,N_1316,N_1502);
and U2284 (N_2284,N_1426,N_1194);
xor U2285 (N_2285,N_1955,N_1042);
nand U2286 (N_2286,N_1452,N_1322);
or U2287 (N_2287,N_1111,N_1741);
nor U2288 (N_2288,N_1601,N_1751);
nor U2289 (N_2289,N_1682,N_1290);
nand U2290 (N_2290,N_1545,N_1737);
and U2291 (N_2291,N_1910,N_1251);
nor U2292 (N_2292,N_1681,N_1123);
or U2293 (N_2293,N_1542,N_1032);
xor U2294 (N_2294,N_1697,N_1565);
or U2295 (N_2295,N_1078,N_1957);
or U2296 (N_2296,N_1454,N_1813);
nand U2297 (N_2297,N_1396,N_1558);
nor U2298 (N_2298,N_1106,N_1495);
nand U2299 (N_2299,N_1128,N_1585);
nor U2300 (N_2300,N_1919,N_1796);
nand U2301 (N_2301,N_1903,N_1749);
and U2302 (N_2302,N_1156,N_1733);
or U2303 (N_2303,N_1889,N_1619);
nor U2304 (N_2304,N_1319,N_1464);
xnor U2305 (N_2305,N_1466,N_1904);
xnor U2306 (N_2306,N_1235,N_1646);
nand U2307 (N_2307,N_1073,N_1310);
xor U2308 (N_2308,N_1673,N_1782);
nor U2309 (N_2309,N_1038,N_1327);
or U2310 (N_2310,N_1818,N_1848);
xnor U2311 (N_2311,N_1797,N_1978);
or U2312 (N_2312,N_1885,N_1039);
nor U2313 (N_2313,N_1909,N_1357);
or U2314 (N_2314,N_1715,N_1986);
xor U2315 (N_2315,N_1160,N_1699);
xor U2316 (N_2316,N_1193,N_1471);
xor U2317 (N_2317,N_1886,N_1187);
xnor U2318 (N_2318,N_1780,N_1016);
and U2319 (N_2319,N_1668,N_1525);
or U2320 (N_2320,N_1811,N_1199);
or U2321 (N_2321,N_1906,N_1566);
nor U2322 (N_2322,N_1581,N_1329);
nor U2323 (N_2323,N_1806,N_1289);
xor U2324 (N_2324,N_1915,N_1939);
nand U2325 (N_2325,N_1661,N_1672);
xor U2326 (N_2326,N_1445,N_1114);
xnor U2327 (N_2327,N_1450,N_1644);
xnor U2328 (N_2328,N_1747,N_1144);
or U2329 (N_2329,N_1922,N_1244);
nor U2330 (N_2330,N_1940,N_1371);
nor U2331 (N_2331,N_1983,N_1826);
or U2332 (N_2332,N_1820,N_1869);
nand U2333 (N_2333,N_1376,N_1175);
or U2334 (N_2334,N_1124,N_1304);
xnor U2335 (N_2335,N_1101,N_1368);
or U2336 (N_2336,N_1481,N_1895);
nand U2337 (N_2337,N_1203,N_1265);
nand U2338 (N_2338,N_1219,N_1059);
and U2339 (N_2339,N_1353,N_1958);
xor U2340 (N_2340,N_1284,N_1208);
nand U2341 (N_2341,N_1980,N_1790);
xnor U2342 (N_2342,N_1772,N_1206);
xor U2343 (N_2343,N_1662,N_1706);
and U2344 (N_2344,N_1146,N_1793);
or U2345 (N_2345,N_1392,N_1395);
and U2346 (N_2346,N_1911,N_1576);
nand U2347 (N_2347,N_1527,N_1647);
nand U2348 (N_2348,N_1595,N_1878);
and U2349 (N_2349,N_1402,N_1401);
and U2350 (N_2350,N_1544,N_1705);
and U2351 (N_2351,N_1801,N_1339);
xnor U2352 (N_2352,N_1995,N_1516);
nand U2353 (N_2353,N_1212,N_1360);
nand U2354 (N_2354,N_1135,N_1997);
nand U2355 (N_2355,N_1098,N_1303);
nor U2356 (N_2356,N_1269,N_1374);
xnor U2357 (N_2357,N_1358,N_1858);
nor U2358 (N_2358,N_1442,N_1037);
and U2359 (N_2359,N_1282,N_1224);
and U2360 (N_2360,N_1925,N_1084);
and U2361 (N_2361,N_1063,N_1131);
nor U2362 (N_2362,N_1258,N_1136);
xor U2363 (N_2363,N_1844,N_1564);
nor U2364 (N_2364,N_1988,N_1070);
nor U2365 (N_2365,N_1854,N_1347);
or U2366 (N_2366,N_1046,N_1791);
nand U2367 (N_2367,N_1611,N_1839);
nor U2368 (N_2368,N_1190,N_1789);
nand U2369 (N_2369,N_1451,N_1272);
nand U2370 (N_2370,N_1449,N_1145);
xor U2371 (N_2371,N_1967,N_1288);
xor U2372 (N_2372,N_1268,N_1239);
nand U2373 (N_2373,N_1280,N_1060);
or U2374 (N_2374,N_1499,N_1541);
nand U2375 (N_2375,N_1927,N_1400);
or U2376 (N_2376,N_1810,N_1314);
and U2377 (N_2377,N_1800,N_1166);
and U2378 (N_2378,N_1579,N_1264);
nor U2379 (N_2379,N_1086,N_1692);
or U2380 (N_2380,N_1686,N_1154);
xor U2381 (N_2381,N_1391,N_1363);
nand U2382 (N_2382,N_1966,N_1383);
nand U2383 (N_2383,N_1603,N_1185);
xor U2384 (N_2384,N_1742,N_1770);
xnor U2385 (N_2385,N_1104,N_1517);
and U2386 (N_2386,N_1428,N_1470);
nand U2387 (N_2387,N_1157,N_1174);
xnor U2388 (N_2388,N_1457,N_1713);
and U2389 (N_2389,N_1232,N_1226);
nor U2390 (N_2390,N_1629,N_1531);
or U2391 (N_2391,N_1021,N_1035);
or U2392 (N_2392,N_1982,N_1684);
and U2393 (N_2393,N_1505,N_1378);
and U2394 (N_2394,N_1080,N_1648);
nor U2395 (N_2395,N_1761,N_1941);
nand U2396 (N_2396,N_1735,N_1947);
xor U2397 (N_2397,N_1483,N_1198);
nor U2398 (N_2398,N_1872,N_1965);
xor U2399 (N_2399,N_1510,N_1946);
nand U2400 (N_2400,N_1589,N_1744);
xor U2401 (N_2401,N_1150,N_1099);
and U2402 (N_2402,N_1028,N_1335);
or U2403 (N_2403,N_1351,N_1484);
nand U2404 (N_2404,N_1816,N_1921);
nor U2405 (N_2405,N_1138,N_1588);
xor U2406 (N_2406,N_1433,N_1173);
nor U2407 (N_2407,N_1556,N_1252);
and U2408 (N_2408,N_1876,N_1332);
nand U2409 (N_2409,N_1068,N_1036);
nand U2410 (N_2410,N_1837,N_1899);
and U2411 (N_2411,N_1794,N_1012);
and U2412 (N_2412,N_1552,N_1607);
xor U2413 (N_2413,N_1559,N_1900);
or U2414 (N_2414,N_1064,N_1137);
nor U2415 (N_2415,N_1563,N_1196);
nand U2416 (N_2416,N_1656,N_1469);
and U2417 (N_2417,N_1867,N_1807);
nor U2418 (N_2418,N_1897,N_1500);
and U2419 (N_2419,N_1352,N_1278);
xor U2420 (N_2420,N_1179,N_1838);
nand U2421 (N_2421,N_1085,N_1066);
nand U2422 (N_2422,N_1926,N_1480);
or U2423 (N_2423,N_1277,N_1056);
nor U2424 (N_2424,N_1970,N_1488);
and U2425 (N_2425,N_1594,N_1528);
and U2426 (N_2426,N_1013,N_1964);
or U2427 (N_2427,N_1406,N_1691);
nor U2428 (N_2428,N_1009,N_1462);
or U2429 (N_2429,N_1007,N_1645);
xnor U2430 (N_2430,N_1109,N_1468);
nand U2431 (N_2431,N_1422,N_1367);
and U2432 (N_2432,N_1651,N_1240);
nor U2433 (N_2433,N_1417,N_1953);
nand U2434 (N_2434,N_1130,N_1286);
or U2435 (N_2435,N_1550,N_1427);
and U2436 (N_2436,N_1223,N_1908);
and U2437 (N_2437,N_1227,N_1584);
nand U2438 (N_2438,N_1802,N_1524);
nor U2439 (N_2439,N_1134,N_1882);
nand U2440 (N_2440,N_1095,N_1976);
nor U2441 (N_2441,N_1081,N_1178);
xor U2442 (N_2442,N_1659,N_1825);
or U2443 (N_2443,N_1708,N_1103);
xor U2444 (N_2444,N_1536,N_1165);
or U2445 (N_2445,N_1711,N_1000);
or U2446 (N_2446,N_1622,N_1689);
and U2447 (N_2447,N_1025,N_1748);
and U2448 (N_2448,N_1479,N_1972);
xor U2449 (N_2449,N_1162,N_1256);
and U2450 (N_2450,N_1211,N_1625);
and U2451 (N_2451,N_1567,N_1843);
nand U2452 (N_2452,N_1430,N_1746);
nor U2453 (N_2453,N_1323,N_1853);
nand U2454 (N_2454,N_1133,N_1554);
nor U2455 (N_2455,N_1143,N_1864);
xnor U2456 (N_2456,N_1213,N_1365);
nand U2457 (N_2457,N_1618,N_1610);
and U2458 (N_2458,N_1423,N_1075);
nor U2459 (N_2459,N_1182,N_1446);
nor U2460 (N_2460,N_1871,N_1973);
or U2461 (N_2461,N_1238,N_1336);
or U2462 (N_2462,N_1096,N_1331);
xor U2463 (N_2463,N_1845,N_1243);
and U2464 (N_2464,N_1605,N_1514);
or U2465 (N_2465,N_1333,N_1655);
nand U2466 (N_2466,N_1453,N_1274);
or U2467 (N_2467,N_1533,N_1755);
nand U2468 (N_2468,N_1788,N_1418);
or U2469 (N_2469,N_1346,N_1503);
nor U2470 (N_2470,N_1296,N_1515);
and U2471 (N_2471,N_1529,N_1292);
xnor U2472 (N_2472,N_1827,N_1459);
nor U2473 (N_2473,N_1257,N_1914);
xnor U2474 (N_2474,N_1731,N_1460);
xor U2475 (N_2475,N_1364,N_1340);
or U2476 (N_2476,N_1090,N_1991);
nand U2477 (N_2477,N_1083,N_1110);
nand U2478 (N_2478,N_1765,N_1560);
nor U2479 (N_2479,N_1892,N_1020);
and U2480 (N_2480,N_1907,N_1977);
or U2481 (N_2481,N_1654,N_1270);
nand U2482 (N_2482,N_1971,N_1467);
and U2483 (N_2483,N_1852,N_1431);
or U2484 (N_2484,N_1003,N_1228);
or U2485 (N_2485,N_1476,N_1511);
nand U2486 (N_2486,N_1002,N_1847);
nor U2487 (N_2487,N_1118,N_1786);
xnor U2488 (N_2488,N_1771,N_1139);
xnor U2489 (N_2489,N_1799,N_1773);
xnor U2490 (N_2490,N_1306,N_1990);
and U2491 (N_2491,N_1435,N_1197);
xor U2492 (N_2492,N_1546,N_1704);
xnor U2493 (N_2493,N_1613,N_1490);
nor U2494 (N_2494,N_1717,N_1404);
or U2495 (N_2495,N_1324,N_1979);
and U2496 (N_2496,N_1494,N_1177);
or U2497 (N_2497,N_1928,N_1674);
xor U2498 (N_2498,N_1271,N_1996);
nand U2499 (N_2499,N_1221,N_1664);
or U2500 (N_2500,N_1155,N_1753);
nand U2501 (N_2501,N_1614,N_1710);
xnor U2502 (N_2502,N_1114,N_1355);
or U2503 (N_2503,N_1015,N_1096);
or U2504 (N_2504,N_1274,N_1946);
and U2505 (N_2505,N_1330,N_1763);
nand U2506 (N_2506,N_1936,N_1107);
xnor U2507 (N_2507,N_1627,N_1298);
or U2508 (N_2508,N_1807,N_1603);
xor U2509 (N_2509,N_1115,N_1465);
xor U2510 (N_2510,N_1460,N_1323);
xnor U2511 (N_2511,N_1602,N_1091);
nand U2512 (N_2512,N_1526,N_1887);
or U2513 (N_2513,N_1076,N_1750);
nand U2514 (N_2514,N_1488,N_1943);
or U2515 (N_2515,N_1040,N_1846);
or U2516 (N_2516,N_1003,N_1464);
nand U2517 (N_2517,N_1161,N_1312);
and U2518 (N_2518,N_1197,N_1858);
nand U2519 (N_2519,N_1672,N_1275);
xnor U2520 (N_2520,N_1945,N_1036);
nand U2521 (N_2521,N_1599,N_1504);
or U2522 (N_2522,N_1899,N_1308);
nor U2523 (N_2523,N_1788,N_1801);
xnor U2524 (N_2524,N_1778,N_1648);
and U2525 (N_2525,N_1001,N_1854);
nand U2526 (N_2526,N_1541,N_1950);
xor U2527 (N_2527,N_1070,N_1009);
or U2528 (N_2528,N_1863,N_1100);
and U2529 (N_2529,N_1545,N_1174);
nand U2530 (N_2530,N_1455,N_1329);
or U2531 (N_2531,N_1520,N_1880);
and U2532 (N_2532,N_1212,N_1685);
nor U2533 (N_2533,N_1306,N_1728);
xor U2534 (N_2534,N_1972,N_1533);
or U2535 (N_2535,N_1069,N_1921);
and U2536 (N_2536,N_1342,N_1843);
or U2537 (N_2537,N_1798,N_1296);
xor U2538 (N_2538,N_1803,N_1952);
or U2539 (N_2539,N_1661,N_1645);
xor U2540 (N_2540,N_1045,N_1617);
and U2541 (N_2541,N_1110,N_1547);
nand U2542 (N_2542,N_1378,N_1959);
nand U2543 (N_2543,N_1936,N_1613);
or U2544 (N_2544,N_1674,N_1516);
nand U2545 (N_2545,N_1177,N_1041);
and U2546 (N_2546,N_1587,N_1260);
nand U2547 (N_2547,N_1500,N_1322);
nor U2548 (N_2548,N_1208,N_1938);
nor U2549 (N_2549,N_1669,N_1147);
nand U2550 (N_2550,N_1859,N_1895);
nor U2551 (N_2551,N_1828,N_1383);
nor U2552 (N_2552,N_1592,N_1763);
nor U2553 (N_2553,N_1060,N_1113);
xnor U2554 (N_2554,N_1380,N_1678);
and U2555 (N_2555,N_1201,N_1205);
and U2556 (N_2556,N_1217,N_1470);
xnor U2557 (N_2557,N_1908,N_1814);
or U2558 (N_2558,N_1181,N_1747);
xnor U2559 (N_2559,N_1094,N_1517);
and U2560 (N_2560,N_1764,N_1894);
or U2561 (N_2561,N_1983,N_1388);
and U2562 (N_2562,N_1069,N_1405);
xnor U2563 (N_2563,N_1083,N_1638);
nor U2564 (N_2564,N_1142,N_1497);
and U2565 (N_2565,N_1181,N_1509);
and U2566 (N_2566,N_1921,N_1880);
or U2567 (N_2567,N_1785,N_1716);
or U2568 (N_2568,N_1198,N_1211);
xor U2569 (N_2569,N_1568,N_1363);
nand U2570 (N_2570,N_1865,N_1840);
and U2571 (N_2571,N_1229,N_1802);
nand U2572 (N_2572,N_1133,N_1268);
and U2573 (N_2573,N_1150,N_1106);
xnor U2574 (N_2574,N_1792,N_1933);
nand U2575 (N_2575,N_1060,N_1666);
xor U2576 (N_2576,N_1559,N_1248);
or U2577 (N_2577,N_1150,N_1283);
and U2578 (N_2578,N_1156,N_1519);
and U2579 (N_2579,N_1582,N_1395);
nor U2580 (N_2580,N_1049,N_1653);
nor U2581 (N_2581,N_1846,N_1527);
and U2582 (N_2582,N_1256,N_1939);
and U2583 (N_2583,N_1111,N_1977);
or U2584 (N_2584,N_1147,N_1110);
or U2585 (N_2585,N_1122,N_1689);
nand U2586 (N_2586,N_1242,N_1672);
nand U2587 (N_2587,N_1071,N_1325);
xnor U2588 (N_2588,N_1921,N_1422);
nand U2589 (N_2589,N_1706,N_1256);
nor U2590 (N_2590,N_1928,N_1082);
or U2591 (N_2591,N_1324,N_1232);
or U2592 (N_2592,N_1870,N_1049);
or U2593 (N_2593,N_1881,N_1168);
and U2594 (N_2594,N_1454,N_1755);
xor U2595 (N_2595,N_1750,N_1710);
nor U2596 (N_2596,N_1449,N_1304);
xor U2597 (N_2597,N_1589,N_1717);
nand U2598 (N_2598,N_1127,N_1467);
xnor U2599 (N_2599,N_1172,N_1808);
or U2600 (N_2600,N_1742,N_1211);
or U2601 (N_2601,N_1455,N_1251);
xnor U2602 (N_2602,N_1300,N_1873);
nor U2603 (N_2603,N_1991,N_1362);
nor U2604 (N_2604,N_1506,N_1108);
nor U2605 (N_2605,N_1260,N_1825);
nor U2606 (N_2606,N_1610,N_1188);
and U2607 (N_2607,N_1252,N_1790);
nand U2608 (N_2608,N_1153,N_1605);
nand U2609 (N_2609,N_1885,N_1171);
or U2610 (N_2610,N_1857,N_1166);
nand U2611 (N_2611,N_1191,N_1092);
nand U2612 (N_2612,N_1531,N_1540);
nor U2613 (N_2613,N_1450,N_1777);
nor U2614 (N_2614,N_1345,N_1462);
nor U2615 (N_2615,N_1406,N_1210);
xnor U2616 (N_2616,N_1408,N_1592);
xor U2617 (N_2617,N_1892,N_1664);
and U2618 (N_2618,N_1641,N_1713);
xor U2619 (N_2619,N_1498,N_1334);
or U2620 (N_2620,N_1105,N_1027);
nor U2621 (N_2621,N_1478,N_1604);
xnor U2622 (N_2622,N_1357,N_1161);
nand U2623 (N_2623,N_1300,N_1393);
nand U2624 (N_2624,N_1343,N_1536);
nand U2625 (N_2625,N_1225,N_1743);
or U2626 (N_2626,N_1066,N_1227);
nand U2627 (N_2627,N_1193,N_1636);
nor U2628 (N_2628,N_1602,N_1606);
nand U2629 (N_2629,N_1111,N_1453);
or U2630 (N_2630,N_1676,N_1318);
and U2631 (N_2631,N_1186,N_1499);
nand U2632 (N_2632,N_1503,N_1713);
and U2633 (N_2633,N_1965,N_1082);
and U2634 (N_2634,N_1857,N_1012);
nor U2635 (N_2635,N_1110,N_1503);
or U2636 (N_2636,N_1119,N_1350);
xor U2637 (N_2637,N_1965,N_1020);
nor U2638 (N_2638,N_1192,N_1173);
xor U2639 (N_2639,N_1352,N_1896);
xor U2640 (N_2640,N_1484,N_1475);
nor U2641 (N_2641,N_1725,N_1741);
nor U2642 (N_2642,N_1042,N_1777);
nor U2643 (N_2643,N_1459,N_1395);
and U2644 (N_2644,N_1059,N_1542);
xor U2645 (N_2645,N_1928,N_1527);
nand U2646 (N_2646,N_1650,N_1746);
nand U2647 (N_2647,N_1938,N_1012);
or U2648 (N_2648,N_1687,N_1346);
nor U2649 (N_2649,N_1489,N_1195);
and U2650 (N_2650,N_1629,N_1460);
or U2651 (N_2651,N_1328,N_1042);
xnor U2652 (N_2652,N_1574,N_1579);
and U2653 (N_2653,N_1017,N_1916);
or U2654 (N_2654,N_1092,N_1962);
nor U2655 (N_2655,N_1492,N_1537);
nand U2656 (N_2656,N_1637,N_1147);
nor U2657 (N_2657,N_1505,N_1358);
or U2658 (N_2658,N_1485,N_1300);
nand U2659 (N_2659,N_1822,N_1254);
and U2660 (N_2660,N_1939,N_1691);
nor U2661 (N_2661,N_1850,N_1037);
or U2662 (N_2662,N_1263,N_1372);
and U2663 (N_2663,N_1090,N_1346);
xor U2664 (N_2664,N_1786,N_1550);
and U2665 (N_2665,N_1077,N_1592);
xor U2666 (N_2666,N_1784,N_1894);
nand U2667 (N_2667,N_1235,N_1482);
or U2668 (N_2668,N_1342,N_1249);
or U2669 (N_2669,N_1916,N_1127);
and U2670 (N_2670,N_1792,N_1652);
nand U2671 (N_2671,N_1700,N_1452);
and U2672 (N_2672,N_1778,N_1625);
nor U2673 (N_2673,N_1744,N_1742);
or U2674 (N_2674,N_1619,N_1725);
xor U2675 (N_2675,N_1037,N_1014);
nor U2676 (N_2676,N_1646,N_1787);
or U2677 (N_2677,N_1571,N_1545);
xnor U2678 (N_2678,N_1247,N_1877);
or U2679 (N_2679,N_1190,N_1229);
xor U2680 (N_2680,N_1999,N_1785);
or U2681 (N_2681,N_1570,N_1367);
and U2682 (N_2682,N_1585,N_1535);
xnor U2683 (N_2683,N_1174,N_1443);
and U2684 (N_2684,N_1600,N_1436);
and U2685 (N_2685,N_1209,N_1805);
and U2686 (N_2686,N_1031,N_1223);
nand U2687 (N_2687,N_1664,N_1350);
xor U2688 (N_2688,N_1545,N_1385);
nor U2689 (N_2689,N_1919,N_1413);
or U2690 (N_2690,N_1889,N_1308);
or U2691 (N_2691,N_1672,N_1055);
or U2692 (N_2692,N_1796,N_1271);
xor U2693 (N_2693,N_1874,N_1315);
and U2694 (N_2694,N_1549,N_1347);
or U2695 (N_2695,N_1440,N_1152);
and U2696 (N_2696,N_1131,N_1627);
nor U2697 (N_2697,N_1923,N_1682);
or U2698 (N_2698,N_1676,N_1190);
xnor U2699 (N_2699,N_1943,N_1929);
nor U2700 (N_2700,N_1081,N_1161);
and U2701 (N_2701,N_1125,N_1740);
xor U2702 (N_2702,N_1603,N_1438);
nor U2703 (N_2703,N_1944,N_1770);
xor U2704 (N_2704,N_1179,N_1811);
nand U2705 (N_2705,N_1812,N_1664);
nor U2706 (N_2706,N_1801,N_1277);
nand U2707 (N_2707,N_1398,N_1490);
or U2708 (N_2708,N_1850,N_1354);
and U2709 (N_2709,N_1172,N_1664);
nor U2710 (N_2710,N_1403,N_1887);
nor U2711 (N_2711,N_1748,N_1020);
nor U2712 (N_2712,N_1828,N_1605);
nor U2713 (N_2713,N_1478,N_1182);
xor U2714 (N_2714,N_1684,N_1947);
nor U2715 (N_2715,N_1727,N_1568);
nor U2716 (N_2716,N_1165,N_1629);
nor U2717 (N_2717,N_1932,N_1337);
nor U2718 (N_2718,N_1003,N_1656);
xor U2719 (N_2719,N_1279,N_1165);
and U2720 (N_2720,N_1709,N_1291);
and U2721 (N_2721,N_1466,N_1308);
nand U2722 (N_2722,N_1610,N_1974);
xnor U2723 (N_2723,N_1559,N_1159);
nor U2724 (N_2724,N_1959,N_1578);
nand U2725 (N_2725,N_1787,N_1582);
or U2726 (N_2726,N_1431,N_1773);
nand U2727 (N_2727,N_1967,N_1545);
nand U2728 (N_2728,N_1759,N_1277);
and U2729 (N_2729,N_1230,N_1123);
or U2730 (N_2730,N_1105,N_1118);
or U2731 (N_2731,N_1340,N_1388);
nor U2732 (N_2732,N_1438,N_1310);
xnor U2733 (N_2733,N_1702,N_1525);
or U2734 (N_2734,N_1508,N_1266);
or U2735 (N_2735,N_1593,N_1122);
nor U2736 (N_2736,N_1030,N_1855);
or U2737 (N_2737,N_1930,N_1612);
xnor U2738 (N_2738,N_1679,N_1542);
and U2739 (N_2739,N_1518,N_1563);
and U2740 (N_2740,N_1781,N_1711);
and U2741 (N_2741,N_1379,N_1850);
nand U2742 (N_2742,N_1816,N_1186);
nor U2743 (N_2743,N_1224,N_1726);
or U2744 (N_2744,N_1986,N_1870);
and U2745 (N_2745,N_1521,N_1676);
xor U2746 (N_2746,N_1524,N_1390);
and U2747 (N_2747,N_1228,N_1200);
nor U2748 (N_2748,N_1975,N_1180);
nor U2749 (N_2749,N_1383,N_1493);
xnor U2750 (N_2750,N_1777,N_1017);
xnor U2751 (N_2751,N_1056,N_1586);
and U2752 (N_2752,N_1794,N_1449);
nand U2753 (N_2753,N_1369,N_1409);
and U2754 (N_2754,N_1431,N_1785);
nor U2755 (N_2755,N_1965,N_1134);
or U2756 (N_2756,N_1845,N_1004);
and U2757 (N_2757,N_1897,N_1349);
xor U2758 (N_2758,N_1283,N_1205);
xor U2759 (N_2759,N_1384,N_1985);
nor U2760 (N_2760,N_1880,N_1489);
nor U2761 (N_2761,N_1585,N_1733);
nand U2762 (N_2762,N_1806,N_1787);
and U2763 (N_2763,N_1225,N_1064);
or U2764 (N_2764,N_1145,N_1858);
and U2765 (N_2765,N_1365,N_1440);
nand U2766 (N_2766,N_1105,N_1160);
xnor U2767 (N_2767,N_1466,N_1211);
xor U2768 (N_2768,N_1135,N_1867);
xor U2769 (N_2769,N_1397,N_1392);
xor U2770 (N_2770,N_1834,N_1800);
nand U2771 (N_2771,N_1317,N_1303);
xor U2772 (N_2772,N_1105,N_1515);
nor U2773 (N_2773,N_1363,N_1782);
nor U2774 (N_2774,N_1874,N_1167);
and U2775 (N_2775,N_1856,N_1604);
and U2776 (N_2776,N_1120,N_1975);
nor U2777 (N_2777,N_1087,N_1302);
and U2778 (N_2778,N_1515,N_1118);
nand U2779 (N_2779,N_1077,N_1600);
and U2780 (N_2780,N_1200,N_1271);
nor U2781 (N_2781,N_1709,N_1092);
or U2782 (N_2782,N_1285,N_1345);
and U2783 (N_2783,N_1829,N_1634);
nor U2784 (N_2784,N_1669,N_1921);
or U2785 (N_2785,N_1430,N_1260);
or U2786 (N_2786,N_1649,N_1518);
or U2787 (N_2787,N_1107,N_1923);
nor U2788 (N_2788,N_1776,N_1106);
and U2789 (N_2789,N_1639,N_1923);
xor U2790 (N_2790,N_1656,N_1445);
or U2791 (N_2791,N_1639,N_1864);
nand U2792 (N_2792,N_1596,N_1200);
nor U2793 (N_2793,N_1659,N_1445);
or U2794 (N_2794,N_1211,N_1706);
nand U2795 (N_2795,N_1440,N_1107);
xnor U2796 (N_2796,N_1627,N_1956);
and U2797 (N_2797,N_1237,N_1414);
nor U2798 (N_2798,N_1164,N_1155);
and U2799 (N_2799,N_1957,N_1732);
nand U2800 (N_2800,N_1101,N_1195);
and U2801 (N_2801,N_1163,N_1110);
nand U2802 (N_2802,N_1436,N_1871);
and U2803 (N_2803,N_1273,N_1611);
nor U2804 (N_2804,N_1484,N_1372);
xor U2805 (N_2805,N_1243,N_1026);
and U2806 (N_2806,N_1384,N_1930);
and U2807 (N_2807,N_1216,N_1995);
nor U2808 (N_2808,N_1305,N_1416);
nand U2809 (N_2809,N_1512,N_1126);
or U2810 (N_2810,N_1503,N_1909);
or U2811 (N_2811,N_1473,N_1373);
and U2812 (N_2812,N_1624,N_1854);
nand U2813 (N_2813,N_1039,N_1825);
and U2814 (N_2814,N_1647,N_1055);
nor U2815 (N_2815,N_1507,N_1114);
and U2816 (N_2816,N_1714,N_1700);
and U2817 (N_2817,N_1432,N_1663);
xnor U2818 (N_2818,N_1149,N_1758);
nand U2819 (N_2819,N_1036,N_1443);
nand U2820 (N_2820,N_1986,N_1726);
nor U2821 (N_2821,N_1790,N_1787);
and U2822 (N_2822,N_1148,N_1903);
xor U2823 (N_2823,N_1609,N_1759);
and U2824 (N_2824,N_1130,N_1409);
nor U2825 (N_2825,N_1648,N_1342);
and U2826 (N_2826,N_1526,N_1838);
xor U2827 (N_2827,N_1205,N_1016);
or U2828 (N_2828,N_1875,N_1649);
or U2829 (N_2829,N_1654,N_1100);
xnor U2830 (N_2830,N_1197,N_1216);
nor U2831 (N_2831,N_1663,N_1815);
or U2832 (N_2832,N_1670,N_1144);
xnor U2833 (N_2833,N_1751,N_1159);
nor U2834 (N_2834,N_1305,N_1016);
xor U2835 (N_2835,N_1963,N_1858);
nand U2836 (N_2836,N_1705,N_1270);
nand U2837 (N_2837,N_1605,N_1316);
nand U2838 (N_2838,N_1545,N_1092);
and U2839 (N_2839,N_1559,N_1166);
or U2840 (N_2840,N_1144,N_1201);
nand U2841 (N_2841,N_1421,N_1975);
and U2842 (N_2842,N_1936,N_1240);
xnor U2843 (N_2843,N_1126,N_1059);
nand U2844 (N_2844,N_1232,N_1661);
nor U2845 (N_2845,N_1857,N_1955);
and U2846 (N_2846,N_1780,N_1203);
nand U2847 (N_2847,N_1377,N_1476);
nor U2848 (N_2848,N_1502,N_1033);
and U2849 (N_2849,N_1424,N_1685);
xnor U2850 (N_2850,N_1329,N_1174);
and U2851 (N_2851,N_1184,N_1725);
or U2852 (N_2852,N_1969,N_1223);
xor U2853 (N_2853,N_1070,N_1671);
nand U2854 (N_2854,N_1410,N_1730);
and U2855 (N_2855,N_1920,N_1747);
xor U2856 (N_2856,N_1635,N_1657);
nor U2857 (N_2857,N_1112,N_1060);
nand U2858 (N_2858,N_1405,N_1345);
and U2859 (N_2859,N_1885,N_1853);
nand U2860 (N_2860,N_1032,N_1056);
nor U2861 (N_2861,N_1782,N_1676);
nand U2862 (N_2862,N_1300,N_1802);
nand U2863 (N_2863,N_1662,N_1533);
nand U2864 (N_2864,N_1108,N_1200);
or U2865 (N_2865,N_1542,N_1605);
and U2866 (N_2866,N_1395,N_1930);
nor U2867 (N_2867,N_1452,N_1333);
nand U2868 (N_2868,N_1052,N_1752);
and U2869 (N_2869,N_1582,N_1211);
nor U2870 (N_2870,N_1342,N_1425);
or U2871 (N_2871,N_1918,N_1007);
xor U2872 (N_2872,N_1360,N_1096);
nand U2873 (N_2873,N_1552,N_1832);
or U2874 (N_2874,N_1172,N_1379);
xor U2875 (N_2875,N_1480,N_1068);
nand U2876 (N_2876,N_1596,N_1475);
xor U2877 (N_2877,N_1724,N_1130);
nor U2878 (N_2878,N_1823,N_1577);
nand U2879 (N_2879,N_1794,N_1677);
nand U2880 (N_2880,N_1264,N_1494);
and U2881 (N_2881,N_1349,N_1979);
or U2882 (N_2882,N_1520,N_1376);
nor U2883 (N_2883,N_1069,N_1391);
or U2884 (N_2884,N_1048,N_1413);
or U2885 (N_2885,N_1146,N_1995);
and U2886 (N_2886,N_1655,N_1848);
nand U2887 (N_2887,N_1303,N_1725);
xor U2888 (N_2888,N_1153,N_1829);
or U2889 (N_2889,N_1141,N_1662);
and U2890 (N_2890,N_1395,N_1307);
and U2891 (N_2891,N_1202,N_1786);
nand U2892 (N_2892,N_1942,N_1227);
xnor U2893 (N_2893,N_1330,N_1540);
xor U2894 (N_2894,N_1634,N_1647);
nand U2895 (N_2895,N_1372,N_1974);
xnor U2896 (N_2896,N_1483,N_1240);
xor U2897 (N_2897,N_1050,N_1220);
xor U2898 (N_2898,N_1222,N_1119);
and U2899 (N_2899,N_1798,N_1885);
xor U2900 (N_2900,N_1449,N_1612);
and U2901 (N_2901,N_1199,N_1978);
and U2902 (N_2902,N_1741,N_1059);
nand U2903 (N_2903,N_1976,N_1981);
or U2904 (N_2904,N_1619,N_1128);
nand U2905 (N_2905,N_1209,N_1586);
nor U2906 (N_2906,N_1162,N_1005);
xor U2907 (N_2907,N_1020,N_1336);
nand U2908 (N_2908,N_1156,N_1478);
and U2909 (N_2909,N_1679,N_1345);
xnor U2910 (N_2910,N_1601,N_1687);
xnor U2911 (N_2911,N_1102,N_1429);
xnor U2912 (N_2912,N_1254,N_1761);
and U2913 (N_2913,N_1630,N_1564);
nor U2914 (N_2914,N_1221,N_1362);
or U2915 (N_2915,N_1116,N_1969);
and U2916 (N_2916,N_1342,N_1990);
nor U2917 (N_2917,N_1648,N_1303);
or U2918 (N_2918,N_1213,N_1752);
xor U2919 (N_2919,N_1618,N_1072);
and U2920 (N_2920,N_1229,N_1230);
and U2921 (N_2921,N_1012,N_1218);
xnor U2922 (N_2922,N_1509,N_1547);
and U2923 (N_2923,N_1845,N_1107);
nand U2924 (N_2924,N_1500,N_1809);
nor U2925 (N_2925,N_1568,N_1551);
and U2926 (N_2926,N_1979,N_1379);
xnor U2927 (N_2927,N_1890,N_1884);
and U2928 (N_2928,N_1599,N_1715);
xor U2929 (N_2929,N_1200,N_1972);
or U2930 (N_2930,N_1420,N_1678);
and U2931 (N_2931,N_1474,N_1072);
xor U2932 (N_2932,N_1829,N_1735);
nor U2933 (N_2933,N_1331,N_1232);
xor U2934 (N_2934,N_1358,N_1838);
xor U2935 (N_2935,N_1355,N_1434);
nand U2936 (N_2936,N_1803,N_1830);
nor U2937 (N_2937,N_1635,N_1289);
and U2938 (N_2938,N_1203,N_1319);
nand U2939 (N_2939,N_1681,N_1799);
or U2940 (N_2940,N_1847,N_1960);
nand U2941 (N_2941,N_1624,N_1107);
nor U2942 (N_2942,N_1879,N_1776);
xor U2943 (N_2943,N_1223,N_1711);
nand U2944 (N_2944,N_1043,N_1772);
xor U2945 (N_2945,N_1088,N_1831);
or U2946 (N_2946,N_1135,N_1369);
and U2947 (N_2947,N_1155,N_1478);
xor U2948 (N_2948,N_1324,N_1532);
nor U2949 (N_2949,N_1007,N_1102);
nor U2950 (N_2950,N_1980,N_1343);
nand U2951 (N_2951,N_1075,N_1694);
nor U2952 (N_2952,N_1482,N_1633);
and U2953 (N_2953,N_1089,N_1248);
xor U2954 (N_2954,N_1677,N_1232);
nor U2955 (N_2955,N_1928,N_1261);
or U2956 (N_2956,N_1464,N_1820);
nand U2957 (N_2957,N_1217,N_1720);
xnor U2958 (N_2958,N_1555,N_1958);
nand U2959 (N_2959,N_1124,N_1829);
or U2960 (N_2960,N_1031,N_1706);
xor U2961 (N_2961,N_1806,N_1895);
nand U2962 (N_2962,N_1172,N_1761);
and U2963 (N_2963,N_1764,N_1518);
or U2964 (N_2964,N_1701,N_1772);
nor U2965 (N_2965,N_1899,N_1414);
and U2966 (N_2966,N_1850,N_1980);
nor U2967 (N_2967,N_1481,N_1676);
xnor U2968 (N_2968,N_1373,N_1241);
or U2969 (N_2969,N_1365,N_1482);
or U2970 (N_2970,N_1159,N_1088);
and U2971 (N_2971,N_1101,N_1100);
and U2972 (N_2972,N_1560,N_1472);
nand U2973 (N_2973,N_1537,N_1632);
and U2974 (N_2974,N_1267,N_1853);
and U2975 (N_2975,N_1382,N_1969);
or U2976 (N_2976,N_1897,N_1506);
nand U2977 (N_2977,N_1370,N_1453);
and U2978 (N_2978,N_1939,N_1353);
or U2979 (N_2979,N_1109,N_1387);
or U2980 (N_2980,N_1509,N_1217);
and U2981 (N_2981,N_1734,N_1038);
nor U2982 (N_2982,N_1840,N_1942);
or U2983 (N_2983,N_1743,N_1152);
or U2984 (N_2984,N_1730,N_1141);
nand U2985 (N_2985,N_1172,N_1120);
nand U2986 (N_2986,N_1669,N_1879);
xor U2987 (N_2987,N_1808,N_1857);
and U2988 (N_2988,N_1429,N_1504);
nor U2989 (N_2989,N_1549,N_1787);
and U2990 (N_2990,N_1343,N_1929);
nand U2991 (N_2991,N_1870,N_1582);
nand U2992 (N_2992,N_1405,N_1197);
nor U2993 (N_2993,N_1539,N_1707);
and U2994 (N_2994,N_1777,N_1696);
nand U2995 (N_2995,N_1207,N_1810);
nor U2996 (N_2996,N_1022,N_1545);
nor U2997 (N_2997,N_1807,N_1982);
xor U2998 (N_2998,N_1869,N_1411);
nor U2999 (N_2999,N_1684,N_1145);
xor U3000 (N_3000,N_2089,N_2717);
or U3001 (N_3001,N_2714,N_2385);
or U3002 (N_3002,N_2427,N_2775);
and U3003 (N_3003,N_2210,N_2457);
and U3004 (N_3004,N_2045,N_2090);
or U3005 (N_3005,N_2443,N_2500);
and U3006 (N_3006,N_2477,N_2339);
xor U3007 (N_3007,N_2699,N_2223);
nor U3008 (N_3008,N_2792,N_2613);
xor U3009 (N_3009,N_2200,N_2087);
or U3010 (N_3010,N_2373,N_2050);
or U3011 (N_3011,N_2317,N_2883);
and U3012 (N_3012,N_2582,N_2215);
xnor U3013 (N_3013,N_2820,N_2763);
xor U3014 (N_3014,N_2845,N_2399);
nor U3015 (N_3015,N_2201,N_2587);
or U3016 (N_3016,N_2798,N_2003);
nor U3017 (N_3017,N_2534,N_2861);
nand U3018 (N_3018,N_2429,N_2138);
nor U3019 (N_3019,N_2451,N_2124);
and U3020 (N_3020,N_2590,N_2471);
and U3021 (N_3021,N_2463,N_2430);
nand U3022 (N_3022,N_2646,N_2356);
xnor U3023 (N_3023,N_2411,N_2418);
nor U3024 (N_3024,N_2135,N_2364);
and U3025 (N_3025,N_2764,N_2868);
nand U3026 (N_3026,N_2597,N_2194);
nor U3027 (N_3027,N_2610,N_2348);
nor U3028 (N_3028,N_2809,N_2494);
xnor U3029 (N_3029,N_2272,N_2332);
nand U3030 (N_3030,N_2746,N_2234);
and U3031 (N_3031,N_2287,N_2986);
nor U3032 (N_3032,N_2640,N_2540);
nor U3033 (N_3033,N_2663,N_2833);
nand U3034 (N_3034,N_2203,N_2366);
nor U3035 (N_3035,N_2354,N_2721);
nor U3036 (N_3036,N_2572,N_2831);
or U3037 (N_3037,N_2658,N_2057);
xnor U3038 (N_3038,N_2678,N_2467);
xnor U3039 (N_3039,N_2794,N_2550);
and U3040 (N_3040,N_2612,N_2183);
nand U3041 (N_3041,N_2144,N_2335);
nor U3042 (N_3042,N_2675,N_2805);
nand U3043 (N_3043,N_2859,N_2575);
or U3044 (N_3044,N_2837,N_2732);
and U3045 (N_3045,N_2823,N_2172);
or U3046 (N_3046,N_2964,N_2403);
and U3047 (N_3047,N_2759,N_2727);
or U3048 (N_3048,N_2322,N_2639);
xor U3049 (N_3049,N_2110,N_2495);
nand U3050 (N_3050,N_2803,N_2520);
or U3051 (N_3051,N_2382,N_2815);
nor U3052 (N_3052,N_2072,N_2434);
xnor U3053 (N_3053,N_2718,N_2188);
xor U3054 (N_3054,N_2175,N_2513);
xnor U3055 (N_3055,N_2554,N_2931);
or U3056 (N_3056,N_2576,N_2093);
nand U3057 (N_3057,N_2165,N_2244);
nand U3058 (N_3058,N_2836,N_2959);
nand U3059 (N_3059,N_2415,N_2114);
xnor U3060 (N_3060,N_2005,N_2207);
nand U3061 (N_3061,N_2168,N_2092);
and U3062 (N_3062,N_2445,N_2543);
and U3063 (N_3063,N_2942,N_2464);
or U3064 (N_3064,N_2519,N_2261);
and U3065 (N_3065,N_2478,N_2007);
nor U3066 (N_3066,N_2967,N_2325);
xor U3067 (N_3067,N_2459,N_2224);
xnor U3068 (N_3068,N_2885,N_2148);
nor U3069 (N_3069,N_2954,N_2031);
xnor U3070 (N_3070,N_2561,N_2372);
or U3071 (N_3071,N_2601,N_2706);
xor U3072 (N_3072,N_2008,N_2501);
and U3073 (N_3073,N_2822,N_2414);
xnor U3074 (N_3074,N_2752,N_2762);
xor U3075 (N_3075,N_2992,N_2687);
xor U3076 (N_3076,N_2644,N_2424);
nand U3077 (N_3077,N_2566,N_2568);
or U3078 (N_3078,N_2839,N_2055);
nand U3079 (N_3079,N_2344,N_2474);
nand U3080 (N_3080,N_2531,N_2692);
or U3081 (N_3081,N_2696,N_2070);
nor U3082 (N_3082,N_2104,N_2130);
nand U3083 (N_3083,N_2788,N_2630);
xnor U3084 (N_3084,N_2901,N_2405);
xor U3085 (N_3085,N_2258,N_2648);
nor U3086 (N_3086,N_2169,N_2064);
nand U3087 (N_3087,N_2984,N_2028);
or U3088 (N_3088,N_2857,N_2862);
or U3089 (N_3089,N_2659,N_2041);
or U3090 (N_3090,N_2591,N_2637);
xnor U3091 (N_3091,N_2012,N_2231);
nor U3092 (N_3092,N_2671,N_2357);
nor U3093 (N_3093,N_2375,N_2480);
nand U3094 (N_3094,N_2017,N_2108);
or U3095 (N_3095,N_2510,N_2131);
nor U3096 (N_3096,N_2290,N_2420);
nand U3097 (N_3097,N_2448,N_2879);
xnor U3098 (N_3098,N_2206,N_2466);
and U3099 (N_3099,N_2887,N_2054);
or U3100 (N_3100,N_2748,N_2359);
nand U3101 (N_3101,N_2565,N_2182);
xnor U3102 (N_3102,N_2940,N_2626);
nor U3103 (N_3103,N_2624,N_2245);
or U3104 (N_3104,N_2199,N_2807);
or U3105 (N_3105,N_2437,N_2242);
xor U3106 (N_3106,N_2402,N_2300);
xor U3107 (N_3107,N_2091,N_2856);
nor U3108 (N_3108,N_2677,N_2056);
or U3109 (N_3109,N_2975,N_2846);
or U3110 (N_3110,N_2256,N_2584);
xnor U3111 (N_3111,N_2878,N_2826);
nand U3112 (N_3112,N_2749,N_2275);
xnor U3113 (N_3113,N_2532,N_2835);
xnor U3114 (N_3114,N_2653,N_2324);
nand U3115 (N_3115,N_2974,N_2439);
or U3116 (N_3116,N_2378,N_2787);
or U3117 (N_3117,N_2512,N_2269);
nand U3118 (N_3118,N_2524,N_2758);
nor U3119 (N_3119,N_2395,N_2580);
and U3120 (N_3120,N_2113,N_2617);
and U3121 (N_3121,N_2987,N_2795);
nor U3122 (N_3122,N_2574,N_2609);
nor U3123 (N_3123,N_2923,N_2834);
xor U3124 (N_3124,N_2810,N_2485);
nor U3125 (N_3125,N_2782,N_2517);
and U3126 (N_3126,N_2394,N_2979);
or U3127 (N_3127,N_2010,N_2783);
or U3128 (N_3128,N_2042,N_2944);
xnor U3129 (N_3129,N_2547,N_2178);
and U3130 (N_3130,N_2291,N_2652);
nor U3131 (N_3131,N_2698,N_2682);
nand U3132 (N_3132,N_2129,N_2595);
and U3133 (N_3133,N_2526,N_2119);
nand U3134 (N_3134,N_2600,N_2268);
nor U3135 (N_3135,N_2473,N_2305);
nor U3136 (N_3136,N_2904,N_2655);
nor U3137 (N_3137,N_2848,N_2981);
nor U3138 (N_3138,N_2622,N_2053);
or U3139 (N_3139,N_2537,N_2674);
xor U3140 (N_3140,N_2440,N_2909);
xnor U3141 (N_3141,N_2867,N_2033);
nor U3142 (N_3142,N_2662,N_2875);
or U3143 (N_3143,N_2755,N_2292);
or U3144 (N_3144,N_2401,N_2866);
or U3145 (N_3145,N_2422,N_2498);
or U3146 (N_3146,N_2227,N_2946);
or U3147 (N_3147,N_2035,N_2465);
nand U3148 (N_3148,N_2232,N_2611);
nand U3149 (N_3149,N_2202,N_2340);
nand U3150 (N_3150,N_2396,N_2013);
and U3151 (N_3151,N_2970,N_2253);
or U3152 (N_3152,N_2529,N_2850);
and U3153 (N_3153,N_2281,N_2163);
or U3154 (N_3154,N_2707,N_2898);
and U3155 (N_3155,N_2973,N_2585);
xor U3156 (N_3156,N_2143,N_2725);
or U3157 (N_3157,N_2939,N_2254);
nor U3158 (N_3158,N_2355,N_2829);
or U3159 (N_3159,N_2100,N_2358);
nor U3160 (N_3160,N_2177,N_2908);
or U3161 (N_3161,N_2799,N_2160);
nand U3162 (N_3162,N_2661,N_2802);
xor U3163 (N_3163,N_2599,N_2628);
or U3164 (N_3164,N_2925,N_2404);
nand U3165 (N_3165,N_2497,N_2535);
xor U3166 (N_3166,N_2078,N_2766);
and U3167 (N_3167,N_2669,N_2650);
nand U3168 (N_3168,N_2487,N_2625);
nand U3169 (N_3169,N_2051,N_2681);
nand U3170 (N_3170,N_2556,N_2059);
nor U3171 (N_3171,N_2731,N_2184);
and U3172 (N_3172,N_2685,N_2310);
nand U3173 (N_3173,N_2225,N_2869);
or U3174 (N_3174,N_2744,N_2907);
or U3175 (N_3175,N_2690,N_2142);
xor U3176 (N_3176,N_2779,N_2761);
nand U3177 (N_3177,N_2813,N_2990);
nor U3178 (N_3178,N_2309,N_2488);
nor U3179 (N_3179,N_2294,N_2623);
and U3180 (N_3180,N_2694,N_2251);
nor U3181 (N_3181,N_2496,N_2873);
xor U3182 (N_3182,N_2830,N_2539);
xnor U3183 (N_3183,N_2930,N_2980);
or U3184 (N_3184,N_2924,N_2740);
nand U3185 (N_3185,N_2765,N_2276);
xor U3186 (N_3186,N_2299,N_2511);
nand U3187 (N_3187,N_2757,N_2971);
nor U3188 (N_3188,N_2893,N_2304);
nor U3189 (N_3189,N_2107,N_2470);
nand U3190 (N_3190,N_2703,N_2337);
or U3191 (N_3191,N_2506,N_2238);
nor U3192 (N_3192,N_2935,N_2071);
nand U3193 (N_3193,N_2193,N_2282);
or U3194 (N_3194,N_2191,N_2111);
nor U3195 (N_3195,N_2295,N_2683);
or U3196 (N_3196,N_2088,N_2011);
and U3197 (N_3197,N_2320,N_2502);
and U3198 (N_3198,N_2336,N_2548);
or U3199 (N_3199,N_2865,N_2001);
nor U3200 (N_3200,N_2647,N_2277);
and U3201 (N_3201,N_2842,N_2505);
nor U3202 (N_3202,N_2314,N_2376);
and U3203 (N_3203,N_2558,N_2723);
nand U3204 (N_3204,N_2492,N_2343);
nor U3205 (N_3205,N_2438,N_2997);
xor U3206 (N_3206,N_2751,N_2668);
and U3207 (N_3207,N_2614,N_2009);
and U3208 (N_3208,N_2265,N_2419);
xor U3209 (N_3209,N_2928,N_2567);
or U3210 (N_3210,N_2918,N_2433);
nor U3211 (N_3211,N_2243,N_2863);
and U3212 (N_3212,N_2722,N_2503);
or U3213 (N_3213,N_2363,N_2991);
and U3214 (N_3214,N_2458,N_2158);
or U3215 (N_3215,N_2298,N_2933);
and U3216 (N_3216,N_2047,N_2937);
nor U3217 (N_3217,N_2881,N_2577);
or U3218 (N_3218,N_2280,N_2482);
or U3219 (N_3219,N_2914,N_2629);
or U3220 (N_3220,N_2246,N_2832);
and U3221 (N_3221,N_2573,N_2593);
xnor U3222 (N_3222,N_2793,N_2077);
nor U3223 (N_3223,N_2801,N_2950);
nand U3224 (N_3224,N_2545,N_2136);
and U3225 (N_3225,N_2301,N_2365);
xor U3226 (N_3226,N_2296,N_2538);
nor U3227 (N_3227,N_2735,N_2333);
xor U3228 (N_3228,N_2384,N_2563);
or U3229 (N_3229,N_2934,N_2627);
nor U3230 (N_3230,N_2407,N_2767);
or U3231 (N_3231,N_2122,N_2369);
nor U3232 (N_3232,N_2578,N_2679);
nor U3233 (N_3233,N_2774,N_2999);
nand U3234 (N_3234,N_2481,N_2781);
or U3235 (N_3235,N_2890,N_2938);
nor U3236 (N_3236,N_2034,N_2441);
xnor U3237 (N_3237,N_2386,N_2150);
xnor U3238 (N_3238,N_2274,N_2022);
xnor U3239 (N_3239,N_2527,N_2444);
or U3240 (N_3240,N_2398,N_2204);
and U3241 (N_3241,N_2360,N_2888);
or U3242 (N_3242,N_2307,N_2852);
nor U3243 (N_3243,N_2021,N_2476);
nor U3244 (N_3244,N_2800,N_2509);
xor U3245 (N_3245,N_2818,N_2952);
nand U3246 (N_3246,N_2770,N_2943);
or U3247 (N_3247,N_2239,N_2279);
xor U3248 (N_3248,N_2213,N_2469);
nor U3249 (N_3249,N_2579,N_2331);
and U3250 (N_3250,N_2367,N_2541);
nor U3251 (N_3251,N_2821,N_2564);
nand U3252 (N_3252,N_2927,N_2976);
and U3253 (N_3253,N_2133,N_2039);
or U3254 (N_3254,N_2392,N_2745);
and U3255 (N_3255,N_2515,N_2174);
nor U3256 (N_3256,N_2328,N_2214);
nor U3257 (N_3257,N_2374,N_2341);
nand U3258 (N_3258,N_2116,N_2004);
xor U3259 (N_3259,N_2257,N_2190);
nand U3260 (N_3260,N_2096,N_2780);
nor U3261 (N_3261,N_2146,N_2075);
and U3262 (N_3262,N_2977,N_2302);
or U3263 (N_3263,N_2181,N_2417);
or U3264 (N_3264,N_2285,N_2472);
or U3265 (N_3265,N_2874,N_2326);
and U3266 (N_3266,N_2052,N_2049);
nor U3267 (N_3267,N_2286,N_2642);
nand U3268 (N_3268,N_2393,N_2080);
xor U3269 (N_3269,N_2120,N_2843);
nor U3270 (N_3270,N_2858,N_2817);
nand U3271 (N_3271,N_2955,N_2633);
and U3272 (N_3272,N_2043,N_2283);
or U3273 (N_3273,N_2270,N_2894);
nor U3274 (N_3274,N_2902,N_2903);
xor U3275 (N_3275,N_2379,N_2074);
xnor U3276 (N_3276,N_2046,N_2164);
or U3277 (N_3277,N_2560,N_2263);
xnor U3278 (N_3278,N_2103,N_2230);
or U3279 (N_3279,N_2872,N_2618);
nor U3280 (N_3280,N_2040,N_2828);
or U3281 (N_3281,N_2330,N_2149);
nor U3282 (N_3282,N_2730,N_2919);
and U3283 (N_3283,N_2086,N_2994);
or U3284 (N_3284,N_2468,N_2185);
or U3285 (N_3285,N_2187,N_2708);
xnor U3286 (N_3286,N_2804,N_2099);
or U3287 (N_3287,N_2029,N_2020);
and U3288 (N_3288,N_2460,N_2596);
nand U3289 (N_3289,N_2691,N_2284);
nand U3290 (N_3290,N_2886,N_2953);
and U3291 (N_3291,N_2428,N_2037);
nor U3292 (N_3292,N_2777,N_2176);
nand U3293 (N_3293,N_2651,N_2095);
nand U3294 (N_3294,N_2643,N_2205);
nand U3295 (N_3295,N_2569,N_2173);
nor U3296 (N_3296,N_2453,N_2729);
nand U3297 (N_3297,N_2186,N_2588);
nand U3298 (N_3298,N_2312,N_2266);
nand U3299 (N_3299,N_2381,N_2211);
or U3300 (N_3300,N_2380,N_2670);
and U3301 (N_3301,N_2347,N_2018);
nor U3302 (N_3302,N_2109,N_2413);
and U3303 (N_3303,N_2960,N_2297);
nand U3304 (N_3304,N_2208,N_2880);
nand U3305 (N_3305,N_2737,N_2657);
nand U3306 (N_3306,N_2068,N_2084);
nand U3307 (N_3307,N_2079,N_2406);
nand U3308 (N_3308,N_2808,N_2447);
nand U3309 (N_3309,N_2267,N_2948);
and U3310 (N_3310,N_2308,N_2956);
and U3311 (N_3311,N_2702,N_2240);
nand U3312 (N_3312,N_2278,N_2860);
nor U3313 (N_3313,N_2978,N_2226);
and U3314 (N_3314,N_2704,N_2542);
and U3315 (N_3315,N_2006,N_2222);
nand U3316 (N_3316,N_2252,N_2137);
nor U3317 (N_3317,N_2559,N_2313);
nand U3318 (N_3318,N_2026,N_2897);
nand U3319 (N_3319,N_2998,N_2570);
nor U3320 (N_3320,N_2212,N_2016);
nand U3321 (N_3321,N_2772,N_2504);
and U3322 (N_3322,N_2632,N_2634);
xnor U3323 (N_3323,N_2705,N_2776);
and U3324 (N_3324,N_2361,N_2132);
or U3325 (N_3325,N_2048,N_2645);
or U3326 (N_3326,N_2724,N_2989);
nor U3327 (N_3327,N_2715,N_2736);
nor U3328 (N_3328,N_2423,N_2156);
or U3329 (N_3329,N_2557,N_2958);
nand U3330 (N_3330,N_2949,N_2247);
xor U3331 (N_3331,N_2889,N_2323);
and U3332 (N_3332,N_2123,N_2786);
and U3333 (N_3333,N_2790,N_2841);
xor U3334 (N_3334,N_2032,N_2228);
nand U3335 (N_3335,N_2877,N_2066);
nand U3336 (N_3336,N_2362,N_2237);
or U3337 (N_3337,N_2260,N_2273);
or U3338 (N_3338,N_2604,N_2271);
and U3339 (N_3339,N_2676,N_2117);
nor U3340 (N_3340,N_2598,N_2025);
xor U3341 (N_3341,N_2996,N_2913);
and U3342 (N_3342,N_2377,N_2638);
nand U3343 (N_3343,N_2002,N_2734);
and U3344 (N_3344,N_2030,N_2063);
or U3345 (N_3345,N_2432,N_2219);
nor U3346 (N_3346,N_2549,N_2555);
nand U3347 (N_3347,N_2391,N_2015);
nand U3348 (N_3348,N_2452,N_2824);
xor U3349 (N_3349,N_2983,N_2179);
nand U3350 (N_3350,N_2825,N_2666);
or U3351 (N_3351,N_2912,N_2533);
xor U3352 (N_3352,N_2636,N_2484);
xor U3353 (N_3353,N_2947,N_2462);
nand U3354 (N_3354,N_2155,N_2667);
nand U3355 (N_3355,N_2499,N_2988);
or U3356 (N_3356,N_2660,N_2289);
or U3357 (N_3357,N_2058,N_2608);
nand U3358 (N_3358,N_2241,N_2789);
nand U3359 (N_3359,N_2654,N_2311);
xor U3360 (N_3360,N_2083,N_2993);
nor U3361 (N_3361,N_2014,N_2635);
nor U3362 (N_3362,N_2450,N_2941);
xor U3363 (N_3363,N_2785,N_2665);
and U3364 (N_3364,N_2250,N_2491);
nand U3365 (N_3365,N_2768,N_2797);
nand U3366 (N_3366,N_2303,N_2159);
and U3367 (N_3367,N_2589,N_2552);
nor U3368 (N_3368,N_2603,N_2456);
nand U3369 (N_3369,N_2921,N_2383);
or U3370 (N_3370,N_2262,N_2352);
nand U3371 (N_3371,N_2838,N_2097);
nor U3372 (N_3372,N_2019,N_2726);
nand U3373 (N_3373,N_2605,N_2689);
nor U3374 (N_3374,N_2038,N_2806);
and U3375 (N_3375,N_2747,N_2400);
or U3376 (N_3376,N_2220,N_2709);
nor U3377 (N_3377,N_2695,N_2743);
xor U3378 (N_3378,N_2085,N_2412);
nand U3379 (N_3379,N_2189,N_2416);
nand U3380 (N_3380,N_2700,N_2528);
xnor U3381 (N_3381,N_2397,N_2170);
nor U3382 (N_3382,N_2854,N_2969);
xnor U3383 (N_3383,N_2390,N_2508);
nand U3384 (N_3384,N_2641,N_2876);
nand U3385 (N_3385,N_2963,N_2082);
and U3386 (N_3386,N_2895,N_2951);
nand U3387 (N_3387,N_2916,N_2192);
and U3388 (N_3388,N_2346,N_2141);
or U3389 (N_3389,N_2139,N_2784);
or U3390 (N_3390,N_2410,N_2349);
xnor U3391 (N_3391,N_2891,N_2522);
nor U3392 (N_3392,N_2446,N_2140);
xnor U3393 (N_3393,N_2811,N_2076);
and U3394 (N_3394,N_2607,N_2306);
nor U3395 (N_3395,N_2435,N_2711);
or U3396 (N_3396,N_2371,N_2686);
nand U3397 (N_3397,N_2932,N_2154);
and U3398 (N_3398,N_2870,N_2945);
xnor U3399 (N_3399,N_2882,N_2844);
nand U3400 (N_3400,N_2728,N_2000);
or U3401 (N_3401,N_2514,N_2530);
or U3402 (N_3402,N_2065,N_2115);
xnor U3403 (N_3403,N_2094,N_2490);
or U3404 (N_3404,N_2216,N_2905);
xnor U3405 (N_3405,N_2370,N_2812);
or U3406 (N_3406,N_2507,N_2345);
nor U3407 (N_3407,N_2024,N_2733);
and U3408 (N_3408,N_2217,N_2684);
or U3409 (N_3409,N_2738,N_2153);
xnor U3410 (N_3410,N_2796,N_2917);
nand U3411 (N_3411,N_2121,N_2483);
and U3412 (N_3412,N_2536,N_2926);
and U3413 (N_3413,N_2760,N_2493);
or U3414 (N_3414,N_2697,N_2544);
xor U3415 (N_3415,N_2649,N_2553);
and U3416 (N_3416,N_2819,N_2368);
or U3417 (N_3417,N_2965,N_2264);
or U3418 (N_3418,N_2847,N_2118);
xor U3419 (N_3419,N_2221,N_2334);
nand U3420 (N_3420,N_2426,N_2218);
or U3421 (N_3421,N_2036,N_2342);
or U3422 (N_3422,N_2387,N_2957);
and U3423 (N_3423,N_2518,N_2920);
or U3424 (N_3424,N_2060,N_2995);
nand U3425 (N_3425,N_2739,N_2102);
nand U3426 (N_3426,N_2840,N_2105);
xor U3427 (N_3427,N_2892,N_2713);
and U3428 (N_3428,N_2409,N_2816);
nor U3429 (N_3429,N_2672,N_2769);
xnor U3430 (N_3430,N_2936,N_2849);
xor U3431 (N_3431,N_2023,N_2436);
and U3432 (N_3432,N_2329,N_2408);
and U3433 (N_3433,N_2151,N_2853);
nand U3434 (N_3434,N_2209,N_2899);
and U3435 (N_3435,N_2710,N_2656);
or U3436 (N_3436,N_2197,N_2198);
nand U3437 (N_3437,N_2098,N_2754);
nor U3438 (N_3438,N_2318,N_2293);
xnor U3439 (N_3439,N_2615,N_2425);
xnor U3440 (N_3440,N_2061,N_2106);
nor U3441 (N_3441,N_2044,N_2431);
or U3442 (N_3442,N_2259,N_2719);
nor U3443 (N_3443,N_2851,N_2756);
or U3444 (N_3444,N_2127,N_2606);
nand U3445 (N_3445,N_2389,N_2753);
and U3446 (N_3446,N_2350,N_2195);
nor U3447 (N_3447,N_2982,N_2961);
nor U3448 (N_3448,N_2516,N_2562);
or U3449 (N_3449,N_2388,N_2966);
or U3450 (N_3450,N_2855,N_2884);
or U3451 (N_3451,N_2631,N_2248);
or U3452 (N_3452,N_2315,N_2985);
nand U3453 (N_3453,N_2621,N_2338);
and U3454 (N_3454,N_2929,N_2166);
nor U3455 (N_3455,N_2814,N_2062);
or U3456 (N_3456,N_2571,N_2479);
nor U3457 (N_3457,N_2664,N_2680);
nand U3458 (N_3458,N_2081,N_2586);
and U3459 (N_3459,N_2619,N_2475);
xor U3460 (N_3460,N_2972,N_2128);
nor U3461 (N_3461,N_2720,N_2791);
or U3462 (N_3462,N_2742,N_2180);
nand U3463 (N_3463,N_2910,N_2351);
or U3464 (N_3464,N_2771,N_2449);
and U3465 (N_3465,N_2229,N_2126);
and U3466 (N_3466,N_2523,N_2171);
xor U3467 (N_3467,N_2288,N_2145);
or U3468 (N_3468,N_2069,N_2233);
nand U3469 (N_3469,N_2461,N_2125);
xor U3470 (N_3470,N_2255,N_2249);
xor U3471 (N_3471,N_2442,N_2602);
nor U3472 (N_3472,N_2906,N_2773);
and U3473 (N_3473,N_2152,N_2067);
nor U3474 (N_3474,N_2693,N_2962);
nand U3475 (N_3475,N_2489,N_2196);
and U3476 (N_3476,N_2147,N_2896);
nand U3477 (N_3477,N_2101,N_2353);
nor U3478 (N_3478,N_2594,N_2620);
nor U3479 (N_3479,N_2716,N_2688);
or U3480 (N_3480,N_2592,N_2581);
nand U3481 (N_3481,N_2167,N_2546);
and U3482 (N_3482,N_2827,N_2922);
nor U3483 (N_3483,N_2236,N_2316);
or U3484 (N_3484,N_2235,N_2525);
xnor U3485 (N_3485,N_2321,N_2701);
and U3486 (N_3486,N_2112,N_2162);
or U3487 (N_3487,N_2455,N_2421);
or U3488 (N_3488,N_2551,N_2134);
nand U3489 (N_3489,N_2027,N_2900);
nand U3490 (N_3490,N_2157,N_2871);
nor U3491 (N_3491,N_2741,N_2968);
xor U3492 (N_3492,N_2319,N_2454);
and U3493 (N_3493,N_2161,N_2911);
nor U3494 (N_3494,N_2521,N_2583);
and U3495 (N_3495,N_2673,N_2486);
xor U3496 (N_3496,N_2915,N_2073);
nand U3497 (N_3497,N_2712,N_2616);
nor U3498 (N_3498,N_2864,N_2750);
and U3499 (N_3499,N_2778,N_2327);
and U3500 (N_3500,N_2935,N_2142);
xor U3501 (N_3501,N_2212,N_2471);
and U3502 (N_3502,N_2816,N_2564);
nand U3503 (N_3503,N_2316,N_2392);
xor U3504 (N_3504,N_2748,N_2205);
and U3505 (N_3505,N_2028,N_2786);
and U3506 (N_3506,N_2740,N_2539);
xor U3507 (N_3507,N_2754,N_2006);
xor U3508 (N_3508,N_2197,N_2037);
xor U3509 (N_3509,N_2729,N_2210);
nand U3510 (N_3510,N_2991,N_2251);
or U3511 (N_3511,N_2715,N_2198);
xor U3512 (N_3512,N_2962,N_2040);
nor U3513 (N_3513,N_2797,N_2043);
or U3514 (N_3514,N_2876,N_2415);
or U3515 (N_3515,N_2012,N_2228);
and U3516 (N_3516,N_2556,N_2755);
or U3517 (N_3517,N_2713,N_2840);
and U3518 (N_3518,N_2211,N_2589);
nor U3519 (N_3519,N_2249,N_2706);
and U3520 (N_3520,N_2263,N_2418);
and U3521 (N_3521,N_2169,N_2104);
nor U3522 (N_3522,N_2150,N_2195);
nand U3523 (N_3523,N_2550,N_2687);
xor U3524 (N_3524,N_2894,N_2786);
nand U3525 (N_3525,N_2319,N_2020);
xnor U3526 (N_3526,N_2142,N_2027);
nand U3527 (N_3527,N_2551,N_2003);
nand U3528 (N_3528,N_2172,N_2003);
or U3529 (N_3529,N_2294,N_2245);
nand U3530 (N_3530,N_2070,N_2447);
nor U3531 (N_3531,N_2940,N_2090);
nor U3532 (N_3532,N_2791,N_2033);
and U3533 (N_3533,N_2990,N_2022);
xnor U3534 (N_3534,N_2778,N_2344);
and U3535 (N_3535,N_2038,N_2489);
or U3536 (N_3536,N_2191,N_2511);
nand U3537 (N_3537,N_2248,N_2359);
xor U3538 (N_3538,N_2015,N_2251);
nor U3539 (N_3539,N_2203,N_2356);
xnor U3540 (N_3540,N_2734,N_2870);
or U3541 (N_3541,N_2372,N_2335);
nor U3542 (N_3542,N_2887,N_2925);
nor U3543 (N_3543,N_2489,N_2965);
or U3544 (N_3544,N_2970,N_2794);
xnor U3545 (N_3545,N_2425,N_2704);
xnor U3546 (N_3546,N_2386,N_2131);
or U3547 (N_3547,N_2430,N_2119);
nand U3548 (N_3548,N_2496,N_2838);
or U3549 (N_3549,N_2878,N_2300);
and U3550 (N_3550,N_2024,N_2687);
nand U3551 (N_3551,N_2794,N_2127);
nand U3552 (N_3552,N_2580,N_2278);
or U3553 (N_3553,N_2462,N_2395);
xnor U3554 (N_3554,N_2223,N_2738);
or U3555 (N_3555,N_2746,N_2910);
nand U3556 (N_3556,N_2715,N_2375);
or U3557 (N_3557,N_2811,N_2689);
nor U3558 (N_3558,N_2329,N_2635);
nand U3559 (N_3559,N_2795,N_2736);
nor U3560 (N_3560,N_2696,N_2941);
or U3561 (N_3561,N_2427,N_2995);
nand U3562 (N_3562,N_2299,N_2088);
nor U3563 (N_3563,N_2597,N_2804);
xor U3564 (N_3564,N_2341,N_2637);
nand U3565 (N_3565,N_2703,N_2117);
nor U3566 (N_3566,N_2237,N_2849);
and U3567 (N_3567,N_2795,N_2151);
and U3568 (N_3568,N_2486,N_2181);
or U3569 (N_3569,N_2780,N_2398);
nor U3570 (N_3570,N_2528,N_2032);
nor U3571 (N_3571,N_2089,N_2802);
and U3572 (N_3572,N_2050,N_2511);
xor U3573 (N_3573,N_2893,N_2005);
or U3574 (N_3574,N_2159,N_2772);
nand U3575 (N_3575,N_2909,N_2281);
xor U3576 (N_3576,N_2317,N_2583);
or U3577 (N_3577,N_2979,N_2818);
and U3578 (N_3578,N_2786,N_2785);
and U3579 (N_3579,N_2288,N_2998);
and U3580 (N_3580,N_2264,N_2261);
or U3581 (N_3581,N_2916,N_2306);
nor U3582 (N_3582,N_2460,N_2498);
nand U3583 (N_3583,N_2384,N_2742);
and U3584 (N_3584,N_2424,N_2139);
or U3585 (N_3585,N_2290,N_2346);
or U3586 (N_3586,N_2459,N_2416);
xnor U3587 (N_3587,N_2928,N_2109);
xor U3588 (N_3588,N_2332,N_2672);
xnor U3589 (N_3589,N_2747,N_2814);
and U3590 (N_3590,N_2536,N_2247);
and U3591 (N_3591,N_2391,N_2380);
or U3592 (N_3592,N_2737,N_2009);
nand U3593 (N_3593,N_2211,N_2532);
nor U3594 (N_3594,N_2974,N_2825);
xnor U3595 (N_3595,N_2007,N_2914);
and U3596 (N_3596,N_2321,N_2687);
nand U3597 (N_3597,N_2450,N_2289);
or U3598 (N_3598,N_2417,N_2712);
xor U3599 (N_3599,N_2403,N_2636);
xnor U3600 (N_3600,N_2435,N_2010);
or U3601 (N_3601,N_2540,N_2379);
or U3602 (N_3602,N_2290,N_2737);
nor U3603 (N_3603,N_2856,N_2057);
or U3604 (N_3604,N_2953,N_2101);
nor U3605 (N_3605,N_2067,N_2512);
or U3606 (N_3606,N_2135,N_2060);
xnor U3607 (N_3607,N_2160,N_2715);
nor U3608 (N_3608,N_2409,N_2129);
xor U3609 (N_3609,N_2550,N_2347);
nand U3610 (N_3610,N_2770,N_2057);
or U3611 (N_3611,N_2775,N_2739);
nor U3612 (N_3612,N_2749,N_2274);
nor U3613 (N_3613,N_2294,N_2746);
and U3614 (N_3614,N_2051,N_2493);
or U3615 (N_3615,N_2781,N_2428);
nand U3616 (N_3616,N_2089,N_2600);
nor U3617 (N_3617,N_2701,N_2765);
nand U3618 (N_3618,N_2415,N_2236);
xor U3619 (N_3619,N_2048,N_2108);
nand U3620 (N_3620,N_2563,N_2766);
and U3621 (N_3621,N_2005,N_2622);
nand U3622 (N_3622,N_2652,N_2547);
nand U3623 (N_3623,N_2440,N_2986);
or U3624 (N_3624,N_2101,N_2804);
or U3625 (N_3625,N_2303,N_2751);
nand U3626 (N_3626,N_2462,N_2379);
nand U3627 (N_3627,N_2299,N_2311);
nand U3628 (N_3628,N_2269,N_2816);
and U3629 (N_3629,N_2884,N_2383);
and U3630 (N_3630,N_2151,N_2929);
and U3631 (N_3631,N_2321,N_2547);
nor U3632 (N_3632,N_2983,N_2876);
nand U3633 (N_3633,N_2619,N_2323);
and U3634 (N_3634,N_2603,N_2500);
nand U3635 (N_3635,N_2674,N_2485);
or U3636 (N_3636,N_2854,N_2637);
nor U3637 (N_3637,N_2101,N_2779);
nor U3638 (N_3638,N_2196,N_2566);
nor U3639 (N_3639,N_2438,N_2732);
or U3640 (N_3640,N_2382,N_2596);
nor U3641 (N_3641,N_2514,N_2775);
and U3642 (N_3642,N_2588,N_2384);
nand U3643 (N_3643,N_2431,N_2474);
nand U3644 (N_3644,N_2428,N_2934);
nor U3645 (N_3645,N_2786,N_2509);
and U3646 (N_3646,N_2027,N_2515);
nor U3647 (N_3647,N_2730,N_2391);
nor U3648 (N_3648,N_2151,N_2142);
nand U3649 (N_3649,N_2983,N_2758);
nand U3650 (N_3650,N_2755,N_2423);
xnor U3651 (N_3651,N_2578,N_2357);
nor U3652 (N_3652,N_2379,N_2453);
nor U3653 (N_3653,N_2206,N_2126);
nor U3654 (N_3654,N_2195,N_2109);
or U3655 (N_3655,N_2675,N_2353);
and U3656 (N_3656,N_2497,N_2103);
and U3657 (N_3657,N_2600,N_2313);
nand U3658 (N_3658,N_2776,N_2726);
nor U3659 (N_3659,N_2763,N_2928);
nor U3660 (N_3660,N_2818,N_2514);
xnor U3661 (N_3661,N_2968,N_2831);
nand U3662 (N_3662,N_2968,N_2777);
or U3663 (N_3663,N_2351,N_2827);
xor U3664 (N_3664,N_2430,N_2705);
nor U3665 (N_3665,N_2260,N_2615);
or U3666 (N_3666,N_2165,N_2721);
nor U3667 (N_3667,N_2103,N_2303);
nor U3668 (N_3668,N_2134,N_2848);
xor U3669 (N_3669,N_2703,N_2294);
and U3670 (N_3670,N_2807,N_2110);
nor U3671 (N_3671,N_2895,N_2160);
nand U3672 (N_3672,N_2498,N_2598);
nor U3673 (N_3673,N_2876,N_2193);
and U3674 (N_3674,N_2536,N_2044);
xnor U3675 (N_3675,N_2863,N_2175);
nor U3676 (N_3676,N_2135,N_2874);
nand U3677 (N_3677,N_2845,N_2658);
nand U3678 (N_3678,N_2863,N_2059);
and U3679 (N_3679,N_2860,N_2530);
or U3680 (N_3680,N_2191,N_2847);
xor U3681 (N_3681,N_2523,N_2600);
or U3682 (N_3682,N_2970,N_2389);
and U3683 (N_3683,N_2247,N_2136);
xnor U3684 (N_3684,N_2877,N_2965);
and U3685 (N_3685,N_2557,N_2478);
nor U3686 (N_3686,N_2063,N_2514);
xnor U3687 (N_3687,N_2739,N_2189);
or U3688 (N_3688,N_2516,N_2361);
or U3689 (N_3689,N_2392,N_2753);
or U3690 (N_3690,N_2965,N_2373);
and U3691 (N_3691,N_2922,N_2819);
xor U3692 (N_3692,N_2841,N_2536);
nor U3693 (N_3693,N_2894,N_2336);
nand U3694 (N_3694,N_2937,N_2206);
xor U3695 (N_3695,N_2764,N_2716);
xnor U3696 (N_3696,N_2876,N_2861);
xnor U3697 (N_3697,N_2425,N_2112);
and U3698 (N_3698,N_2971,N_2421);
or U3699 (N_3699,N_2587,N_2401);
nor U3700 (N_3700,N_2027,N_2961);
nand U3701 (N_3701,N_2066,N_2627);
xnor U3702 (N_3702,N_2227,N_2698);
xor U3703 (N_3703,N_2102,N_2461);
nor U3704 (N_3704,N_2989,N_2644);
and U3705 (N_3705,N_2880,N_2612);
nor U3706 (N_3706,N_2767,N_2248);
and U3707 (N_3707,N_2005,N_2514);
and U3708 (N_3708,N_2792,N_2929);
and U3709 (N_3709,N_2185,N_2107);
or U3710 (N_3710,N_2400,N_2949);
nand U3711 (N_3711,N_2266,N_2741);
or U3712 (N_3712,N_2729,N_2459);
nand U3713 (N_3713,N_2859,N_2576);
or U3714 (N_3714,N_2389,N_2359);
nand U3715 (N_3715,N_2669,N_2024);
or U3716 (N_3716,N_2007,N_2383);
or U3717 (N_3717,N_2811,N_2960);
xnor U3718 (N_3718,N_2175,N_2742);
nor U3719 (N_3719,N_2256,N_2084);
or U3720 (N_3720,N_2793,N_2162);
and U3721 (N_3721,N_2209,N_2966);
nand U3722 (N_3722,N_2740,N_2663);
nor U3723 (N_3723,N_2521,N_2964);
nor U3724 (N_3724,N_2992,N_2891);
xor U3725 (N_3725,N_2510,N_2133);
nor U3726 (N_3726,N_2802,N_2413);
xor U3727 (N_3727,N_2471,N_2360);
nand U3728 (N_3728,N_2122,N_2439);
or U3729 (N_3729,N_2326,N_2960);
nor U3730 (N_3730,N_2450,N_2111);
or U3731 (N_3731,N_2356,N_2716);
and U3732 (N_3732,N_2531,N_2827);
nor U3733 (N_3733,N_2497,N_2718);
xor U3734 (N_3734,N_2420,N_2966);
or U3735 (N_3735,N_2588,N_2130);
and U3736 (N_3736,N_2779,N_2698);
nand U3737 (N_3737,N_2861,N_2065);
or U3738 (N_3738,N_2006,N_2071);
or U3739 (N_3739,N_2471,N_2251);
and U3740 (N_3740,N_2068,N_2988);
nor U3741 (N_3741,N_2395,N_2042);
nor U3742 (N_3742,N_2970,N_2115);
xor U3743 (N_3743,N_2389,N_2428);
and U3744 (N_3744,N_2795,N_2746);
nand U3745 (N_3745,N_2206,N_2585);
nor U3746 (N_3746,N_2458,N_2297);
xor U3747 (N_3747,N_2905,N_2400);
xor U3748 (N_3748,N_2718,N_2937);
and U3749 (N_3749,N_2466,N_2116);
xnor U3750 (N_3750,N_2564,N_2427);
xnor U3751 (N_3751,N_2556,N_2597);
xnor U3752 (N_3752,N_2133,N_2304);
xnor U3753 (N_3753,N_2631,N_2959);
nand U3754 (N_3754,N_2118,N_2412);
nor U3755 (N_3755,N_2089,N_2252);
nand U3756 (N_3756,N_2328,N_2399);
or U3757 (N_3757,N_2891,N_2110);
and U3758 (N_3758,N_2968,N_2948);
or U3759 (N_3759,N_2995,N_2379);
or U3760 (N_3760,N_2942,N_2465);
and U3761 (N_3761,N_2529,N_2844);
nor U3762 (N_3762,N_2213,N_2929);
nand U3763 (N_3763,N_2097,N_2813);
xor U3764 (N_3764,N_2135,N_2611);
nand U3765 (N_3765,N_2208,N_2849);
nand U3766 (N_3766,N_2557,N_2942);
and U3767 (N_3767,N_2718,N_2658);
xnor U3768 (N_3768,N_2603,N_2320);
nand U3769 (N_3769,N_2225,N_2532);
or U3770 (N_3770,N_2304,N_2804);
and U3771 (N_3771,N_2670,N_2520);
nand U3772 (N_3772,N_2548,N_2899);
xnor U3773 (N_3773,N_2681,N_2596);
xor U3774 (N_3774,N_2987,N_2288);
or U3775 (N_3775,N_2735,N_2870);
and U3776 (N_3776,N_2009,N_2340);
and U3777 (N_3777,N_2350,N_2039);
xnor U3778 (N_3778,N_2102,N_2978);
or U3779 (N_3779,N_2548,N_2683);
or U3780 (N_3780,N_2158,N_2742);
xnor U3781 (N_3781,N_2300,N_2898);
and U3782 (N_3782,N_2501,N_2737);
and U3783 (N_3783,N_2936,N_2357);
nor U3784 (N_3784,N_2417,N_2285);
nand U3785 (N_3785,N_2648,N_2297);
or U3786 (N_3786,N_2792,N_2909);
nand U3787 (N_3787,N_2486,N_2122);
nand U3788 (N_3788,N_2928,N_2236);
nand U3789 (N_3789,N_2370,N_2663);
xor U3790 (N_3790,N_2037,N_2485);
xor U3791 (N_3791,N_2892,N_2359);
xnor U3792 (N_3792,N_2667,N_2161);
nor U3793 (N_3793,N_2491,N_2970);
xnor U3794 (N_3794,N_2177,N_2284);
and U3795 (N_3795,N_2044,N_2372);
nand U3796 (N_3796,N_2774,N_2096);
nand U3797 (N_3797,N_2589,N_2905);
or U3798 (N_3798,N_2310,N_2194);
or U3799 (N_3799,N_2454,N_2579);
or U3800 (N_3800,N_2357,N_2057);
and U3801 (N_3801,N_2051,N_2401);
xnor U3802 (N_3802,N_2764,N_2724);
and U3803 (N_3803,N_2233,N_2043);
and U3804 (N_3804,N_2487,N_2039);
nand U3805 (N_3805,N_2431,N_2324);
xnor U3806 (N_3806,N_2484,N_2792);
xnor U3807 (N_3807,N_2478,N_2652);
nor U3808 (N_3808,N_2718,N_2684);
or U3809 (N_3809,N_2536,N_2228);
nand U3810 (N_3810,N_2047,N_2104);
or U3811 (N_3811,N_2472,N_2968);
xor U3812 (N_3812,N_2832,N_2705);
xnor U3813 (N_3813,N_2569,N_2382);
xor U3814 (N_3814,N_2482,N_2397);
xor U3815 (N_3815,N_2045,N_2039);
and U3816 (N_3816,N_2465,N_2843);
nand U3817 (N_3817,N_2814,N_2332);
or U3818 (N_3818,N_2611,N_2717);
xnor U3819 (N_3819,N_2129,N_2713);
and U3820 (N_3820,N_2292,N_2672);
and U3821 (N_3821,N_2216,N_2288);
nor U3822 (N_3822,N_2652,N_2873);
nor U3823 (N_3823,N_2677,N_2146);
xor U3824 (N_3824,N_2382,N_2418);
xnor U3825 (N_3825,N_2805,N_2446);
nand U3826 (N_3826,N_2647,N_2415);
nor U3827 (N_3827,N_2331,N_2824);
or U3828 (N_3828,N_2613,N_2370);
and U3829 (N_3829,N_2833,N_2768);
and U3830 (N_3830,N_2755,N_2403);
nand U3831 (N_3831,N_2545,N_2844);
nor U3832 (N_3832,N_2659,N_2405);
xor U3833 (N_3833,N_2677,N_2299);
or U3834 (N_3834,N_2981,N_2361);
xnor U3835 (N_3835,N_2276,N_2644);
nand U3836 (N_3836,N_2786,N_2820);
and U3837 (N_3837,N_2604,N_2972);
nand U3838 (N_3838,N_2108,N_2798);
nor U3839 (N_3839,N_2515,N_2963);
or U3840 (N_3840,N_2048,N_2656);
or U3841 (N_3841,N_2834,N_2220);
xnor U3842 (N_3842,N_2929,N_2384);
and U3843 (N_3843,N_2938,N_2030);
nor U3844 (N_3844,N_2891,N_2359);
and U3845 (N_3845,N_2688,N_2631);
nand U3846 (N_3846,N_2724,N_2608);
nand U3847 (N_3847,N_2458,N_2174);
nor U3848 (N_3848,N_2429,N_2391);
and U3849 (N_3849,N_2750,N_2880);
and U3850 (N_3850,N_2379,N_2720);
and U3851 (N_3851,N_2221,N_2923);
and U3852 (N_3852,N_2014,N_2786);
and U3853 (N_3853,N_2937,N_2560);
nor U3854 (N_3854,N_2220,N_2461);
or U3855 (N_3855,N_2086,N_2926);
or U3856 (N_3856,N_2698,N_2501);
and U3857 (N_3857,N_2216,N_2554);
nand U3858 (N_3858,N_2045,N_2290);
nand U3859 (N_3859,N_2630,N_2285);
nand U3860 (N_3860,N_2112,N_2512);
and U3861 (N_3861,N_2819,N_2750);
nand U3862 (N_3862,N_2337,N_2095);
nor U3863 (N_3863,N_2427,N_2589);
xor U3864 (N_3864,N_2504,N_2864);
xnor U3865 (N_3865,N_2747,N_2137);
nand U3866 (N_3866,N_2619,N_2838);
nand U3867 (N_3867,N_2055,N_2307);
or U3868 (N_3868,N_2430,N_2652);
xnor U3869 (N_3869,N_2579,N_2427);
and U3870 (N_3870,N_2760,N_2940);
or U3871 (N_3871,N_2686,N_2830);
nor U3872 (N_3872,N_2210,N_2473);
nor U3873 (N_3873,N_2929,N_2055);
or U3874 (N_3874,N_2850,N_2330);
or U3875 (N_3875,N_2836,N_2078);
or U3876 (N_3876,N_2690,N_2562);
nor U3877 (N_3877,N_2136,N_2054);
nor U3878 (N_3878,N_2237,N_2255);
nand U3879 (N_3879,N_2091,N_2972);
nand U3880 (N_3880,N_2157,N_2574);
xnor U3881 (N_3881,N_2366,N_2237);
nand U3882 (N_3882,N_2405,N_2462);
and U3883 (N_3883,N_2897,N_2105);
or U3884 (N_3884,N_2607,N_2959);
or U3885 (N_3885,N_2986,N_2209);
or U3886 (N_3886,N_2713,N_2198);
and U3887 (N_3887,N_2279,N_2186);
or U3888 (N_3888,N_2777,N_2956);
and U3889 (N_3889,N_2761,N_2303);
and U3890 (N_3890,N_2135,N_2552);
or U3891 (N_3891,N_2479,N_2530);
or U3892 (N_3892,N_2322,N_2005);
and U3893 (N_3893,N_2658,N_2139);
and U3894 (N_3894,N_2599,N_2762);
nand U3895 (N_3895,N_2403,N_2563);
nor U3896 (N_3896,N_2987,N_2043);
nand U3897 (N_3897,N_2596,N_2847);
nor U3898 (N_3898,N_2668,N_2873);
nand U3899 (N_3899,N_2899,N_2498);
nand U3900 (N_3900,N_2638,N_2916);
nor U3901 (N_3901,N_2963,N_2753);
or U3902 (N_3902,N_2607,N_2350);
and U3903 (N_3903,N_2624,N_2581);
nor U3904 (N_3904,N_2877,N_2968);
nand U3905 (N_3905,N_2133,N_2036);
nand U3906 (N_3906,N_2588,N_2908);
and U3907 (N_3907,N_2290,N_2515);
or U3908 (N_3908,N_2289,N_2133);
nor U3909 (N_3909,N_2863,N_2762);
nor U3910 (N_3910,N_2163,N_2578);
nor U3911 (N_3911,N_2699,N_2840);
and U3912 (N_3912,N_2990,N_2941);
xor U3913 (N_3913,N_2928,N_2038);
nand U3914 (N_3914,N_2886,N_2394);
xnor U3915 (N_3915,N_2135,N_2095);
nand U3916 (N_3916,N_2450,N_2664);
xor U3917 (N_3917,N_2180,N_2849);
or U3918 (N_3918,N_2619,N_2770);
xnor U3919 (N_3919,N_2530,N_2348);
and U3920 (N_3920,N_2610,N_2597);
xnor U3921 (N_3921,N_2069,N_2987);
or U3922 (N_3922,N_2111,N_2786);
or U3923 (N_3923,N_2762,N_2464);
and U3924 (N_3924,N_2822,N_2932);
or U3925 (N_3925,N_2992,N_2238);
and U3926 (N_3926,N_2924,N_2391);
nand U3927 (N_3927,N_2384,N_2485);
or U3928 (N_3928,N_2850,N_2908);
xnor U3929 (N_3929,N_2532,N_2039);
xnor U3930 (N_3930,N_2183,N_2339);
and U3931 (N_3931,N_2960,N_2950);
or U3932 (N_3932,N_2120,N_2925);
xor U3933 (N_3933,N_2213,N_2525);
nor U3934 (N_3934,N_2974,N_2904);
nor U3935 (N_3935,N_2827,N_2230);
nor U3936 (N_3936,N_2110,N_2392);
and U3937 (N_3937,N_2648,N_2922);
and U3938 (N_3938,N_2812,N_2675);
xor U3939 (N_3939,N_2443,N_2510);
nand U3940 (N_3940,N_2897,N_2836);
xnor U3941 (N_3941,N_2080,N_2313);
xor U3942 (N_3942,N_2969,N_2824);
and U3943 (N_3943,N_2068,N_2533);
xnor U3944 (N_3944,N_2416,N_2445);
nand U3945 (N_3945,N_2966,N_2780);
xnor U3946 (N_3946,N_2950,N_2027);
nand U3947 (N_3947,N_2312,N_2887);
or U3948 (N_3948,N_2644,N_2893);
nand U3949 (N_3949,N_2626,N_2463);
and U3950 (N_3950,N_2772,N_2110);
nand U3951 (N_3951,N_2874,N_2710);
nand U3952 (N_3952,N_2435,N_2063);
or U3953 (N_3953,N_2359,N_2088);
or U3954 (N_3954,N_2749,N_2841);
or U3955 (N_3955,N_2326,N_2930);
nand U3956 (N_3956,N_2495,N_2146);
nand U3957 (N_3957,N_2686,N_2512);
nor U3958 (N_3958,N_2105,N_2940);
nand U3959 (N_3959,N_2414,N_2166);
nand U3960 (N_3960,N_2174,N_2563);
and U3961 (N_3961,N_2949,N_2099);
or U3962 (N_3962,N_2181,N_2003);
xor U3963 (N_3963,N_2780,N_2815);
xnor U3964 (N_3964,N_2988,N_2715);
and U3965 (N_3965,N_2350,N_2598);
and U3966 (N_3966,N_2162,N_2548);
or U3967 (N_3967,N_2542,N_2519);
nand U3968 (N_3968,N_2867,N_2624);
nand U3969 (N_3969,N_2744,N_2048);
nor U3970 (N_3970,N_2575,N_2742);
or U3971 (N_3971,N_2336,N_2237);
nor U3972 (N_3972,N_2305,N_2633);
nand U3973 (N_3973,N_2018,N_2306);
nor U3974 (N_3974,N_2057,N_2347);
and U3975 (N_3975,N_2198,N_2107);
and U3976 (N_3976,N_2246,N_2032);
nand U3977 (N_3977,N_2113,N_2121);
and U3978 (N_3978,N_2914,N_2831);
nor U3979 (N_3979,N_2251,N_2493);
nor U3980 (N_3980,N_2084,N_2958);
xnor U3981 (N_3981,N_2774,N_2918);
nand U3982 (N_3982,N_2273,N_2166);
or U3983 (N_3983,N_2814,N_2442);
xor U3984 (N_3984,N_2779,N_2577);
nand U3985 (N_3985,N_2012,N_2948);
nor U3986 (N_3986,N_2793,N_2983);
nand U3987 (N_3987,N_2665,N_2798);
xor U3988 (N_3988,N_2121,N_2073);
xnor U3989 (N_3989,N_2080,N_2319);
or U3990 (N_3990,N_2976,N_2082);
nand U3991 (N_3991,N_2038,N_2229);
nand U3992 (N_3992,N_2174,N_2163);
nor U3993 (N_3993,N_2831,N_2851);
xor U3994 (N_3994,N_2293,N_2919);
nor U3995 (N_3995,N_2041,N_2417);
and U3996 (N_3996,N_2284,N_2587);
xnor U3997 (N_3997,N_2727,N_2360);
and U3998 (N_3998,N_2295,N_2711);
or U3999 (N_3999,N_2544,N_2870);
or U4000 (N_4000,N_3453,N_3686);
xor U4001 (N_4001,N_3014,N_3905);
and U4002 (N_4002,N_3162,N_3287);
and U4003 (N_4003,N_3090,N_3843);
or U4004 (N_4004,N_3527,N_3044);
nand U4005 (N_4005,N_3349,N_3676);
and U4006 (N_4006,N_3280,N_3168);
xnor U4007 (N_4007,N_3050,N_3248);
nand U4008 (N_4008,N_3845,N_3596);
xnor U4009 (N_4009,N_3996,N_3554);
nand U4010 (N_4010,N_3654,N_3602);
xor U4011 (N_4011,N_3141,N_3723);
or U4012 (N_4012,N_3029,N_3551);
nor U4013 (N_4013,N_3609,N_3655);
or U4014 (N_4014,N_3445,N_3166);
xnor U4015 (N_4015,N_3185,N_3399);
nor U4016 (N_4016,N_3652,N_3765);
nor U4017 (N_4017,N_3754,N_3645);
nor U4018 (N_4018,N_3317,N_3762);
xnor U4019 (N_4019,N_3721,N_3827);
nor U4020 (N_4020,N_3859,N_3129);
nand U4021 (N_4021,N_3742,N_3978);
and U4022 (N_4022,N_3821,N_3989);
xnor U4023 (N_4023,N_3476,N_3359);
or U4024 (N_4024,N_3336,N_3632);
nand U4025 (N_4025,N_3277,N_3255);
xor U4026 (N_4026,N_3131,N_3072);
nand U4027 (N_4027,N_3474,N_3697);
and U4028 (N_4028,N_3954,N_3205);
nand U4029 (N_4029,N_3574,N_3640);
nand U4030 (N_4030,N_3970,N_3600);
or U4031 (N_4031,N_3866,N_3641);
nand U4032 (N_4032,N_3709,N_3824);
nand U4033 (N_4033,N_3296,N_3089);
nor U4034 (N_4034,N_3744,N_3499);
and U4035 (N_4035,N_3545,N_3009);
nor U4036 (N_4036,N_3613,N_3030);
xnor U4037 (N_4037,N_3673,N_3668);
nand U4038 (N_4038,N_3599,N_3663);
xor U4039 (N_4039,N_3148,N_3225);
nor U4040 (N_4040,N_3741,N_3471);
nand U4041 (N_4041,N_3900,N_3828);
or U4042 (N_4042,N_3683,N_3959);
and U4043 (N_4043,N_3812,N_3688);
and U4044 (N_4044,N_3625,N_3962);
and U4045 (N_4045,N_3383,N_3245);
nor U4046 (N_4046,N_3229,N_3036);
xor U4047 (N_4047,N_3795,N_3379);
nand U4048 (N_4048,N_3032,N_3739);
xor U4049 (N_4049,N_3509,N_3059);
and U4050 (N_4050,N_3815,N_3111);
xnor U4051 (N_4051,N_3204,N_3005);
nor U4052 (N_4052,N_3098,N_3000);
nor U4053 (N_4053,N_3950,N_3888);
xnor U4054 (N_4054,N_3736,N_3390);
or U4055 (N_4055,N_3043,N_3764);
xor U4056 (N_4056,N_3882,N_3694);
nor U4057 (N_4057,N_3258,N_3108);
or U4058 (N_4058,N_3137,N_3513);
and U4059 (N_4059,N_3535,N_3187);
or U4060 (N_4060,N_3650,N_3102);
and U4061 (N_4061,N_3196,N_3980);
xnor U4062 (N_4062,N_3822,N_3370);
nand U4063 (N_4063,N_3156,N_3426);
nand U4064 (N_4064,N_3218,N_3594);
or U4065 (N_4065,N_3691,N_3793);
and U4066 (N_4066,N_3175,N_3854);
nand U4067 (N_4067,N_3363,N_3995);
xnor U4068 (N_4068,N_3487,N_3100);
nor U4069 (N_4069,N_3113,N_3027);
xnor U4070 (N_4070,N_3687,N_3885);
nor U4071 (N_4071,N_3716,N_3491);
or U4072 (N_4072,N_3073,N_3095);
nand U4073 (N_4073,N_3227,N_3271);
nand U4074 (N_4074,N_3235,N_3555);
xnor U4075 (N_4075,N_3428,N_3348);
xor U4076 (N_4076,N_3610,N_3105);
nor U4077 (N_4077,N_3203,N_3344);
nor U4078 (N_4078,N_3147,N_3870);
and U4079 (N_4079,N_3434,N_3753);
or U4080 (N_4080,N_3669,N_3731);
nand U4081 (N_4081,N_3540,N_3388);
nor U4082 (N_4082,N_3128,N_3897);
and U4083 (N_4083,N_3468,N_3772);
xnor U4084 (N_4084,N_3523,N_3238);
nor U4085 (N_4085,N_3890,N_3435);
or U4086 (N_4086,N_3389,N_3524);
or U4087 (N_4087,N_3957,N_3661);
and U4088 (N_4088,N_3924,N_3405);
nor U4089 (N_4089,N_3759,N_3288);
and U4090 (N_4090,N_3192,N_3174);
nand U4091 (N_4091,N_3157,N_3717);
and U4092 (N_4092,N_3958,N_3126);
or U4093 (N_4093,N_3743,N_3507);
and U4094 (N_4094,N_3211,N_3586);
or U4095 (N_4095,N_3079,N_3464);
and U4096 (N_4096,N_3024,N_3247);
or U4097 (N_4097,N_3355,N_3581);
xnor U4098 (N_4098,N_3286,N_3322);
nor U4099 (N_4099,N_3403,N_3114);
and U4100 (N_4100,N_3585,N_3366);
nor U4101 (N_4101,N_3463,N_3222);
or U4102 (N_4102,N_3398,N_3053);
nor U4103 (N_4103,N_3022,N_3001);
and U4104 (N_4104,N_3981,N_3994);
nor U4105 (N_4105,N_3851,N_3770);
nor U4106 (N_4106,N_3558,N_3844);
xnor U4107 (N_4107,N_3207,N_3932);
nand U4108 (N_4108,N_3076,N_3480);
nor U4109 (N_4109,N_3023,N_3929);
nand U4110 (N_4110,N_3630,N_3530);
nor U4111 (N_4111,N_3293,N_3689);
or U4112 (N_4112,N_3416,N_3488);
xor U4113 (N_4113,N_3942,N_3587);
and U4114 (N_4114,N_3707,N_3608);
nor U4115 (N_4115,N_3516,N_3703);
nand U4116 (N_4116,N_3145,N_3936);
and U4117 (N_4117,N_3228,N_3504);
nand U4118 (N_4118,N_3922,N_3636);
nand U4119 (N_4119,N_3961,N_3969);
nor U4120 (N_4120,N_3150,N_3629);
nor U4121 (N_4121,N_3603,N_3733);
nor U4122 (N_4122,N_3482,N_3015);
or U4123 (N_4123,N_3552,N_3323);
and U4124 (N_4124,N_3070,N_3345);
and U4125 (N_4125,N_3911,N_3814);
and U4126 (N_4126,N_3439,N_3004);
and U4127 (N_4127,N_3262,N_3976);
xor U4128 (N_4128,N_3261,N_3493);
xnor U4129 (N_4129,N_3944,N_3088);
and U4130 (N_4130,N_3003,N_3461);
nand U4131 (N_4131,N_3011,N_3243);
nor U4132 (N_4132,N_3537,N_3106);
and U4133 (N_4133,N_3294,N_3791);
or U4134 (N_4134,N_3894,N_3028);
and U4135 (N_4135,N_3849,N_3952);
xor U4136 (N_4136,N_3916,N_3928);
xnor U4137 (N_4137,N_3542,N_3171);
xnor U4138 (N_4138,N_3183,N_3873);
nor U4139 (N_4139,N_3906,N_3281);
and U4140 (N_4140,N_3257,N_3649);
or U4141 (N_4141,N_3706,N_3841);
nor U4142 (N_4142,N_3583,N_3877);
nand U4143 (N_4143,N_3184,N_3884);
or U4144 (N_4144,N_3808,N_3013);
nor U4145 (N_4145,N_3202,N_3648);
or U4146 (N_4146,N_3968,N_3677);
and U4147 (N_4147,N_3452,N_3240);
nand U4148 (N_4148,N_3084,N_3146);
or U4149 (N_4149,N_3457,N_3879);
xnor U4150 (N_4150,N_3949,N_3943);
xnor U4151 (N_4151,N_3395,N_3283);
nand U4152 (N_4152,N_3582,N_3685);
or U4153 (N_4153,N_3371,N_3241);
nor U4154 (N_4154,N_3833,N_3621);
nor U4155 (N_4155,N_3749,N_3273);
nor U4156 (N_4156,N_3539,N_3373);
nor U4157 (N_4157,N_3892,N_3667);
or U4158 (N_4158,N_3172,N_3510);
nor U4159 (N_4159,N_3490,N_3276);
nand U4160 (N_4160,N_3357,N_3788);
and U4161 (N_4161,N_3986,N_3699);
or U4162 (N_4162,N_3913,N_3475);
xor U4163 (N_4163,N_3740,N_3138);
nor U4164 (N_4164,N_3564,N_3651);
nand U4165 (N_4165,N_3067,N_3285);
xnor U4166 (N_4166,N_3017,N_3498);
and U4167 (N_4167,N_3107,N_3149);
nand U4168 (N_4168,N_3127,N_3034);
xnor U4169 (N_4169,N_3604,N_3020);
xnor U4170 (N_4170,N_3397,N_3769);
nor U4171 (N_4171,N_3834,N_3289);
or U4172 (N_4172,N_3842,N_3058);
or U4173 (N_4173,N_3016,N_3838);
and U4174 (N_4174,N_3720,N_3186);
and U4175 (N_4175,N_3985,N_3557);
or U4176 (N_4176,N_3372,N_3618);
and U4177 (N_4177,N_3075,N_3459);
nor U4178 (N_4178,N_3454,N_3133);
and U4179 (N_4179,N_3292,N_3934);
nor U4180 (N_4180,N_3696,N_3492);
xor U4181 (N_4181,N_3052,N_3546);
xnor U4182 (N_4182,N_3469,N_3449);
nand U4183 (N_4183,N_3615,N_3899);
nand U4184 (N_4184,N_3099,N_3481);
xnor U4185 (N_4185,N_3501,N_3097);
nand U4186 (N_4186,N_3809,N_3565);
xor U4187 (N_4187,N_3031,N_3628);
or U4188 (N_4188,N_3935,N_3531);
nand U4189 (N_4189,N_3143,N_3974);
and U4190 (N_4190,N_3303,N_3216);
nor U4191 (N_4191,N_3406,N_3642);
xnor U4192 (N_4192,N_3310,N_3049);
or U4193 (N_4193,N_3597,N_3591);
nand U4194 (N_4194,N_3737,N_3619);
and U4195 (N_4195,N_3792,N_3221);
nand U4196 (N_4196,N_3901,N_3252);
and U4197 (N_4197,N_3945,N_3614);
and U4198 (N_4198,N_3466,N_3898);
and U4199 (N_4199,N_3035,N_3037);
or U4200 (N_4200,N_3992,N_3332);
or U4201 (N_4201,N_3589,N_3857);
and U4202 (N_4202,N_3063,N_3291);
xnor U4203 (N_4203,N_3334,N_3069);
nand U4204 (N_4204,N_3239,N_3622);
xor U4205 (N_4205,N_3860,N_3083);
xnor U4206 (N_4206,N_3830,N_3269);
nand U4207 (N_4207,N_3701,N_3693);
nand U4208 (N_4208,N_3246,N_3339);
or U4209 (N_4209,N_3012,N_3964);
nor U4210 (N_4210,N_3253,N_3718);
or U4211 (N_4211,N_3606,N_3467);
nand U4212 (N_4212,N_3473,N_3835);
or U4213 (N_4213,N_3160,N_3647);
xnor U4214 (N_4214,N_3477,N_3983);
or U4215 (N_4215,N_3919,N_3508);
and U4216 (N_4216,N_3726,N_3987);
xnor U4217 (N_4217,N_3495,N_3948);
or U4218 (N_4218,N_3190,N_3401);
nand U4219 (N_4219,N_3767,N_3408);
and U4220 (N_4220,N_3132,N_3447);
nor U4221 (N_4221,N_3364,N_3536);
nand U4222 (N_4222,N_3368,N_3019);
or U4223 (N_4223,N_3085,N_3396);
or U4224 (N_4224,N_3313,N_3456);
xor U4225 (N_4225,N_3979,N_3643);
nand U4226 (N_4226,N_3343,N_3025);
xor U4227 (N_4227,N_3635,N_3951);
and U4228 (N_4228,N_3420,N_3074);
nand U4229 (N_4229,N_3863,N_3908);
and U4230 (N_4230,N_3584,N_3886);
nand U4231 (N_4231,N_3521,N_3250);
nor U4232 (N_4232,N_3955,N_3082);
nand U4233 (N_4233,N_3665,N_3623);
nand U4234 (N_4234,N_3165,N_3352);
nor U4235 (N_4235,N_3249,N_3528);
or U4236 (N_4236,N_3680,N_3776);
nor U4237 (N_4237,N_3350,N_3946);
nand U4238 (N_4238,N_3265,N_3967);
xor U4239 (N_4239,N_3392,N_3158);
nor U4240 (N_4240,N_3093,N_3086);
nand U4241 (N_4241,N_3198,N_3181);
or U4242 (N_4242,N_3080,N_3144);
nor U4243 (N_4243,N_3993,N_3917);
and U4244 (N_4244,N_3064,N_3656);
nand U4245 (N_4245,N_3799,N_3316);
nor U4246 (N_4246,N_3297,N_3071);
xor U4247 (N_4247,N_3279,N_3761);
and U4248 (N_4248,N_3541,N_3805);
and U4249 (N_4249,N_3506,N_3358);
nand U4250 (N_4250,N_3872,N_3394);
xor U4251 (N_4251,N_3662,N_3548);
nor U4252 (N_4252,N_3960,N_3818);
or U4253 (N_4253,N_3829,N_3874);
nand U4254 (N_4254,N_3891,N_3728);
nor U4255 (N_4255,N_3876,N_3790);
and U4256 (N_4256,N_3918,N_3400);
or U4257 (N_4257,N_3007,N_3377);
nand U4258 (N_4258,N_3436,N_3909);
and U4259 (N_4259,N_3927,N_3566);
or U4260 (N_4260,N_3505,N_3549);
xnor U4261 (N_4261,N_3333,N_3732);
xor U4262 (N_4262,N_3061,N_3206);
nand U4263 (N_4263,N_3215,N_3458);
or U4264 (N_4264,N_3750,N_3335);
nand U4265 (N_4265,N_3309,N_3646);
or U4266 (N_4266,N_3778,N_3496);
xnor U4267 (N_4267,N_3757,N_3135);
nand U4268 (N_4268,N_3307,N_3404);
xor U4269 (N_4269,N_3605,N_3010);
nor U4270 (N_4270,N_3538,N_3402);
nand U4271 (N_4271,N_3134,N_3806);
xnor U4272 (N_4272,N_3189,N_3451);
nor U4273 (N_4273,N_3547,N_3375);
and U4274 (N_4274,N_3479,N_3612);
nand U4275 (N_4275,N_3163,N_3638);
or U4276 (N_4276,N_3520,N_3485);
or U4277 (N_4277,N_3381,N_3234);
xor U4278 (N_4278,N_3304,N_3956);
nand U4279 (N_4279,N_3801,N_3411);
xor U4280 (N_4280,N_3299,N_3798);
or U4281 (N_4281,N_3616,N_3515);
xor U4282 (N_4282,N_3494,N_3785);
nand U4283 (N_4283,N_3953,N_3284);
nor U4284 (N_4284,N_3511,N_3991);
or U4285 (N_4285,N_3385,N_3182);
and U4286 (N_4286,N_3220,N_3318);
nand U4287 (N_4287,N_3155,N_3775);
nor U4288 (N_4288,N_3940,N_3272);
nor U4289 (N_4289,N_3826,N_3251);
or U4290 (N_4290,N_3021,N_3231);
or U4291 (N_4291,N_3774,N_3807);
nor U4292 (N_4292,N_3698,N_3997);
or U4293 (N_4293,N_3119,N_3054);
or U4294 (N_4294,N_3329,N_3112);
nor U4295 (N_4295,N_3560,N_3161);
xnor U4296 (N_4296,N_3167,N_3766);
or U4297 (N_4297,N_3965,N_3933);
nand U4298 (N_4298,N_3580,N_3443);
nand U4299 (N_4299,N_3224,N_3941);
nand U4300 (N_4300,N_3244,N_3104);
xnor U4301 (N_4301,N_3056,N_3631);
nor U4302 (N_4302,N_3820,N_3208);
xor U4303 (N_4303,N_3925,N_3382);
nand U4304 (N_4304,N_3633,N_3893);
or U4305 (N_4305,N_3045,N_3529);
xor U4306 (N_4306,N_3412,N_3008);
xnor U4307 (N_4307,N_3556,N_3973);
xor U4308 (N_4308,N_3711,N_3188);
xnor U4309 (N_4309,N_3361,N_3771);
nand U4310 (N_4310,N_3553,N_3627);
nor U4311 (N_4311,N_3675,N_3671);
and U4312 (N_4312,N_3522,N_3300);
and U4313 (N_4313,N_3780,N_3164);
or U4314 (N_4314,N_3236,N_3210);
or U4315 (N_4315,N_3990,N_3789);
nor U4316 (N_4316,N_3006,N_3432);
or U4317 (N_4317,N_3122,N_3092);
xnor U4318 (N_4318,N_3429,N_3972);
and U4319 (N_4319,N_3971,N_3173);
nor U4320 (N_4320,N_3786,N_3042);
xnor U4321 (N_4321,N_3330,N_3077);
nor U4322 (N_4322,N_3340,N_3722);
or U4323 (N_4323,N_3773,N_3170);
or U4324 (N_4324,N_3907,N_3051);
and U4325 (N_4325,N_3176,N_3376);
xor U4326 (N_4326,N_3758,N_3440);
or U4327 (N_4327,N_3571,N_3802);
and U4328 (N_4328,N_3214,N_3200);
or U4329 (N_4329,N_3577,N_3048);
nor U4330 (N_4330,N_3847,N_3486);
or U4331 (N_4331,N_3091,N_3532);
and U4332 (N_4332,N_3378,N_3437);
nand U4333 (N_4333,N_3710,N_3777);
xnor U4334 (N_4334,N_3784,N_3904);
xor U4335 (N_4335,N_3427,N_3518);
nor U4336 (N_4336,N_3139,N_3433);
nor U4337 (N_4337,N_3472,N_3861);
or U4338 (N_4338,N_3018,N_3430);
xor U4339 (N_4339,N_3195,N_3837);
xnor U4340 (N_4340,N_3617,N_3217);
or U4341 (N_4341,N_3926,N_3700);
nor U4342 (N_4342,N_3875,N_3197);
and U4343 (N_4343,N_3855,N_3738);
or U4344 (N_4344,N_3853,N_3517);
and U4345 (N_4345,N_3561,N_3569);
and U4346 (N_4346,N_3351,N_3704);
nor U4347 (N_4347,N_3328,N_3380);
nand U4348 (N_4348,N_3142,N_3768);
xnor U4349 (N_4349,N_3319,N_3568);
xnor U4350 (N_4350,N_3823,N_3678);
and U4351 (N_4351,N_3887,N_3444);
xnor U4352 (N_4352,N_3305,N_3998);
nor U4353 (N_4353,N_3338,N_3760);
nor U4354 (N_4354,N_3484,N_3066);
or U4355 (N_4355,N_3460,N_3282);
or U4356 (N_4356,N_3664,N_3356);
and U4357 (N_4357,N_3260,N_3325);
nor U4358 (N_4358,N_3081,N_3354);
and U4359 (N_4359,N_3797,N_3327);
xnor U4360 (N_4360,N_3931,N_3923);
xor U4361 (N_4361,N_3804,N_3575);
nand U4362 (N_4362,N_3109,N_3223);
and U4363 (N_4363,N_3729,N_3423);
nand U4364 (N_4364,N_3078,N_3803);
or U4365 (N_4365,N_3442,N_3154);
nand U4366 (N_4366,N_3410,N_3424);
nor U4367 (N_4367,N_3624,N_3578);
nor U4368 (N_4368,N_3101,N_3441);
nor U4369 (N_4369,N_3407,N_3512);
nor U4370 (N_4370,N_3415,N_3856);
nor U4371 (N_4371,N_3719,N_3832);
or U4372 (N_4372,N_3026,N_3938);
and U4373 (N_4373,N_3103,N_3588);
xnor U4374 (N_4374,N_3094,N_3057);
nand U4375 (N_4375,N_3233,N_3682);
nor U4376 (N_4376,N_3914,N_3858);
and U4377 (N_4377,N_3254,N_3975);
and U4378 (N_4378,N_3118,N_3966);
nand U4379 (N_4379,N_3462,N_3500);
xor U4380 (N_4380,N_3130,N_3681);
xor U4381 (N_4381,N_3751,N_3570);
xnor U4382 (N_4382,N_3865,N_3193);
xor U4383 (N_4383,N_3748,N_3895);
and U4384 (N_4384,N_3620,N_3576);
xnor U4385 (N_4385,N_3705,N_3840);
nor U4386 (N_4386,N_3353,N_3421);
xnor U4387 (N_4387,N_3337,N_3046);
xnor U4388 (N_4388,N_3180,N_3315);
or U4389 (N_4389,N_3320,N_3115);
or U4390 (N_4390,N_3302,N_3867);
xor U4391 (N_4391,N_3674,N_3783);
and U4392 (N_4392,N_3745,N_3713);
nand U4393 (N_4393,N_3690,N_3672);
xnor U4394 (N_4394,N_3868,N_3947);
and U4395 (N_4395,N_3519,N_3369);
xor U4396 (N_4396,N_3136,N_3562);
nand U4397 (N_4397,N_3915,N_3256);
or U4398 (N_4398,N_3230,N_3242);
nand U4399 (N_4399,N_3747,N_3213);
nand U4400 (N_4400,N_3201,N_3819);
nand U4401 (N_4401,N_3725,N_3159);
nor U4402 (N_4402,N_3425,N_3746);
nor U4403 (N_4403,N_3259,N_3544);
nor U4404 (N_4404,N_3982,N_3525);
nor U4405 (N_4405,N_3695,N_3598);
or U4406 (N_4406,N_3209,N_3409);
xnor U4407 (N_4407,N_3431,N_3047);
or U4408 (N_4408,N_3125,N_3883);
or U4409 (N_4409,N_3194,N_3796);
and U4410 (N_4410,N_3559,N_3503);
nand U4411 (N_4411,N_3543,N_3592);
or U4412 (N_4412,N_3607,N_3489);
and U4413 (N_4413,N_3123,N_3422);
nand U4414 (N_4414,N_3573,N_3177);
xor U4415 (N_4415,N_3878,N_3124);
nor U4416 (N_4416,N_3321,N_3367);
nand U4417 (N_4417,N_3880,N_3414);
nor U4418 (N_4418,N_3497,N_3626);
nand U4419 (N_4419,N_3572,N_3324);
nor U4420 (N_4420,N_3116,N_3178);
nand U4421 (N_4421,N_3593,N_3692);
xor U4422 (N_4422,N_3724,N_3391);
or U4423 (N_4423,N_3362,N_3811);
or U4424 (N_4424,N_3274,N_3151);
and U4425 (N_4425,N_3060,N_3684);
nand U4426 (N_4426,N_3590,N_3831);
nor U4427 (N_4427,N_3752,N_3670);
nor U4428 (N_4428,N_3326,N_3921);
or U4429 (N_4429,N_3903,N_3153);
or U4430 (N_4430,N_3963,N_3290);
nor U4431 (N_4431,N_3526,N_3212);
nor U4432 (N_4432,N_3387,N_3312);
nand U4433 (N_4433,N_3679,N_3930);
and U4434 (N_4434,N_3889,N_3852);
or U4435 (N_4435,N_3817,N_3714);
xor U4436 (N_4436,N_3920,N_3653);
nor U4437 (N_4437,N_3869,N_3413);
or U4438 (N_4438,N_3730,N_3278);
nor U4439 (N_4439,N_3306,N_3910);
nand U4440 (N_4440,N_3787,N_3346);
or U4441 (N_4441,N_3735,N_3040);
nand U4442 (N_4442,N_3341,N_3301);
or U4443 (N_4443,N_3386,N_3595);
and U4444 (N_4444,N_3062,N_3419);
and U4445 (N_4445,N_3839,N_3563);
and U4446 (N_4446,N_3448,N_3483);
or U4447 (N_4447,N_3782,N_3110);
and U4448 (N_4448,N_3611,N_3450);
xnor U4449 (N_4449,N_3311,N_3937);
or U4450 (N_4450,N_3756,N_3881);
nand U4451 (N_4451,N_3660,N_3264);
xor U4452 (N_4452,N_3117,N_3902);
and U4453 (N_4453,N_3199,N_3567);
xnor U4454 (N_4454,N_3871,N_3939);
and U4455 (N_4455,N_3275,N_3846);
nor U4456 (N_4456,N_3864,N_3727);
xor U4457 (N_4457,N_3266,N_3836);
nor U4458 (N_4458,N_3298,N_3658);
xor U4459 (N_4459,N_3755,N_3446);
nor U4460 (N_4460,N_3659,N_3219);
and U4461 (N_4461,N_3999,N_3734);
and U4462 (N_4462,N_3169,N_3191);
and U4463 (N_4463,N_3984,N_3268);
or U4464 (N_4464,N_3232,N_3465);
and U4465 (N_4465,N_3140,N_3708);
or U4466 (N_4466,N_3848,N_3237);
nand U4467 (N_4467,N_3666,N_3550);
xnor U4468 (N_4468,N_3712,N_3039);
and U4469 (N_4469,N_3342,N_3781);
and U4470 (N_4470,N_3810,N_3702);
and U4471 (N_4471,N_3657,N_3896);
xor U4472 (N_4472,N_3977,N_3347);
or U4473 (N_4473,N_3179,N_3637);
or U4474 (N_4474,N_3533,N_3634);
nand U4475 (N_4475,N_3226,N_3763);
and U4476 (N_4476,N_3295,N_3514);
xnor U4477 (N_4477,N_3579,N_3639);
nand U4478 (N_4478,N_3988,N_3152);
nor U4479 (N_4479,N_3850,N_3267);
or U4480 (N_4480,N_3816,N_3644);
and U4481 (N_4481,N_3087,N_3041);
or U4482 (N_4482,N_3038,N_3384);
nor U4483 (N_4483,N_3502,N_3331);
nand U4484 (N_4484,N_3794,N_3601);
nor U4485 (N_4485,N_3800,N_3068);
xnor U4486 (N_4486,N_3270,N_3417);
or U4487 (N_4487,N_3418,N_3374);
xnor U4488 (N_4488,N_3096,N_3121);
or U4489 (N_4489,N_3365,N_3033);
xor U4490 (N_4490,N_3912,N_3308);
xnor U4491 (N_4491,N_3534,N_3393);
nand U4492 (N_4492,N_3360,N_3455);
nor U4493 (N_4493,N_3715,N_3055);
nor U4494 (N_4494,N_3813,N_3065);
xor U4495 (N_4495,N_3438,N_3862);
nor U4496 (N_4496,N_3478,N_3779);
and U4497 (N_4497,N_3120,N_3470);
or U4498 (N_4498,N_3263,N_3825);
nor U4499 (N_4499,N_3002,N_3314);
or U4500 (N_4500,N_3080,N_3769);
xor U4501 (N_4501,N_3172,N_3569);
and U4502 (N_4502,N_3320,N_3844);
or U4503 (N_4503,N_3516,N_3911);
nor U4504 (N_4504,N_3623,N_3237);
xor U4505 (N_4505,N_3317,N_3256);
and U4506 (N_4506,N_3570,N_3760);
nor U4507 (N_4507,N_3601,N_3033);
xor U4508 (N_4508,N_3149,N_3097);
nor U4509 (N_4509,N_3040,N_3551);
nor U4510 (N_4510,N_3619,N_3511);
nor U4511 (N_4511,N_3416,N_3355);
nand U4512 (N_4512,N_3052,N_3890);
or U4513 (N_4513,N_3526,N_3708);
nand U4514 (N_4514,N_3952,N_3789);
or U4515 (N_4515,N_3363,N_3515);
xnor U4516 (N_4516,N_3188,N_3855);
nor U4517 (N_4517,N_3239,N_3760);
nand U4518 (N_4518,N_3465,N_3412);
and U4519 (N_4519,N_3584,N_3581);
or U4520 (N_4520,N_3330,N_3812);
nand U4521 (N_4521,N_3594,N_3751);
nand U4522 (N_4522,N_3541,N_3301);
or U4523 (N_4523,N_3477,N_3110);
or U4524 (N_4524,N_3506,N_3416);
and U4525 (N_4525,N_3445,N_3603);
xor U4526 (N_4526,N_3160,N_3641);
nand U4527 (N_4527,N_3159,N_3195);
and U4528 (N_4528,N_3873,N_3970);
nand U4529 (N_4529,N_3342,N_3889);
nand U4530 (N_4530,N_3438,N_3759);
nor U4531 (N_4531,N_3298,N_3211);
nand U4532 (N_4532,N_3475,N_3487);
or U4533 (N_4533,N_3826,N_3365);
or U4534 (N_4534,N_3975,N_3940);
xor U4535 (N_4535,N_3725,N_3783);
and U4536 (N_4536,N_3218,N_3208);
or U4537 (N_4537,N_3789,N_3472);
nand U4538 (N_4538,N_3558,N_3784);
or U4539 (N_4539,N_3225,N_3252);
and U4540 (N_4540,N_3280,N_3063);
nand U4541 (N_4541,N_3557,N_3229);
or U4542 (N_4542,N_3706,N_3151);
nor U4543 (N_4543,N_3481,N_3238);
nand U4544 (N_4544,N_3505,N_3851);
or U4545 (N_4545,N_3338,N_3954);
nor U4546 (N_4546,N_3566,N_3317);
nand U4547 (N_4547,N_3087,N_3590);
and U4548 (N_4548,N_3086,N_3593);
or U4549 (N_4549,N_3436,N_3078);
xnor U4550 (N_4550,N_3074,N_3669);
nand U4551 (N_4551,N_3904,N_3307);
nor U4552 (N_4552,N_3952,N_3381);
and U4553 (N_4553,N_3819,N_3689);
nor U4554 (N_4554,N_3875,N_3865);
or U4555 (N_4555,N_3159,N_3710);
xnor U4556 (N_4556,N_3098,N_3373);
nor U4557 (N_4557,N_3452,N_3690);
xnor U4558 (N_4558,N_3736,N_3933);
and U4559 (N_4559,N_3351,N_3194);
nand U4560 (N_4560,N_3673,N_3503);
and U4561 (N_4561,N_3220,N_3518);
or U4562 (N_4562,N_3660,N_3344);
and U4563 (N_4563,N_3982,N_3035);
xor U4564 (N_4564,N_3726,N_3753);
nor U4565 (N_4565,N_3242,N_3674);
nor U4566 (N_4566,N_3875,N_3138);
nand U4567 (N_4567,N_3987,N_3006);
or U4568 (N_4568,N_3840,N_3930);
nand U4569 (N_4569,N_3562,N_3835);
nor U4570 (N_4570,N_3707,N_3125);
nor U4571 (N_4571,N_3220,N_3243);
or U4572 (N_4572,N_3249,N_3938);
xor U4573 (N_4573,N_3371,N_3871);
or U4574 (N_4574,N_3405,N_3447);
nor U4575 (N_4575,N_3506,N_3408);
nand U4576 (N_4576,N_3638,N_3504);
or U4577 (N_4577,N_3394,N_3378);
xnor U4578 (N_4578,N_3418,N_3012);
or U4579 (N_4579,N_3977,N_3173);
nor U4580 (N_4580,N_3691,N_3438);
nor U4581 (N_4581,N_3446,N_3726);
or U4582 (N_4582,N_3622,N_3541);
and U4583 (N_4583,N_3252,N_3791);
or U4584 (N_4584,N_3154,N_3061);
nor U4585 (N_4585,N_3110,N_3821);
nand U4586 (N_4586,N_3009,N_3467);
or U4587 (N_4587,N_3984,N_3446);
or U4588 (N_4588,N_3967,N_3254);
or U4589 (N_4589,N_3510,N_3112);
xnor U4590 (N_4590,N_3348,N_3449);
and U4591 (N_4591,N_3215,N_3810);
or U4592 (N_4592,N_3626,N_3551);
nor U4593 (N_4593,N_3553,N_3823);
xor U4594 (N_4594,N_3938,N_3904);
nor U4595 (N_4595,N_3528,N_3911);
nor U4596 (N_4596,N_3628,N_3387);
xor U4597 (N_4597,N_3301,N_3389);
or U4598 (N_4598,N_3562,N_3883);
or U4599 (N_4599,N_3571,N_3430);
nor U4600 (N_4600,N_3630,N_3565);
and U4601 (N_4601,N_3201,N_3865);
nand U4602 (N_4602,N_3021,N_3735);
xor U4603 (N_4603,N_3864,N_3180);
nor U4604 (N_4604,N_3892,N_3472);
nand U4605 (N_4605,N_3665,N_3746);
nand U4606 (N_4606,N_3022,N_3821);
nand U4607 (N_4607,N_3000,N_3612);
nand U4608 (N_4608,N_3361,N_3875);
and U4609 (N_4609,N_3051,N_3108);
and U4610 (N_4610,N_3111,N_3552);
or U4611 (N_4611,N_3555,N_3915);
or U4612 (N_4612,N_3238,N_3842);
or U4613 (N_4613,N_3942,N_3569);
and U4614 (N_4614,N_3091,N_3402);
and U4615 (N_4615,N_3075,N_3341);
nor U4616 (N_4616,N_3842,N_3801);
nand U4617 (N_4617,N_3819,N_3648);
xor U4618 (N_4618,N_3363,N_3021);
xnor U4619 (N_4619,N_3962,N_3248);
and U4620 (N_4620,N_3581,N_3857);
xnor U4621 (N_4621,N_3939,N_3022);
or U4622 (N_4622,N_3767,N_3058);
or U4623 (N_4623,N_3839,N_3598);
xnor U4624 (N_4624,N_3059,N_3499);
nand U4625 (N_4625,N_3438,N_3344);
or U4626 (N_4626,N_3229,N_3530);
xor U4627 (N_4627,N_3754,N_3248);
or U4628 (N_4628,N_3334,N_3961);
nand U4629 (N_4629,N_3912,N_3027);
xnor U4630 (N_4630,N_3809,N_3381);
nor U4631 (N_4631,N_3965,N_3489);
nand U4632 (N_4632,N_3701,N_3425);
nand U4633 (N_4633,N_3809,N_3999);
and U4634 (N_4634,N_3168,N_3264);
nor U4635 (N_4635,N_3947,N_3857);
and U4636 (N_4636,N_3199,N_3033);
nor U4637 (N_4637,N_3795,N_3746);
xnor U4638 (N_4638,N_3448,N_3109);
nand U4639 (N_4639,N_3568,N_3257);
nand U4640 (N_4640,N_3599,N_3221);
or U4641 (N_4641,N_3420,N_3485);
nand U4642 (N_4642,N_3274,N_3227);
nand U4643 (N_4643,N_3324,N_3145);
xor U4644 (N_4644,N_3704,N_3176);
and U4645 (N_4645,N_3185,N_3156);
xor U4646 (N_4646,N_3874,N_3597);
nor U4647 (N_4647,N_3225,N_3978);
and U4648 (N_4648,N_3997,N_3680);
nand U4649 (N_4649,N_3781,N_3685);
nand U4650 (N_4650,N_3153,N_3445);
or U4651 (N_4651,N_3671,N_3826);
or U4652 (N_4652,N_3021,N_3981);
nor U4653 (N_4653,N_3601,N_3929);
xor U4654 (N_4654,N_3477,N_3066);
xnor U4655 (N_4655,N_3234,N_3650);
or U4656 (N_4656,N_3617,N_3781);
nor U4657 (N_4657,N_3637,N_3794);
or U4658 (N_4658,N_3957,N_3106);
xnor U4659 (N_4659,N_3777,N_3480);
nand U4660 (N_4660,N_3941,N_3331);
nand U4661 (N_4661,N_3477,N_3014);
or U4662 (N_4662,N_3792,N_3461);
xnor U4663 (N_4663,N_3821,N_3087);
and U4664 (N_4664,N_3652,N_3120);
and U4665 (N_4665,N_3146,N_3580);
xnor U4666 (N_4666,N_3818,N_3681);
nand U4667 (N_4667,N_3517,N_3333);
or U4668 (N_4668,N_3611,N_3363);
nor U4669 (N_4669,N_3230,N_3984);
xor U4670 (N_4670,N_3573,N_3964);
and U4671 (N_4671,N_3538,N_3014);
and U4672 (N_4672,N_3151,N_3053);
and U4673 (N_4673,N_3352,N_3420);
or U4674 (N_4674,N_3398,N_3108);
or U4675 (N_4675,N_3951,N_3350);
and U4676 (N_4676,N_3653,N_3428);
xor U4677 (N_4677,N_3304,N_3189);
xor U4678 (N_4678,N_3352,N_3140);
or U4679 (N_4679,N_3550,N_3797);
xnor U4680 (N_4680,N_3048,N_3104);
and U4681 (N_4681,N_3187,N_3038);
nor U4682 (N_4682,N_3704,N_3481);
and U4683 (N_4683,N_3818,N_3380);
xnor U4684 (N_4684,N_3778,N_3043);
xor U4685 (N_4685,N_3936,N_3358);
nor U4686 (N_4686,N_3236,N_3116);
nand U4687 (N_4687,N_3564,N_3021);
and U4688 (N_4688,N_3177,N_3733);
and U4689 (N_4689,N_3868,N_3354);
or U4690 (N_4690,N_3719,N_3774);
nor U4691 (N_4691,N_3193,N_3797);
xor U4692 (N_4692,N_3595,N_3970);
nand U4693 (N_4693,N_3646,N_3478);
nor U4694 (N_4694,N_3332,N_3629);
and U4695 (N_4695,N_3575,N_3961);
or U4696 (N_4696,N_3088,N_3858);
or U4697 (N_4697,N_3645,N_3181);
and U4698 (N_4698,N_3922,N_3434);
nor U4699 (N_4699,N_3377,N_3935);
or U4700 (N_4700,N_3218,N_3135);
and U4701 (N_4701,N_3214,N_3189);
xnor U4702 (N_4702,N_3145,N_3339);
and U4703 (N_4703,N_3105,N_3653);
nor U4704 (N_4704,N_3888,N_3788);
nor U4705 (N_4705,N_3564,N_3992);
nor U4706 (N_4706,N_3143,N_3951);
nor U4707 (N_4707,N_3982,N_3710);
or U4708 (N_4708,N_3866,N_3752);
nand U4709 (N_4709,N_3831,N_3655);
nor U4710 (N_4710,N_3392,N_3660);
nor U4711 (N_4711,N_3505,N_3639);
xor U4712 (N_4712,N_3476,N_3625);
or U4713 (N_4713,N_3210,N_3179);
nand U4714 (N_4714,N_3036,N_3043);
nand U4715 (N_4715,N_3726,N_3410);
nor U4716 (N_4716,N_3161,N_3121);
nand U4717 (N_4717,N_3480,N_3534);
or U4718 (N_4718,N_3895,N_3597);
and U4719 (N_4719,N_3402,N_3208);
and U4720 (N_4720,N_3380,N_3084);
and U4721 (N_4721,N_3810,N_3277);
nand U4722 (N_4722,N_3908,N_3962);
xnor U4723 (N_4723,N_3213,N_3663);
xnor U4724 (N_4724,N_3559,N_3747);
nor U4725 (N_4725,N_3692,N_3146);
xor U4726 (N_4726,N_3821,N_3421);
nor U4727 (N_4727,N_3664,N_3949);
and U4728 (N_4728,N_3106,N_3254);
xnor U4729 (N_4729,N_3935,N_3587);
nor U4730 (N_4730,N_3296,N_3032);
or U4731 (N_4731,N_3138,N_3773);
nor U4732 (N_4732,N_3905,N_3182);
nor U4733 (N_4733,N_3065,N_3586);
nand U4734 (N_4734,N_3473,N_3237);
nand U4735 (N_4735,N_3455,N_3887);
or U4736 (N_4736,N_3371,N_3720);
xor U4737 (N_4737,N_3396,N_3350);
nand U4738 (N_4738,N_3816,N_3638);
xnor U4739 (N_4739,N_3613,N_3547);
and U4740 (N_4740,N_3217,N_3692);
xnor U4741 (N_4741,N_3168,N_3479);
nor U4742 (N_4742,N_3788,N_3392);
and U4743 (N_4743,N_3329,N_3813);
and U4744 (N_4744,N_3032,N_3278);
and U4745 (N_4745,N_3161,N_3352);
xor U4746 (N_4746,N_3003,N_3903);
or U4747 (N_4747,N_3125,N_3223);
or U4748 (N_4748,N_3874,N_3143);
nor U4749 (N_4749,N_3666,N_3749);
nand U4750 (N_4750,N_3321,N_3221);
nand U4751 (N_4751,N_3455,N_3691);
nand U4752 (N_4752,N_3147,N_3976);
and U4753 (N_4753,N_3192,N_3175);
or U4754 (N_4754,N_3582,N_3375);
xor U4755 (N_4755,N_3001,N_3091);
and U4756 (N_4756,N_3499,N_3747);
and U4757 (N_4757,N_3567,N_3649);
nor U4758 (N_4758,N_3535,N_3537);
nand U4759 (N_4759,N_3877,N_3538);
nand U4760 (N_4760,N_3017,N_3416);
nand U4761 (N_4761,N_3210,N_3139);
xor U4762 (N_4762,N_3157,N_3022);
nor U4763 (N_4763,N_3708,N_3351);
nand U4764 (N_4764,N_3124,N_3152);
nor U4765 (N_4765,N_3073,N_3760);
nor U4766 (N_4766,N_3318,N_3048);
or U4767 (N_4767,N_3014,N_3517);
xor U4768 (N_4768,N_3613,N_3902);
nand U4769 (N_4769,N_3329,N_3533);
nand U4770 (N_4770,N_3114,N_3479);
nand U4771 (N_4771,N_3588,N_3289);
nand U4772 (N_4772,N_3858,N_3228);
and U4773 (N_4773,N_3611,N_3014);
nand U4774 (N_4774,N_3871,N_3707);
or U4775 (N_4775,N_3776,N_3457);
nor U4776 (N_4776,N_3541,N_3106);
and U4777 (N_4777,N_3635,N_3835);
or U4778 (N_4778,N_3080,N_3444);
nor U4779 (N_4779,N_3863,N_3325);
xor U4780 (N_4780,N_3929,N_3969);
and U4781 (N_4781,N_3520,N_3814);
nor U4782 (N_4782,N_3696,N_3219);
nor U4783 (N_4783,N_3662,N_3563);
xnor U4784 (N_4784,N_3016,N_3313);
nor U4785 (N_4785,N_3538,N_3454);
nand U4786 (N_4786,N_3353,N_3403);
xnor U4787 (N_4787,N_3808,N_3875);
nor U4788 (N_4788,N_3305,N_3358);
nor U4789 (N_4789,N_3379,N_3022);
xnor U4790 (N_4790,N_3153,N_3386);
xor U4791 (N_4791,N_3789,N_3161);
nor U4792 (N_4792,N_3896,N_3750);
xnor U4793 (N_4793,N_3016,N_3648);
nor U4794 (N_4794,N_3005,N_3618);
nor U4795 (N_4795,N_3715,N_3806);
and U4796 (N_4796,N_3398,N_3283);
and U4797 (N_4797,N_3678,N_3116);
nand U4798 (N_4798,N_3976,N_3771);
or U4799 (N_4799,N_3809,N_3539);
nand U4800 (N_4800,N_3684,N_3837);
nor U4801 (N_4801,N_3478,N_3354);
nand U4802 (N_4802,N_3864,N_3462);
and U4803 (N_4803,N_3107,N_3473);
xor U4804 (N_4804,N_3158,N_3942);
or U4805 (N_4805,N_3311,N_3459);
and U4806 (N_4806,N_3343,N_3604);
or U4807 (N_4807,N_3476,N_3850);
nor U4808 (N_4808,N_3788,N_3246);
nor U4809 (N_4809,N_3754,N_3442);
and U4810 (N_4810,N_3402,N_3919);
nand U4811 (N_4811,N_3040,N_3266);
and U4812 (N_4812,N_3760,N_3682);
nand U4813 (N_4813,N_3713,N_3124);
nand U4814 (N_4814,N_3278,N_3793);
xnor U4815 (N_4815,N_3768,N_3634);
nor U4816 (N_4816,N_3855,N_3566);
nand U4817 (N_4817,N_3433,N_3300);
nand U4818 (N_4818,N_3485,N_3588);
nor U4819 (N_4819,N_3558,N_3716);
and U4820 (N_4820,N_3319,N_3850);
nor U4821 (N_4821,N_3818,N_3320);
and U4822 (N_4822,N_3778,N_3215);
nand U4823 (N_4823,N_3796,N_3538);
nor U4824 (N_4824,N_3461,N_3206);
nand U4825 (N_4825,N_3389,N_3275);
or U4826 (N_4826,N_3952,N_3446);
nand U4827 (N_4827,N_3189,N_3457);
xor U4828 (N_4828,N_3088,N_3543);
nor U4829 (N_4829,N_3750,N_3385);
or U4830 (N_4830,N_3490,N_3612);
or U4831 (N_4831,N_3627,N_3695);
and U4832 (N_4832,N_3821,N_3785);
nand U4833 (N_4833,N_3814,N_3036);
nor U4834 (N_4834,N_3797,N_3264);
xor U4835 (N_4835,N_3249,N_3514);
and U4836 (N_4836,N_3428,N_3144);
nor U4837 (N_4837,N_3767,N_3986);
and U4838 (N_4838,N_3099,N_3568);
and U4839 (N_4839,N_3746,N_3601);
nor U4840 (N_4840,N_3601,N_3302);
and U4841 (N_4841,N_3920,N_3684);
nor U4842 (N_4842,N_3058,N_3880);
or U4843 (N_4843,N_3802,N_3435);
and U4844 (N_4844,N_3430,N_3093);
xnor U4845 (N_4845,N_3430,N_3705);
nor U4846 (N_4846,N_3963,N_3395);
nand U4847 (N_4847,N_3892,N_3280);
xor U4848 (N_4848,N_3618,N_3002);
nor U4849 (N_4849,N_3528,N_3999);
or U4850 (N_4850,N_3898,N_3184);
nor U4851 (N_4851,N_3620,N_3110);
or U4852 (N_4852,N_3778,N_3180);
nand U4853 (N_4853,N_3110,N_3394);
nor U4854 (N_4854,N_3247,N_3738);
xnor U4855 (N_4855,N_3791,N_3258);
or U4856 (N_4856,N_3695,N_3664);
or U4857 (N_4857,N_3444,N_3502);
nor U4858 (N_4858,N_3903,N_3923);
or U4859 (N_4859,N_3995,N_3151);
and U4860 (N_4860,N_3016,N_3924);
or U4861 (N_4861,N_3330,N_3098);
nand U4862 (N_4862,N_3337,N_3648);
nor U4863 (N_4863,N_3454,N_3946);
and U4864 (N_4864,N_3836,N_3190);
nand U4865 (N_4865,N_3949,N_3739);
xor U4866 (N_4866,N_3319,N_3177);
nor U4867 (N_4867,N_3707,N_3448);
and U4868 (N_4868,N_3979,N_3272);
xor U4869 (N_4869,N_3957,N_3540);
or U4870 (N_4870,N_3274,N_3564);
xor U4871 (N_4871,N_3925,N_3497);
xnor U4872 (N_4872,N_3599,N_3997);
xnor U4873 (N_4873,N_3077,N_3212);
xor U4874 (N_4874,N_3545,N_3481);
nor U4875 (N_4875,N_3615,N_3058);
nand U4876 (N_4876,N_3297,N_3040);
xnor U4877 (N_4877,N_3976,N_3877);
and U4878 (N_4878,N_3692,N_3864);
xor U4879 (N_4879,N_3836,N_3811);
nor U4880 (N_4880,N_3625,N_3369);
or U4881 (N_4881,N_3310,N_3622);
xor U4882 (N_4882,N_3861,N_3847);
nor U4883 (N_4883,N_3692,N_3026);
xnor U4884 (N_4884,N_3890,N_3019);
nand U4885 (N_4885,N_3580,N_3756);
nor U4886 (N_4886,N_3149,N_3073);
and U4887 (N_4887,N_3096,N_3727);
nand U4888 (N_4888,N_3024,N_3612);
nand U4889 (N_4889,N_3418,N_3248);
xnor U4890 (N_4890,N_3988,N_3737);
or U4891 (N_4891,N_3240,N_3393);
nor U4892 (N_4892,N_3387,N_3391);
xor U4893 (N_4893,N_3673,N_3666);
xnor U4894 (N_4894,N_3741,N_3410);
or U4895 (N_4895,N_3948,N_3898);
nor U4896 (N_4896,N_3958,N_3614);
or U4897 (N_4897,N_3386,N_3472);
nor U4898 (N_4898,N_3398,N_3546);
or U4899 (N_4899,N_3541,N_3372);
nand U4900 (N_4900,N_3076,N_3946);
and U4901 (N_4901,N_3049,N_3202);
and U4902 (N_4902,N_3057,N_3935);
nand U4903 (N_4903,N_3959,N_3624);
nand U4904 (N_4904,N_3081,N_3458);
nor U4905 (N_4905,N_3530,N_3083);
nor U4906 (N_4906,N_3545,N_3365);
and U4907 (N_4907,N_3177,N_3235);
nand U4908 (N_4908,N_3919,N_3000);
nand U4909 (N_4909,N_3602,N_3374);
nor U4910 (N_4910,N_3508,N_3338);
xnor U4911 (N_4911,N_3345,N_3986);
xor U4912 (N_4912,N_3696,N_3135);
nor U4913 (N_4913,N_3956,N_3478);
or U4914 (N_4914,N_3766,N_3885);
xnor U4915 (N_4915,N_3683,N_3562);
or U4916 (N_4916,N_3980,N_3862);
or U4917 (N_4917,N_3197,N_3317);
or U4918 (N_4918,N_3311,N_3729);
xnor U4919 (N_4919,N_3355,N_3672);
or U4920 (N_4920,N_3123,N_3639);
nor U4921 (N_4921,N_3841,N_3336);
nor U4922 (N_4922,N_3390,N_3718);
xnor U4923 (N_4923,N_3902,N_3456);
and U4924 (N_4924,N_3290,N_3460);
and U4925 (N_4925,N_3132,N_3386);
nor U4926 (N_4926,N_3423,N_3910);
or U4927 (N_4927,N_3725,N_3398);
nand U4928 (N_4928,N_3579,N_3833);
or U4929 (N_4929,N_3812,N_3853);
or U4930 (N_4930,N_3983,N_3729);
nand U4931 (N_4931,N_3063,N_3423);
or U4932 (N_4932,N_3478,N_3986);
nand U4933 (N_4933,N_3743,N_3930);
and U4934 (N_4934,N_3826,N_3035);
and U4935 (N_4935,N_3886,N_3695);
nor U4936 (N_4936,N_3485,N_3625);
xor U4937 (N_4937,N_3307,N_3267);
and U4938 (N_4938,N_3900,N_3242);
nand U4939 (N_4939,N_3072,N_3779);
nor U4940 (N_4940,N_3842,N_3832);
and U4941 (N_4941,N_3061,N_3484);
or U4942 (N_4942,N_3694,N_3851);
and U4943 (N_4943,N_3458,N_3201);
nand U4944 (N_4944,N_3627,N_3354);
xnor U4945 (N_4945,N_3711,N_3344);
and U4946 (N_4946,N_3954,N_3499);
xor U4947 (N_4947,N_3723,N_3191);
nor U4948 (N_4948,N_3567,N_3381);
nand U4949 (N_4949,N_3305,N_3111);
or U4950 (N_4950,N_3713,N_3028);
nor U4951 (N_4951,N_3203,N_3220);
nor U4952 (N_4952,N_3407,N_3943);
nor U4953 (N_4953,N_3481,N_3161);
xnor U4954 (N_4954,N_3853,N_3917);
or U4955 (N_4955,N_3902,N_3861);
nor U4956 (N_4956,N_3582,N_3211);
nand U4957 (N_4957,N_3642,N_3716);
and U4958 (N_4958,N_3135,N_3213);
xnor U4959 (N_4959,N_3774,N_3315);
nand U4960 (N_4960,N_3710,N_3122);
nand U4961 (N_4961,N_3334,N_3550);
and U4962 (N_4962,N_3450,N_3234);
xor U4963 (N_4963,N_3584,N_3379);
and U4964 (N_4964,N_3027,N_3797);
xnor U4965 (N_4965,N_3402,N_3450);
or U4966 (N_4966,N_3279,N_3557);
nand U4967 (N_4967,N_3631,N_3589);
or U4968 (N_4968,N_3785,N_3029);
nor U4969 (N_4969,N_3351,N_3923);
nor U4970 (N_4970,N_3177,N_3602);
and U4971 (N_4971,N_3907,N_3352);
nor U4972 (N_4972,N_3594,N_3266);
xnor U4973 (N_4973,N_3897,N_3747);
or U4974 (N_4974,N_3515,N_3145);
or U4975 (N_4975,N_3631,N_3369);
and U4976 (N_4976,N_3947,N_3530);
xor U4977 (N_4977,N_3022,N_3679);
nor U4978 (N_4978,N_3579,N_3720);
xor U4979 (N_4979,N_3047,N_3845);
xor U4980 (N_4980,N_3339,N_3000);
nor U4981 (N_4981,N_3803,N_3907);
nand U4982 (N_4982,N_3129,N_3505);
nor U4983 (N_4983,N_3373,N_3158);
or U4984 (N_4984,N_3636,N_3946);
nor U4985 (N_4985,N_3832,N_3626);
xor U4986 (N_4986,N_3307,N_3386);
xnor U4987 (N_4987,N_3020,N_3744);
or U4988 (N_4988,N_3681,N_3522);
or U4989 (N_4989,N_3526,N_3173);
nand U4990 (N_4990,N_3392,N_3176);
and U4991 (N_4991,N_3608,N_3957);
nand U4992 (N_4992,N_3414,N_3083);
or U4993 (N_4993,N_3235,N_3058);
nor U4994 (N_4994,N_3502,N_3584);
nor U4995 (N_4995,N_3198,N_3093);
and U4996 (N_4996,N_3692,N_3096);
nor U4997 (N_4997,N_3885,N_3274);
nor U4998 (N_4998,N_3219,N_3919);
and U4999 (N_4999,N_3082,N_3908);
nor UO_0 (O_0,N_4061,N_4516);
nor UO_1 (O_1,N_4490,N_4628);
nor UO_2 (O_2,N_4190,N_4481);
and UO_3 (O_3,N_4992,N_4099);
or UO_4 (O_4,N_4984,N_4145);
or UO_5 (O_5,N_4565,N_4188);
xor UO_6 (O_6,N_4557,N_4045);
xnor UO_7 (O_7,N_4588,N_4892);
nor UO_8 (O_8,N_4851,N_4907);
xnor UO_9 (O_9,N_4801,N_4040);
or UO_10 (O_10,N_4142,N_4574);
xor UO_11 (O_11,N_4670,N_4784);
or UO_12 (O_12,N_4882,N_4407);
or UO_13 (O_13,N_4775,N_4589);
nor UO_14 (O_14,N_4173,N_4251);
nand UO_15 (O_15,N_4300,N_4870);
nor UO_16 (O_16,N_4413,N_4336);
nand UO_17 (O_17,N_4414,N_4608);
and UO_18 (O_18,N_4742,N_4046);
nand UO_19 (O_19,N_4586,N_4053);
nand UO_20 (O_20,N_4397,N_4858);
and UO_21 (O_21,N_4845,N_4576);
nor UO_22 (O_22,N_4301,N_4920);
and UO_23 (O_23,N_4482,N_4506);
xnor UO_24 (O_24,N_4857,N_4750);
nand UO_25 (O_25,N_4860,N_4613);
nor UO_26 (O_26,N_4991,N_4060);
nand UO_27 (O_27,N_4694,N_4368);
or UO_28 (O_28,N_4513,N_4256);
and UO_29 (O_29,N_4098,N_4151);
or UO_30 (O_30,N_4197,N_4620);
nor UO_31 (O_31,N_4957,N_4401);
nand UO_32 (O_32,N_4463,N_4829);
and UO_33 (O_33,N_4824,N_4417);
nand UO_34 (O_34,N_4938,N_4479);
and UO_35 (O_35,N_4720,N_4459);
nand UO_36 (O_36,N_4484,N_4217);
nor UO_37 (O_37,N_4525,N_4290);
xnor UO_38 (O_38,N_4929,N_4715);
and UO_39 (O_39,N_4621,N_4392);
nand UO_40 (O_40,N_4675,N_4949);
nand UO_41 (O_41,N_4140,N_4765);
or UO_42 (O_42,N_4072,N_4073);
and UO_43 (O_43,N_4844,N_4612);
and UO_44 (O_44,N_4426,N_4822);
nor UO_45 (O_45,N_4286,N_4896);
nand UO_46 (O_46,N_4831,N_4402);
nor UO_47 (O_47,N_4315,N_4123);
or UO_48 (O_48,N_4320,N_4657);
or UO_49 (O_49,N_4186,N_4755);
nor UO_50 (O_50,N_4213,N_4967);
or UO_51 (O_51,N_4406,N_4554);
or UO_52 (O_52,N_4867,N_4661);
and UO_53 (O_53,N_4356,N_4686);
nand UO_54 (O_54,N_4924,N_4909);
nor UO_55 (O_55,N_4989,N_4887);
nand UO_56 (O_56,N_4047,N_4718);
and UO_57 (O_57,N_4044,N_4833);
or UO_58 (O_58,N_4489,N_4161);
and UO_59 (O_59,N_4879,N_4550);
xnor UO_60 (O_60,N_4185,N_4637);
nand UO_61 (O_61,N_4841,N_4773);
or UO_62 (O_62,N_4312,N_4629);
and UO_63 (O_63,N_4225,N_4010);
xor UO_64 (O_64,N_4708,N_4423);
nand UO_65 (O_65,N_4601,N_4243);
xor UO_66 (O_66,N_4253,N_4355);
or UO_67 (O_67,N_4241,N_4314);
nor UO_68 (O_68,N_4931,N_4208);
xor UO_69 (O_69,N_4227,N_4587);
or UO_70 (O_70,N_4446,N_4058);
and UO_71 (O_71,N_4485,N_4088);
or UO_72 (O_72,N_4902,N_4597);
and UO_73 (O_73,N_4619,N_4007);
xor UO_74 (O_74,N_4877,N_4937);
and UO_75 (O_75,N_4859,N_4034);
nor UO_76 (O_76,N_4714,N_4561);
and UO_77 (O_77,N_4215,N_4717);
or UO_78 (O_78,N_4032,N_4043);
nand UO_79 (O_79,N_4460,N_4434);
nand UO_80 (O_80,N_4329,N_4530);
xnor UO_81 (O_81,N_4848,N_4299);
nor UO_82 (O_82,N_4359,N_4507);
nand UO_83 (O_83,N_4156,N_4866);
and UO_84 (O_84,N_4131,N_4529);
nor UO_85 (O_85,N_4239,N_4634);
or UO_86 (O_86,N_4326,N_4966);
nor UO_87 (O_87,N_4526,N_4724);
or UO_88 (O_88,N_4263,N_4664);
or UO_89 (O_89,N_4956,N_4927);
nor UO_90 (O_90,N_4093,N_4900);
nor UO_91 (O_91,N_4112,N_4672);
or UO_92 (O_92,N_4693,N_4248);
xor UO_93 (O_93,N_4182,N_4497);
xor UO_94 (O_94,N_4050,N_4415);
nand UO_95 (O_95,N_4195,N_4030);
or UO_96 (O_96,N_4847,N_4642);
nor UO_97 (O_97,N_4996,N_4184);
nand UO_98 (O_98,N_4081,N_4641);
nor UO_99 (O_99,N_4494,N_4635);
xor UO_100 (O_100,N_4805,N_4566);
or UO_101 (O_101,N_4676,N_4932);
or UO_102 (O_102,N_4157,N_4544);
and UO_103 (O_103,N_4362,N_4262);
or UO_104 (O_104,N_4654,N_4761);
nand UO_105 (O_105,N_4653,N_4796);
xnor UO_106 (O_106,N_4204,N_4436);
nor UO_107 (O_107,N_4881,N_4577);
nand UO_108 (O_108,N_4293,N_4175);
nor UO_109 (O_109,N_4656,N_4055);
or UO_110 (O_110,N_4644,N_4449);
nor UO_111 (O_111,N_4370,N_4291);
nand UO_112 (O_112,N_4158,N_4385);
nand UO_113 (O_113,N_4639,N_4816);
nor UO_114 (O_114,N_4679,N_4220);
and UO_115 (O_115,N_4268,N_4977);
xor UO_116 (O_116,N_4535,N_4607);
nor UO_117 (O_117,N_4994,N_4071);
xnor UO_118 (O_118,N_4770,N_4231);
nand UO_119 (O_119,N_4008,N_4074);
nor UO_120 (O_120,N_4458,N_4905);
or UO_121 (O_121,N_4467,N_4662);
xnor UO_122 (O_122,N_4687,N_4108);
nand UO_123 (O_123,N_4849,N_4187);
xnor UO_124 (O_124,N_4940,N_4183);
and UO_125 (O_125,N_4165,N_4842);
or UO_126 (O_126,N_4101,N_4017);
and UO_127 (O_127,N_4563,N_4180);
nor UO_128 (O_128,N_4104,N_4983);
xnor UO_129 (O_129,N_4224,N_4388);
and UO_130 (O_130,N_4424,N_4429);
nand UO_131 (O_131,N_4511,N_4432);
nor UO_132 (O_132,N_4127,N_4440);
nor UO_133 (O_133,N_4351,N_4015);
or UO_134 (O_134,N_4020,N_4421);
xor UO_135 (O_135,N_4404,N_4310);
and UO_136 (O_136,N_4332,N_4042);
nand UO_137 (O_137,N_4166,N_4539);
nand UO_138 (O_138,N_4762,N_4922);
or UO_139 (O_139,N_4084,N_4939);
nor UO_140 (O_140,N_4874,N_4041);
nor UO_141 (O_141,N_4825,N_4033);
or UO_142 (O_142,N_4153,N_4681);
xnor UO_143 (O_143,N_4083,N_4445);
and UO_144 (O_144,N_4431,N_4000);
and UO_145 (O_145,N_4496,N_4119);
or UO_146 (O_146,N_4056,N_4592);
or UO_147 (O_147,N_4371,N_4699);
nor UO_148 (O_148,N_4502,N_4547);
nor UO_149 (O_149,N_4945,N_4505);
or UO_150 (O_150,N_4752,N_4384);
xor UO_151 (O_151,N_4466,N_4111);
xor UO_152 (O_152,N_4154,N_4982);
xor UO_153 (O_153,N_4673,N_4645);
or UO_154 (O_154,N_4082,N_4680);
xor UO_155 (O_155,N_4935,N_4564);
nor UO_156 (O_156,N_4808,N_4028);
nor UO_157 (O_157,N_4521,N_4249);
xor UO_158 (O_158,N_4361,N_4572);
or UO_159 (O_159,N_4124,N_4289);
or UO_160 (O_160,N_4660,N_4418);
or UO_161 (O_161,N_4791,N_4476);
nor UO_162 (O_162,N_4094,N_4039);
xnor UO_163 (O_163,N_4692,N_4345);
and UO_164 (O_164,N_4631,N_4487);
xnor UO_165 (O_165,N_4986,N_4096);
or UO_166 (O_166,N_4735,N_4541);
and UO_167 (O_167,N_4579,N_4194);
xor UO_168 (O_168,N_4258,N_4843);
xnor UO_169 (O_169,N_4170,N_4760);
nand UO_170 (O_170,N_4504,N_4177);
or UO_171 (O_171,N_4500,N_4317);
nand UO_172 (O_172,N_4223,N_4558);
and UO_173 (O_173,N_4780,N_4917);
nand UO_174 (O_174,N_4854,N_4062);
xnor UO_175 (O_175,N_4545,N_4453);
or UO_176 (O_176,N_4528,N_4582);
or UO_177 (O_177,N_4292,N_4149);
nor UO_178 (O_178,N_4281,N_4609);
and UO_179 (O_179,N_4830,N_4865);
nor UO_180 (O_180,N_4958,N_4234);
xor UO_181 (O_181,N_4856,N_4520);
nand UO_182 (O_182,N_4553,N_4988);
or UO_183 (O_183,N_4396,N_4552);
nand UO_184 (O_184,N_4075,N_4677);
or UO_185 (O_185,N_4340,N_4538);
nand UO_186 (O_186,N_4428,N_4583);
nor UO_187 (O_187,N_4238,N_4269);
xor UO_188 (O_188,N_4560,N_4943);
and UO_189 (O_189,N_4493,N_4369);
nor UO_190 (O_190,N_4115,N_4952);
and UO_191 (O_191,N_4420,N_4668);
nand UO_192 (O_192,N_4176,N_4793);
nor UO_193 (O_193,N_4985,N_4596);
nand UO_194 (O_194,N_4737,N_4897);
xnor UO_195 (O_195,N_4978,N_4972);
nor UO_196 (O_196,N_4973,N_4462);
xor UO_197 (O_197,N_4132,N_4029);
or UO_198 (O_198,N_4953,N_4105);
nand UO_199 (O_199,N_4838,N_4107);
nor UO_200 (O_200,N_4390,N_4834);
and UO_201 (O_201,N_4019,N_4797);
or UO_202 (O_202,N_4103,N_4210);
nand UO_203 (O_203,N_4556,N_4230);
nand UO_204 (O_204,N_4001,N_4610);
nor UO_205 (O_205,N_4261,N_4378);
and UO_206 (O_206,N_4265,N_4734);
or UO_207 (O_207,N_4522,N_4051);
nor UO_208 (O_208,N_4454,N_4193);
nand UO_209 (O_209,N_4080,N_4813);
and UO_210 (O_210,N_4990,N_4199);
nor UO_211 (O_211,N_4947,N_4551);
nand UO_212 (O_212,N_4002,N_4643);
nand UO_213 (O_213,N_4085,N_4005);
xor UO_214 (O_214,N_4562,N_4179);
nor UO_215 (O_215,N_4471,N_4214);
or UO_216 (O_216,N_4191,N_4745);
or UO_217 (O_217,N_4744,N_4581);
and UO_218 (O_218,N_4658,N_4035);
xor UO_219 (O_219,N_4114,N_4221);
nor UO_220 (O_220,N_4143,N_4405);
or UO_221 (O_221,N_4871,N_4321);
nand UO_222 (O_222,N_4965,N_4725);
xor UO_223 (O_223,N_4537,N_4893);
nor UO_224 (O_224,N_4655,N_4517);
and UO_225 (O_225,N_4646,N_4515);
nand UO_226 (O_226,N_4409,N_4669);
xor UO_227 (O_227,N_4478,N_4995);
or UO_228 (O_228,N_4910,N_4349);
xnor UO_229 (O_229,N_4855,N_4955);
xor UO_230 (O_230,N_4707,N_4323);
xor UO_231 (O_231,N_4689,N_4357);
or UO_232 (O_232,N_4721,N_4732);
or UO_233 (O_233,N_4064,N_4331);
nor UO_234 (O_234,N_4264,N_4534);
nor UO_235 (O_235,N_4287,N_4171);
nor UO_236 (O_236,N_4393,N_4278);
and UO_237 (O_237,N_4852,N_4026);
or UO_238 (O_238,N_4363,N_4811);
xor UO_239 (O_239,N_4727,N_4219);
or UO_240 (O_240,N_4303,N_4800);
or UO_241 (O_241,N_4951,N_4086);
or UO_242 (O_242,N_4782,N_4942);
xnor UO_243 (O_243,N_4884,N_4804);
nor UO_244 (O_244,N_4928,N_4569);
and UO_245 (O_245,N_4464,N_4309);
xnor UO_246 (O_246,N_4704,N_4850);
nor UO_247 (O_247,N_4751,N_4280);
nand UO_248 (O_248,N_4139,N_4427);
nor UO_249 (O_249,N_4394,N_4348);
or UO_250 (O_250,N_4013,N_4063);
nor UO_251 (O_251,N_4381,N_4970);
nand UO_252 (O_252,N_4398,N_4270);
or UO_253 (O_253,N_4508,N_4523);
nor UO_254 (O_254,N_4004,N_4792);
or UO_255 (O_255,N_4731,N_4283);
nand UO_256 (O_256,N_4366,N_4106);
xor UO_257 (O_257,N_4469,N_4533);
nor UO_258 (O_258,N_4488,N_4766);
nand UO_259 (O_259,N_4350,N_4048);
or UO_260 (O_260,N_4665,N_4736);
nor UO_261 (O_261,N_4546,N_4135);
xnor UO_262 (O_262,N_4772,N_4695);
or UO_263 (O_263,N_4781,N_4324);
nor UO_264 (O_264,N_4590,N_4712);
and UO_265 (O_265,N_4122,N_4452);
nand UO_266 (O_266,N_4531,N_4120);
or UO_267 (O_267,N_4740,N_4486);
nor UO_268 (O_268,N_4383,N_4906);
nor UO_269 (O_269,N_4457,N_4330);
or UO_270 (O_270,N_4981,N_4810);
xnor UO_271 (O_271,N_4443,N_4031);
nand UO_272 (O_272,N_4726,N_4748);
and UO_273 (O_273,N_4244,N_4647);
and UO_274 (O_274,N_4618,N_4311);
xor UO_275 (O_275,N_4503,N_4444);
or UO_276 (O_276,N_4602,N_4974);
nand UO_277 (O_277,N_4778,N_4276);
xnor UO_278 (O_278,N_4364,N_4174);
nor UO_279 (O_279,N_4162,N_4701);
and UO_280 (O_280,N_4730,N_4092);
nor UO_281 (O_281,N_4211,N_4163);
xnor UO_282 (O_282,N_4456,N_4820);
xnor UO_283 (O_283,N_4322,N_4279);
or UO_284 (O_284,N_4437,N_4993);
xnor UO_285 (O_285,N_4192,N_4671);
xnor UO_286 (O_286,N_4438,N_4483);
xor UO_287 (O_287,N_4894,N_4346);
xor UO_288 (O_288,N_4284,N_4594);
nor UO_289 (O_289,N_4763,N_4136);
and UO_290 (O_290,N_4749,N_4450);
and UO_291 (O_291,N_4201,N_4605);
xor UO_292 (O_292,N_4304,N_4768);
xnor UO_293 (O_293,N_4172,N_4254);
or UO_294 (O_294,N_4117,N_4963);
xor UO_295 (O_295,N_4872,N_4237);
or UO_296 (O_296,N_4786,N_4069);
nand UO_297 (O_297,N_4059,N_4089);
and UO_298 (O_298,N_4433,N_4313);
xnor UO_299 (O_299,N_4767,N_4674);
nand UO_300 (O_300,N_4626,N_4918);
and UO_301 (O_301,N_4509,N_4477);
or UO_302 (O_302,N_4295,N_4367);
or UO_303 (O_303,N_4876,N_4719);
nor UO_304 (O_304,N_4713,N_4698);
nor UO_305 (O_305,N_4138,N_4376);
nor UO_306 (O_306,N_4474,N_4235);
or UO_307 (O_307,N_4307,N_4391);
or UO_308 (O_308,N_4997,N_4152);
and UO_309 (O_309,N_4333,N_4435);
and UO_310 (O_310,N_4196,N_4022);
nor UO_311 (O_311,N_4400,N_4743);
nor UO_312 (O_312,N_4288,N_4389);
nor UO_313 (O_313,N_4787,N_4422);
nor UO_314 (O_314,N_4116,N_4473);
and UO_315 (O_315,N_4416,N_4568);
nand UO_316 (O_316,N_4595,N_4373);
and UO_317 (O_317,N_4794,N_4334);
nor UO_318 (O_318,N_4979,N_4944);
nor UO_319 (O_319,N_4627,N_4441);
or UO_320 (O_320,N_4439,N_4711);
or UO_321 (O_321,N_4964,N_4571);
nand UO_322 (O_322,N_4512,N_4222);
nor UO_323 (O_323,N_4746,N_4144);
and UO_324 (O_324,N_4226,N_4267);
nand UO_325 (O_325,N_4954,N_4129);
nand UO_326 (O_326,N_4764,N_4066);
nor UO_327 (O_327,N_4987,N_4738);
xor UO_328 (O_328,N_4710,N_4246);
nand UO_329 (O_329,N_4853,N_4837);
and UO_330 (O_330,N_4683,N_4347);
nand UO_331 (O_331,N_4372,N_4861);
or UO_332 (O_332,N_4169,N_4663);
nand UO_333 (O_333,N_4442,N_4065);
or UO_334 (O_334,N_4475,N_4828);
and UO_335 (O_335,N_4339,N_4492);
nor UO_336 (O_336,N_4798,N_4408);
nand UO_337 (O_337,N_4294,N_4023);
or UO_338 (O_338,N_4913,N_4411);
xnor UO_339 (O_339,N_4499,N_4819);
and UO_340 (O_340,N_4790,N_4016);
or UO_341 (O_341,N_4395,N_4250);
nor UO_342 (O_342,N_4277,N_4926);
and UO_343 (O_343,N_4011,N_4399);
and UO_344 (O_344,N_4899,N_4980);
xnor UO_345 (O_345,N_4448,N_4232);
nand UO_346 (O_346,N_4150,N_4818);
and UO_347 (O_347,N_4919,N_4216);
and UO_348 (O_348,N_4134,N_4341);
xnor UO_349 (O_349,N_4971,N_4969);
or UO_350 (O_350,N_4836,N_4527);
or UO_351 (O_351,N_4159,N_4617);
xnor UO_352 (O_352,N_4883,N_4319);
nand UO_353 (O_353,N_4480,N_4864);
nand UO_354 (O_354,N_4110,N_4916);
nor UO_355 (O_355,N_4090,N_4133);
xnor UO_356 (O_356,N_4189,N_4832);
or UO_357 (O_357,N_4274,N_4206);
and UO_358 (O_358,N_4252,N_4706);
nor UO_359 (O_359,N_4946,N_4360);
nand UO_360 (O_360,N_4147,N_4343);
nand UO_361 (O_361,N_4869,N_4109);
nand UO_362 (O_362,N_4638,N_4891);
nor UO_363 (O_363,N_4585,N_4815);
or UO_364 (O_364,N_4593,N_4999);
or UO_365 (O_365,N_4968,N_4904);
nor UO_366 (O_366,N_4901,N_4976);
nand UO_367 (O_367,N_4624,N_4959);
nor UO_368 (O_368,N_4769,N_4911);
and UO_369 (O_369,N_4275,N_4247);
or UO_370 (O_370,N_4447,N_4455);
xor UO_371 (O_371,N_4076,N_4014);
nor UO_372 (O_372,N_4067,N_4282);
nor UO_373 (O_373,N_4961,N_4728);
nand UO_374 (O_374,N_4302,N_4614);
nor UO_375 (O_375,N_4148,N_4603);
nor UO_376 (O_376,N_4049,N_4057);
and UO_377 (O_377,N_4691,N_4242);
xor UO_378 (O_378,N_4164,N_4203);
and UO_379 (O_379,N_4501,N_4933);
xor UO_380 (O_380,N_4412,N_4685);
xnor UO_381 (O_381,N_4365,N_4739);
nor UO_382 (O_382,N_4233,N_4078);
xnor UO_383 (O_383,N_4705,N_4578);
and UO_384 (O_384,N_4121,N_4025);
xnor UO_385 (O_385,N_4344,N_4925);
nand UO_386 (O_386,N_4325,N_4377);
nand UO_387 (O_387,N_4652,N_4354);
or UO_388 (O_388,N_4759,N_4868);
xnor UO_389 (O_389,N_4316,N_4630);
and UO_390 (O_390,N_4379,N_4255);
xnor UO_391 (O_391,N_4783,N_4141);
xor UO_392 (O_392,N_4812,N_4651);
or UO_393 (O_393,N_4606,N_4753);
nor UO_394 (O_394,N_4068,N_4155);
or UO_395 (O_395,N_4102,N_4198);
xor UO_396 (O_396,N_4305,N_4875);
nor UO_397 (O_397,N_4690,N_4636);
nor UO_398 (O_398,N_4809,N_4702);
xnor UO_399 (O_399,N_4741,N_4684);
and UO_400 (O_400,N_4495,N_4077);
nand UO_401 (O_401,N_4259,N_4789);
and UO_402 (O_402,N_4375,N_4009);
nor UO_403 (O_403,N_4327,N_4666);
nand UO_404 (O_404,N_4018,N_4491);
or UO_405 (O_405,N_4168,N_4430);
and UO_406 (O_406,N_4598,N_4229);
xor UO_407 (O_407,N_4387,N_4633);
nand UO_408 (O_408,N_4353,N_4205);
or UO_409 (O_409,N_4567,N_4342);
xnor UO_410 (O_410,N_4839,N_4202);
or UO_411 (O_411,N_4532,N_4930);
or UO_412 (O_412,N_4200,N_4510);
or UO_413 (O_413,N_4054,N_4024);
and UO_414 (O_414,N_4659,N_4650);
nor UO_415 (O_415,N_4540,N_4468);
and UO_416 (O_416,N_4840,N_4543);
xor UO_417 (O_417,N_4632,N_4260);
xor UO_418 (O_418,N_4688,N_4465);
nor UO_419 (O_419,N_4880,N_4318);
nand UO_420 (O_420,N_4814,N_4137);
nand UO_421 (O_421,N_4052,N_4682);
or UO_422 (O_422,N_4006,N_4079);
xor UO_423 (O_423,N_4903,N_4885);
xor UO_424 (O_424,N_4898,N_4771);
nor UO_425 (O_425,N_4027,N_4962);
nor UO_426 (O_426,N_4095,N_4306);
and UO_427 (O_427,N_4273,N_4756);
nor UO_428 (O_428,N_4754,N_4950);
or UO_429 (O_429,N_4498,N_4236);
nor UO_430 (O_430,N_4130,N_4451);
or UO_431 (O_431,N_4519,N_4113);
or UO_432 (O_432,N_4779,N_4625);
or UO_433 (O_433,N_4722,N_4298);
nand UO_434 (O_434,N_4616,N_4228);
nor UO_435 (O_435,N_4806,N_4285);
xnor UO_436 (O_436,N_4678,N_4873);
and UO_437 (O_437,N_4700,N_4863);
nor UO_438 (O_438,N_4272,N_4788);
nor UO_439 (O_439,N_4817,N_4998);
nor UO_440 (O_440,N_4716,N_4821);
nand UO_441 (O_441,N_4380,N_4549);
nor UO_442 (O_442,N_4559,N_4697);
nor UO_443 (O_443,N_4126,N_4245);
xnor UO_444 (O_444,N_4948,N_4723);
and UO_445 (O_445,N_4070,N_4648);
or UO_446 (O_446,N_4886,N_4623);
and UO_447 (O_447,N_4012,N_4036);
nor UO_448 (O_448,N_4923,N_4758);
and UO_449 (O_449,N_4799,N_4374);
or UO_450 (O_450,N_4240,N_4097);
nand UO_451 (O_451,N_4352,N_4795);
nand UO_452 (O_452,N_4461,N_4146);
and UO_453 (O_453,N_4386,N_4555);
or UO_454 (O_454,N_4733,N_4472);
and UO_455 (O_455,N_4167,N_4615);
or UO_456 (O_456,N_4003,N_4181);
nor UO_457 (O_457,N_4709,N_4580);
and UO_458 (O_458,N_4308,N_4328);
nor UO_459 (O_459,N_4912,N_4803);
or UO_460 (O_460,N_4835,N_4846);
nand UO_461 (O_461,N_4297,N_4575);
nand UO_462 (O_462,N_4862,N_4209);
or UO_463 (O_463,N_4890,N_4827);
or UO_464 (O_464,N_4747,N_4640);
nand UO_465 (O_465,N_4021,N_4570);
nor UO_466 (O_466,N_4960,N_4038);
and UO_467 (O_467,N_4908,N_4337);
or UO_468 (O_468,N_4037,N_4703);
or UO_469 (O_469,N_4785,N_4777);
nor UO_470 (O_470,N_4212,N_4178);
xor UO_471 (O_471,N_4802,N_4921);
nor UO_472 (O_472,N_4128,N_4358);
nand UO_473 (O_473,N_4125,N_4667);
or UO_474 (O_474,N_4599,N_4604);
nand UO_475 (O_475,N_4403,N_4338);
nor UO_476 (O_476,N_4518,N_4941);
nand UO_477 (O_477,N_4696,N_4878);
and UO_478 (O_478,N_4524,N_4915);
nand UO_479 (O_479,N_4382,N_4271);
xor UO_480 (O_480,N_4622,N_4611);
nor UO_481 (O_481,N_4207,N_4591);
and UO_482 (O_482,N_4807,N_4934);
and UO_483 (O_483,N_4584,N_4757);
nand UO_484 (O_484,N_4649,N_4914);
and UO_485 (O_485,N_4536,N_4470);
nor UO_486 (O_486,N_4514,N_4218);
xnor UO_487 (O_487,N_4296,N_4160);
xor UO_488 (O_488,N_4573,N_4419);
and UO_489 (O_489,N_4548,N_4888);
xor UO_490 (O_490,N_4774,N_4889);
and UO_491 (O_491,N_4091,N_4118);
nor UO_492 (O_492,N_4600,N_4266);
nand UO_493 (O_493,N_4895,N_4087);
nor UO_494 (O_494,N_4100,N_4823);
or UO_495 (O_495,N_4936,N_4729);
or UO_496 (O_496,N_4776,N_4826);
nand UO_497 (O_497,N_4542,N_4335);
and UO_498 (O_498,N_4425,N_4975);
or UO_499 (O_499,N_4257,N_4410);
nor UO_500 (O_500,N_4696,N_4746);
and UO_501 (O_501,N_4711,N_4747);
nand UO_502 (O_502,N_4415,N_4551);
and UO_503 (O_503,N_4998,N_4774);
nand UO_504 (O_504,N_4263,N_4127);
nand UO_505 (O_505,N_4662,N_4320);
nor UO_506 (O_506,N_4215,N_4122);
xor UO_507 (O_507,N_4286,N_4158);
nor UO_508 (O_508,N_4701,N_4991);
and UO_509 (O_509,N_4977,N_4132);
nor UO_510 (O_510,N_4702,N_4057);
nand UO_511 (O_511,N_4949,N_4959);
or UO_512 (O_512,N_4333,N_4613);
and UO_513 (O_513,N_4866,N_4129);
nand UO_514 (O_514,N_4124,N_4464);
and UO_515 (O_515,N_4315,N_4568);
nand UO_516 (O_516,N_4749,N_4455);
nand UO_517 (O_517,N_4293,N_4265);
nor UO_518 (O_518,N_4425,N_4078);
and UO_519 (O_519,N_4562,N_4064);
and UO_520 (O_520,N_4403,N_4256);
and UO_521 (O_521,N_4896,N_4517);
nor UO_522 (O_522,N_4885,N_4450);
nor UO_523 (O_523,N_4954,N_4628);
or UO_524 (O_524,N_4081,N_4516);
nand UO_525 (O_525,N_4272,N_4065);
nand UO_526 (O_526,N_4903,N_4327);
and UO_527 (O_527,N_4038,N_4972);
nand UO_528 (O_528,N_4294,N_4257);
xor UO_529 (O_529,N_4753,N_4820);
xnor UO_530 (O_530,N_4157,N_4398);
xnor UO_531 (O_531,N_4082,N_4092);
xor UO_532 (O_532,N_4787,N_4733);
xnor UO_533 (O_533,N_4495,N_4445);
and UO_534 (O_534,N_4834,N_4790);
nand UO_535 (O_535,N_4463,N_4278);
xor UO_536 (O_536,N_4873,N_4279);
or UO_537 (O_537,N_4535,N_4589);
nand UO_538 (O_538,N_4845,N_4101);
and UO_539 (O_539,N_4308,N_4709);
nor UO_540 (O_540,N_4880,N_4324);
and UO_541 (O_541,N_4707,N_4052);
xnor UO_542 (O_542,N_4349,N_4603);
or UO_543 (O_543,N_4411,N_4816);
or UO_544 (O_544,N_4515,N_4598);
or UO_545 (O_545,N_4523,N_4177);
nor UO_546 (O_546,N_4981,N_4879);
xor UO_547 (O_547,N_4114,N_4370);
nand UO_548 (O_548,N_4927,N_4740);
nand UO_549 (O_549,N_4779,N_4796);
nor UO_550 (O_550,N_4296,N_4264);
or UO_551 (O_551,N_4645,N_4311);
nand UO_552 (O_552,N_4660,N_4200);
nor UO_553 (O_553,N_4506,N_4526);
nand UO_554 (O_554,N_4378,N_4151);
or UO_555 (O_555,N_4420,N_4480);
or UO_556 (O_556,N_4405,N_4997);
xnor UO_557 (O_557,N_4265,N_4508);
and UO_558 (O_558,N_4393,N_4648);
and UO_559 (O_559,N_4600,N_4746);
or UO_560 (O_560,N_4763,N_4298);
nand UO_561 (O_561,N_4705,N_4854);
nor UO_562 (O_562,N_4402,N_4154);
and UO_563 (O_563,N_4954,N_4683);
and UO_564 (O_564,N_4719,N_4576);
xnor UO_565 (O_565,N_4786,N_4665);
or UO_566 (O_566,N_4805,N_4372);
or UO_567 (O_567,N_4018,N_4950);
xor UO_568 (O_568,N_4869,N_4395);
xnor UO_569 (O_569,N_4927,N_4091);
nor UO_570 (O_570,N_4836,N_4116);
nand UO_571 (O_571,N_4162,N_4916);
xnor UO_572 (O_572,N_4994,N_4025);
xnor UO_573 (O_573,N_4660,N_4196);
and UO_574 (O_574,N_4595,N_4950);
or UO_575 (O_575,N_4996,N_4096);
xnor UO_576 (O_576,N_4991,N_4986);
xor UO_577 (O_577,N_4342,N_4945);
or UO_578 (O_578,N_4511,N_4329);
nor UO_579 (O_579,N_4519,N_4128);
xor UO_580 (O_580,N_4191,N_4098);
or UO_581 (O_581,N_4001,N_4003);
or UO_582 (O_582,N_4027,N_4888);
xnor UO_583 (O_583,N_4137,N_4876);
or UO_584 (O_584,N_4940,N_4988);
xor UO_585 (O_585,N_4843,N_4817);
and UO_586 (O_586,N_4860,N_4462);
or UO_587 (O_587,N_4346,N_4193);
or UO_588 (O_588,N_4702,N_4461);
and UO_589 (O_589,N_4471,N_4114);
nand UO_590 (O_590,N_4559,N_4781);
nor UO_591 (O_591,N_4483,N_4070);
nor UO_592 (O_592,N_4639,N_4838);
and UO_593 (O_593,N_4231,N_4037);
xor UO_594 (O_594,N_4185,N_4172);
nand UO_595 (O_595,N_4066,N_4917);
nor UO_596 (O_596,N_4959,N_4958);
xor UO_597 (O_597,N_4583,N_4419);
xnor UO_598 (O_598,N_4029,N_4957);
and UO_599 (O_599,N_4656,N_4179);
or UO_600 (O_600,N_4803,N_4725);
nand UO_601 (O_601,N_4457,N_4166);
nand UO_602 (O_602,N_4333,N_4852);
nor UO_603 (O_603,N_4079,N_4250);
and UO_604 (O_604,N_4150,N_4645);
and UO_605 (O_605,N_4297,N_4377);
nand UO_606 (O_606,N_4544,N_4467);
and UO_607 (O_607,N_4194,N_4204);
and UO_608 (O_608,N_4556,N_4131);
nor UO_609 (O_609,N_4462,N_4885);
nor UO_610 (O_610,N_4207,N_4883);
and UO_611 (O_611,N_4649,N_4819);
and UO_612 (O_612,N_4911,N_4509);
xnor UO_613 (O_613,N_4553,N_4790);
nand UO_614 (O_614,N_4838,N_4417);
and UO_615 (O_615,N_4229,N_4042);
and UO_616 (O_616,N_4052,N_4825);
nand UO_617 (O_617,N_4097,N_4803);
xnor UO_618 (O_618,N_4655,N_4057);
and UO_619 (O_619,N_4917,N_4627);
and UO_620 (O_620,N_4887,N_4190);
nand UO_621 (O_621,N_4682,N_4584);
or UO_622 (O_622,N_4779,N_4304);
xor UO_623 (O_623,N_4243,N_4730);
xor UO_624 (O_624,N_4679,N_4406);
nor UO_625 (O_625,N_4712,N_4511);
and UO_626 (O_626,N_4870,N_4758);
nand UO_627 (O_627,N_4248,N_4482);
or UO_628 (O_628,N_4653,N_4620);
or UO_629 (O_629,N_4500,N_4324);
or UO_630 (O_630,N_4703,N_4280);
or UO_631 (O_631,N_4119,N_4340);
nor UO_632 (O_632,N_4269,N_4184);
xor UO_633 (O_633,N_4430,N_4973);
nand UO_634 (O_634,N_4607,N_4473);
and UO_635 (O_635,N_4103,N_4181);
xor UO_636 (O_636,N_4026,N_4854);
nand UO_637 (O_637,N_4304,N_4525);
or UO_638 (O_638,N_4455,N_4918);
nand UO_639 (O_639,N_4423,N_4703);
xnor UO_640 (O_640,N_4992,N_4893);
nor UO_641 (O_641,N_4102,N_4571);
or UO_642 (O_642,N_4733,N_4761);
xor UO_643 (O_643,N_4695,N_4083);
xnor UO_644 (O_644,N_4305,N_4163);
nand UO_645 (O_645,N_4364,N_4954);
nor UO_646 (O_646,N_4793,N_4029);
nor UO_647 (O_647,N_4908,N_4272);
nand UO_648 (O_648,N_4605,N_4460);
and UO_649 (O_649,N_4200,N_4151);
and UO_650 (O_650,N_4313,N_4800);
or UO_651 (O_651,N_4894,N_4464);
nor UO_652 (O_652,N_4948,N_4126);
nor UO_653 (O_653,N_4150,N_4835);
nand UO_654 (O_654,N_4918,N_4392);
nand UO_655 (O_655,N_4783,N_4600);
and UO_656 (O_656,N_4961,N_4616);
and UO_657 (O_657,N_4405,N_4732);
and UO_658 (O_658,N_4643,N_4428);
xnor UO_659 (O_659,N_4043,N_4062);
and UO_660 (O_660,N_4007,N_4709);
and UO_661 (O_661,N_4364,N_4824);
nand UO_662 (O_662,N_4735,N_4503);
xnor UO_663 (O_663,N_4718,N_4003);
xor UO_664 (O_664,N_4645,N_4564);
xor UO_665 (O_665,N_4448,N_4886);
or UO_666 (O_666,N_4517,N_4378);
nor UO_667 (O_667,N_4410,N_4300);
and UO_668 (O_668,N_4850,N_4384);
nor UO_669 (O_669,N_4691,N_4790);
and UO_670 (O_670,N_4230,N_4254);
and UO_671 (O_671,N_4778,N_4623);
nor UO_672 (O_672,N_4320,N_4075);
nor UO_673 (O_673,N_4519,N_4853);
and UO_674 (O_674,N_4169,N_4337);
or UO_675 (O_675,N_4355,N_4294);
xor UO_676 (O_676,N_4467,N_4794);
and UO_677 (O_677,N_4260,N_4840);
xor UO_678 (O_678,N_4675,N_4348);
nand UO_679 (O_679,N_4454,N_4682);
xor UO_680 (O_680,N_4041,N_4270);
nand UO_681 (O_681,N_4682,N_4511);
or UO_682 (O_682,N_4317,N_4548);
or UO_683 (O_683,N_4426,N_4945);
nor UO_684 (O_684,N_4095,N_4960);
and UO_685 (O_685,N_4391,N_4313);
xor UO_686 (O_686,N_4445,N_4210);
or UO_687 (O_687,N_4876,N_4896);
or UO_688 (O_688,N_4418,N_4222);
nand UO_689 (O_689,N_4156,N_4988);
or UO_690 (O_690,N_4450,N_4119);
xor UO_691 (O_691,N_4330,N_4923);
xor UO_692 (O_692,N_4862,N_4711);
and UO_693 (O_693,N_4247,N_4332);
nand UO_694 (O_694,N_4267,N_4097);
nand UO_695 (O_695,N_4445,N_4257);
nor UO_696 (O_696,N_4888,N_4630);
or UO_697 (O_697,N_4603,N_4789);
nor UO_698 (O_698,N_4965,N_4905);
nor UO_699 (O_699,N_4987,N_4967);
xor UO_700 (O_700,N_4057,N_4616);
xnor UO_701 (O_701,N_4065,N_4359);
xor UO_702 (O_702,N_4880,N_4457);
nand UO_703 (O_703,N_4256,N_4316);
xnor UO_704 (O_704,N_4920,N_4062);
xnor UO_705 (O_705,N_4050,N_4630);
nand UO_706 (O_706,N_4848,N_4644);
nand UO_707 (O_707,N_4000,N_4911);
or UO_708 (O_708,N_4088,N_4161);
xor UO_709 (O_709,N_4625,N_4670);
and UO_710 (O_710,N_4878,N_4828);
nor UO_711 (O_711,N_4160,N_4743);
nand UO_712 (O_712,N_4192,N_4275);
nand UO_713 (O_713,N_4095,N_4999);
and UO_714 (O_714,N_4075,N_4588);
nand UO_715 (O_715,N_4763,N_4253);
xnor UO_716 (O_716,N_4746,N_4284);
xnor UO_717 (O_717,N_4485,N_4288);
or UO_718 (O_718,N_4166,N_4956);
and UO_719 (O_719,N_4975,N_4922);
nand UO_720 (O_720,N_4100,N_4489);
nand UO_721 (O_721,N_4391,N_4805);
nand UO_722 (O_722,N_4633,N_4400);
or UO_723 (O_723,N_4715,N_4097);
nor UO_724 (O_724,N_4389,N_4031);
nand UO_725 (O_725,N_4413,N_4135);
and UO_726 (O_726,N_4626,N_4071);
xnor UO_727 (O_727,N_4034,N_4747);
or UO_728 (O_728,N_4872,N_4740);
xnor UO_729 (O_729,N_4285,N_4311);
and UO_730 (O_730,N_4046,N_4300);
or UO_731 (O_731,N_4517,N_4002);
and UO_732 (O_732,N_4794,N_4992);
and UO_733 (O_733,N_4057,N_4691);
xnor UO_734 (O_734,N_4550,N_4175);
xnor UO_735 (O_735,N_4142,N_4998);
xnor UO_736 (O_736,N_4256,N_4009);
or UO_737 (O_737,N_4110,N_4389);
and UO_738 (O_738,N_4453,N_4393);
and UO_739 (O_739,N_4729,N_4243);
nor UO_740 (O_740,N_4692,N_4721);
nand UO_741 (O_741,N_4164,N_4254);
and UO_742 (O_742,N_4326,N_4174);
and UO_743 (O_743,N_4769,N_4565);
xor UO_744 (O_744,N_4225,N_4159);
xor UO_745 (O_745,N_4565,N_4767);
and UO_746 (O_746,N_4336,N_4419);
xnor UO_747 (O_747,N_4083,N_4964);
or UO_748 (O_748,N_4803,N_4344);
nor UO_749 (O_749,N_4103,N_4720);
or UO_750 (O_750,N_4796,N_4384);
and UO_751 (O_751,N_4648,N_4008);
xor UO_752 (O_752,N_4875,N_4277);
or UO_753 (O_753,N_4909,N_4021);
or UO_754 (O_754,N_4655,N_4851);
xnor UO_755 (O_755,N_4630,N_4200);
xnor UO_756 (O_756,N_4939,N_4955);
nand UO_757 (O_757,N_4482,N_4207);
nand UO_758 (O_758,N_4925,N_4920);
or UO_759 (O_759,N_4956,N_4553);
xor UO_760 (O_760,N_4748,N_4794);
or UO_761 (O_761,N_4277,N_4660);
xor UO_762 (O_762,N_4422,N_4678);
nand UO_763 (O_763,N_4219,N_4846);
nor UO_764 (O_764,N_4314,N_4841);
and UO_765 (O_765,N_4616,N_4638);
or UO_766 (O_766,N_4238,N_4524);
nand UO_767 (O_767,N_4923,N_4749);
xnor UO_768 (O_768,N_4955,N_4644);
and UO_769 (O_769,N_4548,N_4770);
nor UO_770 (O_770,N_4642,N_4573);
xor UO_771 (O_771,N_4364,N_4193);
xnor UO_772 (O_772,N_4538,N_4552);
or UO_773 (O_773,N_4612,N_4548);
nor UO_774 (O_774,N_4430,N_4723);
or UO_775 (O_775,N_4610,N_4939);
nor UO_776 (O_776,N_4333,N_4412);
nor UO_777 (O_777,N_4859,N_4758);
nand UO_778 (O_778,N_4618,N_4045);
nor UO_779 (O_779,N_4197,N_4872);
nand UO_780 (O_780,N_4824,N_4752);
or UO_781 (O_781,N_4201,N_4645);
nor UO_782 (O_782,N_4823,N_4256);
nor UO_783 (O_783,N_4232,N_4893);
and UO_784 (O_784,N_4155,N_4564);
nor UO_785 (O_785,N_4806,N_4550);
or UO_786 (O_786,N_4859,N_4943);
or UO_787 (O_787,N_4000,N_4633);
xor UO_788 (O_788,N_4263,N_4035);
nor UO_789 (O_789,N_4175,N_4328);
or UO_790 (O_790,N_4378,N_4880);
nand UO_791 (O_791,N_4964,N_4817);
nor UO_792 (O_792,N_4230,N_4420);
nand UO_793 (O_793,N_4237,N_4860);
xor UO_794 (O_794,N_4023,N_4853);
nand UO_795 (O_795,N_4926,N_4689);
nor UO_796 (O_796,N_4798,N_4135);
nand UO_797 (O_797,N_4250,N_4962);
or UO_798 (O_798,N_4737,N_4341);
nor UO_799 (O_799,N_4282,N_4789);
xnor UO_800 (O_800,N_4276,N_4859);
or UO_801 (O_801,N_4670,N_4049);
and UO_802 (O_802,N_4667,N_4061);
xor UO_803 (O_803,N_4725,N_4234);
xor UO_804 (O_804,N_4281,N_4486);
xnor UO_805 (O_805,N_4527,N_4993);
or UO_806 (O_806,N_4035,N_4627);
nor UO_807 (O_807,N_4736,N_4996);
nand UO_808 (O_808,N_4639,N_4419);
or UO_809 (O_809,N_4802,N_4020);
nand UO_810 (O_810,N_4319,N_4181);
and UO_811 (O_811,N_4235,N_4031);
and UO_812 (O_812,N_4720,N_4986);
or UO_813 (O_813,N_4035,N_4467);
nand UO_814 (O_814,N_4293,N_4912);
nor UO_815 (O_815,N_4124,N_4152);
or UO_816 (O_816,N_4583,N_4397);
nand UO_817 (O_817,N_4198,N_4522);
and UO_818 (O_818,N_4576,N_4083);
xnor UO_819 (O_819,N_4286,N_4933);
or UO_820 (O_820,N_4846,N_4156);
or UO_821 (O_821,N_4654,N_4345);
nor UO_822 (O_822,N_4156,N_4117);
or UO_823 (O_823,N_4601,N_4429);
nor UO_824 (O_824,N_4251,N_4757);
nand UO_825 (O_825,N_4956,N_4456);
nor UO_826 (O_826,N_4174,N_4666);
nor UO_827 (O_827,N_4831,N_4914);
nand UO_828 (O_828,N_4579,N_4606);
and UO_829 (O_829,N_4585,N_4412);
or UO_830 (O_830,N_4886,N_4855);
nand UO_831 (O_831,N_4341,N_4478);
and UO_832 (O_832,N_4860,N_4641);
nand UO_833 (O_833,N_4884,N_4611);
or UO_834 (O_834,N_4182,N_4853);
xor UO_835 (O_835,N_4342,N_4978);
xor UO_836 (O_836,N_4469,N_4812);
xor UO_837 (O_837,N_4968,N_4387);
and UO_838 (O_838,N_4544,N_4948);
nand UO_839 (O_839,N_4543,N_4301);
xnor UO_840 (O_840,N_4135,N_4699);
or UO_841 (O_841,N_4274,N_4323);
xnor UO_842 (O_842,N_4343,N_4245);
nor UO_843 (O_843,N_4969,N_4898);
nand UO_844 (O_844,N_4876,N_4518);
nor UO_845 (O_845,N_4361,N_4598);
xor UO_846 (O_846,N_4000,N_4684);
and UO_847 (O_847,N_4573,N_4662);
nand UO_848 (O_848,N_4237,N_4615);
nand UO_849 (O_849,N_4593,N_4395);
and UO_850 (O_850,N_4813,N_4588);
nor UO_851 (O_851,N_4897,N_4764);
and UO_852 (O_852,N_4348,N_4123);
nand UO_853 (O_853,N_4238,N_4170);
nor UO_854 (O_854,N_4716,N_4105);
or UO_855 (O_855,N_4785,N_4745);
and UO_856 (O_856,N_4032,N_4249);
xor UO_857 (O_857,N_4401,N_4232);
xor UO_858 (O_858,N_4306,N_4831);
nor UO_859 (O_859,N_4110,N_4359);
nand UO_860 (O_860,N_4467,N_4949);
and UO_861 (O_861,N_4867,N_4770);
and UO_862 (O_862,N_4032,N_4219);
nand UO_863 (O_863,N_4199,N_4066);
or UO_864 (O_864,N_4833,N_4718);
nor UO_865 (O_865,N_4261,N_4708);
and UO_866 (O_866,N_4933,N_4046);
nor UO_867 (O_867,N_4223,N_4204);
or UO_868 (O_868,N_4952,N_4658);
nor UO_869 (O_869,N_4041,N_4528);
xnor UO_870 (O_870,N_4253,N_4746);
or UO_871 (O_871,N_4385,N_4919);
nand UO_872 (O_872,N_4849,N_4651);
and UO_873 (O_873,N_4282,N_4028);
nand UO_874 (O_874,N_4754,N_4522);
and UO_875 (O_875,N_4160,N_4726);
xor UO_876 (O_876,N_4135,N_4076);
xnor UO_877 (O_877,N_4011,N_4322);
nor UO_878 (O_878,N_4381,N_4068);
or UO_879 (O_879,N_4450,N_4921);
xor UO_880 (O_880,N_4191,N_4086);
and UO_881 (O_881,N_4540,N_4776);
xnor UO_882 (O_882,N_4863,N_4812);
nor UO_883 (O_883,N_4875,N_4862);
or UO_884 (O_884,N_4431,N_4675);
or UO_885 (O_885,N_4412,N_4285);
nor UO_886 (O_886,N_4787,N_4260);
or UO_887 (O_887,N_4337,N_4215);
xor UO_888 (O_888,N_4421,N_4278);
nand UO_889 (O_889,N_4634,N_4784);
or UO_890 (O_890,N_4112,N_4071);
xor UO_891 (O_891,N_4139,N_4777);
nor UO_892 (O_892,N_4628,N_4159);
nand UO_893 (O_893,N_4042,N_4687);
nor UO_894 (O_894,N_4767,N_4612);
nor UO_895 (O_895,N_4911,N_4085);
and UO_896 (O_896,N_4803,N_4671);
nand UO_897 (O_897,N_4311,N_4626);
and UO_898 (O_898,N_4723,N_4448);
nor UO_899 (O_899,N_4364,N_4297);
xor UO_900 (O_900,N_4856,N_4108);
xnor UO_901 (O_901,N_4760,N_4921);
and UO_902 (O_902,N_4889,N_4708);
and UO_903 (O_903,N_4359,N_4554);
and UO_904 (O_904,N_4419,N_4486);
nand UO_905 (O_905,N_4975,N_4267);
or UO_906 (O_906,N_4285,N_4727);
xnor UO_907 (O_907,N_4806,N_4955);
or UO_908 (O_908,N_4944,N_4814);
or UO_909 (O_909,N_4205,N_4152);
nand UO_910 (O_910,N_4514,N_4812);
nand UO_911 (O_911,N_4323,N_4819);
nor UO_912 (O_912,N_4875,N_4416);
or UO_913 (O_913,N_4749,N_4437);
xor UO_914 (O_914,N_4069,N_4325);
or UO_915 (O_915,N_4925,N_4394);
xnor UO_916 (O_916,N_4871,N_4889);
xor UO_917 (O_917,N_4535,N_4267);
xnor UO_918 (O_918,N_4084,N_4907);
and UO_919 (O_919,N_4710,N_4396);
or UO_920 (O_920,N_4687,N_4680);
nor UO_921 (O_921,N_4870,N_4565);
and UO_922 (O_922,N_4671,N_4394);
or UO_923 (O_923,N_4965,N_4919);
nor UO_924 (O_924,N_4576,N_4971);
and UO_925 (O_925,N_4929,N_4933);
nor UO_926 (O_926,N_4131,N_4177);
and UO_927 (O_927,N_4910,N_4329);
or UO_928 (O_928,N_4098,N_4680);
nor UO_929 (O_929,N_4139,N_4611);
and UO_930 (O_930,N_4911,N_4722);
nand UO_931 (O_931,N_4890,N_4914);
nor UO_932 (O_932,N_4222,N_4132);
xor UO_933 (O_933,N_4199,N_4420);
xor UO_934 (O_934,N_4041,N_4943);
nor UO_935 (O_935,N_4882,N_4157);
and UO_936 (O_936,N_4208,N_4716);
xor UO_937 (O_937,N_4668,N_4127);
nor UO_938 (O_938,N_4576,N_4360);
and UO_939 (O_939,N_4835,N_4296);
nand UO_940 (O_940,N_4485,N_4003);
xnor UO_941 (O_941,N_4743,N_4241);
xnor UO_942 (O_942,N_4164,N_4946);
xor UO_943 (O_943,N_4907,N_4759);
xnor UO_944 (O_944,N_4147,N_4268);
and UO_945 (O_945,N_4495,N_4821);
nand UO_946 (O_946,N_4757,N_4697);
or UO_947 (O_947,N_4107,N_4360);
and UO_948 (O_948,N_4464,N_4493);
or UO_949 (O_949,N_4179,N_4748);
xor UO_950 (O_950,N_4791,N_4792);
or UO_951 (O_951,N_4763,N_4908);
xnor UO_952 (O_952,N_4274,N_4935);
nor UO_953 (O_953,N_4641,N_4850);
xor UO_954 (O_954,N_4061,N_4099);
nand UO_955 (O_955,N_4663,N_4065);
nor UO_956 (O_956,N_4221,N_4192);
or UO_957 (O_957,N_4225,N_4103);
nand UO_958 (O_958,N_4744,N_4926);
or UO_959 (O_959,N_4447,N_4844);
xnor UO_960 (O_960,N_4925,N_4924);
or UO_961 (O_961,N_4113,N_4091);
and UO_962 (O_962,N_4265,N_4853);
and UO_963 (O_963,N_4887,N_4062);
or UO_964 (O_964,N_4927,N_4170);
xnor UO_965 (O_965,N_4055,N_4781);
xor UO_966 (O_966,N_4095,N_4578);
or UO_967 (O_967,N_4661,N_4648);
nand UO_968 (O_968,N_4127,N_4005);
xnor UO_969 (O_969,N_4097,N_4024);
nor UO_970 (O_970,N_4285,N_4306);
nor UO_971 (O_971,N_4406,N_4192);
nor UO_972 (O_972,N_4539,N_4953);
nor UO_973 (O_973,N_4852,N_4674);
nand UO_974 (O_974,N_4519,N_4500);
xor UO_975 (O_975,N_4969,N_4675);
nand UO_976 (O_976,N_4982,N_4068);
nand UO_977 (O_977,N_4463,N_4378);
or UO_978 (O_978,N_4254,N_4717);
and UO_979 (O_979,N_4072,N_4488);
nor UO_980 (O_980,N_4135,N_4600);
nor UO_981 (O_981,N_4123,N_4171);
and UO_982 (O_982,N_4461,N_4225);
or UO_983 (O_983,N_4433,N_4178);
nand UO_984 (O_984,N_4327,N_4061);
nand UO_985 (O_985,N_4275,N_4585);
nor UO_986 (O_986,N_4357,N_4935);
xnor UO_987 (O_987,N_4044,N_4225);
or UO_988 (O_988,N_4471,N_4181);
nand UO_989 (O_989,N_4691,N_4299);
or UO_990 (O_990,N_4476,N_4562);
and UO_991 (O_991,N_4960,N_4535);
and UO_992 (O_992,N_4809,N_4357);
xor UO_993 (O_993,N_4950,N_4885);
xor UO_994 (O_994,N_4998,N_4792);
nor UO_995 (O_995,N_4407,N_4834);
nand UO_996 (O_996,N_4666,N_4177);
or UO_997 (O_997,N_4733,N_4593);
nand UO_998 (O_998,N_4036,N_4480);
nand UO_999 (O_999,N_4147,N_4434);
endmodule