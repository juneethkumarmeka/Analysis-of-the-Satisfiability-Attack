module basic_500_3000_500_15_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_211,In_109);
and U1 (N_1,In_120,In_427);
nand U2 (N_2,In_466,In_116);
and U3 (N_3,In_451,In_429);
nor U4 (N_4,In_374,In_391);
and U5 (N_5,In_212,In_275);
or U6 (N_6,In_157,In_117);
nor U7 (N_7,In_218,In_335);
xor U8 (N_8,In_119,In_165);
xor U9 (N_9,In_303,In_144);
nor U10 (N_10,In_497,In_70);
nor U11 (N_11,In_168,In_122);
nand U12 (N_12,In_395,In_27);
and U13 (N_13,In_184,In_356);
nand U14 (N_14,In_469,In_201);
nor U15 (N_15,In_464,In_5);
and U16 (N_16,In_200,In_219);
or U17 (N_17,In_204,In_25);
nand U18 (N_18,In_258,In_452);
and U19 (N_19,In_36,In_189);
or U20 (N_20,In_493,In_48);
nand U21 (N_21,In_312,In_454);
nand U22 (N_22,In_156,In_419);
xnor U23 (N_23,In_309,In_73);
and U24 (N_24,In_248,In_118);
nor U25 (N_25,In_345,In_185);
and U26 (N_26,In_237,In_351);
nor U27 (N_27,In_447,In_14);
nor U28 (N_28,In_271,In_132);
or U29 (N_29,In_193,In_438);
and U30 (N_30,In_197,In_114);
or U31 (N_31,In_364,In_333);
or U32 (N_32,In_477,In_272);
xnor U33 (N_33,In_79,In_456);
nand U34 (N_34,In_423,In_255);
nand U35 (N_35,In_16,In_32);
or U36 (N_36,In_56,In_3);
or U37 (N_37,In_485,In_76);
and U38 (N_38,In_100,In_394);
or U39 (N_39,In_318,In_232);
xnor U40 (N_40,In_11,In_435);
nand U41 (N_41,In_418,In_472);
and U42 (N_42,In_177,In_260);
and U43 (N_43,In_243,In_146);
nor U44 (N_44,In_236,In_289);
nand U45 (N_45,In_62,In_327);
and U46 (N_46,In_393,In_142);
or U47 (N_47,In_229,In_107);
or U48 (N_48,In_499,In_251);
nor U49 (N_49,In_360,In_199);
nor U50 (N_50,In_152,In_214);
and U51 (N_51,In_491,In_257);
nor U52 (N_52,In_145,In_96);
and U53 (N_53,In_421,In_473);
xor U54 (N_54,In_227,In_127);
nand U55 (N_55,In_131,In_247);
nand U56 (N_56,In_476,In_319);
or U57 (N_57,In_398,In_479);
and U58 (N_58,In_481,In_354);
or U59 (N_59,In_102,In_47);
nand U60 (N_60,In_325,In_431);
nand U61 (N_61,In_471,In_112);
or U62 (N_62,In_375,In_175);
or U63 (N_63,In_372,In_140);
nor U64 (N_64,In_183,In_254);
nor U65 (N_65,In_162,In_176);
nand U66 (N_66,In_361,In_344);
nand U67 (N_67,In_313,In_392);
and U68 (N_68,In_163,In_34);
or U69 (N_69,In_483,In_252);
nand U70 (N_70,In_170,In_337);
and U71 (N_71,In_383,In_77);
and U72 (N_72,In_40,In_274);
nand U73 (N_73,In_234,In_424);
nor U74 (N_74,In_305,In_71);
or U75 (N_75,In_437,In_215);
nand U76 (N_76,In_126,In_386);
or U77 (N_77,In_24,In_461);
or U78 (N_78,In_291,In_378);
nand U79 (N_79,In_26,In_6);
and U80 (N_80,In_94,In_192);
and U81 (N_81,In_217,In_203);
and U82 (N_82,In_329,In_417);
nor U83 (N_83,In_495,In_18);
nor U84 (N_84,In_206,In_230);
and U85 (N_85,In_113,In_180);
nor U86 (N_86,In_89,In_349);
and U87 (N_87,In_433,In_110);
nand U88 (N_88,In_8,In_85);
nor U89 (N_89,In_178,In_480);
nand U90 (N_90,In_450,In_53);
nand U91 (N_91,In_91,In_101);
nand U92 (N_92,In_388,In_64);
xnor U93 (N_93,In_128,In_324);
and U94 (N_94,In_151,In_428);
nor U95 (N_95,In_39,In_409);
nand U96 (N_96,In_288,In_256);
nand U97 (N_97,In_460,In_164);
or U98 (N_98,In_357,In_88);
nand U99 (N_99,In_339,In_346);
nand U100 (N_100,In_323,In_238);
or U101 (N_101,In_420,In_262);
and U102 (N_102,In_86,In_68);
or U103 (N_103,In_328,In_80);
nor U104 (N_104,In_441,In_396);
or U105 (N_105,In_434,In_382);
nand U106 (N_106,In_35,In_23);
or U107 (N_107,In_367,In_225);
and U108 (N_108,In_331,In_496);
or U109 (N_109,In_224,In_10);
nor U110 (N_110,In_366,In_83);
or U111 (N_111,In_261,In_415);
nand U112 (N_112,In_103,In_241);
nand U113 (N_113,In_336,In_202);
nor U114 (N_114,In_442,In_93);
nand U115 (N_115,In_81,In_332);
nand U116 (N_116,In_368,In_381);
and U117 (N_117,In_463,In_84);
or U118 (N_118,In_376,In_124);
nor U119 (N_119,In_209,In_194);
and U120 (N_120,In_279,In_121);
and U121 (N_121,In_266,In_486);
or U122 (N_122,In_426,In_154);
nor U123 (N_123,In_150,In_67);
and U124 (N_124,In_61,In_51);
nor U125 (N_125,In_208,In_195);
nand U126 (N_126,In_158,In_92);
or U127 (N_127,In_66,In_467);
or U128 (N_128,In_408,In_444);
nand U129 (N_129,In_414,In_311);
or U130 (N_130,In_359,In_348);
nand U131 (N_131,In_384,In_205);
or U132 (N_132,In_182,In_355);
and U133 (N_133,In_138,In_422);
nor U134 (N_134,In_173,In_167);
nand U135 (N_135,In_377,In_264);
and U136 (N_136,In_432,In_342);
or U137 (N_137,In_406,In_489);
and U138 (N_138,In_457,In_78);
nor U139 (N_139,In_317,In_465);
nor U140 (N_140,In_314,In_304);
and U141 (N_141,In_407,In_49);
or U142 (N_142,In_397,In_181);
and U143 (N_143,In_226,In_322);
nand U144 (N_144,In_478,In_196);
or U145 (N_145,In_136,In_296);
nor U146 (N_146,In_37,In_446);
nand U147 (N_147,In_403,In_231);
nand U148 (N_148,In_468,In_448);
nor U149 (N_149,In_307,In_290);
nor U150 (N_150,In_60,In_380);
nand U151 (N_151,In_123,In_240);
nor U152 (N_152,In_405,In_353);
and U153 (N_153,In_220,In_166);
nand U154 (N_154,In_293,In_43);
or U155 (N_155,In_347,In_74);
or U156 (N_156,In_172,In_470);
nand U157 (N_157,In_15,In_244);
nor U158 (N_158,In_487,In_270);
xor U159 (N_159,In_90,In_436);
nor U160 (N_160,In_213,In_20);
nand U161 (N_161,In_31,In_28);
nor U162 (N_162,In_416,In_410);
or U163 (N_163,In_280,In_259);
nor U164 (N_164,In_135,In_340);
nor U165 (N_165,In_263,In_155);
or U166 (N_166,In_320,In_462);
nor U167 (N_167,In_169,In_250);
nor U168 (N_168,In_57,In_153);
nand U169 (N_169,In_38,In_190);
or U170 (N_170,In_282,In_341);
nand U171 (N_171,In_330,In_298);
nor U172 (N_172,In_242,In_498);
nor U173 (N_173,In_458,In_46);
and U174 (N_174,In_19,In_453);
nor U175 (N_175,In_297,In_315);
nor U176 (N_176,In_334,In_283);
or U177 (N_177,In_97,In_186);
nor U178 (N_178,In_149,In_95);
nand U179 (N_179,In_294,In_111);
nand U180 (N_180,In_54,In_302);
and U181 (N_181,In_358,In_268);
nand U182 (N_182,In_228,In_161);
nand U183 (N_183,In_482,In_338);
nor U184 (N_184,In_370,In_308);
or U185 (N_185,In_75,In_267);
or U186 (N_186,In_44,In_239);
and U187 (N_187,In_321,In_385);
and U188 (N_188,In_17,In_171);
and U189 (N_189,In_425,In_9);
and U190 (N_190,In_411,In_379);
and U191 (N_191,In_390,In_160);
nand U192 (N_192,In_369,In_4);
and U193 (N_193,In_265,In_445);
nor U194 (N_194,In_475,In_187);
and U195 (N_195,In_105,In_129);
nor U196 (N_196,In_41,In_141);
and U197 (N_197,In_299,In_253);
nand U198 (N_198,In_281,In_389);
nand U199 (N_199,In_130,In_58);
nor U200 (N_200,N_148,N_89);
nand U201 (N_201,In_459,In_50);
nand U202 (N_202,N_121,N_112);
or U203 (N_203,In_310,N_24);
nor U204 (N_204,N_77,N_170);
nor U205 (N_205,N_196,N_192);
nor U206 (N_206,N_189,N_75);
nand U207 (N_207,N_177,In_488);
nor U208 (N_208,N_171,In_300);
nand U209 (N_209,In_222,N_47);
and U210 (N_210,In_474,N_98);
and U211 (N_211,N_185,N_99);
or U212 (N_212,N_168,N_97);
nor U213 (N_213,In_72,N_101);
or U214 (N_214,In_295,N_23);
nor U215 (N_215,N_90,N_1);
or U216 (N_216,In_33,N_64);
xnor U217 (N_217,In_278,N_15);
nor U218 (N_218,N_116,N_163);
nand U219 (N_219,N_186,N_107);
and U220 (N_220,In_401,N_73);
nor U221 (N_221,N_162,In_42);
nand U222 (N_222,In_1,N_9);
xnor U223 (N_223,N_48,N_174);
nand U224 (N_224,N_31,N_55);
and U225 (N_225,In_284,N_133);
or U226 (N_226,N_33,N_149);
and U227 (N_227,N_114,In_286);
nor U228 (N_228,N_43,In_12);
nor U229 (N_229,N_132,In_221);
nand U230 (N_230,N_105,In_22);
nor U231 (N_231,N_36,N_169);
nand U232 (N_232,N_20,N_70);
nor U233 (N_233,N_29,N_51);
and U234 (N_234,In_147,In_449);
nor U235 (N_235,N_46,In_371);
nand U236 (N_236,N_156,N_79);
nor U237 (N_237,In_148,In_65);
nand U238 (N_238,In_52,In_174);
and U239 (N_239,N_69,In_207);
and U240 (N_240,N_4,In_484);
and U241 (N_241,N_137,N_198);
and U242 (N_242,N_50,N_27);
and U243 (N_243,N_13,In_292);
and U244 (N_244,In_55,In_82);
nor U245 (N_245,In_404,N_142);
nor U246 (N_246,In_492,In_13);
xor U247 (N_247,N_124,N_80);
nand U248 (N_248,N_94,In_21);
or U249 (N_249,N_130,In_2);
or U250 (N_250,In_235,N_88);
and U251 (N_251,N_143,In_108);
and U252 (N_252,N_187,N_123);
nor U253 (N_253,N_176,In_115);
nor U254 (N_254,N_66,N_76);
nor U255 (N_255,N_135,N_115);
nand U256 (N_256,In_285,N_128);
nand U257 (N_257,N_117,N_11);
nor U258 (N_258,In_399,In_316);
and U259 (N_259,N_182,N_58);
nor U260 (N_260,In_455,N_59);
xor U261 (N_261,N_72,In_223);
and U262 (N_262,In_99,In_87);
and U263 (N_263,N_44,In_412);
nand U264 (N_264,N_188,N_52);
and U265 (N_265,In_365,In_69);
nand U266 (N_266,N_158,N_53);
or U267 (N_267,N_147,In_490);
nor U268 (N_268,In_387,In_350);
or U269 (N_269,N_157,N_197);
nand U270 (N_270,N_159,In_362);
nand U271 (N_271,N_106,N_141);
nor U272 (N_272,N_7,N_42);
nand U273 (N_273,N_195,In_63);
nand U274 (N_274,N_10,In_443);
or U275 (N_275,In_45,N_193);
and U276 (N_276,N_67,N_62);
or U277 (N_277,N_34,N_184);
or U278 (N_278,N_38,N_3);
nor U279 (N_279,N_45,In_137);
nor U280 (N_280,In_159,In_7);
nand U281 (N_281,In_277,In_249);
and U282 (N_282,N_199,In_233);
and U283 (N_283,N_96,In_273);
or U284 (N_284,N_68,N_71);
nand U285 (N_285,N_93,N_30);
or U286 (N_286,N_154,N_6);
nand U287 (N_287,N_63,N_25);
and U288 (N_288,N_183,In_139);
and U289 (N_289,N_19,N_153);
nor U290 (N_290,N_111,N_166);
nor U291 (N_291,N_16,N_160);
and U292 (N_292,In_269,N_18);
and U293 (N_293,N_95,In_106);
nand U294 (N_294,N_81,N_57);
or U295 (N_295,N_180,N_191);
or U296 (N_296,In_59,In_276);
and U297 (N_297,In_188,N_129);
nand U298 (N_298,N_28,N_92);
nor U299 (N_299,In_216,N_78);
nand U300 (N_300,N_145,N_179);
nand U301 (N_301,N_126,In_343);
and U302 (N_302,In_430,In_198);
or U303 (N_303,N_8,N_164);
nor U304 (N_304,N_120,N_131);
xor U305 (N_305,In_287,N_41);
or U306 (N_306,In_326,N_175);
or U307 (N_307,N_74,N_190);
nor U308 (N_308,N_161,N_17);
xor U309 (N_309,In_245,N_150);
and U310 (N_310,N_144,In_133);
xnor U311 (N_311,N_56,N_100);
and U312 (N_312,In_402,N_140);
nand U313 (N_313,N_110,N_60);
and U314 (N_314,N_54,N_151);
nor U315 (N_315,N_102,In_363);
nor U316 (N_316,In_400,In_352);
and U317 (N_317,N_12,N_173);
or U318 (N_318,N_125,In_301);
or U319 (N_319,N_134,In_134);
or U320 (N_320,N_155,In_439);
nand U321 (N_321,In_143,In_30);
or U322 (N_322,N_118,N_136);
or U323 (N_323,N_5,N_165);
nand U324 (N_324,In_125,N_152);
nand U325 (N_325,In_373,N_21);
nand U326 (N_326,N_108,N_39);
nand U327 (N_327,N_84,N_32);
and U328 (N_328,N_127,In_104);
nor U329 (N_329,In_494,In_440);
nand U330 (N_330,In_306,N_26);
and U331 (N_331,N_109,N_65);
nand U332 (N_332,N_194,In_191);
nand U333 (N_333,In_0,N_91);
and U334 (N_334,N_181,N_37);
nand U335 (N_335,N_172,N_104);
nor U336 (N_336,N_122,In_179);
nand U337 (N_337,N_85,N_83);
nand U338 (N_338,N_82,N_0);
nor U339 (N_339,In_413,N_2);
nand U340 (N_340,N_87,In_29);
nand U341 (N_341,N_40,N_35);
nand U342 (N_342,N_113,N_167);
nor U343 (N_343,N_119,In_210);
or U344 (N_344,N_139,N_86);
and U345 (N_345,N_103,N_138);
or U346 (N_346,N_178,In_246);
or U347 (N_347,N_61,In_98);
and U348 (N_348,N_14,N_49);
and U349 (N_349,N_22,N_146);
and U350 (N_350,N_2,N_93);
nor U351 (N_351,In_42,In_12);
nand U352 (N_352,N_9,N_63);
nand U353 (N_353,N_75,N_151);
nor U354 (N_354,In_7,In_287);
or U355 (N_355,N_13,N_115);
and U356 (N_356,N_136,In_125);
or U357 (N_357,In_82,In_284);
nand U358 (N_358,N_81,N_45);
or U359 (N_359,In_455,N_128);
or U360 (N_360,In_12,N_154);
and U361 (N_361,In_492,N_140);
and U362 (N_362,N_132,In_216);
nor U363 (N_363,In_125,In_439);
nor U364 (N_364,N_163,N_146);
and U365 (N_365,N_179,In_0);
nand U366 (N_366,N_154,N_50);
nand U367 (N_367,In_207,N_30);
and U368 (N_368,N_160,In_295);
nor U369 (N_369,N_1,In_69);
or U370 (N_370,In_30,In_108);
or U371 (N_371,In_287,N_162);
nand U372 (N_372,N_55,N_92);
or U373 (N_373,In_210,N_2);
and U374 (N_374,In_269,N_184);
nand U375 (N_375,N_138,N_139);
nor U376 (N_376,In_207,N_168);
nor U377 (N_377,N_9,In_443);
xnor U378 (N_378,In_365,N_59);
nand U379 (N_379,N_69,In_269);
xor U380 (N_380,N_144,N_117);
xnor U381 (N_381,N_77,N_135);
or U382 (N_382,In_45,In_306);
nor U383 (N_383,N_158,In_72);
xor U384 (N_384,N_92,N_111);
and U385 (N_385,In_30,N_123);
or U386 (N_386,In_413,N_3);
nand U387 (N_387,N_172,In_207);
and U388 (N_388,In_21,N_149);
and U389 (N_389,N_65,In_125);
or U390 (N_390,N_163,N_121);
and U391 (N_391,N_31,N_84);
nor U392 (N_392,N_190,N_112);
or U393 (N_393,N_102,In_439);
nand U394 (N_394,N_14,N_16);
and U395 (N_395,N_96,N_147);
and U396 (N_396,N_47,N_134);
or U397 (N_397,N_199,N_111);
nor U398 (N_398,In_286,In_474);
or U399 (N_399,N_90,In_413);
nand U400 (N_400,N_252,N_368);
and U401 (N_401,N_328,N_387);
nand U402 (N_402,N_343,N_347);
nand U403 (N_403,N_396,N_237);
xnor U404 (N_404,N_314,N_238);
nand U405 (N_405,N_259,N_287);
or U406 (N_406,N_253,N_215);
or U407 (N_407,N_234,N_205);
or U408 (N_408,N_263,N_383);
and U409 (N_409,N_214,N_364);
nand U410 (N_410,N_291,N_351);
nand U411 (N_411,N_294,N_369);
nand U412 (N_412,N_227,N_255);
nor U413 (N_413,N_338,N_266);
or U414 (N_414,N_318,N_262);
nor U415 (N_415,N_281,N_204);
or U416 (N_416,N_340,N_374);
nor U417 (N_417,N_394,N_304);
nor U418 (N_418,N_282,N_203);
and U419 (N_419,N_319,N_244);
nor U420 (N_420,N_366,N_295);
xor U421 (N_421,N_327,N_276);
nand U422 (N_422,N_359,N_218);
nor U423 (N_423,N_321,N_251);
nor U424 (N_424,N_283,N_337);
nand U425 (N_425,N_247,N_308);
nor U426 (N_426,N_322,N_326);
or U427 (N_427,N_375,N_230);
nor U428 (N_428,N_209,N_334);
and U429 (N_429,N_286,N_267);
or U430 (N_430,N_280,N_225);
or U431 (N_431,N_219,N_278);
and U432 (N_432,N_370,N_277);
or U433 (N_433,N_339,N_279);
nor U434 (N_434,N_305,N_246);
nand U435 (N_435,N_332,N_329);
xnor U436 (N_436,N_210,N_330);
nand U437 (N_437,N_222,N_272);
and U438 (N_438,N_381,N_254);
nand U439 (N_439,N_354,N_208);
and U440 (N_440,N_315,N_206);
or U441 (N_441,N_233,N_216);
or U442 (N_442,N_213,N_229);
xnor U443 (N_443,N_290,N_323);
nand U444 (N_444,N_273,N_243);
and U445 (N_445,N_235,N_299);
and U446 (N_446,N_382,N_249);
or U447 (N_447,N_211,N_324);
xor U448 (N_448,N_200,N_392);
nand U449 (N_449,N_344,N_207);
nand U450 (N_450,N_371,N_312);
and U451 (N_451,N_333,N_316);
nand U452 (N_452,N_223,N_264);
or U453 (N_453,N_306,N_212);
and U454 (N_454,N_367,N_248);
nor U455 (N_455,N_399,N_377);
or U456 (N_456,N_220,N_217);
nor U457 (N_457,N_355,N_391);
and U458 (N_458,N_384,N_257);
or U459 (N_459,N_297,N_202);
or U460 (N_460,N_336,N_240);
nand U461 (N_461,N_242,N_388);
nand U462 (N_462,N_228,N_357);
nand U463 (N_463,N_268,N_310);
nand U464 (N_464,N_361,N_231);
nor U465 (N_465,N_362,N_307);
or U466 (N_466,N_298,N_258);
and U467 (N_467,N_358,N_260);
nor U468 (N_468,N_397,N_345);
or U469 (N_469,N_224,N_353);
nor U470 (N_470,N_320,N_389);
and U471 (N_471,N_341,N_303);
nand U472 (N_472,N_313,N_311);
and U473 (N_473,N_379,N_386);
nand U474 (N_474,N_265,N_372);
or U475 (N_475,N_346,N_342);
nor U476 (N_476,N_331,N_245);
nor U477 (N_477,N_356,N_348);
or U478 (N_478,N_296,N_241);
nor U479 (N_479,N_292,N_275);
nand U480 (N_480,N_271,N_378);
nor U481 (N_481,N_335,N_393);
or U482 (N_482,N_395,N_239);
or U483 (N_483,N_226,N_274);
and U484 (N_484,N_285,N_236);
nor U485 (N_485,N_363,N_288);
and U486 (N_486,N_380,N_385);
nand U487 (N_487,N_390,N_232);
and U488 (N_488,N_250,N_270);
nand U489 (N_489,N_365,N_352);
and U490 (N_490,N_309,N_256);
nor U491 (N_491,N_398,N_293);
nor U492 (N_492,N_201,N_376);
nor U493 (N_493,N_289,N_350);
nor U494 (N_494,N_261,N_317);
or U495 (N_495,N_360,N_300);
and U496 (N_496,N_221,N_269);
or U497 (N_497,N_325,N_301);
nor U498 (N_498,N_349,N_302);
nor U499 (N_499,N_373,N_284);
nor U500 (N_500,N_340,N_283);
or U501 (N_501,N_371,N_266);
and U502 (N_502,N_262,N_309);
nor U503 (N_503,N_301,N_225);
and U504 (N_504,N_353,N_291);
nand U505 (N_505,N_314,N_233);
nand U506 (N_506,N_318,N_314);
and U507 (N_507,N_272,N_292);
nand U508 (N_508,N_314,N_356);
nand U509 (N_509,N_304,N_353);
and U510 (N_510,N_215,N_213);
and U511 (N_511,N_368,N_211);
nand U512 (N_512,N_379,N_234);
nor U513 (N_513,N_212,N_220);
nand U514 (N_514,N_226,N_276);
nor U515 (N_515,N_357,N_229);
and U516 (N_516,N_326,N_330);
nor U517 (N_517,N_375,N_251);
and U518 (N_518,N_250,N_206);
nand U519 (N_519,N_235,N_353);
and U520 (N_520,N_293,N_253);
and U521 (N_521,N_343,N_265);
and U522 (N_522,N_340,N_302);
or U523 (N_523,N_242,N_248);
nand U524 (N_524,N_277,N_259);
nor U525 (N_525,N_345,N_214);
or U526 (N_526,N_384,N_348);
nand U527 (N_527,N_310,N_261);
or U528 (N_528,N_241,N_262);
and U529 (N_529,N_351,N_392);
or U530 (N_530,N_360,N_229);
and U531 (N_531,N_291,N_213);
nor U532 (N_532,N_313,N_364);
and U533 (N_533,N_212,N_371);
nor U534 (N_534,N_376,N_222);
or U535 (N_535,N_232,N_329);
nand U536 (N_536,N_268,N_380);
and U537 (N_537,N_218,N_391);
xor U538 (N_538,N_223,N_205);
or U539 (N_539,N_329,N_284);
nand U540 (N_540,N_298,N_324);
nor U541 (N_541,N_388,N_325);
and U542 (N_542,N_262,N_250);
nand U543 (N_543,N_258,N_311);
nand U544 (N_544,N_329,N_369);
and U545 (N_545,N_216,N_320);
and U546 (N_546,N_216,N_249);
or U547 (N_547,N_305,N_201);
and U548 (N_548,N_347,N_295);
nand U549 (N_549,N_375,N_372);
and U550 (N_550,N_223,N_309);
nand U551 (N_551,N_316,N_205);
and U552 (N_552,N_362,N_378);
and U553 (N_553,N_366,N_249);
and U554 (N_554,N_351,N_397);
nand U555 (N_555,N_285,N_306);
nor U556 (N_556,N_328,N_311);
nor U557 (N_557,N_286,N_388);
xnor U558 (N_558,N_284,N_209);
nor U559 (N_559,N_321,N_271);
nand U560 (N_560,N_235,N_348);
nor U561 (N_561,N_343,N_312);
or U562 (N_562,N_326,N_245);
nand U563 (N_563,N_349,N_281);
or U564 (N_564,N_302,N_325);
nor U565 (N_565,N_256,N_327);
nand U566 (N_566,N_297,N_261);
or U567 (N_567,N_344,N_244);
and U568 (N_568,N_302,N_390);
nand U569 (N_569,N_203,N_290);
nand U570 (N_570,N_230,N_364);
and U571 (N_571,N_394,N_302);
and U572 (N_572,N_358,N_203);
and U573 (N_573,N_207,N_375);
or U574 (N_574,N_389,N_306);
nand U575 (N_575,N_273,N_361);
nor U576 (N_576,N_225,N_320);
nor U577 (N_577,N_267,N_394);
or U578 (N_578,N_355,N_324);
or U579 (N_579,N_251,N_237);
nand U580 (N_580,N_266,N_251);
nand U581 (N_581,N_333,N_202);
nand U582 (N_582,N_324,N_361);
and U583 (N_583,N_393,N_253);
nand U584 (N_584,N_270,N_321);
or U585 (N_585,N_201,N_304);
nor U586 (N_586,N_389,N_312);
nand U587 (N_587,N_365,N_343);
nand U588 (N_588,N_238,N_384);
or U589 (N_589,N_205,N_312);
nand U590 (N_590,N_279,N_389);
nand U591 (N_591,N_212,N_308);
nor U592 (N_592,N_269,N_248);
or U593 (N_593,N_209,N_299);
or U594 (N_594,N_396,N_296);
or U595 (N_595,N_311,N_361);
and U596 (N_596,N_285,N_234);
or U597 (N_597,N_220,N_325);
or U598 (N_598,N_244,N_364);
and U599 (N_599,N_353,N_281);
nor U600 (N_600,N_547,N_437);
nand U601 (N_601,N_535,N_405);
and U602 (N_602,N_512,N_411);
nor U603 (N_603,N_451,N_426);
nand U604 (N_604,N_574,N_508);
and U605 (N_605,N_497,N_414);
nor U606 (N_606,N_469,N_517);
nor U607 (N_607,N_514,N_511);
nor U608 (N_608,N_513,N_433);
and U609 (N_609,N_457,N_431);
or U610 (N_610,N_586,N_596);
nor U611 (N_611,N_595,N_505);
nand U612 (N_612,N_550,N_554);
or U613 (N_613,N_453,N_500);
and U614 (N_614,N_441,N_518);
or U615 (N_615,N_459,N_576);
and U616 (N_616,N_585,N_502);
nor U617 (N_617,N_587,N_532);
nand U618 (N_618,N_556,N_592);
and U619 (N_619,N_403,N_476);
and U620 (N_620,N_570,N_466);
and U621 (N_621,N_536,N_493);
or U622 (N_622,N_425,N_479);
nor U623 (N_623,N_424,N_427);
and U624 (N_624,N_446,N_471);
nor U625 (N_625,N_452,N_551);
nand U626 (N_626,N_454,N_438);
nand U627 (N_627,N_489,N_488);
nor U628 (N_628,N_523,N_448);
or U629 (N_629,N_491,N_584);
nor U630 (N_630,N_402,N_423);
and U631 (N_631,N_559,N_460);
or U632 (N_632,N_510,N_546);
and U633 (N_633,N_516,N_591);
and U634 (N_634,N_429,N_468);
nand U635 (N_635,N_499,N_565);
and U636 (N_636,N_544,N_524);
nand U637 (N_637,N_447,N_569);
nand U638 (N_638,N_567,N_412);
and U639 (N_639,N_478,N_597);
nor U640 (N_640,N_539,N_475);
or U641 (N_641,N_571,N_545);
and U642 (N_642,N_407,N_417);
nand U643 (N_643,N_549,N_404);
and U644 (N_644,N_590,N_495);
or U645 (N_645,N_498,N_579);
nor U646 (N_646,N_435,N_480);
or U647 (N_647,N_542,N_430);
and U648 (N_648,N_477,N_530);
or U649 (N_649,N_563,N_436);
nor U650 (N_650,N_538,N_409);
nor U651 (N_651,N_558,N_577);
nand U652 (N_652,N_520,N_525);
nand U653 (N_653,N_548,N_521);
nor U654 (N_654,N_434,N_494);
xnor U655 (N_655,N_526,N_474);
or U656 (N_656,N_566,N_519);
or U657 (N_657,N_557,N_504);
or U658 (N_658,N_575,N_555);
nand U659 (N_659,N_462,N_482);
or U660 (N_660,N_537,N_439);
and U661 (N_661,N_473,N_506);
xor U662 (N_662,N_487,N_588);
nand U663 (N_663,N_580,N_583);
nand U664 (N_664,N_470,N_507);
or U665 (N_665,N_598,N_484);
or U666 (N_666,N_496,N_422);
or U667 (N_667,N_455,N_444);
and U668 (N_668,N_568,N_467);
nor U669 (N_669,N_456,N_533);
and U670 (N_670,N_593,N_415);
and U671 (N_671,N_492,N_582);
and U672 (N_672,N_522,N_419);
or U673 (N_673,N_408,N_501);
and U674 (N_674,N_406,N_534);
nand U675 (N_675,N_450,N_540);
or U676 (N_676,N_527,N_458);
or U677 (N_677,N_413,N_573);
or U678 (N_678,N_486,N_561);
nor U679 (N_679,N_440,N_552);
nor U680 (N_680,N_421,N_564);
nand U681 (N_681,N_464,N_420);
and U682 (N_682,N_449,N_594);
nor U683 (N_683,N_543,N_509);
nor U684 (N_684,N_463,N_445);
nand U685 (N_685,N_416,N_581);
nor U686 (N_686,N_428,N_442);
and U687 (N_687,N_578,N_465);
nand U688 (N_688,N_503,N_432);
or U689 (N_689,N_490,N_481);
nor U690 (N_690,N_483,N_562);
and U691 (N_691,N_529,N_485);
or U692 (N_692,N_401,N_553);
nand U693 (N_693,N_589,N_541);
nor U694 (N_694,N_400,N_560);
or U695 (N_695,N_472,N_531);
nor U696 (N_696,N_418,N_528);
nand U697 (N_697,N_515,N_410);
or U698 (N_698,N_599,N_572);
and U699 (N_699,N_461,N_443);
or U700 (N_700,N_487,N_584);
nand U701 (N_701,N_452,N_585);
and U702 (N_702,N_587,N_537);
nand U703 (N_703,N_565,N_503);
nor U704 (N_704,N_550,N_596);
nor U705 (N_705,N_414,N_435);
or U706 (N_706,N_599,N_505);
nand U707 (N_707,N_507,N_444);
or U708 (N_708,N_576,N_580);
nor U709 (N_709,N_534,N_487);
nor U710 (N_710,N_477,N_502);
nor U711 (N_711,N_426,N_512);
and U712 (N_712,N_534,N_423);
and U713 (N_713,N_473,N_519);
xor U714 (N_714,N_519,N_488);
and U715 (N_715,N_402,N_486);
and U716 (N_716,N_445,N_441);
nor U717 (N_717,N_486,N_415);
nor U718 (N_718,N_475,N_582);
and U719 (N_719,N_575,N_484);
nor U720 (N_720,N_568,N_430);
and U721 (N_721,N_482,N_552);
nor U722 (N_722,N_437,N_436);
or U723 (N_723,N_547,N_411);
nor U724 (N_724,N_529,N_502);
nand U725 (N_725,N_483,N_424);
nor U726 (N_726,N_571,N_483);
and U727 (N_727,N_553,N_447);
nand U728 (N_728,N_589,N_493);
nor U729 (N_729,N_598,N_404);
nand U730 (N_730,N_528,N_588);
nand U731 (N_731,N_448,N_430);
and U732 (N_732,N_516,N_583);
nor U733 (N_733,N_424,N_563);
nand U734 (N_734,N_579,N_523);
and U735 (N_735,N_449,N_412);
nor U736 (N_736,N_582,N_500);
nor U737 (N_737,N_447,N_409);
nor U738 (N_738,N_445,N_548);
and U739 (N_739,N_441,N_438);
nor U740 (N_740,N_554,N_521);
nand U741 (N_741,N_528,N_466);
nand U742 (N_742,N_548,N_476);
nand U743 (N_743,N_598,N_536);
or U744 (N_744,N_545,N_499);
nand U745 (N_745,N_584,N_453);
nor U746 (N_746,N_411,N_535);
nand U747 (N_747,N_537,N_524);
nor U748 (N_748,N_475,N_432);
and U749 (N_749,N_403,N_522);
and U750 (N_750,N_407,N_576);
xor U751 (N_751,N_479,N_494);
nor U752 (N_752,N_431,N_521);
or U753 (N_753,N_412,N_561);
nand U754 (N_754,N_418,N_467);
or U755 (N_755,N_425,N_546);
or U756 (N_756,N_425,N_404);
nand U757 (N_757,N_582,N_510);
nor U758 (N_758,N_495,N_444);
nor U759 (N_759,N_456,N_571);
or U760 (N_760,N_486,N_585);
nand U761 (N_761,N_567,N_499);
nor U762 (N_762,N_436,N_415);
and U763 (N_763,N_538,N_513);
nor U764 (N_764,N_405,N_469);
nand U765 (N_765,N_562,N_598);
and U766 (N_766,N_543,N_488);
or U767 (N_767,N_419,N_430);
nand U768 (N_768,N_510,N_524);
nand U769 (N_769,N_548,N_455);
and U770 (N_770,N_566,N_425);
nor U771 (N_771,N_522,N_525);
or U772 (N_772,N_446,N_542);
nor U773 (N_773,N_544,N_518);
nand U774 (N_774,N_411,N_452);
nor U775 (N_775,N_430,N_482);
nand U776 (N_776,N_511,N_590);
nor U777 (N_777,N_557,N_577);
and U778 (N_778,N_510,N_444);
and U779 (N_779,N_533,N_429);
or U780 (N_780,N_564,N_460);
nand U781 (N_781,N_499,N_480);
nand U782 (N_782,N_434,N_534);
and U783 (N_783,N_500,N_412);
and U784 (N_784,N_590,N_427);
and U785 (N_785,N_533,N_535);
and U786 (N_786,N_508,N_406);
nor U787 (N_787,N_556,N_454);
nor U788 (N_788,N_450,N_471);
xnor U789 (N_789,N_477,N_433);
and U790 (N_790,N_554,N_534);
nand U791 (N_791,N_543,N_599);
nor U792 (N_792,N_466,N_578);
nor U793 (N_793,N_536,N_505);
or U794 (N_794,N_570,N_414);
nand U795 (N_795,N_584,N_519);
nor U796 (N_796,N_581,N_418);
xor U797 (N_797,N_590,N_465);
nor U798 (N_798,N_559,N_576);
or U799 (N_799,N_554,N_499);
nor U800 (N_800,N_667,N_752);
nand U801 (N_801,N_726,N_749);
or U802 (N_802,N_717,N_678);
nor U803 (N_803,N_642,N_727);
or U804 (N_804,N_694,N_619);
or U805 (N_805,N_637,N_771);
nand U806 (N_806,N_705,N_611);
or U807 (N_807,N_769,N_788);
nand U808 (N_808,N_766,N_765);
or U809 (N_809,N_670,N_745);
nand U810 (N_810,N_790,N_700);
nand U811 (N_811,N_608,N_675);
and U812 (N_812,N_721,N_639);
or U813 (N_813,N_793,N_662);
or U814 (N_814,N_695,N_647);
and U815 (N_815,N_653,N_648);
or U816 (N_816,N_724,N_699);
and U817 (N_817,N_644,N_686);
xor U818 (N_818,N_677,N_605);
and U819 (N_819,N_621,N_767);
and U820 (N_820,N_685,N_778);
and U821 (N_821,N_691,N_618);
nand U822 (N_822,N_748,N_761);
nor U823 (N_823,N_645,N_676);
nand U824 (N_824,N_751,N_663);
nand U825 (N_825,N_607,N_733);
nand U826 (N_826,N_616,N_776);
or U827 (N_827,N_603,N_711);
or U828 (N_828,N_697,N_696);
nor U829 (N_829,N_782,N_630);
or U830 (N_830,N_713,N_635);
or U831 (N_831,N_680,N_651);
nand U832 (N_832,N_660,N_720);
nand U833 (N_833,N_683,N_757);
nor U834 (N_834,N_643,N_764);
nand U835 (N_835,N_785,N_780);
nor U836 (N_836,N_789,N_715);
nor U837 (N_837,N_728,N_617);
or U838 (N_838,N_734,N_736);
and U839 (N_839,N_796,N_656);
or U840 (N_840,N_710,N_661);
or U841 (N_841,N_792,N_755);
and U842 (N_842,N_763,N_681);
nor U843 (N_843,N_669,N_640);
nor U844 (N_844,N_768,N_772);
nor U845 (N_845,N_673,N_627);
and U846 (N_846,N_799,N_629);
and U847 (N_847,N_604,N_707);
or U848 (N_848,N_610,N_716);
and U849 (N_849,N_774,N_787);
nand U850 (N_850,N_701,N_730);
nor U851 (N_851,N_714,N_623);
xnor U852 (N_852,N_665,N_703);
nor U853 (N_853,N_758,N_798);
nand U854 (N_854,N_746,N_668);
nand U855 (N_855,N_739,N_698);
and U856 (N_856,N_738,N_797);
and U857 (N_857,N_614,N_631);
nor U858 (N_858,N_600,N_641);
nor U859 (N_859,N_652,N_636);
nand U860 (N_860,N_620,N_754);
nor U861 (N_861,N_679,N_612);
nor U862 (N_862,N_659,N_646);
nor U863 (N_863,N_781,N_775);
and U864 (N_864,N_747,N_756);
and U865 (N_865,N_773,N_784);
or U866 (N_866,N_795,N_672);
nor U867 (N_867,N_649,N_657);
nor U868 (N_868,N_750,N_622);
or U869 (N_869,N_712,N_682);
or U870 (N_870,N_737,N_744);
and U871 (N_871,N_729,N_634);
or U872 (N_872,N_615,N_741);
nor U873 (N_873,N_740,N_777);
nor U874 (N_874,N_654,N_719);
and U875 (N_875,N_783,N_602);
nand U876 (N_876,N_786,N_625);
or U877 (N_877,N_638,N_628);
and U878 (N_878,N_671,N_674);
and U879 (N_879,N_762,N_601);
or U880 (N_880,N_731,N_609);
nand U881 (N_881,N_658,N_693);
nor U882 (N_882,N_702,N_735);
and U883 (N_883,N_794,N_770);
nand U884 (N_884,N_624,N_655);
and U885 (N_885,N_791,N_753);
nand U886 (N_886,N_759,N_742);
or U887 (N_887,N_760,N_633);
nor U888 (N_888,N_650,N_706);
and U889 (N_889,N_689,N_723);
nand U890 (N_890,N_709,N_664);
nand U891 (N_891,N_606,N_704);
or U892 (N_892,N_687,N_732);
nor U893 (N_893,N_626,N_690);
nand U894 (N_894,N_708,N_688);
nand U895 (N_895,N_692,N_613);
or U896 (N_896,N_666,N_722);
and U897 (N_897,N_684,N_779);
nor U898 (N_898,N_718,N_725);
nand U899 (N_899,N_743,N_632);
nand U900 (N_900,N_764,N_748);
nand U901 (N_901,N_638,N_766);
and U902 (N_902,N_767,N_704);
and U903 (N_903,N_769,N_665);
and U904 (N_904,N_732,N_741);
and U905 (N_905,N_653,N_691);
nor U906 (N_906,N_661,N_794);
xnor U907 (N_907,N_683,N_639);
and U908 (N_908,N_713,N_744);
nor U909 (N_909,N_781,N_790);
nand U910 (N_910,N_798,N_794);
nand U911 (N_911,N_794,N_744);
or U912 (N_912,N_636,N_788);
nand U913 (N_913,N_764,N_772);
and U914 (N_914,N_660,N_728);
or U915 (N_915,N_761,N_631);
or U916 (N_916,N_784,N_780);
or U917 (N_917,N_658,N_751);
and U918 (N_918,N_709,N_711);
and U919 (N_919,N_736,N_626);
xnor U920 (N_920,N_759,N_690);
nor U921 (N_921,N_613,N_677);
nor U922 (N_922,N_798,N_762);
nor U923 (N_923,N_644,N_652);
nor U924 (N_924,N_629,N_725);
nor U925 (N_925,N_687,N_792);
nand U926 (N_926,N_653,N_769);
or U927 (N_927,N_654,N_789);
or U928 (N_928,N_635,N_614);
and U929 (N_929,N_720,N_706);
nand U930 (N_930,N_653,N_645);
or U931 (N_931,N_685,N_650);
or U932 (N_932,N_725,N_639);
or U933 (N_933,N_635,N_624);
or U934 (N_934,N_603,N_665);
or U935 (N_935,N_749,N_785);
nor U936 (N_936,N_690,N_610);
nor U937 (N_937,N_774,N_650);
and U938 (N_938,N_654,N_713);
nor U939 (N_939,N_677,N_629);
and U940 (N_940,N_771,N_777);
or U941 (N_941,N_637,N_601);
or U942 (N_942,N_776,N_656);
nand U943 (N_943,N_755,N_796);
and U944 (N_944,N_781,N_642);
or U945 (N_945,N_732,N_704);
nor U946 (N_946,N_634,N_665);
nand U947 (N_947,N_785,N_720);
or U948 (N_948,N_688,N_619);
nand U949 (N_949,N_757,N_628);
and U950 (N_950,N_785,N_683);
and U951 (N_951,N_797,N_693);
nor U952 (N_952,N_743,N_790);
nand U953 (N_953,N_658,N_634);
and U954 (N_954,N_608,N_612);
and U955 (N_955,N_659,N_691);
nor U956 (N_956,N_676,N_781);
nor U957 (N_957,N_655,N_770);
nor U958 (N_958,N_672,N_702);
nand U959 (N_959,N_703,N_693);
nand U960 (N_960,N_622,N_663);
nor U961 (N_961,N_603,N_730);
or U962 (N_962,N_704,N_682);
and U963 (N_963,N_617,N_705);
or U964 (N_964,N_739,N_781);
nor U965 (N_965,N_786,N_601);
nor U966 (N_966,N_761,N_714);
nand U967 (N_967,N_642,N_719);
and U968 (N_968,N_715,N_610);
or U969 (N_969,N_671,N_609);
nand U970 (N_970,N_667,N_652);
nand U971 (N_971,N_774,N_707);
or U972 (N_972,N_707,N_740);
nor U973 (N_973,N_744,N_700);
or U974 (N_974,N_655,N_788);
and U975 (N_975,N_759,N_760);
nand U976 (N_976,N_664,N_748);
and U977 (N_977,N_728,N_627);
nor U978 (N_978,N_697,N_648);
and U979 (N_979,N_705,N_740);
nor U980 (N_980,N_730,N_720);
nand U981 (N_981,N_776,N_754);
nor U982 (N_982,N_715,N_636);
or U983 (N_983,N_604,N_754);
nand U984 (N_984,N_773,N_647);
and U985 (N_985,N_601,N_763);
or U986 (N_986,N_643,N_736);
or U987 (N_987,N_673,N_711);
or U988 (N_988,N_769,N_640);
nand U989 (N_989,N_645,N_659);
nand U990 (N_990,N_774,N_662);
and U991 (N_991,N_662,N_799);
or U992 (N_992,N_787,N_642);
or U993 (N_993,N_695,N_612);
or U994 (N_994,N_639,N_710);
or U995 (N_995,N_716,N_619);
nand U996 (N_996,N_603,N_695);
nand U997 (N_997,N_642,N_744);
nand U998 (N_998,N_627,N_619);
nand U999 (N_999,N_754,N_648);
nand U1000 (N_1000,N_992,N_931);
nor U1001 (N_1001,N_848,N_991);
or U1002 (N_1002,N_954,N_858);
or U1003 (N_1003,N_953,N_946);
xor U1004 (N_1004,N_868,N_889);
or U1005 (N_1005,N_828,N_920);
or U1006 (N_1006,N_820,N_812);
or U1007 (N_1007,N_813,N_964);
and U1008 (N_1008,N_918,N_869);
and U1009 (N_1009,N_923,N_938);
nor U1010 (N_1010,N_926,N_961);
nand U1011 (N_1011,N_883,N_891);
nand U1012 (N_1012,N_811,N_925);
and U1013 (N_1013,N_943,N_841);
nor U1014 (N_1014,N_885,N_928);
nor U1015 (N_1015,N_949,N_838);
nand U1016 (N_1016,N_871,N_998);
nand U1017 (N_1017,N_963,N_945);
and U1018 (N_1018,N_944,N_922);
nand U1019 (N_1019,N_906,N_888);
or U1020 (N_1020,N_849,N_932);
nand U1021 (N_1021,N_912,N_836);
nor U1022 (N_1022,N_965,N_853);
and U1023 (N_1023,N_977,N_984);
and U1024 (N_1024,N_893,N_892);
and U1025 (N_1025,N_894,N_911);
nor U1026 (N_1026,N_987,N_983);
or U1027 (N_1027,N_956,N_887);
xnor U1028 (N_1028,N_942,N_916);
nand U1029 (N_1029,N_840,N_978);
and U1030 (N_1030,N_855,N_835);
nor U1031 (N_1031,N_872,N_933);
xor U1032 (N_1032,N_900,N_952);
nor U1033 (N_1033,N_880,N_846);
and U1034 (N_1034,N_966,N_814);
nand U1035 (N_1035,N_962,N_817);
nand U1036 (N_1036,N_851,N_809);
nand U1037 (N_1037,N_986,N_873);
nand U1038 (N_1038,N_903,N_951);
and U1039 (N_1039,N_860,N_822);
nor U1040 (N_1040,N_821,N_971);
nor U1041 (N_1041,N_985,N_877);
nor U1042 (N_1042,N_833,N_973);
xor U1043 (N_1043,N_898,N_806);
and U1044 (N_1044,N_831,N_957);
nand U1045 (N_1045,N_913,N_930);
or U1046 (N_1046,N_874,N_847);
nor U1047 (N_1047,N_968,N_994);
and U1048 (N_1048,N_999,N_852);
or U1049 (N_1049,N_832,N_910);
nand U1050 (N_1050,N_967,N_854);
or U1051 (N_1051,N_830,N_870);
nand U1052 (N_1052,N_807,N_936);
nand U1053 (N_1053,N_878,N_879);
or U1054 (N_1054,N_884,N_881);
and U1055 (N_1055,N_917,N_907);
nor U1056 (N_1056,N_914,N_929);
nand U1057 (N_1057,N_864,N_842);
nand U1058 (N_1058,N_866,N_934);
or U1059 (N_1059,N_975,N_808);
nor U1060 (N_1060,N_805,N_800);
nor U1061 (N_1061,N_935,N_950);
nand U1062 (N_1062,N_988,N_958);
and U1063 (N_1063,N_982,N_976);
nand U1064 (N_1064,N_837,N_823);
or U1065 (N_1065,N_895,N_801);
nor U1066 (N_1066,N_827,N_989);
or U1067 (N_1067,N_886,N_927);
nor U1068 (N_1068,N_981,N_850);
nor U1069 (N_1069,N_921,N_824);
or U1070 (N_1070,N_859,N_919);
and U1071 (N_1071,N_845,N_844);
and U1072 (N_1072,N_959,N_905);
or U1073 (N_1073,N_897,N_834);
and U1074 (N_1074,N_810,N_899);
nor U1075 (N_1075,N_825,N_826);
or U1076 (N_1076,N_862,N_819);
nor U1077 (N_1077,N_909,N_867);
or U1078 (N_1078,N_815,N_856);
nor U1079 (N_1079,N_901,N_882);
and U1080 (N_1080,N_876,N_863);
or U1081 (N_1081,N_839,N_947);
nor U1082 (N_1082,N_995,N_960);
or U1083 (N_1083,N_843,N_969);
and U1084 (N_1084,N_818,N_857);
nand U1085 (N_1085,N_875,N_974);
nor U1086 (N_1086,N_896,N_970);
nor U1087 (N_1087,N_804,N_990);
and U1088 (N_1088,N_861,N_937);
nand U1089 (N_1089,N_902,N_979);
nand U1090 (N_1090,N_908,N_924);
and U1091 (N_1091,N_915,N_996);
nand U1092 (N_1092,N_941,N_939);
nand U1093 (N_1093,N_948,N_904);
nand U1094 (N_1094,N_980,N_802);
and U1095 (N_1095,N_940,N_829);
nor U1096 (N_1096,N_993,N_997);
nor U1097 (N_1097,N_890,N_803);
and U1098 (N_1098,N_865,N_972);
or U1099 (N_1099,N_955,N_816);
nor U1100 (N_1100,N_811,N_828);
or U1101 (N_1101,N_815,N_946);
nand U1102 (N_1102,N_822,N_963);
or U1103 (N_1103,N_987,N_845);
nand U1104 (N_1104,N_991,N_934);
or U1105 (N_1105,N_913,N_819);
nand U1106 (N_1106,N_997,N_937);
and U1107 (N_1107,N_833,N_841);
nor U1108 (N_1108,N_931,N_831);
and U1109 (N_1109,N_827,N_805);
nor U1110 (N_1110,N_881,N_929);
nand U1111 (N_1111,N_836,N_896);
nor U1112 (N_1112,N_919,N_826);
or U1113 (N_1113,N_831,N_988);
or U1114 (N_1114,N_966,N_937);
and U1115 (N_1115,N_918,N_921);
nand U1116 (N_1116,N_997,N_836);
nand U1117 (N_1117,N_889,N_829);
nand U1118 (N_1118,N_971,N_805);
and U1119 (N_1119,N_920,N_962);
nor U1120 (N_1120,N_923,N_865);
or U1121 (N_1121,N_964,N_917);
and U1122 (N_1122,N_993,N_949);
and U1123 (N_1123,N_976,N_871);
nand U1124 (N_1124,N_852,N_963);
and U1125 (N_1125,N_833,N_886);
and U1126 (N_1126,N_923,N_930);
nand U1127 (N_1127,N_820,N_960);
nand U1128 (N_1128,N_861,N_913);
and U1129 (N_1129,N_900,N_956);
or U1130 (N_1130,N_939,N_870);
nand U1131 (N_1131,N_834,N_896);
and U1132 (N_1132,N_975,N_892);
or U1133 (N_1133,N_951,N_999);
nor U1134 (N_1134,N_957,N_877);
and U1135 (N_1135,N_962,N_901);
nor U1136 (N_1136,N_962,N_806);
nor U1137 (N_1137,N_941,N_812);
or U1138 (N_1138,N_810,N_974);
nor U1139 (N_1139,N_900,N_920);
and U1140 (N_1140,N_855,N_977);
nor U1141 (N_1141,N_838,N_915);
nor U1142 (N_1142,N_942,N_935);
and U1143 (N_1143,N_981,N_911);
nor U1144 (N_1144,N_903,N_923);
or U1145 (N_1145,N_903,N_813);
nor U1146 (N_1146,N_869,N_819);
or U1147 (N_1147,N_927,N_823);
nor U1148 (N_1148,N_902,N_930);
or U1149 (N_1149,N_964,N_832);
or U1150 (N_1150,N_917,N_885);
nand U1151 (N_1151,N_812,N_996);
or U1152 (N_1152,N_820,N_822);
and U1153 (N_1153,N_992,N_828);
or U1154 (N_1154,N_822,N_845);
nand U1155 (N_1155,N_840,N_996);
nand U1156 (N_1156,N_866,N_956);
and U1157 (N_1157,N_929,N_836);
or U1158 (N_1158,N_881,N_996);
nor U1159 (N_1159,N_926,N_936);
or U1160 (N_1160,N_834,N_977);
xor U1161 (N_1161,N_861,N_943);
or U1162 (N_1162,N_932,N_812);
nor U1163 (N_1163,N_885,N_820);
and U1164 (N_1164,N_991,N_866);
nand U1165 (N_1165,N_979,N_831);
nor U1166 (N_1166,N_909,N_832);
nor U1167 (N_1167,N_837,N_940);
or U1168 (N_1168,N_872,N_900);
nand U1169 (N_1169,N_819,N_839);
nand U1170 (N_1170,N_905,N_972);
nand U1171 (N_1171,N_991,N_926);
nor U1172 (N_1172,N_918,N_855);
or U1173 (N_1173,N_952,N_996);
nand U1174 (N_1174,N_896,N_955);
nand U1175 (N_1175,N_938,N_874);
nand U1176 (N_1176,N_983,N_853);
nor U1177 (N_1177,N_991,N_833);
nor U1178 (N_1178,N_880,N_867);
or U1179 (N_1179,N_864,N_936);
or U1180 (N_1180,N_879,N_997);
nand U1181 (N_1181,N_853,N_989);
and U1182 (N_1182,N_871,N_823);
nor U1183 (N_1183,N_836,N_962);
nor U1184 (N_1184,N_815,N_990);
nor U1185 (N_1185,N_895,N_965);
nand U1186 (N_1186,N_825,N_840);
and U1187 (N_1187,N_934,N_946);
or U1188 (N_1188,N_914,N_825);
nor U1189 (N_1189,N_952,N_932);
nand U1190 (N_1190,N_904,N_918);
or U1191 (N_1191,N_990,N_897);
or U1192 (N_1192,N_851,N_939);
nand U1193 (N_1193,N_986,N_954);
or U1194 (N_1194,N_973,N_819);
and U1195 (N_1195,N_838,N_934);
and U1196 (N_1196,N_975,N_954);
or U1197 (N_1197,N_941,N_866);
nor U1198 (N_1198,N_913,N_887);
or U1199 (N_1199,N_818,N_834);
or U1200 (N_1200,N_1179,N_1193);
nor U1201 (N_1201,N_1153,N_1137);
or U1202 (N_1202,N_1104,N_1030);
xor U1203 (N_1203,N_1186,N_1132);
or U1204 (N_1204,N_1065,N_1053);
and U1205 (N_1205,N_1199,N_1139);
and U1206 (N_1206,N_1176,N_1189);
and U1207 (N_1207,N_1047,N_1088);
and U1208 (N_1208,N_1067,N_1172);
nor U1209 (N_1209,N_1049,N_1026);
or U1210 (N_1210,N_1093,N_1009);
nand U1211 (N_1211,N_1044,N_1023);
and U1212 (N_1212,N_1197,N_1083);
and U1213 (N_1213,N_1099,N_1050);
nor U1214 (N_1214,N_1151,N_1159);
and U1215 (N_1215,N_1143,N_1059);
nor U1216 (N_1216,N_1000,N_1082);
nor U1217 (N_1217,N_1100,N_1149);
and U1218 (N_1218,N_1055,N_1058);
nor U1219 (N_1219,N_1070,N_1190);
and U1220 (N_1220,N_1074,N_1158);
nor U1221 (N_1221,N_1195,N_1106);
nand U1222 (N_1222,N_1124,N_1028);
nor U1223 (N_1223,N_1021,N_1069);
nor U1224 (N_1224,N_1146,N_1107);
and U1225 (N_1225,N_1123,N_1043);
nand U1226 (N_1226,N_1012,N_1001);
and U1227 (N_1227,N_1181,N_1163);
and U1228 (N_1228,N_1174,N_1184);
nand U1229 (N_1229,N_1118,N_1114);
nand U1230 (N_1230,N_1024,N_1084);
nand U1231 (N_1231,N_1007,N_1052);
or U1232 (N_1232,N_1073,N_1161);
nor U1233 (N_1233,N_1060,N_1034);
or U1234 (N_1234,N_1020,N_1138);
or U1235 (N_1235,N_1033,N_1041);
nor U1236 (N_1236,N_1017,N_1177);
or U1237 (N_1237,N_1006,N_1131);
nand U1238 (N_1238,N_1182,N_1188);
or U1239 (N_1239,N_1096,N_1031);
or U1240 (N_1240,N_1010,N_1013);
nor U1241 (N_1241,N_1126,N_1016);
and U1242 (N_1242,N_1101,N_1076);
nor U1243 (N_1243,N_1078,N_1122);
nand U1244 (N_1244,N_1160,N_1037);
nand U1245 (N_1245,N_1168,N_1025);
nor U1246 (N_1246,N_1102,N_1022);
and U1247 (N_1247,N_1018,N_1165);
and U1248 (N_1248,N_1135,N_1048);
or U1249 (N_1249,N_1154,N_1064);
nand U1250 (N_1250,N_1117,N_1185);
nor U1251 (N_1251,N_1140,N_1162);
nor U1252 (N_1252,N_1008,N_1136);
or U1253 (N_1253,N_1166,N_1108);
or U1254 (N_1254,N_1128,N_1054);
nand U1255 (N_1255,N_1147,N_1157);
or U1256 (N_1256,N_1068,N_1167);
xor U1257 (N_1257,N_1061,N_1094);
or U1258 (N_1258,N_1175,N_1063);
or U1259 (N_1259,N_1194,N_1192);
nor U1260 (N_1260,N_1112,N_1027);
nand U1261 (N_1261,N_1005,N_1086);
or U1262 (N_1262,N_1040,N_1142);
nor U1263 (N_1263,N_1183,N_1198);
and U1264 (N_1264,N_1089,N_1075);
and U1265 (N_1265,N_1097,N_1191);
or U1266 (N_1266,N_1072,N_1098);
and U1267 (N_1267,N_1056,N_1011);
nand U1268 (N_1268,N_1113,N_1014);
or U1269 (N_1269,N_1103,N_1087);
nand U1270 (N_1270,N_1170,N_1171);
or U1271 (N_1271,N_1071,N_1057);
or U1272 (N_1272,N_1120,N_1145);
nand U1273 (N_1273,N_1111,N_1178);
and U1274 (N_1274,N_1051,N_1127);
and U1275 (N_1275,N_1116,N_1150);
nand U1276 (N_1276,N_1144,N_1085);
nor U1277 (N_1277,N_1019,N_1156);
or U1278 (N_1278,N_1046,N_1134);
nor U1279 (N_1279,N_1105,N_1129);
nor U1280 (N_1280,N_1119,N_1090);
and U1281 (N_1281,N_1148,N_1042);
nand U1282 (N_1282,N_1109,N_1091);
and U1283 (N_1283,N_1173,N_1152);
nor U1284 (N_1284,N_1035,N_1141);
nor U1285 (N_1285,N_1130,N_1164);
nor U1286 (N_1286,N_1077,N_1039);
or U1287 (N_1287,N_1187,N_1029);
nor U1288 (N_1288,N_1045,N_1121);
or U1289 (N_1289,N_1015,N_1092);
or U1290 (N_1290,N_1080,N_1095);
and U1291 (N_1291,N_1079,N_1155);
nand U1292 (N_1292,N_1196,N_1133);
nor U1293 (N_1293,N_1002,N_1169);
nand U1294 (N_1294,N_1038,N_1036);
nor U1295 (N_1295,N_1004,N_1032);
or U1296 (N_1296,N_1110,N_1081);
and U1297 (N_1297,N_1062,N_1066);
or U1298 (N_1298,N_1180,N_1003);
or U1299 (N_1299,N_1125,N_1115);
nand U1300 (N_1300,N_1182,N_1076);
or U1301 (N_1301,N_1111,N_1012);
nand U1302 (N_1302,N_1083,N_1189);
nor U1303 (N_1303,N_1070,N_1030);
nor U1304 (N_1304,N_1144,N_1076);
nand U1305 (N_1305,N_1128,N_1110);
nand U1306 (N_1306,N_1150,N_1152);
or U1307 (N_1307,N_1032,N_1030);
nand U1308 (N_1308,N_1096,N_1158);
and U1309 (N_1309,N_1078,N_1148);
nor U1310 (N_1310,N_1191,N_1137);
xnor U1311 (N_1311,N_1187,N_1152);
or U1312 (N_1312,N_1042,N_1117);
nor U1313 (N_1313,N_1159,N_1184);
nor U1314 (N_1314,N_1130,N_1064);
nand U1315 (N_1315,N_1027,N_1154);
and U1316 (N_1316,N_1111,N_1148);
and U1317 (N_1317,N_1047,N_1004);
and U1318 (N_1318,N_1053,N_1068);
nor U1319 (N_1319,N_1156,N_1134);
nor U1320 (N_1320,N_1090,N_1193);
or U1321 (N_1321,N_1099,N_1066);
and U1322 (N_1322,N_1115,N_1132);
nor U1323 (N_1323,N_1173,N_1052);
nor U1324 (N_1324,N_1155,N_1009);
nor U1325 (N_1325,N_1182,N_1116);
nand U1326 (N_1326,N_1065,N_1088);
and U1327 (N_1327,N_1029,N_1020);
and U1328 (N_1328,N_1002,N_1176);
or U1329 (N_1329,N_1082,N_1175);
and U1330 (N_1330,N_1073,N_1049);
or U1331 (N_1331,N_1095,N_1165);
and U1332 (N_1332,N_1021,N_1172);
nand U1333 (N_1333,N_1116,N_1117);
or U1334 (N_1334,N_1029,N_1132);
and U1335 (N_1335,N_1146,N_1081);
and U1336 (N_1336,N_1121,N_1111);
and U1337 (N_1337,N_1111,N_1133);
nor U1338 (N_1338,N_1099,N_1177);
nor U1339 (N_1339,N_1053,N_1152);
and U1340 (N_1340,N_1109,N_1045);
and U1341 (N_1341,N_1194,N_1102);
nand U1342 (N_1342,N_1120,N_1163);
and U1343 (N_1343,N_1154,N_1151);
and U1344 (N_1344,N_1077,N_1050);
nand U1345 (N_1345,N_1004,N_1037);
and U1346 (N_1346,N_1170,N_1082);
nand U1347 (N_1347,N_1039,N_1122);
and U1348 (N_1348,N_1111,N_1101);
and U1349 (N_1349,N_1153,N_1100);
nand U1350 (N_1350,N_1072,N_1029);
nor U1351 (N_1351,N_1036,N_1183);
and U1352 (N_1352,N_1065,N_1160);
nand U1353 (N_1353,N_1010,N_1083);
and U1354 (N_1354,N_1016,N_1132);
and U1355 (N_1355,N_1035,N_1000);
nor U1356 (N_1356,N_1182,N_1083);
and U1357 (N_1357,N_1135,N_1046);
and U1358 (N_1358,N_1109,N_1039);
and U1359 (N_1359,N_1096,N_1177);
or U1360 (N_1360,N_1130,N_1022);
and U1361 (N_1361,N_1168,N_1035);
and U1362 (N_1362,N_1128,N_1051);
and U1363 (N_1363,N_1164,N_1042);
nor U1364 (N_1364,N_1015,N_1159);
and U1365 (N_1365,N_1173,N_1048);
and U1366 (N_1366,N_1184,N_1106);
nor U1367 (N_1367,N_1001,N_1152);
or U1368 (N_1368,N_1116,N_1003);
nand U1369 (N_1369,N_1066,N_1054);
nor U1370 (N_1370,N_1001,N_1032);
nand U1371 (N_1371,N_1119,N_1122);
nand U1372 (N_1372,N_1060,N_1184);
or U1373 (N_1373,N_1187,N_1079);
nor U1374 (N_1374,N_1078,N_1025);
and U1375 (N_1375,N_1116,N_1178);
or U1376 (N_1376,N_1115,N_1153);
nor U1377 (N_1377,N_1164,N_1119);
or U1378 (N_1378,N_1030,N_1188);
nor U1379 (N_1379,N_1150,N_1026);
and U1380 (N_1380,N_1095,N_1174);
or U1381 (N_1381,N_1025,N_1076);
nand U1382 (N_1382,N_1066,N_1029);
xor U1383 (N_1383,N_1028,N_1003);
and U1384 (N_1384,N_1029,N_1133);
and U1385 (N_1385,N_1008,N_1141);
and U1386 (N_1386,N_1076,N_1108);
and U1387 (N_1387,N_1187,N_1173);
nand U1388 (N_1388,N_1177,N_1178);
nor U1389 (N_1389,N_1005,N_1008);
or U1390 (N_1390,N_1163,N_1108);
or U1391 (N_1391,N_1001,N_1093);
or U1392 (N_1392,N_1080,N_1035);
nor U1393 (N_1393,N_1139,N_1188);
and U1394 (N_1394,N_1014,N_1131);
nand U1395 (N_1395,N_1160,N_1121);
or U1396 (N_1396,N_1170,N_1173);
nand U1397 (N_1397,N_1142,N_1148);
nand U1398 (N_1398,N_1024,N_1096);
nand U1399 (N_1399,N_1088,N_1184);
and U1400 (N_1400,N_1236,N_1331);
nor U1401 (N_1401,N_1365,N_1358);
and U1402 (N_1402,N_1217,N_1354);
and U1403 (N_1403,N_1283,N_1207);
nand U1404 (N_1404,N_1306,N_1270);
and U1405 (N_1405,N_1262,N_1254);
nand U1406 (N_1406,N_1322,N_1332);
and U1407 (N_1407,N_1258,N_1221);
xnor U1408 (N_1408,N_1351,N_1269);
and U1409 (N_1409,N_1321,N_1203);
and U1410 (N_1410,N_1388,N_1230);
nor U1411 (N_1411,N_1211,N_1256);
nor U1412 (N_1412,N_1391,N_1293);
nand U1413 (N_1413,N_1349,N_1288);
nand U1414 (N_1414,N_1341,N_1375);
or U1415 (N_1415,N_1225,N_1235);
or U1416 (N_1416,N_1264,N_1357);
and U1417 (N_1417,N_1324,N_1342);
nor U1418 (N_1418,N_1205,N_1278);
nor U1419 (N_1419,N_1376,N_1366);
nand U1420 (N_1420,N_1316,N_1347);
and U1421 (N_1421,N_1260,N_1378);
or U1422 (N_1422,N_1394,N_1267);
nor U1423 (N_1423,N_1281,N_1265);
or U1424 (N_1424,N_1218,N_1244);
or U1425 (N_1425,N_1319,N_1370);
and U1426 (N_1426,N_1364,N_1372);
nand U1427 (N_1427,N_1362,N_1263);
and U1428 (N_1428,N_1336,N_1215);
and U1429 (N_1429,N_1317,N_1382);
or U1430 (N_1430,N_1326,N_1299);
and U1431 (N_1431,N_1333,N_1222);
and U1432 (N_1432,N_1295,N_1202);
and U1433 (N_1433,N_1253,N_1204);
and U1434 (N_1434,N_1240,N_1396);
nand U1435 (N_1435,N_1355,N_1219);
and U1436 (N_1436,N_1398,N_1252);
nand U1437 (N_1437,N_1369,N_1356);
and U1438 (N_1438,N_1289,N_1329);
and U1439 (N_1439,N_1259,N_1395);
and U1440 (N_1440,N_1373,N_1310);
and U1441 (N_1441,N_1352,N_1387);
nand U1442 (N_1442,N_1266,N_1246);
xor U1443 (N_1443,N_1249,N_1330);
nor U1444 (N_1444,N_1384,N_1314);
or U1445 (N_1445,N_1379,N_1383);
or U1446 (N_1446,N_1271,N_1241);
nand U1447 (N_1447,N_1208,N_1298);
nand U1448 (N_1448,N_1210,N_1304);
nor U1449 (N_1449,N_1377,N_1232);
or U1450 (N_1450,N_1346,N_1272);
or U1451 (N_1451,N_1292,N_1247);
and U1452 (N_1452,N_1325,N_1327);
or U1453 (N_1453,N_1226,N_1268);
and U1454 (N_1454,N_1276,N_1374);
and U1455 (N_1455,N_1243,N_1296);
nand U1456 (N_1456,N_1360,N_1233);
or U1457 (N_1457,N_1335,N_1200);
xnor U1458 (N_1458,N_1274,N_1255);
nor U1459 (N_1459,N_1371,N_1303);
nor U1460 (N_1460,N_1216,N_1353);
nor U1461 (N_1461,N_1343,N_1345);
nand U1462 (N_1462,N_1328,N_1284);
or U1463 (N_1463,N_1359,N_1239);
and U1464 (N_1464,N_1337,N_1250);
nand U1465 (N_1465,N_1311,N_1399);
and U1466 (N_1466,N_1390,N_1285);
and U1467 (N_1467,N_1242,N_1386);
or U1468 (N_1468,N_1231,N_1287);
nand U1469 (N_1469,N_1273,N_1229);
or U1470 (N_1470,N_1368,N_1261);
and U1471 (N_1471,N_1393,N_1313);
or U1472 (N_1472,N_1340,N_1380);
or U1473 (N_1473,N_1397,N_1214);
or U1474 (N_1474,N_1385,N_1251);
nand U1475 (N_1475,N_1275,N_1318);
or U1476 (N_1476,N_1334,N_1257);
and U1477 (N_1477,N_1213,N_1301);
and U1478 (N_1478,N_1320,N_1350);
nand U1479 (N_1479,N_1308,N_1361);
and U1480 (N_1480,N_1279,N_1201);
and U1481 (N_1481,N_1339,N_1302);
nor U1482 (N_1482,N_1323,N_1297);
and U1483 (N_1483,N_1282,N_1227);
and U1484 (N_1484,N_1228,N_1280);
nor U1485 (N_1485,N_1238,N_1392);
nor U1486 (N_1486,N_1245,N_1223);
nor U1487 (N_1487,N_1237,N_1224);
or U1488 (N_1488,N_1290,N_1381);
nand U1489 (N_1489,N_1348,N_1315);
or U1490 (N_1490,N_1212,N_1305);
xnor U1491 (N_1491,N_1307,N_1234);
xnor U1492 (N_1492,N_1338,N_1367);
nor U1493 (N_1493,N_1206,N_1300);
and U1494 (N_1494,N_1248,N_1209);
xor U1495 (N_1495,N_1294,N_1220);
nor U1496 (N_1496,N_1344,N_1291);
or U1497 (N_1497,N_1312,N_1286);
nand U1498 (N_1498,N_1277,N_1389);
or U1499 (N_1499,N_1363,N_1309);
and U1500 (N_1500,N_1294,N_1289);
nor U1501 (N_1501,N_1252,N_1222);
or U1502 (N_1502,N_1241,N_1311);
and U1503 (N_1503,N_1217,N_1388);
and U1504 (N_1504,N_1342,N_1280);
and U1505 (N_1505,N_1251,N_1380);
nor U1506 (N_1506,N_1208,N_1288);
or U1507 (N_1507,N_1349,N_1203);
nand U1508 (N_1508,N_1305,N_1304);
nor U1509 (N_1509,N_1359,N_1324);
and U1510 (N_1510,N_1239,N_1210);
nor U1511 (N_1511,N_1310,N_1292);
and U1512 (N_1512,N_1275,N_1235);
nand U1513 (N_1513,N_1346,N_1377);
and U1514 (N_1514,N_1228,N_1311);
and U1515 (N_1515,N_1216,N_1211);
and U1516 (N_1516,N_1364,N_1278);
or U1517 (N_1517,N_1217,N_1257);
nor U1518 (N_1518,N_1232,N_1310);
and U1519 (N_1519,N_1318,N_1295);
or U1520 (N_1520,N_1206,N_1282);
or U1521 (N_1521,N_1242,N_1380);
nand U1522 (N_1522,N_1276,N_1317);
or U1523 (N_1523,N_1392,N_1207);
or U1524 (N_1524,N_1336,N_1349);
or U1525 (N_1525,N_1295,N_1353);
nand U1526 (N_1526,N_1370,N_1375);
nand U1527 (N_1527,N_1320,N_1318);
and U1528 (N_1528,N_1340,N_1363);
or U1529 (N_1529,N_1390,N_1361);
nor U1530 (N_1530,N_1307,N_1274);
nor U1531 (N_1531,N_1217,N_1328);
nor U1532 (N_1532,N_1371,N_1297);
and U1533 (N_1533,N_1357,N_1390);
or U1534 (N_1534,N_1200,N_1264);
xor U1535 (N_1535,N_1398,N_1255);
or U1536 (N_1536,N_1343,N_1212);
nor U1537 (N_1537,N_1269,N_1239);
and U1538 (N_1538,N_1325,N_1315);
or U1539 (N_1539,N_1351,N_1295);
and U1540 (N_1540,N_1377,N_1331);
or U1541 (N_1541,N_1231,N_1370);
nor U1542 (N_1542,N_1373,N_1336);
or U1543 (N_1543,N_1235,N_1315);
or U1544 (N_1544,N_1369,N_1214);
or U1545 (N_1545,N_1335,N_1246);
nor U1546 (N_1546,N_1345,N_1370);
nor U1547 (N_1547,N_1211,N_1301);
or U1548 (N_1548,N_1271,N_1219);
nand U1549 (N_1549,N_1313,N_1368);
nor U1550 (N_1550,N_1342,N_1230);
or U1551 (N_1551,N_1263,N_1334);
or U1552 (N_1552,N_1284,N_1286);
or U1553 (N_1553,N_1342,N_1257);
or U1554 (N_1554,N_1286,N_1309);
and U1555 (N_1555,N_1359,N_1293);
nand U1556 (N_1556,N_1213,N_1310);
or U1557 (N_1557,N_1329,N_1242);
nor U1558 (N_1558,N_1300,N_1301);
nor U1559 (N_1559,N_1376,N_1244);
or U1560 (N_1560,N_1218,N_1255);
xor U1561 (N_1561,N_1251,N_1209);
and U1562 (N_1562,N_1310,N_1369);
or U1563 (N_1563,N_1390,N_1380);
or U1564 (N_1564,N_1311,N_1306);
nand U1565 (N_1565,N_1200,N_1372);
nand U1566 (N_1566,N_1344,N_1314);
or U1567 (N_1567,N_1201,N_1211);
nand U1568 (N_1568,N_1249,N_1231);
nand U1569 (N_1569,N_1306,N_1251);
or U1570 (N_1570,N_1286,N_1298);
nor U1571 (N_1571,N_1321,N_1216);
nor U1572 (N_1572,N_1366,N_1374);
nand U1573 (N_1573,N_1287,N_1385);
nor U1574 (N_1574,N_1200,N_1222);
or U1575 (N_1575,N_1344,N_1332);
and U1576 (N_1576,N_1247,N_1248);
nand U1577 (N_1577,N_1271,N_1374);
or U1578 (N_1578,N_1348,N_1218);
nand U1579 (N_1579,N_1218,N_1257);
or U1580 (N_1580,N_1204,N_1393);
and U1581 (N_1581,N_1313,N_1264);
and U1582 (N_1582,N_1222,N_1208);
and U1583 (N_1583,N_1383,N_1349);
xor U1584 (N_1584,N_1373,N_1347);
nor U1585 (N_1585,N_1322,N_1218);
or U1586 (N_1586,N_1294,N_1357);
or U1587 (N_1587,N_1387,N_1317);
or U1588 (N_1588,N_1392,N_1326);
nor U1589 (N_1589,N_1337,N_1304);
or U1590 (N_1590,N_1253,N_1289);
or U1591 (N_1591,N_1280,N_1254);
or U1592 (N_1592,N_1384,N_1219);
or U1593 (N_1593,N_1290,N_1263);
nand U1594 (N_1594,N_1289,N_1352);
and U1595 (N_1595,N_1396,N_1223);
nand U1596 (N_1596,N_1398,N_1321);
or U1597 (N_1597,N_1237,N_1280);
nor U1598 (N_1598,N_1393,N_1248);
nand U1599 (N_1599,N_1263,N_1342);
and U1600 (N_1600,N_1520,N_1598);
and U1601 (N_1601,N_1545,N_1517);
nor U1602 (N_1602,N_1479,N_1472);
nor U1603 (N_1603,N_1585,N_1469);
nor U1604 (N_1604,N_1418,N_1578);
or U1605 (N_1605,N_1411,N_1522);
or U1606 (N_1606,N_1549,N_1551);
nand U1607 (N_1607,N_1535,N_1519);
and U1608 (N_1608,N_1471,N_1496);
or U1609 (N_1609,N_1476,N_1534);
nor U1610 (N_1610,N_1499,N_1502);
nor U1611 (N_1611,N_1468,N_1581);
nand U1612 (N_1612,N_1402,N_1452);
nand U1613 (N_1613,N_1547,N_1554);
nor U1614 (N_1614,N_1435,N_1597);
nand U1615 (N_1615,N_1481,N_1407);
and U1616 (N_1616,N_1459,N_1580);
nor U1617 (N_1617,N_1512,N_1406);
nand U1618 (N_1618,N_1445,N_1492);
or U1619 (N_1619,N_1414,N_1465);
and U1620 (N_1620,N_1579,N_1446);
nand U1621 (N_1621,N_1582,N_1555);
nand U1622 (N_1622,N_1436,N_1498);
nor U1623 (N_1623,N_1576,N_1574);
nor U1624 (N_1624,N_1557,N_1569);
and U1625 (N_1625,N_1403,N_1430);
nor U1626 (N_1626,N_1490,N_1537);
nand U1627 (N_1627,N_1477,N_1428);
nor U1628 (N_1628,N_1521,N_1575);
xnor U1629 (N_1629,N_1475,N_1412);
and U1630 (N_1630,N_1586,N_1480);
nand U1631 (N_1631,N_1592,N_1553);
and U1632 (N_1632,N_1536,N_1437);
nor U1633 (N_1633,N_1530,N_1563);
xnor U1634 (N_1634,N_1462,N_1599);
nor U1635 (N_1635,N_1429,N_1419);
nor U1636 (N_1636,N_1516,N_1506);
or U1637 (N_1637,N_1415,N_1421);
nand U1638 (N_1638,N_1562,N_1556);
and U1639 (N_1639,N_1482,N_1489);
or U1640 (N_1640,N_1433,N_1432);
or U1641 (N_1641,N_1427,N_1561);
xnor U1642 (N_1642,N_1588,N_1447);
and U1643 (N_1643,N_1552,N_1596);
and U1644 (N_1644,N_1423,N_1441);
or U1645 (N_1645,N_1526,N_1457);
and U1646 (N_1646,N_1495,N_1568);
or U1647 (N_1647,N_1509,N_1449);
and U1648 (N_1648,N_1529,N_1484);
nand U1649 (N_1649,N_1400,N_1500);
nand U1650 (N_1650,N_1405,N_1450);
nor U1651 (N_1651,N_1528,N_1464);
nor U1652 (N_1652,N_1542,N_1525);
nor U1653 (N_1653,N_1571,N_1497);
or U1654 (N_1654,N_1548,N_1559);
or U1655 (N_1655,N_1453,N_1558);
or U1656 (N_1656,N_1514,N_1560);
nor U1657 (N_1657,N_1461,N_1417);
and U1658 (N_1658,N_1513,N_1463);
nand U1659 (N_1659,N_1404,N_1564);
nand U1660 (N_1660,N_1456,N_1587);
nor U1661 (N_1661,N_1572,N_1511);
and U1662 (N_1662,N_1584,N_1420);
nor U1663 (N_1663,N_1487,N_1422);
nor U1664 (N_1664,N_1533,N_1409);
nand U1665 (N_1665,N_1458,N_1442);
or U1666 (N_1666,N_1425,N_1493);
and U1667 (N_1667,N_1505,N_1508);
xnor U1668 (N_1668,N_1485,N_1532);
and U1669 (N_1669,N_1410,N_1455);
nand U1670 (N_1670,N_1518,N_1565);
or U1671 (N_1671,N_1538,N_1444);
nand U1672 (N_1672,N_1591,N_1590);
or U1673 (N_1673,N_1491,N_1573);
nand U1674 (N_1674,N_1589,N_1546);
and U1675 (N_1675,N_1583,N_1577);
and U1676 (N_1676,N_1474,N_1570);
and U1677 (N_1677,N_1567,N_1544);
nor U1678 (N_1678,N_1466,N_1540);
nand U1679 (N_1679,N_1467,N_1594);
and U1680 (N_1680,N_1454,N_1443);
or U1681 (N_1681,N_1483,N_1448);
nand U1682 (N_1682,N_1523,N_1501);
or U1683 (N_1683,N_1527,N_1504);
nor U1684 (N_1684,N_1470,N_1541);
and U1685 (N_1685,N_1478,N_1440);
or U1686 (N_1686,N_1595,N_1550);
nand U1687 (N_1687,N_1416,N_1401);
nor U1688 (N_1688,N_1531,N_1543);
nor U1689 (N_1689,N_1515,N_1494);
xnor U1690 (N_1690,N_1413,N_1431);
or U1691 (N_1691,N_1507,N_1438);
nor U1692 (N_1692,N_1451,N_1424);
nor U1693 (N_1693,N_1473,N_1439);
nor U1694 (N_1694,N_1408,N_1426);
nor U1695 (N_1695,N_1593,N_1488);
nand U1696 (N_1696,N_1503,N_1566);
or U1697 (N_1697,N_1486,N_1524);
and U1698 (N_1698,N_1434,N_1460);
or U1699 (N_1699,N_1510,N_1539);
nor U1700 (N_1700,N_1563,N_1568);
nor U1701 (N_1701,N_1581,N_1446);
or U1702 (N_1702,N_1419,N_1502);
or U1703 (N_1703,N_1405,N_1436);
nand U1704 (N_1704,N_1483,N_1579);
nor U1705 (N_1705,N_1555,N_1527);
nor U1706 (N_1706,N_1425,N_1551);
nor U1707 (N_1707,N_1486,N_1551);
nor U1708 (N_1708,N_1594,N_1413);
or U1709 (N_1709,N_1475,N_1426);
nand U1710 (N_1710,N_1452,N_1519);
nor U1711 (N_1711,N_1495,N_1490);
nand U1712 (N_1712,N_1498,N_1486);
nand U1713 (N_1713,N_1502,N_1525);
or U1714 (N_1714,N_1451,N_1433);
or U1715 (N_1715,N_1565,N_1569);
nor U1716 (N_1716,N_1477,N_1487);
nand U1717 (N_1717,N_1571,N_1512);
nor U1718 (N_1718,N_1402,N_1496);
and U1719 (N_1719,N_1595,N_1434);
and U1720 (N_1720,N_1412,N_1503);
nand U1721 (N_1721,N_1494,N_1498);
nand U1722 (N_1722,N_1431,N_1509);
xnor U1723 (N_1723,N_1474,N_1547);
and U1724 (N_1724,N_1564,N_1516);
nor U1725 (N_1725,N_1423,N_1466);
nand U1726 (N_1726,N_1537,N_1581);
and U1727 (N_1727,N_1436,N_1403);
or U1728 (N_1728,N_1464,N_1523);
and U1729 (N_1729,N_1442,N_1497);
nand U1730 (N_1730,N_1585,N_1461);
xnor U1731 (N_1731,N_1535,N_1400);
nand U1732 (N_1732,N_1528,N_1502);
and U1733 (N_1733,N_1502,N_1510);
or U1734 (N_1734,N_1442,N_1436);
nor U1735 (N_1735,N_1576,N_1513);
and U1736 (N_1736,N_1590,N_1423);
and U1737 (N_1737,N_1587,N_1420);
nand U1738 (N_1738,N_1439,N_1467);
nand U1739 (N_1739,N_1414,N_1516);
nand U1740 (N_1740,N_1554,N_1431);
nor U1741 (N_1741,N_1431,N_1534);
nor U1742 (N_1742,N_1520,N_1477);
nor U1743 (N_1743,N_1548,N_1530);
nor U1744 (N_1744,N_1541,N_1464);
nor U1745 (N_1745,N_1589,N_1567);
xnor U1746 (N_1746,N_1536,N_1564);
and U1747 (N_1747,N_1480,N_1524);
or U1748 (N_1748,N_1530,N_1419);
nor U1749 (N_1749,N_1428,N_1441);
nor U1750 (N_1750,N_1438,N_1411);
or U1751 (N_1751,N_1470,N_1454);
nand U1752 (N_1752,N_1521,N_1478);
or U1753 (N_1753,N_1570,N_1409);
and U1754 (N_1754,N_1454,N_1576);
and U1755 (N_1755,N_1428,N_1548);
or U1756 (N_1756,N_1481,N_1484);
nor U1757 (N_1757,N_1500,N_1549);
nand U1758 (N_1758,N_1484,N_1431);
and U1759 (N_1759,N_1442,N_1481);
and U1760 (N_1760,N_1414,N_1447);
nor U1761 (N_1761,N_1442,N_1433);
or U1762 (N_1762,N_1450,N_1493);
nor U1763 (N_1763,N_1527,N_1482);
and U1764 (N_1764,N_1556,N_1436);
nand U1765 (N_1765,N_1521,N_1435);
nand U1766 (N_1766,N_1441,N_1470);
or U1767 (N_1767,N_1542,N_1494);
and U1768 (N_1768,N_1513,N_1554);
or U1769 (N_1769,N_1474,N_1443);
nand U1770 (N_1770,N_1412,N_1429);
and U1771 (N_1771,N_1534,N_1537);
nand U1772 (N_1772,N_1422,N_1434);
nor U1773 (N_1773,N_1403,N_1545);
nor U1774 (N_1774,N_1445,N_1407);
or U1775 (N_1775,N_1470,N_1419);
nand U1776 (N_1776,N_1538,N_1470);
or U1777 (N_1777,N_1505,N_1543);
or U1778 (N_1778,N_1479,N_1572);
or U1779 (N_1779,N_1497,N_1552);
and U1780 (N_1780,N_1547,N_1473);
and U1781 (N_1781,N_1500,N_1557);
or U1782 (N_1782,N_1598,N_1591);
and U1783 (N_1783,N_1413,N_1448);
nand U1784 (N_1784,N_1521,N_1546);
or U1785 (N_1785,N_1568,N_1447);
or U1786 (N_1786,N_1510,N_1537);
or U1787 (N_1787,N_1574,N_1468);
and U1788 (N_1788,N_1596,N_1577);
nand U1789 (N_1789,N_1544,N_1546);
and U1790 (N_1790,N_1511,N_1440);
or U1791 (N_1791,N_1451,N_1508);
or U1792 (N_1792,N_1528,N_1530);
and U1793 (N_1793,N_1497,N_1551);
and U1794 (N_1794,N_1524,N_1444);
or U1795 (N_1795,N_1590,N_1427);
nand U1796 (N_1796,N_1427,N_1598);
or U1797 (N_1797,N_1448,N_1555);
nor U1798 (N_1798,N_1571,N_1509);
nand U1799 (N_1799,N_1572,N_1431);
nand U1800 (N_1800,N_1625,N_1757);
nor U1801 (N_1801,N_1751,N_1613);
nand U1802 (N_1802,N_1748,N_1752);
nand U1803 (N_1803,N_1687,N_1614);
nand U1804 (N_1804,N_1643,N_1727);
or U1805 (N_1805,N_1698,N_1713);
nand U1806 (N_1806,N_1773,N_1780);
nand U1807 (N_1807,N_1769,N_1641);
or U1808 (N_1808,N_1674,N_1671);
nor U1809 (N_1809,N_1706,N_1718);
or U1810 (N_1810,N_1694,N_1646);
nand U1811 (N_1811,N_1719,N_1663);
or U1812 (N_1812,N_1654,N_1606);
nand U1813 (N_1813,N_1618,N_1605);
or U1814 (N_1814,N_1729,N_1631);
nor U1815 (N_1815,N_1709,N_1699);
nor U1816 (N_1816,N_1602,N_1695);
and U1817 (N_1817,N_1610,N_1622);
or U1818 (N_1818,N_1788,N_1761);
and U1819 (N_1819,N_1783,N_1647);
nand U1820 (N_1820,N_1691,N_1794);
nor U1821 (N_1821,N_1630,N_1796);
nor U1822 (N_1822,N_1722,N_1658);
nor U1823 (N_1823,N_1735,N_1707);
or U1824 (N_1824,N_1758,N_1710);
and U1825 (N_1825,N_1638,N_1633);
nor U1826 (N_1826,N_1798,N_1785);
nor U1827 (N_1827,N_1669,N_1664);
xor U1828 (N_1828,N_1702,N_1704);
or U1829 (N_1829,N_1790,N_1701);
nor U1830 (N_1830,N_1665,N_1697);
and U1831 (N_1831,N_1730,N_1755);
nor U1832 (N_1832,N_1734,N_1717);
and U1833 (N_1833,N_1703,N_1753);
nand U1834 (N_1834,N_1608,N_1648);
or U1835 (N_1835,N_1771,N_1635);
nor U1836 (N_1836,N_1637,N_1781);
or U1837 (N_1837,N_1711,N_1675);
or U1838 (N_1838,N_1624,N_1672);
nor U1839 (N_1839,N_1720,N_1607);
nand U1840 (N_1840,N_1793,N_1621);
nor U1841 (N_1841,N_1600,N_1673);
nor U1842 (N_1842,N_1705,N_1726);
or U1843 (N_1843,N_1666,N_1649);
nor U1844 (N_1844,N_1745,N_1740);
nor U1845 (N_1845,N_1682,N_1733);
nand U1846 (N_1846,N_1723,N_1668);
and U1847 (N_1847,N_1779,N_1656);
and U1848 (N_1848,N_1689,N_1609);
nor U1849 (N_1849,N_1746,N_1728);
or U1850 (N_1850,N_1651,N_1667);
and U1851 (N_1851,N_1775,N_1679);
nor U1852 (N_1852,N_1678,N_1712);
nor U1853 (N_1853,N_1677,N_1611);
and U1854 (N_1854,N_1716,N_1708);
and U1855 (N_1855,N_1741,N_1604);
or U1856 (N_1856,N_1736,N_1767);
nand U1857 (N_1857,N_1670,N_1680);
nand U1858 (N_1858,N_1778,N_1784);
and U1859 (N_1859,N_1636,N_1681);
nor U1860 (N_1860,N_1685,N_1714);
nor U1861 (N_1861,N_1776,N_1661);
or U1862 (N_1862,N_1616,N_1747);
or U1863 (N_1863,N_1766,N_1696);
nor U1864 (N_1864,N_1615,N_1688);
and U1865 (N_1865,N_1692,N_1676);
or U1866 (N_1866,N_1744,N_1617);
nand U1867 (N_1867,N_1652,N_1662);
nor U1868 (N_1868,N_1655,N_1626);
nor U1869 (N_1869,N_1645,N_1724);
nand U1870 (N_1870,N_1737,N_1619);
and U1871 (N_1871,N_1690,N_1777);
nor U1872 (N_1872,N_1759,N_1772);
nor U1873 (N_1873,N_1686,N_1763);
nor U1874 (N_1874,N_1715,N_1725);
nor U1875 (N_1875,N_1623,N_1693);
nand U1876 (N_1876,N_1603,N_1762);
and U1877 (N_1877,N_1743,N_1756);
or U1878 (N_1878,N_1650,N_1639);
nand U1879 (N_1879,N_1601,N_1742);
nor U1880 (N_1880,N_1774,N_1731);
and U1881 (N_1881,N_1732,N_1786);
or U1882 (N_1882,N_1765,N_1754);
nor U1883 (N_1883,N_1684,N_1739);
nor U1884 (N_1884,N_1789,N_1787);
nor U1885 (N_1885,N_1683,N_1760);
and U1886 (N_1886,N_1797,N_1640);
or U1887 (N_1887,N_1612,N_1749);
and U1888 (N_1888,N_1792,N_1620);
or U1889 (N_1889,N_1764,N_1795);
and U1890 (N_1890,N_1642,N_1627);
or U1891 (N_1891,N_1659,N_1653);
nand U1892 (N_1892,N_1738,N_1632);
nand U1893 (N_1893,N_1750,N_1768);
nor U1894 (N_1894,N_1628,N_1629);
or U1895 (N_1895,N_1660,N_1782);
nor U1896 (N_1896,N_1770,N_1700);
and U1897 (N_1897,N_1791,N_1721);
nand U1898 (N_1898,N_1634,N_1657);
or U1899 (N_1899,N_1644,N_1799);
or U1900 (N_1900,N_1657,N_1724);
nand U1901 (N_1901,N_1758,N_1675);
and U1902 (N_1902,N_1775,N_1742);
and U1903 (N_1903,N_1747,N_1738);
or U1904 (N_1904,N_1777,N_1615);
and U1905 (N_1905,N_1785,N_1743);
or U1906 (N_1906,N_1650,N_1670);
and U1907 (N_1907,N_1646,N_1664);
nor U1908 (N_1908,N_1664,N_1625);
and U1909 (N_1909,N_1696,N_1622);
or U1910 (N_1910,N_1634,N_1770);
and U1911 (N_1911,N_1785,N_1654);
nor U1912 (N_1912,N_1793,N_1771);
and U1913 (N_1913,N_1765,N_1712);
nor U1914 (N_1914,N_1745,N_1624);
nor U1915 (N_1915,N_1729,N_1675);
nor U1916 (N_1916,N_1619,N_1769);
or U1917 (N_1917,N_1658,N_1709);
and U1918 (N_1918,N_1637,N_1654);
and U1919 (N_1919,N_1643,N_1750);
nor U1920 (N_1920,N_1790,N_1669);
nor U1921 (N_1921,N_1728,N_1768);
or U1922 (N_1922,N_1613,N_1606);
nand U1923 (N_1923,N_1658,N_1747);
nor U1924 (N_1924,N_1738,N_1798);
and U1925 (N_1925,N_1788,N_1717);
nor U1926 (N_1926,N_1723,N_1664);
or U1927 (N_1927,N_1765,N_1745);
nor U1928 (N_1928,N_1718,N_1756);
or U1929 (N_1929,N_1682,N_1606);
or U1930 (N_1930,N_1734,N_1635);
or U1931 (N_1931,N_1610,N_1745);
nand U1932 (N_1932,N_1749,N_1668);
and U1933 (N_1933,N_1624,N_1768);
and U1934 (N_1934,N_1778,N_1613);
or U1935 (N_1935,N_1670,N_1616);
nand U1936 (N_1936,N_1715,N_1686);
nand U1937 (N_1937,N_1791,N_1607);
and U1938 (N_1938,N_1616,N_1606);
or U1939 (N_1939,N_1665,N_1612);
and U1940 (N_1940,N_1750,N_1625);
and U1941 (N_1941,N_1627,N_1658);
nand U1942 (N_1942,N_1694,N_1751);
xnor U1943 (N_1943,N_1675,N_1683);
xor U1944 (N_1944,N_1625,N_1718);
and U1945 (N_1945,N_1791,N_1744);
nor U1946 (N_1946,N_1701,N_1631);
nor U1947 (N_1947,N_1741,N_1792);
or U1948 (N_1948,N_1736,N_1777);
nor U1949 (N_1949,N_1697,N_1620);
nand U1950 (N_1950,N_1601,N_1664);
and U1951 (N_1951,N_1786,N_1668);
nor U1952 (N_1952,N_1764,N_1746);
or U1953 (N_1953,N_1659,N_1795);
nand U1954 (N_1954,N_1747,N_1603);
and U1955 (N_1955,N_1644,N_1697);
and U1956 (N_1956,N_1728,N_1790);
nor U1957 (N_1957,N_1789,N_1726);
and U1958 (N_1958,N_1678,N_1759);
nand U1959 (N_1959,N_1609,N_1657);
nand U1960 (N_1960,N_1784,N_1634);
and U1961 (N_1961,N_1610,N_1629);
nor U1962 (N_1962,N_1738,N_1613);
or U1963 (N_1963,N_1633,N_1731);
or U1964 (N_1964,N_1790,N_1680);
or U1965 (N_1965,N_1618,N_1667);
or U1966 (N_1966,N_1639,N_1691);
nor U1967 (N_1967,N_1621,N_1664);
or U1968 (N_1968,N_1723,N_1666);
or U1969 (N_1969,N_1682,N_1711);
nand U1970 (N_1970,N_1685,N_1705);
or U1971 (N_1971,N_1762,N_1731);
nand U1972 (N_1972,N_1726,N_1718);
nand U1973 (N_1973,N_1671,N_1630);
nor U1974 (N_1974,N_1712,N_1621);
and U1975 (N_1975,N_1728,N_1722);
nor U1976 (N_1976,N_1729,N_1706);
and U1977 (N_1977,N_1731,N_1643);
or U1978 (N_1978,N_1615,N_1651);
nor U1979 (N_1979,N_1619,N_1799);
or U1980 (N_1980,N_1797,N_1657);
and U1981 (N_1981,N_1690,N_1602);
nand U1982 (N_1982,N_1690,N_1672);
or U1983 (N_1983,N_1699,N_1798);
and U1984 (N_1984,N_1610,N_1683);
and U1985 (N_1985,N_1737,N_1611);
nand U1986 (N_1986,N_1786,N_1736);
nor U1987 (N_1987,N_1618,N_1631);
nor U1988 (N_1988,N_1759,N_1679);
xor U1989 (N_1989,N_1664,N_1697);
nor U1990 (N_1990,N_1777,N_1694);
nand U1991 (N_1991,N_1614,N_1698);
and U1992 (N_1992,N_1728,N_1719);
nor U1993 (N_1993,N_1796,N_1661);
nor U1994 (N_1994,N_1796,N_1705);
nor U1995 (N_1995,N_1739,N_1617);
nor U1996 (N_1996,N_1714,N_1630);
nand U1997 (N_1997,N_1686,N_1657);
nand U1998 (N_1998,N_1623,N_1694);
or U1999 (N_1999,N_1611,N_1675);
nor U2000 (N_2000,N_1812,N_1985);
and U2001 (N_2001,N_1900,N_1882);
or U2002 (N_2002,N_1859,N_1866);
and U2003 (N_2003,N_1967,N_1902);
nand U2004 (N_2004,N_1935,N_1818);
or U2005 (N_2005,N_1986,N_1861);
nand U2006 (N_2006,N_1903,N_1981);
or U2007 (N_2007,N_1850,N_1845);
and U2008 (N_2008,N_1831,N_1933);
nand U2009 (N_2009,N_1885,N_1990);
nand U2010 (N_2010,N_1929,N_1855);
and U2011 (N_2011,N_1854,N_1833);
and U2012 (N_2012,N_1946,N_1975);
nor U2013 (N_2013,N_1901,N_1931);
nor U2014 (N_2014,N_1846,N_1991);
or U2015 (N_2015,N_1844,N_1879);
nand U2016 (N_2016,N_1955,N_1875);
and U2017 (N_2017,N_1966,N_1948);
and U2018 (N_2018,N_1964,N_1880);
nor U2019 (N_2019,N_1994,N_1807);
nand U2020 (N_2020,N_1883,N_1957);
nor U2021 (N_2021,N_1837,N_1814);
or U2022 (N_2022,N_1950,N_1830);
and U2023 (N_2023,N_1801,N_1871);
nor U2024 (N_2024,N_1851,N_1932);
or U2025 (N_2025,N_1965,N_1840);
or U2026 (N_2026,N_1881,N_1978);
nand U2027 (N_2027,N_1824,N_1984);
nand U2028 (N_2028,N_1823,N_1825);
nor U2029 (N_2029,N_1916,N_1813);
and U2030 (N_2030,N_1923,N_1888);
and U2031 (N_2031,N_1977,N_1834);
xnor U2032 (N_2032,N_1887,N_1805);
or U2033 (N_2033,N_1853,N_1997);
nand U2034 (N_2034,N_1951,N_1921);
xor U2035 (N_2035,N_1826,N_1872);
or U2036 (N_2036,N_1922,N_1918);
or U2037 (N_2037,N_1877,N_1941);
nand U2038 (N_2038,N_1940,N_1949);
nand U2039 (N_2039,N_1862,N_1827);
or U2040 (N_2040,N_1804,N_1962);
or U2041 (N_2041,N_1927,N_1856);
xnor U2042 (N_2042,N_1808,N_1863);
nand U2043 (N_2043,N_1996,N_1947);
nand U2044 (N_2044,N_1806,N_1852);
or U2045 (N_2045,N_1843,N_1904);
or U2046 (N_2046,N_1954,N_1884);
or U2047 (N_2047,N_1993,N_1820);
nand U2048 (N_2048,N_1868,N_1809);
or U2049 (N_2049,N_1930,N_1971);
and U2050 (N_2050,N_1972,N_1945);
and U2051 (N_2051,N_1956,N_1810);
and U2052 (N_2052,N_1998,N_1889);
nand U2053 (N_2053,N_1995,N_1928);
and U2054 (N_2054,N_1961,N_1802);
nor U2055 (N_2055,N_1944,N_1829);
and U2056 (N_2056,N_1943,N_1913);
nor U2057 (N_2057,N_1867,N_1937);
nand U2058 (N_2058,N_1987,N_1907);
nor U2059 (N_2059,N_1963,N_1917);
nand U2060 (N_2060,N_1980,N_1847);
xnor U2061 (N_2061,N_1910,N_1999);
and U2062 (N_2062,N_1973,N_1870);
nor U2063 (N_2063,N_1878,N_1938);
or U2064 (N_2064,N_1969,N_1970);
nor U2065 (N_2065,N_1894,N_1936);
nand U2066 (N_2066,N_1815,N_1925);
and U2067 (N_2067,N_1912,N_1821);
xor U2068 (N_2068,N_1968,N_1836);
or U2069 (N_2069,N_1899,N_1891);
and U2070 (N_2070,N_1895,N_1819);
nand U2071 (N_2071,N_1890,N_1828);
nand U2072 (N_2072,N_1911,N_1835);
nor U2073 (N_2073,N_1905,N_1893);
or U2074 (N_2074,N_1974,N_1915);
nor U2075 (N_2075,N_1838,N_1920);
or U2076 (N_2076,N_1934,N_1869);
and U2077 (N_2077,N_1816,N_1839);
xor U2078 (N_2078,N_1860,N_1926);
or U2079 (N_2079,N_1857,N_1989);
nor U2080 (N_2080,N_1960,N_1992);
nand U2081 (N_2081,N_1886,N_1953);
nand U2082 (N_2082,N_1873,N_1924);
nand U2083 (N_2083,N_1909,N_1803);
nor U2084 (N_2084,N_1914,N_1892);
and U2085 (N_2085,N_1874,N_1939);
or U2086 (N_2086,N_1919,N_1876);
or U2087 (N_2087,N_1842,N_1952);
and U2088 (N_2088,N_1822,N_1908);
nand U2089 (N_2089,N_1959,N_1976);
nand U2090 (N_2090,N_1942,N_1906);
and U2091 (N_2091,N_1988,N_1848);
nor U2092 (N_2092,N_1958,N_1898);
and U2093 (N_2093,N_1841,N_1811);
nand U2094 (N_2094,N_1858,N_1865);
or U2095 (N_2095,N_1983,N_1817);
or U2096 (N_2096,N_1896,N_1864);
and U2097 (N_2097,N_1849,N_1979);
nand U2098 (N_2098,N_1832,N_1982);
or U2099 (N_2099,N_1897,N_1800);
and U2100 (N_2100,N_1822,N_1846);
or U2101 (N_2101,N_1818,N_1902);
or U2102 (N_2102,N_1905,N_1924);
or U2103 (N_2103,N_1856,N_1833);
nor U2104 (N_2104,N_1821,N_1865);
nor U2105 (N_2105,N_1984,N_1845);
and U2106 (N_2106,N_1830,N_1834);
and U2107 (N_2107,N_1943,N_1813);
or U2108 (N_2108,N_1839,N_1937);
and U2109 (N_2109,N_1942,N_1979);
and U2110 (N_2110,N_1880,N_1819);
or U2111 (N_2111,N_1974,N_1885);
and U2112 (N_2112,N_1826,N_1828);
and U2113 (N_2113,N_1862,N_1861);
nor U2114 (N_2114,N_1809,N_1941);
nand U2115 (N_2115,N_1986,N_1923);
and U2116 (N_2116,N_1998,N_1919);
nand U2117 (N_2117,N_1907,N_1802);
nand U2118 (N_2118,N_1909,N_1964);
and U2119 (N_2119,N_1984,N_1865);
or U2120 (N_2120,N_1987,N_1867);
nand U2121 (N_2121,N_1875,N_1969);
and U2122 (N_2122,N_1924,N_1964);
nand U2123 (N_2123,N_1936,N_1811);
nor U2124 (N_2124,N_1919,N_1831);
nor U2125 (N_2125,N_1830,N_1852);
or U2126 (N_2126,N_1878,N_1894);
nor U2127 (N_2127,N_1922,N_1823);
nor U2128 (N_2128,N_1859,N_1854);
or U2129 (N_2129,N_1802,N_1973);
nand U2130 (N_2130,N_1841,N_1981);
and U2131 (N_2131,N_1915,N_1883);
and U2132 (N_2132,N_1936,N_1907);
nor U2133 (N_2133,N_1881,N_1845);
nor U2134 (N_2134,N_1932,N_1808);
and U2135 (N_2135,N_1837,N_1877);
and U2136 (N_2136,N_1917,N_1970);
and U2137 (N_2137,N_1842,N_1828);
and U2138 (N_2138,N_1811,N_1900);
or U2139 (N_2139,N_1979,N_1994);
and U2140 (N_2140,N_1937,N_1979);
nor U2141 (N_2141,N_1840,N_1918);
or U2142 (N_2142,N_1961,N_1868);
and U2143 (N_2143,N_1877,N_1893);
nor U2144 (N_2144,N_1927,N_1853);
nand U2145 (N_2145,N_1935,N_1805);
or U2146 (N_2146,N_1910,N_1822);
nor U2147 (N_2147,N_1836,N_1996);
nor U2148 (N_2148,N_1858,N_1877);
nand U2149 (N_2149,N_1861,N_1867);
and U2150 (N_2150,N_1907,N_1949);
and U2151 (N_2151,N_1922,N_1911);
nand U2152 (N_2152,N_1829,N_1978);
nor U2153 (N_2153,N_1930,N_1803);
nand U2154 (N_2154,N_1959,N_1940);
nor U2155 (N_2155,N_1847,N_1866);
and U2156 (N_2156,N_1811,N_1802);
nor U2157 (N_2157,N_1996,N_1949);
and U2158 (N_2158,N_1993,N_1969);
and U2159 (N_2159,N_1942,N_1953);
and U2160 (N_2160,N_1862,N_1963);
and U2161 (N_2161,N_1934,N_1874);
or U2162 (N_2162,N_1814,N_1848);
and U2163 (N_2163,N_1934,N_1952);
nand U2164 (N_2164,N_1809,N_1900);
nor U2165 (N_2165,N_1819,N_1949);
nor U2166 (N_2166,N_1827,N_1868);
or U2167 (N_2167,N_1911,N_1865);
nor U2168 (N_2168,N_1990,N_1936);
nand U2169 (N_2169,N_1865,N_1944);
nor U2170 (N_2170,N_1931,N_1883);
and U2171 (N_2171,N_1971,N_1922);
nand U2172 (N_2172,N_1958,N_1815);
or U2173 (N_2173,N_1906,N_1809);
nand U2174 (N_2174,N_1908,N_1818);
nand U2175 (N_2175,N_1969,N_1914);
nand U2176 (N_2176,N_1969,N_1846);
nor U2177 (N_2177,N_1982,N_1860);
and U2178 (N_2178,N_1992,N_1816);
and U2179 (N_2179,N_1996,N_1908);
nor U2180 (N_2180,N_1869,N_1961);
and U2181 (N_2181,N_1845,N_1947);
nor U2182 (N_2182,N_1881,N_1973);
nand U2183 (N_2183,N_1908,N_1945);
and U2184 (N_2184,N_1963,N_1845);
xnor U2185 (N_2185,N_1877,N_1927);
nor U2186 (N_2186,N_1836,N_1870);
and U2187 (N_2187,N_1851,N_1806);
or U2188 (N_2188,N_1948,N_1980);
or U2189 (N_2189,N_1989,N_1923);
and U2190 (N_2190,N_1990,N_1835);
nand U2191 (N_2191,N_1912,N_1998);
nor U2192 (N_2192,N_1902,N_1889);
or U2193 (N_2193,N_1894,N_1832);
nand U2194 (N_2194,N_1949,N_1982);
or U2195 (N_2195,N_1884,N_1883);
or U2196 (N_2196,N_1884,N_1843);
nand U2197 (N_2197,N_1908,N_1956);
or U2198 (N_2198,N_1952,N_1887);
or U2199 (N_2199,N_1886,N_1968);
nor U2200 (N_2200,N_2010,N_2124);
nand U2201 (N_2201,N_2028,N_2067);
or U2202 (N_2202,N_2096,N_2163);
or U2203 (N_2203,N_2042,N_2035);
nand U2204 (N_2204,N_2036,N_2185);
and U2205 (N_2205,N_2105,N_2136);
nand U2206 (N_2206,N_2117,N_2143);
nand U2207 (N_2207,N_2012,N_2087);
and U2208 (N_2208,N_2044,N_2190);
nand U2209 (N_2209,N_2016,N_2169);
nor U2210 (N_2210,N_2155,N_2106);
nand U2211 (N_2211,N_2005,N_2186);
or U2212 (N_2212,N_2138,N_2085);
nand U2213 (N_2213,N_2064,N_2183);
and U2214 (N_2214,N_2058,N_2068);
nor U2215 (N_2215,N_2111,N_2008);
nor U2216 (N_2216,N_2041,N_2131);
nor U2217 (N_2217,N_2081,N_2188);
nand U2218 (N_2218,N_2056,N_2071);
nor U2219 (N_2219,N_2059,N_2025);
and U2220 (N_2220,N_2001,N_2161);
nor U2221 (N_2221,N_2133,N_2139);
and U2222 (N_2222,N_2156,N_2108);
nor U2223 (N_2223,N_2069,N_2130);
nand U2224 (N_2224,N_2088,N_2160);
nor U2225 (N_2225,N_2014,N_2029);
or U2226 (N_2226,N_2097,N_2094);
and U2227 (N_2227,N_2062,N_2026);
and U2228 (N_2228,N_2151,N_2004);
and U2229 (N_2229,N_2034,N_2015);
nor U2230 (N_2230,N_2137,N_2061);
nor U2231 (N_2231,N_2132,N_2189);
nor U2232 (N_2232,N_2089,N_2075);
or U2233 (N_2233,N_2002,N_2184);
nor U2234 (N_2234,N_2178,N_2120);
nor U2235 (N_2235,N_2127,N_2022);
and U2236 (N_2236,N_2141,N_2037);
and U2237 (N_2237,N_2073,N_2048);
and U2238 (N_2238,N_2070,N_2198);
or U2239 (N_2239,N_2128,N_2021);
or U2240 (N_2240,N_2135,N_2027);
nor U2241 (N_2241,N_2082,N_2159);
nand U2242 (N_2242,N_2045,N_2119);
and U2243 (N_2243,N_2121,N_2074);
nor U2244 (N_2244,N_2182,N_2177);
nor U2245 (N_2245,N_2174,N_2083);
and U2246 (N_2246,N_2145,N_2146);
and U2247 (N_2247,N_2144,N_2157);
or U2248 (N_2248,N_2172,N_2149);
nand U2249 (N_2249,N_2003,N_2154);
nor U2250 (N_2250,N_2153,N_2040);
or U2251 (N_2251,N_2107,N_2013);
or U2252 (N_2252,N_2115,N_2019);
and U2253 (N_2253,N_2162,N_2104);
nand U2254 (N_2254,N_2140,N_2171);
nand U2255 (N_2255,N_2020,N_2179);
and U2256 (N_2256,N_2122,N_2170);
and U2257 (N_2257,N_2055,N_2168);
and U2258 (N_2258,N_2091,N_2100);
or U2259 (N_2259,N_2147,N_2009);
and U2260 (N_2260,N_2125,N_2018);
nor U2261 (N_2261,N_2197,N_2116);
nor U2262 (N_2262,N_2193,N_2011);
and U2263 (N_2263,N_2113,N_2077);
nor U2264 (N_2264,N_2038,N_2114);
nand U2265 (N_2265,N_2043,N_2109);
and U2266 (N_2266,N_2057,N_2031);
or U2267 (N_2267,N_2092,N_2080);
nand U2268 (N_2268,N_2134,N_2191);
or U2269 (N_2269,N_2187,N_2007);
nor U2270 (N_2270,N_2194,N_2090);
nor U2271 (N_2271,N_2158,N_2192);
nand U2272 (N_2272,N_2053,N_2195);
or U2273 (N_2273,N_2099,N_2199);
nand U2274 (N_2274,N_2165,N_2150);
and U2275 (N_2275,N_2173,N_2102);
and U2276 (N_2276,N_2196,N_2054);
and U2277 (N_2277,N_2006,N_2129);
nand U2278 (N_2278,N_2101,N_2030);
or U2279 (N_2279,N_2166,N_2084);
or U2280 (N_2280,N_2032,N_2024);
or U2281 (N_2281,N_2050,N_2110);
or U2282 (N_2282,N_2098,N_2123);
nor U2283 (N_2283,N_2181,N_2052);
nor U2284 (N_2284,N_2142,N_2072);
or U2285 (N_2285,N_2126,N_2175);
and U2286 (N_2286,N_2086,N_2112);
nand U2287 (N_2287,N_2148,N_2103);
and U2288 (N_2288,N_2093,N_2000);
xor U2289 (N_2289,N_2047,N_2065);
nand U2290 (N_2290,N_2079,N_2046);
and U2291 (N_2291,N_2152,N_2078);
and U2292 (N_2292,N_2167,N_2076);
nand U2293 (N_2293,N_2063,N_2164);
or U2294 (N_2294,N_2176,N_2180);
nor U2295 (N_2295,N_2118,N_2033);
and U2296 (N_2296,N_2066,N_2095);
nor U2297 (N_2297,N_2049,N_2051);
nor U2298 (N_2298,N_2023,N_2060);
and U2299 (N_2299,N_2039,N_2017);
nand U2300 (N_2300,N_2163,N_2050);
nand U2301 (N_2301,N_2033,N_2195);
nor U2302 (N_2302,N_2010,N_2189);
nand U2303 (N_2303,N_2117,N_2150);
nor U2304 (N_2304,N_2115,N_2191);
nand U2305 (N_2305,N_2043,N_2101);
nand U2306 (N_2306,N_2054,N_2008);
nor U2307 (N_2307,N_2173,N_2037);
and U2308 (N_2308,N_2030,N_2009);
nor U2309 (N_2309,N_2064,N_2146);
and U2310 (N_2310,N_2108,N_2155);
nand U2311 (N_2311,N_2052,N_2165);
and U2312 (N_2312,N_2176,N_2040);
or U2313 (N_2313,N_2172,N_2111);
nor U2314 (N_2314,N_2079,N_2186);
nor U2315 (N_2315,N_2067,N_2039);
xor U2316 (N_2316,N_2073,N_2097);
and U2317 (N_2317,N_2023,N_2030);
and U2318 (N_2318,N_2142,N_2148);
nor U2319 (N_2319,N_2082,N_2180);
and U2320 (N_2320,N_2067,N_2145);
xor U2321 (N_2321,N_2120,N_2191);
and U2322 (N_2322,N_2162,N_2068);
nor U2323 (N_2323,N_2161,N_2027);
or U2324 (N_2324,N_2132,N_2078);
nand U2325 (N_2325,N_2065,N_2136);
nand U2326 (N_2326,N_2082,N_2124);
or U2327 (N_2327,N_2046,N_2124);
and U2328 (N_2328,N_2169,N_2189);
nand U2329 (N_2329,N_2123,N_2024);
and U2330 (N_2330,N_2144,N_2013);
or U2331 (N_2331,N_2166,N_2113);
nor U2332 (N_2332,N_2153,N_2099);
nand U2333 (N_2333,N_2080,N_2165);
nor U2334 (N_2334,N_2060,N_2142);
nor U2335 (N_2335,N_2190,N_2196);
and U2336 (N_2336,N_2139,N_2116);
or U2337 (N_2337,N_2097,N_2177);
and U2338 (N_2338,N_2018,N_2094);
and U2339 (N_2339,N_2035,N_2066);
nand U2340 (N_2340,N_2017,N_2048);
and U2341 (N_2341,N_2177,N_2082);
nand U2342 (N_2342,N_2158,N_2149);
or U2343 (N_2343,N_2126,N_2038);
nand U2344 (N_2344,N_2011,N_2120);
or U2345 (N_2345,N_2172,N_2117);
nor U2346 (N_2346,N_2171,N_2136);
nor U2347 (N_2347,N_2166,N_2036);
nand U2348 (N_2348,N_2093,N_2140);
or U2349 (N_2349,N_2058,N_2168);
nand U2350 (N_2350,N_2009,N_2192);
nor U2351 (N_2351,N_2195,N_2158);
or U2352 (N_2352,N_2159,N_2076);
nor U2353 (N_2353,N_2135,N_2151);
nor U2354 (N_2354,N_2061,N_2005);
or U2355 (N_2355,N_2004,N_2197);
nand U2356 (N_2356,N_2152,N_2067);
nor U2357 (N_2357,N_2114,N_2056);
nor U2358 (N_2358,N_2048,N_2096);
and U2359 (N_2359,N_2155,N_2172);
nor U2360 (N_2360,N_2042,N_2091);
nand U2361 (N_2361,N_2059,N_2082);
nor U2362 (N_2362,N_2006,N_2002);
and U2363 (N_2363,N_2125,N_2110);
nor U2364 (N_2364,N_2004,N_2052);
or U2365 (N_2365,N_2009,N_2089);
nor U2366 (N_2366,N_2129,N_2157);
or U2367 (N_2367,N_2191,N_2158);
and U2368 (N_2368,N_2191,N_2140);
nand U2369 (N_2369,N_2081,N_2135);
nand U2370 (N_2370,N_2021,N_2172);
and U2371 (N_2371,N_2063,N_2089);
nand U2372 (N_2372,N_2130,N_2141);
or U2373 (N_2373,N_2006,N_2015);
nand U2374 (N_2374,N_2128,N_2154);
nand U2375 (N_2375,N_2176,N_2120);
xor U2376 (N_2376,N_2045,N_2051);
and U2377 (N_2377,N_2147,N_2083);
nor U2378 (N_2378,N_2057,N_2093);
or U2379 (N_2379,N_2106,N_2101);
nand U2380 (N_2380,N_2198,N_2193);
nor U2381 (N_2381,N_2182,N_2058);
nand U2382 (N_2382,N_2050,N_2048);
and U2383 (N_2383,N_2011,N_2002);
nand U2384 (N_2384,N_2046,N_2075);
xnor U2385 (N_2385,N_2180,N_2117);
xnor U2386 (N_2386,N_2025,N_2055);
or U2387 (N_2387,N_2143,N_2119);
nand U2388 (N_2388,N_2062,N_2194);
or U2389 (N_2389,N_2111,N_2126);
and U2390 (N_2390,N_2175,N_2078);
or U2391 (N_2391,N_2092,N_2172);
nor U2392 (N_2392,N_2061,N_2067);
nand U2393 (N_2393,N_2078,N_2147);
and U2394 (N_2394,N_2143,N_2061);
and U2395 (N_2395,N_2010,N_2097);
nor U2396 (N_2396,N_2045,N_2111);
and U2397 (N_2397,N_2084,N_2126);
nand U2398 (N_2398,N_2001,N_2158);
and U2399 (N_2399,N_2141,N_2142);
nand U2400 (N_2400,N_2348,N_2387);
nor U2401 (N_2401,N_2314,N_2212);
nand U2402 (N_2402,N_2217,N_2274);
nand U2403 (N_2403,N_2395,N_2245);
and U2404 (N_2404,N_2200,N_2390);
nor U2405 (N_2405,N_2377,N_2281);
nor U2406 (N_2406,N_2209,N_2346);
and U2407 (N_2407,N_2389,N_2256);
or U2408 (N_2408,N_2367,N_2218);
or U2409 (N_2409,N_2250,N_2296);
nor U2410 (N_2410,N_2297,N_2391);
and U2411 (N_2411,N_2290,N_2321);
nand U2412 (N_2412,N_2319,N_2360);
nor U2413 (N_2413,N_2313,N_2222);
and U2414 (N_2414,N_2324,N_2268);
nor U2415 (N_2415,N_2304,N_2328);
nor U2416 (N_2416,N_2275,N_2345);
or U2417 (N_2417,N_2271,N_2237);
nand U2418 (N_2418,N_2272,N_2287);
and U2419 (N_2419,N_2386,N_2259);
nand U2420 (N_2420,N_2246,N_2206);
or U2421 (N_2421,N_2234,N_2322);
and U2422 (N_2422,N_2388,N_2249);
nand U2423 (N_2423,N_2341,N_2219);
nor U2424 (N_2424,N_2374,N_2393);
or U2425 (N_2425,N_2226,N_2251);
or U2426 (N_2426,N_2302,N_2361);
or U2427 (N_2427,N_2370,N_2210);
or U2428 (N_2428,N_2349,N_2383);
nor U2429 (N_2429,N_2356,N_2265);
xor U2430 (N_2430,N_2330,N_2225);
and U2431 (N_2431,N_2359,N_2352);
and U2432 (N_2432,N_2310,N_2207);
nor U2433 (N_2433,N_2267,N_2295);
or U2434 (N_2434,N_2230,N_2331);
or U2435 (N_2435,N_2224,N_2340);
nand U2436 (N_2436,N_2255,N_2334);
and U2437 (N_2437,N_2220,N_2381);
and U2438 (N_2438,N_2286,N_2253);
and U2439 (N_2439,N_2247,N_2293);
and U2440 (N_2440,N_2364,N_2369);
or U2441 (N_2441,N_2357,N_2235);
or U2442 (N_2442,N_2298,N_2337);
or U2443 (N_2443,N_2240,N_2291);
or U2444 (N_2444,N_2236,N_2283);
nand U2445 (N_2445,N_2316,N_2371);
and U2446 (N_2446,N_2327,N_2320);
or U2447 (N_2447,N_2312,N_2354);
nand U2448 (N_2448,N_2284,N_2227);
or U2449 (N_2449,N_2292,N_2289);
nand U2450 (N_2450,N_2299,N_2335);
or U2451 (N_2451,N_2373,N_2343);
nor U2452 (N_2452,N_2303,N_2338);
nor U2453 (N_2453,N_2294,N_2211);
nand U2454 (N_2454,N_2363,N_2308);
and U2455 (N_2455,N_2232,N_2325);
and U2456 (N_2456,N_2201,N_2311);
nor U2457 (N_2457,N_2257,N_2254);
or U2458 (N_2458,N_2384,N_2396);
and U2459 (N_2459,N_2355,N_2215);
nor U2460 (N_2460,N_2288,N_2329);
or U2461 (N_2461,N_2379,N_2205);
or U2462 (N_2462,N_2203,N_2368);
nand U2463 (N_2463,N_2277,N_2305);
or U2464 (N_2464,N_2266,N_2344);
and U2465 (N_2465,N_2399,N_2204);
nor U2466 (N_2466,N_2242,N_2276);
and U2467 (N_2467,N_2333,N_2243);
or U2468 (N_2468,N_2248,N_2262);
nor U2469 (N_2469,N_2397,N_2336);
nor U2470 (N_2470,N_2280,N_2339);
or U2471 (N_2471,N_2260,N_2350);
nand U2472 (N_2472,N_2332,N_2382);
nand U2473 (N_2473,N_2375,N_2231);
or U2474 (N_2474,N_2353,N_2239);
and U2475 (N_2475,N_2326,N_2365);
nor U2476 (N_2476,N_2282,N_2398);
and U2477 (N_2477,N_2306,N_2323);
and U2478 (N_2478,N_2244,N_2221);
nor U2479 (N_2479,N_2229,N_2238);
and U2480 (N_2480,N_2362,N_2223);
or U2481 (N_2481,N_2264,N_2216);
nor U2482 (N_2482,N_2285,N_2351);
nand U2483 (N_2483,N_2278,N_2261);
and U2484 (N_2484,N_2233,N_2315);
and U2485 (N_2485,N_2347,N_2258);
nand U2486 (N_2486,N_2366,N_2273);
xor U2487 (N_2487,N_2269,N_2358);
or U2488 (N_2488,N_2252,N_2309);
or U2489 (N_2489,N_2241,N_2380);
xor U2490 (N_2490,N_2202,N_2307);
or U2491 (N_2491,N_2317,N_2279);
nand U2492 (N_2492,N_2342,N_2214);
and U2493 (N_2493,N_2301,N_2228);
or U2494 (N_2494,N_2372,N_2213);
or U2495 (N_2495,N_2378,N_2270);
or U2496 (N_2496,N_2318,N_2394);
or U2497 (N_2497,N_2376,N_2300);
nand U2498 (N_2498,N_2263,N_2208);
nor U2499 (N_2499,N_2392,N_2385);
nor U2500 (N_2500,N_2321,N_2314);
nor U2501 (N_2501,N_2329,N_2212);
nor U2502 (N_2502,N_2333,N_2350);
or U2503 (N_2503,N_2211,N_2369);
xnor U2504 (N_2504,N_2222,N_2339);
nand U2505 (N_2505,N_2396,N_2264);
and U2506 (N_2506,N_2274,N_2279);
nand U2507 (N_2507,N_2291,N_2200);
and U2508 (N_2508,N_2354,N_2336);
nand U2509 (N_2509,N_2328,N_2231);
and U2510 (N_2510,N_2388,N_2378);
xnor U2511 (N_2511,N_2363,N_2254);
nor U2512 (N_2512,N_2320,N_2330);
or U2513 (N_2513,N_2276,N_2212);
or U2514 (N_2514,N_2342,N_2205);
nor U2515 (N_2515,N_2388,N_2327);
or U2516 (N_2516,N_2218,N_2266);
nand U2517 (N_2517,N_2383,N_2225);
nand U2518 (N_2518,N_2311,N_2380);
and U2519 (N_2519,N_2309,N_2229);
nor U2520 (N_2520,N_2212,N_2241);
or U2521 (N_2521,N_2333,N_2330);
nor U2522 (N_2522,N_2232,N_2286);
xor U2523 (N_2523,N_2354,N_2200);
nor U2524 (N_2524,N_2341,N_2201);
nor U2525 (N_2525,N_2298,N_2313);
nor U2526 (N_2526,N_2238,N_2372);
or U2527 (N_2527,N_2373,N_2234);
or U2528 (N_2528,N_2386,N_2232);
nand U2529 (N_2529,N_2235,N_2358);
nand U2530 (N_2530,N_2226,N_2270);
nor U2531 (N_2531,N_2224,N_2330);
nand U2532 (N_2532,N_2275,N_2272);
and U2533 (N_2533,N_2362,N_2309);
or U2534 (N_2534,N_2326,N_2274);
or U2535 (N_2535,N_2383,N_2384);
or U2536 (N_2536,N_2340,N_2310);
and U2537 (N_2537,N_2216,N_2225);
nand U2538 (N_2538,N_2323,N_2280);
and U2539 (N_2539,N_2242,N_2214);
nor U2540 (N_2540,N_2311,N_2253);
or U2541 (N_2541,N_2379,N_2385);
or U2542 (N_2542,N_2343,N_2292);
and U2543 (N_2543,N_2235,N_2234);
or U2544 (N_2544,N_2225,N_2375);
or U2545 (N_2545,N_2262,N_2237);
and U2546 (N_2546,N_2262,N_2209);
or U2547 (N_2547,N_2310,N_2261);
nor U2548 (N_2548,N_2219,N_2359);
and U2549 (N_2549,N_2235,N_2226);
nor U2550 (N_2550,N_2349,N_2299);
nor U2551 (N_2551,N_2297,N_2347);
nand U2552 (N_2552,N_2344,N_2338);
or U2553 (N_2553,N_2238,N_2227);
or U2554 (N_2554,N_2381,N_2236);
nor U2555 (N_2555,N_2229,N_2215);
and U2556 (N_2556,N_2388,N_2237);
nand U2557 (N_2557,N_2324,N_2387);
nor U2558 (N_2558,N_2389,N_2219);
or U2559 (N_2559,N_2294,N_2370);
nand U2560 (N_2560,N_2383,N_2355);
nor U2561 (N_2561,N_2299,N_2248);
or U2562 (N_2562,N_2265,N_2226);
nand U2563 (N_2563,N_2391,N_2313);
nor U2564 (N_2564,N_2282,N_2397);
nand U2565 (N_2565,N_2336,N_2203);
nor U2566 (N_2566,N_2246,N_2391);
or U2567 (N_2567,N_2238,N_2384);
or U2568 (N_2568,N_2302,N_2286);
or U2569 (N_2569,N_2327,N_2286);
nor U2570 (N_2570,N_2244,N_2342);
nand U2571 (N_2571,N_2371,N_2395);
nor U2572 (N_2572,N_2203,N_2343);
nor U2573 (N_2573,N_2360,N_2269);
or U2574 (N_2574,N_2213,N_2227);
nand U2575 (N_2575,N_2254,N_2264);
and U2576 (N_2576,N_2308,N_2372);
and U2577 (N_2577,N_2386,N_2392);
nand U2578 (N_2578,N_2369,N_2216);
xnor U2579 (N_2579,N_2372,N_2346);
nor U2580 (N_2580,N_2211,N_2396);
nor U2581 (N_2581,N_2253,N_2352);
nand U2582 (N_2582,N_2333,N_2378);
and U2583 (N_2583,N_2224,N_2287);
nor U2584 (N_2584,N_2277,N_2240);
nor U2585 (N_2585,N_2367,N_2360);
and U2586 (N_2586,N_2293,N_2225);
nor U2587 (N_2587,N_2306,N_2267);
nor U2588 (N_2588,N_2351,N_2241);
and U2589 (N_2589,N_2366,N_2236);
or U2590 (N_2590,N_2260,N_2283);
and U2591 (N_2591,N_2258,N_2290);
nand U2592 (N_2592,N_2320,N_2257);
nor U2593 (N_2593,N_2386,N_2339);
nand U2594 (N_2594,N_2373,N_2341);
and U2595 (N_2595,N_2360,N_2310);
nand U2596 (N_2596,N_2203,N_2350);
nor U2597 (N_2597,N_2217,N_2351);
or U2598 (N_2598,N_2281,N_2269);
and U2599 (N_2599,N_2312,N_2390);
nor U2600 (N_2600,N_2538,N_2468);
nor U2601 (N_2601,N_2555,N_2473);
and U2602 (N_2602,N_2417,N_2478);
nand U2603 (N_2603,N_2431,N_2501);
or U2604 (N_2604,N_2598,N_2491);
or U2605 (N_2605,N_2400,N_2449);
nand U2606 (N_2606,N_2488,N_2452);
or U2607 (N_2607,N_2521,N_2525);
nand U2608 (N_2608,N_2524,N_2539);
or U2609 (N_2609,N_2585,N_2593);
or U2610 (N_2610,N_2564,N_2535);
or U2611 (N_2611,N_2416,N_2408);
and U2612 (N_2612,N_2546,N_2595);
or U2613 (N_2613,N_2407,N_2497);
and U2614 (N_2614,N_2415,N_2437);
or U2615 (N_2615,N_2581,N_2550);
nor U2616 (N_2616,N_2561,N_2493);
or U2617 (N_2617,N_2511,N_2515);
or U2618 (N_2618,N_2577,N_2574);
or U2619 (N_2619,N_2494,N_2553);
nand U2620 (N_2620,N_2476,N_2448);
nand U2621 (N_2621,N_2500,N_2441);
nand U2622 (N_2622,N_2444,N_2519);
nand U2623 (N_2623,N_2460,N_2483);
xnor U2624 (N_2624,N_2498,N_2482);
nand U2625 (N_2625,N_2462,N_2549);
or U2626 (N_2626,N_2461,N_2474);
or U2627 (N_2627,N_2590,N_2544);
nand U2628 (N_2628,N_2418,N_2499);
and U2629 (N_2629,N_2438,N_2570);
and U2630 (N_2630,N_2432,N_2430);
or U2631 (N_2631,N_2424,N_2455);
and U2632 (N_2632,N_2413,N_2496);
nand U2633 (N_2633,N_2443,N_2588);
or U2634 (N_2634,N_2536,N_2467);
or U2635 (N_2635,N_2412,N_2560);
nor U2636 (N_2636,N_2596,N_2409);
and U2637 (N_2637,N_2517,N_2470);
nor U2638 (N_2638,N_2589,N_2547);
and U2639 (N_2639,N_2558,N_2484);
nand U2640 (N_2640,N_2422,N_2587);
or U2641 (N_2641,N_2583,N_2486);
nor U2642 (N_2642,N_2551,N_2453);
nor U2643 (N_2643,N_2402,N_2423);
nand U2644 (N_2644,N_2428,N_2512);
nor U2645 (N_2645,N_2427,N_2472);
xnor U2646 (N_2646,N_2404,N_2563);
nor U2647 (N_2647,N_2419,N_2533);
nand U2648 (N_2648,N_2505,N_2548);
and U2649 (N_2649,N_2485,N_2456);
nand U2650 (N_2650,N_2411,N_2506);
or U2651 (N_2651,N_2523,N_2507);
and U2652 (N_2652,N_2557,N_2463);
nand U2653 (N_2653,N_2526,N_2454);
xor U2654 (N_2654,N_2464,N_2573);
nand U2655 (N_2655,N_2459,N_2514);
and U2656 (N_2656,N_2599,N_2410);
nor U2657 (N_2657,N_2425,N_2554);
and U2658 (N_2658,N_2552,N_2445);
and U2659 (N_2659,N_2540,N_2545);
and U2660 (N_2660,N_2591,N_2481);
nand U2661 (N_2661,N_2578,N_2421);
or U2662 (N_2662,N_2527,N_2580);
nand U2663 (N_2663,N_2489,N_2576);
or U2664 (N_2664,N_2513,N_2508);
and U2665 (N_2665,N_2490,N_2528);
and U2666 (N_2666,N_2439,N_2531);
nand U2667 (N_2667,N_2442,N_2565);
nand U2668 (N_2668,N_2433,N_2492);
and U2669 (N_2669,N_2469,N_2566);
nor U2670 (N_2670,N_2503,N_2405);
nand U2671 (N_2671,N_2542,N_2575);
nor U2672 (N_2672,N_2529,N_2434);
nor U2673 (N_2673,N_2495,N_2569);
nand U2674 (N_2674,N_2436,N_2592);
and U2675 (N_2675,N_2440,N_2582);
and U2676 (N_2676,N_2471,N_2522);
nor U2677 (N_2677,N_2567,N_2556);
and U2678 (N_2678,N_2584,N_2504);
nor U2679 (N_2679,N_2518,N_2520);
and U2680 (N_2680,N_2457,N_2414);
or U2681 (N_2681,N_2516,N_2426);
nor U2682 (N_2682,N_2530,N_2502);
nand U2683 (N_2683,N_2532,N_2466);
and U2684 (N_2684,N_2479,N_2435);
nor U2685 (N_2685,N_2403,N_2446);
or U2686 (N_2686,N_2420,N_2543);
and U2687 (N_2687,N_2537,N_2579);
or U2688 (N_2688,N_2541,N_2465);
nand U2689 (N_2689,N_2458,N_2487);
or U2690 (N_2690,N_2571,N_2475);
or U2691 (N_2691,N_2572,N_2429);
nor U2692 (N_2692,N_2510,N_2568);
nand U2693 (N_2693,N_2562,N_2586);
and U2694 (N_2694,N_2447,N_2534);
or U2695 (N_2695,N_2477,N_2451);
or U2696 (N_2696,N_2597,N_2559);
nand U2697 (N_2697,N_2401,N_2509);
and U2698 (N_2698,N_2450,N_2406);
or U2699 (N_2699,N_2480,N_2594);
or U2700 (N_2700,N_2422,N_2416);
xnor U2701 (N_2701,N_2442,N_2492);
or U2702 (N_2702,N_2517,N_2536);
nand U2703 (N_2703,N_2518,N_2403);
or U2704 (N_2704,N_2466,N_2401);
nand U2705 (N_2705,N_2494,N_2598);
and U2706 (N_2706,N_2568,N_2548);
or U2707 (N_2707,N_2475,N_2579);
and U2708 (N_2708,N_2489,N_2410);
or U2709 (N_2709,N_2476,N_2520);
nand U2710 (N_2710,N_2495,N_2584);
nand U2711 (N_2711,N_2520,N_2456);
or U2712 (N_2712,N_2513,N_2583);
xnor U2713 (N_2713,N_2427,N_2591);
nor U2714 (N_2714,N_2400,N_2467);
and U2715 (N_2715,N_2415,N_2427);
and U2716 (N_2716,N_2433,N_2580);
or U2717 (N_2717,N_2569,N_2424);
or U2718 (N_2718,N_2540,N_2486);
xnor U2719 (N_2719,N_2461,N_2505);
nand U2720 (N_2720,N_2593,N_2589);
nand U2721 (N_2721,N_2577,N_2417);
and U2722 (N_2722,N_2589,N_2417);
nor U2723 (N_2723,N_2417,N_2511);
nor U2724 (N_2724,N_2441,N_2474);
nor U2725 (N_2725,N_2448,N_2417);
or U2726 (N_2726,N_2506,N_2530);
nand U2727 (N_2727,N_2583,N_2476);
nor U2728 (N_2728,N_2410,N_2563);
or U2729 (N_2729,N_2472,N_2596);
and U2730 (N_2730,N_2440,N_2580);
nand U2731 (N_2731,N_2490,N_2437);
nor U2732 (N_2732,N_2432,N_2591);
or U2733 (N_2733,N_2431,N_2570);
nand U2734 (N_2734,N_2439,N_2561);
nand U2735 (N_2735,N_2502,N_2544);
or U2736 (N_2736,N_2546,N_2463);
nor U2737 (N_2737,N_2525,N_2430);
nor U2738 (N_2738,N_2560,N_2410);
nand U2739 (N_2739,N_2457,N_2532);
nor U2740 (N_2740,N_2533,N_2460);
nor U2741 (N_2741,N_2582,N_2444);
and U2742 (N_2742,N_2571,N_2427);
and U2743 (N_2743,N_2576,N_2548);
nand U2744 (N_2744,N_2412,N_2481);
nand U2745 (N_2745,N_2559,N_2437);
and U2746 (N_2746,N_2476,N_2409);
nand U2747 (N_2747,N_2591,N_2560);
and U2748 (N_2748,N_2573,N_2400);
nand U2749 (N_2749,N_2545,N_2519);
and U2750 (N_2750,N_2554,N_2535);
nand U2751 (N_2751,N_2581,N_2545);
nand U2752 (N_2752,N_2584,N_2570);
nor U2753 (N_2753,N_2562,N_2469);
or U2754 (N_2754,N_2502,N_2523);
nand U2755 (N_2755,N_2486,N_2541);
nor U2756 (N_2756,N_2487,N_2478);
xor U2757 (N_2757,N_2553,N_2534);
nand U2758 (N_2758,N_2505,N_2430);
and U2759 (N_2759,N_2409,N_2491);
nor U2760 (N_2760,N_2539,N_2513);
nor U2761 (N_2761,N_2549,N_2525);
or U2762 (N_2762,N_2429,N_2405);
nand U2763 (N_2763,N_2583,N_2515);
nand U2764 (N_2764,N_2484,N_2431);
and U2765 (N_2765,N_2549,N_2424);
nor U2766 (N_2766,N_2464,N_2564);
nand U2767 (N_2767,N_2498,N_2461);
nor U2768 (N_2768,N_2482,N_2550);
or U2769 (N_2769,N_2403,N_2428);
nand U2770 (N_2770,N_2431,N_2548);
nor U2771 (N_2771,N_2473,N_2593);
nor U2772 (N_2772,N_2476,N_2584);
nor U2773 (N_2773,N_2414,N_2578);
nand U2774 (N_2774,N_2571,N_2445);
nand U2775 (N_2775,N_2479,N_2545);
nor U2776 (N_2776,N_2509,N_2564);
and U2777 (N_2777,N_2579,N_2577);
nor U2778 (N_2778,N_2557,N_2403);
and U2779 (N_2779,N_2412,N_2450);
xnor U2780 (N_2780,N_2462,N_2457);
nor U2781 (N_2781,N_2536,N_2530);
or U2782 (N_2782,N_2576,N_2499);
nor U2783 (N_2783,N_2437,N_2549);
or U2784 (N_2784,N_2491,N_2545);
nand U2785 (N_2785,N_2404,N_2431);
or U2786 (N_2786,N_2513,N_2466);
nand U2787 (N_2787,N_2474,N_2464);
and U2788 (N_2788,N_2568,N_2416);
nand U2789 (N_2789,N_2468,N_2471);
nor U2790 (N_2790,N_2551,N_2512);
nor U2791 (N_2791,N_2599,N_2439);
nor U2792 (N_2792,N_2450,N_2596);
and U2793 (N_2793,N_2431,N_2464);
nand U2794 (N_2794,N_2473,N_2496);
and U2795 (N_2795,N_2410,N_2406);
nor U2796 (N_2796,N_2568,N_2533);
nor U2797 (N_2797,N_2496,N_2569);
nand U2798 (N_2798,N_2536,N_2423);
nand U2799 (N_2799,N_2451,N_2555);
or U2800 (N_2800,N_2695,N_2669);
xor U2801 (N_2801,N_2626,N_2710);
nand U2802 (N_2802,N_2684,N_2744);
and U2803 (N_2803,N_2656,N_2799);
nand U2804 (N_2804,N_2784,N_2625);
nand U2805 (N_2805,N_2700,N_2611);
and U2806 (N_2806,N_2725,N_2740);
and U2807 (N_2807,N_2792,N_2655);
or U2808 (N_2808,N_2603,N_2765);
nor U2809 (N_2809,N_2658,N_2750);
nor U2810 (N_2810,N_2670,N_2758);
nand U2811 (N_2811,N_2693,N_2754);
or U2812 (N_2812,N_2604,N_2650);
nand U2813 (N_2813,N_2640,N_2652);
or U2814 (N_2814,N_2606,N_2668);
nor U2815 (N_2815,N_2764,N_2600);
nor U2816 (N_2816,N_2634,N_2676);
nor U2817 (N_2817,N_2622,N_2616);
nor U2818 (N_2818,N_2649,N_2718);
and U2819 (N_2819,N_2760,N_2618);
or U2820 (N_2820,N_2797,N_2749);
or U2821 (N_2821,N_2722,N_2644);
or U2822 (N_2822,N_2686,N_2787);
and U2823 (N_2823,N_2778,N_2709);
or U2824 (N_2824,N_2673,N_2752);
nand U2825 (N_2825,N_2796,N_2780);
or U2826 (N_2826,N_2687,N_2653);
nor U2827 (N_2827,N_2646,N_2748);
and U2828 (N_2828,N_2729,N_2761);
nand U2829 (N_2829,N_2737,N_2636);
and U2830 (N_2830,N_2753,N_2769);
or U2831 (N_2831,N_2621,N_2741);
nor U2832 (N_2832,N_2619,N_2654);
nor U2833 (N_2833,N_2648,N_2763);
and U2834 (N_2834,N_2691,N_2708);
nand U2835 (N_2835,N_2713,N_2759);
nor U2836 (N_2836,N_2746,N_2671);
or U2837 (N_2837,N_2793,N_2743);
nand U2838 (N_2838,N_2630,N_2633);
and U2839 (N_2839,N_2627,N_2624);
and U2840 (N_2840,N_2608,N_2731);
and U2841 (N_2841,N_2772,N_2637);
nand U2842 (N_2842,N_2711,N_2775);
nand U2843 (N_2843,N_2755,N_2661);
nor U2844 (N_2844,N_2790,N_2664);
nand U2845 (N_2845,N_2738,N_2766);
and U2846 (N_2846,N_2703,N_2771);
or U2847 (N_2847,N_2666,N_2774);
and U2848 (N_2848,N_2727,N_2660);
or U2849 (N_2849,N_2675,N_2694);
nor U2850 (N_2850,N_2629,N_2742);
nand U2851 (N_2851,N_2662,N_2614);
or U2852 (N_2852,N_2623,N_2798);
nand U2853 (N_2853,N_2732,N_2723);
and U2854 (N_2854,N_2719,N_2701);
or U2855 (N_2855,N_2714,N_2781);
and U2856 (N_2856,N_2638,N_2699);
xor U2857 (N_2857,N_2751,N_2779);
or U2858 (N_2858,N_2706,N_2683);
and U2859 (N_2859,N_2663,N_2692);
or U2860 (N_2860,N_2685,N_2734);
nand U2861 (N_2861,N_2651,N_2688);
and U2862 (N_2862,N_2647,N_2788);
xnor U2863 (N_2863,N_2712,N_2715);
and U2864 (N_2864,N_2770,N_2605);
or U2865 (N_2865,N_2674,N_2667);
or U2866 (N_2866,N_2717,N_2786);
nor U2867 (N_2867,N_2782,N_2678);
nor U2868 (N_2868,N_2601,N_2602);
nand U2869 (N_2869,N_2726,N_2659);
nor U2870 (N_2870,N_2607,N_2696);
and U2871 (N_2871,N_2768,N_2720);
nand U2872 (N_2872,N_2767,N_2756);
nand U2873 (N_2873,N_2609,N_2641);
and U2874 (N_2874,N_2739,N_2735);
and U2875 (N_2875,N_2724,N_2690);
or U2876 (N_2876,N_2707,N_2615);
or U2877 (N_2877,N_2762,N_2612);
or U2878 (N_2878,N_2665,N_2777);
nand U2879 (N_2879,N_2736,N_2791);
and U2880 (N_2880,N_2733,N_2721);
nand U2881 (N_2881,N_2642,N_2645);
and U2882 (N_2882,N_2698,N_2704);
nor U2883 (N_2883,N_2620,N_2794);
nor U2884 (N_2884,N_2672,N_2702);
and U2885 (N_2885,N_2639,N_2635);
nor U2886 (N_2886,N_2682,N_2697);
nor U2887 (N_2887,N_2705,N_2632);
nand U2888 (N_2888,N_2783,N_2680);
nor U2889 (N_2889,N_2610,N_2716);
nand U2890 (N_2890,N_2613,N_2745);
nand U2891 (N_2891,N_2776,N_2643);
nor U2892 (N_2892,N_2795,N_2679);
nand U2893 (N_2893,N_2617,N_2728);
nand U2894 (N_2894,N_2631,N_2747);
or U2895 (N_2895,N_2757,N_2628);
nand U2896 (N_2896,N_2657,N_2681);
nor U2897 (N_2897,N_2789,N_2773);
nand U2898 (N_2898,N_2677,N_2785);
nand U2899 (N_2899,N_2689,N_2730);
nand U2900 (N_2900,N_2781,N_2743);
xor U2901 (N_2901,N_2683,N_2635);
or U2902 (N_2902,N_2709,N_2771);
or U2903 (N_2903,N_2670,N_2778);
or U2904 (N_2904,N_2770,N_2725);
nand U2905 (N_2905,N_2740,N_2755);
nor U2906 (N_2906,N_2697,N_2614);
and U2907 (N_2907,N_2778,N_2704);
nand U2908 (N_2908,N_2783,N_2790);
and U2909 (N_2909,N_2720,N_2647);
xnor U2910 (N_2910,N_2757,N_2639);
or U2911 (N_2911,N_2707,N_2733);
nand U2912 (N_2912,N_2718,N_2706);
or U2913 (N_2913,N_2733,N_2694);
nor U2914 (N_2914,N_2787,N_2684);
nand U2915 (N_2915,N_2629,N_2657);
and U2916 (N_2916,N_2758,N_2660);
nor U2917 (N_2917,N_2683,N_2771);
or U2918 (N_2918,N_2708,N_2781);
nand U2919 (N_2919,N_2638,N_2659);
xnor U2920 (N_2920,N_2612,N_2679);
nor U2921 (N_2921,N_2763,N_2661);
nand U2922 (N_2922,N_2709,N_2624);
and U2923 (N_2923,N_2678,N_2739);
nand U2924 (N_2924,N_2621,N_2786);
xor U2925 (N_2925,N_2767,N_2663);
nand U2926 (N_2926,N_2732,N_2784);
nor U2927 (N_2927,N_2792,N_2790);
nand U2928 (N_2928,N_2621,N_2704);
nor U2929 (N_2929,N_2755,N_2610);
and U2930 (N_2930,N_2767,N_2672);
nand U2931 (N_2931,N_2738,N_2653);
nor U2932 (N_2932,N_2680,N_2723);
nor U2933 (N_2933,N_2702,N_2624);
xnor U2934 (N_2934,N_2747,N_2625);
nand U2935 (N_2935,N_2647,N_2690);
nand U2936 (N_2936,N_2670,N_2642);
or U2937 (N_2937,N_2645,N_2615);
or U2938 (N_2938,N_2623,N_2747);
or U2939 (N_2939,N_2770,N_2635);
and U2940 (N_2940,N_2745,N_2701);
or U2941 (N_2941,N_2601,N_2622);
and U2942 (N_2942,N_2727,N_2674);
nand U2943 (N_2943,N_2714,N_2645);
or U2944 (N_2944,N_2780,N_2608);
nor U2945 (N_2945,N_2604,N_2638);
nand U2946 (N_2946,N_2680,N_2767);
nor U2947 (N_2947,N_2637,N_2739);
nor U2948 (N_2948,N_2619,N_2635);
and U2949 (N_2949,N_2632,N_2637);
or U2950 (N_2950,N_2761,N_2754);
nor U2951 (N_2951,N_2635,N_2733);
nand U2952 (N_2952,N_2776,N_2641);
or U2953 (N_2953,N_2630,N_2703);
and U2954 (N_2954,N_2672,N_2613);
or U2955 (N_2955,N_2738,N_2787);
nor U2956 (N_2956,N_2754,N_2753);
or U2957 (N_2957,N_2652,N_2737);
nand U2958 (N_2958,N_2764,N_2705);
and U2959 (N_2959,N_2673,N_2614);
nand U2960 (N_2960,N_2680,N_2657);
nand U2961 (N_2961,N_2605,N_2637);
or U2962 (N_2962,N_2698,N_2694);
or U2963 (N_2963,N_2653,N_2633);
or U2964 (N_2964,N_2608,N_2728);
and U2965 (N_2965,N_2706,N_2636);
or U2966 (N_2966,N_2643,N_2769);
nand U2967 (N_2967,N_2674,N_2751);
or U2968 (N_2968,N_2673,N_2774);
nor U2969 (N_2969,N_2659,N_2784);
nand U2970 (N_2970,N_2742,N_2777);
nand U2971 (N_2971,N_2745,N_2712);
or U2972 (N_2972,N_2690,N_2689);
nand U2973 (N_2973,N_2726,N_2653);
nand U2974 (N_2974,N_2686,N_2665);
nand U2975 (N_2975,N_2715,N_2772);
or U2976 (N_2976,N_2707,N_2620);
or U2977 (N_2977,N_2684,N_2649);
nand U2978 (N_2978,N_2705,N_2700);
nand U2979 (N_2979,N_2775,N_2746);
nor U2980 (N_2980,N_2678,N_2767);
or U2981 (N_2981,N_2699,N_2786);
nand U2982 (N_2982,N_2660,N_2601);
nand U2983 (N_2983,N_2732,N_2686);
and U2984 (N_2984,N_2758,N_2763);
xnor U2985 (N_2985,N_2622,N_2735);
or U2986 (N_2986,N_2704,N_2650);
nand U2987 (N_2987,N_2717,N_2623);
nor U2988 (N_2988,N_2731,N_2697);
or U2989 (N_2989,N_2639,N_2791);
or U2990 (N_2990,N_2636,N_2640);
or U2991 (N_2991,N_2744,N_2769);
or U2992 (N_2992,N_2639,N_2724);
nor U2993 (N_2993,N_2615,N_2619);
nor U2994 (N_2994,N_2785,N_2618);
and U2995 (N_2995,N_2669,N_2698);
nor U2996 (N_2996,N_2780,N_2629);
nand U2997 (N_2997,N_2615,N_2767);
nand U2998 (N_2998,N_2653,N_2700);
and U2999 (N_2999,N_2753,N_2686);
nor UO_0 (O_0,N_2969,N_2990);
nand UO_1 (O_1,N_2885,N_2810);
or UO_2 (O_2,N_2832,N_2916);
or UO_3 (O_3,N_2918,N_2847);
or UO_4 (O_4,N_2880,N_2839);
or UO_5 (O_5,N_2935,N_2961);
nor UO_6 (O_6,N_2915,N_2970);
and UO_7 (O_7,N_2884,N_2879);
nand UO_8 (O_8,N_2930,N_2952);
and UO_9 (O_9,N_2841,N_2825);
nor UO_10 (O_10,N_2967,N_2908);
xnor UO_11 (O_11,N_2936,N_2983);
or UO_12 (O_12,N_2833,N_2831);
nand UO_13 (O_13,N_2817,N_2933);
xor UO_14 (O_14,N_2972,N_2902);
nor UO_15 (O_15,N_2939,N_2876);
nand UO_16 (O_16,N_2962,N_2843);
and UO_17 (O_17,N_2920,N_2907);
nor UO_18 (O_18,N_2844,N_2824);
or UO_19 (O_19,N_2888,N_2974);
nand UO_20 (O_20,N_2955,N_2973);
nand UO_21 (O_21,N_2906,N_2875);
or UO_22 (O_22,N_2945,N_2904);
nand UO_23 (O_23,N_2956,N_2861);
nor UO_24 (O_24,N_2851,N_2984);
or UO_25 (O_25,N_2889,N_2997);
and UO_26 (O_26,N_2900,N_2807);
nor UO_27 (O_27,N_2995,N_2856);
and UO_28 (O_28,N_2850,N_2865);
nor UO_29 (O_29,N_2836,N_2985);
nor UO_30 (O_30,N_2813,N_2919);
or UO_31 (O_31,N_2924,N_2968);
or UO_32 (O_32,N_2835,N_2815);
nand UO_33 (O_33,N_2975,N_2914);
or UO_34 (O_34,N_2801,N_2863);
or UO_35 (O_35,N_2887,N_2982);
nand UO_36 (O_36,N_2822,N_2896);
and UO_37 (O_37,N_2966,N_2987);
nor UO_38 (O_38,N_2871,N_2855);
and UO_39 (O_39,N_2808,N_2944);
nand UO_40 (O_40,N_2834,N_2866);
nor UO_41 (O_41,N_2951,N_2811);
and UO_42 (O_42,N_2864,N_2910);
nand UO_43 (O_43,N_2960,N_2852);
nor UO_44 (O_44,N_2826,N_2846);
xor UO_45 (O_45,N_2954,N_2988);
nand UO_46 (O_46,N_2814,N_2909);
nand UO_47 (O_47,N_2860,N_2827);
and UO_48 (O_48,N_2823,N_2898);
nor UO_49 (O_49,N_2858,N_2840);
and UO_50 (O_50,N_2996,N_2977);
or UO_51 (O_51,N_2809,N_2940);
or UO_52 (O_52,N_2901,N_2941);
nor UO_53 (O_53,N_2803,N_2928);
nand UO_54 (O_54,N_2949,N_2965);
nor UO_55 (O_55,N_2927,N_2838);
and UO_56 (O_56,N_2842,N_2854);
nor UO_57 (O_57,N_2893,N_2829);
nand UO_58 (O_58,N_2883,N_2971);
nor UO_59 (O_59,N_2862,N_2926);
or UO_60 (O_60,N_2964,N_2867);
nand UO_61 (O_61,N_2819,N_2950);
or UO_62 (O_62,N_2905,N_2849);
nor UO_63 (O_63,N_2837,N_2937);
nor UO_64 (O_64,N_2925,N_2948);
nand UO_65 (O_65,N_2989,N_2891);
nor UO_66 (O_66,N_2991,N_2943);
and UO_67 (O_67,N_2886,N_2806);
or UO_68 (O_68,N_2932,N_2899);
nand UO_69 (O_69,N_2903,N_2959);
nor UO_70 (O_70,N_2877,N_2942);
nand UO_71 (O_71,N_2857,N_2878);
nor UO_72 (O_72,N_2882,N_2957);
and UO_73 (O_73,N_2947,N_2820);
and UO_74 (O_74,N_2830,N_2895);
nand UO_75 (O_75,N_2859,N_2998);
nor UO_76 (O_76,N_2881,N_2921);
nor UO_77 (O_77,N_2828,N_2853);
nor UO_78 (O_78,N_2870,N_2912);
and UO_79 (O_79,N_2818,N_2868);
or UO_80 (O_80,N_2805,N_2978);
or UO_81 (O_81,N_2845,N_2917);
nor UO_82 (O_82,N_2804,N_2872);
nand UO_83 (O_83,N_2873,N_2897);
or UO_84 (O_84,N_2980,N_2800);
and UO_85 (O_85,N_2812,N_2979);
nor UO_86 (O_86,N_2981,N_2934);
and UO_87 (O_87,N_2994,N_2816);
xnor UO_88 (O_88,N_2986,N_2802);
nor UO_89 (O_89,N_2869,N_2929);
nand UO_90 (O_90,N_2892,N_2923);
xnor UO_91 (O_91,N_2938,N_2946);
or UO_92 (O_92,N_2922,N_2890);
nor UO_93 (O_93,N_2963,N_2911);
nand UO_94 (O_94,N_2993,N_2953);
and UO_95 (O_95,N_2913,N_2848);
nor UO_96 (O_96,N_2894,N_2874);
nand UO_97 (O_97,N_2976,N_2992);
or UO_98 (O_98,N_2999,N_2931);
and UO_99 (O_99,N_2821,N_2958);
or UO_100 (O_100,N_2816,N_2856);
nand UO_101 (O_101,N_2992,N_2964);
and UO_102 (O_102,N_2912,N_2810);
and UO_103 (O_103,N_2923,N_2838);
or UO_104 (O_104,N_2976,N_2856);
and UO_105 (O_105,N_2882,N_2844);
nand UO_106 (O_106,N_2970,N_2953);
and UO_107 (O_107,N_2938,N_2832);
nor UO_108 (O_108,N_2932,N_2839);
or UO_109 (O_109,N_2835,N_2881);
nand UO_110 (O_110,N_2812,N_2868);
nand UO_111 (O_111,N_2995,N_2928);
and UO_112 (O_112,N_2947,N_2921);
or UO_113 (O_113,N_2964,N_2983);
nand UO_114 (O_114,N_2961,N_2949);
and UO_115 (O_115,N_2813,N_2874);
or UO_116 (O_116,N_2955,N_2833);
xnor UO_117 (O_117,N_2943,N_2941);
xor UO_118 (O_118,N_2954,N_2931);
nand UO_119 (O_119,N_2917,N_2954);
or UO_120 (O_120,N_2909,N_2977);
and UO_121 (O_121,N_2801,N_2872);
or UO_122 (O_122,N_2890,N_2821);
xor UO_123 (O_123,N_2827,N_2995);
and UO_124 (O_124,N_2868,N_2883);
or UO_125 (O_125,N_2936,N_2935);
nor UO_126 (O_126,N_2919,N_2998);
nor UO_127 (O_127,N_2857,N_2814);
and UO_128 (O_128,N_2936,N_2933);
or UO_129 (O_129,N_2996,N_2848);
or UO_130 (O_130,N_2874,N_2834);
nor UO_131 (O_131,N_2955,N_2814);
nor UO_132 (O_132,N_2982,N_2948);
nand UO_133 (O_133,N_2934,N_2852);
nor UO_134 (O_134,N_2994,N_2810);
nand UO_135 (O_135,N_2962,N_2912);
nand UO_136 (O_136,N_2941,N_2812);
nand UO_137 (O_137,N_2857,N_2911);
or UO_138 (O_138,N_2992,N_2952);
nand UO_139 (O_139,N_2891,N_2833);
or UO_140 (O_140,N_2842,N_2974);
nor UO_141 (O_141,N_2916,N_2978);
nand UO_142 (O_142,N_2926,N_2953);
nor UO_143 (O_143,N_2985,N_2891);
nor UO_144 (O_144,N_2864,N_2817);
and UO_145 (O_145,N_2800,N_2891);
nand UO_146 (O_146,N_2909,N_2940);
and UO_147 (O_147,N_2973,N_2838);
or UO_148 (O_148,N_2907,N_2820);
or UO_149 (O_149,N_2877,N_2991);
nand UO_150 (O_150,N_2836,N_2823);
nand UO_151 (O_151,N_2872,N_2937);
or UO_152 (O_152,N_2815,N_2823);
nand UO_153 (O_153,N_2929,N_2917);
or UO_154 (O_154,N_2827,N_2809);
nor UO_155 (O_155,N_2895,N_2956);
and UO_156 (O_156,N_2976,N_2988);
nor UO_157 (O_157,N_2878,N_2872);
xnor UO_158 (O_158,N_2822,N_2880);
nor UO_159 (O_159,N_2808,N_2884);
and UO_160 (O_160,N_2818,N_2889);
nand UO_161 (O_161,N_2895,N_2849);
nor UO_162 (O_162,N_2841,N_2933);
or UO_163 (O_163,N_2904,N_2962);
or UO_164 (O_164,N_2946,N_2921);
xnor UO_165 (O_165,N_2834,N_2846);
or UO_166 (O_166,N_2968,N_2900);
nand UO_167 (O_167,N_2950,N_2973);
and UO_168 (O_168,N_2995,N_2885);
and UO_169 (O_169,N_2847,N_2871);
nor UO_170 (O_170,N_2905,N_2987);
nor UO_171 (O_171,N_2858,N_2851);
and UO_172 (O_172,N_2879,N_2831);
and UO_173 (O_173,N_2825,N_2943);
and UO_174 (O_174,N_2971,N_2926);
or UO_175 (O_175,N_2975,N_2840);
nor UO_176 (O_176,N_2963,N_2828);
nand UO_177 (O_177,N_2929,N_2878);
nor UO_178 (O_178,N_2879,N_2821);
or UO_179 (O_179,N_2826,N_2897);
nor UO_180 (O_180,N_2992,N_2993);
or UO_181 (O_181,N_2821,N_2934);
nand UO_182 (O_182,N_2808,N_2980);
nand UO_183 (O_183,N_2892,N_2951);
nor UO_184 (O_184,N_2889,N_2844);
or UO_185 (O_185,N_2888,N_2844);
or UO_186 (O_186,N_2929,N_2930);
and UO_187 (O_187,N_2848,N_2987);
nand UO_188 (O_188,N_2876,N_2827);
and UO_189 (O_189,N_2889,N_2865);
nand UO_190 (O_190,N_2900,N_2949);
or UO_191 (O_191,N_2867,N_2854);
nor UO_192 (O_192,N_2800,N_2802);
and UO_193 (O_193,N_2890,N_2818);
or UO_194 (O_194,N_2915,N_2955);
nor UO_195 (O_195,N_2847,N_2912);
nand UO_196 (O_196,N_2951,N_2959);
nand UO_197 (O_197,N_2954,N_2992);
nor UO_198 (O_198,N_2806,N_2991);
and UO_199 (O_199,N_2905,N_2827);
and UO_200 (O_200,N_2870,N_2882);
or UO_201 (O_201,N_2911,N_2960);
nand UO_202 (O_202,N_2926,N_2863);
and UO_203 (O_203,N_2826,N_2887);
or UO_204 (O_204,N_2829,N_2925);
and UO_205 (O_205,N_2810,N_2906);
or UO_206 (O_206,N_2925,N_2964);
nor UO_207 (O_207,N_2941,N_2912);
and UO_208 (O_208,N_2992,N_2881);
and UO_209 (O_209,N_2956,N_2921);
nor UO_210 (O_210,N_2857,N_2869);
nor UO_211 (O_211,N_2918,N_2902);
nor UO_212 (O_212,N_2804,N_2956);
and UO_213 (O_213,N_2948,N_2952);
nand UO_214 (O_214,N_2857,N_2892);
and UO_215 (O_215,N_2843,N_2818);
or UO_216 (O_216,N_2948,N_2861);
and UO_217 (O_217,N_2935,N_2945);
and UO_218 (O_218,N_2831,N_2844);
and UO_219 (O_219,N_2993,N_2914);
nor UO_220 (O_220,N_2875,N_2966);
and UO_221 (O_221,N_2945,N_2844);
and UO_222 (O_222,N_2946,N_2917);
nand UO_223 (O_223,N_2919,N_2825);
and UO_224 (O_224,N_2856,N_2830);
nor UO_225 (O_225,N_2893,N_2872);
xor UO_226 (O_226,N_2923,N_2884);
nand UO_227 (O_227,N_2988,N_2862);
and UO_228 (O_228,N_2899,N_2826);
or UO_229 (O_229,N_2802,N_2950);
and UO_230 (O_230,N_2809,N_2964);
and UO_231 (O_231,N_2942,N_2914);
nor UO_232 (O_232,N_2922,N_2999);
or UO_233 (O_233,N_2904,N_2935);
or UO_234 (O_234,N_2914,N_2855);
and UO_235 (O_235,N_2804,N_2884);
nor UO_236 (O_236,N_2917,N_2975);
nor UO_237 (O_237,N_2956,N_2897);
or UO_238 (O_238,N_2895,N_2805);
or UO_239 (O_239,N_2974,N_2884);
or UO_240 (O_240,N_2994,N_2849);
or UO_241 (O_241,N_2964,N_2871);
and UO_242 (O_242,N_2936,N_2866);
nor UO_243 (O_243,N_2904,N_2882);
and UO_244 (O_244,N_2952,N_2976);
nor UO_245 (O_245,N_2868,N_2949);
nor UO_246 (O_246,N_2801,N_2820);
or UO_247 (O_247,N_2957,N_2983);
nand UO_248 (O_248,N_2999,N_2801);
nor UO_249 (O_249,N_2882,N_2893);
nand UO_250 (O_250,N_2855,N_2886);
nor UO_251 (O_251,N_2913,N_2826);
nor UO_252 (O_252,N_2958,N_2845);
or UO_253 (O_253,N_2964,N_2957);
nand UO_254 (O_254,N_2931,N_2922);
nand UO_255 (O_255,N_2859,N_2964);
nor UO_256 (O_256,N_2934,N_2866);
or UO_257 (O_257,N_2928,N_2866);
or UO_258 (O_258,N_2920,N_2810);
or UO_259 (O_259,N_2866,N_2996);
nor UO_260 (O_260,N_2861,N_2944);
nor UO_261 (O_261,N_2966,N_2963);
nand UO_262 (O_262,N_2945,N_2814);
nand UO_263 (O_263,N_2966,N_2992);
nand UO_264 (O_264,N_2907,N_2886);
nor UO_265 (O_265,N_2960,N_2846);
and UO_266 (O_266,N_2819,N_2908);
nor UO_267 (O_267,N_2828,N_2960);
or UO_268 (O_268,N_2900,N_2849);
nor UO_269 (O_269,N_2926,N_2860);
and UO_270 (O_270,N_2831,N_2814);
xor UO_271 (O_271,N_2805,N_2847);
or UO_272 (O_272,N_2897,N_2950);
nor UO_273 (O_273,N_2987,N_2883);
nand UO_274 (O_274,N_2957,N_2910);
nor UO_275 (O_275,N_2836,N_2830);
nor UO_276 (O_276,N_2968,N_2832);
nand UO_277 (O_277,N_2842,N_2812);
nand UO_278 (O_278,N_2816,N_2876);
nor UO_279 (O_279,N_2851,N_2848);
and UO_280 (O_280,N_2869,N_2922);
and UO_281 (O_281,N_2826,N_2868);
or UO_282 (O_282,N_2969,N_2815);
nand UO_283 (O_283,N_2899,N_2822);
nand UO_284 (O_284,N_2833,N_2804);
nor UO_285 (O_285,N_2869,N_2873);
or UO_286 (O_286,N_2870,N_2923);
or UO_287 (O_287,N_2803,N_2989);
nand UO_288 (O_288,N_2814,N_2898);
nor UO_289 (O_289,N_2958,N_2977);
and UO_290 (O_290,N_2938,N_2897);
or UO_291 (O_291,N_2987,N_2809);
nor UO_292 (O_292,N_2867,N_2863);
or UO_293 (O_293,N_2996,N_2897);
nand UO_294 (O_294,N_2818,N_2926);
nand UO_295 (O_295,N_2910,N_2978);
and UO_296 (O_296,N_2941,N_2810);
nor UO_297 (O_297,N_2859,N_2883);
nor UO_298 (O_298,N_2935,N_2838);
nor UO_299 (O_299,N_2908,N_2968);
and UO_300 (O_300,N_2954,N_2990);
and UO_301 (O_301,N_2883,N_2886);
nand UO_302 (O_302,N_2893,N_2861);
nand UO_303 (O_303,N_2834,N_2879);
and UO_304 (O_304,N_2810,N_2892);
or UO_305 (O_305,N_2809,N_2917);
or UO_306 (O_306,N_2892,N_2897);
and UO_307 (O_307,N_2867,N_2991);
nor UO_308 (O_308,N_2862,N_2949);
and UO_309 (O_309,N_2816,N_2969);
and UO_310 (O_310,N_2902,N_2885);
nand UO_311 (O_311,N_2864,N_2870);
nor UO_312 (O_312,N_2930,N_2949);
and UO_313 (O_313,N_2960,N_2831);
or UO_314 (O_314,N_2825,N_2880);
and UO_315 (O_315,N_2985,N_2851);
or UO_316 (O_316,N_2823,N_2818);
and UO_317 (O_317,N_2969,N_2941);
or UO_318 (O_318,N_2839,N_2941);
nand UO_319 (O_319,N_2980,N_2889);
or UO_320 (O_320,N_2832,N_2982);
or UO_321 (O_321,N_2903,N_2803);
nand UO_322 (O_322,N_2825,N_2827);
and UO_323 (O_323,N_2825,N_2961);
nand UO_324 (O_324,N_2937,N_2877);
nor UO_325 (O_325,N_2936,N_2953);
nand UO_326 (O_326,N_2904,N_2889);
nand UO_327 (O_327,N_2852,N_2996);
or UO_328 (O_328,N_2916,N_2966);
and UO_329 (O_329,N_2976,N_2824);
nand UO_330 (O_330,N_2899,N_2894);
or UO_331 (O_331,N_2964,N_2869);
or UO_332 (O_332,N_2936,N_2820);
and UO_333 (O_333,N_2815,N_2971);
or UO_334 (O_334,N_2924,N_2849);
nor UO_335 (O_335,N_2876,N_2979);
nor UO_336 (O_336,N_2848,N_2993);
nand UO_337 (O_337,N_2862,N_2914);
and UO_338 (O_338,N_2853,N_2896);
nor UO_339 (O_339,N_2884,N_2943);
and UO_340 (O_340,N_2867,N_2970);
nor UO_341 (O_341,N_2873,N_2953);
nand UO_342 (O_342,N_2841,N_2878);
nand UO_343 (O_343,N_2811,N_2962);
nor UO_344 (O_344,N_2930,N_2862);
or UO_345 (O_345,N_2890,N_2980);
and UO_346 (O_346,N_2951,N_2916);
nor UO_347 (O_347,N_2933,N_2814);
or UO_348 (O_348,N_2999,N_2961);
nor UO_349 (O_349,N_2998,N_2921);
or UO_350 (O_350,N_2979,N_2924);
nor UO_351 (O_351,N_2904,N_2975);
nor UO_352 (O_352,N_2978,N_2963);
nand UO_353 (O_353,N_2836,N_2963);
or UO_354 (O_354,N_2952,N_2957);
nor UO_355 (O_355,N_2901,N_2827);
nor UO_356 (O_356,N_2814,N_2900);
nand UO_357 (O_357,N_2960,N_2957);
nand UO_358 (O_358,N_2870,N_2973);
or UO_359 (O_359,N_2841,N_2888);
nand UO_360 (O_360,N_2807,N_2869);
or UO_361 (O_361,N_2930,N_2907);
and UO_362 (O_362,N_2951,N_2917);
nor UO_363 (O_363,N_2940,N_2918);
and UO_364 (O_364,N_2998,N_2962);
nand UO_365 (O_365,N_2974,N_2892);
nor UO_366 (O_366,N_2858,N_2818);
nand UO_367 (O_367,N_2960,N_2997);
and UO_368 (O_368,N_2835,N_2921);
or UO_369 (O_369,N_2881,N_2855);
nand UO_370 (O_370,N_2933,N_2804);
nor UO_371 (O_371,N_2834,N_2937);
nand UO_372 (O_372,N_2861,N_2882);
nand UO_373 (O_373,N_2825,N_2906);
and UO_374 (O_374,N_2953,N_2840);
nand UO_375 (O_375,N_2824,N_2966);
nand UO_376 (O_376,N_2849,N_2995);
nand UO_377 (O_377,N_2803,N_2897);
nor UO_378 (O_378,N_2878,N_2955);
xor UO_379 (O_379,N_2849,N_2922);
or UO_380 (O_380,N_2924,N_2811);
nand UO_381 (O_381,N_2826,N_2830);
nor UO_382 (O_382,N_2828,N_2834);
and UO_383 (O_383,N_2807,N_2934);
or UO_384 (O_384,N_2886,N_2978);
nand UO_385 (O_385,N_2875,N_2817);
xor UO_386 (O_386,N_2936,N_2802);
or UO_387 (O_387,N_2962,N_2896);
nand UO_388 (O_388,N_2962,N_2837);
nor UO_389 (O_389,N_2887,N_2859);
and UO_390 (O_390,N_2986,N_2823);
and UO_391 (O_391,N_2838,N_2839);
nor UO_392 (O_392,N_2888,N_2937);
nor UO_393 (O_393,N_2869,N_2803);
nor UO_394 (O_394,N_2929,N_2984);
nor UO_395 (O_395,N_2869,N_2997);
nor UO_396 (O_396,N_2862,N_2977);
or UO_397 (O_397,N_2916,N_2868);
nand UO_398 (O_398,N_2830,N_2971);
nor UO_399 (O_399,N_2889,N_2973);
nand UO_400 (O_400,N_2951,N_2899);
and UO_401 (O_401,N_2859,N_2844);
and UO_402 (O_402,N_2889,N_2908);
and UO_403 (O_403,N_2894,N_2986);
and UO_404 (O_404,N_2993,N_2905);
xor UO_405 (O_405,N_2908,N_2905);
and UO_406 (O_406,N_2881,N_2826);
nand UO_407 (O_407,N_2843,N_2834);
nor UO_408 (O_408,N_2853,N_2930);
nand UO_409 (O_409,N_2897,N_2877);
nand UO_410 (O_410,N_2900,N_2970);
nor UO_411 (O_411,N_2887,N_2831);
nand UO_412 (O_412,N_2970,N_2847);
and UO_413 (O_413,N_2995,N_2889);
and UO_414 (O_414,N_2982,N_2980);
or UO_415 (O_415,N_2936,N_2844);
nor UO_416 (O_416,N_2944,N_2970);
nor UO_417 (O_417,N_2830,N_2959);
nand UO_418 (O_418,N_2956,N_2972);
nand UO_419 (O_419,N_2993,N_2876);
nand UO_420 (O_420,N_2825,N_2975);
xnor UO_421 (O_421,N_2845,N_2863);
and UO_422 (O_422,N_2907,N_2877);
nand UO_423 (O_423,N_2842,N_2990);
xor UO_424 (O_424,N_2883,N_2996);
nor UO_425 (O_425,N_2899,N_2977);
nand UO_426 (O_426,N_2992,N_2810);
and UO_427 (O_427,N_2843,N_2855);
nand UO_428 (O_428,N_2864,N_2868);
and UO_429 (O_429,N_2912,N_2857);
nor UO_430 (O_430,N_2969,N_2964);
and UO_431 (O_431,N_2922,N_2954);
nor UO_432 (O_432,N_2806,N_2959);
nand UO_433 (O_433,N_2842,N_2892);
or UO_434 (O_434,N_2957,N_2858);
or UO_435 (O_435,N_2987,N_2929);
and UO_436 (O_436,N_2923,N_2806);
or UO_437 (O_437,N_2879,N_2863);
nor UO_438 (O_438,N_2911,N_2884);
and UO_439 (O_439,N_2838,N_2825);
and UO_440 (O_440,N_2979,N_2984);
xor UO_441 (O_441,N_2811,N_2805);
and UO_442 (O_442,N_2926,N_2802);
and UO_443 (O_443,N_2863,N_2935);
nor UO_444 (O_444,N_2894,N_2998);
nor UO_445 (O_445,N_2909,N_2837);
nand UO_446 (O_446,N_2830,N_2944);
nand UO_447 (O_447,N_2930,N_2846);
and UO_448 (O_448,N_2909,N_2944);
or UO_449 (O_449,N_2944,N_2993);
nand UO_450 (O_450,N_2996,N_2833);
or UO_451 (O_451,N_2891,N_2972);
or UO_452 (O_452,N_2840,N_2813);
and UO_453 (O_453,N_2815,N_2983);
and UO_454 (O_454,N_2873,N_2822);
and UO_455 (O_455,N_2936,N_2848);
nand UO_456 (O_456,N_2912,N_2920);
nor UO_457 (O_457,N_2847,N_2974);
and UO_458 (O_458,N_2809,N_2861);
nand UO_459 (O_459,N_2848,N_2868);
xnor UO_460 (O_460,N_2907,N_2972);
nand UO_461 (O_461,N_2982,N_2830);
or UO_462 (O_462,N_2856,N_2940);
nand UO_463 (O_463,N_2903,N_2885);
nand UO_464 (O_464,N_2801,N_2904);
or UO_465 (O_465,N_2947,N_2822);
and UO_466 (O_466,N_2891,N_2842);
nand UO_467 (O_467,N_2982,N_2936);
or UO_468 (O_468,N_2908,N_2864);
or UO_469 (O_469,N_2836,N_2984);
and UO_470 (O_470,N_2928,N_2885);
or UO_471 (O_471,N_2971,N_2861);
nor UO_472 (O_472,N_2869,N_2876);
and UO_473 (O_473,N_2959,N_2927);
nor UO_474 (O_474,N_2871,N_2901);
or UO_475 (O_475,N_2966,N_2908);
or UO_476 (O_476,N_2950,N_2817);
nand UO_477 (O_477,N_2854,N_2949);
and UO_478 (O_478,N_2961,N_2966);
nor UO_479 (O_479,N_2895,N_2920);
or UO_480 (O_480,N_2943,N_2939);
or UO_481 (O_481,N_2956,N_2849);
nor UO_482 (O_482,N_2886,N_2890);
and UO_483 (O_483,N_2871,N_2881);
and UO_484 (O_484,N_2896,N_2872);
and UO_485 (O_485,N_2995,N_2954);
nor UO_486 (O_486,N_2942,N_2948);
and UO_487 (O_487,N_2839,N_2993);
nand UO_488 (O_488,N_2977,N_2800);
or UO_489 (O_489,N_2808,N_2940);
nand UO_490 (O_490,N_2973,N_2989);
nand UO_491 (O_491,N_2837,N_2920);
and UO_492 (O_492,N_2918,N_2826);
or UO_493 (O_493,N_2867,N_2979);
nor UO_494 (O_494,N_2918,N_2990);
and UO_495 (O_495,N_2988,N_2872);
or UO_496 (O_496,N_2829,N_2844);
nand UO_497 (O_497,N_2978,N_2896);
nand UO_498 (O_498,N_2965,N_2801);
or UO_499 (O_499,N_2917,N_2873);
endmodule