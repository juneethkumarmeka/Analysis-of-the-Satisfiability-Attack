module basic_1500_15000_2000_20_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1269,In_940);
nand U1 (N_1,In_1472,In_563);
xnor U2 (N_2,In_1156,In_938);
nor U3 (N_3,In_554,In_248);
nor U4 (N_4,In_1370,In_787);
nand U5 (N_5,In_1401,In_1356);
nand U6 (N_6,In_756,In_1237);
nand U7 (N_7,In_1015,In_883);
or U8 (N_8,In_813,In_1268);
and U9 (N_9,In_906,In_183);
and U10 (N_10,In_1173,In_1137);
nor U11 (N_11,In_1079,In_305);
and U12 (N_12,In_1481,In_1125);
and U13 (N_13,In_1376,In_1064);
nor U14 (N_14,In_535,In_247);
or U15 (N_15,In_1053,In_1328);
nand U16 (N_16,In_406,In_362);
nand U17 (N_17,In_1458,In_503);
and U18 (N_18,In_23,In_594);
or U19 (N_19,In_221,In_489);
nand U20 (N_20,In_346,In_1442);
nand U21 (N_21,In_1367,In_433);
and U22 (N_22,In_359,In_1469);
nand U23 (N_23,In_1341,In_1478);
or U24 (N_24,In_292,In_916);
nand U25 (N_25,In_479,In_157);
nand U26 (N_26,In_799,In_1228);
and U27 (N_27,In_1017,In_77);
nand U28 (N_28,In_807,In_439);
nand U29 (N_29,In_1194,In_715);
or U30 (N_30,In_261,In_899);
and U31 (N_31,In_1471,In_1062);
and U32 (N_32,In_354,In_925);
or U33 (N_33,In_901,In_605);
nand U34 (N_34,In_1362,In_403);
nor U35 (N_35,In_431,In_1084);
xnor U36 (N_36,In_198,In_910);
nand U37 (N_37,In_919,In_720);
or U38 (N_38,In_1457,In_1135);
nand U39 (N_39,In_487,In_1291);
and U40 (N_40,In_1298,In_338);
nor U41 (N_41,In_161,In_735);
nor U42 (N_42,In_397,In_254);
nand U43 (N_43,In_1300,In_131);
or U44 (N_44,In_709,In_747);
nand U45 (N_45,In_805,In_1495);
and U46 (N_46,In_1180,In_1212);
and U47 (N_47,In_381,In_1290);
and U48 (N_48,In_231,In_360);
nand U49 (N_49,In_852,In_591);
nand U50 (N_50,In_33,In_57);
and U51 (N_51,In_1490,In_669);
and U52 (N_52,In_1106,In_267);
and U53 (N_53,In_417,In_1468);
or U54 (N_54,In_998,In_323);
or U55 (N_55,In_1359,In_481);
nor U56 (N_56,In_507,In_20);
or U57 (N_57,In_956,In_301);
and U58 (N_58,In_1092,In_1216);
and U59 (N_59,In_763,In_19);
and U60 (N_60,In_789,In_1195);
nor U61 (N_61,In_449,In_544);
and U62 (N_62,In_1201,In_628);
or U63 (N_63,In_1229,In_56);
nand U64 (N_64,In_2,In_1455);
nand U65 (N_65,In_1494,In_136);
and U66 (N_66,In_376,In_1444);
or U67 (N_67,In_964,In_336);
nor U68 (N_68,In_436,In_378);
nor U69 (N_69,In_55,In_818);
or U70 (N_70,In_1060,In_643);
xnor U71 (N_71,In_1040,In_526);
nand U72 (N_72,In_275,In_559);
nand U73 (N_73,In_438,In_918);
nor U74 (N_74,In_38,In_114);
or U75 (N_75,In_861,In_86);
or U76 (N_76,In_92,In_1235);
and U77 (N_77,In_802,In_42);
nor U78 (N_78,In_686,In_877);
and U79 (N_79,In_636,In_1221);
or U80 (N_80,In_281,In_1334);
nor U81 (N_81,In_164,In_537);
nand U82 (N_82,In_350,In_600);
and U83 (N_83,In_1012,In_566);
nor U84 (N_84,In_592,In_59);
and U85 (N_85,In_1406,In_966);
or U86 (N_86,In_105,In_768);
xnor U87 (N_87,In_493,In_97);
or U88 (N_88,In_188,In_478);
nor U89 (N_89,In_588,In_147);
nor U90 (N_90,In_837,In_200);
and U91 (N_91,In_0,In_1282);
xor U92 (N_92,In_1332,In_210);
nor U93 (N_93,In_945,In_1355);
xnor U94 (N_94,In_1166,In_662);
nor U95 (N_95,In_93,In_490);
or U96 (N_96,In_150,In_72);
or U97 (N_97,In_538,In_485);
nand U98 (N_98,In_99,In_1473);
or U99 (N_99,In_345,In_1072);
nor U100 (N_100,In_1151,In_262);
or U101 (N_101,In_1435,In_1443);
nand U102 (N_102,In_313,In_1417);
and U103 (N_103,In_1105,In_408);
and U104 (N_104,In_108,In_565);
nand U105 (N_105,In_604,In_1198);
and U106 (N_106,In_1054,In_280);
xnor U107 (N_107,In_1134,In_829);
nor U108 (N_108,In_295,In_671);
nor U109 (N_109,In_981,In_238);
and U110 (N_110,In_415,In_933);
or U111 (N_111,In_1096,In_50);
and U112 (N_112,In_218,In_923);
xor U113 (N_113,In_355,In_1424);
and U114 (N_114,In_285,In_865);
or U115 (N_115,In_1460,In_911);
and U116 (N_116,In_1144,In_920);
nor U117 (N_117,In_1475,In_539);
nand U118 (N_118,In_995,In_251);
or U119 (N_119,In_637,In_297);
nand U120 (N_120,In_767,In_759);
nor U121 (N_121,In_95,In_1391);
xnor U122 (N_122,In_755,In_1489);
nor U123 (N_123,In_53,In_371);
xor U124 (N_124,In_1496,In_508);
nor U125 (N_125,In_991,In_1085);
nor U126 (N_126,In_340,In_731);
or U127 (N_127,In_639,In_894);
and U128 (N_128,In_1352,In_309);
or U129 (N_129,In_1372,In_1465);
nand U130 (N_130,In_722,In_326);
nand U131 (N_131,In_575,In_927);
nand U132 (N_132,In_265,In_1462);
or U133 (N_133,In_402,In_445);
nor U134 (N_134,In_1030,In_1021);
nand U135 (N_135,In_973,In_178);
nand U136 (N_136,In_546,In_1175);
or U137 (N_137,In_548,In_830);
xnor U138 (N_138,In_1243,In_1075);
or U139 (N_139,In_723,In_458);
and U140 (N_140,In_252,In_1093);
nor U141 (N_141,In_1078,In_881);
or U142 (N_142,In_1108,In_66);
nor U143 (N_143,In_68,In_838);
nand U144 (N_144,In_62,In_528);
or U145 (N_145,In_74,In_393);
nor U146 (N_146,In_1178,In_989);
nor U147 (N_147,In_388,In_851);
or U148 (N_148,In_957,In_848);
or U149 (N_149,In_1218,In_1209);
nor U150 (N_150,In_692,In_176);
nor U151 (N_151,In_844,In_1052);
or U152 (N_152,In_840,In_680);
or U153 (N_153,In_1095,In_219);
nand U154 (N_154,In_1136,In_587);
or U155 (N_155,In_1147,In_513);
xor U156 (N_156,In_929,In_687);
and U157 (N_157,In_1275,In_1110);
nor U158 (N_158,In_1142,In_1239);
xor U159 (N_159,In_629,In_1009);
or U160 (N_160,In_540,In_125);
xnor U161 (N_161,In_703,In_810);
or U162 (N_162,In_1326,In_761);
nor U163 (N_163,In_660,In_373);
or U164 (N_164,In_812,In_199);
nand U165 (N_165,In_902,In_542);
xor U166 (N_166,In_1338,In_1283);
and U167 (N_167,In_1348,In_1279);
nand U168 (N_168,In_578,In_205);
or U169 (N_169,In_650,In_843);
xnor U170 (N_170,In_886,In_1187);
nand U171 (N_171,In_6,In_1396);
or U172 (N_172,In_98,In_783);
nor U173 (N_173,In_1158,In_1482);
nand U174 (N_174,In_530,In_800);
nand U175 (N_175,In_1028,In_1407);
xor U176 (N_176,In_633,In_12);
or U177 (N_177,In_1033,In_704);
nor U178 (N_178,In_1224,In_1385);
or U179 (N_179,In_612,In_1247);
xnor U180 (N_180,In_987,In_480);
or U181 (N_181,In_863,In_127);
and U182 (N_182,In_889,In_120);
or U183 (N_183,In_1265,In_524);
and U184 (N_184,In_873,In_651);
or U185 (N_185,In_483,In_593);
or U186 (N_186,In_970,In_377);
and U187 (N_187,In_646,In_884);
nand U188 (N_188,In_774,In_366);
nor U189 (N_189,In_182,In_517);
nand U190 (N_190,In_1303,In_616);
and U191 (N_191,In_472,In_197);
nand U192 (N_192,In_369,In_240);
or U193 (N_193,In_208,In_1335);
nand U194 (N_194,In_888,In_1321);
xnor U195 (N_195,In_745,In_522);
and U196 (N_196,In_809,In_1313);
nand U197 (N_197,In_1358,In_908);
nand U198 (N_198,In_1289,In_220);
and U199 (N_199,In_85,In_795);
or U200 (N_200,In_892,In_241);
or U201 (N_201,In_1382,In_443);
or U202 (N_202,In_440,In_1309);
and U203 (N_203,In_728,In_4);
nor U204 (N_204,In_597,In_1488);
and U205 (N_205,In_337,In_342);
nand U206 (N_206,In_214,In_1434);
nor U207 (N_207,In_1467,In_316);
nand U208 (N_208,In_1422,In_287);
and U209 (N_209,In_1154,In_124);
and U210 (N_210,In_678,In_574);
and U211 (N_211,In_425,In_893);
or U212 (N_212,In_1423,In_794);
and U213 (N_213,In_60,In_1034);
nor U214 (N_214,In_571,In_765);
or U215 (N_215,In_1246,In_1206);
nand U216 (N_216,In_54,In_24);
nand U217 (N_217,In_414,In_1199);
nand U218 (N_218,In_151,In_1409);
nand U219 (N_219,In_630,In_1403);
or U220 (N_220,In_103,In_567);
nand U221 (N_221,In_467,In_963);
xnor U222 (N_222,In_132,In_1013);
or U223 (N_223,In_341,In_428);
nand U224 (N_224,In_882,In_1447);
or U225 (N_225,In_333,In_652);
xnor U226 (N_226,In_1055,In_519);
nor U227 (N_227,In_885,In_90);
and U228 (N_228,In_1164,In_1076);
nand U229 (N_229,In_259,In_1416);
xor U230 (N_230,In_642,In_1051);
nor U231 (N_231,In_798,In_714);
xor U232 (N_232,In_497,In_1306);
or U233 (N_233,In_1018,In_613);
nor U234 (N_234,In_321,In_96);
nand U235 (N_235,In_1254,In_1296);
nor U236 (N_236,In_43,In_1128);
or U237 (N_237,In_107,In_717);
nand U238 (N_238,In_654,In_895);
and U239 (N_239,In_627,In_831);
nand U240 (N_240,In_1251,In_121);
nor U241 (N_241,In_368,In_435);
nor U242 (N_242,In_1188,In_1253);
or U243 (N_243,In_191,In_904);
xnor U244 (N_244,In_974,In_1207);
nand U245 (N_245,In_781,In_780);
nand U246 (N_246,In_585,In_1077);
and U247 (N_247,In_1412,In_1477);
and U248 (N_248,In_734,In_282);
or U249 (N_249,In_769,In_444);
or U250 (N_250,In_1058,In_772);
nor U251 (N_251,In_1420,In_1167);
and U252 (N_252,In_398,In_1091);
and U253 (N_253,In_931,In_1157);
nor U254 (N_254,In_665,In_1171);
and U255 (N_255,In_1205,In_1162);
and U256 (N_256,In_793,In_1336);
or U257 (N_257,In_803,In_1386);
or U258 (N_258,In_502,In_1257);
nand U259 (N_259,In_1418,In_471);
nor U260 (N_260,In_101,In_460);
nand U261 (N_261,In_641,In_1);
and U262 (N_262,In_367,In_169);
nand U263 (N_263,In_739,In_782);
or U264 (N_264,In_201,In_160);
nor U265 (N_265,In_317,In_1193);
xnor U266 (N_266,In_422,In_1446);
nand U267 (N_267,In_527,In_328);
or U268 (N_268,In_283,In_73);
and U269 (N_269,In_79,In_580);
or U270 (N_270,In_999,In_534);
or U271 (N_271,In_626,In_119);
nand U272 (N_272,In_832,In_356);
and U273 (N_273,In_1031,In_757);
xnor U274 (N_274,In_145,In_590);
nor U275 (N_275,In_977,In_318);
and U276 (N_276,In_1181,In_1320);
nor U277 (N_277,In_1003,In_579);
nor U278 (N_278,In_1277,In_1274);
nor U279 (N_279,In_155,In_615);
nor U280 (N_280,In_673,In_421);
xor U281 (N_281,In_82,In_1324);
or U282 (N_282,In_13,In_1002);
nor U283 (N_283,In_635,In_335);
nor U284 (N_284,In_196,In_1057);
nand U285 (N_285,In_1441,In_63);
and U286 (N_286,In_212,In_1450);
nor U287 (N_287,In_250,In_1059);
nor U288 (N_288,In_1360,In_18);
nand U289 (N_289,In_903,In_410);
and U290 (N_290,In_1448,In_1264);
or U291 (N_291,In_496,In_1429);
nand U292 (N_292,In_1163,In_608);
and U293 (N_293,In_348,In_162);
and U294 (N_294,In_744,In_239);
nor U295 (N_295,In_937,In_1067);
xor U296 (N_296,In_330,In_917);
nor U297 (N_297,In_405,In_584);
xnor U298 (N_298,In_1208,In_984);
xor U299 (N_299,In_972,In_1350);
or U300 (N_300,In_1089,In_1025);
nor U301 (N_301,In_1373,In_1349);
and U302 (N_302,In_1153,In_531);
and U303 (N_303,In_666,In_953);
or U304 (N_304,In_1214,In_117);
nor U305 (N_305,In_694,In_1252);
nor U306 (N_306,In_272,In_543);
xor U307 (N_307,In_29,In_1318);
nand U308 (N_308,In_1408,In_40);
xnor U309 (N_309,In_1241,In_839);
or U310 (N_310,In_257,In_568);
or U311 (N_311,In_1392,In_320);
or U312 (N_312,In_1314,In_1400);
or U313 (N_313,In_549,In_374);
nor U314 (N_314,In_1184,In_10);
or U315 (N_315,In_1232,In_1046);
nand U316 (N_316,In_1043,In_175);
and U317 (N_317,In_946,In_1389);
nor U318 (N_318,In_944,In_674);
and U319 (N_319,In_1363,In_299);
nor U320 (N_320,In_707,In_510);
and U321 (N_321,In_1056,In_951);
nor U322 (N_322,In_1019,In_187);
and U323 (N_323,In_557,In_258);
nor U324 (N_324,In_1319,In_1159);
nor U325 (N_325,In_1236,In_603);
nor U326 (N_326,In_791,In_142);
and U327 (N_327,In_558,In_907);
nor U328 (N_328,In_514,In_296);
nand U329 (N_329,In_1189,In_1172);
nand U330 (N_330,In_833,In_1127);
xor U331 (N_331,In_1215,In_475);
nor U332 (N_332,In_1222,In_311);
xor U333 (N_333,In_244,In_137);
and U334 (N_334,In_749,In_1393);
nor U335 (N_335,In_488,In_961);
nor U336 (N_336,In_1177,In_228);
or U337 (N_337,In_1390,In_994);
nand U338 (N_338,In_1087,In_180);
nor U339 (N_339,In_658,In_1197);
and U340 (N_340,In_1001,In_21);
nand U341 (N_341,In_766,In_1345);
nor U342 (N_342,In_820,In_1285);
and U343 (N_343,In_876,In_771);
nor U344 (N_344,In_1433,In_112);
and U345 (N_345,In_857,In_122);
and U346 (N_346,In_599,In_491);
or U347 (N_347,In_1061,In_1068);
nand U348 (N_348,In_1427,In_1259);
nor U349 (N_349,In_869,In_203);
or U350 (N_350,In_391,In_75);
or U351 (N_351,In_1383,In_35);
xnor U352 (N_352,In_1404,In_319);
or U353 (N_353,In_1016,In_968);
or U354 (N_354,In_100,In_610);
nand U355 (N_355,In_456,In_790);
or U356 (N_356,In_1452,In_154);
nand U357 (N_357,In_733,In_1398);
nand U358 (N_358,In_15,In_675);
or U359 (N_359,In_466,In_828);
xor U360 (N_360,In_1364,In_454);
nand U361 (N_361,In_255,In_1027);
nand U362 (N_362,In_382,In_1463);
or U363 (N_363,In_279,In_740);
nor U364 (N_364,In_1331,In_486);
nor U365 (N_365,In_506,In_1032);
nor U366 (N_366,In_236,In_695);
and U367 (N_367,In_80,In_1491);
and U368 (N_368,In_725,In_1413);
nand U369 (N_369,In_814,In_773);
nor U370 (N_370,In_511,In_389);
nor U371 (N_371,In_1371,In_606);
nand U372 (N_372,In_880,In_817);
nor U373 (N_373,In_484,In_195);
and U374 (N_374,In_8,In_291);
nand U375 (N_375,In_455,In_609);
nor U376 (N_376,In_343,In_801);
nor U377 (N_377,In_560,In_1453);
nor U378 (N_378,In_332,In_862);
or U379 (N_379,In_173,In_181);
or U380 (N_380,In_249,In_1288);
nand U381 (N_381,In_1007,In_589);
or U382 (N_382,In_777,In_1354);
xor U383 (N_383,In_290,In_1036);
and U384 (N_384,In_1168,In_515);
or U385 (N_385,In_947,In_632);
and U386 (N_386,In_1081,In_668);
or U387 (N_387,In_583,In_845);
xnor U388 (N_388,In_648,In_1459);
nor U389 (N_389,In_909,In_1339);
nor U390 (N_390,In_1273,In_457);
nor U391 (N_391,In_1483,In_811);
xor U392 (N_392,In_1185,In_1063);
nor U393 (N_393,In_732,In_891);
nor U394 (N_394,In_225,In_380);
nor U395 (N_395,In_1299,In_1148);
and U396 (N_396,In_217,In_143);
and U397 (N_397,In_268,In_582);
nand U398 (N_398,In_303,In_165);
or U399 (N_399,In_1486,In_1100);
or U400 (N_400,In_992,In_640);
or U401 (N_401,In_806,In_743);
nand U402 (N_402,In_1297,In_1261);
or U403 (N_403,In_213,In_516);
and U404 (N_404,In_14,In_1426);
and U405 (N_405,In_278,In_1026);
nor U406 (N_406,In_1124,In_270);
or U407 (N_407,In_1470,In_1461);
nand U408 (N_408,In_713,In_102);
nor U409 (N_409,In_499,In_357);
and U410 (N_410,In_437,In_624);
or U411 (N_411,In_1112,In_409);
nand U412 (N_412,In_363,In_158);
nand U413 (N_413,In_1113,In_1022);
or U414 (N_414,In_847,In_1484);
and U415 (N_415,In_1118,In_685);
nand U416 (N_416,In_1329,In_140);
and U417 (N_417,In_276,In_928);
and U418 (N_418,In_1226,In_392);
nor U419 (N_419,In_495,In_1161);
nor U420 (N_420,In_1301,In_741);
nand U421 (N_421,In_498,In_688);
nor U422 (N_422,In_206,In_962);
or U423 (N_423,In_504,In_61);
nand U424 (N_424,In_215,In_352);
or U425 (N_425,In_1248,In_407);
or U426 (N_426,In_1107,In_1141);
or U427 (N_427,In_1263,In_958);
or U428 (N_428,In_1451,In_1238);
nand U429 (N_429,In_778,In_1456);
and U430 (N_430,In_706,In_78);
or U431 (N_431,In_1430,In_693);
nor U432 (N_432,In_395,In_148);
nand U433 (N_433,In_420,In_174);
and U434 (N_434,In_1333,In_1109);
nor U435 (N_435,In_1271,In_816);
nor U436 (N_436,In_618,In_1365);
and U437 (N_437,In_1280,In_752);
or U438 (N_438,In_664,In_94);
and U439 (N_439,In_1270,In_264);
or U440 (N_440,In_647,In_598);
and U441 (N_441,In_266,In_1316);
and U442 (N_442,In_533,In_116);
or U443 (N_443,In_1449,In_1351);
nor U444 (N_444,In_1287,In_7);
or U445 (N_445,In_727,In_1381);
or U446 (N_446,In_941,In_39);
or U447 (N_447,In_1311,In_705);
or U448 (N_448,In_413,In_1049);
nor U449 (N_449,In_224,In_1202);
and U450 (N_450,In_737,In_602);
nor U451 (N_451,In_596,In_1074);
or U452 (N_452,In_1099,In_430);
and U453 (N_453,In_172,In_620);
xor U454 (N_454,In_625,In_564);
and U455 (N_455,In_726,In_211);
and U456 (N_456,In_163,In_28);
or U457 (N_457,In_1244,In_1070);
or U458 (N_458,In_943,In_520);
or U459 (N_459,In_509,In_361);
or U460 (N_460,In_325,In_912);
and U461 (N_461,In_1405,In_146);
and U462 (N_462,In_1284,In_835);
or U463 (N_463,In_846,In_450);
and U464 (N_464,In_1230,In_1262);
nand U465 (N_465,In_860,In_521);
and U466 (N_466,In_327,In_27);
nor U467 (N_467,In_89,In_1485);
nand U468 (N_468,In_1256,In_135);
or U469 (N_469,In_83,In_677);
nand U470 (N_470,In_1010,In_1117);
xnor U471 (N_471,In_1191,In_1304);
and U472 (N_472,In_1170,In_447);
nand U473 (N_473,In_1139,In_952);
and U474 (N_474,In_1425,In_84);
and U475 (N_475,In_879,In_1375);
nand U476 (N_476,In_271,In_1169);
and U477 (N_477,In_37,In_379);
or U478 (N_478,In_128,In_253);
nand U479 (N_479,In_1323,In_474);
or U480 (N_480,In_915,In_1384);
nor U481 (N_481,In_314,In_47);
and U482 (N_482,In_1366,In_286);
or U483 (N_483,In_1152,In_1165);
or U484 (N_484,In_45,In_87);
nor U485 (N_485,In_302,In_1006);
or U486 (N_486,In_1088,In_708);
and U487 (N_487,In_711,In_996);
and U488 (N_488,In_729,In_1103);
nor U489 (N_489,In_1097,In_193);
and U490 (N_490,In_670,In_227);
and U491 (N_491,In_661,In_553);
or U492 (N_492,In_611,In_1149);
and U493 (N_493,In_1213,In_1278);
and U494 (N_494,In_716,In_190);
xnor U495 (N_495,In_432,In_601);
and U496 (N_496,In_573,In_468);
or U497 (N_497,In_1104,In_788);
nor U498 (N_498,In_1227,In_1024);
and U499 (N_499,In_1102,In_969);
or U500 (N_500,In_289,In_934);
nand U501 (N_501,In_260,In_1122);
nor U502 (N_502,In_322,In_505);
nor U503 (N_503,In_166,In_825);
nand U504 (N_504,In_1120,In_887);
or U505 (N_505,In_230,In_1260);
or U506 (N_506,In_1415,In_742);
or U507 (N_507,In_1242,In_653);
and U508 (N_508,In_1044,In_858);
nand U509 (N_509,In_753,In_1037);
nor U510 (N_510,In_736,In_1000);
or U511 (N_511,In_1203,In_3);
or U512 (N_512,In_896,In_866);
or U513 (N_513,In_469,In_149);
xnor U514 (N_514,In_70,In_1042);
and U515 (N_515,In_1369,In_1307);
and U516 (N_516,In_1344,In_1234);
nand U517 (N_517,In_470,In_294);
or U518 (N_518,In_797,In_905);
and U519 (N_519,In_91,In_1126);
nor U520 (N_520,In_898,In_914);
and U521 (N_521,In_1292,In_1445);
and U522 (N_522,In_932,In_463);
xor U523 (N_523,In_856,In_1245);
or U524 (N_524,In_1123,In_855);
nor U525 (N_525,In_1387,In_1065);
or U526 (N_526,In_1421,In_1397);
xor U527 (N_527,In_288,In_922);
and U528 (N_528,In_69,In_532);
and U529 (N_529,In_1498,In_245);
nor U530 (N_530,In_523,In_1431);
nand U531 (N_531,In_26,In_353);
nand U532 (N_532,In_17,In_1272);
nor U533 (N_533,In_207,In_383);
and U534 (N_534,In_339,In_1402);
and U535 (N_535,In_298,In_775);
nor U536 (N_536,In_1295,In_1183);
xnor U537 (N_537,In_11,In_1454);
nor U538 (N_538,In_482,In_134);
nand U539 (N_539,In_690,In_1132);
nor U540 (N_540,In_418,In_141);
or U541 (N_541,In_784,In_1432);
nor U542 (N_542,In_1308,In_529);
nand U543 (N_543,In_1394,In_65);
and U544 (N_544,In_667,In_948);
or U545 (N_545,In_139,In_1305);
xor U546 (N_546,In_1150,In_751);
xnor U547 (N_547,In_955,In_1240);
nor U548 (N_548,In_386,In_426);
nand U549 (N_549,In_525,In_698);
nor U550 (N_550,In_1347,In_477);
or U551 (N_551,In_1281,In_785);
nor U552 (N_552,In_1330,In_442);
nand U553 (N_553,In_209,In_644);
nor U554 (N_554,In_451,In_1499);
nor U555 (N_555,In_1090,In_129);
nor U556 (N_556,In_1436,In_5);
xnor U557 (N_557,In_1176,In_779);
xor U558 (N_558,In_949,In_461);
and U559 (N_559,In_171,In_459);
and U560 (N_560,In_700,In_1121);
nor U561 (N_561,In_351,In_619);
and U562 (N_562,In_699,In_1050);
nor U563 (N_563,In_545,In_1302);
and U564 (N_564,In_144,In_555);
nor U565 (N_565,In_344,In_758);
nand U566 (N_566,In_547,In_1145);
or U567 (N_567,In_234,In_364);
nor U568 (N_568,In_126,In_1266);
xnor U569 (N_569,In_36,In_168);
and U570 (N_570,In_419,In_821);
nor U571 (N_571,In_1492,In_304);
nor U572 (N_572,In_315,In_394);
nor U573 (N_573,In_1439,In_390);
nor U574 (N_574,In_649,In_446);
nor U575 (N_575,In_384,In_1337);
nand U576 (N_576,In_192,In_153);
nand U577 (N_577,In_256,In_978);
or U578 (N_578,In_233,In_277);
and U579 (N_579,In_853,In_997);
or U580 (N_580,In_1038,In_1190);
and U581 (N_581,In_659,In_577);
nor U582 (N_582,In_1428,In_1476);
or U583 (N_583,In_111,In_656);
and U584 (N_584,In_681,In_827);
xor U585 (N_585,In_399,In_1143);
and U586 (N_586,In_494,In_1155);
or U587 (N_587,In_1379,In_1111);
nor U588 (N_588,In_536,In_645);
nand U589 (N_589,In_476,In_819);
nand U590 (N_590,In_1293,In_1023);
or U591 (N_591,In_81,In_926);
or U592 (N_592,In_130,In_1410);
nand U593 (N_593,In_76,In_746);
or U594 (N_594,In_1114,In_1497);
xnor U595 (N_595,In_71,In_263);
xnor U596 (N_596,In_246,In_808);
nor U597 (N_597,In_712,In_550);
or U598 (N_598,In_1438,In_684);
or U599 (N_599,In_1479,In_501);
and U600 (N_600,In_387,In_942);
nor U601 (N_601,In_1116,In_672);
and U602 (N_602,In_1069,In_25);
and U603 (N_603,In_1211,In_1045);
or U604 (N_604,In_570,In_243);
and U605 (N_605,In_864,In_561);
nand U606 (N_606,In_1294,In_324);
nor U607 (N_607,In_1094,In_935);
nand U608 (N_608,In_1325,In_617);
nor U609 (N_609,In_512,In_1310);
nand U610 (N_610,In_416,In_223);
or U611 (N_611,In_412,In_123);
nand U612 (N_612,In_194,In_754);
nand U613 (N_613,In_576,In_133);
xnor U614 (N_614,In_473,In_300);
xnor U615 (N_615,In_427,In_138);
or U616 (N_616,In_796,In_980);
nand U617 (N_617,In_312,In_1493);
and U618 (N_618,In_448,In_657);
and U619 (N_619,In_836,In_115);
nor U620 (N_620,In_1014,In_106);
xor U621 (N_621,In_874,In_965);
nor U622 (N_622,In_202,In_1411);
xor U623 (N_623,In_1255,In_1474);
nor U624 (N_624,In_1131,In_434);
nand U625 (N_625,In_631,In_872);
nor U626 (N_626,In_738,In_1220);
nor U627 (N_627,In_623,In_696);
or U628 (N_628,In_760,In_1440);
nand U629 (N_629,In_170,In_971);
nand U630 (N_630,In_556,In_1217);
or U631 (N_631,In_823,In_179);
xnor U632 (N_632,In_1182,In_1174);
and U633 (N_633,In_16,In_1098);
nand U634 (N_634,In_1039,In_762);
and U635 (N_635,In_307,In_184);
or U636 (N_636,In_1029,In_1342);
or U637 (N_637,In_993,In_1437);
and U638 (N_638,In_1200,In_424);
nor U639 (N_639,In_423,In_982);
and U640 (N_640,In_1080,In_834);
or U641 (N_641,In_867,In_216);
nand U642 (N_642,In_691,In_358);
nor U643 (N_643,In_1267,In_702);
or U644 (N_644,In_152,In_465);
and U645 (N_645,In_1317,In_959);
nand U646 (N_646,In_569,In_1041);
or U647 (N_647,In_770,In_46);
nor U648 (N_648,In_921,In_110);
nand U649 (N_649,In_1388,In_1146);
nor U650 (N_650,In_167,In_1011);
and U651 (N_651,In_385,In_638);
or U652 (N_652,In_375,In_518);
nor U653 (N_653,In_159,In_697);
or U654 (N_654,In_32,In_900);
nand U655 (N_655,In_655,In_1225);
or U656 (N_656,In_764,In_939);
nand U657 (N_657,In_1129,In_308);
and U658 (N_658,In_235,In_51);
or U659 (N_659,In_1276,In_1249);
or U660 (N_660,In_683,In_1340);
nand U661 (N_661,In_1082,In_22);
and U662 (N_662,In_222,In_1419);
and U663 (N_663,In_441,In_274);
and U664 (N_664,In_185,In_1374);
and U665 (N_665,In_1115,In_986);
nor U666 (N_666,In_748,In_329);
and U667 (N_667,In_1322,In_1101);
nor U668 (N_668,In_229,In_1250);
nor U669 (N_669,In_242,In_411);
nand U670 (N_670,In_871,In_1192);
nor U671 (N_671,In_551,In_824);
xor U672 (N_672,In_967,In_1140);
nand U673 (N_673,In_983,In_634);
and U674 (N_674,In_1005,In_988);
nor U675 (N_675,In_595,In_730);
and U676 (N_676,In_1286,In_1377);
or U677 (N_677,In_365,In_1231);
or U678 (N_678,In_306,In_750);
nand U679 (N_679,In_189,In_310);
or U680 (N_680,In_607,In_293);
nor U681 (N_681,In_1047,In_701);
and U682 (N_682,In_1219,In_269);
or U683 (N_683,In_710,In_859);
or U684 (N_684,In_118,In_49);
nand U685 (N_685,In_453,In_372);
and U686 (N_686,In_1130,In_822);
nor U687 (N_687,In_67,In_1466);
and U688 (N_688,In_1071,In_776);
or U689 (N_689,In_890,In_492);
and U690 (N_690,In_682,In_48);
nand U691 (N_691,In_815,In_44);
nand U692 (N_692,In_1378,In_1210);
nand U693 (N_693,In_826,In_718);
nor U694 (N_694,In_1368,In_347);
xor U695 (N_695,In_841,In_88);
or U696 (N_696,In_950,In_52);
nand U697 (N_697,In_273,In_990);
xor U698 (N_698,In_1133,In_1035);
and U699 (N_699,In_1086,In_452);
nand U700 (N_700,In_1004,In_1464);
and U701 (N_701,In_724,In_232);
nand U702 (N_702,In_1357,In_1223);
nand U703 (N_703,In_719,In_1312);
and U704 (N_704,In_58,In_177);
or U705 (N_705,In_572,In_237);
and U706 (N_706,In_850,In_870);
and U707 (N_707,In_614,In_1343);
xnor U708 (N_708,In_109,In_804);
and U709 (N_709,In_462,In_1346);
or U710 (N_710,In_1353,In_464);
or U711 (N_711,In_541,In_979);
nand U712 (N_712,In_1186,In_334);
nor U713 (N_713,In_396,In_924);
and U714 (N_714,In_875,In_401);
and U715 (N_715,In_930,In_1380);
nand U716 (N_716,In_30,In_1048);
and U717 (N_717,In_1179,In_721);
or U718 (N_718,In_500,In_9);
nor U719 (N_719,In_400,In_113);
nor U720 (N_720,In_1361,In_622);
and U721 (N_721,In_689,In_1083);
or U722 (N_722,In_854,In_849);
or U723 (N_723,In_581,In_1066);
nor U724 (N_724,In_1204,In_985);
or U725 (N_725,In_621,In_1233);
nand U726 (N_726,In_786,In_186);
and U727 (N_727,In_586,In_204);
nand U728 (N_728,In_676,In_104);
and U729 (N_729,In_41,In_878);
nor U730 (N_730,In_552,In_1487);
nor U731 (N_731,In_1327,In_954);
nor U732 (N_732,In_349,In_1196);
nor U733 (N_733,In_936,In_1258);
nor U734 (N_734,In_1395,In_663);
and U735 (N_735,In_404,In_1020);
or U736 (N_736,In_31,In_960);
xor U737 (N_737,In_975,In_976);
nor U738 (N_738,In_842,In_331);
and U739 (N_739,In_226,In_370);
xor U740 (N_740,In_1160,In_284);
or U741 (N_741,In_897,In_1073);
xnor U742 (N_742,In_1414,In_792);
nand U743 (N_743,In_562,In_429);
and U744 (N_744,In_34,In_868);
xor U745 (N_745,In_1138,In_156);
and U746 (N_746,In_679,In_1119);
and U747 (N_747,In_1008,In_913);
nand U748 (N_748,In_1480,In_64);
nand U749 (N_749,In_1399,In_1315);
nor U750 (N_750,N_665,N_372);
xor U751 (N_751,N_87,N_607);
nand U752 (N_752,N_582,N_219);
nor U753 (N_753,N_42,N_37);
or U754 (N_754,N_73,N_2);
or U755 (N_755,N_100,N_405);
or U756 (N_756,N_355,N_214);
and U757 (N_757,N_555,N_378);
or U758 (N_758,N_367,N_552);
and U759 (N_759,N_174,N_554);
nor U760 (N_760,N_308,N_616);
nand U761 (N_761,N_589,N_318);
nand U762 (N_762,N_585,N_510);
or U763 (N_763,N_29,N_319);
and U764 (N_764,N_579,N_720);
or U765 (N_765,N_606,N_639);
or U766 (N_766,N_627,N_519);
or U767 (N_767,N_124,N_374);
and U768 (N_768,N_584,N_691);
nor U769 (N_769,N_343,N_697);
nand U770 (N_770,N_310,N_186);
or U771 (N_771,N_126,N_497);
nor U772 (N_772,N_89,N_22);
nor U773 (N_773,N_24,N_201);
nand U774 (N_774,N_479,N_229);
or U775 (N_775,N_409,N_12);
nor U776 (N_776,N_134,N_425);
nor U777 (N_777,N_599,N_439);
xor U778 (N_778,N_400,N_713);
or U779 (N_779,N_456,N_94);
nand U780 (N_780,N_162,N_339);
or U781 (N_781,N_385,N_362);
nand U782 (N_782,N_568,N_569);
nor U783 (N_783,N_347,N_705);
and U784 (N_784,N_43,N_323);
or U785 (N_785,N_447,N_36);
or U786 (N_786,N_641,N_517);
nand U787 (N_787,N_596,N_509);
or U788 (N_788,N_441,N_290);
nand U789 (N_789,N_445,N_361);
or U790 (N_790,N_390,N_149);
nor U791 (N_791,N_233,N_131);
or U792 (N_792,N_285,N_560);
nand U793 (N_793,N_593,N_438);
nand U794 (N_794,N_139,N_413);
or U795 (N_795,N_414,N_474);
nand U796 (N_796,N_740,N_255);
nor U797 (N_797,N_199,N_230);
nand U798 (N_798,N_289,N_288);
nand U799 (N_799,N_156,N_685);
xnor U800 (N_800,N_222,N_693);
and U801 (N_801,N_689,N_631);
and U802 (N_802,N_518,N_386);
xor U803 (N_803,N_198,N_603);
and U804 (N_804,N_734,N_181);
nor U805 (N_805,N_403,N_442);
and U806 (N_806,N_745,N_562);
or U807 (N_807,N_648,N_63);
or U808 (N_808,N_31,N_59);
or U809 (N_809,N_415,N_292);
nand U810 (N_810,N_663,N_3);
nand U811 (N_811,N_541,N_498);
or U812 (N_812,N_215,N_695);
or U813 (N_813,N_244,N_264);
nand U814 (N_814,N_530,N_180);
nand U815 (N_815,N_428,N_184);
nand U816 (N_816,N_591,N_117);
nand U817 (N_817,N_528,N_628);
or U818 (N_818,N_283,N_743);
and U819 (N_819,N_505,N_209);
or U820 (N_820,N_249,N_470);
or U821 (N_821,N_331,N_389);
nand U822 (N_822,N_95,N_500);
nor U823 (N_823,N_398,N_563);
or U824 (N_824,N_306,N_575);
nand U825 (N_825,N_392,N_657);
nor U826 (N_826,N_189,N_618);
nand U827 (N_827,N_39,N_128);
nand U828 (N_828,N_161,N_449);
nand U829 (N_829,N_56,N_330);
or U830 (N_830,N_267,N_531);
xnor U831 (N_831,N_246,N_614);
and U832 (N_832,N_130,N_9);
or U833 (N_833,N_658,N_512);
nand U834 (N_834,N_223,N_363);
xor U835 (N_835,N_687,N_513);
nor U836 (N_836,N_723,N_231);
and U837 (N_837,N_666,N_507);
nand U838 (N_838,N_268,N_598);
or U839 (N_839,N_110,N_276);
or U840 (N_840,N_340,N_625);
and U841 (N_841,N_459,N_178);
and U842 (N_842,N_206,N_580);
nand U843 (N_843,N_356,N_321);
nor U844 (N_844,N_305,N_698);
and U845 (N_845,N_662,N_160);
or U846 (N_846,N_26,N_27);
or U847 (N_847,N_113,N_481);
or U848 (N_848,N_699,N_342);
or U849 (N_849,N_696,N_67);
and U850 (N_850,N_349,N_74);
nand U851 (N_851,N_708,N_592);
nand U852 (N_852,N_679,N_643);
nor U853 (N_853,N_686,N_213);
or U854 (N_854,N_477,N_402);
xnor U855 (N_855,N_287,N_533);
or U856 (N_856,N_25,N_454);
nand U857 (N_857,N_433,N_434);
nor U858 (N_858,N_382,N_119);
and U859 (N_859,N_655,N_701);
nand U860 (N_860,N_647,N_550);
nand U861 (N_861,N_182,N_573);
nor U862 (N_862,N_391,N_738);
nor U863 (N_863,N_51,N_672);
or U864 (N_864,N_544,N_153);
nand U865 (N_865,N_86,N_604);
and U866 (N_866,N_116,N_265);
nand U867 (N_867,N_247,N_432);
xnor U868 (N_868,N_17,N_646);
nor U869 (N_869,N_300,N_379);
and U870 (N_870,N_45,N_144);
or U871 (N_871,N_193,N_190);
nor U872 (N_872,N_661,N_669);
nand U873 (N_873,N_320,N_532);
and U874 (N_874,N_270,N_727);
nand U875 (N_875,N_478,N_674);
or U876 (N_876,N_393,N_396);
or U877 (N_877,N_138,N_313);
nor U878 (N_878,N_387,N_350);
or U879 (N_879,N_96,N_633);
and U880 (N_880,N_47,N_601);
or U881 (N_881,N_261,N_348);
and U882 (N_882,N_577,N_424);
xnor U883 (N_883,N_203,N_325);
nand U884 (N_884,N_630,N_680);
or U885 (N_885,N_467,N_650);
nor U886 (N_886,N_324,N_397);
or U887 (N_887,N_238,N_380);
nand U888 (N_888,N_32,N_158);
nand U889 (N_889,N_430,N_163);
nor U890 (N_890,N_561,N_104);
and U891 (N_891,N_165,N_399);
nor U892 (N_892,N_511,N_464);
nor U893 (N_893,N_462,N_538);
nor U894 (N_894,N_337,N_351);
and U895 (N_895,N_105,N_60);
nand U896 (N_896,N_84,N_704);
xnor U897 (N_897,N_307,N_352);
and U898 (N_898,N_426,N_83);
nor U899 (N_899,N_613,N_458);
or U900 (N_900,N_711,N_252);
or U901 (N_901,N_44,N_677);
or U902 (N_902,N_684,N_502);
or U903 (N_903,N_133,N_151);
and U904 (N_904,N_617,N_717);
or U905 (N_905,N_480,N_702);
and U906 (N_906,N_277,N_654);
nor U907 (N_907,N_615,N_465);
and U908 (N_908,N_377,N_728);
nor U909 (N_909,N_317,N_642);
and U910 (N_910,N_749,N_383);
xor U911 (N_911,N_99,N_673);
and U912 (N_912,N_681,N_463);
and U913 (N_913,N_291,N_494);
nand U914 (N_914,N_543,N_521);
or U915 (N_915,N_72,N_653);
nor U916 (N_916,N_281,N_659);
or U917 (N_917,N_241,N_314);
and U918 (N_918,N_602,N_260);
nand U919 (N_919,N_49,N_54);
nand U920 (N_920,N_312,N_62);
nor U921 (N_921,N_173,N_731);
and U922 (N_922,N_644,N_394);
xnor U923 (N_923,N_217,N_545);
nor U924 (N_924,N_730,N_177);
nand U925 (N_925,N_301,N_197);
nor U926 (N_926,N_504,N_141);
nor U927 (N_927,N_417,N_472);
xor U928 (N_928,N_64,N_407);
nand U929 (N_929,N_81,N_656);
or U930 (N_930,N_537,N_612);
nand U931 (N_931,N_623,N_485);
nor U932 (N_932,N_91,N_475);
xor U933 (N_933,N_443,N_50);
nor U934 (N_934,N_735,N_609);
nand U935 (N_935,N_594,N_316);
xor U936 (N_936,N_132,N_28);
nand U937 (N_937,N_7,N_236);
and U938 (N_938,N_499,N_714);
and U939 (N_939,N_102,N_489);
nand U940 (N_940,N_376,N_5);
or U941 (N_941,N_92,N_712);
or U942 (N_942,N_106,N_540);
or U943 (N_943,N_707,N_329);
nor U944 (N_944,N_488,N_237);
nor U945 (N_945,N_457,N_58);
nand U946 (N_946,N_448,N_295);
and U947 (N_947,N_297,N_460);
nor U948 (N_948,N_228,N_640);
xor U949 (N_949,N_194,N_668);
and U950 (N_950,N_188,N_66);
nor U951 (N_951,N_737,N_221);
nor U952 (N_952,N_234,N_183);
nand U953 (N_953,N_38,N_423);
nor U954 (N_954,N_476,N_142);
nand U955 (N_955,N_46,N_278);
nor U956 (N_956,N_482,N_53);
nor U957 (N_957,N_484,N_595);
and U958 (N_958,N_280,N_311);
and U959 (N_959,N_610,N_581);
nor U960 (N_960,N_468,N_416);
or U961 (N_961,N_250,N_522);
and U962 (N_962,N_358,N_157);
xor U963 (N_963,N_514,N_729);
xnor U964 (N_964,N_109,N_61);
xnor U965 (N_965,N_200,N_210);
nand U966 (N_966,N_16,N_239);
nand U967 (N_967,N_303,N_76);
xor U968 (N_968,N_101,N_676);
nor U969 (N_969,N_263,N_664);
nor U970 (N_970,N_195,N_520);
nor U971 (N_971,N_539,N_700);
and U972 (N_972,N_21,N_240);
and U973 (N_973,N_401,N_251);
xnor U974 (N_974,N_286,N_258);
and U975 (N_975,N_167,N_486);
and U976 (N_976,N_586,N_282);
nor U977 (N_977,N_719,N_332);
and U978 (N_978,N_716,N_440);
and U979 (N_979,N_275,N_176);
nor U980 (N_980,N_638,N_97);
and U981 (N_981,N_140,N_490);
xor U982 (N_982,N_15,N_619);
nor U983 (N_983,N_567,N_410);
nand U984 (N_984,N_166,N_469);
and U985 (N_985,N_108,N_18);
nand U986 (N_986,N_322,N_262);
and U987 (N_987,N_304,N_451);
and U988 (N_988,N_148,N_4);
or U989 (N_989,N_115,N_559);
and U990 (N_990,N_726,N_473);
and U991 (N_991,N_395,N_205);
nand U992 (N_992,N_272,N_8);
nor U993 (N_993,N_651,N_578);
nor U994 (N_994,N_245,N_649);
or U995 (N_995,N_344,N_253);
and U996 (N_996,N_80,N_373);
nor U997 (N_997,N_254,N_65);
or U998 (N_998,N_576,N_381);
or U999 (N_999,N_293,N_690);
nor U1000 (N_1000,N_436,N_721);
or U1001 (N_1001,N_274,N_146);
or U1002 (N_1002,N_493,N_6);
or U1003 (N_1003,N_341,N_626);
nor U1004 (N_1004,N_412,N_123);
or U1005 (N_1005,N_23,N_572);
nor U1006 (N_1006,N_435,N_127);
and U1007 (N_1007,N_529,N_327);
nor U1008 (N_1008,N_526,N_137);
and U1009 (N_1009,N_709,N_667);
nand U1010 (N_1010,N_112,N_365);
nand U1011 (N_1011,N_742,N_556);
or U1012 (N_1012,N_629,N_558);
or U1013 (N_1013,N_52,N_79);
nor U1014 (N_1014,N_411,N_227);
and U1015 (N_1015,N_455,N_1);
or U1016 (N_1016,N_77,N_524);
and U1017 (N_1017,N_170,N_688);
nand U1018 (N_1018,N_55,N_40);
nor U1019 (N_1019,N_491,N_35);
or U1020 (N_1020,N_159,N_645);
nand U1021 (N_1021,N_143,N_620);
and U1022 (N_1022,N_431,N_164);
and U1023 (N_1023,N_418,N_527);
nand U1024 (N_1024,N_334,N_279);
nand U1025 (N_1025,N_453,N_471);
and U1026 (N_1026,N_444,N_694);
nor U1027 (N_1027,N_671,N_747);
nand U1028 (N_1028,N_273,N_624);
and U1029 (N_1029,N_706,N_501);
nor U1030 (N_1030,N_145,N_450);
or U1031 (N_1031,N_506,N_13);
and U1032 (N_1032,N_670,N_461);
and U1033 (N_1033,N_406,N_375);
nand U1034 (N_1034,N_359,N_225);
xor U1035 (N_1035,N_574,N_336);
and U1036 (N_1036,N_269,N_683);
nand U1037 (N_1037,N_78,N_243);
or U1038 (N_1038,N_736,N_384);
nor U1039 (N_1039,N_611,N_335);
and U1040 (N_1040,N_404,N_364);
nand U1041 (N_1041,N_187,N_408);
xnor U1042 (N_1042,N_710,N_637);
xnor U1043 (N_1043,N_583,N_284);
or U1044 (N_1044,N_366,N_175);
nor U1045 (N_1045,N_370,N_715);
nor U1046 (N_1046,N_114,N_536);
or U1047 (N_1047,N_271,N_678);
and U1048 (N_1048,N_692,N_120);
nor U1049 (N_1049,N_82,N_388);
or U1050 (N_1050,N_420,N_535);
or U1051 (N_1051,N_309,N_600);
nand U1052 (N_1052,N_547,N_542);
nor U1053 (N_1053,N_732,N_452);
nor U1054 (N_1054,N_48,N_212);
or U1055 (N_1055,N_549,N_622);
and U1056 (N_1056,N_523,N_179);
xor U1057 (N_1057,N_147,N_360);
nor U1058 (N_1058,N_93,N_571);
nand U1059 (N_1059,N_733,N_196);
nor U1060 (N_1060,N_294,N_525);
xnor U1061 (N_1061,N_437,N_608);
nor U1062 (N_1062,N_224,N_70);
and U1063 (N_1063,N_226,N_590);
nor U1064 (N_1064,N_11,N_33);
nor U1065 (N_1065,N_636,N_660);
nand U1066 (N_1066,N_111,N_635);
and U1067 (N_1067,N_218,N_487);
nand U1068 (N_1068,N_90,N_328);
nand U1069 (N_1069,N_354,N_632);
and U1070 (N_1070,N_429,N_257);
or U1071 (N_1071,N_588,N_368);
or U1072 (N_1072,N_19,N_152);
and U1073 (N_1073,N_171,N_202);
nor U1074 (N_1074,N_98,N_155);
nor U1075 (N_1075,N_725,N_516);
or U1076 (N_1076,N_150,N_204);
or U1077 (N_1077,N_621,N_242);
and U1078 (N_1078,N_515,N_0);
xnor U1079 (N_1079,N_496,N_71);
and U1080 (N_1080,N_718,N_724);
or U1081 (N_1081,N_168,N_207);
and U1082 (N_1082,N_605,N_192);
nand U1083 (N_1083,N_353,N_125);
or U1084 (N_1084,N_682,N_118);
or U1085 (N_1085,N_357,N_346);
nor U1086 (N_1086,N_211,N_326);
nor U1087 (N_1087,N_333,N_256);
or U1088 (N_1088,N_741,N_68);
and U1089 (N_1089,N_597,N_508);
nor U1090 (N_1090,N_169,N_546);
nor U1091 (N_1091,N_57,N_299);
and U1092 (N_1092,N_20,N_587);
or U1093 (N_1093,N_103,N_744);
nor U1094 (N_1094,N_302,N_557);
or U1095 (N_1095,N_566,N_534);
and U1096 (N_1096,N_248,N_30);
nand U1097 (N_1097,N_739,N_652);
nor U1098 (N_1098,N_136,N_266);
nor U1099 (N_1099,N_565,N_232);
and U1100 (N_1100,N_553,N_570);
nand U1101 (N_1101,N_722,N_220);
nor U1102 (N_1102,N_122,N_495);
or U1103 (N_1103,N_492,N_172);
and U1104 (N_1104,N_634,N_421);
and U1105 (N_1105,N_129,N_746);
and U1106 (N_1106,N_422,N_446);
nand U1107 (N_1107,N_69,N_564);
nor U1108 (N_1108,N_296,N_235);
and U1109 (N_1109,N_675,N_185);
nand U1110 (N_1110,N_338,N_191);
nor U1111 (N_1111,N_88,N_107);
nor U1112 (N_1112,N_345,N_208);
and U1113 (N_1113,N_315,N_483);
nor U1114 (N_1114,N_551,N_85);
or U1115 (N_1115,N_419,N_748);
or U1116 (N_1116,N_41,N_34);
nand U1117 (N_1117,N_548,N_216);
nand U1118 (N_1118,N_503,N_371);
nand U1119 (N_1119,N_466,N_14);
or U1120 (N_1120,N_703,N_427);
nand U1121 (N_1121,N_259,N_298);
xnor U1122 (N_1122,N_10,N_369);
or U1123 (N_1123,N_135,N_75);
nor U1124 (N_1124,N_154,N_121);
nor U1125 (N_1125,N_173,N_122);
or U1126 (N_1126,N_435,N_558);
or U1127 (N_1127,N_551,N_35);
and U1128 (N_1128,N_434,N_366);
nor U1129 (N_1129,N_58,N_497);
or U1130 (N_1130,N_292,N_557);
or U1131 (N_1131,N_324,N_700);
or U1132 (N_1132,N_7,N_443);
or U1133 (N_1133,N_430,N_261);
nor U1134 (N_1134,N_299,N_117);
nor U1135 (N_1135,N_402,N_37);
xnor U1136 (N_1136,N_189,N_131);
and U1137 (N_1137,N_25,N_367);
xor U1138 (N_1138,N_497,N_742);
nand U1139 (N_1139,N_560,N_496);
nor U1140 (N_1140,N_604,N_548);
nor U1141 (N_1141,N_513,N_312);
nor U1142 (N_1142,N_606,N_356);
or U1143 (N_1143,N_27,N_543);
nor U1144 (N_1144,N_324,N_2);
xor U1145 (N_1145,N_661,N_80);
and U1146 (N_1146,N_25,N_348);
nor U1147 (N_1147,N_745,N_237);
xnor U1148 (N_1148,N_511,N_387);
nor U1149 (N_1149,N_376,N_452);
nand U1150 (N_1150,N_205,N_738);
or U1151 (N_1151,N_667,N_503);
nand U1152 (N_1152,N_117,N_107);
or U1153 (N_1153,N_446,N_163);
nand U1154 (N_1154,N_355,N_642);
and U1155 (N_1155,N_152,N_14);
or U1156 (N_1156,N_120,N_163);
and U1157 (N_1157,N_228,N_414);
xnor U1158 (N_1158,N_405,N_152);
or U1159 (N_1159,N_435,N_429);
and U1160 (N_1160,N_35,N_284);
nand U1161 (N_1161,N_601,N_425);
or U1162 (N_1162,N_249,N_224);
nor U1163 (N_1163,N_653,N_106);
and U1164 (N_1164,N_114,N_517);
nand U1165 (N_1165,N_325,N_419);
nor U1166 (N_1166,N_672,N_424);
nand U1167 (N_1167,N_576,N_336);
and U1168 (N_1168,N_352,N_480);
nand U1169 (N_1169,N_543,N_492);
and U1170 (N_1170,N_55,N_64);
or U1171 (N_1171,N_405,N_496);
or U1172 (N_1172,N_509,N_554);
nand U1173 (N_1173,N_262,N_385);
or U1174 (N_1174,N_476,N_624);
nor U1175 (N_1175,N_545,N_129);
nand U1176 (N_1176,N_569,N_83);
or U1177 (N_1177,N_509,N_599);
and U1178 (N_1178,N_312,N_624);
and U1179 (N_1179,N_327,N_15);
and U1180 (N_1180,N_7,N_5);
nand U1181 (N_1181,N_152,N_700);
nand U1182 (N_1182,N_172,N_331);
or U1183 (N_1183,N_607,N_618);
nor U1184 (N_1184,N_134,N_412);
or U1185 (N_1185,N_125,N_344);
or U1186 (N_1186,N_688,N_732);
nor U1187 (N_1187,N_186,N_324);
or U1188 (N_1188,N_620,N_705);
or U1189 (N_1189,N_430,N_368);
nor U1190 (N_1190,N_503,N_507);
or U1191 (N_1191,N_39,N_203);
or U1192 (N_1192,N_155,N_342);
or U1193 (N_1193,N_491,N_149);
xnor U1194 (N_1194,N_396,N_146);
and U1195 (N_1195,N_480,N_363);
and U1196 (N_1196,N_471,N_480);
nor U1197 (N_1197,N_159,N_732);
or U1198 (N_1198,N_603,N_717);
or U1199 (N_1199,N_7,N_165);
or U1200 (N_1200,N_75,N_85);
nand U1201 (N_1201,N_560,N_420);
xor U1202 (N_1202,N_644,N_278);
nor U1203 (N_1203,N_137,N_34);
nand U1204 (N_1204,N_236,N_157);
or U1205 (N_1205,N_218,N_709);
nor U1206 (N_1206,N_516,N_196);
xor U1207 (N_1207,N_197,N_562);
nor U1208 (N_1208,N_393,N_504);
nor U1209 (N_1209,N_359,N_462);
and U1210 (N_1210,N_49,N_602);
nand U1211 (N_1211,N_455,N_426);
nand U1212 (N_1212,N_496,N_235);
or U1213 (N_1213,N_270,N_84);
nand U1214 (N_1214,N_179,N_666);
nand U1215 (N_1215,N_667,N_245);
xor U1216 (N_1216,N_441,N_523);
and U1217 (N_1217,N_575,N_512);
nand U1218 (N_1218,N_93,N_632);
nor U1219 (N_1219,N_409,N_616);
nand U1220 (N_1220,N_746,N_119);
or U1221 (N_1221,N_436,N_143);
and U1222 (N_1222,N_657,N_708);
nand U1223 (N_1223,N_342,N_174);
nor U1224 (N_1224,N_504,N_82);
and U1225 (N_1225,N_547,N_273);
or U1226 (N_1226,N_329,N_485);
or U1227 (N_1227,N_588,N_620);
and U1228 (N_1228,N_583,N_645);
or U1229 (N_1229,N_224,N_76);
and U1230 (N_1230,N_678,N_528);
nand U1231 (N_1231,N_588,N_337);
nand U1232 (N_1232,N_430,N_363);
and U1233 (N_1233,N_408,N_381);
or U1234 (N_1234,N_471,N_196);
nand U1235 (N_1235,N_648,N_351);
nand U1236 (N_1236,N_211,N_185);
and U1237 (N_1237,N_651,N_291);
nand U1238 (N_1238,N_529,N_649);
and U1239 (N_1239,N_697,N_628);
or U1240 (N_1240,N_483,N_631);
and U1241 (N_1241,N_83,N_367);
or U1242 (N_1242,N_106,N_682);
xor U1243 (N_1243,N_284,N_607);
or U1244 (N_1244,N_274,N_616);
nor U1245 (N_1245,N_292,N_567);
or U1246 (N_1246,N_241,N_109);
nand U1247 (N_1247,N_15,N_590);
nand U1248 (N_1248,N_632,N_502);
nor U1249 (N_1249,N_377,N_575);
xor U1250 (N_1250,N_112,N_606);
or U1251 (N_1251,N_319,N_733);
nand U1252 (N_1252,N_195,N_716);
or U1253 (N_1253,N_521,N_488);
or U1254 (N_1254,N_125,N_220);
nor U1255 (N_1255,N_493,N_405);
nand U1256 (N_1256,N_585,N_79);
and U1257 (N_1257,N_250,N_691);
or U1258 (N_1258,N_37,N_554);
nand U1259 (N_1259,N_671,N_317);
or U1260 (N_1260,N_483,N_392);
and U1261 (N_1261,N_566,N_263);
or U1262 (N_1262,N_204,N_129);
and U1263 (N_1263,N_711,N_18);
xnor U1264 (N_1264,N_665,N_506);
xnor U1265 (N_1265,N_43,N_118);
nand U1266 (N_1266,N_166,N_283);
and U1267 (N_1267,N_719,N_247);
nand U1268 (N_1268,N_608,N_284);
xor U1269 (N_1269,N_568,N_504);
or U1270 (N_1270,N_131,N_641);
nand U1271 (N_1271,N_82,N_404);
and U1272 (N_1272,N_625,N_284);
and U1273 (N_1273,N_506,N_593);
nor U1274 (N_1274,N_190,N_277);
nand U1275 (N_1275,N_553,N_41);
xnor U1276 (N_1276,N_377,N_744);
and U1277 (N_1277,N_564,N_259);
xor U1278 (N_1278,N_684,N_490);
nand U1279 (N_1279,N_194,N_613);
nor U1280 (N_1280,N_634,N_646);
nor U1281 (N_1281,N_228,N_266);
nand U1282 (N_1282,N_269,N_414);
nor U1283 (N_1283,N_516,N_230);
xnor U1284 (N_1284,N_55,N_700);
nand U1285 (N_1285,N_80,N_286);
nand U1286 (N_1286,N_345,N_138);
or U1287 (N_1287,N_264,N_470);
and U1288 (N_1288,N_666,N_366);
nand U1289 (N_1289,N_712,N_542);
and U1290 (N_1290,N_78,N_614);
and U1291 (N_1291,N_707,N_599);
and U1292 (N_1292,N_445,N_6);
or U1293 (N_1293,N_398,N_408);
nor U1294 (N_1294,N_201,N_82);
nand U1295 (N_1295,N_551,N_597);
nor U1296 (N_1296,N_302,N_389);
and U1297 (N_1297,N_216,N_664);
or U1298 (N_1298,N_504,N_417);
nor U1299 (N_1299,N_169,N_403);
and U1300 (N_1300,N_576,N_747);
nor U1301 (N_1301,N_740,N_634);
nor U1302 (N_1302,N_88,N_153);
xnor U1303 (N_1303,N_394,N_519);
nor U1304 (N_1304,N_669,N_262);
and U1305 (N_1305,N_301,N_269);
nor U1306 (N_1306,N_738,N_282);
and U1307 (N_1307,N_586,N_420);
nor U1308 (N_1308,N_415,N_749);
and U1309 (N_1309,N_278,N_260);
nand U1310 (N_1310,N_134,N_218);
nor U1311 (N_1311,N_172,N_50);
or U1312 (N_1312,N_21,N_65);
or U1313 (N_1313,N_505,N_571);
or U1314 (N_1314,N_191,N_71);
nand U1315 (N_1315,N_188,N_216);
nand U1316 (N_1316,N_667,N_619);
nor U1317 (N_1317,N_298,N_145);
nor U1318 (N_1318,N_271,N_664);
nor U1319 (N_1319,N_325,N_440);
or U1320 (N_1320,N_318,N_407);
and U1321 (N_1321,N_466,N_28);
or U1322 (N_1322,N_561,N_537);
nand U1323 (N_1323,N_253,N_626);
nor U1324 (N_1324,N_23,N_132);
nand U1325 (N_1325,N_45,N_419);
and U1326 (N_1326,N_377,N_557);
and U1327 (N_1327,N_577,N_361);
nand U1328 (N_1328,N_671,N_342);
and U1329 (N_1329,N_734,N_414);
nand U1330 (N_1330,N_451,N_733);
nand U1331 (N_1331,N_77,N_624);
nand U1332 (N_1332,N_642,N_154);
nor U1333 (N_1333,N_276,N_289);
nand U1334 (N_1334,N_642,N_179);
and U1335 (N_1335,N_21,N_411);
nor U1336 (N_1336,N_556,N_585);
and U1337 (N_1337,N_301,N_612);
and U1338 (N_1338,N_268,N_290);
xor U1339 (N_1339,N_467,N_279);
nand U1340 (N_1340,N_13,N_658);
nor U1341 (N_1341,N_696,N_292);
and U1342 (N_1342,N_511,N_118);
nand U1343 (N_1343,N_491,N_187);
or U1344 (N_1344,N_683,N_159);
or U1345 (N_1345,N_647,N_717);
and U1346 (N_1346,N_414,N_432);
xor U1347 (N_1347,N_138,N_417);
xor U1348 (N_1348,N_249,N_449);
nand U1349 (N_1349,N_77,N_657);
and U1350 (N_1350,N_319,N_519);
or U1351 (N_1351,N_557,N_579);
or U1352 (N_1352,N_663,N_160);
or U1353 (N_1353,N_202,N_302);
or U1354 (N_1354,N_302,N_645);
and U1355 (N_1355,N_564,N_709);
and U1356 (N_1356,N_203,N_748);
xor U1357 (N_1357,N_196,N_192);
nand U1358 (N_1358,N_216,N_566);
and U1359 (N_1359,N_686,N_645);
or U1360 (N_1360,N_435,N_427);
nand U1361 (N_1361,N_120,N_478);
nand U1362 (N_1362,N_558,N_353);
and U1363 (N_1363,N_470,N_336);
nor U1364 (N_1364,N_256,N_562);
or U1365 (N_1365,N_245,N_359);
nor U1366 (N_1366,N_599,N_658);
and U1367 (N_1367,N_199,N_737);
and U1368 (N_1368,N_51,N_161);
nor U1369 (N_1369,N_518,N_401);
or U1370 (N_1370,N_553,N_467);
and U1371 (N_1371,N_98,N_708);
nor U1372 (N_1372,N_198,N_491);
or U1373 (N_1373,N_134,N_477);
and U1374 (N_1374,N_352,N_193);
xnor U1375 (N_1375,N_22,N_680);
nor U1376 (N_1376,N_152,N_608);
nor U1377 (N_1377,N_514,N_404);
and U1378 (N_1378,N_340,N_14);
or U1379 (N_1379,N_90,N_505);
and U1380 (N_1380,N_163,N_694);
nand U1381 (N_1381,N_255,N_744);
or U1382 (N_1382,N_38,N_81);
and U1383 (N_1383,N_636,N_350);
or U1384 (N_1384,N_231,N_184);
or U1385 (N_1385,N_737,N_735);
nand U1386 (N_1386,N_177,N_53);
or U1387 (N_1387,N_484,N_5);
and U1388 (N_1388,N_665,N_358);
nor U1389 (N_1389,N_343,N_678);
nor U1390 (N_1390,N_133,N_181);
or U1391 (N_1391,N_185,N_303);
and U1392 (N_1392,N_229,N_512);
nor U1393 (N_1393,N_444,N_485);
nand U1394 (N_1394,N_229,N_366);
nor U1395 (N_1395,N_337,N_690);
nand U1396 (N_1396,N_41,N_141);
and U1397 (N_1397,N_544,N_637);
nand U1398 (N_1398,N_447,N_553);
and U1399 (N_1399,N_485,N_218);
nand U1400 (N_1400,N_652,N_23);
nand U1401 (N_1401,N_567,N_713);
nor U1402 (N_1402,N_351,N_617);
or U1403 (N_1403,N_514,N_109);
and U1404 (N_1404,N_181,N_322);
or U1405 (N_1405,N_418,N_471);
xnor U1406 (N_1406,N_176,N_710);
nand U1407 (N_1407,N_73,N_241);
nor U1408 (N_1408,N_84,N_511);
or U1409 (N_1409,N_100,N_157);
or U1410 (N_1410,N_262,N_423);
xnor U1411 (N_1411,N_160,N_624);
or U1412 (N_1412,N_307,N_386);
xor U1413 (N_1413,N_675,N_121);
xor U1414 (N_1414,N_276,N_290);
nor U1415 (N_1415,N_241,N_573);
and U1416 (N_1416,N_692,N_43);
nand U1417 (N_1417,N_69,N_734);
nor U1418 (N_1418,N_603,N_327);
nand U1419 (N_1419,N_14,N_739);
and U1420 (N_1420,N_238,N_370);
or U1421 (N_1421,N_245,N_515);
xor U1422 (N_1422,N_65,N_201);
nand U1423 (N_1423,N_290,N_603);
and U1424 (N_1424,N_536,N_388);
nand U1425 (N_1425,N_647,N_173);
nor U1426 (N_1426,N_694,N_305);
nor U1427 (N_1427,N_149,N_699);
and U1428 (N_1428,N_557,N_39);
nor U1429 (N_1429,N_412,N_582);
and U1430 (N_1430,N_124,N_541);
or U1431 (N_1431,N_38,N_132);
xor U1432 (N_1432,N_168,N_71);
and U1433 (N_1433,N_595,N_223);
nor U1434 (N_1434,N_311,N_497);
and U1435 (N_1435,N_21,N_51);
or U1436 (N_1436,N_591,N_461);
or U1437 (N_1437,N_189,N_393);
or U1438 (N_1438,N_163,N_550);
nand U1439 (N_1439,N_623,N_115);
nand U1440 (N_1440,N_635,N_140);
nand U1441 (N_1441,N_403,N_250);
nor U1442 (N_1442,N_748,N_357);
nand U1443 (N_1443,N_76,N_28);
and U1444 (N_1444,N_542,N_623);
nor U1445 (N_1445,N_307,N_581);
or U1446 (N_1446,N_633,N_247);
nor U1447 (N_1447,N_354,N_41);
and U1448 (N_1448,N_747,N_426);
or U1449 (N_1449,N_31,N_665);
or U1450 (N_1450,N_556,N_480);
nor U1451 (N_1451,N_675,N_408);
or U1452 (N_1452,N_399,N_246);
nand U1453 (N_1453,N_577,N_395);
nand U1454 (N_1454,N_595,N_747);
nand U1455 (N_1455,N_580,N_384);
and U1456 (N_1456,N_464,N_411);
or U1457 (N_1457,N_678,N_616);
nand U1458 (N_1458,N_494,N_369);
or U1459 (N_1459,N_654,N_656);
nor U1460 (N_1460,N_329,N_226);
nand U1461 (N_1461,N_563,N_646);
nand U1462 (N_1462,N_675,N_106);
nand U1463 (N_1463,N_338,N_478);
nand U1464 (N_1464,N_108,N_200);
and U1465 (N_1465,N_522,N_229);
nor U1466 (N_1466,N_90,N_281);
nand U1467 (N_1467,N_13,N_708);
xnor U1468 (N_1468,N_223,N_736);
nand U1469 (N_1469,N_29,N_172);
nand U1470 (N_1470,N_691,N_700);
nor U1471 (N_1471,N_602,N_579);
nand U1472 (N_1472,N_335,N_193);
or U1473 (N_1473,N_396,N_375);
xor U1474 (N_1474,N_647,N_401);
xnor U1475 (N_1475,N_172,N_416);
or U1476 (N_1476,N_310,N_274);
xor U1477 (N_1477,N_134,N_468);
xor U1478 (N_1478,N_103,N_18);
nor U1479 (N_1479,N_349,N_616);
nand U1480 (N_1480,N_156,N_333);
nand U1481 (N_1481,N_107,N_349);
nand U1482 (N_1482,N_475,N_520);
nand U1483 (N_1483,N_164,N_17);
or U1484 (N_1484,N_629,N_271);
nand U1485 (N_1485,N_687,N_549);
or U1486 (N_1486,N_152,N_533);
nor U1487 (N_1487,N_143,N_470);
or U1488 (N_1488,N_45,N_70);
and U1489 (N_1489,N_206,N_62);
xor U1490 (N_1490,N_53,N_733);
and U1491 (N_1491,N_488,N_297);
xor U1492 (N_1492,N_249,N_28);
or U1493 (N_1493,N_43,N_557);
nor U1494 (N_1494,N_383,N_158);
and U1495 (N_1495,N_110,N_239);
and U1496 (N_1496,N_670,N_138);
nor U1497 (N_1497,N_717,N_725);
or U1498 (N_1498,N_197,N_618);
and U1499 (N_1499,N_352,N_737);
nand U1500 (N_1500,N_1219,N_1056);
xnor U1501 (N_1501,N_1498,N_1216);
or U1502 (N_1502,N_806,N_1112);
nand U1503 (N_1503,N_905,N_1097);
and U1504 (N_1504,N_1207,N_1188);
nor U1505 (N_1505,N_1284,N_991);
nor U1506 (N_1506,N_1131,N_1159);
nand U1507 (N_1507,N_956,N_1302);
nor U1508 (N_1508,N_960,N_930);
and U1509 (N_1509,N_1166,N_1205);
or U1510 (N_1510,N_1297,N_1433);
nand U1511 (N_1511,N_1497,N_768);
nor U1512 (N_1512,N_1173,N_1103);
nand U1513 (N_1513,N_1094,N_853);
or U1514 (N_1514,N_1061,N_984);
and U1515 (N_1515,N_1352,N_1336);
nor U1516 (N_1516,N_1037,N_1024);
or U1517 (N_1517,N_1314,N_1218);
nand U1518 (N_1518,N_938,N_1235);
nor U1519 (N_1519,N_1398,N_1105);
nor U1520 (N_1520,N_1451,N_1099);
or U1521 (N_1521,N_1100,N_1458);
nor U1522 (N_1522,N_1281,N_1265);
nor U1523 (N_1523,N_898,N_830);
nand U1524 (N_1524,N_940,N_1138);
xnor U1525 (N_1525,N_1347,N_921);
nand U1526 (N_1526,N_992,N_1456);
nor U1527 (N_1527,N_1483,N_873);
nor U1528 (N_1528,N_1454,N_1298);
and U1529 (N_1529,N_883,N_1035);
and U1530 (N_1530,N_1135,N_1369);
nor U1531 (N_1531,N_1424,N_1434);
nor U1532 (N_1532,N_1272,N_1130);
or U1533 (N_1533,N_1109,N_807);
xnor U1534 (N_1534,N_1200,N_786);
nand U1535 (N_1535,N_1279,N_790);
or U1536 (N_1536,N_1170,N_841);
and U1537 (N_1537,N_875,N_810);
or U1538 (N_1538,N_911,N_1041);
or U1539 (N_1539,N_1441,N_772);
and U1540 (N_1540,N_1491,N_1315);
or U1541 (N_1541,N_1139,N_843);
nor U1542 (N_1542,N_1176,N_804);
nand U1543 (N_1543,N_1348,N_1078);
nand U1544 (N_1544,N_1006,N_922);
nor U1545 (N_1545,N_1289,N_1419);
or U1546 (N_1546,N_1335,N_935);
nor U1547 (N_1547,N_978,N_754);
nor U1548 (N_1548,N_1417,N_1102);
or U1549 (N_1549,N_1285,N_1113);
nand U1550 (N_1550,N_1384,N_1212);
or U1551 (N_1551,N_1372,N_840);
nand U1552 (N_1552,N_1440,N_1310);
or U1553 (N_1553,N_864,N_1088);
xnor U1554 (N_1554,N_762,N_881);
nand U1555 (N_1555,N_1196,N_1146);
nand U1556 (N_1556,N_1343,N_782);
nand U1557 (N_1557,N_1472,N_958);
nor U1558 (N_1558,N_1154,N_1082);
nor U1559 (N_1559,N_1333,N_1437);
and U1560 (N_1560,N_990,N_1363);
xnor U1561 (N_1561,N_1072,N_1390);
or U1562 (N_1562,N_1052,N_1098);
and U1563 (N_1563,N_1358,N_1446);
nor U1564 (N_1564,N_886,N_847);
and U1565 (N_1565,N_1340,N_1048);
or U1566 (N_1566,N_818,N_966);
xor U1567 (N_1567,N_1476,N_1237);
nor U1568 (N_1568,N_1420,N_904);
nand U1569 (N_1569,N_986,N_1484);
and U1570 (N_1570,N_1079,N_1385);
or U1571 (N_1571,N_1224,N_1167);
and U1572 (N_1572,N_1300,N_1186);
and U1573 (N_1573,N_1194,N_950);
or U1574 (N_1574,N_1323,N_1496);
nand U1575 (N_1575,N_1288,N_1256);
or U1576 (N_1576,N_1287,N_1026);
nand U1577 (N_1577,N_775,N_1059);
or U1578 (N_1578,N_777,N_931);
xnor U1579 (N_1579,N_1487,N_1397);
and U1580 (N_1580,N_828,N_1263);
nor U1581 (N_1581,N_1180,N_1202);
nor U1582 (N_1582,N_1334,N_761);
nor U1583 (N_1583,N_907,N_973);
and U1584 (N_1584,N_1391,N_1198);
nand U1585 (N_1585,N_767,N_809);
nor U1586 (N_1586,N_1060,N_1355);
nor U1587 (N_1587,N_1253,N_1039);
xor U1588 (N_1588,N_1295,N_1000);
nand U1589 (N_1589,N_1273,N_1337);
nor U1590 (N_1590,N_1303,N_833);
nor U1591 (N_1591,N_784,N_1234);
and U1592 (N_1592,N_1007,N_1312);
and U1593 (N_1593,N_1293,N_1044);
nand U1594 (N_1594,N_1066,N_1242);
and U1595 (N_1595,N_953,N_1003);
nor U1596 (N_1596,N_1283,N_1459);
or U1597 (N_1597,N_1020,N_1277);
nand U1598 (N_1598,N_1104,N_893);
or U1599 (N_1599,N_1428,N_1244);
and U1600 (N_1600,N_1402,N_927);
nor U1601 (N_1601,N_1399,N_801);
nor U1602 (N_1602,N_839,N_832);
nor U1603 (N_1603,N_1158,N_1490);
nand U1604 (N_1604,N_998,N_957);
nand U1605 (N_1605,N_1479,N_795);
nand U1606 (N_1606,N_1262,N_1432);
and U1607 (N_1607,N_1322,N_816);
xnor U1608 (N_1608,N_955,N_1439);
xor U1609 (N_1609,N_988,N_1258);
nand U1610 (N_1610,N_1249,N_1423);
or U1611 (N_1611,N_867,N_1469);
nor U1612 (N_1612,N_1115,N_1199);
nand U1613 (N_1613,N_803,N_1266);
xor U1614 (N_1614,N_1259,N_1032);
and U1615 (N_1615,N_1069,N_1381);
nand U1616 (N_1616,N_1030,N_1238);
nand U1617 (N_1617,N_1033,N_849);
and U1618 (N_1618,N_1089,N_770);
nor U1619 (N_1619,N_897,N_796);
and U1620 (N_1620,N_794,N_1408);
nand U1621 (N_1621,N_1425,N_1243);
nand U1622 (N_1622,N_1444,N_771);
nand U1623 (N_1623,N_769,N_1380);
xnor U1624 (N_1624,N_887,N_1370);
or U1625 (N_1625,N_1144,N_1450);
and U1626 (N_1626,N_902,N_1461);
or U1627 (N_1627,N_1296,N_791);
nand U1628 (N_1628,N_822,N_1429);
and U1629 (N_1629,N_1350,N_1093);
or U1630 (N_1630,N_788,N_1148);
nor U1631 (N_1631,N_766,N_1053);
or U1632 (N_1632,N_1489,N_892);
xnor U1633 (N_1633,N_1276,N_1270);
or U1634 (N_1634,N_1083,N_774);
nand U1635 (N_1635,N_1405,N_1046);
and U1636 (N_1636,N_1017,N_1204);
nor U1637 (N_1637,N_760,N_1076);
or U1638 (N_1638,N_965,N_1382);
nor U1639 (N_1639,N_932,N_1108);
or U1640 (N_1640,N_912,N_1002);
or U1641 (N_1641,N_1366,N_985);
or U1642 (N_1642,N_1246,N_778);
nor U1643 (N_1643,N_1021,N_1137);
nand U1644 (N_1644,N_972,N_899);
or U1645 (N_1645,N_941,N_757);
nor U1646 (N_1646,N_1229,N_987);
nand U1647 (N_1647,N_1360,N_1403);
and U1648 (N_1648,N_865,N_1201);
and U1649 (N_1649,N_982,N_1043);
nand U1650 (N_1650,N_1211,N_1004);
nor U1651 (N_1651,N_1404,N_1318);
and U1652 (N_1652,N_845,N_1058);
or U1653 (N_1653,N_1257,N_1379);
nand U1654 (N_1654,N_1174,N_1077);
and U1655 (N_1655,N_834,N_1463);
and U1656 (N_1656,N_813,N_1413);
and U1657 (N_1657,N_980,N_1010);
nand U1658 (N_1658,N_1495,N_884);
nand U1659 (N_1659,N_1431,N_933);
or U1660 (N_1660,N_901,N_1477);
nor U1661 (N_1661,N_1261,N_752);
and U1662 (N_1662,N_1050,N_1448);
and U1663 (N_1663,N_948,N_1019);
nor U1664 (N_1664,N_776,N_1025);
nor U1665 (N_1665,N_835,N_1172);
nor U1666 (N_1666,N_1001,N_1354);
xor U1667 (N_1667,N_1195,N_1421);
nand U1668 (N_1668,N_1435,N_1321);
and U1669 (N_1669,N_975,N_989);
xor U1670 (N_1670,N_753,N_1455);
nor U1671 (N_1671,N_756,N_1367);
or U1672 (N_1672,N_1269,N_969);
or U1673 (N_1673,N_1470,N_758);
and U1674 (N_1674,N_1275,N_1409);
or U1675 (N_1675,N_1177,N_1427);
nor U1676 (N_1676,N_936,N_1473);
nor U1677 (N_1677,N_1143,N_908);
and U1678 (N_1678,N_1449,N_1065);
xor U1679 (N_1679,N_1254,N_787);
and U1680 (N_1680,N_1416,N_997);
and U1681 (N_1681,N_1213,N_811);
xor U1682 (N_1682,N_1418,N_909);
nor U1683 (N_1683,N_860,N_1414);
and U1684 (N_1684,N_1124,N_871);
nor U1685 (N_1685,N_1274,N_914);
and U1686 (N_1686,N_1075,N_1457);
and U1687 (N_1687,N_876,N_1387);
nand U1688 (N_1688,N_1412,N_1231);
or U1689 (N_1689,N_1407,N_1307);
or U1690 (N_1690,N_844,N_1197);
nor U1691 (N_1691,N_1400,N_981);
or U1692 (N_1692,N_763,N_1045);
nand U1693 (N_1693,N_1164,N_1221);
xor U1694 (N_1694,N_962,N_1190);
and U1695 (N_1695,N_1031,N_1325);
nor U1696 (N_1696,N_1482,N_1327);
or U1697 (N_1697,N_1080,N_1471);
nor U1698 (N_1698,N_829,N_1395);
nor U1699 (N_1699,N_977,N_802);
or U1700 (N_1700,N_910,N_937);
nand U1701 (N_1701,N_1264,N_1294);
or U1702 (N_1702,N_1107,N_1055);
or U1703 (N_1703,N_799,N_1156);
and U1704 (N_1704,N_814,N_827);
nor U1705 (N_1705,N_916,N_1236);
nor U1706 (N_1706,N_1392,N_1305);
nand U1707 (N_1707,N_888,N_856);
nor U1708 (N_1708,N_1071,N_793);
and U1709 (N_1709,N_1064,N_1341);
xor U1710 (N_1710,N_1084,N_1415);
nand U1711 (N_1711,N_1443,N_1324);
nand U1712 (N_1712,N_1248,N_1227);
nand U1713 (N_1713,N_1233,N_1442);
and U1714 (N_1714,N_1191,N_959);
xnor U1715 (N_1715,N_1015,N_1153);
or U1716 (N_1716,N_961,N_1073);
or U1717 (N_1717,N_798,N_1319);
nand U1718 (N_1718,N_1127,N_1304);
or U1719 (N_1719,N_837,N_923);
nor U1720 (N_1720,N_1068,N_852);
or U1721 (N_1721,N_1160,N_1394);
and U1722 (N_1722,N_1086,N_783);
or U1723 (N_1723,N_850,N_1478);
nor U1724 (N_1724,N_1332,N_1036);
and U1725 (N_1725,N_1309,N_1151);
nand U1726 (N_1726,N_869,N_1027);
nor U1727 (N_1727,N_1331,N_913);
and U1728 (N_1728,N_781,N_1465);
xor U1729 (N_1729,N_889,N_1317);
or U1730 (N_1730,N_1203,N_1049);
or U1731 (N_1731,N_1018,N_1123);
nand U1732 (N_1732,N_951,N_1426);
or U1733 (N_1733,N_1168,N_1375);
and U1734 (N_1734,N_879,N_1128);
nand U1735 (N_1735,N_915,N_1165);
nand U1736 (N_1736,N_1040,N_836);
and U1737 (N_1737,N_1493,N_900);
or U1738 (N_1738,N_947,N_1393);
nand U1739 (N_1739,N_1481,N_1022);
or U1740 (N_1740,N_1268,N_1184);
nand U1741 (N_1741,N_1014,N_1492);
or U1742 (N_1742,N_1377,N_1241);
and U1743 (N_1743,N_1430,N_885);
and U1744 (N_1744,N_1125,N_1223);
and U1745 (N_1745,N_918,N_819);
nor U1746 (N_1746,N_868,N_1117);
nor U1747 (N_1747,N_1013,N_866);
nor U1748 (N_1748,N_971,N_1122);
nand U1749 (N_1749,N_1499,N_1386);
nand U1750 (N_1750,N_1271,N_755);
nand U1751 (N_1751,N_894,N_1299);
nor U1752 (N_1752,N_1311,N_1150);
and U1753 (N_1753,N_970,N_1356);
nor U1754 (N_1754,N_751,N_1023);
or U1755 (N_1755,N_1121,N_825);
nor U1756 (N_1756,N_917,N_1445);
nand U1757 (N_1757,N_785,N_1182);
nand U1758 (N_1758,N_1016,N_1120);
or U1759 (N_1759,N_773,N_1193);
and U1760 (N_1760,N_1038,N_823);
nor U1761 (N_1761,N_1353,N_821);
or U1762 (N_1762,N_1316,N_1005);
nor U1763 (N_1763,N_797,N_896);
nor U1764 (N_1764,N_942,N_999);
nand U1765 (N_1765,N_854,N_1087);
and U1766 (N_1766,N_808,N_1133);
xor U1767 (N_1767,N_863,N_1245);
nand U1768 (N_1768,N_1090,N_1054);
or U1769 (N_1769,N_1157,N_1362);
nand U1770 (N_1770,N_1411,N_824);
nor U1771 (N_1771,N_1183,N_1132);
nor U1772 (N_1772,N_800,N_877);
or U1773 (N_1773,N_1009,N_1371);
xor U1774 (N_1774,N_1376,N_878);
nand U1775 (N_1775,N_1228,N_1251);
nand U1776 (N_1776,N_882,N_1267);
nand U1777 (N_1777,N_1438,N_1175);
nor U1778 (N_1778,N_848,N_1339);
nand U1779 (N_1779,N_1152,N_1282);
and U1780 (N_1780,N_1474,N_963);
xnor U1781 (N_1781,N_1255,N_1396);
nand U1782 (N_1782,N_934,N_1206);
nand U1783 (N_1783,N_861,N_1126);
xor U1784 (N_1784,N_1320,N_1468);
or U1785 (N_1785,N_929,N_1214);
xor U1786 (N_1786,N_792,N_949);
nand U1787 (N_1787,N_1208,N_1142);
or U1788 (N_1788,N_1436,N_1081);
and U1789 (N_1789,N_1301,N_1178);
nand U1790 (N_1790,N_820,N_1169);
nor U1791 (N_1791,N_851,N_995);
nand U1792 (N_1792,N_944,N_1091);
or U1793 (N_1793,N_1485,N_1260);
nor U1794 (N_1794,N_964,N_1351);
nor U1795 (N_1795,N_1406,N_779);
nor U1796 (N_1796,N_1106,N_874);
and U1797 (N_1797,N_945,N_1291);
and U1798 (N_1798,N_1110,N_1179);
nand U1799 (N_1799,N_1239,N_1215);
nor U1800 (N_1800,N_924,N_1111);
xor U1801 (N_1801,N_954,N_1119);
or U1802 (N_1802,N_1240,N_1368);
and U1803 (N_1803,N_1134,N_1306);
or U1804 (N_1804,N_1357,N_805);
and U1805 (N_1805,N_1359,N_983);
and U1806 (N_1806,N_1092,N_1342);
and U1807 (N_1807,N_1464,N_855);
nand U1808 (N_1808,N_1313,N_1147);
or U1809 (N_1809,N_1141,N_1095);
nor U1810 (N_1810,N_1140,N_1192);
nor U1811 (N_1811,N_1326,N_870);
and U1812 (N_1812,N_1222,N_1062);
xnor U1813 (N_1813,N_764,N_1388);
nor U1814 (N_1814,N_1494,N_1209);
nand U1815 (N_1815,N_903,N_1486);
or U1816 (N_1816,N_976,N_1057);
nor U1817 (N_1817,N_872,N_1475);
nand U1818 (N_1818,N_1187,N_812);
and U1819 (N_1819,N_838,N_890);
nand U1820 (N_1820,N_789,N_765);
xor U1821 (N_1821,N_1292,N_1217);
and U1822 (N_1822,N_1096,N_974);
and U1823 (N_1823,N_928,N_1466);
and U1824 (N_1824,N_859,N_1226);
nand U1825 (N_1825,N_1042,N_1185);
nand U1826 (N_1826,N_1063,N_858);
or U1827 (N_1827,N_1488,N_1034);
nor U1828 (N_1828,N_1345,N_967);
xor U1829 (N_1829,N_1210,N_979);
nand U1830 (N_1830,N_1462,N_1364);
nor U1831 (N_1831,N_1346,N_906);
nand U1832 (N_1832,N_1012,N_1118);
and U1833 (N_1833,N_1028,N_1401);
nor U1834 (N_1834,N_1452,N_926);
and U1835 (N_1835,N_1070,N_1171);
or U1836 (N_1836,N_1361,N_759);
nand U1837 (N_1837,N_1480,N_994);
nor U1838 (N_1838,N_1230,N_895);
nor U1839 (N_1839,N_1225,N_919);
or U1840 (N_1840,N_1365,N_1374);
and U1841 (N_1841,N_1422,N_1278);
nor U1842 (N_1842,N_1145,N_1389);
nor U1843 (N_1843,N_920,N_1252);
or U1844 (N_1844,N_1116,N_1008);
nor U1845 (N_1845,N_1338,N_993);
and U1846 (N_1846,N_1344,N_1349);
nand U1847 (N_1847,N_880,N_891);
and U1848 (N_1848,N_1114,N_831);
nor U1849 (N_1849,N_1250,N_1155);
and U1850 (N_1850,N_1161,N_1051);
or U1851 (N_1851,N_815,N_857);
and U1852 (N_1852,N_1029,N_1220);
nor U1853 (N_1853,N_1067,N_1460);
or U1854 (N_1854,N_1136,N_1085);
nor U1855 (N_1855,N_1232,N_968);
xnor U1856 (N_1856,N_1467,N_1330);
and U1857 (N_1857,N_1011,N_1280);
xor U1858 (N_1858,N_1189,N_1378);
nand U1859 (N_1859,N_780,N_1181);
nand U1860 (N_1860,N_817,N_925);
nor U1861 (N_1861,N_1163,N_1453);
xnor U1862 (N_1862,N_1129,N_1162);
xor U1863 (N_1863,N_939,N_1047);
nand U1864 (N_1864,N_1074,N_1329);
nor U1865 (N_1865,N_1383,N_1290);
or U1866 (N_1866,N_750,N_842);
nand U1867 (N_1867,N_1247,N_996);
and U1868 (N_1868,N_946,N_952);
and U1869 (N_1869,N_943,N_1447);
and U1870 (N_1870,N_862,N_1328);
or U1871 (N_1871,N_1101,N_1149);
xor U1872 (N_1872,N_1373,N_1308);
nand U1873 (N_1873,N_1410,N_1286);
nand U1874 (N_1874,N_826,N_846);
xor U1875 (N_1875,N_1076,N_1385);
nor U1876 (N_1876,N_869,N_1424);
and U1877 (N_1877,N_803,N_1323);
nand U1878 (N_1878,N_1223,N_757);
and U1879 (N_1879,N_792,N_898);
nand U1880 (N_1880,N_1020,N_1366);
and U1881 (N_1881,N_1149,N_1170);
nand U1882 (N_1882,N_1113,N_866);
or U1883 (N_1883,N_1224,N_1187);
xor U1884 (N_1884,N_1137,N_778);
or U1885 (N_1885,N_937,N_752);
nor U1886 (N_1886,N_1288,N_974);
and U1887 (N_1887,N_1339,N_850);
and U1888 (N_1888,N_787,N_1205);
and U1889 (N_1889,N_1450,N_834);
nor U1890 (N_1890,N_791,N_758);
and U1891 (N_1891,N_1441,N_1322);
or U1892 (N_1892,N_854,N_1125);
nand U1893 (N_1893,N_1383,N_1043);
nor U1894 (N_1894,N_1028,N_1021);
nor U1895 (N_1895,N_877,N_1258);
and U1896 (N_1896,N_1315,N_789);
or U1897 (N_1897,N_1166,N_835);
or U1898 (N_1898,N_1126,N_1463);
nor U1899 (N_1899,N_1200,N_1274);
nor U1900 (N_1900,N_1380,N_971);
nand U1901 (N_1901,N_1455,N_991);
nand U1902 (N_1902,N_1323,N_1147);
nor U1903 (N_1903,N_1443,N_1353);
nand U1904 (N_1904,N_850,N_824);
or U1905 (N_1905,N_1183,N_1479);
nor U1906 (N_1906,N_1379,N_1217);
nor U1907 (N_1907,N_1394,N_844);
and U1908 (N_1908,N_1320,N_1176);
or U1909 (N_1909,N_866,N_1416);
nand U1910 (N_1910,N_1283,N_1267);
and U1911 (N_1911,N_1382,N_1234);
or U1912 (N_1912,N_1290,N_1286);
nor U1913 (N_1913,N_830,N_920);
nand U1914 (N_1914,N_966,N_806);
and U1915 (N_1915,N_1147,N_1476);
and U1916 (N_1916,N_911,N_1076);
or U1917 (N_1917,N_1045,N_1183);
and U1918 (N_1918,N_1370,N_1206);
or U1919 (N_1919,N_1138,N_1037);
xnor U1920 (N_1920,N_1341,N_1069);
nand U1921 (N_1921,N_935,N_1391);
and U1922 (N_1922,N_1467,N_1328);
and U1923 (N_1923,N_882,N_988);
nand U1924 (N_1924,N_1300,N_1013);
nand U1925 (N_1925,N_1319,N_1136);
or U1926 (N_1926,N_861,N_1103);
nor U1927 (N_1927,N_1107,N_982);
nand U1928 (N_1928,N_1446,N_1283);
nand U1929 (N_1929,N_1255,N_981);
and U1930 (N_1930,N_1002,N_1396);
or U1931 (N_1931,N_1287,N_1056);
nor U1932 (N_1932,N_874,N_1384);
and U1933 (N_1933,N_1314,N_1174);
or U1934 (N_1934,N_1113,N_897);
nand U1935 (N_1935,N_1317,N_1403);
xor U1936 (N_1936,N_825,N_1344);
and U1937 (N_1937,N_801,N_1057);
or U1938 (N_1938,N_1070,N_872);
or U1939 (N_1939,N_1283,N_1098);
or U1940 (N_1940,N_1276,N_1150);
or U1941 (N_1941,N_1494,N_1307);
nor U1942 (N_1942,N_918,N_1359);
nand U1943 (N_1943,N_964,N_1120);
nor U1944 (N_1944,N_1026,N_1353);
nor U1945 (N_1945,N_1305,N_827);
and U1946 (N_1946,N_1015,N_753);
nand U1947 (N_1947,N_802,N_1131);
nor U1948 (N_1948,N_886,N_1077);
nor U1949 (N_1949,N_1484,N_776);
or U1950 (N_1950,N_1126,N_777);
and U1951 (N_1951,N_849,N_1147);
and U1952 (N_1952,N_1243,N_1133);
or U1953 (N_1953,N_1032,N_955);
nor U1954 (N_1954,N_1496,N_1187);
xor U1955 (N_1955,N_1295,N_1133);
and U1956 (N_1956,N_1253,N_1485);
nand U1957 (N_1957,N_867,N_1357);
nand U1958 (N_1958,N_827,N_1332);
or U1959 (N_1959,N_1026,N_1211);
nor U1960 (N_1960,N_993,N_837);
nand U1961 (N_1961,N_1269,N_926);
nor U1962 (N_1962,N_841,N_959);
or U1963 (N_1963,N_1260,N_947);
and U1964 (N_1964,N_1372,N_1443);
xnor U1965 (N_1965,N_1291,N_987);
nor U1966 (N_1966,N_942,N_823);
nor U1967 (N_1967,N_1218,N_949);
or U1968 (N_1968,N_886,N_911);
or U1969 (N_1969,N_764,N_808);
nor U1970 (N_1970,N_1295,N_1007);
nor U1971 (N_1971,N_1283,N_1273);
and U1972 (N_1972,N_997,N_971);
nand U1973 (N_1973,N_1456,N_1152);
nor U1974 (N_1974,N_1013,N_1066);
and U1975 (N_1975,N_1487,N_1262);
or U1976 (N_1976,N_773,N_1330);
nand U1977 (N_1977,N_1069,N_1145);
nor U1978 (N_1978,N_1357,N_912);
or U1979 (N_1979,N_1045,N_798);
and U1980 (N_1980,N_983,N_1114);
nor U1981 (N_1981,N_1426,N_1256);
and U1982 (N_1982,N_1012,N_990);
xnor U1983 (N_1983,N_997,N_1458);
nand U1984 (N_1984,N_1389,N_1397);
nand U1985 (N_1985,N_1029,N_1378);
nand U1986 (N_1986,N_1117,N_1105);
and U1987 (N_1987,N_941,N_893);
nand U1988 (N_1988,N_1399,N_1189);
nand U1989 (N_1989,N_1141,N_1284);
and U1990 (N_1990,N_1279,N_1120);
nand U1991 (N_1991,N_812,N_1409);
or U1992 (N_1992,N_956,N_1458);
nand U1993 (N_1993,N_1233,N_1165);
or U1994 (N_1994,N_1062,N_1256);
xnor U1995 (N_1995,N_1453,N_834);
and U1996 (N_1996,N_1323,N_1258);
or U1997 (N_1997,N_796,N_1017);
and U1998 (N_1998,N_1040,N_1382);
and U1999 (N_1999,N_784,N_1431);
or U2000 (N_2000,N_1477,N_1406);
and U2001 (N_2001,N_867,N_878);
or U2002 (N_2002,N_1121,N_1329);
and U2003 (N_2003,N_1415,N_1030);
nor U2004 (N_2004,N_848,N_1070);
xnor U2005 (N_2005,N_826,N_862);
and U2006 (N_2006,N_1179,N_892);
nor U2007 (N_2007,N_964,N_809);
nand U2008 (N_2008,N_1246,N_1353);
xor U2009 (N_2009,N_783,N_1171);
nor U2010 (N_2010,N_980,N_875);
nand U2011 (N_2011,N_1196,N_1045);
nand U2012 (N_2012,N_1396,N_897);
nand U2013 (N_2013,N_1099,N_1203);
nor U2014 (N_2014,N_1217,N_801);
nand U2015 (N_2015,N_856,N_1146);
xnor U2016 (N_2016,N_1320,N_841);
or U2017 (N_2017,N_906,N_867);
or U2018 (N_2018,N_971,N_1412);
or U2019 (N_2019,N_1328,N_830);
nand U2020 (N_2020,N_1068,N_968);
and U2021 (N_2021,N_852,N_1292);
or U2022 (N_2022,N_1357,N_996);
or U2023 (N_2023,N_1093,N_1180);
nor U2024 (N_2024,N_895,N_1341);
or U2025 (N_2025,N_913,N_1362);
and U2026 (N_2026,N_876,N_1492);
nor U2027 (N_2027,N_1415,N_789);
nand U2028 (N_2028,N_1304,N_1232);
or U2029 (N_2029,N_1366,N_1189);
nor U2030 (N_2030,N_843,N_1324);
or U2031 (N_2031,N_1332,N_1490);
nor U2032 (N_2032,N_952,N_1344);
nand U2033 (N_2033,N_833,N_1362);
and U2034 (N_2034,N_877,N_1170);
nor U2035 (N_2035,N_902,N_966);
or U2036 (N_2036,N_840,N_1111);
nor U2037 (N_2037,N_1300,N_863);
and U2038 (N_2038,N_873,N_1334);
and U2039 (N_2039,N_1273,N_841);
or U2040 (N_2040,N_1003,N_1401);
nand U2041 (N_2041,N_1066,N_1386);
or U2042 (N_2042,N_1033,N_874);
and U2043 (N_2043,N_1110,N_973);
nor U2044 (N_2044,N_1227,N_1357);
nand U2045 (N_2045,N_1126,N_941);
xor U2046 (N_2046,N_1261,N_1073);
and U2047 (N_2047,N_1318,N_958);
and U2048 (N_2048,N_1184,N_1446);
nand U2049 (N_2049,N_1207,N_875);
and U2050 (N_2050,N_1326,N_1273);
or U2051 (N_2051,N_1062,N_917);
or U2052 (N_2052,N_1238,N_966);
nor U2053 (N_2053,N_1424,N_1221);
xor U2054 (N_2054,N_848,N_1369);
and U2055 (N_2055,N_1475,N_756);
nor U2056 (N_2056,N_1070,N_887);
nand U2057 (N_2057,N_943,N_1220);
and U2058 (N_2058,N_1174,N_1178);
xor U2059 (N_2059,N_1110,N_1487);
nor U2060 (N_2060,N_777,N_1145);
nand U2061 (N_2061,N_1345,N_1356);
nor U2062 (N_2062,N_1227,N_1150);
and U2063 (N_2063,N_752,N_1474);
and U2064 (N_2064,N_1103,N_961);
or U2065 (N_2065,N_781,N_1313);
or U2066 (N_2066,N_842,N_1289);
nor U2067 (N_2067,N_1047,N_1357);
nor U2068 (N_2068,N_1258,N_1455);
nor U2069 (N_2069,N_955,N_1020);
and U2070 (N_2070,N_1059,N_799);
nor U2071 (N_2071,N_794,N_1271);
nor U2072 (N_2072,N_1419,N_1262);
and U2073 (N_2073,N_1392,N_1024);
and U2074 (N_2074,N_1136,N_1417);
nand U2075 (N_2075,N_965,N_1082);
and U2076 (N_2076,N_861,N_1494);
and U2077 (N_2077,N_804,N_1412);
and U2078 (N_2078,N_1135,N_1426);
xnor U2079 (N_2079,N_829,N_1478);
nor U2080 (N_2080,N_1320,N_1331);
or U2081 (N_2081,N_1006,N_1250);
and U2082 (N_2082,N_1189,N_1383);
nand U2083 (N_2083,N_1246,N_844);
nor U2084 (N_2084,N_1044,N_1030);
nand U2085 (N_2085,N_1348,N_1280);
and U2086 (N_2086,N_815,N_1043);
nor U2087 (N_2087,N_1372,N_1044);
nor U2088 (N_2088,N_818,N_1362);
or U2089 (N_2089,N_800,N_1157);
and U2090 (N_2090,N_1233,N_1222);
nor U2091 (N_2091,N_1193,N_1435);
xor U2092 (N_2092,N_973,N_835);
or U2093 (N_2093,N_1410,N_958);
or U2094 (N_2094,N_1148,N_1253);
and U2095 (N_2095,N_1187,N_1386);
nand U2096 (N_2096,N_906,N_859);
xor U2097 (N_2097,N_1235,N_1122);
or U2098 (N_2098,N_1394,N_1271);
nand U2099 (N_2099,N_756,N_1150);
nand U2100 (N_2100,N_1066,N_910);
nor U2101 (N_2101,N_898,N_1213);
and U2102 (N_2102,N_1346,N_979);
nand U2103 (N_2103,N_1011,N_1130);
or U2104 (N_2104,N_769,N_1163);
and U2105 (N_2105,N_820,N_935);
nor U2106 (N_2106,N_1404,N_1312);
or U2107 (N_2107,N_1381,N_1386);
nand U2108 (N_2108,N_887,N_901);
nor U2109 (N_2109,N_838,N_1033);
or U2110 (N_2110,N_1459,N_1336);
xor U2111 (N_2111,N_1111,N_1209);
nand U2112 (N_2112,N_1070,N_1367);
and U2113 (N_2113,N_1201,N_1265);
nand U2114 (N_2114,N_1118,N_1389);
nand U2115 (N_2115,N_1335,N_1186);
or U2116 (N_2116,N_1235,N_1191);
nor U2117 (N_2117,N_1284,N_952);
and U2118 (N_2118,N_752,N_1111);
and U2119 (N_2119,N_1467,N_1097);
nand U2120 (N_2120,N_1155,N_1384);
nand U2121 (N_2121,N_765,N_1239);
nand U2122 (N_2122,N_1412,N_1361);
nand U2123 (N_2123,N_982,N_1327);
and U2124 (N_2124,N_1069,N_884);
nor U2125 (N_2125,N_1111,N_962);
nand U2126 (N_2126,N_924,N_1071);
and U2127 (N_2127,N_1125,N_1110);
nor U2128 (N_2128,N_1206,N_1040);
or U2129 (N_2129,N_808,N_1475);
nand U2130 (N_2130,N_1255,N_760);
nand U2131 (N_2131,N_1404,N_974);
or U2132 (N_2132,N_1264,N_1123);
or U2133 (N_2133,N_1287,N_1430);
nor U2134 (N_2134,N_1095,N_831);
nand U2135 (N_2135,N_1295,N_1243);
nand U2136 (N_2136,N_1420,N_1104);
and U2137 (N_2137,N_1269,N_1468);
nand U2138 (N_2138,N_1114,N_1496);
and U2139 (N_2139,N_870,N_1110);
nand U2140 (N_2140,N_766,N_1175);
nand U2141 (N_2141,N_858,N_1028);
nand U2142 (N_2142,N_966,N_928);
nor U2143 (N_2143,N_988,N_1475);
nor U2144 (N_2144,N_929,N_1260);
nor U2145 (N_2145,N_1271,N_883);
nor U2146 (N_2146,N_1107,N_1471);
nand U2147 (N_2147,N_1305,N_989);
nor U2148 (N_2148,N_885,N_1171);
nor U2149 (N_2149,N_818,N_1267);
nand U2150 (N_2150,N_1204,N_992);
and U2151 (N_2151,N_1134,N_1465);
or U2152 (N_2152,N_1078,N_1345);
or U2153 (N_2153,N_981,N_1067);
nand U2154 (N_2154,N_1108,N_1059);
and U2155 (N_2155,N_997,N_1272);
nor U2156 (N_2156,N_1204,N_792);
or U2157 (N_2157,N_984,N_963);
nand U2158 (N_2158,N_1238,N_1311);
and U2159 (N_2159,N_1355,N_1236);
and U2160 (N_2160,N_1275,N_1455);
and U2161 (N_2161,N_1491,N_1035);
and U2162 (N_2162,N_834,N_751);
xnor U2163 (N_2163,N_754,N_846);
and U2164 (N_2164,N_1036,N_1388);
nand U2165 (N_2165,N_1263,N_908);
nor U2166 (N_2166,N_982,N_1307);
and U2167 (N_2167,N_768,N_1392);
and U2168 (N_2168,N_1491,N_946);
nand U2169 (N_2169,N_1191,N_1063);
nor U2170 (N_2170,N_1168,N_1461);
nand U2171 (N_2171,N_834,N_1076);
and U2172 (N_2172,N_844,N_1305);
and U2173 (N_2173,N_1119,N_1202);
nor U2174 (N_2174,N_1412,N_1188);
nand U2175 (N_2175,N_1449,N_1324);
or U2176 (N_2176,N_833,N_1309);
xor U2177 (N_2177,N_831,N_1060);
or U2178 (N_2178,N_1072,N_1224);
nor U2179 (N_2179,N_876,N_1187);
and U2180 (N_2180,N_1070,N_1000);
xor U2181 (N_2181,N_794,N_880);
nand U2182 (N_2182,N_1485,N_975);
nand U2183 (N_2183,N_1123,N_1219);
nand U2184 (N_2184,N_953,N_1119);
or U2185 (N_2185,N_1147,N_1110);
xor U2186 (N_2186,N_812,N_857);
or U2187 (N_2187,N_1335,N_1438);
nand U2188 (N_2188,N_1388,N_1363);
nand U2189 (N_2189,N_768,N_797);
nor U2190 (N_2190,N_990,N_798);
nand U2191 (N_2191,N_1020,N_1488);
nand U2192 (N_2192,N_1142,N_983);
or U2193 (N_2193,N_780,N_1254);
or U2194 (N_2194,N_1411,N_1092);
or U2195 (N_2195,N_1054,N_1240);
nand U2196 (N_2196,N_1131,N_1337);
and U2197 (N_2197,N_1148,N_852);
and U2198 (N_2198,N_1240,N_1294);
and U2199 (N_2199,N_1210,N_1449);
nand U2200 (N_2200,N_1329,N_1258);
and U2201 (N_2201,N_979,N_1325);
and U2202 (N_2202,N_917,N_1344);
and U2203 (N_2203,N_1376,N_1126);
and U2204 (N_2204,N_1434,N_1184);
or U2205 (N_2205,N_882,N_1382);
nor U2206 (N_2206,N_1153,N_1122);
xor U2207 (N_2207,N_1080,N_786);
xor U2208 (N_2208,N_1447,N_1213);
nand U2209 (N_2209,N_1370,N_1261);
or U2210 (N_2210,N_1275,N_773);
nand U2211 (N_2211,N_1110,N_1181);
or U2212 (N_2212,N_1274,N_952);
nand U2213 (N_2213,N_769,N_1211);
and U2214 (N_2214,N_837,N_1371);
and U2215 (N_2215,N_1254,N_1273);
nand U2216 (N_2216,N_1047,N_961);
or U2217 (N_2217,N_1277,N_969);
nor U2218 (N_2218,N_1021,N_824);
xor U2219 (N_2219,N_1414,N_1405);
or U2220 (N_2220,N_999,N_1072);
nor U2221 (N_2221,N_813,N_905);
nor U2222 (N_2222,N_1062,N_766);
nand U2223 (N_2223,N_1498,N_1105);
or U2224 (N_2224,N_1491,N_1297);
nand U2225 (N_2225,N_1252,N_819);
xor U2226 (N_2226,N_1164,N_1209);
or U2227 (N_2227,N_1390,N_1144);
or U2228 (N_2228,N_1465,N_1317);
nand U2229 (N_2229,N_1080,N_1475);
xor U2230 (N_2230,N_1321,N_1046);
nand U2231 (N_2231,N_1140,N_904);
xnor U2232 (N_2232,N_1373,N_1098);
nand U2233 (N_2233,N_914,N_1058);
nand U2234 (N_2234,N_960,N_1044);
and U2235 (N_2235,N_1453,N_1144);
nor U2236 (N_2236,N_1383,N_1039);
or U2237 (N_2237,N_1279,N_1026);
nor U2238 (N_2238,N_1390,N_1119);
and U2239 (N_2239,N_1006,N_792);
or U2240 (N_2240,N_1211,N_994);
or U2241 (N_2241,N_1317,N_1483);
and U2242 (N_2242,N_999,N_975);
or U2243 (N_2243,N_1166,N_1283);
or U2244 (N_2244,N_1441,N_785);
nand U2245 (N_2245,N_936,N_1299);
nor U2246 (N_2246,N_1180,N_1088);
and U2247 (N_2247,N_1010,N_1420);
nor U2248 (N_2248,N_1287,N_964);
or U2249 (N_2249,N_1200,N_1085);
nand U2250 (N_2250,N_1630,N_2056);
or U2251 (N_2251,N_1885,N_1677);
or U2252 (N_2252,N_1523,N_1957);
or U2253 (N_2253,N_2230,N_1644);
nor U2254 (N_2254,N_1655,N_1937);
nand U2255 (N_2255,N_2128,N_1809);
nor U2256 (N_2256,N_1807,N_1618);
and U2257 (N_2257,N_1609,N_1726);
nand U2258 (N_2258,N_1782,N_2028);
nor U2259 (N_2259,N_1679,N_1989);
nand U2260 (N_2260,N_1963,N_1821);
nor U2261 (N_2261,N_2108,N_1769);
nand U2262 (N_2262,N_2084,N_1858);
nand U2263 (N_2263,N_1999,N_2159);
xor U2264 (N_2264,N_1949,N_1757);
or U2265 (N_2265,N_1518,N_1725);
nor U2266 (N_2266,N_1990,N_1827);
and U2267 (N_2267,N_2175,N_1527);
or U2268 (N_2268,N_2190,N_1952);
nand U2269 (N_2269,N_2143,N_1652);
nor U2270 (N_2270,N_2112,N_2122);
and U2271 (N_2271,N_2186,N_1673);
or U2272 (N_2272,N_2129,N_1699);
or U2273 (N_2273,N_2031,N_2200);
xor U2274 (N_2274,N_1992,N_1773);
or U2275 (N_2275,N_1997,N_2106);
nor U2276 (N_2276,N_1903,N_2168);
nand U2277 (N_2277,N_1832,N_2064);
and U2278 (N_2278,N_2038,N_1824);
or U2279 (N_2279,N_2243,N_2061);
nor U2280 (N_2280,N_2119,N_2057);
and U2281 (N_2281,N_2059,N_1507);
and U2282 (N_2282,N_1660,N_1765);
nand U2283 (N_2283,N_2209,N_1982);
nor U2284 (N_2284,N_1927,N_1887);
nor U2285 (N_2285,N_1570,N_1924);
nand U2286 (N_2286,N_1939,N_1615);
nor U2287 (N_2287,N_1598,N_1863);
and U2288 (N_2288,N_1857,N_1948);
nand U2289 (N_2289,N_1607,N_2234);
nor U2290 (N_2290,N_1995,N_1503);
xor U2291 (N_2291,N_1713,N_2166);
nand U2292 (N_2292,N_2009,N_1859);
and U2293 (N_2293,N_1951,N_2094);
nor U2294 (N_2294,N_2051,N_1822);
xnor U2295 (N_2295,N_2073,N_1543);
nand U2296 (N_2296,N_2070,N_2172);
nand U2297 (N_2297,N_1978,N_1522);
and U2298 (N_2298,N_2184,N_2034);
or U2299 (N_2299,N_1826,N_1753);
and U2300 (N_2300,N_1813,N_2029);
or U2301 (N_2301,N_1623,N_2179);
nor U2302 (N_2302,N_1833,N_1945);
xnor U2303 (N_2303,N_1986,N_2077);
and U2304 (N_2304,N_1682,N_1843);
or U2305 (N_2305,N_1915,N_2016);
and U2306 (N_2306,N_1529,N_2237);
nor U2307 (N_2307,N_1834,N_1587);
nand U2308 (N_2308,N_1900,N_1720);
or U2309 (N_2309,N_1555,N_1818);
and U2310 (N_2310,N_2217,N_2127);
nand U2311 (N_2311,N_1586,N_1691);
and U2312 (N_2312,N_1576,N_2071);
nand U2313 (N_2313,N_2130,N_2219);
nand U2314 (N_2314,N_2080,N_2215);
nor U2315 (N_2315,N_1519,N_1916);
or U2316 (N_2316,N_2203,N_1983);
nor U2317 (N_2317,N_1538,N_1697);
nand U2318 (N_2318,N_1844,N_1902);
nor U2319 (N_2319,N_1793,N_1798);
or U2320 (N_2320,N_1656,N_1977);
nor U2321 (N_2321,N_1582,N_1645);
and U2322 (N_2322,N_2114,N_2185);
nor U2323 (N_2323,N_1906,N_1875);
and U2324 (N_2324,N_1705,N_1692);
and U2325 (N_2325,N_2150,N_1671);
nand U2326 (N_2326,N_1628,N_2220);
or U2327 (N_2327,N_2105,N_1647);
xnor U2328 (N_2328,N_1974,N_1800);
and U2329 (N_2329,N_1756,N_2148);
and U2330 (N_2330,N_1605,N_2082);
and U2331 (N_2331,N_2044,N_1931);
or U2332 (N_2332,N_1953,N_1544);
nand U2333 (N_2333,N_2235,N_1779);
and U2334 (N_2334,N_2183,N_1878);
and U2335 (N_2335,N_1583,N_1524);
and U2336 (N_2336,N_1867,N_2246);
nand U2337 (N_2337,N_1959,N_1721);
or U2338 (N_2338,N_1802,N_1954);
or U2339 (N_2339,N_2102,N_1670);
or U2340 (N_2340,N_2060,N_1817);
nor U2341 (N_2341,N_2205,N_2093);
and U2342 (N_2342,N_1661,N_1734);
nor U2343 (N_2343,N_2227,N_1861);
xor U2344 (N_2344,N_1577,N_2170);
nand U2345 (N_2345,N_1899,N_1530);
or U2346 (N_2346,N_1685,N_1556);
nand U2347 (N_2347,N_1636,N_1780);
and U2348 (N_2348,N_2229,N_2096);
or U2349 (N_2349,N_1996,N_1701);
nand U2350 (N_2350,N_1758,N_1790);
or U2351 (N_2351,N_2196,N_1872);
or U2352 (N_2352,N_1745,N_1898);
and U2353 (N_2353,N_1551,N_1847);
nand U2354 (N_2354,N_2189,N_2037);
or U2355 (N_2355,N_1869,N_2171);
or U2356 (N_2356,N_1508,N_1512);
and U2357 (N_2357,N_1526,N_1629);
nand U2358 (N_2358,N_1666,N_1866);
xor U2359 (N_2359,N_1568,N_1755);
and U2360 (N_2360,N_2055,N_2008);
nor U2361 (N_2361,N_2192,N_1921);
nand U2362 (N_2362,N_1525,N_2025);
or U2363 (N_2363,N_1668,N_2083);
nand U2364 (N_2364,N_1804,N_1676);
and U2365 (N_2365,N_2015,N_1542);
nand U2366 (N_2366,N_2231,N_2019);
nand U2367 (N_2367,N_2245,N_2117);
or U2368 (N_2368,N_1515,N_2144);
or U2369 (N_2369,N_2240,N_2221);
xnor U2370 (N_2370,N_1856,N_2027);
xnor U2371 (N_2371,N_2052,N_1942);
nor U2372 (N_2372,N_2075,N_2158);
nor U2373 (N_2373,N_1553,N_1766);
nor U2374 (N_2374,N_1751,N_2004);
nor U2375 (N_2375,N_1998,N_1830);
and U2376 (N_2376,N_1740,N_1894);
nand U2377 (N_2377,N_2062,N_2050);
nor U2378 (N_2378,N_1747,N_2123);
nor U2379 (N_2379,N_2091,N_2174);
or U2380 (N_2380,N_1729,N_1588);
and U2381 (N_2381,N_1723,N_1579);
nor U2382 (N_2382,N_1820,N_2046);
nand U2383 (N_2383,N_1981,N_1783);
nand U2384 (N_2384,N_2247,N_1732);
xnor U2385 (N_2385,N_2198,N_2173);
and U2386 (N_2386,N_1738,N_2089);
nor U2387 (N_2387,N_1781,N_2099);
nand U2388 (N_2388,N_2023,N_1606);
xnor U2389 (N_2389,N_1988,N_1626);
nand U2390 (N_2390,N_2022,N_1801);
nand U2391 (N_2391,N_1510,N_2239);
or U2392 (N_2392,N_2078,N_2156);
xor U2393 (N_2393,N_1689,N_2208);
and U2394 (N_2394,N_1509,N_1960);
or U2395 (N_2395,N_2041,N_1967);
or U2396 (N_2396,N_1908,N_1620);
and U2397 (N_2397,N_1882,N_2026);
or U2398 (N_2398,N_2012,N_1557);
xor U2399 (N_2399,N_1966,N_1639);
nand U2400 (N_2400,N_2118,N_1559);
or U2401 (N_2401,N_2216,N_2067);
and U2402 (N_2402,N_2151,N_2167);
or U2403 (N_2403,N_2146,N_1584);
nor U2404 (N_2404,N_2090,N_1835);
xor U2405 (N_2405,N_1654,N_2109);
or U2406 (N_2406,N_1502,N_1565);
and U2407 (N_2407,N_2201,N_1643);
nand U2408 (N_2408,N_1838,N_2104);
or U2409 (N_2409,N_1663,N_1973);
nand U2410 (N_2410,N_1961,N_2066);
nor U2411 (N_2411,N_2098,N_1597);
and U2412 (N_2412,N_1855,N_1575);
or U2413 (N_2413,N_1578,N_1547);
nand U2414 (N_2414,N_2054,N_1870);
nand U2415 (N_2415,N_1625,N_2202);
and U2416 (N_2416,N_2017,N_1760);
or U2417 (N_2417,N_2136,N_1562);
or U2418 (N_2418,N_1823,N_1871);
nand U2419 (N_2419,N_2191,N_1516);
nand U2420 (N_2420,N_1846,N_2107);
nand U2421 (N_2421,N_1651,N_2032);
nand U2422 (N_2422,N_2103,N_2135);
or U2423 (N_2423,N_2236,N_1560);
and U2424 (N_2424,N_1631,N_1836);
or U2425 (N_2425,N_1595,N_2018);
nor U2426 (N_2426,N_2228,N_1956);
nand U2427 (N_2427,N_1860,N_2030);
xor U2428 (N_2428,N_1828,N_1980);
or U2429 (N_2429,N_1710,N_2132);
and U2430 (N_2430,N_1714,N_1744);
nor U2431 (N_2431,N_1569,N_1864);
nand U2432 (N_2432,N_2048,N_1657);
xor U2433 (N_2433,N_1594,N_1994);
or U2434 (N_2434,N_1554,N_1501);
nand U2435 (N_2435,N_1791,N_2125);
and U2436 (N_2436,N_1923,N_1561);
nand U2437 (N_2437,N_1777,N_1684);
and U2438 (N_2438,N_2176,N_1612);
nor U2439 (N_2439,N_1593,N_2163);
or U2440 (N_2440,N_1795,N_1640);
nor U2441 (N_2441,N_1571,N_1500);
and U2442 (N_2442,N_1698,N_2131);
or U2443 (N_2443,N_1648,N_1881);
nor U2444 (N_2444,N_1849,N_1752);
nor U2445 (N_2445,N_1619,N_2120);
or U2446 (N_2446,N_1669,N_1541);
xor U2447 (N_2447,N_1778,N_1742);
xor U2448 (N_2448,N_2006,N_1922);
nand U2449 (N_2449,N_1808,N_2193);
or U2450 (N_2450,N_1914,N_2021);
nand U2451 (N_2451,N_1514,N_1733);
nand U2452 (N_2452,N_1536,N_1563);
nand U2453 (N_2453,N_2065,N_1877);
and U2454 (N_2454,N_1805,N_1520);
and U2455 (N_2455,N_1616,N_1944);
nand U2456 (N_2456,N_1789,N_2020);
or U2457 (N_2457,N_1581,N_1892);
or U2458 (N_2458,N_1947,N_1511);
and U2459 (N_2459,N_1506,N_1854);
nand U2460 (N_2460,N_1718,N_1950);
or U2461 (N_2461,N_2110,N_1969);
nor U2462 (N_2462,N_1589,N_1775);
or U2463 (N_2463,N_1750,N_1737);
nor U2464 (N_2464,N_1848,N_1600);
xnor U2465 (N_2465,N_1558,N_2223);
and U2466 (N_2466,N_1929,N_2002);
nand U2467 (N_2467,N_1935,N_1905);
nand U2468 (N_2468,N_1932,N_1816);
xor U2469 (N_2469,N_1591,N_1886);
and U2470 (N_2470,N_1614,N_1611);
xor U2471 (N_2471,N_1741,N_2047);
nor U2472 (N_2472,N_1608,N_1764);
nand U2473 (N_2473,N_1761,N_2072);
xor U2474 (N_2474,N_1604,N_2194);
or U2475 (N_2475,N_2141,N_1727);
xor U2476 (N_2476,N_2233,N_1984);
or U2477 (N_2477,N_1641,N_2182);
and U2478 (N_2478,N_1646,N_1672);
nand U2479 (N_2479,N_1624,N_1962);
or U2480 (N_2480,N_2133,N_1930);
and U2481 (N_2481,N_1938,N_2115);
nor U2482 (N_2482,N_1716,N_1549);
or U2483 (N_2483,N_2211,N_1674);
nor U2484 (N_2484,N_1889,N_2138);
and U2485 (N_2485,N_1683,N_1853);
or U2486 (N_2486,N_1724,N_1664);
or U2487 (N_2487,N_2005,N_1603);
nor U2488 (N_2488,N_2162,N_1715);
xor U2489 (N_2489,N_1888,N_1772);
nor U2490 (N_2490,N_2043,N_1896);
and U2491 (N_2491,N_1876,N_1814);
or U2492 (N_2492,N_1891,N_1993);
or U2493 (N_2493,N_2207,N_1776);
nor U2494 (N_2494,N_2111,N_1890);
or U2495 (N_2495,N_1552,N_1762);
nand U2496 (N_2496,N_1531,N_2232);
or U2497 (N_2497,N_1678,N_1601);
xnor U2498 (N_2498,N_1667,N_2042);
nor U2499 (N_2499,N_2188,N_1979);
or U2500 (N_2500,N_2014,N_1968);
or U2501 (N_2501,N_1943,N_1521);
nand U2502 (N_2502,N_1919,N_1545);
or U2503 (N_2503,N_1613,N_2181);
xnor U2504 (N_2504,N_1686,N_1596);
nor U2505 (N_2505,N_1786,N_1884);
nor U2506 (N_2506,N_1829,N_1774);
and U2507 (N_2507,N_2101,N_1627);
or U2508 (N_2508,N_2204,N_2213);
and U2509 (N_2509,N_1540,N_2137);
or U2510 (N_2510,N_1799,N_2079);
nor U2511 (N_2511,N_2160,N_1722);
xnor U2512 (N_2512,N_1653,N_1771);
nor U2513 (N_2513,N_2013,N_1650);
nor U2514 (N_2514,N_1632,N_1879);
xor U2515 (N_2515,N_1690,N_2214);
and U2516 (N_2516,N_2058,N_1706);
nand U2517 (N_2517,N_1880,N_1852);
and U2518 (N_2518,N_2036,N_2113);
and U2519 (N_2519,N_1926,N_1839);
nand U2520 (N_2520,N_2069,N_1748);
xor U2521 (N_2521,N_1895,N_1987);
or U2522 (N_2522,N_2092,N_1785);
nand U2523 (N_2523,N_1910,N_2199);
and U2524 (N_2524,N_1635,N_1633);
nor U2525 (N_2525,N_2157,N_1573);
nand U2526 (N_2526,N_1970,N_2076);
nor U2527 (N_2527,N_2081,N_1788);
or U2528 (N_2528,N_1688,N_2074);
or U2529 (N_2529,N_2153,N_1592);
xnor U2530 (N_2530,N_1976,N_1703);
nand U2531 (N_2531,N_1599,N_2124);
nand U2532 (N_2532,N_1546,N_1743);
and U2533 (N_2533,N_1504,N_1909);
nand U2534 (N_2534,N_2169,N_1911);
or U2535 (N_2535,N_1700,N_1680);
nand U2536 (N_2536,N_2241,N_1958);
or U2537 (N_2537,N_1746,N_1602);
or U2538 (N_2538,N_1711,N_1694);
nand U2539 (N_2539,N_2126,N_1675);
nand U2540 (N_2540,N_1649,N_1803);
and U2541 (N_2541,N_1897,N_1964);
or U2542 (N_2542,N_2007,N_2040);
and U2543 (N_2543,N_2155,N_1907);
and U2544 (N_2544,N_2039,N_1971);
xnor U2545 (N_2545,N_1883,N_1928);
nor U2546 (N_2546,N_1985,N_1768);
nand U2547 (N_2547,N_1787,N_1659);
nand U2548 (N_2548,N_1917,N_1893);
and U2549 (N_2549,N_2164,N_1505);
or U2550 (N_2550,N_1850,N_1810);
nor U2551 (N_2551,N_2033,N_1702);
and U2552 (N_2552,N_2085,N_2087);
xor U2553 (N_2553,N_2222,N_1638);
nand U2554 (N_2554,N_1831,N_1794);
and U2555 (N_2555,N_1658,N_2149);
or U2556 (N_2556,N_1566,N_1837);
or U2557 (N_2557,N_1851,N_2134);
xnor U2558 (N_2558,N_2000,N_1537);
nor U2559 (N_2559,N_1806,N_1572);
or U2560 (N_2560,N_1842,N_1585);
nor U2561 (N_2561,N_1717,N_2001);
or U2562 (N_2562,N_1840,N_1812);
or U2563 (N_2563,N_1532,N_2088);
nor U2564 (N_2564,N_1712,N_2242);
nand U2565 (N_2565,N_1622,N_1913);
or U2566 (N_2566,N_2049,N_1873);
and U2567 (N_2567,N_2024,N_1841);
xnor U2568 (N_2568,N_2086,N_1811);
or U2569 (N_2569,N_1634,N_2249);
or U2570 (N_2570,N_2053,N_1865);
and U2571 (N_2571,N_2152,N_1925);
xnor U2572 (N_2572,N_1533,N_1874);
or U2573 (N_2573,N_1972,N_2145);
and U2574 (N_2574,N_1617,N_2011);
or U2575 (N_2575,N_2063,N_1687);
or U2576 (N_2576,N_1610,N_2097);
nor U2577 (N_2577,N_1528,N_1567);
nand U2578 (N_2578,N_2121,N_2180);
and U2579 (N_2579,N_1735,N_1736);
or U2580 (N_2580,N_1792,N_1550);
nand U2581 (N_2581,N_2224,N_2218);
nand U2582 (N_2582,N_2177,N_1535);
nand U2583 (N_2583,N_1707,N_1719);
nor U2584 (N_2584,N_1590,N_1819);
nand U2585 (N_2585,N_2068,N_1797);
or U2586 (N_2586,N_1621,N_1796);
and U2587 (N_2587,N_2197,N_1946);
or U2588 (N_2588,N_1739,N_1564);
or U2589 (N_2589,N_1770,N_1934);
nor U2590 (N_2590,N_2100,N_2165);
or U2591 (N_2591,N_1642,N_1637);
nor U2592 (N_2592,N_1708,N_1825);
nor U2593 (N_2593,N_1696,N_1580);
xnor U2594 (N_2594,N_2244,N_2178);
and U2595 (N_2595,N_1539,N_1862);
and U2596 (N_2596,N_1681,N_1517);
nand U2597 (N_2597,N_1784,N_2226);
and U2598 (N_2598,N_1759,N_2161);
nand U2599 (N_2599,N_1709,N_1991);
nor U2600 (N_2600,N_1704,N_1920);
nand U2601 (N_2601,N_2003,N_2206);
nand U2602 (N_2602,N_2212,N_2210);
nand U2603 (N_2603,N_1662,N_1936);
nand U2604 (N_2604,N_1904,N_1763);
nand U2605 (N_2605,N_1534,N_2140);
or U2606 (N_2606,N_1815,N_1574);
xor U2607 (N_2607,N_1749,N_2225);
and U2608 (N_2608,N_1941,N_2142);
xor U2609 (N_2609,N_2195,N_2238);
and U2610 (N_2610,N_2248,N_1731);
nand U2611 (N_2611,N_2045,N_2116);
and U2612 (N_2612,N_2147,N_2010);
nor U2613 (N_2613,N_1868,N_2154);
nor U2614 (N_2614,N_1693,N_1767);
and U2615 (N_2615,N_1901,N_2095);
nor U2616 (N_2616,N_1513,N_1665);
or U2617 (N_2617,N_1975,N_2035);
nand U2618 (N_2618,N_1845,N_2139);
nor U2619 (N_2619,N_1912,N_1754);
and U2620 (N_2620,N_1918,N_1548);
or U2621 (N_2621,N_1933,N_1730);
nand U2622 (N_2622,N_1965,N_2187);
or U2623 (N_2623,N_1955,N_1695);
xnor U2624 (N_2624,N_1728,N_1940);
and U2625 (N_2625,N_1815,N_2222);
xnor U2626 (N_2626,N_2154,N_1553);
nor U2627 (N_2627,N_1592,N_2094);
xnor U2628 (N_2628,N_2082,N_1749);
and U2629 (N_2629,N_1740,N_2137);
nor U2630 (N_2630,N_1907,N_2086);
nand U2631 (N_2631,N_1941,N_1742);
xor U2632 (N_2632,N_2094,N_1638);
xnor U2633 (N_2633,N_1717,N_1657);
or U2634 (N_2634,N_2098,N_1920);
or U2635 (N_2635,N_2214,N_1876);
or U2636 (N_2636,N_1615,N_1577);
nor U2637 (N_2637,N_2249,N_1614);
or U2638 (N_2638,N_2134,N_2177);
nor U2639 (N_2639,N_1518,N_2046);
nand U2640 (N_2640,N_1586,N_1547);
nor U2641 (N_2641,N_2180,N_1573);
and U2642 (N_2642,N_2224,N_1686);
and U2643 (N_2643,N_1927,N_1716);
nor U2644 (N_2644,N_2053,N_2015);
nor U2645 (N_2645,N_2120,N_1807);
and U2646 (N_2646,N_2178,N_1591);
nand U2647 (N_2647,N_1868,N_1579);
and U2648 (N_2648,N_1925,N_1852);
xnor U2649 (N_2649,N_2220,N_1681);
nor U2650 (N_2650,N_2162,N_1573);
nor U2651 (N_2651,N_2079,N_1586);
or U2652 (N_2652,N_1669,N_1911);
nand U2653 (N_2653,N_2202,N_1512);
and U2654 (N_2654,N_2205,N_1556);
nand U2655 (N_2655,N_1669,N_1935);
and U2656 (N_2656,N_1709,N_2101);
nor U2657 (N_2657,N_1886,N_2222);
xnor U2658 (N_2658,N_1623,N_1672);
or U2659 (N_2659,N_1771,N_1683);
or U2660 (N_2660,N_1867,N_1934);
and U2661 (N_2661,N_2079,N_1836);
nor U2662 (N_2662,N_1725,N_2054);
nor U2663 (N_2663,N_1641,N_1891);
or U2664 (N_2664,N_1947,N_1780);
and U2665 (N_2665,N_2179,N_2240);
nor U2666 (N_2666,N_2004,N_1709);
and U2667 (N_2667,N_1560,N_1618);
nand U2668 (N_2668,N_2197,N_1897);
and U2669 (N_2669,N_2160,N_1681);
and U2670 (N_2670,N_1504,N_1584);
nand U2671 (N_2671,N_1863,N_1752);
and U2672 (N_2672,N_2192,N_1818);
nand U2673 (N_2673,N_1816,N_1642);
or U2674 (N_2674,N_1539,N_1880);
or U2675 (N_2675,N_2137,N_2040);
or U2676 (N_2676,N_1549,N_2081);
and U2677 (N_2677,N_1631,N_2086);
and U2678 (N_2678,N_1982,N_2061);
and U2679 (N_2679,N_2105,N_1618);
xor U2680 (N_2680,N_1552,N_2111);
nor U2681 (N_2681,N_1688,N_1944);
nand U2682 (N_2682,N_1619,N_1965);
or U2683 (N_2683,N_2091,N_2161);
nor U2684 (N_2684,N_1705,N_2209);
nand U2685 (N_2685,N_1605,N_2096);
nor U2686 (N_2686,N_2010,N_1791);
and U2687 (N_2687,N_1977,N_1525);
nand U2688 (N_2688,N_1638,N_1693);
nor U2689 (N_2689,N_1890,N_1995);
nor U2690 (N_2690,N_1805,N_2031);
nor U2691 (N_2691,N_1664,N_1832);
or U2692 (N_2692,N_1833,N_1673);
or U2693 (N_2693,N_2151,N_1665);
nor U2694 (N_2694,N_1938,N_1537);
or U2695 (N_2695,N_1604,N_1937);
nand U2696 (N_2696,N_1721,N_1565);
xor U2697 (N_2697,N_2132,N_1745);
nand U2698 (N_2698,N_1848,N_1553);
nor U2699 (N_2699,N_1503,N_1934);
or U2700 (N_2700,N_1841,N_1767);
nand U2701 (N_2701,N_1604,N_1830);
nor U2702 (N_2702,N_1801,N_1841);
xnor U2703 (N_2703,N_1773,N_1859);
nor U2704 (N_2704,N_2241,N_2197);
nand U2705 (N_2705,N_1902,N_1718);
and U2706 (N_2706,N_1724,N_2067);
or U2707 (N_2707,N_2195,N_2185);
xor U2708 (N_2708,N_1547,N_2113);
or U2709 (N_2709,N_2108,N_2015);
and U2710 (N_2710,N_2031,N_1542);
or U2711 (N_2711,N_2237,N_2159);
or U2712 (N_2712,N_1583,N_1945);
or U2713 (N_2713,N_1988,N_1550);
or U2714 (N_2714,N_2166,N_1523);
nand U2715 (N_2715,N_2209,N_2048);
nand U2716 (N_2716,N_2128,N_1754);
nand U2717 (N_2717,N_2209,N_1584);
or U2718 (N_2718,N_1629,N_1706);
and U2719 (N_2719,N_2044,N_1563);
nand U2720 (N_2720,N_1769,N_2234);
and U2721 (N_2721,N_1638,N_2246);
nor U2722 (N_2722,N_1915,N_2182);
nand U2723 (N_2723,N_2136,N_2179);
xnor U2724 (N_2724,N_1829,N_1614);
and U2725 (N_2725,N_1950,N_1942);
or U2726 (N_2726,N_1937,N_1694);
nand U2727 (N_2727,N_2172,N_2236);
and U2728 (N_2728,N_1619,N_1615);
or U2729 (N_2729,N_2180,N_1963);
and U2730 (N_2730,N_1635,N_1686);
nand U2731 (N_2731,N_2117,N_1725);
nor U2732 (N_2732,N_1871,N_1551);
or U2733 (N_2733,N_2214,N_1886);
nand U2734 (N_2734,N_1915,N_1883);
xnor U2735 (N_2735,N_1563,N_2228);
nand U2736 (N_2736,N_2067,N_1907);
nand U2737 (N_2737,N_2053,N_1800);
xor U2738 (N_2738,N_1916,N_2033);
or U2739 (N_2739,N_1690,N_2206);
nand U2740 (N_2740,N_1939,N_2172);
and U2741 (N_2741,N_1777,N_2211);
or U2742 (N_2742,N_1781,N_2201);
nand U2743 (N_2743,N_1507,N_1892);
or U2744 (N_2744,N_1528,N_2184);
nand U2745 (N_2745,N_1858,N_1946);
nand U2746 (N_2746,N_1875,N_1583);
and U2747 (N_2747,N_2228,N_1824);
xor U2748 (N_2748,N_1505,N_2035);
nand U2749 (N_2749,N_1748,N_1923);
or U2750 (N_2750,N_2133,N_1559);
nand U2751 (N_2751,N_1753,N_1880);
or U2752 (N_2752,N_1531,N_1881);
or U2753 (N_2753,N_2176,N_1562);
nand U2754 (N_2754,N_2218,N_1544);
xnor U2755 (N_2755,N_1560,N_1574);
xor U2756 (N_2756,N_1574,N_2142);
nor U2757 (N_2757,N_1856,N_2034);
and U2758 (N_2758,N_2204,N_1537);
or U2759 (N_2759,N_2162,N_1843);
nand U2760 (N_2760,N_2138,N_1718);
xnor U2761 (N_2761,N_1593,N_1848);
nor U2762 (N_2762,N_1933,N_2031);
nand U2763 (N_2763,N_1957,N_2102);
nand U2764 (N_2764,N_1652,N_1943);
and U2765 (N_2765,N_1767,N_1515);
nand U2766 (N_2766,N_1818,N_1923);
or U2767 (N_2767,N_1959,N_2026);
nand U2768 (N_2768,N_2006,N_2142);
xnor U2769 (N_2769,N_2236,N_1519);
nor U2770 (N_2770,N_1818,N_2141);
nor U2771 (N_2771,N_2020,N_1710);
and U2772 (N_2772,N_1989,N_2064);
nand U2773 (N_2773,N_2001,N_1583);
nand U2774 (N_2774,N_2155,N_2107);
nand U2775 (N_2775,N_1857,N_1598);
and U2776 (N_2776,N_1710,N_2043);
nand U2777 (N_2777,N_2106,N_2207);
nand U2778 (N_2778,N_1892,N_2136);
or U2779 (N_2779,N_1647,N_1632);
nor U2780 (N_2780,N_2148,N_1545);
xnor U2781 (N_2781,N_1721,N_2179);
and U2782 (N_2782,N_1965,N_1892);
nor U2783 (N_2783,N_1599,N_1682);
or U2784 (N_2784,N_1545,N_1710);
or U2785 (N_2785,N_1595,N_1614);
nand U2786 (N_2786,N_1954,N_1627);
nand U2787 (N_2787,N_2140,N_1895);
or U2788 (N_2788,N_1706,N_1659);
or U2789 (N_2789,N_1717,N_1757);
and U2790 (N_2790,N_1594,N_1711);
nor U2791 (N_2791,N_1869,N_1897);
and U2792 (N_2792,N_1922,N_2246);
and U2793 (N_2793,N_2021,N_1736);
nand U2794 (N_2794,N_1809,N_1527);
or U2795 (N_2795,N_1740,N_1707);
nand U2796 (N_2796,N_2171,N_2164);
or U2797 (N_2797,N_1540,N_1669);
and U2798 (N_2798,N_1575,N_1865);
xnor U2799 (N_2799,N_2079,N_1855);
xnor U2800 (N_2800,N_1540,N_2141);
nand U2801 (N_2801,N_2140,N_2134);
and U2802 (N_2802,N_2212,N_1644);
and U2803 (N_2803,N_2221,N_2169);
nor U2804 (N_2804,N_1662,N_2182);
and U2805 (N_2805,N_2201,N_2235);
nor U2806 (N_2806,N_1568,N_1947);
nor U2807 (N_2807,N_1794,N_1887);
or U2808 (N_2808,N_1765,N_2040);
nor U2809 (N_2809,N_1713,N_1748);
xnor U2810 (N_2810,N_1853,N_1881);
and U2811 (N_2811,N_2142,N_2123);
nand U2812 (N_2812,N_1776,N_1629);
or U2813 (N_2813,N_1847,N_1694);
nand U2814 (N_2814,N_2113,N_2066);
and U2815 (N_2815,N_1804,N_1571);
nor U2816 (N_2816,N_1870,N_1824);
nand U2817 (N_2817,N_1872,N_1731);
and U2818 (N_2818,N_2024,N_2134);
nor U2819 (N_2819,N_2205,N_2102);
or U2820 (N_2820,N_1535,N_1892);
and U2821 (N_2821,N_2169,N_2061);
nand U2822 (N_2822,N_1819,N_1597);
and U2823 (N_2823,N_2067,N_1628);
nor U2824 (N_2824,N_1788,N_1737);
nor U2825 (N_2825,N_1946,N_1925);
or U2826 (N_2826,N_2030,N_1734);
and U2827 (N_2827,N_1663,N_1861);
nor U2828 (N_2828,N_1988,N_2136);
nand U2829 (N_2829,N_1550,N_2138);
and U2830 (N_2830,N_1652,N_2069);
xnor U2831 (N_2831,N_1868,N_2106);
and U2832 (N_2832,N_1628,N_1612);
and U2833 (N_2833,N_2073,N_1687);
xor U2834 (N_2834,N_1850,N_1883);
or U2835 (N_2835,N_1741,N_2169);
and U2836 (N_2836,N_1657,N_1528);
nand U2837 (N_2837,N_1873,N_2043);
nand U2838 (N_2838,N_1867,N_1568);
and U2839 (N_2839,N_1867,N_1647);
or U2840 (N_2840,N_1901,N_1692);
nand U2841 (N_2841,N_1712,N_2172);
nor U2842 (N_2842,N_1890,N_2224);
nor U2843 (N_2843,N_1731,N_2048);
nand U2844 (N_2844,N_2077,N_1595);
nor U2845 (N_2845,N_1701,N_1828);
xnor U2846 (N_2846,N_2138,N_1554);
nor U2847 (N_2847,N_1897,N_1958);
or U2848 (N_2848,N_1895,N_2160);
and U2849 (N_2849,N_1809,N_1760);
and U2850 (N_2850,N_1520,N_2013);
and U2851 (N_2851,N_2167,N_1776);
and U2852 (N_2852,N_1898,N_1757);
nor U2853 (N_2853,N_2142,N_1505);
nand U2854 (N_2854,N_1815,N_2237);
and U2855 (N_2855,N_2102,N_2198);
nand U2856 (N_2856,N_2170,N_2032);
and U2857 (N_2857,N_1929,N_2118);
and U2858 (N_2858,N_2235,N_2066);
and U2859 (N_2859,N_2216,N_1838);
nor U2860 (N_2860,N_1975,N_1563);
nor U2861 (N_2861,N_1717,N_1834);
nand U2862 (N_2862,N_1784,N_1989);
nand U2863 (N_2863,N_1699,N_2161);
or U2864 (N_2864,N_1900,N_1872);
xnor U2865 (N_2865,N_2029,N_1535);
nand U2866 (N_2866,N_2015,N_1929);
or U2867 (N_2867,N_2190,N_1972);
xnor U2868 (N_2868,N_1950,N_1898);
and U2869 (N_2869,N_1745,N_1974);
and U2870 (N_2870,N_1716,N_1755);
or U2871 (N_2871,N_1890,N_1765);
or U2872 (N_2872,N_2106,N_1561);
and U2873 (N_2873,N_1615,N_2216);
or U2874 (N_2874,N_1651,N_1745);
nor U2875 (N_2875,N_2034,N_1638);
nor U2876 (N_2876,N_2192,N_1965);
nand U2877 (N_2877,N_1526,N_1833);
or U2878 (N_2878,N_1716,N_1977);
and U2879 (N_2879,N_1610,N_2213);
xor U2880 (N_2880,N_1960,N_2204);
and U2881 (N_2881,N_2220,N_2175);
nor U2882 (N_2882,N_2064,N_1502);
nand U2883 (N_2883,N_2239,N_1998);
xor U2884 (N_2884,N_1503,N_2056);
nor U2885 (N_2885,N_1931,N_2207);
or U2886 (N_2886,N_2043,N_1647);
nand U2887 (N_2887,N_1975,N_2031);
nand U2888 (N_2888,N_1624,N_1801);
nand U2889 (N_2889,N_1909,N_2220);
nor U2890 (N_2890,N_1590,N_2181);
nor U2891 (N_2891,N_1525,N_1570);
nor U2892 (N_2892,N_1624,N_1733);
or U2893 (N_2893,N_2013,N_2225);
xnor U2894 (N_2894,N_2234,N_1889);
nor U2895 (N_2895,N_2225,N_2156);
and U2896 (N_2896,N_2219,N_1550);
nand U2897 (N_2897,N_1730,N_1823);
nand U2898 (N_2898,N_1697,N_1751);
xor U2899 (N_2899,N_1824,N_1732);
nor U2900 (N_2900,N_1808,N_2081);
or U2901 (N_2901,N_2121,N_1617);
or U2902 (N_2902,N_1500,N_2105);
nand U2903 (N_2903,N_1527,N_2081);
nand U2904 (N_2904,N_1935,N_1801);
nand U2905 (N_2905,N_1664,N_1927);
xor U2906 (N_2906,N_2023,N_2129);
nor U2907 (N_2907,N_1610,N_1817);
and U2908 (N_2908,N_2246,N_1519);
and U2909 (N_2909,N_1712,N_1858);
nor U2910 (N_2910,N_1771,N_1869);
and U2911 (N_2911,N_1627,N_1600);
xor U2912 (N_2912,N_1513,N_2010);
nor U2913 (N_2913,N_1826,N_1861);
nor U2914 (N_2914,N_1912,N_1826);
nor U2915 (N_2915,N_2019,N_2151);
nor U2916 (N_2916,N_1980,N_1695);
and U2917 (N_2917,N_1607,N_1765);
nor U2918 (N_2918,N_1810,N_1610);
or U2919 (N_2919,N_2233,N_1520);
or U2920 (N_2920,N_1685,N_1933);
and U2921 (N_2921,N_1757,N_1997);
and U2922 (N_2922,N_1942,N_2014);
or U2923 (N_2923,N_1848,N_1787);
and U2924 (N_2924,N_1713,N_1743);
nor U2925 (N_2925,N_2240,N_1853);
nor U2926 (N_2926,N_2096,N_1912);
nand U2927 (N_2927,N_1652,N_2156);
xor U2928 (N_2928,N_1568,N_1681);
and U2929 (N_2929,N_1842,N_1549);
nor U2930 (N_2930,N_2245,N_1802);
and U2931 (N_2931,N_1573,N_2224);
nand U2932 (N_2932,N_1634,N_1560);
or U2933 (N_2933,N_1553,N_1507);
nor U2934 (N_2934,N_1556,N_1861);
and U2935 (N_2935,N_1838,N_2080);
nor U2936 (N_2936,N_1660,N_1931);
and U2937 (N_2937,N_1624,N_1872);
xor U2938 (N_2938,N_1550,N_2032);
and U2939 (N_2939,N_2002,N_2187);
or U2940 (N_2940,N_2222,N_2185);
or U2941 (N_2941,N_1522,N_2173);
nor U2942 (N_2942,N_2128,N_2038);
or U2943 (N_2943,N_2068,N_1766);
or U2944 (N_2944,N_2228,N_1764);
or U2945 (N_2945,N_2012,N_1602);
nor U2946 (N_2946,N_2000,N_2232);
nand U2947 (N_2947,N_2173,N_2145);
and U2948 (N_2948,N_1563,N_1715);
xnor U2949 (N_2949,N_2213,N_2203);
nor U2950 (N_2950,N_1616,N_1738);
nor U2951 (N_2951,N_2006,N_2081);
nor U2952 (N_2952,N_2142,N_1779);
nor U2953 (N_2953,N_1955,N_2161);
nor U2954 (N_2954,N_1874,N_1708);
and U2955 (N_2955,N_2224,N_1703);
or U2956 (N_2956,N_1515,N_1724);
nand U2957 (N_2957,N_1902,N_2011);
or U2958 (N_2958,N_1734,N_1736);
nand U2959 (N_2959,N_2112,N_1737);
nand U2960 (N_2960,N_1720,N_2195);
or U2961 (N_2961,N_1948,N_2026);
or U2962 (N_2962,N_1796,N_2097);
or U2963 (N_2963,N_1556,N_1928);
xnor U2964 (N_2964,N_2028,N_2113);
nor U2965 (N_2965,N_2202,N_2119);
or U2966 (N_2966,N_1902,N_2017);
nor U2967 (N_2967,N_1907,N_2115);
or U2968 (N_2968,N_1708,N_1929);
and U2969 (N_2969,N_2075,N_1855);
and U2970 (N_2970,N_1973,N_1736);
or U2971 (N_2971,N_2215,N_1972);
xnor U2972 (N_2972,N_1725,N_1747);
xnor U2973 (N_2973,N_1973,N_2095);
and U2974 (N_2974,N_1763,N_2185);
or U2975 (N_2975,N_1989,N_1958);
nand U2976 (N_2976,N_2060,N_1950);
xnor U2977 (N_2977,N_1796,N_1640);
nand U2978 (N_2978,N_1716,N_2101);
nor U2979 (N_2979,N_2063,N_1783);
or U2980 (N_2980,N_1858,N_1535);
or U2981 (N_2981,N_1647,N_1543);
and U2982 (N_2982,N_1757,N_1747);
and U2983 (N_2983,N_1663,N_1908);
or U2984 (N_2984,N_2242,N_2017);
nand U2985 (N_2985,N_1803,N_1554);
and U2986 (N_2986,N_1704,N_1573);
nand U2987 (N_2987,N_2184,N_1885);
and U2988 (N_2988,N_1766,N_1543);
nand U2989 (N_2989,N_1686,N_1937);
or U2990 (N_2990,N_1696,N_1720);
and U2991 (N_2991,N_1884,N_2152);
or U2992 (N_2992,N_2165,N_1671);
nand U2993 (N_2993,N_2040,N_2220);
or U2994 (N_2994,N_1684,N_1965);
and U2995 (N_2995,N_1737,N_2115);
or U2996 (N_2996,N_1644,N_1659);
nand U2997 (N_2997,N_1969,N_1844);
nand U2998 (N_2998,N_1589,N_1764);
nor U2999 (N_2999,N_1885,N_2036);
nand U3000 (N_3000,N_2304,N_2776);
nand U3001 (N_3001,N_2489,N_2950);
or U3002 (N_3002,N_2826,N_2696);
nor U3003 (N_3003,N_2428,N_2889);
and U3004 (N_3004,N_2447,N_2453);
or U3005 (N_3005,N_2600,N_2700);
nor U3006 (N_3006,N_2669,N_2295);
xnor U3007 (N_3007,N_2260,N_2637);
nor U3008 (N_3008,N_2909,N_2482);
nor U3009 (N_3009,N_2467,N_2866);
nand U3010 (N_3010,N_2606,N_2317);
or U3011 (N_3011,N_2426,N_2855);
nand U3012 (N_3012,N_2901,N_2570);
and U3013 (N_3013,N_2661,N_2346);
and U3014 (N_3014,N_2995,N_2778);
nor U3015 (N_3015,N_2290,N_2664);
xnor U3016 (N_3016,N_2843,N_2974);
or U3017 (N_3017,N_2867,N_2477);
nor U3018 (N_3018,N_2964,N_2398);
xor U3019 (N_3019,N_2734,N_2391);
nand U3020 (N_3020,N_2438,N_2801);
or U3021 (N_3021,N_2720,N_2299);
and U3022 (N_3022,N_2535,N_2825);
xnor U3023 (N_3023,N_2937,N_2797);
nand U3024 (N_3024,N_2455,N_2989);
and U3025 (N_3025,N_2717,N_2803);
nor U3026 (N_3026,N_2279,N_2822);
or U3027 (N_3027,N_2832,N_2422);
nor U3028 (N_3028,N_2993,N_2860);
nor U3029 (N_3029,N_2774,N_2283);
xor U3030 (N_3030,N_2508,N_2417);
or U3031 (N_3031,N_2620,N_2973);
nand U3032 (N_3032,N_2448,N_2367);
nand U3033 (N_3033,N_2436,N_2285);
or U3034 (N_3034,N_2492,N_2543);
nor U3035 (N_3035,N_2882,N_2737);
nor U3036 (N_3036,N_2975,N_2782);
nor U3037 (N_3037,N_2705,N_2357);
nor U3038 (N_3038,N_2938,N_2271);
and U3039 (N_3039,N_2847,N_2445);
xor U3040 (N_3040,N_2597,N_2651);
nand U3041 (N_3041,N_2565,N_2942);
or U3042 (N_3042,N_2821,N_2377);
xnor U3043 (N_3043,N_2786,N_2890);
or U3044 (N_3044,N_2320,N_2675);
or U3045 (N_3045,N_2525,N_2931);
and U3046 (N_3046,N_2878,N_2442);
or U3047 (N_3047,N_2614,N_2439);
or U3048 (N_3048,N_2491,N_2310);
nor U3049 (N_3049,N_2864,N_2941);
nand U3050 (N_3050,N_2899,N_2433);
nor U3051 (N_3051,N_2642,N_2876);
nand U3052 (N_3052,N_2587,N_2735);
xor U3053 (N_3053,N_2400,N_2714);
and U3054 (N_3054,N_2785,N_2567);
xnor U3055 (N_3055,N_2356,N_2753);
or U3056 (N_3056,N_2990,N_2951);
and U3057 (N_3057,N_2498,N_2384);
nand U3058 (N_3058,N_2392,N_2738);
xnor U3059 (N_3059,N_2721,N_2683);
nand U3060 (N_3060,N_2773,N_2898);
nor U3061 (N_3061,N_2731,N_2934);
and U3062 (N_3062,N_2560,N_2680);
nor U3063 (N_3063,N_2393,N_2814);
nor U3064 (N_3064,N_2596,N_2744);
or U3065 (N_3065,N_2517,N_2634);
or U3066 (N_3066,N_2590,N_2454);
nor U3067 (N_3067,N_2531,N_2338);
nand U3068 (N_3068,N_2799,N_2854);
and U3069 (N_3069,N_2981,N_2910);
and U3070 (N_3070,N_2547,N_2834);
nand U3071 (N_3071,N_2791,N_2552);
or U3072 (N_3072,N_2293,N_2354);
and U3073 (N_3073,N_2630,N_2336);
and U3074 (N_3074,N_2330,N_2345);
and U3075 (N_3075,N_2471,N_2877);
nor U3076 (N_3076,N_2968,N_2674);
nor U3077 (N_3077,N_2595,N_2965);
xor U3078 (N_3078,N_2533,N_2324);
nand U3079 (N_3079,N_2564,N_2385);
nor U3080 (N_3080,N_2879,N_2494);
nand U3081 (N_3081,N_2390,N_2263);
or U3082 (N_3082,N_2611,N_2274);
or U3083 (N_3083,N_2311,N_2955);
nand U3084 (N_3084,N_2906,N_2677);
nor U3085 (N_3085,N_2430,N_2539);
xor U3086 (N_3086,N_2687,N_2852);
or U3087 (N_3087,N_2657,N_2796);
nand U3088 (N_3088,N_2710,N_2413);
nand U3089 (N_3089,N_2730,N_2980);
and U3090 (N_3090,N_2399,N_2256);
xnor U3091 (N_3091,N_2419,N_2551);
and U3092 (N_3092,N_2459,N_2591);
or U3093 (N_3093,N_2312,N_2586);
nor U3094 (N_3094,N_2521,N_2954);
nand U3095 (N_3095,N_2402,N_2513);
nor U3096 (N_3096,N_2575,N_2309);
nor U3097 (N_3097,N_2523,N_2837);
and U3098 (N_3098,N_2308,N_2701);
nand U3099 (N_3099,N_2540,N_2986);
nor U3100 (N_3100,N_2457,N_2431);
nand U3101 (N_3101,N_2380,N_2631);
nand U3102 (N_3102,N_2418,N_2808);
nor U3103 (N_3103,N_2662,N_2992);
and U3104 (N_3104,N_2755,N_2999);
nand U3105 (N_3105,N_2649,N_2887);
nand U3106 (N_3106,N_2758,N_2421);
or U3107 (N_3107,N_2365,N_2676);
and U3108 (N_3108,N_2613,N_2281);
nand U3109 (N_3109,N_2555,N_2793);
or U3110 (N_3110,N_2895,N_2646);
nor U3111 (N_3111,N_2915,N_2949);
and U3112 (N_3112,N_2255,N_2893);
xnor U3113 (N_3113,N_2819,N_2914);
or U3114 (N_3114,N_2952,N_2333);
or U3115 (N_3115,N_2722,N_2960);
nor U3116 (N_3116,N_2351,N_2561);
and U3117 (N_3117,N_2994,N_2538);
or U3118 (N_3118,N_2764,N_2405);
and U3119 (N_3119,N_2542,N_2569);
nor U3120 (N_3120,N_2483,N_2660);
nor U3121 (N_3121,N_2379,N_2788);
or U3122 (N_3122,N_2881,N_2568);
nand U3123 (N_3123,N_2865,N_2956);
or U3124 (N_3124,N_2655,N_2532);
nor U3125 (N_3125,N_2766,N_2451);
and U3126 (N_3126,N_2982,N_2997);
nand U3127 (N_3127,N_2362,N_2603);
or U3128 (N_3128,N_2315,N_2548);
or U3129 (N_3129,N_2516,N_2850);
and U3130 (N_3130,N_2472,N_2610);
and U3131 (N_3131,N_2647,N_2967);
nor U3132 (N_3132,N_2358,N_2724);
and U3133 (N_3133,N_2728,N_2327);
nor U3134 (N_3134,N_2976,N_2301);
nand U3135 (N_3135,N_2894,N_2804);
nor U3136 (N_3136,N_2427,N_2971);
nand U3137 (N_3137,N_2395,N_2874);
xor U3138 (N_3138,N_2578,N_2623);
nor U3139 (N_3139,N_2605,N_2679);
xnor U3140 (N_3140,N_2820,N_2585);
xnor U3141 (N_3141,N_2337,N_2780);
xnor U3142 (N_3142,N_2562,N_2886);
xor U3143 (N_3143,N_2468,N_2440);
or U3144 (N_3144,N_2715,N_2618);
nand U3145 (N_3145,N_2607,N_2497);
nand U3146 (N_3146,N_2269,N_2718);
xor U3147 (N_3147,N_2505,N_2828);
nor U3148 (N_3148,N_2340,N_2353);
or U3149 (N_3149,N_2948,N_2287);
or U3150 (N_3150,N_2707,N_2708);
xor U3151 (N_3151,N_2411,N_2963);
nand U3152 (N_3152,N_2318,N_2946);
nand U3153 (N_3153,N_2795,N_2783);
nor U3154 (N_3154,N_2781,N_2643);
xnor U3155 (N_3155,N_2692,N_2806);
and U3156 (N_3156,N_2550,N_2593);
or U3157 (N_3157,N_2348,N_2888);
nor U3158 (N_3158,N_2479,N_2838);
nand U3159 (N_3159,N_2686,N_2500);
and U3160 (N_3160,N_2370,N_2487);
nand U3161 (N_3161,N_2302,N_2342);
nand U3162 (N_3162,N_2920,N_2969);
and U3163 (N_3163,N_2601,N_2944);
nor U3164 (N_3164,N_2933,N_2917);
nand U3165 (N_3165,N_2652,N_2475);
nand U3166 (N_3166,N_2784,N_2831);
nor U3167 (N_3167,N_2689,N_2856);
nand U3168 (N_3168,N_2699,N_2844);
or U3169 (N_3169,N_2979,N_2251);
nand U3170 (N_3170,N_2485,N_2469);
xor U3171 (N_3171,N_2464,N_2711);
nor U3172 (N_3172,N_2761,N_2684);
or U3173 (N_3173,N_2849,N_2493);
nor U3174 (N_3174,N_2507,N_2627);
or U3175 (N_3175,N_2522,N_2815);
or U3176 (N_3176,N_2703,N_2970);
nand U3177 (N_3177,N_2861,N_2863);
nor U3178 (N_3178,N_2266,N_2261);
or U3179 (N_3179,N_2463,N_2347);
or U3180 (N_3180,N_2499,N_2919);
nand U3181 (N_3181,N_2732,N_2510);
nand U3182 (N_3182,N_2387,N_2300);
nor U3183 (N_3183,N_2885,N_2672);
nor U3184 (N_3184,N_2818,N_2667);
or U3185 (N_3185,N_2388,N_2871);
nor U3186 (N_3186,N_2297,N_2374);
nor U3187 (N_3187,N_2742,N_2292);
xnor U3188 (N_3188,N_2404,N_2836);
or U3189 (N_3189,N_2389,N_2289);
xor U3190 (N_3190,N_2918,N_2811);
nor U3191 (N_3191,N_2905,N_2759);
xor U3192 (N_3192,N_2927,N_2534);
nand U3193 (N_3193,N_2577,N_2789);
and U3194 (N_3194,N_2966,N_2685);
or U3195 (N_3195,N_2739,N_2695);
nand U3196 (N_3196,N_2829,N_2681);
or U3197 (N_3197,N_2458,N_2698);
xnor U3198 (N_3198,N_2410,N_2432);
nor U3199 (N_3199,N_2644,N_2288);
or U3200 (N_3200,N_2896,N_2368);
and U3201 (N_3201,N_2653,N_2749);
xor U3202 (N_3202,N_2277,N_2977);
nor U3203 (N_3203,N_2792,N_2394);
nand U3204 (N_3204,N_2371,N_2305);
and U3205 (N_3205,N_2619,N_2682);
nand U3206 (N_3206,N_2633,N_2823);
nand U3207 (N_3207,N_2845,N_2363);
xor U3208 (N_3208,N_2923,N_2557);
and U3209 (N_3209,N_2434,N_2713);
nand U3210 (N_3210,N_2252,N_2412);
or U3211 (N_3211,N_2827,N_2361);
nand U3212 (N_3212,N_2908,N_2880);
nor U3213 (N_3213,N_2943,N_2840);
xor U3214 (N_3214,N_2663,N_2546);
or U3215 (N_3215,N_2461,N_2873);
nor U3216 (N_3216,N_2648,N_2930);
and U3217 (N_3217,N_2519,N_2763);
nand U3218 (N_3218,N_2736,N_2268);
xor U3219 (N_3219,N_2284,N_2907);
nor U3220 (N_3220,N_2449,N_2706);
nor U3221 (N_3221,N_2996,N_2359);
nor U3222 (N_3222,N_2884,N_2563);
nor U3223 (N_3223,N_2857,N_2429);
or U3224 (N_3224,N_2892,N_2868);
nand U3225 (N_3225,N_2509,N_2869);
nor U3226 (N_3226,N_2258,N_2328);
or U3227 (N_3227,N_2262,N_2645);
nor U3228 (N_3228,N_2903,N_2306);
nand U3229 (N_3229,N_2512,N_2959);
nor U3230 (N_3230,N_2846,N_2924);
and U3231 (N_3231,N_2665,N_2545);
and U3232 (N_3232,N_2729,N_2875);
or U3233 (N_3233,N_2291,N_2303);
nor U3234 (N_3234,N_2900,N_2922);
or U3235 (N_3235,N_2382,N_2702);
nor U3236 (N_3236,N_2423,N_2566);
nand U3237 (N_3237,N_2574,N_2501);
nor U3238 (N_3238,N_2641,N_2372);
or U3239 (N_3239,N_2556,N_2929);
nor U3240 (N_3240,N_2771,N_2940);
and U3241 (N_3241,N_2571,N_2511);
or U3242 (N_3242,N_2343,N_2957);
nor U3243 (N_3243,N_2858,N_2848);
and U3244 (N_3244,N_2656,N_2527);
nor U3245 (N_3245,N_2916,N_2790);
or U3246 (N_3246,N_2958,N_2381);
nand U3247 (N_3247,N_2465,N_2747);
nand U3248 (N_3248,N_2444,N_2622);
nor U3249 (N_3249,N_2670,N_2580);
or U3250 (N_3250,N_2553,N_2396);
nor U3251 (N_3251,N_2925,N_2765);
nor U3252 (N_3252,N_2639,N_2767);
xnor U3253 (N_3253,N_2750,N_2452);
or U3254 (N_3254,N_2748,N_2369);
nor U3255 (N_3255,N_2425,N_2339);
and U3256 (N_3256,N_2988,N_2488);
nand U3257 (N_3257,N_2514,N_2375);
nand U3258 (N_3258,N_2688,N_2830);
nor U3259 (N_3259,N_2816,N_2480);
and U3260 (N_3260,N_2344,N_2842);
or U3261 (N_3261,N_2629,N_2697);
or U3262 (N_3262,N_2625,N_2267);
nor U3263 (N_3263,N_2529,N_2579);
and U3264 (N_3264,N_2298,N_2294);
nor U3265 (N_3265,N_2953,N_2280);
or U3266 (N_3266,N_2802,N_2588);
xnor U3267 (N_3267,N_2859,N_2594);
nand U3268 (N_3268,N_2787,N_2559);
and U3269 (N_3269,N_2544,N_2466);
xor U3270 (N_3270,N_2528,N_2694);
and U3271 (N_3271,N_2599,N_2709);
and U3272 (N_3272,N_2987,N_2407);
nand U3273 (N_3273,N_2321,N_2817);
nand U3274 (N_3274,N_2504,N_2350);
xnor U3275 (N_3275,N_2666,N_2604);
and U3276 (N_3276,N_2460,N_2450);
nand U3277 (N_3277,N_2424,N_2862);
or U3278 (N_3278,N_2360,N_2264);
nand U3279 (N_3279,N_2441,N_2470);
nand U3280 (N_3280,N_2636,N_2671);
nand U3281 (N_3281,N_2364,N_2926);
or U3282 (N_3282,N_2257,N_2592);
nor U3283 (N_3283,N_2608,N_2366);
nor U3284 (N_3284,N_2443,N_2406);
xnor U3285 (N_3285,N_2853,N_2276);
and U3286 (N_3286,N_2921,N_2332);
nand U3287 (N_3287,N_2355,N_2904);
nor U3288 (N_3288,N_2397,N_2420);
and U3289 (N_3289,N_2573,N_2998);
or U3290 (N_3290,N_2537,N_2770);
nor U3291 (N_3291,N_2481,N_2602);
or U3292 (N_3292,N_2496,N_2668);
and U3293 (N_3293,N_2978,N_2704);
nor U3294 (N_3294,N_2401,N_2947);
and U3295 (N_3295,N_2983,N_2913);
nand U3296 (N_3296,N_2270,N_2549);
nor U3297 (N_3297,N_2326,N_2807);
or U3298 (N_3298,N_2476,N_2741);
nor U3299 (N_3299,N_2473,N_2762);
nor U3300 (N_3300,N_2530,N_2751);
nand U3301 (N_3301,N_2833,N_2416);
nor U3302 (N_3302,N_2581,N_2726);
nor U3303 (N_3303,N_2754,N_2349);
xnor U3304 (N_3304,N_2414,N_2628);
or U3305 (N_3305,N_2779,N_2911);
nor U3306 (N_3306,N_2912,N_2250);
and U3307 (N_3307,N_2809,N_2812);
nor U3308 (N_3308,N_2712,N_2939);
or U3309 (N_3309,N_2462,N_2278);
nand U3310 (N_3310,N_2386,N_2640);
nor U3311 (N_3311,N_2598,N_2589);
and U3312 (N_3312,N_2659,N_2282);
nand U3313 (N_3313,N_2841,N_2824);
nor U3314 (N_3314,N_2484,N_2961);
or U3315 (N_3315,N_2690,N_2678);
xor U3316 (N_3316,N_2632,N_2638);
nor U3317 (N_3317,N_2518,N_2673);
and U3318 (N_3318,N_2502,N_2446);
xnor U3319 (N_3319,N_2408,N_2409);
nand U3320 (N_3320,N_2932,N_2746);
xor U3321 (N_3321,N_2733,N_2936);
nand U3322 (N_3322,N_2658,N_2621);
nor U3323 (N_3323,N_2945,N_2506);
xnor U3324 (N_3324,N_2985,N_2928);
nor U3325 (N_3325,N_2839,N_2768);
nor U3326 (N_3326,N_2772,N_2296);
or U3327 (N_3327,N_2962,N_2609);
nand U3328 (N_3328,N_2743,N_2329);
nor U3329 (N_3329,N_2272,N_2756);
nor U3330 (N_3330,N_2319,N_2800);
and U3331 (N_3331,N_2495,N_2275);
or U3332 (N_3332,N_2835,N_2810);
or U3333 (N_3333,N_2341,N_2383);
nand U3334 (N_3334,N_2752,N_2322);
and U3335 (N_3335,N_2617,N_2725);
xnor U3336 (N_3336,N_2972,N_2654);
and U3337 (N_3337,N_2757,N_2456);
nor U3338 (N_3338,N_2984,N_2719);
nor U3339 (N_3339,N_2870,N_2259);
or U3340 (N_3340,N_2478,N_2760);
or U3341 (N_3341,N_2584,N_2554);
and U3342 (N_3342,N_2745,N_2435);
nor U3343 (N_3343,N_2897,N_2805);
nor U3344 (N_3344,N_2798,N_2883);
and U3345 (N_3345,N_2253,N_2524);
nor U3346 (N_3346,N_2872,N_2254);
nor U3347 (N_3347,N_2307,N_2851);
and U3348 (N_3348,N_2378,N_2991);
or U3349 (N_3349,N_2313,N_2769);
nor U3350 (N_3350,N_2891,N_2526);
nand U3351 (N_3351,N_2520,N_2813);
nor U3352 (N_3352,N_2740,N_2777);
and U3353 (N_3353,N_2624,N_2536);
nand U3354 (N_3354,N_2572,N_2582);
nor U3355 (N_3355,N_2314,N_2273);
nand U3356 (N_3356,N_2286,N_2265);
nand U3357 (N_3357,N_2376,N_2352);
and U3358 (N_3358,N_2723,N_2437);
xor U3359 (N_3359,N_2541,N_2331);
and U3360 (N_3360,N_2935,N_2727);
nand U3361 (N_3361,N_2615,N_2316);
or U3362 (N_3362,N_2323,N_2635);
and U3363 (N_3363,N_2503,N_2335);
nor U3364 (N_3364,N_2576,N_2415);
xnor U3365 (N_3365,N_2515,N_2794);
xor U3366 (N_3366,N_2403,N_2334);
nand U3367 (N_3367,N_2583,N_2716);
and U3368 (N_3368,N_2486,N_2612);
nor U3369 (N_3369,N_2902,N_2650);
nor U3370 (N_3370,N_2325,N_2474);
nor U3371 (N_3371,N_2691,N_2693);
nor U3372 (N_3372,N_2373,N_2616);
nor U3373 (N_3373,N_2626,N_2490);
nand U3374 (N_3374,N_2775,N_2558);
or U3375 (N_3375,N_2528,N_2453);
and U3376 (N_3376,N_2693,N_2787);
or U3377 (N_3377,N_2321,N_2252);
xnor U3378 (N_3378,N_2661,N_2833);
or U3379 (N_3379,N_2809,N_2369);
and U3380 (N_3380,N_2378,N_2455);
nand U3381 (N_3381,N_2773,N_2965);
or U3382 (N_3382,N_2412,N_2527);
or U3383 (N_3383,N_2316,N_2279);
or U3384 (N_3384,N_2967,N_2334);
or U3385 (N_3385,N_2307,N_2555);
nand U3386 (N_3386,N_2872,N_2439);
nand U3387 (N_3387,N_2265,N_2998);
nor U3388 (N_3388,N_2383,N_2856);
or U3389 (N_3389,N_2826,N_2422);
nor U3390 (N_3390,N_2410,N_2770);
nor U3391 (N_3391,N_2700,N_2530);
or U3392 (N_3392,N_2799,N_2389);
and U3393 (N_3393,N_2739,N_2742);
and U3394 (N_3394,N_2275,N_2436);
xnor U3395 (N_3395,N_2987,N_2504);
xnor U3396 (N_3396,N_2969,N_2607);
and U3397 (N_3397,N_2989,N_2848);
or U3398 (N_3398,N_2939,N_2644);
nor U3399 (N_3399,N_2692,N_2705);
nor U3400 (N_3400,N_2729,N_2418);
or U3401 (N_3401,N_2977,N_2323);
nand U3402 (N_3402,N_2448,N_2757);
or U3403 (N_3403,N_2556,N_2597);
nand U3404 (N_3404,N_2385,N_2859);
nand U3405 (N_3405,N_2800,N_2513);
xor U3406 (N_3406,N_2623,N_2895);
and U3407 (N_3407,N_2813,N_2654);
and U3408 (N_3408,N_2669,N_2316);
nor U3409 (N_3409,N_2635,N_2925);
and U3410 (N_3410,N_2948,N_2872);
or U3411 (N_3411,N_2797,N_2252);
and U3412 (N_3412,N_2735,N_2706);
nand U3413 (N_3413,N_2845,N_2730);
and U3414 (N_3414,N_2742,N_2492);
and U3415 (N_3415,N_2641,N_2538);
or U3416 (N_3416,N_2687,N_2963);
nor U3417 (N_3417,N_2788,N_2863);
and U3418 (N_3418,N_2971,N_2285);
nand U3419 (N_3419,N_2958,N_2440);
nor U3420 (N_3420,N_2920,N_2992);
xnor U3421 (N_3421,N_2472,N_2502);
or U3422 (N_3422,N_2845,N_2360);
nor U3423 (N_3423,N_2556,N_2457);
and U3424 (N_3424,N_2283,N_2980);
nor U3425 (N_3425,N_2730,N_2975);
nor U3426 (N_3426,N_2940,N_2407);
nor U3427 (N_3427,N_2742,N_2418);
nand U3428 (N_3428,N_2622,N_2327);
or U3429 (N_3429,N_2871,N_2255);
and U3430 (N_3430,N_2278,N_2528);
or U3431 (N_3431,N_2435,N_2710);
or U3432 (N_3432,N_2775,N_2766);
nor U3433 (N_3433,N_2542,N_2952);
xor U3434 (N_3434,N_2442,N_2503);
or U3435 (N_3435,N_2799,N_2969);
and U3436 (N_3436,N_2627,N_2500);
nand U3437 (N_3437,N_2623,N_2547);
nand U3438 (N_3438,N_2523,N_2933);
nand U3439 (N_3439,N_2399,N_2448);
nand U3440 (N_3440,N_2366,N_2353);
nand U3441 (N_3441,N_2933,N_2851);
and U3442 (N_3442,N_2379,N_2281);
nor U3443 (N_3443,N_2867,N_2543);
nand U3444 (N_3444,N_2703,N_2995);
nand U3445 (N_3445,N_2553,N_2475);
and U3446 (N_3446,N_2345,N_2669);
nand U3447 (N_3447,N_2290,N_2951);
xnor U3448 (N_3448,N_2862,N_2439);
nand U3449 (N_3449,N_2525,N_2567);
nor U3450 (N_3450,N_2915,N_2582);
nand U3451 (N_3451,N_2500,N_2662);
xnor U3452 (N_3452,N_2359,N_2586);
nor U3453 (N_3453,N_2296,N_2873);
nand U3454 (N_3454,N_2456,N_2955);
nand U3455 (N_3455,N_2481,N_2393);
nand U3456 (N_3456,N_2960,N_2900);
or U3457 (N_3457,N_2707,N_2343);
or U3458 (N_3458,N_2275,N_2501);
or U3459 (N_3459,N_2877,N_2984);
nand U3460 (N_3460,N_2256,N_2829);
nand U3461 (N_3461,N_2384,N_2912);
nor U3462 (N_3462,N_2856,N_2394);
nand U3463 (N_3463,N_2372,N_2477);
nand U3464 (N_3464,N_2274,N_2319);
and U3465 (N_3465,N_2975,N_2529);
or U3466 (N_3466,N_2942,N_2934);
nor U3467 (N_3467,N_2901,N_2981);
nor U3468 (N_3468,N_2964,N_2972);
and U3469 (N_3469,N_2618,N_2419);
and U3470 (N_3470,N_2473,N_2402);
xnor U3471 (N_3471,N_2339,N_2508);
and U3472 (N_3472,N_2465,N_2819);
and U3473 (N_3473,N_2868,N_2656);
or U3474 (N_3474,N_2933,N_2939);
and U3475 (N_3475,N_2274,N_2971);
and U3476 (N_3476,N_2728,N_2367);
nand U3477 (N_3477,N_2678,N_2761);
nor U3478 (N_3478,N_2273,N_2366);
nand U3479 (N_3479,N_2299,N_2744);
nor U3480 (N_3480,N_2451,N_2897);
or U3481 (N_3481,N_2509,N_2319);
and U3482 (N_3482,N_2875,N_2952);
xor U3483 (N_3483,N_2699,N_2302);
nor U3484 (N_3484,N_2856,N_2921);
nand U3485 (N_3485,N_2817,N_2576);
xnor U3486 (N_3486,N_2818,N_2278);
xnor U3487 (N_3487,N_2947,N_2292);
nor U3488 (N_3488,N_2620,N_2263);
nand U3489 (N_3489,N_2736,N_2621);
xnor U3490 (N_3490,N_2478,N_2560);
or U3491 (N_3491,N_2925,N_2902);
nand U3492 (N_3492,N_2942,N_2252);
and U3493 (N_3493,N_2905,N_2833);
nor U3494 (N_3494,N_2601,N_2693);
or U3495 (N_3495,N_2776,N_2855);
or U3496 (N_3496,N_2630,N_2494);
or U3497 (N_3497,N_2968,N_2619);
nor U3498 (N_3498,N_2860,N_2283);
nand U3499 (N_3499,N_2884,N_2407);
and U3500 (N_3500,N_2897,N_2691);
or U3501 (N_3501,N_2728,N_2814);
nor U3502 (N_3502,N_2394,N_2273);
nor U3503 (N_3503,N_2736,N_2507);
and U3504 (N_3504,N_2878,N_2604);
or U3505 (N_3505,N_2918,N_2473);
or U3506 (N_3506,N_2637,N_2818);
or U3507 (N_3507,N_2326,N_2828);
and U3508 (N_3508,N_2298,N_2485);
nor U3509 (N_3509,N_2534,N_2567);
nor U3510 (N_3510,N_2741,N_2251);
nor U3511 (N_3511,N_2503,N_2457);
xor U3512 (N_3512,N_2605,N_2467);
or U3513 (N_3513,N_2628,N_2774);
xor U3514 (N_3514,N_2374,N_2853);
nand U3515 (N_3515,N_2986,N_2484);
nand U3516 (N_3516,N_2861,N_2884);
nand U3517 (N_3517,N_2577,N_2950);
and U3518 (N_3518,N_2323,N_2862);
or U3519 (N_3519,N_2313,N_2676);
and U3520 (N_3520,N_2777,N_2873);
nand U3521 (N_3521,N_2278,N_2912);
nor U3522 (N_3522,N_2312,N_2855);
or U3523 (N_3523,N_2834,N_2525);
or U3524 (N_3524,N_2518,N_2259);
and U3525 (N_3525,N_2565,N_2495);
and U3526 (N_3526,N_2774,N_2885);
or U3527 (N_3527,N_2947,N_2414);
nand U3528 (N_3528,N_2657,N_2257);
and U3529 (N_3529,N_2699,N_2931);
or U3530 (N_3530,N_2366,N_2371);
xor U3531 (N_3531,N_2438,N_2305);
nand U3532 (N_3532,N_2252,N_2927);
xnor U3533 (N_3533,N_2564,N_2516);
nand U3534 (N_3534,N_2359,N_2573);
nor U3535 (N_3535,N_2656,N_2389);
and U3536 (N_3536,N_2906,N_2555);
or U3537 (N_3537,N_2932,N_2380);
or U3538 (N_3538,N_2364,N_2350);
or U3539 (N_3539,N_2464,N_2598);
and U3540 (N_3540,N_2440,N_2409);
nand U3541 (N_3541,N_2513,N_2816);
nand U3542 (N_3542,N_2841,N_2982);
and U3543 (N_3543,N_2512,N_2822);
and U3544 (N_3544,N_2559,N_2694);
nand U3545 (N_3545,N_2979,N_2313);
and U3546 (N_3546,N_2866,N_2875);
or U3547 (N_3547,N_2319,N_2745);
nand U3548 (N_3548,N_2281,N_2960);
nand U3549 (N_3549,N_2817,N_2396);
nor U3550 (N_3550,N_2869,N_2715);
or U3551 (N_3551,N_2534,N_2458);
xnor U3552 (N_3552,N_2340,N_2274);
nand U3553 (N_3553,N_2756,N_2815);
nor U3554 (N_3554,N_2428,N_2854);
nand U3555 (N_3555,N_2921,N_2438);
nor U3556 (N_3556,N_2946,N_2294);
nand U3557 (N_3557,N_2742,N_2779);
or U3558 (N_3558,N_2334,N_2525);
nor U3559 (N_3559,N_2529,N_2493);
and U3560 (N_3560,N_2661,N_2514);
nor U3561 (N_3561,N_2515,N_2615);
nor U3562 (N_3562,N_2927,N_2351);
or U3563 (N_3563,N_2649,N_2554);
nand U3564 (N_3564,N_2936,N_2365);
xor U3565 (N_3565,N_2736,N_2614);
and U3566 (N_3566,N_2925,N_2689);
nand U3567 (N_3567,N_2687,N_2617);
nor U3568 (N_3568,N_2379,N_2538);
nor U3569 (N_3569,N_2260,N_2341);
and U3570 (N_3570,N_2806,N_2708);
nor U3571 (N_3571,N_2528,N_2969);
nand U3572 (N_3572,N_2760,N_2858);
or U3573 (N_3573,N_2517,N_2552);
xnor U3574 (N_3574,N_2830,N_2374);
nand U3575 (N_3575,N_2711,N_2693);
or U3576 (N_3576,N_2267,N_2995);
nand U3577 (N_3577,N_2949,N_2530);
or U3578 (N_3578,N_2885,N_2959);
and U3579 (N_3579,N_2958,N_2536);
nand U3580 (N_3580,N_2959,N_2272);
nor U3581 (N_3581,N_2276,N_2560);
xor U3582 (N_3582,N_2589,N_2856);
nor U3583 (N_3583,N_2540,N_2992);
nor U3584 (N_3584,N_2738,N_2796);
xor U3585 (N_3585,N_2257,N_2577);
xnor U3586 (N_3586,N_2525,N_2740);
nand U3587 (N_3587,N_2328,N_2743);
nor U3588 (N_3588,N_2323,N_2671);
nand U3589 (N_3589,N_2530,N_2335);
or U3590 (N_3590,N_2820,N_2431);
xor U3591 (N_3591,N_2620,N_2285);
nand U3592 (N_3592,N_2504,N_2632);
nand U3593 (N_3593,N_2654,N_2413);
nand U3594 (N_3594,N_2284,N_2903);
nand U3595 (N_3595,N_2629,N_2904);
nor U3596 (N_3596,N_2542,N_2314);
and U3597 (N_3597,N_2643,N_2871);
and U3598 (N_3598,N_2317,N_2523);
xor U3599 (N_3599,N_2882,N_2551);
nor U3600 (N_3600,N_2779,N_2712);
and U3601 (N_3601,N_2903,N_2616);
or U3602 (N_3602,N_2640,N_2377);
nand U3603 (N_3603,N_2536,N_2382);
nor U3604 (N_3604,N_2414,N_2771);
nand U3605 (N_3605,N_2988,N_2652);
or U3606 (N_3606,N_2339,N_2708);
nand U3607 (N_3607,N_2839,N_2514);
nor U3608 (N_3608,N_2817,N_2914);
nor U3609 (N_3609,N_2271,N_2811);
and U3610 (N_3610,N_2384,N_2530);
nand U3611 (N_3611,N_2865,N_2654);
nor U3612 (N_3612,N_2675,N_2577);
nor U3613 (N_3613,N_2411,N_2672);
nand U3614 (N_3614,N_2766,N_2552);
nand U3615 (N_3615,N_2251,N_2840);
nand U3616 (N_3616,N_2302,N_2683);
or U3617 (N_3617,N_2552,N_2906);
and U3618 (N_3618,N_2912,N_2838);
and U3619 (N_3619,N_2884,N_2430);
and U3620 (N_3620,N_2437,N_2501);
or U3621 (N_3621,N_2401,N_2984);
or U3622 (N_3622,N_2971,N_2551);
nand U3623 (N_3623,N_2527,N_2514);
xor U3624 (N_3624,N_2824,N_2344);
nand U3625 (N_3625,N_2945,N_2449);
and U3626 (N_3626,N_2900,N_2460);
nor U3627 (N_3627,N_2866,N_2998);
xnor U3628 (N_3628,N_2352,N_2575);
xnor U3629 (N_3629,N_2634,N_2627);
nand U3630 (N_3630,N_2261,N_2822);
xnor U3631 (N_3631,N_2470,N_2388);
or U3632 (N_3632,N_2744,N_2457);
and U3633 (N_3633,N_2605,N_2313);
xor U3634 (N_3634,N_2865,N_2974);
and U3635 (N_3635,N_2280,N_2312);
nand U3636 (N_3636,N_2559,N_2444);
or U3637 (N_3637,N_2398,N_2790);
xnor U3638 (N_3638,N_2432,N_2786);
nor U3639 (N_3639,N_2532,N_2785);
nor U3640 (N_3640,N_2508,N_2875);
or U3641 (N_3641,N_2577,N_2714);
or U3642 (N_3642,N_2718,N_2904);
nand U3643 (N_3643,N_2763,N_2594);
xnor U3644 (N_3644,N_2636,N_2506);
nor U3645 (N_3645,N_2374,N_2468);
and U3646 (N_3646,N_2537,N_2852);
or U3647 (N_3647,N_2379,N_2254);
or U3648 (N_3648,N_2320,N_2842);
or U3649 (N_3649,N_2657,N_2987);
and U3650 (N_3650,N_2437,N_2780);
nor U3651 (N_3651,N_2251,N_2684);
or U3652 (N_3652,N_2916,N_2479);
and U3653 (N_3653,N_2952,N_2761);
or U3654 (N_3654,N_2468,N_2383);
nand U3655 (N_3655,N_2732,N_2976);
and U3656 (N_3656,N_2719,N_2850);
xnor U3657 (N_3657,N_2436,N_2933);
nand U3658 (N_3658,N_2561,N_2982);
and U3659 (N_3659,N_2705,N_2628);
or U3660 (N_3660,N_2587,N_2495);
nor U3661 (N_3661,N_2301,N_2550);
nor U3662 (N_3662,N_2915,N_2644);
nor U3663 (N_3663,N_2701,N_2258);
or U3664 (N_3664,N_2274,N_2412);
and U3665 (N_3665,N_2481,N_2819);
or U3666 (N_3666,N_2843,N_2365);
nor U3667 (N_3667,N_2656,N_2325);
nor U3668 (N_3668,N_2742,N_2692);
or U3669 (N_3669,N_2998,N_2715);
and U3670 (N_3670,N_2284,N_2509);
and U3671 (N_3671,N_2817,N_2466);
xor U3672 (N_3672,N_2507,N_2273);
and U3673 (N_3673,N_2666,N_2769);
nand U3674 (N_3674,N_2825,N_2437);
nand U3675 (N_3675,N_2777,N_2381);
nor U3676 (N_3676,N_2739,N_2816);
nor U3677 (N_3677,N_2281,N_2721);
or U3678 (N_3678,N_2918,N_2645);
and U3679 (N_3679,N_2921,N_2281);
nor U3680 (N_3680,N_2986,N_2994);
and U3681 (N_3681,N_2885,N_2479);
nor U3682 (N_3682,N_2795,N_2579);
nand U3683 (N_3683,N_2799,N_2566);
xnor U3684 (N_3684,N_2617,N_2341);
or U3685 (N_3685,N_2904,N_2889);
or U3686 (N_3686,N_2937,N_2518);
nand U3687 (N_3687,N_2980,N_2442);
nand U3688 (N_3688,N_2682,N_2588);
nor U3689 (N_3689,N_2714,N_2929);
nand U3690 (N_3690,N_2826,N_2465);
nor U3691 (N_3691,N_2933,N_2448);
nand U3692 (N_3692,N_2994,N_2677);
or U3693 (N_3693,N_2908,N_2808);
or U3694 (N_3694,N_2705,N_2252);
nand U3695 (N_3695,N_2438,N_2288);
xnor U3696 (N_3696,N_2724,N_2397);
and U3697 (N_3697,N_2363,N_2957);
nor U3698 (N_3698,N_2834,N_2818);
nor U3699 (N_3699,N_2899,N_2278);
nor U3700 (N_3700,N_2460,N_2735);
and U3701 (N_3701,N_2335,N_2710);
nand U3702 (N_3702,N_2391,N_2967);
nand U3703 (N_3703,N_2262,N_2605);
nand U3704 (N_3704,N_2696,N_2272);
or U3705 (N_3705,N_2792,N_2728);
nand U3706 (N_3706,N_2597,N_2787);
nand U3707 (N_3707,N_2478,N_2411);
or U3708 (N_3708,N_2352,N_2942);
and U3709 (N_3709,N_2824,N_2260);
nor U3710 (N_3710,N_2891,N_2268);
or U3711 (N_3711,N_2438,N_2977);
nand U3712 (N_3712,N_2646,N_2591);
nand U3713 (N_3713,N_2547,N_2852);
and U3714 (N_3714,N_2461,N_2998);
nand U3715 (N_3715,N_2503,N_2719);
nor U3716 (N_3716,N_2875,N_2744);
or U3717 (N_3717,N_2980,N_2477);
nand U3718 (N_3718,N_2337,N_2474);
or U3719 (N_3719,N_2297,N_2646);
nor U3720 (N_3720,N_2920,N_2904);
xnor U3721 (N_3721,N_2978,N_2992);
and U3722 (N_3722,N_2833,N_2757);
nor U3723 (N_3723,N_2792,N_2503);
nor U3724 (N_3724,N_2912,N_2546);
nand U3725 (N_3725,N_2762,N_2958);
and U3726 (N_3726,N_2302,N_2448);
or U3727 (N_3727,N_2822,N_2418);
nor U3728 (N_3728,N_2313,N_2777);
nand U3729 (N_3729,N_2765,N_2637);
or U3730 (N_3730,N_2809,N_2461);
or U3731 (N_3731,N_2831,N_2648);
and U3732 (N_3732,N_2697,N_2887);
and U3733 (N_3733,N_2450,N_2388);
and U3734 (N_3734,N_2857,N_2597);
or U3735 (N_3735,N_2256,N_2527);
nand U3736 (N_3736,N_2384,N_2822);
nand U3737 (N_3737,N_2678,N_2579);
nand U3738 (N_3738,N_2797,N_2724);
nand U3739 (N_3739,N_2601,N_2362);
and U3740 (N_3740,N_2973,N_2961);
nor U3741 (N_3741,N_2633,N_2913);
and U3742 (N_3742,N_2572,N_2371);
nor U3743 (N_3743,N_2996,N_2553);
nand U3744 (N_3744,N_2334,N_2930);
nor U3745 (N_3745,N_2531,N_2448);
xor U3746 (N_3746,N_2485,N_2316);
and U3747 (N_3747,N_2436,N_2804);
nor U3748 (N_3748,N_2910,N_2786);
nand U3749 (N_3749,N_2328,N_2993);
and U3750 (N_3750,N_3741,N_3330);
nand U3751 (N_3751,N_3390,N_3018);
and U3752 (N_3752,N_3538,N_3347);
or U3753 (N_3753,N_3176,N_3544);
and U3754 (N_3754,N_3582,N_3216);
or U3755 (N_3755,N_3065,N_3572);
and U3756 (N_3756,N_3139,N_3644);
nand U3757 (N_3757,N_3120,N_3668);
and U3758 (N_3758,N_3612,N_3170);
or U3759 (N_3759,N_3740,N_3081);
nor U3760 (N_3760,N_3445,N_3415);
nor U3761 (N_3761,N_3541,N_3332);
xnor U3762 (N_3762,N_3031,N_3632);
and U3763 (N_3763,N_3517,N_3697);
nor U3764 (N_3764,N_3063,N_3472);
and U3765 (N_3765,N_3079,N_3102);
and U3766 (N_3766,N_3097,N_3345);
or U3767 (N_3767,N_3026,N_3490);
nand U3768 (N_3768,N_3615,N_3092);
and U3769 (N_3769,N_3314,N_3640);
and U3770 (N_3770,N_3308,N_3211);
xnor U3771 (N_3771,N_3661,N_3462);
and U3772 (N_3772,N_3013,N_3224);
and U3773 (N_3773,N_3007,N_3525);
nor U3774 (N_3774,N_3496,N_3564);
or U3775 (N_3775,N_3125,N_3484);
xor U3776 (N_3776,N_3208,N_3118);
nor U3777 (N_3777,N_3707,N_3112);
xnor U3778 (N_3778,N_3491,N_3685);
nor U3779 (N_3779,N_3128,N_3482);
or U3780 (N_3780,N_3457,N_3570);
nand U3781 (N_3781,N_3610,N_3519);
or U3782 (N_3782,N_3161,N_3248);
and U3783 (N_3783,N_3639,N_3736);
and U3784 (N_3784,N_3521,N_3718);
or U3785 (N_3785,N_3704,N_3160);
and U3786 (N_3786,N_3368,N_3370);
and U3787 (N_3787,N_3188,N_3237);
or U3788 (N_3788,N_3398,N_3158);
xor U3789 (N_3789,N_3738,N_3713);
nor U3790 (N_3790,N_3503,N_3015);
nor U3791 (N_3791,N_3405,N_3372);
or U3792 (N_3792,N_3399,N_3413);
nand U3793 (N_3793,N_3074,N_3645);
nand U3794 (N_3794,N_3705,N_3284);
or U3795 (N_3795,N_3289,N_3614);
nand U3796 (N_3796,N_3137,N_3367);
or U3797 (N_3797,N_3229,N_3191);
and U3798 (N_3798,N_3606,N_3146);
nor U3799 (N_3799,N_3657,N_3017);
xor U3800 (N_3800,N_3028,N_3362);
or U3801 (N_3801,N_3667,N_3194);
or U3802 (N_3802,N_3396,N_3428);
nor U3803 (N_3803,N_3662,N_3327);
nor U3804 (N_3804,N_3649,N_3604);
nor U3805 (N_3805,N_3300,N_3673);
nand U3806 (N_3806,N_3566,N_3551);
or U3807 (N_3807,N_3175,N_3545);
nand U3808 (N_3808,N_3556,N_3285);
nand U3809 (N_3809,N_3524,N_3595);
or U3810 (N_3810,N_3051,N_3322);
nor U3811 (N_3811,N_3058,N_3231);
nor U3812 (N_3812,N_3302,N_3268);
or U3813 (N_3813,N_3388,N_3217);
and U3814 (N_3814,N_3167,N_3195);
or U3815 (N_3815,N_3077,N_3351);
or U3816 (N_3816,N_3111,N_3493);
nand U3817 (N_3817,N_3041,N_3312);
or U3818 (N_3818,N_3497,N_3076);
and U3819 (N_3819,N_3676,N_3392);
and U3820 (N_3820,N_3528,N_3295);
nand U3821 (N_3821,N_3546,N_3559);
xor U3822 (N_3822,N_3173,N_3215);
nand U3823 (N_3823,N_3671,N_3547);
xor U3824 (N_3824,N_3591,N_3131);
nor U3825 (N_3825,N_3720,N_3068);
and U3826 (N_3826,N_3476,N_3350);
or U3827 (N_3827,N_3316,N_3333);
nor U3828 (N_3828,N_3230,N_3091);
nor U3829 (N_3829,N_3393,N_3653);
and U3830 (N_3830,N_3261,N_3425);
and U3831 (N_3831,N_3729,N_3067);
nand U3832 (N_3832,N_3672,N_3204);
nand U3833 (N_3833,N_3679,N_3107);
nor U3834 (N_3834,N_3200,N_3179);
nand U3835 (N_3835,N_3353,N_3470);
nand U3836 (N_3836,N_3123,N_3394);
or U3837 (N_3837,N_3724,N_3071);
or U3838 (N_3838,N_3127,N_3562);
and U3839 (N_3839,N_3287,N_3294);
and U3840 (N_3840,N_3417,N_3296);
or U3841 (N_3841,N_3335,N_3590);
or U3842 (N_3842,N_3611,N_3251);
or U3843 (N_3843,N_3600,N_3499);
or U3844 (N_3844,N_3433,N_3070);
and U3845 (N_3845,N_3605,N_3737);
or U3846 (N_3846,N_3592,N_3563);
or U3847 (N_3847,N_3078,N_3492);
nand U3848 (N_3848,N_3168,N_3747);
and U3849 (N_3849,N_3714,N_3011);
nor U3850 (N_3850,N_3607,N_3648);
or U3851 (N_3851,N_3010,N_3549);
nor U3852 (N_3852,N_3043,N_3723);
nand U3853 (N_3853,N_3133,N_3603);
nor U3854 (N_3854,N_3371,N_3523);
nor U3855 (N_3855,N_3317,N_3171);
nor U3856 (N_3856,N_3505,N_3203);
or U3857 (N_3857,N_3637,N_3522);
nor U3858 (N_3858,N_3042,N_3656);
and U3859 (N_3859,N_3197,N_3337);
and U3860 (N_3860,N_3264,N_3084);
and U3861 (N_3861,N_3000,N_3543);
nand U3862 (N_3862,N_3282,N_3647);
nor U3863 (N_3863,N_3708,N_3373);
or U3864 (N_3864,N_3022,N_3374);
nand U3865 (N_3865,N_3029,N_3530);
nor U3866 (N_3866,N_3735,N_3004);
nor U3867 (N_3867,N_3354,N_3400);
nand U3868 (N_3868,N_3222,N_3002);
and U3869 (N_3869,N_3620,N_3432);
and U3870 (N_3870,N_3115,N_3085);
and U3871 (N_3871,N_3186,N_3542);
and U3872 (N_3872,N_3514,N_3508);
nor U3873 (N_3873,N_3243,N_3658);
and U3874 (N_3874,N_3536,N_3193);
or U3875 (N_3875,N_3693,N_3087);
nand U3876 (N_3876,N_3655,N_3181);
nor U3877 (N_3877,N_3323,N_3096);
and U3878 (N_3878,N_3262,N_3424);
or U3879 (N_3879,N_3165,N_3512);
and U3880 (N_3880,N_3421,N_3006);
and U3881 (N_3881,N_3040,N_3739);
or U3882 (N_3882,N_3478,N_3275);
and U3883 (N_3883,N_3280,N_3108);
nand U3884 (N_3884,N_3721,N_3369);
nand U3885 (N_3885,N_3257,N_3054);
nand U3886 (N_3886,N_3122,N_3250);
nand U3887 (N_3887,N_3613,N_3162);
nand U3888 (N_3888,N_3682,N_3587);
nand U3889 (N_3889,N_3474,N_3397);
and U3890 (N_3890,N_3520,N_3526);
xor U3891 (N_3891,N_3716,N_3357);
nor U3892 (N_3892,N_3409,N_3539);
nand U3893 (N_3893,N_3691,N_3252);
nor U3894 (N_3894,N_3325,N_3489);
and U3895 (N_3895,N_3745,N_3192);
or U3896 (N_3896,N_3279,N_3410);
nand U3897 (N_3897,N_3164,N_3328);
xnor U3898 (N_3898,N_3598,N_3038);
or U3899 (N_3899,N_3638,N_3073);
nor U3900 (N_3900,N_3385,N_3451);
xnor U3901 (N_3901,N_3419,N_3273);
and U3902 (N_3902,N_3646,N_3660);
and U3903 (N_3903,N_3293,N_3298);
nand U3904 (N_3904,N_3456,N_3113);
and U3905 (N_3905,N_3339,N_3225);
nand U3906 (N_3906,N_3575,N_3185);
or U3907 (N_3907,N_3506,N_3448);
xnor U3908 (N_3908,N_3555,N_3731);
and U3909 (N_3909,N_3310,N_3386);
nand U3910 (N_3910,N_3001,N_3453);
nand U3911 (N_3911,N_3288,N_3364);
nand U3912 (N_3912,N_3597,N_3098);
or U3913 (N_3913,N_3036,N_3683);
nor U3914 (N_3914,N_3182,N_3481);
and U3915 (N_3915,N_3654,N_3381);
and U3916 (N_3916,N_3291,N_3553);
nand U3917 (N_3917,N_3046,N_3232);
and U3918 (N_3918,N_3458,N_3035);
or U3919 (N_3919,N_3151,N_3062);
or U3920 (N_3920,N_3408,N_3548);
xor U3921 (N_3921,N_3636,N_3343);
xnor U3922 (N_3922,N_3272,N_3190);
xnor U3923 (N_3923,N_3064,N_3665);
and U3924 (N_3924,N_3114,N_3037);
or U3925 (N_3925,N_3246,N_3675);
nor U3926 (N_3926,N_3473,N_3196);
or U3927 (N_3927,N_3532,N_3550);
or U3928 (N_3928,N_3075,N_3053);
nor U3929 (N_3929,N_3320,N_3044);
nor U3930 (N_3930,N_3465,N_3341);
nor U3931 (N_3931,N_3579,N_3034);
nor U3932 (N_3932,N_3699,N_3309);
nor U3933 (N_3933,N_3283,N_3609);
or U3934 (N_3934,N_3659,N_3663);
and U3935 (N_3935,N_3256,N_3177);
nor U3936 (N_3936,N_3263,N_3677);
and U3937 (N_3937,N_3460,N_3634);
nand U3938 (N_3938,N_3558,N_3576);
or U3939 (N_3939,N_3578,N_3728);
and U3940 (N_3940,N_3537,N_3265);
nor U3941 (N_3941,N_3121,N_3702);
and U3942 (N_3942,N_3441,N_3206);
nor U3943 (N_3943,N_3395,N_3163);
nor U3944 (N_3944,N_3223,N_3346);
and U3945 (N_3945,N_3239,N_3515);
nand U3946 (N_3946,N_3746,N_3055);
nor U3947 (N_3947,N_3141,N_3418);
and U3948 (N_3948,N_3082,N_3266);
and U3949 (N_3949,N_3694,N_3535);
nand U3950 (N_3950,N_3406,N_3743);
or U3951 (N_3951,N_3387,N_3726);
nor U3952 (N_3952,N_3153,N_3389);
nor U3953 (N_3953,N_3749,N_3129);
nor U3954 (N_3954,N_3226,N_3375);
and U3955 (N_3955,N_3502,N_3414);
or U3956 (N_3956,N_3500,N_3089);
nand U3957 (N_3957,N_3241,N_3233);
or U3958 (N_3958,N_3618,N_3733);
and U3959 (N_3959,N_3305,N_3198);
and U3960 (N_3960,N_3379,N_3099);
and U3961 (N_3961,N_3722,N_3643);
and U3962 (N_3962,N_3416,N_3292);
nand U3963 (N_3963,N_3688,N_3003);
or U3964 (N_3964,N_3147,N_3355);
or U3965 (N_3965,N_3422,N_3495);
or U3966 (N_3966,N_3411,N_3577);
nor U3967 (N_3967,N_3259,N_3510);
or U3968 (N_3968,N_3629,N_3331);
nor U3969 (N_3969,N_3380,N_3623);
nand U3970 (N_3970,N_3471,N_3023);
or U3971 (N_3971,N_3130,N_3650);
or U3972 (N_3972,N_3719,N_3156);
xor U3973 (N_3973,N_3104,N_3533);
and U3974 (N_3974,N_3069,N_3219);
or U3975 (N_3975,N_3365,N_3338);
nand U3976 (N_3976,N_3318,N_3468);
and U3977 (N_3977,N_3218,N_3686);
and U3978 (N_3978,N_3106,N_3446);
or U3979 (N_3979,N_3254,N_3593);
and U3980 (N_3980,N_3205,N_3270);
nand U3981 (N_3981,N_3617,N_3286);
nand U3982 (N_3982,N_3336,N_3701);
nand U3983 (N_3983,N_3080,N_3485);
nand U3984 (N_3984,N_3596,N_3630);
and U3985 (N_3985,N_3150,N_3455);
nand U3986 (N_3986,N_3260,N_3119);
nand U3987 (N_3987,N_3569,N_3678);
nand U3988 (N_3988,N_3621,N_3066);
and U3989 (N_3989,N_3083,N_3124);
and U3990 (N_3990,N_3625,N_3635);
or U3991 (N_3991,N_3689,N_3202);
nand U3992 (N_3992,N_3450,N_3420);
nor U3993 (N_3993,N_3507,N_3384);
or U3994 (N_3994,N_3172,N_3238);
xnor U3995 (N_3995,N_3602,N_3475);
or U3996 (N_3996,N_3437,N_3401);
or U3997 (N_3997,N_3024,N_3624);
and U3998 (N_3998,N_3047,N_3435);
xor U3999 (N_3999,N_3383,N_3090);
or U4000 (N_4000,N_3692,N_3711);
nand U4001 (N_4001,N_3477,N_3324);
nand U4002 (N_4002,N_3152,N_3690);
and U4003 (N_4003,N_3531,N_3267);
nor U4004 (N_4004,N_3178,N_3014);
and U4005 (N_4005,N_3454,N_3511);
nor U4006 (N_4006,N_3431,N_3277);
or U4007 (N_4007,N_3027,N_3715);
nor U4008 (N_4008,N_3377,N_3666);
and U4009 (N_4009,N_3391,N_3641);
nor U4010 (N_4010,N_3366,N_3321);
and U4011 (N_4011,N_3571,N_3594);
nor U4012 (N_4012,N_3568,N_3005);
xnor U4013 (N_4013,N_3479,N_3221);
nor U4014 (N_4014,N_3050,N_3360);
nand U4015 (N_4015,N_3340,N_3651);
or U4016 (N_4016,N_3378,N_3466);
nor U4017 (N_4017,N_3313,N_3142);
nor U4018 (N_4018,N_3138,N_3616);
or U4019 (N_4019,N_3297,N_3169);
or U4020 (N_4020,N_3467,N_3463);
or U4021 (N_4021,N_3363,N_3274);
and U4022 (N_4022,N_3627,N_3599);
nor U4023 (N_4023,N_3601,N_3326);
and U4024 (N_4024,N_3464,N_3235);
nor U4025 (N_4025,N_3744,N_3516);
xnor U4026 (N_4026,N_3444,N_3086);
or U4027 (N_4027,N_3669,N_3376);
or U4028 (N_4028,N_3244,N_3201);
nand U4029 (N_4029,N_3404,N_3228);
nor U4030 (N_4030,N_3032,N_3271);
nor U4031 (N_4031,N_3427,N_3342);
nand U4032 (N_4032,N_3144,N_3717);
nor U4033 (N_4033,N_3154,N_3057);
and U4034 (N_4034,N_3469,N_3429);
or U4035 (N_4035,N_3748,N_3586);
and U4036 (N_4036,N_3356,N_3025);
and U4037 (N_4037,N_3434,N_3242);
and U4038 (N_4038,N_3443,N_3573);
and U4039 (N_4039,N_3407,N_3487);
nor U4040 (N_4040,N_3220,N_3207);
xor U4041 (N_4041,N_3132,N_3301);
or U4042 (N_4042,N_3608,N_3253);
or U4043 (N_4043,N_3180,N_3136);
nor U4044 (N_4044,N_3019,N_3430);
nor U4045 (N_4045,N_3276,N_3258);
nand U4046 (N_4046,N_3134,N_3567);
or U4047 (N_4047,N_3020,N_3712);
or U4048 (N_4048,N_3101,N_3403);
nand U4049 (N_4049,N_3311,N_3299);
and U4050 (N_4050,N_3212,N_3008);
xor U4051 (N_4051,N_3695,N_3583);
or U4052 (N_4052,N_3382,N_3059);
and U4053 (N_4053,N_3199,N_3249);
nor U4054 (N_4054,N_3157,N_3358);
nand U4055 (N_4055,N_3359,N_3245);
xnor U4056 (N_4056,N_3110,N_3278);
and U4057 (N_4057,N_3227,N_3652);
nor U4058 (N_4058,N_3440,N_3329);
nor U4059 (N_4059,N_3449,N_3045);
nor U4060 (N_4060,N_3269,N_3725);
xor U4061 (N_4061,N_3094,N_3426);
and U4062 (N_4062,N_3145,N_3633);
nor U4063 (N_4063,N_3631,N_3174);
nor U4064 (N_4064,N_3060,N_3439);
or U4065 (N_4065,N_3509,N_3436);
and U4066 (N_4066,N_3412,N_3109);
and U4067 (N_4067,N_3732,N_3304);
and U4068 (N_4068,N_3438,N_3095);
or U4069 (N_4069,N_3684,N_3159);
and U4070 (N_4070,N_3518,N_3494);
nand U4071 (N_4071,N_3213,N_3642);
and U4072 (N_4072,N_3072,N_3116);
or U4073 (N_4073,N_3210,N_3483);
nand U4074 (N_4074,N_3187,N_3140);
and U4075 (N_4075,N_3247,N_3710);
nor U4076 (N_4076,N_3189,N_3009);
nand U4077 (N_4077,N_3021,N_3349);
and U4078 (N_4078,N_3135,N_3700);
nand U4079 (N_4079,N_3670,N_3461);
and U4080 (N_4080,N_3016,N_3459);
nor U4081 (N_4081,N_3480,N_3565);
nand U4082 (N_4082,N_3117,N_3734);
nor U4083 (N_4083,N_3581,N_3100);
nand U4084 (N_4084,N_3049,N_3255);
nor U4085 (N_4085,N_3727,N_3103);
nand U4086 (N_4086,N_3214,N_3184);
and U4087 (N_4087,N_3504,N_3628);
or U4088 (N_4088,N_3498,N_3557);
nor U4089 (N_4089,N_3166,N_3088);
and U4090 (N_4090,N_3240,N_3149);
nor U4091 (N_4091,N_3030,N_3501);
or U4092 (N_4092,N_3709,N_3307);
and U4093 (N_4093,N_3447,N_3742);
nand U4094 (N_4094,N_3698,N_3352);
nand U4095 (N_4095,N_3319,N_3209);
or U4096 (N_4096,N_3585,N_3552);
nor U4097 (N_4097,N_3361,N_3488);
nor U4098 (N_4098,N_3234,N_3703);
nand U4099 (N_4099,N_3143,N_3561);
nand U4100 (N_4100,N_3056,N_3344);
or U4101 (N_4101,N_3486,N_3534);
nor U4102 (N_4102,N_3674,N_3281);
and U4103 (N_4103,N_3061,N_3334);
or U4104 (N_4104,N_3527,N_3033);
nand U4105 (N_4105,N_3589,N_3315);
nand U4106 (N_4106,N_3588,N_3580);
and U4107 (N_4107,N_3554,N_3513);
nand U4108 (N_4108,N_3680,N_3687);
or U4109 (N_4109,N_3093,N_3348);
xor U4110 (N_4110,N_3290,N_3155);
nand U4111 (N_4111,N_3540,N_3529);
nor U4112 (N_4112,N_3664,N_3048);
nand U4113 (N_4113,N_3584,N_3730);
nor U4114 (N_4114,N_3126,N_3626);
nand U4115 (N_4115,N_3619,N_3452);
nand U4116 (N_4116,N_3622,N_3402);
and U4117 (N_4117,N_3560,N_3052);
or U4118 (N_4118,N_3574,N_3442);
nor U4119 (N_4119,N_3183,N_3236);
or U4120 (N_4120,N_3696,N_3105);
nand U4121 (N_4121,N_3681,N_3039);
nand U4122 (N_4122,N_3148,N_3012);
nand U4123 (N_4123,N_3306,N_3423);
or U4124 (N_4124,N_3706,N_3303);
and U4125 (N_4125,N_3318,N_3562);
nor U4126 (N_4126,N_3510,N_3500);
nand U4127 (N_4127,N_3711,N_3501);
and U4128 (N_4128,N_3595,N_3180);
or U4129 (N_4129,N_3488,N_3226);
and U4130 (N_4130,N_3145,N_3339);
nand U4131 (N_4131,N_3014,N_3540);
xor U4132 (N_4132,N_3123,N_3389);
and U4133 (N_4133,N_3714,N_3122);
xor U4134 (N_4134,N_3155,N_3440);
and U4135 (N_4135,N_3417,N_3528);
nand U4136 (N_4136,N_3740,N_3039);
nor U4137 (N_4137,N_3653,N_3741);
nor U4138 (N_4138,N_3642,N_3550);
nand U4139 (N_4139,N_3054,N_3269);
nor U4140 (N_4140,N_3732,N_3172);
nand U4141 (N_4141,N_3478,N_3238);
nand U4142 (N_4142,N_3093,N_3027);
or U4143 (N_4143,N_3029,N_3464);
and U4144 (N_4144,N_3339,N_3298);
or U4145 (N_4145,N_3527,N_3632);
nand U4146 (N_4146,N_3460,N_3443);
or U4147 (N_4147,N_3293,N_3663);
nor U4148 (N_4148,N_3719,N_3575);
and U4149 (N_4149,N_3000,N_3732);
and U4150 (N_4150,N_3450,N_3593);
nand U4151 (N_4151,N_3493,N_3339);
and U4152 (N_4152,N_3251,N_3617);
and U4153 (N_4153,N_3249,N_3715);
nor U4154 (N_4154,N_3107,N_3351);
or U4155 (N_4155,N_3272,N_3281);
and U4156 (N_4156,N_3314,N_3678);
and U4157 (N_4157,N_3272,N_3624);
nand U4158 (N_4158,N_3441,N_3503);
nor U4159 (N_4159,N_3103,N_3194);
nor U4160 (N_4160,N_3126,N_3549);
and U4161 (N_4161,N_3465,N_3620);
and U4162 (N_4162,N_3135,N_3573);
or U4163 (N_4163,N_3695,N_3585);
nor U4164 (N_4164,N_3231,N_3198);
nand U4165 (N_4165,N_3598,N_3629);
nor U4166 (N_4166,N_3285,N_3519);
nor U4167 (N_4167,N_3315,N_3149);
nor U4168 (N_4168,N_3045,N_3402);
and U4169 (N_4169,N_3073,N_3331);
or U4170 (N_4170,N_3209,N_3089);
nor U4171 (N_4171,N_3241,N_3338);
and U4172 (N_4172,N_3735,N_3388);
or U4173 (N_4173,N_3070,N_3570);
nand U4174 (N_4174,N_3216,N_3436);
nor U4175 (N_4175,N_3333,N_3172);
nor U4176 (N_4176,N_3534,N_3399);
nand U4177 (N_4177,N_3586,N_3738);
nand U4178 (N_4178,N_3250,N_3654);
nor U4179 (N_4179,N_3738,N_3099);
nor U4180 (N_4180,N_3242,N_3605);
and U4181 (N_4181,N_3182,N_3672);
nor U4182 (N_4182,N_3092,N_3635);
nor U4183 (N_4183,N_3434,N_3239);
and U4184 (N_4184,N_3557,N_3251);
or U4185 (N_4185,N_3346,N_3565);
or U4186 (N_4186,N_3355,N_3069);
nor U4187 (N_4187,N_3268,N_3355);
nand U4188 (N_4188,N_3165,N_3288);
and U4189 (N_4189,N_3390,N_3036);
or U4190 (N_4190,N_3128,N_3749);
and U4191 (N_4191,N_3530,N_3116);
nor U4192 (N_4192,N_3238,N_3184);
xnor U4193 (N_4193,N_3105,N_3398);
nor U4194 (N_4194,N_3208,N_3406);
nor U4195 (N_4195,N_3267,N_3366);
nand U4196 (N_4196,N_3604,N_3680);
nand U4197 (N_4197,N_3049,N_3729);
nor U4198 (N_4198,N_3241,N_3317);
nand U4199 (N_4199,N_3281,N_3172);
nor U4200 (N_4200,N_3312,N_3492);
xnor U4201 (N_4201,N_3354,N_3408);
nor U4202 (N_4202,N_3274,N_3538);
and U4203 (N_4203,N_3526,N_3651);
xnor U4204 (N_4204,N_3687,N_3547);
nor U4205 (N_4205,N_3406,N_3011);
xnor U4206 (N_4206,N_3335,N_3595);
nand U4207 (N_4207,N_3460,N_3398);
nor U4208 (N_4208,N_3256,N_3636);
nor U4209 (N_4209,N_3476,N_3196);
and U4210 (N_4210,N_3293,N_3370);
and U4211 (N_4211,N_3504,N_3734);
nand U4212 (N_4212,N_3357,N_3453);
and U4213 (N_4213,N_3603,N_3260);
nor U4214 (N_4214,N_3599,N_3325);
and U4215 (N_4215,N_3691,N_3528);
or U4216 (N_4216,N_3264,N_3291);
or U4217 (N_4217,N_3687,N_3302);
or U4218 (N_4218,N_3087,N_3128);
nand U4219 (N_4219,N_3017,N_3555);
and U4220 (N_4220,N_3742,N_3137);
nor U4221 (N_4221,N_3091,N_3636);
or U4222 (N_4222,N_3030,N_3198);
or U4223 (N_4223,N_3692,N_3319);
nand U4224 (N_4224,N_3249,N_3649);
nand U4225 (N_4225,N_3126,N_3147);
or U4226 (N_4226,N_3104,N_3474);
nor U4227 (N_4227,N_3429,N_3706);
nand U4228 (N_4228,N_3266,N_3148);
or U4229 (N_4229,N_3247,N_3168);
or U4230 (N_4230,N_3387,N_3588);
nand U4231 (N_4231,N_3435,N_3457);
and U4232 (N_4232,N_3435,N_3188);
or U4233 (N_4233,N_3017,N_3550);
xor U4234 (N_4234,N_3277,N_3464);
nor U4235 (N_4235,N_3180,N_3485);
or U4236 (N_4236,N_3648,N_3135);
nor U4237 (N_4237,N_3360,N_3249);
or U4238 (N_4238,N_3065,N_3599);
nand U4239 (N_4239,N_3537,N_3309);
xnor U4240 (N_4240,N_3114,N_3344);
and U4241 (N_4241,N_3218,N_3557);
nor U4242 (N_4242,N_3304,N_3744);
nand U4243 (N_4243,N_3304,N_3469);
and U4244 (N_4244,N_3714,N_3087);
or U4245 (N_4245,N_3357,N_3719);
and U4246 (N_4246,N_3072,N_3133);
xnor U4247 (N_4247,N_3655,N_3275);
and U4248 (N_4248,N_3562,N_3057);
or U4249 (N_4249,N_3676,N_3430);
nor U4250 (N_4250,N_3289,N_3661);
or U4251 (N_4251,N_3146,N_3142);
xor U4252 (N_4252,N_3512,N_3424);
xnor U4253 (N_4253,N_3695,N_3388);
and U4254 (N_4254,N_3326,N_3529);
nand U4255 (N_4255,N_3499,N_3642);
and U4256 (N_4256,N_3460,N_3339);
and U4257 (N_4257,N_3668,N_3497);
and U4258 (N_4258,N_3673,N_3497);
or U4259 (N_4259,N_3530,N_3052);
or U4260 (N_4260,N_3237,N_3455);
nand U4261 (N_4261,N_3216,N_3079);
nand U4262 (N_4262,N_3734,N_3207);
xnor U4263 (N_4263,N_3255,N_3104);
and U4264 (N_4264,N_3477,N_3734);
xor U4265 (N_4265,N_3335,N_3462);
nand U4266 (N_4266,N_3375,N_3457);
and U4267 (N_4267,N_3478,N_3225);
and U4268 (N_4268,N_3502,N_3591);
and U4269 (N_4269,N_3518,N_3619);
and U4270 (N_4270,N_3049,N_3327);
nand U4271 (N_4271,N_3511,N_3435);
nand U4272 (N_4272,N_3413,N_3233);
nor U4273 (N_4273,N_3354,N_3675);
nand U4274 (N_4274,N_3167,N_3350);
and U4275 (N_4275,N_3255,N_3389);
nand U4276 (N_4276,N_3472,N_3362);
xnor U4277 (N_4277,N_3732,N_3309);
or U4278 (N_4278,N_3322,N_3163);
or U4279 (N_4279,N_3627,N_3444);
and U4280 (N_4280,N_3570,N_3057);
nor U4281 (N_4281,N_3241,N_3605);
and U4282 (N_4282,N_3021,N_3118);
or U4283 (N_4283,N_3366,N_3059);
and U4284 (N_4284,N_3487,N_3747);
or U4285 (N_4285,N_3200,N_3558);
nand U4286 (N_4286,N_3434,N_3367);
nor U4287 (N_4287,N_3733,N_3028);
or U4288 (N_4288,N_3036,N_3141);
or U4289 (N_4289,N_3374,N_3169);
or U4290 (N_4290,N_3440,N_3107);
or U4291 (N_4291,N_3451,N_3398);
xnor U4292 (N_4292,N_3172,N_3606);
nand U4293 (N_4293,N_3108,N_3355);
nor U4294 (N_4294,N_3217,N_3285);
nand U4295 (N_4295,N_3396,N_3643);
nand U4296 (N_4296,N_3391,N_3215);
xnor U4297 (N_4297,N_3230,N_3159);
and U4298 (N_4298,N_3316,N_3427);
or U4299 (N_4299,N_3740,N_3361);
nand U4300 (N_4300,N_3615,N_3478);
nor U4301 (N_4301,N_3399,N_3663);
nor U4302 (N_4302,N_3522,N_3135);
nor U4303 (N_4303,N_3081,N_3730);
nand U4304 (N_4304,N_3461,N_3359);
or U4305 (N_4305,N_3711,N_3262);
and U4306 (N_4306,N_3409,N_3498);
and U4307 (N_4307,N_3304,N_3146);
xnor U4308 (N_4308,N_3389,N_3240);
or U4309 (N_4309,N_3494,N_3297);
nor U4310 (N_4310,N_3315,N_3200);
nand U4311 (N_4311,N_3531,N_3358);
nand U4312 (N_4312,N_3730,N_3066);
xnor U4313 (N_4313,N_3282,N_3028);
and U4314 (N_4314,N_3579,N_3654);
or U4315 (N_4315,N_3040,N_3076);
and U4316 (N_4316,N_3715,N_3257);
and U4317 (N_4317,N_3215,N_3259);
nor U4318 (N_4318,N_3194,N_3137);
nand U4319 (N_4319,N_3320,N_3000);
or U4320 (N_4320,N_3114,N_3688);
xnor U4321 (N_4321,N_3356,N_3194);
nand U4322 (N_4322,N_3603,N_3612);
nor U4323 (N_4323,N_3294,N_3167);
and U4324 (N_4324,N_3075,N_3538);
and U4325 (N_4325,N_3592,N_3743);
nand U4326 (N_4326,N_3077,N_3507);
nor U4327 (N_4327,N_3351,N_3304);
nand U4328 (N_4328,N_3172,N_3650);
or U4329 (N_4329,N_3563,N_3180);
nor U4330 (N_4330,N_3092,N_3159);
nor U4331 (N_4331,N_3332,N_3665);
and U4332 (N_4332,N_3225,N_3524);
nand U4333 (N_4333,N_3535,N_3446);
nand U4334 (N_4334,N_3270,N_3603);
or U4335 (N_4335,N_3461,N_3041);
nand U4336 (N_4336,N_3289,N_3456);
and U4337 (N_4337,N_3028,N_3216);
nor U4338 (N_4338,N_3244,N_3507);
or U4339 (N_4339,N_3443,N_3361);
nor U4340 (N_4340,N_3183,N_3006);
or U4341 (N_4341,N_3405,N_3225);
nor U4342 (N_4342,N_3456,N_3155);
and U4343 (N_4343,N_3104,N_3114);
and U4344 (N_4344,N_3051,N_3499);
or U4345 (N_4345,N_3305,N_3370);
nand U4346 (N_4346,N_3113,N_3603);
nor U4347 (N_4347,N_3067,N_3526);
or U4348 (N_4348,N_3279,N_3234);
xor U4349 (N_4349,N_3014,N_3270);
nand U4350 (N_4350,N_3125,N_3450);
and U4351 (N_4351,N_3220,N_3510);
and U4352 (N_4352,N_3660,N_3667);
nand U4353 (N_4353,N_3480,N_3648);
or U4354 (N_4354,N_3494,N_3270);
and U4355 (N_4355,N_3211,N_3416);
and U4356 (N_4356,N_3438,N_3319);
nand U4357 (N_4357,N_3261,N_3015);
and U4358 (N_4358,N_3610,N_3230);
xor U4359 (N_4359,N_3678,N_3589);
nand U4360 (N_4360,N_3596,N_3464);
nand U4361 (N_4361,N_3582,N_3128);
and U4362 (N_4362,N_3146,N_3712);
nand U4363 (N_4363,N_3722,N_3002);
or U4364 (N_4364,N_3158,N_3436);
nand U4365 (N_4365,N_3079,N_3286);
or U4366 (N_4366,N_3097,N_3003);
nor U4367 (N_4367,N_3362,N_3315);
nor U4368 (N_4368,N_3053,N_3153);
nand U4369 (N_4369,N_3429,N_3347);
and U4370 (N_4370,N_3306,N_3080);
nand U4371 (N_4371,N_3744,N_3715);
nand U4372 (N_4372,N_3362,N_3350);
nand U4373 (N_4373,N_3204,N_3526);
and U4374 (N_4374,N_3556,N_3037);
xor U4375 (N_4375,N_3238,N_3138);
nand U4376 (N_4376,N_3094,N_3518);
nand U4377 (N_4377,N_3306,N_3166);
nand U4378 (N_4378,N_3722,N_3428);
and U4379 (N_4379,N_3419,N_3684);
or U4380 (N_4380,N_3009,N_3049);
nor U4381 (N_4381,N_3181,N_3322);
or U4382 (N_4382,N_3515,N_3290);
xor U4383 (N_4383,N_3632,N_3723);
nand U4384 (N_4384,N_3134,N_3660);
nor U4385 (N_4385,N_3591,N_3223);
nand U4386 (N_4386,N_3598,N_3391);
nand U4387 (N_4387,N_3083,N_3523);
or U4388 (N_4388,N_3548,N_3284);
and U4389 (N_4389,N_3520,N_3177);
and U4390 (N_4390,N_3558,N_3639);
or U4391 (N_4391,N_3531,N_3342);
nor U4392 (N_4392,N_3613,N_3128);
xnor U4393 (N_4393,N_3224,N_3650);
nand U4394 (N_4394,N_3294,N_3266);
or U4395 (N_4395,N_3478,N_3452);
or U4396 (N_4396,N_3702,N_3241);
or U4397 (N_4397,N_3328,N_3586);
or U4398 (N_4398,N_3361,N_3289);
nand U4399 (N_4399,N_3093,N_3365);
or U4400 (N_4400,N_3354,N_3551);
or U4401 (N_4401,N_3259,N_3420);
nand U4402 (N_4402,N_3356,N_3663);
or U4403 (N_4403,N_3476,N_3279);
or U4404 (N_4404,N_3234,N_3389);
or U4405 (N_4405,N_3714,N_3394);
xor U4406 (N_4406,N_3551,N_3681);
or U4407 (N_4407,N_3481,N_3598);
nor U4408 (N_4408,N_3548,N_3387);
and U4409 (N_4409,N_3641,N_3687);
or U4410 (N_4410,N_3436,N_3681);
and U4411 (N_4411,N_3631,N_3375);
nand U4412 (N_4412,N_3015,N_3693);
nor U4413 (N_4413,N_3490,N_3603);
or U4414 (N_4414,N_3080,N_3024);
nand U4415 (N_4415,N_3313,N_3040);
nor U4416 (N_4416,N_3145,N_3672);
or U4417 (N_4417,N_3259,N_3000);
nor U4418 (N_4418,N_3437,N_3588);
nor U4419 (N_4419,N_3171,N_3595);
and U4420 (N_4420,N_3527,N_3279);
and U4421 (N_4421,N_3388,N_3686);
or U4422 (N_4422,N_3691,N_3610);
nand U4423 (N_4423,N_3137,N_3155);
and U4424 (N_4424,N_3131,N_3401);
and U4425 (N_4425,N_3445,N_3061);
xnor U4426 (N_4426,N_3310,N_3565);
nor U4427 (N_4427,N_3497,N_3069);
nand U4428 (N_4428,N_3574,N_3633);
nor U4429 (N_4429,N_3021,N_3496);
nor U4430 (N_4430,N_3645,N_3133);
and U4431 (N_4431,N_3528,N_3429);
nor U4432 (N_4432,N_3637,N_3311);
nand U4433 (N_4433,N_3002,N_3500);
or U4434 (N_4434,N_3743,N_3279);
xor U4435 (N_4435,N_3088,N_3544);
nor U4436 (N_4436,N_3294,N_3707);
nand U4437 (N_4437,N_3731,N_3458);
nor U4438 (N_4438,N_3189,N_3467);
or U4439 (N_4439,N_3663,N_3412);
nand U4440 (N_4440,N_3611,N_3289);
or U4441 (N_4441,N_3005,N_3208);
and U4442 (N_4442,N_3314,N_3436);
and U4443 (N_4443,N_3524,N_3146);
nand U4444 (N_4444,N_3480,N_3286);
nor U4445 (N_4445,N_3008,N_3235);
nand U4446 (N_4446,N_3342,N_3476);
and U4447 (N_4447,N_3429,N_3671);
nor U4448 (N_4448,N_3003,N_3303);
and U4449 (N_4449,N_3192,N_3631);
nand U4450 (N_4450,N_3702,N_3474);
xnor U4451 (N_4451,N_3702,N_3009);
nand U4452 (N_4452,N_3182,N_3247);
or U4453 (N_4453,N_3384,N_3288);
and U4454 (N_4454,N_3075,N_3332);
nor U4455 (N_4455,N_3156,N_3501);
nand U4456 (N_4456,N_3629,N_3164);
nand U4457 (N_4457,N_3044,N_3083);
nand U4458 (N_4458,N_3177,N_3179);
xnor U4459 (N_4459,N_3173,N_3730);
nor U4460 (N_4460,N_3180,N_3173);
nor U4461 (N_4461,N_3237,N_3464);
nor U4462 (N_4462,N_3062,N_3321);
and U4463 (N_4463,N_3170,N_3037);
nor U4464 (N_4464,N_3358,N_3100);
xnor U4465 (N_4465,N_3230,N_3507);
xnor U4466 (N_4466,N_3450,N_3126);
or U4467 (N_4467,N_3744,N_3740);
nor U4468 (N_4468,N_3069,N_3287);
nor U4469 (N_4469,N_3537,N_3597);
nor U4470 (N_4470,N_3208,N_3313);
and U4471 (N_4471,N_3467,N_3588);
and U4472 (N_4472,N_3188,N_3462);
nor U4473 (N_4473,N_3531,N_3570);
and U4474 (N_4474,N_3037,N_3341);
or U4475 (N_4475,N_3000,N_3657);
or U4476 (N_4476,N_3705,N_3360);
xor U4477 (N_4477,N_3677,N_3228);
or U4478 (N_4478,N_3497,N_3349);
and U4479 (N_4479,N_3596,N_3451);
or U4480 (N_4480,N_3141,N_3593);
or U4481 (N_4481,N_3175,N_3202);
nor U4482 (N_4482,N_3580,N_3133);
or U4483 (N_4483,N_3341,N_3338);
or U4484 (N_4484,N_3217,N_3431);
nor U4485 (N_4485,N_3571,N_3159);
nor U4486 (N_4486,N_3052,N_3219);
nor U4487 (N_4487,N_3600,N_3296);
nor U4488 (N_4488,N_3371,N_3102);
xor U4489 (N_4489,N_3711,N_3226);
or U4490 (N_4490,N_3548,N_3209);
or U4491 (N_4491,N_3414,N_3519);
nand U4492 (N_4492,N_3128,N_3438);
nand U4493 (N_4493,N_3487,N_3528);
nor U4494 (N_4494,N_3386,N_3289);
and U4495 (N_4495,N_3620,N_3288);
and U4496 (N_4496,N_3623,N_3706);
xor U4497 (N_4497,N_3093,N_3648);
nor U4498 (N_4498,N_3103,N_3389);
and U4499 (N_4499,N_3291,N_3310);
nand U4500 (N_4500,N_4447,N_3966);
nand U4501 (N_4501,N_4158,N_4286);
nor U4502 (N_4502,N_4202,N_4009);
nand U4503 (N_4503,N_4124,N_4425);
or U4504 (N_4504,N_4255,N_4275);
and U4505 (N_4505,N_4274,N_4182);
nand U4506 (N_4506,N_4085,N_3773);
xor U4507 (N_4507,N_4317,N_4114);
nand U4508 (N_4508,N_3907,N_3780);
xor U4509 (N_4509,N_3892,N_3865);
or U4510 (N_4510,N_3790,N_4087);
xnor U4511 (N_4511,N_4363,N_4373);
or U4512 (N_4512,N_3847,N_3854);
and U4513 (N_4513,N_3950,N_4306);
or U4514 (N_4514,N_4352,N_4134);
nand U4515 (N_4515,N_3855,N_4184);
or U4516 (N_4516,N_4485,N_3868);
and U4517 (N_4517,N_3846,N_4066);
and U4518 (N_4518,N_4357,N_4028);
or U4519 (N_4519,N_4307,N_4246);
xnor U4520 (N_4520,N_4101,N_4208);
nor U4521 (N_4521,N_3893,N_4375);
nand U4522 (N_4522,N_4126,N_3861);
nor U4523 (N_4523,N_4461,N_3848);
or U4524 (N_4524,N_4444,N_3879);
and U4525 (N_4525,N_4106,N_4016);
nor U4526 (N_4526,N_4284,N_4350);
nand U4527 (N_4527,N_4043,N_4044);
and U4528 (N_4528,N_3962,N_4457);
nor U4529 (N_4529,N_4304,N_3774);
nor U4530 (N_4530,N_4390,N_4001);
and U4531 (N_4531,N_3810,N_4073);
or U4532 (N_4532,N_3984,N_4269);
nor U4533 (N_4533,N_4216,N_4088);
and U4534 (N_4534,N_3964,N_4418);
or U4535 (N_4535,N_3942,N_3838);
xor U4536 (N_4536,N_4256,N_4260);
xnor U4537 (N_4537,N_4039,N_4019);
nor U4538 (N_4538,N_3985,N_3806);
nand U4539 (N_4539,N_3993,N_4492);
and U4540 (N_4540,N_3763,N_4366);
nor U4541 (N_4541,N_4408,N_3822);
nor U4542 (N_4542,N_4163,N_3781);
nor U4543 (N_4543,N_4400,N_4151);
and U4544 (N_4544,N_3902,N_4293);
nand U4545 (N_4545,N_4041,N_4230);
nand U4546 (N_4546,N_3811,N_4113);
and U4547 (N_4547,N_4007,N_3786);
nand U4548 (N_4548,N_4078,N_3880);
xnor U4549 (N_4549,N_3851,N_4467);
or U4550 (N_4550,N_3949,N_3963);
nor U4551 (N_4551,N_3812,N_4416);
nor U4552 (N_4552,N_4322,N_4263);
nor U4553 (N_4553,N_3997,N_4038);
nor U4554 (N_4554,N_3795,N_4148);
or U4555 (N_4555,N_4086,N_4448);
and U4556 (N_4556,N_3759,N_4225);
nand U4557 (N_4557,N_4480,N_4091);
xnor U4558 (N_4558,N_4226,N_4292);
or U4559 (N_4559,N_4242,N_3989);
or U4560 (N_4560,N_4190,N_4189);
or U4561 (N_4561,N_3946,N_3927);
nor U4562 (N_4562,N_3986,N_4167);
xor U4563 (N_4563,N_3890,N_4445);
nor U4564 (N_4564,N_4334,N_3793);
nor U4565 (N_4565,N_3776,N_4470);
or U4566 (N_4566,N_4213,N_3955);
or U4567 (N_4567,N_3863,N_4254);
and U4568 (N_4568,N_4179,N_4355);
xnor U4569 (N_4569,N_4339,N_4077);
xor U4570 (N_4570,N_3754,N_4156);
nand U4571 (N_4571,N_4344,N_3778);
nand U4572 (N_4572,N_4389,N_4268);
or U4573 (N_4573,N_4396,N_4205);
and U4574 (N_4574,N_4080,N_4360);
nand U4575 (N_4575,N_4237,N_4311);
nand U4576 (N_4576,N_4098,N_4055);
nor U4577 (N_4577,N_4048,N_3850);
and U4578 (N_4578,N_4384,N_3978);
nor U4579 (N_4579,N_4361,N_4183);
and U4580 (N_4580,N_3899,N_4435);
or U4581 (N_4581,N_4328,N_4329);
and U4582 (N_4582,N_3797,N_4267);
nand U4583 (N_4583,N_4116,N_4280);
nor U4584 (N_4584,N_4288,N_3869);
or U4585 (N_4585,N_4207,N_3923);
or U4586 (N_4586,N_4194,N_3929);
xor U4587 (N_4587,N_4460,N_3906);
or U4588 (N_4588,N_4118,N_4025);
or U4589 (N_4589,N_4380,N_4325);
nor U4590 (N_4590,N_4424,N_4315);
nand U4591 (N_4591,N_4067,N_3836);
nand U4592 (N_4592,N_4115,N_3756);
and U4593 (N_4593,N_4450,N_4128);
and U4594 (N_4594,N_4359,N_4026);
or U4595 (N_4595,N_3867,N_4250);
xor U4596 (N_4596,N_3947,N_4111);
or U4597 (N_4597,N_4266,N_4058);
or U4598 (N_4598,N_4449,N_4229);
or U4599 (N_4599,N_4137,N_3829);
xnor U4600 (N_4600,N_4439,N_3901);
and U4601 (N_4601,N_4364,N_4348);
nor U4602 (N_4602,N_4238,N_4374);
and U4603 (N_4603,N_4013,N_4402);
or U4604 (N_4604,N_3877,N_3820);
or U4605 (N_4605,N_4217,N_4343);
or U4606 (N_4606,N_4321,N_3996);
or U4607 (N_4607,N_3948,N_4046);
nor U4608 (N_4608,N_4426,N_3991);
nand U4609 (N_4609,N_4022,N_3909);
and U4610 (N_4610,N_4429,N_3944);
xor U4611 (N_4611,N_4175,N_3956);
nor U4612 (N_4612,N_3804,N_4180);
and U4613 (N_4613,N_4029,N_4141);
xor U4614 (N_4614,N_4451,N_3803);
nand U4615 (N_4615,N_4309,N_3762);
or U4616 (N_4616,N_3925,N_4443);
and U4617 (N_4617,N_4469,N_4168);
nand U4618 (N_4618,N_4100,N_4428);
and U4619 (N_4619,N_3913,N_3826);
nand U4620 (N_4620,N_4056,N_4383);
or U4621 (N_4621,N_3873,N_4484);
nand U4622 (N_4622,N_4464,N_4232);
nand U4623 (N_4623,N_4104,N_3798);
and U4624 (N_4624,N_4102,N_3945);
xor U4625 (N_4625,N_4051,N_3788);
nor U4626 (N_4626,N_4454,N_4385);
xor U4627 (N_4627,N_3853,N_4161);
nor U4628 (N_4628,N_4214,N_3981);
or U4629 (N_4629,N_4365,N_3755);
or U4630 (N_4630,N_3932,N_4323);
nand U4631 (N_4631,N_3910,N_4024);
nand U4632 (N_4632,N_4169,N_4005);
or U4633 (N_4633,N_4412,N_4219);
nor U4634 (N_4634,N_4174,N_4145);
and U4635 (N_4635,N_4228,N_4171);
or U4636 (N_4636,N_3784,N_4218);
or U4637 (N_4637,N_4298,N_4079);
or U4638 (N_4638,N_4112,N_4065);
or U4639 (N_4639,N_4064,N_4082);
nor U4640 (N_4640,N_4291,N_3782);
nor U4641 (N_4641,N_3922,N_4072);
nand U4642 (N_4642,N_3878,N_3823);
nor U4643 (N_4643,N_3862,N_4040);
or U4644 (N_4644,N_4477,N_4057);
nor U4645 (N_4645,N_4089,N_4018);
nand U4646 (N_4646,N_4132,N_4392);
nor U4647 (N_4647,N_3887,N_4305);
nor U4648 (N_4648,N_4249,N_3939);
or U4649 (N_4649,N_3834,N_3957);
nand U4650 (N_4650,N_3919,N_4062);
nor U4651 (N_4651,N_3814,N_3928);
nor U4652 (N_4652,N_4473,N_4313);
and U4653 (N_4653,N_4209,N_3976);
and U4654 (N_4654,N_4068,N_4187);
nor U4655 (N_4655,N_4002,N_4281);
xnor U4656 (N_4656,N_3938,N_4204);
nand U4657 (N_4657,N_4060,N_3926);
or U4658 (N_4658,N_4369,N_4397);
xnor U4659 (N_4659,N_4481,N_4076);
and U4660 (N_4660,N_3915,N_4300);
and U4661 (N_4661,N_4338,N_3994);
or U4662 (N_4662,N_4493,N_4144);
and U4663 (N_4663,N_3783,N_4423);
nand U4664 (N_4664,N_4178,N_4193);
nand U4665 (N_4665,N_4422,N_4090);
xor U4666 (N_4666,N_4420,N_4020);
and U4667 (N_4667,N_3839,N_4410);
nor U4668 (N_4668,N_4170,N_4404);
or U4669 (N_4669,N_3785,N_4459);
and U4670 (N_4670,N_4053,N_4388);
or U4671 (N_4671,N_4192,N_4434);
xnor U4672 (N_4672,N_3882,N_4409);
xnor U4673 (N_4673,N_3914,N_4386);
nor U4674 (N_4674,N_3771,N_4117);
or U4675 (N_4675,N_4096,N_4143);
or U4676 (N_4676,N_3807,N_4149);
nor U4677 (N_4677,N_4346,N_4150);
nand U4678 (N_4678,N_4494,N_4059);
xnor U4679 (N_4679,N_4283,N_4047);
xor U4680 (N_4680,N_4395,N_4136);
nand U4681 (N_4681,N_3852,N_4382);
and U4682 (N_4682,N_3813,N_3886);
nor U4683 (N_4683,N_4140,N_4131);
or U4684 (N_4684,N_4071,N_4405);
nand U4685 (N_4685,N_3760,N_4463);
and U4686 (N_4686,N_4160,N_3982);
and U4687 (N_4687,N_4061,N_4378);
nand U4688 (N_4688,N_3970,N_4452);
xor U4689 (N_4689,N_4127,N_4456);
xor U4690 (N_4690,N_4474,N_3936);
or U4691 (N_4691,N_4004,N_3951);
nand U4692 (N_4692,N_3903,N_4271);
and U4693 (N_4693,N_3999,N_4153);
nand U4694 (N_4694,N_4475,N_3958);
or U4695 (N_4695,N_4272,N_4037);
and U4696 (N_4696,N_4109,N_4146);
or U4697 (N_4697,N_4222,N_3988);
nor U4698 (N_4698,N_3972,N_4406);
nor U4699 (N_4699,N_4121,N_3842);
nand U4700 (N_4700,N_4265,N_4239);
and U4701 (N_4701,N_3987,N_3832);
nand U4702 (N_4702,N_4133,N_3941);
or U4703 (N_4703,N_3775,N_3983);
or U4704 (N_4704,N_4027,N_4398);
nor U4705 (N_4705,N_3844,N_4297);
xor U4706 (N_4706,N_3897,N_4017);
and U4707 (N_4707,N_4310,N_3884);
nor U4708 (N_4708,N_4314,N_3753);
and U4709 (N_4709,N_3849,N_3874);
xor U4710 (N_4710,N_3857,N_4231);
or U4711 (N_4711,N_3905,N_4212);
and U4712 (N_4712,N_4342,N_4419);
and U4713 (N_4713,N_3864,N_4489);
xor U4714 (N_4714,N_3841,N_3750);
and U4715 (N_4715,N_3787,N_4433);
xor U4716 (N_4716,N_4142,N_3995);
or U4717 (N_4717,N_3881,N_4414);
and U4718 (N_4718,N_3791,N_4030);
or U4719 (N_4719,N_4277,N_4436);
nand U4720 (N_4720,N_3895,N_4496);
xor U4721 (N_4721,N_4279,N_3965);
xnor U4722 (N_4722,N_4221,N_4084);
nor U4723 (N_4723,N_3931,N_3830);
and U4724 (N_4724,N_3843,N_3770);
nand U4725 (N_4725,N_4455,N_4335);
nand U4726 (N_4726,N_4210,N_4251);
or U4727 (N_4727,N_4497,N_4036);
and U4728 (N_4728,N_4165,N_4241);
xnor U4729 (N_4729,N_4427,N_3967);
and U4730 (N_4730,N_4223,N_4401);
xnor U4731 (N_4731,N_4033,N_3889);
nand U4732 (N_4732,N_4248,N_4287);
and U4733 (N_4733,N_4370,N_4393);
xnor U4734 (N_4734,N_4308,N_3828);
or U4735 (N_4735,N_3757,N_4093);
and U4736 (N_4736,N_4139,N_3973);
or U4737 (N_4737,N_4302,N_4327);
nor U4738 (N_4738,N_4403,N_4159);
nand U4739 (N_4739,N_3917,N_4407);
and U4740 (N_4740,N_4472,N_4301);
or U4741 (N_4741,N_4495,N_4129);
nand U4742 (N_4742,N_4166,N_4276);
nand U4743 (N_4743,N_4234,N_4353);
or U4744 (N_4744,N_4176,N_3998);
nand U4745 (N_4745,N_4413,N_4188);
nor U4746 (N_4746,N_4379,N_4295);
and U4747 (N_4747,N_3959,N_4157);
nor U4748 (N_4748,N_4000,N_4391);
nand U4749 (N_4749,N_4356,N_3954);
nor U4750 (N_4750,N_4122,N_4340);
nor U4751 (N_4751,N_4482,N_4337);
nand U4752 (N_4752,N_4326,N_3870);
and U4753 (N_4753,N_3866,N_3856);
and U4754 (N_4754,N_4316,N_4367);
nor U4755 (N_4755,N_4432,N_4471);
or U4756 (N_4756,N_4211,N_3975);
and U4757 (N_4757,N_4012,N_4438);
nand U4758 (N_4758,N_4008,N_3875);
nand U4759 (N_4759,N_4490,N_4417);
and U4760 (N_4760,N_3827,N_4486);
xor U4761 (N_4761,N_3768,N_3819);
nor U4762 (N_4762,N_3960,N_4105);
or U4763 (N_4763,N_3896,N_3921);
nor U4764 (N_4764,N_3824,N_3968);
and U4765 (N_4765,N_3796,N_4487);
and U4766 (N_4766,N_4446,N_4362);
and U4767 (N_4767,N_3815,N_4282);
nand U4768 (N_4768,N_4345,N_4125);
nor U4769 (N_4769,N_3831,N_4387);
or U4770 (N_4770,N_4381,N_4240);
nor U4771 (N_4771,N_4319,N_4253);
xnor U4772 (N_4772,N_4011,N_4333);
nand U4773 (N_4773,N_4197,N_3908);
nand U4774 (N_4774,N_3801,N_4107);
or U4775 (N_4775,N_4154,N_4336);
nor U4776 (N_4776,N_4083,N_3920);
nand U4777 (N_4777,N_4247,N_4119);
xor U4778 (N_4778,N_4453,N_4050);
and U4779 (N_4779,N_4135,N_4479);
or U4780 (N_4780,N_4324,N_4354);
or U4781 (N_4781,N_4465,N_3833);
nand U4782 (N_4782,N_4172,N_3940);
or U4783 (N_4783,N_4262,N_4220);
nand U4784 (N_4784,N_4195,N_4476);
or U4785 (N_4785,N_4488,N_3952);
nor U4786 (N_4786,N_4185,N_3992);
xor U4787 (N_4787,N_3858,N_4014);
nand U4788 (N_4788,N_4290,N_3916);
or U4789 (N_4789,N_3953,N_3761);
and U4790 (N_4790,N_3794,N_4273);
or U4791 (N_4791,N_4318,N_4200);
nor U4792 (N_4792,N_4152,N_4270);
nor U4793 (N_4793,N_3800,N_4010);
and U4794 (N_4794,N_4094,N_4332);
or U4795 (N_4795,N_4289,N_4006);
nor U4796 (N_4796,N_3979,N_4070);
nor U4797 (N_4797,N_4458,N_4173);
nor U4798 (N_4798,N_4264,N_4349);
xnor U4799 (N_4799,N_3816,N_4162);
and U4800 (N_4800,N_3943,N_4278);
and U4801 (N_4801,N_4069,N_4035);
nand U4802 (N_4802,N_3751,N_4296);
nand U4803 (N_4803,N_4498,N_4442);
nor U4804 (N_4804,N_3980,N_3872);
nor U4805 (N_4805,N_4466,N_4063);
or U4806 (N_4806,N_4312,N_4206);
xor U4807 (N_4807,N_4331,N_4462);
nand U4808 (N_4808,N_4196,N_4372);
nor U4809 (N_4809,N_3752,N_4233);
or U4810 (N_4810,N_3918,N_4499);
and U4811 (N_4811,N_3825,N_4440);
or U4812 (N_4812,N_3792,N_4320);
nand U4813 (N_4813,N_3969,N_4478);
or U4814 (N_4814,N_4351,N_3990);
and U4815 (N_4815,N_4483,N_4181);
or U4816 (N_4816,N_3911,N_3817);
nor U4817 (N_4817,N_3779,N_4399);
and U4818 (N_4818,N_3924,N_4243);
nand U4819 (N_4819,N_4258,N_3758);
and U4820 (N_4820,N_4092,N_4034);
or U4821 (N_4821,N_3799,N_4252);
xor U4822 (N_4822,N_3809,N_4015);
or U4823 (N_4823,N_4468,N_4245);
and U4824 (N_4824,N_4186,N_4099);
or U4825 (N_4825,N_4377,N_4095);
nor U4826 (N_4826,N_4147,N_3937);
nand U4827 (N_4827,N_3766,N_4227);
nor U4828 (N_4828,N_3871,N_4358);
nand U4829 (N_4829,N_4376,N_3885);
nor U4830 (N_4830,N_3835,N_3845);
xor U4831 (N_4831,N_4074,N_4110);
and U4832 (N_4832,N_4120,N_3894);
xor U4833 (N_4833,N_4415,N_3805);
or U4834 (N_4834,N_4430,N_3802);
xnor U4835 (N_4835,N_4191,N_4054);
or U4836 (N_4836,N_4130,N_3935);
or U4837 (N_4837,N_4368,N_4123);
and U4838 (N_4838,N_4042,N_4003);
nand U4839 (N_4839,N_4032,N_4261);
nand U4840 (N_4840,N_4199,N_3961);
xor U4841 (N_4841,N_3840,N_4177);
and U4842 (N_4842,N_4441,N_4164);
nand U4843 (N_4843,N_4371,N_4299);
nor U4844 (N_4844,N_4437,N_3904);
nand U4845 (N_4845,N_3898,N_3974);
and U4846 (N_4846,N_4108,N_3912);
or U4847 (N_4847,N_3777,N_3764);
and U4848 (N_4848,N_3765,N_3821);
and U4849 (N_4849,N_4235,N_4303);
or U4850 (N_4850,N_4075,N_4201);
and U4851 (N_4851,N_3789,N_4491);
and U4852 (N_4852,N_4421,N_4081);
nand U4853 (N_4853,N_4155,N_3888);
and U4854 (N_4854,N_4052,N_4259);
xor U4855 (N_4855,N_3933,N_3818);
nor U4856 (N_4856,N_3837,N_4138);
or U4857 (N_4857,N_4244,N_4294);
or U4858 (N_4858,N_3808,N_3767);
nand U4859 (N_4859,N_3977,N_3859);
nand U4860 (N_4860,N_4198,N_4097);
xor U4861 (N_4861,N_4031,N_3971);
nand U4862 (N_4862,N_3934,N_4023);
nor U4863 (N_4863,N_3772,N_3769);
and U4864 (N_4864,N_4224,N_4049);
xor U4865 (N_4865,N_4236,N_3900);
xor U4866 (N_4866,N_3860,N_4341);
nand U4867 (N_4867,N_4257,N_3930);
nor U4868 (N_4868,N_4021,N_4394);
and U4869 (N_4869,N_4431,N_4411);
and U4870 (N_4870,N_4045,N_4103);
and U4871 (N_4871,N_4330,N_3876);
xnor U4872 (N_4872,N_4215,N_4285);
nand U4873 (N_4873,N_3891,N_4203);
nor U4874 (N_4874,N_4347,N_3883);
or U4875 (N_4875,N_4428,N_3815);
nand U4876 (N_4876,N_3827,N_4317);
or U4877 (N_4877,N_4397,N_3761);
and U4878 (N_4878,N_3833,N_4147);
or U4879 (N_4879,N_4044,N_3846);
and U4880 (N_4880,N_4487,N_4497);
nor U4881 (N_4881,N_4323,N_3750);
nand U4882 (N_4882,N_3909,N_3752);
or U4883 (N_4883,N_4415,N_3995);
and U4884 (N_4884,N_3803,N_4415);
nand U4885 (N_4885,N_4375,N_4419);
or U4886 (N_4886,N_3816,N_4209);
or U4887 (N_4887,N_4308,N_3985);
xor U4888 (N_4888,N_4362,N_3781);
xnor U4889 (N_4889,N_3778,N_4276);
nand U4890 (N_4890,N_3757,N_4417);
nand U4891 (N_4891,N_3918,N_3984);
and U4892 (N_4892,N_4485,N_3856);
nor U4893 (N_4893,N_3901,N_4366);
xnor U4894 (N_4894,N_4083,N_4310);
nand U4895 (N_4895,N_3849,N_3792);
or U4896 (N_4896,N_4190,N_4334);
and U4897 (N_4897,N_3806,N_4104);
and U4898 (N_4898,N_4278,N_3833);
or U4899 (N_4899,N_4344,N_4458);
nor U4900 (N_4900,N_4220,N_4295);
and U4901 (N_4901,N_4160,N_3936);
nor U4902 (N_4902,N_4353,N_3849);
nor U4903 (N_4903,N_3890,N_4314);
nand U4904 (N_4904,N_3772,N_3989);
nand U4905 (N_4905,N_4219,N_3996);
or U4906 (N_4906,N_3831,N_4375);
and U4907 (N_4907,N_3849,N_4102);
and U4908 (N_4908,N_4286,N_3951);
xor U4909 (N_4909,N_4321,N_4345);
xnor U4910 (N_4910,N_4134,N_4035);
nor U4911 (N_4911,N_4152,N_4084);
nor U4912 (N_4912,N_3827,N_4094);
or U4913 (N_4913,N_4005,N_3946);
nand U4914 (N_4914,N_4074,N_3751);
or U4915 (N_4915,N_4498,N_4448);
nor U4916 (N_4916,N_3806,N_4422);
xor U4917 (N_4917,N_3925,N_3911);
and U4918 (N_4918,N_3786,N_4290);
and U4919 (N_4919,N_4077,N_3837);
nand U4920 (N_4920,N_4132,N_4186);
nor U4921 (N_4921,N_4193,N_4472);
nand U4922 (N_4922,N_4010,N_3780);
nand U4923 (N_4923,N_3867,N_4230);
or U4924 (N_4924,N_3758,N_4143);
nor U4925 (N_4925,N_4083,N_4224);
xor U4926 (N_4926,N_3919,N_3778);
nand U4927 (N_4927,N_4311,N_4084);
and U4928 (N_4928,N_4165,N_3985);
xnor U4929 (N_4929,N_4210,N_4052);
nor U4930 (N_4930,N_4217,N_4028);
and U4931 (N_4931,N_3864,N_4033);
xor U4932 (N_4932,N_4373,N_4430);
and U4933 (N_4933,N_4483,N_4142);
nor U4934 (N_4934,N_3907,N_4082);
or U4935 (N_4935,N_4337,N_3987);
nor U4936 (N_4936,N_4013,N_4428);
nor U4937 (N_4937,N_4281,N_3929);
xor U4938 (N_4938,N_4285,N_3971);
or U4939 (N_4939,N_4364,N_3863);
or U4940 (N_4940,N_4172,N_3845);
nor U4941 (N_4941,N_4326,N_3988);
or U4942 (N_4942,N_4265,N_4459);
nand U4943 (N_4943,N_4181,N_4332);
nand U4944 (N_4944,N_3877,N_4179);
nor U4945 (N_4945,N_4362,N_3838);
xor U4946 (N_4946,N_4403,N_4457);
and U4947 (N_4947,N_3929,N_4185);
nand U4948 (N_4948,N_4098,N_3866);
and U4949 (N_4949,N_4318,N_4049);
nand U4950 (N_4950,N_4401,N_4464);
or U4951 (N_4951,N_4332,N_4490);
and U4952 (N_4952,N_4044,N_4187);
and U4953 (N_4953,N_4360,N_3815);
or U4954 (N_4954,N_4196,N_3955);
nand U4955 (N_4955,N_3916,N_4432);
or U4956 (N_4956,N_4012,N_3910);
and U4957 (N_4957,N_3981,N_4005);
nor U4958 (N_4958,N_3974,N_3792);
and U4959 (N_4959,N_4061,N_3854);
and U4960 (N_4960,N_4197,N_4355);
nand U4961 (N_4961,N_3752,N_3794);
nor U4962 (N_4962,N_3810,N_3998);
nand U4963 (N_4963,N_4167,N_4267);
nor U4964 (N_4964,N_3798,N_4075);
or U4965 (N_4965,N_3886,N_3775);
nor U4966 (N_4966,N_3984,N_4335);
nor U4967 (N_4967,N_4122,N_4321);
and U4968 (N_4968,N_3849,N_4267);
xnor U4969 (N_4969,N_4109,N_3753);
nand U4970 (N_4970,N_4393,N_4190);
nor U4971 (N_4971,N_4175,N_3915);
or U4972 (N_4972,N_4342,N_4251);
nand U4973 (N_4973,N_4212,N_3755);
nand U4974 (N_4974,N_4025,N_3840);
nand U4975 (N_4975,N_3981,N_3974);
nand U4976 (N_4976,N_4057,N_4389);
nand U4977 (N_4977,N_4359,N_4061);
nor U4978 (N_4978,N_4359,N_4363);
and U4979 (N_4979,N_3808,N_4181);
nor U4980 (N_4980,N_4009,N_3785);
or U4981 (N_4981,N_4001,N_4290);
xor U4982 (N_4982,N_4089,N_3915);
nor U4983 (N_4983,N_3859,N_4071);
nand U4984 (N_4984,N_4337,N_4452);
nand U4985 (N_4985,N_4283,N_3897);
or U4986 (N_4986,N_4107,N_4194);
and U4987 (N_4987,N_4383,N_3959);
nand U4988 (N_4988,N_4274,N_3943);
and U4989 (N_4989,N_4143,N_4374);
nand U4990 (N_4990,N_4085,N_3934);
nand U4991 (N_4991,N_4125,N_4203);
or U4992 (N_4992,N_4282,N_4243);
nand U4993 (N_4993,N_4469,N_4253);
nor U4994 (N_4994,N_3999,N_3968);
nor U4995 (N_4995,N_4246,N_4160);
or U4996 (N_4996,N_3818,N_4118);
nand U4997 (N_4997,N_4417,N_3987);
and U4998 (N_4998,N_4455,N_3974);
xnor U4999 (N_4999,N_4232,N_4359);
and U5000 (N_5000,N_4245,N_3769);
nor U5001 (N_5001,N_4307,N_4432);
nor U5002 (N_5002,N_4316,N_4448);
and U5003 (N_5003,N_4121,N_4302);
and U5004 (N_5004,N_3847,N_3756);
or U5005 (N_5005,N_4351,N_3865);
xnor U5006 (N_5006,N_3769,N_3784);
and U5007 (N_5007,N_4030,N_4097);
nand U5008 (N_5008,N_4351,N_4125);
xnor U5009 (N_5009,N_4192,N_4343);
nor U5010 (N_5010,N_4137,N_4243);
or U5011 (N_5011,N_4093,N_4275);
nand U5012 (N_5012,N_3926,N_4250);
or U5013 (N_5013,N_4021,N_4182);
or U5014 (N_5014,N_3925,N_3871);
or U5015 (N_5015,N_3797,N_4487);
and U5016 (N_5016,N_3932,N_3854);
nand U5017 (N_5017,N_4166,N_3966);
nand U5018 (N_5018,N_4370,N_3929);
or U5019 (N_5019,N_4325,N_3871);
xor U5020 (N_5020,N_4082,N_4375);
nand U5021 (N_5021,N_4403,N_4324);
nor U5022 (N_5022,N_4117,N_4062);
or U5023 (N_5023,N_4358,N_4339);
nor U5024 (N_5024,N_4444,N_3868);
nor U5025 (N_5025,N_4358,N_4248);
xnor U5026 (N_5026,N_4116,N_3841);
nand U5027 (N_5027,N_4327,N_3791);
nor U5028 (N_5028,N_3984,N_4401);
and U5029 (N_5029,N_3994,N_4335);
nand U5030 (N_5030,N_3956,N_3810);
and U5031 (N_5031,N_3960,N_4420);
and U5032 (N_5032,N_4434,N_4161);
or U5033 (N_5033,N_4217,N_4063);
nor U5034 (N_5034,N_4449,N_3974);
xor U5035 (N_5035,N_4298,N_4436);
and U5036 (N_5036,N_4293,N_4406);
nand U5037 (N_5037,N_4037,N_4310);
or U5038 (N_5038,N_3879,N_3983);
nand U5039 (N_5039,N_3841,N_4304);
nand U5040 (N_5040,N_4109,N_4009);
and U5041 (N_5041,N_4159,N_4182);
xor U5042 (N_5042,N_3936,N_3814);
xnor U5043 (N_5043,N_4248,N_4402);
and U5044 (N_5044,N_3826,N_3811);
nand U5045 (N_5045,N_4298,N_4159);
nand U5046 (N_5046,N_4379,N_4204);
and U5047 (N_5047,N_3851,N_4069);
xnor U5048 (N_5048,N_4310,N_3963);
nand U5049 (N_5049,N_4233,N_3758);
xor U5050 (N_5050,N_4430,N_3892);
and U5051 (N_5051,N_3974,N_3778);
or U5052 (N_5052,N_3967,N_3760);
and U5053 (N_5053,N_4298,N_3889);
nand U5054 (N_5054,N_4288,N_3751);
and U5055 (N_5055,N_4182,N_4451);
and U5056 (N_5056,N_4015,N_4246);
xor U5057 (N_5057,N_3956,N_3900);
or U5058 (N_5058,N_4001,N_4227);
nand U5059 (N_5059,N_3863,N_3878);
xor U5060 (N_5060,N_4219,N_3759);
nand U5061 (N_5061,N_4410,N_4431);
and U5062 (N_5062,N_3851,N_3965);
xnor U5063 (N_5063,N_4296,N_4147);
nor U5064 (N_5064,N_4096,N_4339);
and U5065 (N_5065,N_4204,N_3890);
nand U5066 (N_5066,N_3804,N_4478);
xnor U5067 (N_5067,N_4131,N_4255);
or U5068 (N_5068,N_4055,N_3826);
and U5069 (N_5069,N_4128,N_4048);
nand U5070 (N_5070,N_4449,N_3899);
nor U5071 (N_5071,N_3900,N_3974);
and U5072 (N_5072,N_3755,N_3913);
or U5073 (N_5073,N_4433,N_4174);
nand U5074 (N_5074,N_4443,N_3911);
and U5075 (N_5075,N_4171,N_3913);
nor U5076 (N_5076,N_4102,N_4247);
nand U5077 (N_5077,N_3960,N_4279);
or U5078 (N_5078,N_4087,N_4201);
and U5079 (N_5079,N_4432,N_4294);
or U5080 (N_5080,N_4370,N_4444);
nor U5081 (N_5081,N_4204,N_3856);
nor U5082 (N_5082,N_4359,N_4296);
nor U5083 (N_5083,N_4021,N_3770);
or U5084 (N_5084,N_4345,N_4411);
or U5085 (N_5085,N_4466,N_3908);
nand U5086 (N_5086,N_3810,N_4336);
or U5087 (N_5087,N_4209,N_3896);
and U5088 (N_5088,N_4349,N_3854);
or U5089 (N_5089,N_4391,N_4223);
and U5090 (N_5090,N_4443,N_4132);
nand U5091 (N_5091,N_3762,N_4247);
nand U5092 (N_5092,N_3946,N_3959);
nor U5093 (N_5093,N_3778,N_3910);
or U5094 (N_5094,N_3911,N_3755);
nor U5095 (N_5095,N_4167,N_4336);
nor U5096 (N_5096,N_4224,N_4017);
xor U5097 (N_5097,N_3916,N_4490);
and U5098 (N_5098,N_4284,N_4022);
nor U5099 (N_5099,N_4219,N_3962);
or U5100 (N_5100,N_4197,N_4494);
nand U5101 (N_5101,N_4099,N_3882);
or U5102 (N_5102,N_4101,N_3911);
or U5103 (N_5103,N_4405,N_3797);
nand U5104 (N_5104,N_4261,N_3976);
xnor U5105 (N_5105,N_4049,N_4408);
nor U5106 (N_5106,N_4155,N_4435);
or U5107 (N_5107,N_3919,N_4375);
nor U5108 (N_5108,N_3803,N_3804);
and U5109 (N_5109,N_4037,N_3815);
xnor U5110 (N_5110,N_3772,N_4348);
or U5111 (N_5111,N_4044,N_4210);
nor U5112 (N_5112,N_4020,N_4343);
or U5113 (N_5113,N_3856,N_4262);
or U5114 (N_5114,N_4102,N_3992);
and U5115 (N_5115,N_4090,N_4094);
or U5116 (N_5116,N_4297,N_4455);
nand U5117 (N_5117,N_4006,N_3849);
nand U5118 (N_5118,N_4489,N_4229);
nor U5119 (N_5119,N_3881,N_4351);
or U5120 (N_5120,N_4010,N_4219);
nand U5121 (N_5121,N_4143,N_4327);
and U5122 (N_5122,N_3965,N_3972);
and U5123 (N_5123,N_4217,N_4106);
and U5124 (N_5124,N_4097,N_4186);
nor U5125 (N_5125,N_4178,N_3837);
nor U5126 (N_5126,N_4175,N_4403);
nor U5127 (N_5127,N_4401,N_4494);
or U5128 (N_5128,N_4314,N_4049);
or U5129 (N_5129,N_3891,N_4111);
or U5130 (N_5130,N_4232,N_3844);
or U5131 (N_5131,N_3833,N_3863);
nand U5132 (N_5132,N_4460,N_4027);
nor U5133 (N_5133,N_4265,N_3939);
nor U5134 (N_5134,N_4442,N_4057);
and U5135 (N_5135,N_4278,N_3991);
nand U5136 (N_5136,N_4389,N_4018);
nor U5137 (N_5137,N_3874,N_4060);
nand U5138 (N_5138,N_3855,N_4354);
and U5139 (N_5139,N_4256,N_3961);
xnor U5140 (N_5140,N_3777,N_4274);
xor U5141 (N_5141,N_3837,N_4231);
and U5142 (N_5142,N_3772,N_4491);
nand U5143 (N_5143,N_4001,N_3797);
nor U5144 (N_5144,N_3923,N_3982);
nand U5145 (N_5145,N_4207,N_4114);
or U5146 (N_5146,N_3887,N_4232);
nand U5147 (N_5147,N_3794,N_3919);
and U5148 (N_5148,N_3881,N_4475);
and U5149 (N_5149,N_3890,N_4226);
or U5150 (N_5150,N_3935,N_4255);
nor U5151 (N_5151,N_3955,N_4304);
or U5152 (N_5152,N_4178,N_3775);
xnor U5153 (N_5153,N_4192,N_4175);
or U5154 (N_5154,N_3889,N_3780);
xor U5155 (N_5155,N_4365,N_4194);
or U5156 (N_5156,N_4411,N_3935);
nand U5157 (N_5157,N_3949,N_4062);
xor U5158 (N_5158,N_4428,N_3926);
and U5159 (N_5159,N_4116,N_4453);
or U5160 (N_5160,N_3876,N_4071);
nand U5161 (N_5161,N_4434,N_4325);
nand U5162 (N_5162,N_3751,N_4255);
or U5163 (N_5163,N_4344,N_4336);
and U5164 (N_5164,N_4322,N_3827);
and U5165 (N_5165,N_3969,N_4129);
nor U5166 (N_5166,N_4090,N_4336);
nand U5167 (N_5167,N_3958,N_4337);
and U5168 (N_5168,N_4163,N_4039);
or U5169 (N_5169,N_4246,N_4437);
nand U5170 (N_5170,N_4207,N_4069);
nand U5171 (N_5171,N_4187,N_4392);
or U5172 (N_5172,N_4485,N_4428);
nand U5173 (N_5173,N_3760,N_4002);
or U5174 (N_5174,N_4400,N_3840);
and U5175 (N_5175,N_4465,N_4036);
xnor U5176 (N_5176,N_4383,N_3900);
nand U5177 (N_5177,N_4381,N_4256);
nand U5178 (N_5178,N_3835,N_4038);
or U5179 (N_5179,N_3839,N_4227);
xnor U5180 (N_5180,N_4108,N_4455);
and U5181 (N_5181,N_3754,N_4314);
nor U5182 (N_5182,N_4139,N_3911);
nor U5183 (N_5183,N_3872,N_3856);
and U5184 (N_5184,N_3793,N_4280);
nor U5185 (N_5185,N_4109,N_3762);
xor U5186 (N_5186,N_4033,N_3937);
xnor U5187 (N_5187,N_4432,N_4475);
nor U5188 (N_5188,N_4443,N_4108);
nor U5189 (N_5189,N_4478,N_3918);
xor U5190 (N_5190,N_4238,N_4365);
and U5191 (N_5191,N_3869,N_3921);
or U5192 (N_5192,N_4034,N_3763);
nor U5193 (N_5193,N_4070,N_4270);
nor U5194 (N_5194,N_4065,N_4238);
nand U5195 (N_5195,N_4461,N_4449);
or U5196 (N_5196,N_4302,N_3766);
nand U5197 (N_5197,N_4430,N_4253);
and U5198 (N_5198,N_4200,N_3881);
nor U5199 (N_5199,N_3752,N_3753);
nor U5200 (N_5200,N_4059,N_3773);
or U5201 (N_5201,N_4157,N_4411);
or U5202 (N_5202,N_4292,N_4238);
and U5203 (N_5203,N_4143,N_3792);
nand U5204 (N_5204,N_4198,N_3923);
or U5205 (N_5205,N_4439,N_3792);
or U5206 (N_5206,N_4162,N_4113);
nor U5207 (N_5207,N_4136,N_4370);
nand U5208 (N_5208,N_4206,N_4038);
and U5209 (N_5209,N_4346,N_4060);
nor U5210 (N_5210,N_3799,N_3938);
nand U5211 (N_5211,N_3753,N_4432);
nor U5212 (N_5212,N_3796,N_3857);
and U5213 (N_5213,N_3936,N_3799);
nor U5214 (N_5214,N_4334,N_3901);
nand U5215 (N_5215,N_4144,N_3969);
nor U5216 (N_5216,N_3794,N_4345);
xor U5217 (N_5217,N_4008,N_4043);
xor U5218 (N_5218,N_3755,N_4000);
xnor U5219 (N_5219,N_3845,N_3961);
nand U5220 (N_5220,N_4371,N_4044);
and U5221 (N_5221,N_4347,N_3773);
or U5222 (N_5222,N_4464,N_4228);
nand U5223 (N_5223,N_4237,N_4443);
and U5224 (N_5224,N_3757,N_4219);
nor U5225 (N_5225,N_4249,N_4452);
xor U5226 (N_5226,N_4372,N_4074);
nand U5227 (N_5227,N_4433,N_3943);
nand U5228 (N_5228,N_4017,N_3924);
or U5229 (N_5229,N_3860,N_4010);
nor U5230 (N_5230,N_4222,N_4485);
nor U5231 (N_5231,N_4093,N_4168);
nor U5232 (N_5232,N_4183,N_3815);
and U5233 (N_5233,N_3854,N_4208);
nand U5234 (N_5234,N_4068,N_4260);
nand U5235 (N_5235,N_4322,N_4183);
and U5236 (N_5236,N_4334,N_4023);
nor U5237 (N_5237,N_4212,N_3943);
and U5238 (N_5238,N_4257,N_3762);
or U5239 (N_5239,N_3895,N_4215);
nor U5240 (N_5240,N_4243,N_4253);
nor U5241 (N_5241,N_3898,N_3866);
nor U5242 (N_5242,N_3936,N_3885);
nor U5243 (N_5243,N_4453,N_3891);
and U5244 (N_5244,N_3865,N_3853);
and U5245 (N_5245,N_4424,N_4401);
and U5246 (N_5246,N_4154,N_4253);
nand U5247 (N_5247,N_4293,N_4434);
or U5248 (N_5248,N_4461,N_3952);
nor U5249 (N_5249,N_4452,N_4311);
or U5250 (N_5250,N_4982,N_4624);
or U5251 (N_5251,N_5172,N_4645);
nor U5252 (N_5252,N_4844,N_5042);
nor U5253 (N_5253,N_5175,N_5048);
and U5254 (N_5254,N_5068,N_5064);
or U5255 (N_5255,N_5237,N_5101);
or U5256 (N_5256,N_5055,N_5173);
xnor U5257 (N_5257,N_4551,N_4590);
nand U5258 (N_5258,N_5244,N_4566);
or U5259 (N_5259,N_4570,N_4751);
nand U5260 (N_5260,N_4858,N_4579);
or U5261 (N_5261,N_4887,N_5009);
and U5262 (N_5262,N_4674,N_4602);
and U5263 (N_5263,N_5123,N_4730);
nand U5264 (N_5264,N_5032,N_4866);
and U5265 (N_5265,N_5243,N_4560);
and U5266 (N_5266,N_4512,N_4733);
nor U5267 (N_5267,N_4930,N_4665);
nor U5268 (N_5268,N_4817,N_4799);
nand U5269 (N_5269,N_4716,N_4905);
nand U5270 (N_5270,N_4564,N_4683);
nor U5271 (N_5271,N_4811,N_4500);
nand U5272 (N_5272,N_4853,N_5037);
nand U5273 (N_5273,N_4790,N_5211);
or U5274 (N_5274,N_4881,N_5215);
nor U5275 (N_5275,N_4802,N_4915);
nor U5276 (N_5276,N_4623,N_5153);
nand U5277 (N_5277,N_5223,N_4757);
or U5278 (N_5278,N_4535,N_4890);
nand U5279 (N_5279,N_5058,N_4876);
nand U5280 (N_5280,N_4552,N_4586);
nand U5281 (N_5281,N_4699,N_4988);
nand U5282 (N_5282,N_4949,N_4756);
nor U5283 (N_5283,N_4654,N_5246);
or U5284 (N_5284,N_4826,N_5219);
and U5285 (N_5285,N_5003,N_4720);
or U5286 (N_5286,N_4986,N_4712);
nand U5287 (N_5287,N_5231,N_4531);
and U5288 (N_5288,N_5072,N_5240);
xor U5289 (N_5289,N_4614,N_5146);
nand U5290 (N_5290,N_5004,N_4771);
xnor U5291 (N_5291,N_4565,N_4813);
nand U5292 (N_5292,N_4944,N_4837);
nor U5293 (N_5293,N_4934,N_4509);
and U5294 (N_5294,N_5018,N_4598);
and U5295 (N_5295,N_5171,N_4877);
or U5296 (N_5296,N_5029,N_5245);
and U5297 (N_5297,N_4774,N_4685);
nand U5298 (N_5298,N_5093,N_5138);
nand U5299 (N_5299,N_4516,N_4928);
nand U5300 (N_5300,N_4514,N_5145);
and U5301 (N_5301,N_4530,N_4554);
nand U5302 (N_5302,N_4873,N_4739);
and U5303 (N_5303,N_4687,N_5133);
nand U5304 (N_5304,N_4767,N_4561);
nand U5305 (N_5305,N_4798,N_5163);
or U5306 (N_5306,N_4763,N_4973);
nand U5307 (N_5307,N_4599,N_4562);
and U5308 (N_5308,N_5232,N_4611);
or U5309 (N_5309,N_5118,N_5141);
or U5310 (N_5310,N_5023,N_4888);
nor U5311 (N_5311,N_4882,N_4983);
xor U5312 (N_5312,N_4940,N_4929);
nor U5313 (N_5313,N_5155,N_5199);
and U5314 (N_5314,N_5229,N_5043);
or U5315 (N_5315,N_5051,N_5081);
or U5316 (N_5316,N_4825,N_4950);
and U5317 (N_5317,N_4926,N_4897);
xnor U5318 (N_5318,N_4854,N_4875);
xnor U5319 (N_5319,N_5082,N_5095);
nand U5320 (N_5320,N_4847,N_5194);
xor U5321 (N_5321,N_4738,N_5239);
and U5322 (N_5322,N_4886,N_4870);
xnor U5323 (N_5323,N_4996,N_4542);
nor U5324 (N_5324,N_5174,N_4960);
nand U5325 (N_5325,N_5247,N_5170);
and U5326 (N_5326,N_5184,N_4842);
nor U5327 (N_5327,N_5125,N_4852);
or U5328 (N_5328,N_4731,N_4839);
and U5329 (N_5329,N_4816,N_4613);
or U5330 (N_5330,N_5191,N_5067);
or U5331 (N_5331,N_4788,N_4723);
nor U5332 (N_5332,N_5120,N_4903);
nor U5333 (N_5333,N_5070,N_5022);
nor U5334 (N_5334,N_4504,N_4697);
nor U5335 (N_5335,N_4959,N_4804);
nor U5336 (N_5336,N_4513,N_4729);
nor U5337 (N_5337,N_4506,N_4834);
and U5338 (N_5338,N_4917,N_5090);
nor U5339 (N_5339,N_5063,N_4503);
and U5340 (N_5340,N_5096,N_4991);
nor U5341 (N_5341,N_4860,N_5105);
nor U5342 (N_5342,N_4908,N_4748);
or U5343 (N_5343,N_5135,N_5014);
or U5344 (N_5344,N_5012,N_4728);
nor U5345 (N_5345,N_4622,N_5080);
nand U5346 (N_5346,N_4750,N_5097);
nand U5347 (N_5347,N_4732,N_4688);
nand U5348 (N_5348,N_4931,N_5034);
or U5349 (N_5349,N_4898,N_4692);
nor U5350 (N_5350,N_5102,N_4533);
and U5351 (N_5351,N_5059,N_4544);
nor U5352 (N_5352,N_5179,N_4855);
and U5353 (N_5353,N_5234,N_5226);
nor U5354 (N_5354,N_4806,N_4777);
xnor U5355 (N_5355,N_5074,N_4810);
and U5356 (N_5356,N_4657,N_4938);
nor U5357 (N_5357,N_4606,N_4814);
nor U5358 (N_5358,N_4595,N_4902);
nand U5359 (N_5359,N_4721,N_4961);
nand U5360 (N_5360,N_4984,N_5188);
xor U5361 (N_5361,N_4563,N_4541);
nand U5362 (N_5362,N_4580,N_4828);
or U5363 (N_5363,N_4690,N_5176);
nor U5364 (N_5364,N_5186,N_4880);
nor U5365 (N_5365,N_4529,N_5006);
nand U5366 (N_5366,N_5001,N_4746);
or U5367 (N_5367,N_5065,N_4609);
xor U5368 (N_5368,N_5249,N_5156);
xnor U5369 (N_5369,N_5000,N_4724);
nor U5370 (N_5370,N_4762,N_5129);
nor U5371 (N_5371,N_5189,N_4936);
and U5372 (N_5372,N_5164,N_5121);
and U5373 (N_5373,N_5127,N_4608);
or U5374 (N_5374,N_5204,N_4753);
or U5375 (N_5375,N_4698,N_4987);
nor U5376 (N_5376,N_4523,N_4869);
nand U5377 (N_5377,N_4850,N_4932);
and U5378 (N_5378,N_4953,N_5166);
nor U5379 (N_5379,N_5104,N_4650);
nand U5380 (N_5380,N_4981,N_4964);
nand U5381 (N_5381,N_4913,N_5079);
or U5382 (N_5382,N_4838,N_4717);
nand U5383 (N_5383,N_4846,N_5106);
nand U5384 (N_5384,N_5036,N_4899);
xor U5385 (N_5385,N_4778,N_4643);
or U5386 (N_5386,N_4508,N_5035);
and U5387 (N_5387,N_4587,N_5002);
nor U5388 (N_5388,N_4768,N_5140);
or U5389 (N_5389,N_4661,N_5167);
nand U5390 (N_5390,N_4785,N_4822);
nand U5391 (N_5391,N_5196,N_4660);
or U5392 (N_5392,N_5057,N_5026);
and U5393 (N_5393,N_4628,N_4572);
and U5394 (N_5394,N_5033,N_4999);
or U5395 (N_5395,N_4998,N_4809);
or U5396 (N_5396,N_4710,N_5109);
or U5397 (N_5397,N_5031,N_4749);
nand U5398 (N_5398,N_4861,N_4689);
or U5399 (N_5399,N_4946,N_4911);
nand U5400 (N_5400,N_4947,N_5091);
nor U5401 (N_5401,N_4948,N_4555);
nor U5402 (N_5402,N_5132,N_5050);
nor U5403 (N_5403,N_4780,N_5152);
nor U5404 (N_5404,N_4863,N_4752);
nand U5405 (N_5405,N_4581,N_4968);
nand U5406 (N_5406,N_4538,N_4593);
and U5407 (N_5407,N_5200,N_4843);
or U5408 (N_5408,N_4795,N_4821);
or U5409 (N_5409,N_5025,N_4755);
nor U5410 (N_5410,N_4972,N_4568);
nand U5411 (N_5411,N_5089,N_4819);
nand U5412 (N_5412,N_5221,N_4528);
xnor U5413 (N_5413,N_4703,N_5021);
xor U5414 (N_5414,N_5078,N_4941);
nand U5415 (N_5415,N_4904,N_4620);
or U5416 (N_5416,N_4585,N_4640);
or U5417 (N_5417,N_5117,N_4823);
nor U5418 (N_5418,N_4607,N_4718);
nand U5419 (N_5419,N_5017,N_4715);
nor U5420 (N_5420,N_5169,N_4977);
nor U5421 (N_5421,N_4656,N_4994);
or U5422 (N_5422,N_4600,N_5061);
or U5423 (N_5423,N_4912,N_5128);
and U5424 (N_5424,N_5143,N_4796);
and U5425 (N_5425,N_5016,N_5147);
xor U5426 (N_5426,N_4740,N_4594);
or U5427 (N_5427,N_4652,N_4781);
nand U5428 (N_5428,N_5119,N_4651);
nand U5429 (N_5429,N_4833,N_4696);
nor U5430 (N_5430,N_4727,N_5041);
or U5431 (N_5431,N_5030,N_4976);
nand U5432 (N_5432,N_5013,N_5180);
or U5433 (N_5433,N_4965,N_5046);
nor U5434 (N_5434,N_4848,N_5149);
nand U5435 (N_5435,N_4889,N_4933);
and U5436 (N_5436,N_4558,N_5011);
nor U5437 (N_5437,N_4603,N_4922);
nor U5438 (N_5438,N_4663,N_4772);
nor U5439 (N_5439,N_4507,N_4942);
nor U5440 (N_5440,N_5069,N_4952);
or U5441 (N_5441,N_4575,N_4559);
nand U5442 (N_5442,N_4801,N_5040);
and U5443 (N_5443,N_4962,N_4537);
or U5444 (N_5444,N_5192,N_4662);
nand U5445 (N_5445,N_5183,N_5113);
or U5446 (N_5446,N_5075,N_4629);
or U5447 (N_5447,N_5224,N_4510);
nand U5448 (N_5448,N_4896,N_4892);
or U5449 (N_5449,N_5007,N_4631);
nand U5450 (N_5450,N_4787,N_5195);
and U5451 (N_5451,N_4671,N_4556);
nor U5452 (N_5452,N_4626,N_5098);
nor U5453 (N_5453,N_4879,N_5182);
nor U5454 (N_5454,N_4673,N_4666);
nand U5455 (N_5455,N_4857,N_4546);
nor U5456 (N_5456,N_4840,N_4789);
nor U5457 (N_5457,N_4805,N_4618);
or U5458 (N_5458,N_5187,N_5134);
or U5459 (N_5459,N_4951,N_5020);
nand U5460 (N_5460,N_4539,N_5136);
xor U5461 (N_5461,N_4784,N_4636);
nand U5462 (N_5462,N_4719,N_4578);
or U5463 (N_5463,N_4707,N_4792);
nor U5464 (N_5464,N_5197,N_4742);
or U5465 (N_5465,N_5099,N_4737);
and U5466 (N_5466,N_5100,N_4831);
and U5467 (N_5467,N_4791,N_5162);
nor U5468 (N_5468,N_4711,N_5216);
nand U5469 (N_5469,N_4591,N_5092);
xnor U5470 (N_5470,N_5227,N_4612);
or U5471 (N_5471,N_4963,N_4818);
and U5472 (N_5472,N_4734,N_4637);
or U5473 (N_5473,N_4970,N_4808);
and U5474 (N_5474,N_4937,N_5202);
or U5475 (N_5475,N_4989,N_4985);
nor U5476 (N_5476,N_5242,N_4759);
and U5477 (N_5477,N_5238,N_5203);
nand U5478 (N_5478,N_4701,N_4604);
and U5479 (N_5479,N_4865,N_4694);
xnor U5480 (N_5480,N_5193,N_4693);
or U5481 (N_5481,N_4829,N_5024);
nand U5482 (N_5482,N_4655,N_4522);
and U5483 (N_5483,N_4971,N_4681);
nor U5484 (N_5484,N_4680,N_4549);
nand U5485 (N_5485,N_5087,N_5045);
and U5486 (N_5486,N_5111,N_4800);
and U5487 (N_5487,N_4754,N_4534);
nor U5488 (N_5488,N_4916,N_4980);
nand U5489 (N_5489,N_4803,N_4874);
nand U5490 (N_5490,N_4573,N_4867);
nor U5491 (N_5491,N_5235,N_5178);
nor U5492 (N_5492,N_4764,N_5073);
xor U5493 (N_5493,N_4576,N_5124);
nor U5494 (N_5494,N_4939,N_4525);
nor U5495 (N_5495,N_5157,N_4884);
and U5496 (N_5496,N_4502,N_5177);
and U5497 (N_5497,N_4895,N_5206);
and U5498 (N_5498,N_5213,N_4668);
and U5499 (N_5499,N_4627,N_5233);
nand U5500 (N_5500,N_4747,N_5116);
nor U5501 (N_5501,N_4993,N_4862);
xor U5502 (N_5502,N_5112,N_4761);
nor U5503 (N_5503,N_4684,N_5148);
nand U5504 (N_5504,N_4505,N_4923);
nor U5505 (N_5505,N_4592,N_4894);
nor U5506 (N_5506,N_4616,N_4914);
nor U5507 (N_5507,N_4646,N_4871);
or U5508 (N_5508,N_4511,N_4649);
nor U5509 (N_5509,N_4714,N_4885);
nor U5510 (N_5510,N_4856,N_4659);
nand U5511 (N_5511,N_5010,N_5103);
and U5512 (N_5512,N_4824,N_4995);
nor U5513 (N_5513,N_4676,N_4954);
nand U5514 (N_5514,N_4550,N_4605);
nor U5515 (N_5515,N_5053,N_5160);
nor U5516 (N_5516,N_5208,N_4967);
or U5517 (N_5517,N_4569,N_5139);
nand U5518 (N_5518,N_4518,N_4519);
or U5519 (N_5519,N_5212,N_4807);
and U5520 (N_5520,N_5142,N_5114);
or U5521 (N_5521,N_5076,N_4708);
and U5522 (N_5522,N_4695,N_5218);
xor U5523 (N_5523,N_4625,N_5158);
or U5524 (N_5524,N_5060,N_4943);
nor U5525 (N_5525,N_4744,N_5062);
nor U5526 (N_5526,N_4969,N_4589);
or U5527 (N_5527,N_5052,N_4633);
or U5528 (N_5528,N_4935,N_4820);
and U5529 (N_5529,N_4582,N_5044);
and U5530 (N_5530,N_4526,N_4675);
or U5531 (N_5531,N_4957,N_5071);
nor U5532 (N_5532,N_4812,N_4638);
nor U5533 (N_5533,N_4864,N_4743);
or U5534 (N_5534,N_5094,N_4545);
nand U5535 (N_5535,N_4634,N_4849);
or U5536 (N_5536,N_4891,N_4722);
or U5537 (N_5537,N_4770,N_4765);
nand U5538 (N_5538,N_4745,N_4647);
nor U5539 (N_5539,N_4548,N_4900);
xnor U5540 (N_5540,N_4705,N_4691);
or U5541 (N_5541,N_5122,N_4540);
and U5542 (N_5542,N_4653,N_4845);
nand U5543 (N_5543,N_5110,N_4709);
nand U5544 (N_5544,N_5248,N_4741);
nand U5545 (N_5545,N_4735,N_5086);
nor U5546 (N_5546,N_4527,N_4678);
nand U5547 (N_5547,N_5056,N_5108);
xor U5548 (N_5548,N_5205,N_5115);
or U5549 (N_5549,N_4521,N_5154);
or U5550 (N_5550,N_4974,N_5126);
nor U5551 (N_5551,N_4966,N_4669);
nor U5552 (N_5552,N_5130,N_4793);
or U5553 (N_5553,N_4827,N_5054);
and U5554 (N_5554,N_4557,N_4574);
xnor U5555 (N_5555,N_5144,N_4520);
and U5556 (N_5556,N_5207,N_4658);
or U5557 (N_5557,N_4672,N_4990);
or U5558 (N_5558,N_4997,N_4664);
nand U5559 (N_5559,N_5161,N_4918);
nand U5560 (N_5560,N_4630,N_4677);
nand U5561 (N_5561,N_4835,N_4992);
nand U5562 (N_5562,N_4766,N_5159);
nand U5563 (N_5563,N_4584,N_5198);
or U5564 (N_5564,N_5083,N_4706);
xnor U5565 (N_5565,N_4776,N_4713);
or U5566 (N_5566,N_5201,N_4632);
or U5567 (N_5567,N_4920,N_5210);
xnor U5568 (N_5568,N_4515,N_5015);
nand U5569 (N_5569,N_4601,N_4883);
or U5570 (N_5570,N_5209,N_4779);
nand U5571 (N_5571,N_4567,N_4832);
nor U5572 (N_5572,N_4667,N_5049);
nand U5573 (N_5573,N_5088,N_5038);
and U5574 (N_5574,N_4919,N_4704);
nand U5575 (N_5575,N_4610,N_4958);
nor U5576 (N_5576,N_4644,N_4524);
xnor U5577 (N_5577,N_5220,N_4726);
nor U5578 (N_5578,N_4621,N_4830);
and U5579 (N_5579,N_4955,N_4925);
or U5580 (N_5580,N_4615,N_4682);
nand U5581 (N_5581,N_4725,N_5137);
xnor U5582 (N_5582,N_4909,N_5039);
xor U5583 (N_5583,N_4543,N_4769);
or U5584 (N_5584,N_4921,N_4907);
or U5585 (N_5585,N_4547,N_4872);
nand U5586 (N_5586,N_4670,N_4783);
and U5587 (N_5587,N_4786,N_4517);
or U5588 (N_5588,N_4906,N_4797);
xnor U5589 (N_5589,N_5228,N_4700);
nand U5590 (N_5590,N_4859,N_5084);
or U5591 (N_5591,N_4851,N_4841);
nand U5592 (N_5592,N_5028,N_5085);
nand U5593 (N_5593,N_5241,N_5230);
and U5594 (N_5594,N_4901,N_4760);
or U5595 (N_5595,N_4893,N_4639);
nand U5596 (N_5596,N_4583,N_4619);
nor U5597 (N_5597,N_5019,N_5008);
nor U5598 (N_5598,N_4775,N_4782);
xnor U5599 (N_5599,N_4577,N_5190);
nand U5600 (N_5600,N_4975,N_4956);
and U5601 (N_5601,N_5168,N_4553);
nor U5602 (N_5602,N_5107,N_4597);
and U5603 (N_5603,N_4815,N_4868);
nand U5604 (N_5604,N_4910,N_5185);
nor U5605 (N_5605,N_4617,N_5222);
xor U5606 (N_5606,N_4836,N_4532);
xor U5607 (N_5607,N_4635,N_5131);
or U5608 (N_5608,N_4927,N_4758);
and U5609 (N_5609,N_4773,N_5066);
and U5610 (N_5610,N_5165,N_5225);
nor U5611 (N_5611,N_5005,N_4571);
nor U5612 (N_5612,N_5236,N_4702);
or U5613 (N_5613,N_4978,N_4679);
nand U5614 (N_5614,N_5151,N_4588);
xnor U5615 (N_5615,N_5047,N_4686);
or U5616 (N_5616,N_5027,N_4878);
nor U5617 (N_5617,N_4536,N_5217);
or U5618 (N_5618,N_4924,N_4641);
nand U5619 (N_5619,N_5150,N_4979);
nand U5620 (N_5620,N_4596,N_5181);
nor U5621 (N_5621,N_4648,N_4945);
and U5622 (N_5622,N_5214,N_4736);
or U5623 (N_5623,N_4794,N_4642);
and U5624 (N_5624,N_5077,N_4501);
and U5625 (N_5625,N_5147,N_5010);
nand U5626 (N_5626,N_4991,N_4724);
nand U5627 (N_5627,N_5204,N_5205);
or U5628 (N_5628,N_4711,N_5043);
nand U5629 (N_5629,N_4756,N_4903);
or U5630 (N_5630,N_5030,N_4899);
and U5631 (N_5631,N_4648,N_5177);
nand U5632 (N_5632,N_4723,N_4702);
or U5633 (N_5633,N_4829,N_4681);
xnor U5634 (N_5634,N_5227,N_5171);
xor U5635 (N_5635,N_4820,N_4949);
and U5636 (N_5636,N_4867,N_4931);
nand U5637 (N_5637,N_4653,N_5227);
or U5638 (N_5638,N_4678,N_5164);
xor U5639 (N_5639,N_5125,N_4997);
or U5640 (N_5640,N_5148,N_4886);
xor U5641 (N_5641,N_4723,N_5148);
and U5642 (N_5642,N_5079,N_4501);
nand U5643 (N_5643,N_4792,N_4757);
and U5644 (N_5644,N_5100,N_5088);
xnor U5645 (N_5645,N_5234,N_4597);
or U5646 (N_5646,N_4649,N_4611);
and U5647 (N_5647,N_4870,N_4969);
nor U5648 (N_5648,N_5013,N_4802);
and U5649 (N_5649,N_5096,N_4800);
or U5650 (N_5650,N_4518,N_5192);
nand U5651 (N_5651,N_4870,N_4520);
nand U5652 (N_5652,N_5176,N_4768);
and U5653 (N_5653,N_4691,N_4964);
and U5654 (N_5654,N_4640,N_4834);
or U5655 (N_5655,N_4616,N_4757);
nor U5656 (N_5656,N_4952,N_4515);
nand U5657 (N_5657,N_4803,N_4973);
and U5658 (N_5658,N_5211,N_4888);
or U5659 (N_5659,N_5228,N_5046);
or U5660 (N_5660,N_4920,N_5045);
or U5661 (N_5661,N_4722,N_4994);
and U5662 (N_5662,N_4542,N_4828);
nor U5663 (N_5663,N_4823,N_4901);
nand U5664 (N_5664,N_5143,N_5097);
nand U5665 (N_5665,N_4998,N_4984);
xnor U5666 (N_5666,N_4925,N_5030);
nand U5667 (N_5667,N_4893,N_4621);
and U5668 (N_5668,N_5040,N_4642);
and U5669 (N_5669,N_4651,N_5081);
nor U5670 (N_5670,N_4671,N_4707);
nor U5671 (N_5671,N_4867,N_4651);
or U5672 (N_5672,N_5061,N_5012);
and U5673 (N_5673,N_5238,N_4846);
and U5674 (N_5674,N_4564,N_4970);
and U5675 (N_5675,N_5177,N_4952);
nor U5676 (N_5676,N_4963,N_4682);
or U5677 (N_5677,N_5189,N_4654);
and U5678 (N_5678,N_4696,N_4736);
nand U5679 (N_5679,N_5029,N_5189);
or U5680 (N_5680,N_5180,N_4917);
xnor U5681 (N_5681,N_5127,N_5025);
or U5682 (N_5682,N_4680,N_4646);
and U5683 (N_5683,N_4649,N_4633);
nand U5684 (N_5684,N_5192,N_4919);
and U5685 (N_5685,N_5027,N_4836);
or U5686 (N_5686,N_4888,N_4851);
or U5687 (N_5687,N_4683,N_4716);
or U5688 (N_5688,N_4535,N_4742);
and U5689 (N_5689,N_4628,N_5000);
nand U5690 (N_5690,N_5174,N_4732);
nor U5691 (N_5691,N_4960,N_4938);
or U5692 (N_5692,N_4846,N_4852);
or U5693 (N_5693,N_5036,N_4623);
xnor U5694 (N_5694,N_4764,N_4892);
xnor U5695 (N_5695,N_4738,N_5012);
nand U5696 (N_5696,N_4534,N_4710);
or U5697 (N_5697,N_4559,N_4502);
nor U5698 (N_5698,N_4609,N_5185);
nand U5699 (N_5699,N_4757,N_5247);
or U5700 (N_5700,N_5201,N_4530);
or U5701 (N_5701,N_4567,N_4889);
xor U5702 (N_5702,N_5070,N_4804);
and U5703 (N_5703,N_5199,N_4527);
and U5704 (N_5704,N_5086,N_4968);
nand U5705 (N_5705,N_4813,N_4659);
or U5706 (N_5706,N_5145,N_4891);
and U5707 (N_5707,N_4505,N_4906);
or U5708 (N_5708,N_4791,N_5030);
or U5709 (N_5709,N_4626,N_4908);
or U5710 (N_5710,N_5244,N_4512);
or U5711 (N_5711,N_5053,N_4981);
nor U5712 (N_5712,N_4506,N_5022);
or U5713 (N_5713,N_4501,N_5127);
or U5714 (N_5714,N_4883,N_5025);
or U5715 (N_5715,N_4981,N_5183);
or U5716 (N_5716,N_5204,N_4977);
nand U5717 (N_5717,N_4533,N_4886);
and U5718 (N_5718,N_4794,N_4557);
nor U5719 (N_5719,N_4641,N_4777);
nand U5720 (N_5720,N_5070,N_4777);
nor U5721 (N_5721,N_4778,N_4909);
nand U5722 (N_5722,N_4696,N_4843);
xnor U5723 (N_5723,N_4961,N_4945);
or U5724 (N_5724,N_5055,N_4801);
and U5725 (N_5725,N_4604,N_5092);
nand U5726 (N_5726,N_4800,N_5110);
nor U5727 (N_5727,N_4549,N_5215);
nand U5728 (N_5728,N_4577,N_4733);
nand U5729 (N_5729,N_5140,N_5230);
nor U5730 (N_5730,N_4552,N_5027);
or U5731 (N_5731,N_5051,N_4648);
nand U5732 (N_5732,N_5119,N_4788);
and U5733 (N_5733,N_4802,N_4572);
or U5734 (N_5734,N_5177,N_4733);
xor U5735 (N_5735,N_5191,N_5081);
and U5736 (N_5736,N_5104,N_5003);
or U5737 (N_5737,N_4705,N_4750);
nand U5738 (N_5738,N_4745,N_4792);
or U5739 (N_5739,N_5187,N_5192);
or U5740 (N_5740,N_4926,N_4656);
and U5741 (N_5741,N_4517,N_4584);
and U5742 (N_5742,N_5135,N_5244);
nor U5743 (N_5743,N_4649,N_4817);
and U5744 (N_5744,N_5042,N_4787);
and U5745 (N_5745,N_5046,N_4702);
and U5746 (N_5746,N_4862,N_4601);
and U5747 (N_5747,N_4767,N_4746);
nand U5748 (N_5748,N_5185,N_5104);
nand U5749 (N_5749,N_5248,N_5037);
and U5750 (N_5750,N_5022,N_4909);
nand U5751 (N_5751,N_4807,N_4727);
nand U5752 (N_5752,N_5110,N_5189);
nor U5753 (N_5753,N_4981,N_4890);
xnor U5754 (N_5754,N_5185,N_4908);
or U5755 (N_5755,N_5163,N_4710);
and U5756 (N_5756,N_4523,N_4688);
nand U5757 (N_5757,N_4998,N_5179);
or U5758 (N_5758,N_4673,N_4638);
nor U5759 (N_5759,N_5168,N_5097);
nand U5760 (N_5760,N_4715,N_4532);
and U5761 (N_5761,N_4681,N_4570);
nor U5762 (N_5762,N_4735,N_4602);
and U5763 (N_5763,N_5091,N_4933);
nor U5764 (N_5764,N_5105,N_5203);
nor U5765 (N_5765,N_4541,N_4688);
and U5766 (N_5766,N_5200,N_5009);
nor U5767 (N_5767,N_5229,N_5163);
nor U5768 (N_5768,N_4870,N_4762);
nand U5769 (N_5769,N_4664,N_4943);
xor U5770 (N_5770,N_4506,N_4529);
nand U5771 (N_5771,N_5040,N_4666);
or U5772 (N_5772,N_5179,N_4971);
xnor U5773 (N_5773,N_4979,N_4804);
nand U5774 (N_5774,N_5101,N_4733);
xnor U5775 (N_5775,N_4803,N_4926);
nor U5776 (N_5776,N_4573,N_5063);
xnor U5777 (N_5777,N_4541,N_4896);
nand U5778 (N_5778,N_4792,N_4848);
and U5779 (N_5779,N_4626,N_4815);
or U5780 (N_5780,N_5054,N_4869);
nor U5781 (N_5781,N_4634,N_4868);
nor U5782 (N_5782,N_4724,N_4566);
nand U5783 (N_5783,N_4863,N_4791);
nand U5784 (N_5784,N_4568,N_5017);
nand U5785 (N_5785,N_5150,N_4737);
nor U5786 (N_5786,N_5066,N_4820);
or U5787 (N_5787,N_4583,N_5149);
nor U5788 (N_5788,N_4896,N_4794);
xor U5789 (N_5789,N_4912,N_4811);
nor U5790 (N_5790,N_5173,N_4575);
nand U5791 (N_5791,N_4800,N_5200);
nor U5792 (N_5792,N_5091,N_4790);
nor U5793 (N_5793,N_4780,N_4633);
nor U5794 (N_5794,N_5249,N_5120);
nand U5795 (N_5795,N_4657,N_4769);
and U5796 (N_5796,N_4887,N_4738);
xor U5797 (N_5797,N_5019,N_5142);
nor U5798 (N_5798,N_4830,N_5217);
xnor U5799 (N_5799,N_5030,N_5039);
nor U5800 (N_5800,N_5188,N_4955);
nand U5801 (N_5801,N_5209,N_5191);
and U5802 (N_5802,N_5151,N_4744);
nor U5803 (N_5803,N_4859,N_5091);
and U5804 (N_5804,N_4572,N_4622);
or U5805 (N_5805,N_5184,N_4675);
nand U5806 (N_5806,N_4513,N_4924);
nor U5807 (N_5807,N_4798,N_4513);
nor U5808 (N_5808,N_4698,N_4717);
nand U5809 (N_5809,N_5074,N_4891);
nand U5810 (N_5810,N_4774,N_4656);
or U5811 (N_5811,N_4521,N_4544);
nor U5812 (N_5812,N_4799,N_5081);
nor U5813 (N_5813,N_4806,N_5001);
nor U5814 (N_5814,N_4569,N_4825);
nor U5815 (N_5815,N_5215,N_5121);
nand U5816 (N_5816,N_4517,N_4914);
nand U5817 (N_5817,N_5205,N_5126);
or U5818 (N_5818,N_5053,N_5221);
or U5819 (N_5819,N_5076,N_5169);
nor U5820 (N_5820,N_4638,N_4980);
xor U5821 (N_5821,N_5237,N_4924);
nand U5822 (N_5822,N_4884,N_4807);
nand U5823 (N_5823,N_5113,N_4947);
and U5824 (N_5824,N_4799,N_4509);
nor U5825 (N_5825,N_4511,N_4578);
nand U5826 (N_5826,N_4692,N_5155);
nor U5827 (N_5827,N_5147,N_4549);
or U5828 (N_5828,N_5072,N_4624);
nand U5829 (N_5829,N_4644,N_4835);
and U5830 (N_5830,N_5247,N_4834);
nor U5831 (N_5831,N_4617,N_4914);
and U5832 (N_5832,N_4567,N_5147);
nand U5833 (N_5833,N_5138,N_4718);
and U5834 (N_5834,N_4755,N_4968);
and U5835 (N_5835,N_4514,N_4854);
nor U5836 (N_5836,N_4558,N_5106);
nor U5837 (N_5837,N_4951,N_5022);
nor U5838 (N_5838,N_4958,N_4912);
or U5839 (N_5839,N_5173,N_5156);
and U5840 (N_5840,N_4724,N_4678);
and U5841 (N_5841,N_5160,N_4643);
xor U5842 (N_5842,N_4732,N_4783);
nand U5843 (N_5843,N_4542,N_4789);
nor U5844 (N_5844,N_5077,N_4733);
nor U5845 (N_5845,N_4762,N_5151);
and U5846 (N_5846,N_4856,N_5070);
xor U5847 (N_5847,N_4551,N_4528);
nand U5848 (N_5848,N_5069,N_4864);
xnor U5849 (N_5849,N_5076,N_4706);
and U5850 (N_5850,N_5181,N_5174);
xor U5851 (N_5851,N_5104,N_4604);
and U5852 (N_5852,N_4515,N_5222);
xnor U5853 (N_5853,N_4838,N_4692);
or U5854 (N_5854,N_4994,N_4885);
xnor U5855 (N_5855,N_5093,N_4922);
nand U5856 (N_5856,N_4814,N_4635);
and U5857 (N_5857,N_4763,N_4737);
nor U5858 (N_5858,N_4684,N_5044);
or U5859 (N_5859,N_5209,N_5127);
or U5860 (N_5860,N_4796,N_5023);
nand U5861 (N_5861,N_4569,N_4573);
or U5862 (N_5862,N_5136,N_4854);
nor U5863 (N_5863,N_5170,N_4986);
nand U5864 (N_5864,N_4686,N_4518);
or U5865 (N_5865,N_4842,N_5008);
xnor U5866 (N_5866,N_5124,N_4958);
and U5867 (N_5867,N_5061,N_4852);
nand U5868 (N_5868,N_4869,N_4837);
or U5869 (N_5869,N_4849,N_5022);
or U5870 (N_5870,N_4971,N_4926);
and U5871 (N_5871,N_5109,N_4912);
and U5872 (N_5872,N_4516,N_4730);
nor U5873 (N_5873,N_4697,N_5149);
and U5874 (N_5874,N_5208,N_4871);
nand U5875 (N_5875,N_4765,N_5040);
or U5876 (N_5876,N_5030,N_5103);
nor U5877 (N_5877,N_4565,N_4821);
or U5878 (N_5878,N_4850,N_5030);
and U5879 (N_5879,N_5130,N_4852);
nor U5880 (N_5880,N_4876,N_5098);
and U5881 (N_5881,N_4630,N_4818);
nand U5882 (N_5882,N_4912,N_5033);
and U5883 (N_5883,N_5050,N_5024);
xnor U5884 (N_5884,N_4502,N_5114);
or U5885 (N_5885,N_4515,N_5115);
nand U5886 (N_5886,N_4665,N_4999);
xor U5887 (N_5887,N_5130,N_4564);
nor U5888 (N_5888,N_4624,N_4663);
and U5889 (N_5889,N_4598,N_4940);
nand U5890 (N_5890,N_5137,N_5206);
or U5891 (N_5891,N_4964,N_5045);
nand U5892 (N_5892,N_4577,N_5067);
xnor U5893 (N_5893,N_4968,N_4946);
or U5894 (N_5894,N_5080,N_5208);
xor U5895 (N_5895,N_4727,N_4662);
and U5896 (N_5896,N_4844,N_5065);
or U5897 (N_5897,N_4694,N_4905);
nand U5898 (N_5898,N_4588,N_5047);
nand U5899 (N_5899,N_4847,N_4799);
xnor U5900 (N_5900,N_5015,N_4669);
and U5901 (N_5901,N_4935,N_4951);
or U5902 (N_5902,N_4517,N_5094);
nor U5903 (N_5903,N_4690,N_5169);
and U5904 (N_5904,N_5057,N_5106);
nand U5905 (N_5905,N_4813,N_4651);
or U5906 (N_5906,N_5163,N_5136);
nor U5907 (N_5907,N_4932,N_4937);
xnor U5908 (N_5908,N_4866,N_4933);
xor U5909 (N_5909,N_4564,N_4733);
or U5910 (N_5910,N_4532,N_4753);
or U5911 (N_5911,N_4877,N_4577);
nand U5912 (N_5912,N_4569,N_5239);
xnor U5913 (N_5913,N_4557,N_4618);
nand U5914 (N_5914,N_5232,N_5169);
or U5915 (N_5915,N_5128,N_5004);
nor U5916 (N_5916,N_5147,N_5101);
nor U5917 (N_5917,N_4584,N_4841);
or U5918 (N_5918,N_4805,N_4870);
nand U5919 (N_5919,N_4569,N_4512);
or U5920 (N_5920,N_4851,N_4606);
nor U5921 (N_5921,N_4737,N_5116);
nand U5922 (N_5922,N_4783,N_5159);
nand U5923 (N_5923,N_4751,N_4785);
or U5924 (N_5924,N_5106,N_4906);
or U5925 (N_5925,N_4977,N_5097);
and U5926 (N_5926,N_4882,N_5035);
and U5927 (N_5927,N_5234,N_5152);
nor U5928 (N_5928,N_5204,N_4736);
or U5929 (N_5929,N_5035,N_5026);
nor U5930 (N_5930,N_4604,N_5086);
or U5931 (N_5931,N_4658,N_4522);
and U5932 (N_5932,N_5224,N_5025);
or U5933 (N_5933,N_4555,N_5076);
nor U5934 (N_5934,N_4927,N_4928);
and U5935 (N_5935,N_4969,N_4951);
nor U5936 (N_5936,N_4521,N_4543);
and U5937 (N_5937,N_5180,N_4708);
nor U5938 (N_5938,N_5227,N_4520);
nor U5939 (N_5939,N_4936,N_5080);
or U5940 (N_5940,N_4571,N_5066);
nor U5941 (N_5941,N_4529,N_4986);
or U5942 (N_5942,N_5101,N_4689);
xor U5943 (N_5943,N_4952,N_4587);
nand U5944 (N_5944,N_4516,N_4576);
nand U5945 (N_5945,N_4577,N_4811);
nor U5946 (N_5946,N_4989,N_4678);
nor U5947 (N_5947,N_5094,N_4554);
nor U5948 (N_5948,N_5189,N_5158);
nor U5949 (N_5949,N_4522,N_4597);
nor U5950 (N_5950,N_5015,N_4689);
xor U5951 (N_5951,N_5141,N_5109);
or U5952 (N_5952,N_4902,N_4869);
nor U5953 (N_5953,N_4972,N_4503);
xor U5954 (N_5954,N_4642,N_5025);
or U5955 (N_5955,N_4594,N_4716);
nand U5956 (N_5956,N_4884,N_4773);
or U5957 (N_5957,N_4904,N_4960);
or U5958 (N_5958,N_4984,N_5078);
xor U5959 (N_5959,N_4985,N_4906);
nor U5960 (N_5960,N_4512,N_4600);
or U5961 (N_5961,N_4553,N_5132);
nor U5962 (N_5962,N_5112,N_4814);
or U5963 (N_5963,N_4620,N_5144);
and U5964 (N_5964,N_4998,N_4686);
nand U5965 (N_5965,N_4831,N_4990);
nand U5966 (N_5966,N_5013,N_4515);
nand U5967 (N_5967,N_4725,N_4927);
and U5968 (N_5968,N_5189,N_4562);
and U5969 (N_5969,N_4674,N_4741);
nor U5970 (N_5970,N_4508,N_4857);
and U5971 (N_5971,N_4559,N_4872);
nor U5972 (N_5972,N_4954,N_4670);
xnor U5973 (N_5973,N_5205,N_5090);
or U5974 (N_5974,N_5124,N_5133);
and U5975 (N_5975,N_4681,N_4763);
and U5976 (N_5976,N_4823,N_4870);
nand U5977 (N_5977,N_4686,N_4989);
and U5978 (N_5978,N_4627,N_5118);
xnor U5979 (N_5979,N_4692,N_4508);
nand U5980 (N_5980,N_4531,N_4913);
nand U5981 (N_5981,N_5246,N_4596);
or U5982 (N_5982,N_4532,N_4771);
and U5983 (N_5983,N_4550,N_4960);
or U5984 (N_5984,N_4550,N_5170);
and U5985 (N_5985,N_4571,N_4559);
nand U5986 (N_5986,N_5196,N_5242);
nand U5987 (N_5987,N_5143,N_4671);
nor U5988 (N_5988,N_4698,N_5084);
or U5989 (N_5989,N_5041,N_4910);
or U5990 (N_5990,N_5016,N_5177);
and U5991 (N_5991,N_4764,N_4751);
nand U5992 (N_5992,N_4755,N_5135);
nor U5993 (N_5993,N_4743,N_4695);
nand U5994 (N_5994,N_4825,N_4529);
or U5995 (N_5995,N_5097,N_4662);
and U5996 (N_5996,N_4787,N_4993);
nor U5997 (N_5997,N_4814,N_4555);
nand U5998 (N_5998,N_4692,N_4950);
and U5999 (N_5999,N_5048,N_4560);
nor U6000 (N_6000,N_5786,N_5366);
and U6001 (N_6001,N_5765,N_5337);
or U6002 (N_6002,N_5349,N_5450);
xor U6003 (N_6003,N_5359,N_5660);
xnor U6004 (N_6004,N_5288,N_5296);
or U6005 (N_6005,N_5913,N_5512);
or U6006 (N_6006,N_5332,N_5980);
xor U6007 (N_6007,N_5603,N_5517);
nand U6008 (N_6008,N_5614,N_5827);
and U6009 (N_6009,N_5302,N_5292);
nand U6010 (N_6010,N_5942,N_5963);
nor U6011 (N_6011,N_5848,N_5283);
nand U6012 (N_6012,N_5699,N_5306);
and U6013 (N_6013,N_5350,N_5729);
or U6014 (N_6014,N_5979,N_5816);
nor U6015 (N_6015,N_5944,N_5489);
nand U6016 (N_6016,N_5703,N_5429);
xnor U6017 (N_6017,N_5537,N_5987);
nand U6018 (N_6018,N_5319,N_5281);
nor U6019 (N_6019,N_5778,N_5661);
or U6020 (N_6020,N_5779,N_5293);
nand U6021 (N_6021,N_5620,N_5635);
and U6022 (N_6022,N_5822,N_5863);
nand U6023 (N_6023,N_5839,N_5871);
and U6024 (N_6024,N_5356,N_5821);
and U6025 (N_6025,N_5462,N_5672);
and U6026 (N_6026,N_5837,N_5346);
and U6027 (N_6027,N_5738,N_5644);
nand U6028 (N_6028,N_5756,N_5955);
xnor U6029 (N_6029,N_5470,N_5485);
and U6030 (N_6030,N_5968,N_5448);
nor U6031 (N_6031,N_5264,N_5971);
or U6032 (N_6032,N_5618,N_5726);
and U6033 (N_6033,N_5745,N_5737);
nor U6034 (N_6034,N_5819,N_5328);
and U6035 (N_6035,N_5664,N_5555);
xor U6036 (N_6036,N_5425,N_5731);
or U6037 (N_6037,N_5803,N_5949);
or U6038 (N_6038,N_5565,N_5749);
xor U6039 (N_6039,N_5793,N_5289);
and U6040 (N_6040,N_5312,N_5260);
xnor U6041 (N_6041,N_5443,N_5627);
or U6042 (N_6042,N_5342,N_5970);
or U6043 (N_6043,N_5391,N_5585);
xor U6044 (N_6044,N_5907,N_5771);
nor U6045 (N_6045,N_5399,N_5277);
and U6046 (N_6046,N_5390,N_5624);
nand U6047 (N_6047,N_5256,N_5719);
or U6048 (N_6048,N_5297,N_5747);
and U6049 (N_6049,N_5453,N_5488);
or U6050 (N_6050,N_5958,N_5862);
and U6051 (N_6051,N_5788,N_5780);
nand U6052 (N_6052,N_5505,N_5768);
and U6053 (N_6053,N_5960,N_5322);
xnor U6054 (N_6054,N_5602,N_5697);
or U6055 (N_6055,N_5553,N_5683);
xor U6056 (N_6056,N_5910,N_5455);
or U6057 (N_6057,N_5835,N_5478);
nor U6058 (N_6058,N_5964,N_5886);
nor U6059 (N_6059,N_5690,N_5872);
nor U6060 (N_6060,N_5393,N_5671);
and U6061 (N_6061,N_5781,N_5647);
xnor U6062 (N_6062,N_5520,N_5906);
nand U6063 (N_6063,N_5305,N_5571);
nand U6064 (N_6064,N_5564,N_5775);
nand U6065 (N_6065,N_5414,N_5466);
nand U6066 (N_6066,N_5957,N_5344);
nor U6067 (N_6067,N_5576,N_5769);
nor U6068 (N_6068,N_5417,N_5789);
and U6069 (N_6069,N_5570,N_5665);
nand U6070 (N_6070,N_5891,N_5475);
xnor U6071 (N_6071,N_5885,N_5257);
nor U6072 (N_6072,N_5917,N_5654);
xor U6073 (N_6073,N_5606,N_5262);
or U6074 (N_6074,N_5392,N_5477);
and U6075 (N_6075,N_5834,N_5625);
nor U6076 (N_6076,N_5802,N_5945);
or U6077 (N_6077,N_5723,N_5557);
nand U6078 (N_6078,N_5687,N_5521);
xnor U6079 (N_6079,N_5996,N_5347);
nand U6080 (N_6080,N_5473,N_5762);
xor U6081 (N_6081,N_5932,N_5901);
nor U6082 (N_6082,N_5490,N_5432);
and U6083 (N_6083,N_5704,N_5330);
nand U6084 (N_6084,N_5852,N_5530);
nor U6085 (N_6085,N_5449,N_5652);
nand U6086 (N_6086,N_5582,N_5286);
and U6087 (N_6087,N_5298,N_5763);
nor U6088 (N_6088,N_5628,N_5975);
nand U6089 (N_6089,N_5377,N_5313);
xnor U6090 (N_6090,N_5799,N_5951);
xor U6091 (N_6091,N_5284,N_5581);
nor U6092 (N_6092,N_5501,N_5411);
nor U6093 (N_6093,N_5593,N_5572);
nand U6094 (N_6094,N_5589,N_5597);
nand U6095 (N_6095,N_5688,N_5609);
or U6096 (N_6096,N_5405,N_5755);
and U6097 (N_6097,N_5846,N_5373);
or U6098 (N_6098,N_5916,N_5977);
nor U6099 (N_6099,N_5875,N_5267);
nor U6100 (N_6100,N_5334,N_5805);
nor U6101 (N_6101,N_5685,N_5607);
and U6102 (N_6102,N_5725,N_5721);
or U6103 (N_6103,N_5587,N_5493);
nand U6104 (N_6104,N_5542,N_5543);
nand U6105 (N_6105,N_5989,N_5421);
and U6106 (N_6106,N_5546,N_5435);
nand U6107 (N_6107,N_5828,N_5985);
nor U6108 (N_6108,N_5577,N_5545);
or U6109 (N_6109,N_5991,N_5777);
or U6110 (N_6110,N_5732,N_5867);
or U6111 (N_6111,N_5526,N_5383);
and U6112 (N_6112,N_5472,N_5430);
nand U6113 (N_6113,N_5903,N_5634);
nand U6114 (N_6114,N_5919,N_5534);
or U6115 (N_6115,N_5608,N_5959);
and U6116 (N_6116,N_5622,N_5667);
and U6117 (N_6117,N_5743,N_5578);
or U6118 (N_6118,N_5908,N_5679);
nor U6119 (N_6119,N_5818,N_5295);
nand U6120 (N_6120,N_5385,N_5815);
nand U6121 (N_6121,N_5528,N_5981);
nand U6122 (N_6122,N_5255,N_5406);
and U6123 (N_6123,N_5573,N_5879);
xor U6124 (N_6124,N_5894,N_5857);
nand U6125 (N_6125,N_5533,N_5838);
nor U6126 (N_6126,N_5730,N_5978);
nand U6127 (N_6127,N_5809,N_5689);
nor U6128 (N_6128,N_5881,N_5454);
or U6129 (N_6129,N_5360,N_5817);
or U6130 (N_6130,N_5878,N_5317);
or U6131 (N_6131,N_5476,N_5965);
nor U6132 (N_6132,N_5870,N_5648);
nor U6133 (N_6133,N_5923,N_5850);
xor U6134 (N_6134,N_5860,N_5795);
nor U6135 (N_6135,N_5561,N_5351);
and U6136 (N_6136,N_5370,N_5403);
nor U6137 (N_6137,N_5586,N_5880);
nand U6138 (N_6138,N_5378,N_5864);
nor U6139 (N_6139,N_5458,N_5469);
and U6140 (N_6140,N_5794,N_5339);
or U6141 (N_6141,N_5630,N_5909);
and U6142 (N_6142,N_5467,N_5995);
xnor U6143 (N_6143,N_5890,N_5532);
nand U6144 (N_6144,N_5408,N_5540);
nor U6145 (N_6145,N_5251,N_5943);
nor U6146 (N_6146,N_5904,N_5278);
nor U6147 (N_6147,N_5365,N_5253);
xnor U6148 (N_6148,N_5952,N_5282);
nand U6149 (N_6149,N_5670,N_5424);
nor U6150 (N_6150,N_5820,N_5439);
nand U6151 (N_6151,N_5858,N_5927);
or U6152 (N_6152,N_5826,N_5669);
xor U6153 (N_6153,N_5787,N_5524);
and U6154 (N_6154,N_5736,N_5518);
nor U6155 (N_6155,N_5442,N_5426);
nor U6156 (N_6156,N_5568,N_5343);
nor U6157 (N_6157,N_5333,N_5633);
or U6158 (N_6158,N_5928,N_5479);
nand U6159 (N_6159,N_5836,N_5931);
xor U6160 (N_6160,N_5427,N_5884);
or U6161 (N_6161,N_5735,N_5642);
xor U6162 (N_6162,N_5559,N_5619);
nor U6163 (N_6163,N_5659,N_5481);
or U6164 (N_6164,N_5655,N_5937);
nor U6165 (N_6165,N_5722,N_5918);
xnor U6166 (N_6166,N_5324,N_5547);
nand U6167 (N_6167,N_5291,N_5601);
or U6168 (N_6168,N_5386,N_5680);
and U6169 (N_6169,N_5759,N_5536);
nor U6170 (N_6170,N_5861,N_5596);
and U6171 (N_6171,N_5428,N_5746);
nor U6172 (N_6172,N_5384,N_5700);
and U6173 (N_6173,N_5474,N_5847);
nor U6174 (N_6174,N_5259,N_5309);
and U6175 (N_6175,N_5357,N_5389);
nand U6176 (N_6176,N_5897,N_5849);
xnor U6177 (N_6177,N_5716,N_5701);
xor U6178 (N_6178,N_5315,N_5468);
nand U6179 (N_6179,N_5783,N_5832);
xnor U6180 (N_6180,N_5588,N_5420);
and U6181 (N_6181,N_5776,N_5668);
and U6182 (N_6182,N_5640,N_5329);
or U6183 (N_6183,N_5922,N_5492);
xnor U6184 (N_6184,N_5560,N_5280);
xnor U6185 (N_6185,N_5463,N_5465);
or U6186 (N_6186,N_5415,N_5967);
xnor U6187 (N_6187,N_5326,N_5446);
or U6188 (N_6188,N_5926,N_5705);
or U6189 (N_6189,N_5263,N_5696);
and U6190 (N_6190,N_5503,N_5623);
nand U6191 (N_6191,N_5869,N_5791);
nand U6192 (N_6192,N_5613,N_5912);
nor U6193 (N_6193,N_5767,N_5308);
or U6194 (N_6194,N_5374,N_5873);
xor U6195 (N_6195,N_5921,N_5760);
or U6196 (N_6196,N_5754,N_5375);
and U6197 (N_6197,N_5531,N_5814);
xnor U6198 (N_6198,N_5947,N_5484);
nor U6199 (N_6199,N_5720,N_5457);
or U6200 (N_6200,N_5676,N_5398);
nand U6201 (N_6201,N_5254,N_5973);
and U6202 (N_6202,N_5639,N_5591);
nand U6203 (N_6203,N_5341,N_5379);
and U6204 (N_6204,N_5303,N_5636);
nand U6205 (N_6205,N_5956,N_5632);
nand U6206 (N_6206,N_5666,N_5831);
nand U6207 (N_6207,N_5742,N_5480);
or U6208 (N_6208,N_5495,N_5395);
and U6209 (N_6209,N_5681,N_5686);
xor U6210 (N_6210,N_5452,N_5434);
and U6211 (N_6211,N_5482,N_5539);
and U6212 (N_6212,N_5372,N_5707);
nor U6213 (N_6213,N_5500,N_5299);
or U6214 (N_6214,N_5272,N_5615);
nand U6215 (N_6215,N_5962,N_5276);
or U6216 (N_6216,N_5840,N_5810);
or U6217 (N_6217,N_5724,N_5311);
nor U6218 (N_6218,N_5905,N_5519);
nand U6219 (N_6219,N_5829,N_5307);
or U6220 (N_6220,N_5874,N_5999);
xor U6221 (N_6221,N_5715,N_5400);
or U6222 (N_6222,N_5527,N_5456);
xor U6223 (N_6223,N_5662,N_5833);
or U6224 (N_6224,N_5274,N_5290);
nor U6225 (N_6225,N_5785,N_5541);
and U6226 (N_6226,N_5883,N_5300);
nand U6227 (N_6227,N_5656,N_5711);
nand U6228 (N_6228,N_5764,N_5580);
nor U6229 (N_6229,N_5914,N_5790);
and U6230 (N_6230,N_5598,N_5510);
nand U6231 (N_6231,N_5961,N_5604);
xor U6232 (N_6232,N_5948,N_5807);
and U6233 (N_6233,N_5562,N_5388);
nor U6234 (N_6234,N_5859,N_5695);
nand U6235 (N_6235,N_5507,N_5674);
nor U6236 (N_6236,N_5325,N_5751);
or U6237 (N_6237,N_5605,N_5407);
or U6238 (N_6238,N_5354,N_5941);
nor U6239 (N_6239,N_5946,N_5516);
and U6240 (N_6240,N_5853,N_5486);
xor U6241 (N_6241,N_5447,N_5953);
or U6242 (N_6242,N_5892,N_5252);
and U6243 (N_6243,N_5766,N_5250);
nand U6244 (N_6244,N_5461,N_5882);
or U6245 (N_6245,N_5929,N_5772);
or U6246 (N_6246,N_5369,N_5525);
or U6247 (N_6247,N_5631,N_5784);
and U6248 (N_6248,N_5851,N_5898);
nor U6249 (N_6249,N_5992,N_5436);
or U6250 (N_6250,N_5397,N_5899);
xor U6251 (N_6251,N_5323,N_5331);
or U6252 (N_6252,N_5800,N_5595);
or U6253 (N_6253,N_5413,N_5287);
and U6254 (N_6254,N_5544,N_5404);
nand U6255 (N_6255,N_5431,N_5646);
nand U6256 (N_6256,N_5896,N_5352);
nor U6257 (N_6257,N_5739,N_5804);
and U6258 (N_6258,N_5362,N_5511);
or U6259 (N_6259,N_5645,N_5499);
or U6260 (N_6260,N_5855,N_5717);
or U6261 (N_6261,N_5502,N_5900);
nor U6262 (N_6262,N_5693,N_5782);
or U6263 (N_6263,N_5529,N_5911);
nand U6264 (N_6264,N_5998,N_5355);
and U6265 (N_6265,N_5677,N_5638);
and U6266 (N_6266,N_5269,N_5651);
or U6267 (N_6267,N_5550,N_5773);
and U6268 (N_6268,N_5423,N_5552);
or U6269 (N_6269,N_5844,N_5574);
or U6270 (N_6270,N_5318,N_5514);
and U6271 (N_6271,N_5774,N_5364);
xnor U6272 (N_6272,N_5641,N_5994);
nor U6273 (N_6273,N_5348,N_5509);
and U6274 (N_6274,N_5753,N_5925);
nor U6275 (N_6275,N_5265,N_5702);
nor U6276 (N_6276,N_5438,N_5444);
or U6277 (N_6277,N_5433,N_5744);
nor U6278 (N_6278,N_5491,N_5865);
nand U6279 (N_6279,N_5441,N_5376);
or U6280 (N_6280,N_5361,N_5599);
and U6281 (N_6281,N_5902,N_5549);
nand U6282 (N_6282,N_5682,N_5498);
and U6283 (N_6283,N_5611,N_5437);
nand U6284 (N_6284,N_5972,N_5506);
and U6285 (N_6285,N_5841,N_5924);
nand U6286 (N_6286,N_5842,N_5445);
nor U6287 (N_6287,N_5401,N_5367);
or U6288 (N_6288,N_5757,N_5321);
nand U6289 (N_6289,N_5584,N_5983);
and U6290 (N_6290,N_5740,N_5460);
nand U6291 (N_6291,N_5694,N_5915);
xor U6292 (N_6292,N_5824,N_5387);
or U6293 (N_6293,N_5513,N_5380);
and U6294 (N_6294,N_5988,N_5273);
or U6295 (N_6295,N_5984,N_5416);
nand U6296 (N_6296,N_5974,N_5698);
nor U6297 (N_6297,N_5930,N_5600);
nor U6298 (N_6298,N_5617,N_5410);
and U6299 (N_6299,N_5653,N_5637);
xnor U6300 (N_6300,N_5830,N_5275);
nand U6301 (N_6301,N_5718,N_5396);
or U6302 (N_6302,N_5806,N_5320);
and U6303 (N_6303,N_5657,N_5658);
xor U6304 (N_6304,N_5797,N_5579);
nor U6305 (N_6305,N_5451,N_5301);
nand U6306 (N_6306,N_5621,N_5798);
or U6307 (N_6307,N_5515,N_5304);
or U6308 (N_6308,N_5548,N_5792);
nor U6309 (N_6309,N_5394,N_5440);
xnor U6310 (N_6310,N_5338,N_5535);
or U6311 (N_6311,N_5261,N_5340);
or U6312 (N_6312,N_5496,N_5990);
xor U6313 (N_6313,N_5734,N_5643);
xnor U6314 (N_6314,N_5649,N_5728);
nand U6315 (N_6315,N_5748,N_5663);
nor U6316 (N_6316,N_5368,N_5310);
nor U6317 (N_6317,N_5629,N_5418);
nand U6318 (N_6318,N_5583,N_5856);
or U6319 (N_6319,N_5678,N_5712);
nor U6320 (N_6320,N_5402,N_5626);
and U6321 (N_6321,N_5692,N_5345);
xor U6322 (N_6322,N_5887,N_5522);
nor U6323 (N_6323,N_5268,N_5866);
or U6324 (N_6324,N_5616,N_5733);
or U6325 (N_6325,N_5675,N_5854);
nor U6326 (N_6326,N_5314,N_5808);
nand U6327 (N_6327,N_5982,N_5868);
and U6328 (N_6328,N_5327,N_5936);
nand U6329 (N_6329,N_5270,N_5706);
or U6330 (N_6330,N_5567,N_5483);
or U6331 (N_6331,N_5823,N_5710);
nand U6332 (N_6332,N_5566,N_5538);
or U6333 (N_6333,N_5714,N_5487);
or U6334 (N_6334,N_5813,N_5294);
and U6335 (N_6335,N_5812,N_5523);
and U6336 (N_6336,N_5708,N_5895);
xor U6337 (N_6337,N_5508,N_5494);
or U6338 (N_6338,N_5563,N_5336);
xnor U6339 (N_6339,N_5876,N_5843);
nor U6340 (N_6340,N_5612,N_5569);
or U6341 (N_6341,N_5825,N_5684);
or U6342 (N_6342,N_5422,N_5993);
nor U6343 (N_6343,N_5471,N_5933);
nand U6344 (N_6344,N_5419,N_5575);
and U6345 (N_6345,N_5381,N_5382);
nand U6346 (N_6346,N_5558,N_5363);
nor U6347 (N_6347,N_5371,N_5889);
nor U6348 (N_6348,N_5940,N_5412);
and U6349 (N_6349,N_5741,N_5969);
xor U6350 (N_6350,N_5594,N_5770);
and U6351 (N_6351,N_5279,N_5258);
or U6352 (N_6352,N_5650,N_5920);
nand U6353 (N_6353,N_5554,N_5758);
or U6354 (N_6354,N_5504,N_5888);
nand U6355 (N_6355,N_5590,N_5335);
nand U6356 (N_6356,N_5709,N_5845);
and U6357 (N_6357,N_5939,N_5464);
nand U6358 (N_6358,N_5935,N_5592);
or U6359 (N_6359,N_5752,N_5691);
and U6360 (N_6360,N_5976,N_5497);
and U6361 (N_6361,N_5938,N_5727);
nor U6362 (N_6362,N_5893,N_5358);
nor U6363 (N_6363,N_5610,N_5551);
xnor U6364 (N_6364,N_5811,N_5966);
or U6365 (N_6365,N_5409,N_5801);
nand U6366 (N_6366,N_5877,N_5761);
nor U6367 (N_6367,N_5266,N_5459);
xor U6368 (N_6368,N_5353,N_5796);
nand U6369 (N_6369,N_5986,N_5285);
and U6370 (N_6370,N_5934,N_5954);
nand U6371 (N_6371,N_5997,N_5750);
or U6372 (N_6372,N_5316,N_5950);
and U6373 (N_6373,N_5556,N_5713);
and U6374 (N_6374,N_5271,N_5673);
or U6375 (N_6375,N_5369,N_5664);
or U6376 (N_6376,N_5471,N_5430);
xnor U6377 (N_6377,N_5479,N_5450);
and U6378 (N_6378,N_5967,N_5857);
nor U6379 (N_6379,N_5947,N_5823);
or U6380 (N_6380,N_5446,N_5364);
or U6381 (N_6381,N_5900,N_5447);
nand U6382 (N_6382,N_5352,N_5444);
nor U6383 (N_6383,N_5450,N_5453);
nand U6384 (N_6384,N_5773,N_5827);
nand U6385 (N_6385,N_5684,N_5918);
nand U6386 (N_6386,N_5458,N_5541);
and U6387 (N_6387,N_5877,N_5779);
and U6388 (N_6388,N_5409,N_5811);
and U6389 (N_6389,N_5721,N_5958);
or U6390 (N_6390,N_5371,N_5852);
xor U6391 (N_6391,N_5484,N_5327);
nand U6392 (N_6392,N_5707,N_5673);
nor U6393 (N_6393,N_5732,N_5905);
or U6394 (N_6394,N_5401,N_5458);
xor U6395 (N_6395,N_5275,N_5878);
and U6396 (N_6396,N_5550,N_5743);
nor U6397 (N_6397,N_5467,N_5648);
xnor U6398 (N_6398,N_5339,N_5671);
and U6399 (N_6399,N_5307,N_5642);
xor U6400 (N_6400,N_5687,N_5267);
and U6401 (N_6401,N_5907,N_5708);
nor U6402 (N_6402,N_5488,N_5877);
and U6403 (N_6403,N_5783,N_5432);
or U6404 (N_6404,N_5954,N_5553);
nand U6405 (N_6405,N_5376,N_5806);
or U6406 (N_6406,N_5507,N_5329);
nand U6407 (N_6407,N_5635,N_5611);
nand U6408 (N_6408,N_5995,N_5663);
nand U6409 (N_6409,N_5452,N_5284);
nand U6410 (N_6410,N_5489,N_5605);
nand U6411 (N_6411,N_5673,N_5768);
xnor U6412 (N_6412,N_5441,N_5693);
and U6413 (N_6413,N_5814,N_5691);
nor U6414 (N_6414,N_5752,N_5366);
and U6415 (N_6415,N_5558,N_5523);
nand U6416 (N_6416,N_5361,N_5461);
or U6417 (N_6417,N_5840,N_5323);
and U6418 (N_6418,N_5818,N_5532);
and U6419 (N_6419,N_5766,N_5849);
or U6420 (N_6420,N_5413,N_5272);
nand U6421 (N_6421,N_5611,N_5782);
or U6422 (N_6422,N_5775,N_5733);
or U6423 (N_6423,N_5946,N_5290);
and U6424 (N_6424,N_5649,N_5925);
or U6425 (N_6425,N_5314,N_5667);
and U6426 (N_6426,N_5783,N_5758);
or U6427 (N_6427,N_5853,N_5498);
and U6428 (N_6428,N_5569,N_5381);
nor U6429 (N_6429,N_5587,N_5774);
xor U6430 (N_6430,N_5440,N_5672);
or U6431 (N_6431,N_5497,N_5653);
xor U6432 (N_6432,N_5736,N_5982);
nand U6433 (N_6433,N_5490,N_5911);
nor U6434 (N_6434,N_5665,N_5299);
nor U6435 (N_6435,N_5866,N_5781);
or U6436 (N_6436,N_5688,N_5530);
nand U6437 (N_6437,N_5672,N_5847);
nand U6438 (N_6438,N_5836,N_5678);
or U6439 (N_6439,N_5340,N_5526);
nand U6440 (N_6440,N_5512,N_5793);
nor U6441 (N_6441,N_5292,N_5774);
xor U6442 (N_6442,N_5742,N_5558);
or U6443 (N_6443,N_5316,N_5489);
or U6444 (N_6444,N_5333,N_5319);
or U6445 (N_6445,N_5859,N_5900);
nand U6446 (N_6446,N_5375,N_5653);
nor U6447 (N_6447,N_5864,N_5806);
nand U6448 (N_6448,N_5884,N_5706);
xor U6449 (N_6449,N_5420,N_5914);
xnor U6450 (N_6450,N_5671,N_5298);
xnor U6451 (N_6451,N_5787,N_5824);
xnor U6452 (N_6452,N_5286,N_5546);
and U6453 (N_6453,N_5970,N_5540);
xnor U6454 (N_6454,N_5537,N_5374);
nor U6455 (N_6455,N_5740,N_5647);
xor U6456 (N_6456,N_5712,N_5547);
and U6457 (N_6457,N_5492,N_5599);
or U6458 (N_6458,N_5460,N_5910);
nand U6459 (N_6459,N_5509,N_5879);
and U6460 (N_6460,N_5919,N_5536);
nor U6461 (N_6461,N_5702,N_5624);
xor U6462 (N_6462,N_5663,N_5972);
xnor U6463 (N_6463,N_5717,N_5930);
or U6464 (N_6464,N_5314,N_5473);
or U6465 (N_6465,N_5847,N_5923);
or U6466 (N_6466,N_5528,N_5742);
nor U6467 (N_6467,N_5389,N_5256);
nand U6468 (N_6468,N_5450,N_5701);
nand U6469 (N_6469,N_5711,N_5946);
xnor U6470 (N_6470,N_5309,N_5926);
and U6471 (N_6471,N_5524,N_5300);
and U6472 (N_6472,N_5571,N_5963);
nand U6473 (N_6473,N_5593,N_5282);
or U6474 (N_6474,N_5676,N_5669);
xor U6475 (N_6475,N_5626,N_5891);
nand U6476 (N_6476,N_5829,N_5505);
nor U6477 (N_6477,N_5500,N_5750);
xor U6478 (N_6478,N_5324,N_5934);
nand U6479 (N_6479,N_5559,N_5810);
nand U6480 (N_6480,N_5747,N_5991);
and U6481 (N_6481,N_5533,N_5853);
or U6482 (N_6482,N_5856,N_5250);
or U6483 (N_6483,N_5746,N_5620);
nor U6484 (N_6484,N_5909,N_5620);
and U6485 (N_6485,N_5762,N_5616);
nand U6486 (N_6486,N_5468,N_5794);
and U6487 (N_6487,N_5893,N_5965);
nor U6488 (N_6488,N_5305,N_5783);
nand U6489 (N_6489,N_5881,N_5834);
or U6490 (N_6490,N_5363,N_5282);
nor U6491 (N_6491,N_5281,N_5336);
nand U6492 (N_6492,N_5858,N_5798);
xnor U6493 (N_6493,N_5887,N_5886);
nand U6494 (N_6494,N_5927,N_5575);
and U6495 (N_6495,N_5910,N_5827);
xor U6496 (N_6496,N_5679,N_5614);
xor U6497 (N_6497,N_5560,N_5668);
nand U6498 (N_6498,N_5276,N_5572);
and U6499 (N_6499,N_5885,N_5665);
nand U6500 (N_6500,N_5917,N_5974);
or U6501 (N_6501,N_5868,N_5451);
or U6502 (N_6502,N_5803,N_5732);
or U6503 (N_6503,N_5599,N_5473);
nand U6504 (N_6504,N_5899,N_5918);
and U6505 (N_6505,N_5325,N_5640);
or U6506 (N_6506,N_5420,N_5312);
and U6507 (N_6507,N_5470,N_5940);
and U6508 (N_6508,N_5491,N_5396);
or U6509 (N_6509,N_5529,N_5277);
and U6510 (N_6510,N_5909,N_5855);
nor U6511 (N_6511,N_5926,N_5693);
nand U6512 (N_6512,N_5632,N_5289);
or U6513 (N_6513,N_5752,N_5739);
or U6514 (N_6514,N_5442,N_5666);
and U6515 (N_6515,N_5336,N_5763);
and U6516 (N_6516,N_5447,N_5698);
xnor U6517 (N_6517,N_5882,N_5589);
xor U6518 (N_6518,N_5622,N_5605);
and U6519 (N_6519,N_5951,N_5953);
nor U6520 (N_6520,N_5978,N_5610);
and U6521 (N_6521,N_5830,N_5356);
nor U6522 (N_6522,N_5668,N_5683);
or U6523 (N_6523,N_5769,N_5714);
or U6524 (N_6524,N_5570,N_5349);
and U6525 (N_6525,N_5790,N_5574);
nor U6526 (N_6526,N_5268,N_5960);
nor U6527 (N_6527,N_5772,N_5874);
and U6528 (N_6528,N_5949,N_5927);
or U6529 (N_6529,N_5301,N_5615);
nor U6530 (N_6530,N_5841,N_5972);
xnor U6531 (N_6531,N_5690,N_5328);
nand U6532 (N_6532,N_5368,N_5978);
nor U6533 (N_6533,N_5713,N_5805);
and U6534 (N_6534,N_5589,N_5264);
or U6535 (N_6535,N_5400,N_5627);
nor U6536 (N_6536,N_5491,N_5709);
or U6537 (N_6537,N_5273,N_5940);
nand U6538 (N_6538,N_5606,N_5342);
xnor U6539 (N_6539,N_5459,N_5964);
nand U6540 (N_6540,N_5562,N_5524);
xor U6541 (N_6541,N_5964,N_5265);
nor U6542 (N_6542,N_5793,N_5659);
nor U6543 (N_6543,N_5313,N_5842);
nor U6544 (N_6544,N_5948,N_5694);
nand U6545 (N_6545,N_5323,N_5938);
xor U6546 (N_6546,N_5418,N_5432);
or U6547 (N_6547,N_5416,N_5260);
and U6548 (N_6548,N_5327,N_5920);
or U6549 (N_6549,N_5839,N_5757);
xor U6550 (N_6550,N_5499,N_5712);
nand U6551 (N_6551,N_5400,N_5961);
and U6552 (N_6552,N_5345,N_5854);
or U6553 (N_6553,N_5999,N_5902);
nor U6554 (N_6554,N_5678,N_5294);
or U6555 (N_6555,N_5443,N_5638);
nor U6556 (N_6556,N_5943,N_5314);
or U6557 (N_6557,N_5990,N_5266);
nand U6558 (N_6558,N_5430,N_5494);
and U6559 (N_6559,N_5406,N_5385);
or U6560 (N_6560,N_5881,N_5919);
nand U6561 (N_6561,N_5781,N_5560);
or U6562 (N_6562,N_5860,N_5662);
nand U6563 (N_6563,N_5399,N_5964);
nand U6564 (N_6564,N_5262,N_5678);
or U6565 (N_6565,N_5640,N_5615);
nand U6566 (N_6566,N_5661,N_5874);
xor U6567 (N_6567,N_5736,N_5309);
nand U6568 (N_6568,N_5474,N_5804);
nor U6569 (N_6569,N_5334,N_5680);
and U6570 (N_6570,N_5475,N_5976);
xor U6571 (N_6571,N_5743,N_5336);
nand U6572 (N_6572,N_5943,N_5687);
nor U6573 (N_6573,N_5546,N_5337);
nor U6574 (N_6574,N_5847,N_5925);
or U6575 (N_6575,N_5810,N_5528);
or U6576 (N_6576,N_5353,N_5448);
or U6577 (N_6577,N_5360,N_5877);
and U6578 (N_6578,N_5636,N_5500);
and U6579 (N_6579,N_5347,N_5999);
or U6580 (N_6580,N_5789,N_5475);
nand U6581 (N_6581,N_5896,N_5385);
nand U6582 (N_6582,N_5265,N_5724);
and U6583 (N_6583,N_5480,N_5406);
and U6584 (N_6584,N_5273,N_5777);
and U6585 (N_6585,N_5373,N_5678);
nand U6586 (N_6586,N_5856,N_5620);
nor U6587 (N_6587,N_5326,N_5817);
nand U6588 (N_6588,N_5828,N_5656);
nor U6589 (N_6589,N_5432,N_5784);
and U6590 (N_6590,N_5373,N_5575);
nand U6591 (N_6591,N_5731,N_5523);
nor U6592 (N_6592,N_5583,N_5348);
nor U6593 (N_6593,N_5810,N_5530);
nor U6594 (N_6594,N_5289,N_5830);
nor U6595 (N_6595,N_5496,N_5282);
and U6596 (N_6596,N_5775,N_5950);
nor U6597 (N_6597,N_5443,N_5690);
and U6598 (N_6598,N_5542,N_5828);
nor U6599 (N_6599,N_5709,N_5563);
and U6600 (N_6600,N_5263,N_5634);
nor U6601 (N_6601,N_5710,N_5985);
nor U6602 (N_6602,N_5320,N_5586);
nand U6603 (N_6603,N_5674,N_5278);
or U6604 (N_6604,N_5801,N_5604);
xor U6605 (N_6605,N_5548,N_5278);
and U6606 (N_6606,N_5908,N_5648);
or U6607 (N_6607,N_5299,N_5292);
nor U6608 (N_6608,N_5621,N_5801);
nand U6609 (N_6609,N_5767,N_5751);
nor U6610 (N_6610,N_5707,N_5598);
or U6611 (N_6611,N_5783,N_5807);
nand U6612 (N_6612,N_5368,N_5659);
nor U6613 (N_6613,N_5486,N_5494);
or U6614 (N_6614,N_5514,N_5591);
and U6615 (N_6615,N_5927,N_5914);
or U6616 (N_6616,N_5659,N_5868);
and U6617 (N_6617,N_5746,N_5554);
nor U6618 (N_6618,N_5789,N_5911);
and U6619 (N_6619,N_5384,N_5996);
xor U6620 (N_6620,N_5725,N_5517);
or U6621 (N_6621,N_5681,N_5494);
nor U6622 (N_6622,N_5469,N_5719);
and U6623 (N_6623,N_5547,N_5339);
nand U6624 (N_6624,N_5995,N_5554);
nor U6625 (N_6625,N_5720,N_5758);
nor U6626 (N_6626,N_5791,N_5897);
nor U6627 (N_6627,N_5859,N_5926);
or U6628 (N_6628,N_5379,N_5700);
nor U6629 (N_6629,N_5905,N_5535);
and U6630 (N_6630,N_5264,N_5560);
or U6631 (N_6631,N_5464,N_5365);
nand U6632 (N_6632,N_5597,N_5342);
nand U6633 (N_6633,N_5806,N_5888);
nand U6634 (N_6634,N_5349,N_5897);
or U6635 (N_6635,N_5775,N_5964);
nand U6636 (N_6636,N_5805,N_5614);
nand U6637 (N_6637,N_5304,N_5848);
or U6638 (N_6638,N_5604,N_5342);
and U6639 (N_6639,N_5974,N_5925);
nor U6640 (N_6640,N_5967,N_5907);
nor U6641 (N_6641,N_5516,N_5644);
nor U6642 (N_6642,N_5377,N_5505);
and U6643 (N_6643,N_5336,N_5289);
nor U6644 (N_6644,N_5901,N_5441);
and U6645 (N_6645,N_5878,N_5955);
nor U6646 (N_6646,N_5277,N_5478);
or U6647 (N_6647,N_5538,N_5470);
nor U6648 (N_6648,N_5590,N_5613);
nand U6649 (N_6649,N_5762,N_5837);
nand U6650 (N_6650,N_5342,N_5301);
and U6651 (N_6651,N_5831,N_5384);
and U6652 (N_6652,N_5255,N_5632);
nand U6653 (N_6653,N_5523,N_5687);
nor U6654 (N_6654,N_5263,N_5483);
or U6655 (N_6655,N_5494,N_5650);
nand U6656 (N_6656,N_5939,N_5802);
and U6657 (N_6657,N_5477,N_5263);
nor U6658 (N_6658,N_5676,N_5570);
nand U6659 (N_6659,N_5290,N_5255);
and U6660 (N_6660,N_5505,N_5627);
xnor U6661 (N_6661,N_5966,N_5367);
nor U6662 (N_6662,N_5811,N_5939);
nor U6663 (N_6663,N_5878,N_5529);
xor U6664 (N_6664,N_5771,N_5288);
nand U6665 (N_6665,N_5746,N_5305);
and U6666 (N_6666,N_5533,N_5384);
or U6667 (N_6667,N_5950,N_5595);
and U6668 (N_6668,N_5880,N_5628);
nand U6669 (N_6669,N_5419,N_5309);
nand U6670 (N_6670,N_5828,N_5833);
or U6671 (N_6671,N_5515,N_5822);
nand U6672 (N_6672,N_5442,N_5622);
and U6673 (N_6673,N_5821,N_5323);
nor U6674 (N_6674,N_5473,N_5423);
nor U6675 (N_6675,N_5934,N_5840);
and U6676 (N_6676,N_5963,N_5445);
nand U6677 (N_6677,N_5963,N_5669);
or U6678 (N_6678,N_5372,N_5281);
and U6679 (N_6679,N_5573,N_5518);
nand U6680 (N_6680,N_5831,N_5366);
nand U6681 (N_6681,N_5452,N_5629);
or U6682 (N_6682,N_5679,N_5300);
nor U6683 (N_6683,N_5928,N_5328);
or U6684 (N_6684,N_5931,N_5826);
nor U6685 (N_6685,N_5732,N_5321);
or U6686 (N_6686,N_5836,N_5266);
and U6687 (N_6687,N_5263,N_5636);
and U6688 (N_6688,N_5485,N_5665);
or U6689 (N_6689,N_5771,N_5264);
nor U6690 (N_6690,N_5908,N_5820);
nand U6691 (N_6691,N_5864,N_5855);
or U6692 (N_6692,N_5496,N_5254);
nand U6693 (N_6693,N_5816,N_5887);
xor U6694 (N_6694,N_5597,N_5784);
nor U6695 (N_6695,N_5973,N_5541);
and U6696 (N_6696,N_5988,N_5766);
nand U6697 (N_6697,N_5485,N_5611);
nand U6698 (N_6698,N_5519,N_5633);
or U6699 (N_6699,N_5548,N_5946);
nand U6700 (N_6700,N_5251,N_5388);
and U6701 (N_6701,N_5457,N_5739);
nor U6702 (N_6702,N_5267,N_5719);
and U6703 (N_6703,N_5703,N_5509);
or U6704 (N_6704,N_5531,N_5741);
xnor U6705 (N_6705,N_5296,N_5568);
and U6706 (N_6706,N_5742,N_5265);
nor U6707 (N_6707,N_5257,N_5263);
nor U6708 (N_6708,N_5283,N_5376);
nand U6709 (N_6709,N_5520,N_5897);
and U6710 (N_6710,N_5437,N_5472);
and U6711 (N_6711,N_5871,N_5396);
nand U6712 (N_6712,N_5645,N_5721);
or U6713 (N_6713,N_5841,N_5620);
nand U6714 (N_6714,N_5451,N_5727);
nor U6715 (N_6715,N_5619,N_5376);
and U6716 (N_6716,N_5831,N_5810);
or U6717 (N_6717,N_5567,N_5445);
or U6718 (N_6718,N_5298,N_5394);
or U6719 (N_6719,N_5979,N_5725);
nor U6720 (N_6720,N_5696,N_5270);
or U6721 (N_6721,N_5756,N_5684);
nor U6722 (N_6722,N_5826,N_5883);
nor U6723 (N_6723,N_5589,N_5586);
nor U6724 (N_6724,N_5584,N_5953);
or U6725 (N_6725,N_5645,N_5425);
nand U6726 (N_6726,N_5757,N_5322);
nor U6727 (N_6727,N_5302,N_5556);
nor U6728 (N_6728,N_5566,N_5646);
nand U6729 (N_6729,N_5391,N_5287);
or U6730 (N_6730,N_5968,N_5656);
nand U6731 (N_6731,N_5868,N_5825);
or U6732 (N_6732,N_5304,N_5805);
nand U6733 (N_6733,N_5327,N_5395);
nor U6734 (N_6734,N_5893,N_5867);
and U6735 (N_6735,N_5567,N_5421);
and U6736 (N_6736,N_5856,N_5966);
xnor U6737 (N_6737,N_5749,N_5857);
nand U6738 (N_6738,N_5476,N_5885);
and U6739 (N_6739,N_5488,N_5379);
and U6740 (N_6740,N_5655,N_5971);
nand U6741 (N_6741,N_5659,N_5516);
nor U6742 (N_6742,N_5656,N_5473);
nand U6743 (N_6743,N_5515,N_5880);
nand U6744 (N_6744,N_5925,N_5645);
nor U6745 (N_6745,N_5603,N_5371);
nand U6746 (N_6746,N_5357,N_5586);
nor U6747 (N_6747,N_5765,N_5732);
nor U6748 (N_6748,N_5968,N_5702);
nand U6749 (N_6749,N_5260,N_5836);
and U6750 (N_6750,N_6696,N_6204);
or U6751 (N_6751,N_6176,N_6488);
or U6752 (N_6752,N_6654,N_6317);
nand U6753 (N_6753,N_6743,N_6609);
nor U6754 (N_6754,N_6699,N_6022);
and U6755 (N_6755,N_6080,N_6132);
or U6756 (N_6756,N_6619,N_6029);
nand U6757 (N_6757,N_6073,N_6649);
xor U6758 (N_6758,N_6718,N_6498);
xnor U6759 (N_6759,N_6087,N_6578);
or U6760 (N_6760,N_6378,N_6044);
xor U6761 (N_6761,N_6479,N_6269);
nor U6762 (N_6762,N_6615,N_6723);
or U6763 (N_6763,N_6362,N_6257);
nor U6764 (N_6764,N_6556,N_6147);
nor U6765 (N_6765,N_6031,N_6559);
or U6766 (N_6766,N_6746,N_6105);
nor U6767 (N_6767,N_6681,N_6507);
and U6768 (N_6768,N_6316,N_6118);
or U6769 (N_6769,N_6700,N_6625);
nand U6770 (N_6770,N_6156,N_6177);
and U6771 (N_6771,N_6116,N_6344);
and U6772 (N_6772,N_6091,N_6076);
xor U6773 (N_6773,N_6096,N_6385);
and U6774 (N_6774,N_6013,N_6023);
and U6775 (N_6775,N_6030,N_6747);
nor U6776 (N_6776,N_6386,N_6701);
or U6777 (N_6777,N_6237,N_6028);
xnor U6778 (N_6778,N_6259,N_6202);
and U6779 (N_6779,N_6138,N_6705);
or U6780 (N_6780,N_6651,N_6060);
and U6781 (N_6781,N_6196,N_6579);
or U6782 (N_6782,N_6337,N_6695);
nor U6783 (N_6783,N_6387,N_6140);
and U6784 (N_6784,N_6338,N_6302);
nor U6785 (N_6785,N_6124,N_6424);
or U6786 (N_6786,N_6347,N_6444);
nor U6787 (N_6787,N_6465,N_6329);
xnor U6788 (N_6788,N_6602,N_6068);
or U6789 (N_6789,N_6352,N_6224);
nand U6790 (N_6790,N_6744,N_6351);
nand U6791 (N_6791,N_6405,N_6320);
and U6792 (N_6792,N_6219,N_6055);
xnor U6793 (N_6793,N_6595,N_6078);
xor U6794 (N_6794,N_6016,N_6130);
or U6795 (N_6795,N_6340,N_6165);
nor U6796 (N_6796,N_6518,N_6453);
nor U6797 (N_6797,N_6141,N_6353);
or U6798 (N_6798,N_6460,N_6228);
xnor U6799 (N_6799,N_6180,N_6006);
and U6800 (N_6800,N_6153,N_6547);
and U6801 (N_6801,N_6562,N_6135);
nand U6802 (N_6802,N_6402,N_6238);
and U6803 (N_6803,N_6631,N_6635);
nand U6804 (N_6804,N_6077,N_6706);
and U6805 (N_6805,N_6443,N_6371);
nand U6806 (N_6806,N_6647,N_6439);
nand U6807 (N_6807,N_6208,N_6494);
nor U6808 (N_6808,N_6611,N_6169);
nor U6809 (N_6809,N_6531,N_6232);
xnor U6810 (N_6810,N_6532,N_6104);
nor U6811 (N_6811,N_6117,N_6571);
nand U6812 (N_6812,N_6382,N_6653);
and U6813 (N_6813,N_6283,N_6624);
nand U6814 (N_6814,N_6564,N_6027);
or U6815 (N_6815,N_6021,N_6423);
and U6816 (N_6816,N_6291,N_6497);
or U6817 (N_6817,N_6721,N_6473);
or U6818 (N_6818,N_6039,N_6324);
nor U6819 (N_6819,N_6704,N_6644);
or U6820 (N_6820,N_6363,N_6582);
nand U6821 (N_6821,N_6430,N_6729);
or U6822 (N_6822,N_6639,N_6737);
nor U6823 (N_6823,N_6209,N_6081);
or U6824 (N_6824,N_6446,N_6476);
nand U6825 (N_6825,N_6420,N_6300);
or U6826 (N_6826,N_6409,N_6724);
nor U6827 (N_6827,N_6484,N_6728);
or U6828 (N_6828,N_6590,N_6384);
nor U6829 (N_6829,N_6419,N_6145);
and U6830 (N_6830,N_6440,N_6436);
or U6831 (N_6831,N_6563,N_6711);
nand U6832 (N_6832,N_6535,N_6416);
or U6833 (N_6833,N_6134,N_6489);
nor U6834 (N_6834,N_6233,N_6033);
xnor U6835 (N_6835,N_6062,N_6061);
and U6836 (N_6836,N_6358,N_6434);
xnor U6837 (N_6837,N_6574,N_6053);
and U6838 (N_6838,N_6152,N_6458);
nor U6839 (N_6839,N_6015,N_6425);
nor U6840 (N_6840,N_6139,N_6464);
xnor U6841 (N_6841,N_6236,N_6048);
nor U6842 (N_6842,N_6702,N_6207);
and U6843 (N_6843,N_6738,N_6401);
nand U6844 (N_6844,N_6586,N_6070);
or U6845 (N_6845,N_6311,N_6457);
or U6846 (N_6846,N_6618,N_6066);
or U6847 (N_6847,N_6171,N_6067);
nand U6848 (N_6848,N_6332,N_6273);
or U6849 (N_6849,N_6075,N_6100);
and U6850 (N_6850,N_6486,N_6530);
nand U6851 (N_6851,N_6242,N_6495);
nand U6852 (N_6852,N_6720,N_6265);
and U6853 (N_6853,N_6054,N_6356);
nand U6854 (N_6854,N_6266,N_6674);
or U6855 (N_6855,N_6297,N_6534);
or U6856 (N_6856,N_6375,N_6550);
and U6857 (N_6857,N_6575,N_6648);
nand U6858 (N_6858,N_6391,N_6435);
and U6859 (N_6859,N_6018,N_6043);
nor U6860 (N_6860,N_6278,N_6005);
nor U6861 (N_6861,N_6240,N_6111);
and U6862 (N_6862,N_6042,N_6052);
xor U6863 (N_6863,N_6071,N_6703);
xnor U6864 (N_6864,N_6113,N_6357);
or U6865 (N_6865,N_6692,N_6355);
nor U6866 (N_6866,N_6000,N_6241);
xor U6867 (N_6867,N_6119,N_6331);
nand U6868 (N_6868,N_6270,N_6577);
or U6869 (N_6869,N_6628,N_6088);
or U6870 (N_6870,N_6736,N_6157);
or U6871 (N_6871,N_6292,N_6432);
nor U6872 (N_6872,N_6576,N_6212);
or U6873 (N_6873,N_6438,N_6643);
or U6874 (N_6874,N_6741,N_6256);
or U6875 (N_6875,N_6682,N_6710);
or U6876 (N_6876,N_6588,N_6093);
xnor U6877 (N_6877,N_6129,N_6244);
nand U6878 (N_6878,N_6698,N_6040);
or U6879 (N_6879,N_6306,N_6065);
xor U6880 (N_6880,N_6086,N_6400);
and U6881 (N_6881,N_6468,N_6646);
and U6882 (N_6882,N_6677,N_6678);
nor U6883 (N_6883,N_6211,N_6634);
nand U6884 (N_6884,N_6217,N_6707);
nor U6885 (N_6885,N_6336,N_6395);
or U6886 (N_6886,N_6330,N_6557);
nor U6887 (N_6887,N_6731,N_6187);
nor U6888 (N_6888,N_6543,N_6657);
and U6889 (N_6889,N_6520,N_6200);
xor U6890 (N_6890,N_6669,N_6001);
nand U6891 (N_6891,N_6448,N_6636);
xnor U6892 (N_6892,N_6660,N_6144);
nor U6893 (N_6893,N_6414,N_6299);
nor U6894 (N_6894,N_6218,N_6629);
and U6895 (N_6895,N_6020,N_6342);
xor U6896 (N_6896,N_6449,N_6389);
or U6897 (N_6897,N_6663,N_6626);
nor U6898 (N_6898,N_6418,N_6148);
nand U6899 (N_6899,N_6540,N_6083);
and U6900 (N_6900,N_6687,N_6641);
xnor U6901 (N_6901,N_6255,N_6315);
or U6902 (N_6902,N_6490,N_6733);
nor U6903 (N_6903,N_6110,N_6505);
nand U6904 (N_6904,N_6133,N_6549);
nor U6905 (N_6905,N_6509,N_6412);
or U6906 (N_6906,N_6693,N_6496);
xnor U6907 (N_6907,N_6348,N_6570);
nand U6908 (N_6908,N_6295,N_6034);
and U6909 (N_6909,N_6098,N_6094);
xnor U6910 (N_6910,N_6474,N_6084);
nand U6911 (N_6911,N_6456,N_6193);
xnor U6912 (N_6912,N_6676,N_6154);
xor U6913 (N_6913,N_6126,N_6665);
nor U6914 (N_6914,N_6056,N_6229);
nor U6915 (N_6915,N_6099,N_6179);
nand U6916 (N_6916,N_6343,N_6069);
nor U6917 (N_6917,N_6442,N_6003);
xor U6918 (N_6918,N_6210,N_6587);
nand U6919 (N_6919,N_6554,N_6271);
and U6920 (N_6920,N_6514,N_6106);
or U6921 (N_6921,N_6573,N_6136);
or U6922 (N_6922,N_6280,N_6074);
nor U6923 (N_6923,N_6581,N_6666);
nor U6924 (N_6924,N_6607,N_6417);
nor U6925 (N_6925,N_6592,N_6230);
or U6926 (N_6926,N_6234,N_6477);
nor U6927 (N_6927,N_6115,N_6227);
nand U6928 (N_6928,N_6719,N_6725);
or U6929 (N_6929,N_6471,N_6112);
or U6930 (N_6930,N_6321,N_6679);
nor U6931 (N_6931,N_6103,N_6181);
xnor U6932 (N_6932,N_6404,N_6325);
nor U6933 (N_6933,N_6500,N_6092);
nor U6934 (N_6934,N_6307,N_6263);
nor U6935 (N_6935,N_6726,N_6305);
or U6936 (N_6936,N_6441,N_6183);
nand U6937 (N_6937,N_6732,N_6735);
nor U6938 (N_6938,N_6328,N_6604);
xnor U6939 (N_6939,N_6254,N_6533);
nand U6940 (N_6940,N_6668,N_6007);
nand U6941 (N_6941,N_6287,N_6369);
and U6942 (N_6942,N_6716,N_6637);
nand U6943 (N_6943,N_6184,N_6608);
nor U6944 (N_6944,N_6014,N_6407);
or U6945 (N_6945,N_6308,N_6279);
nor U6946 (N_6946,N_6481,N_6394);
or U6947 (N_6947,N_6516,N_6174);
and U6948 (N_6948,N_6286,N_6312);
nand U6949 (N_6949,N_6206,N_6047);
and U6950 (N_6950,N_6569,N_6482);
nor U6951 (N_6951,N_6551,N_6715);
and U6952 (N_6952,N_6216,N_6341);
and U6953 (N_6953,N_6131,N_6742);
nand U6954 (N_6954,N_6526,N_6319);
or U6955 (N_6955,N_6194,N_6722);
xor U6956 (N_6956,N_6215,N_6222);
or U6957 (N_6957,N_6235,N_6463);
nor U6958 (N_6958,N_6428,N_6597);
or U6959 (N_6959,N_6655,N_6612);
xor U6960 (N_6960,N_6289,N_6593);
and U6961 (N_6961,N_6008,N_6504);
or U6962 (N_6962,N_6192,N_6349);
or U6963 (N_6963,N_6584,N_6510);
xor U6964 (N_6964,N_6290,N_6598);
and U6965 (N_6965,N_6301,N_6617);
nor U6966 (N_6966,N_6127,N_6381);
and U6967 (N_6967,N_6431,N_6149);
nor U6968 (N_6968,N_6709,N_6050);
nor U6969 (N_6969,N_6261,N_6525);
nand U6970 (N_6970,N_6642,N_6383);
xor U6971 (N_6971,N_6010,N_6645);
nand U6972 (N_6972,N_6396,N_6580);
nor U6973 (N_6973,N_6281,N_6390);
nor U6974 (N_6974,N_6189,N_6346);
or U6975 (N_6975,N_6026,N_6175);
nor U6976 (N_6976,N_6045,N_6262);
nand U6977 (N_6977,N_6231,N_6499);
or U6978 (N_6978,N_6025,N_6452);
nand U6979 (N_6979,N_6466,N_6168);
and U6980 (N_6980,N_6178,N_6675);
and U6981 (N_6981,N_6258,N_6661);
and U6982 (N_6982,N_6650,N_6101);
or U6983 (N_6983,N_6277,N_6367);
or U6984 (N_6984,N_6223,N_6555);
nor U6985 (N_6985,N_6561,N_6246);
xor U6986 (N_6986,N_6122,N_6513);
nor U6987 (N_6987,N_6195,N_6051);
nor U6988 (N_6988,N_6511,N_6372);
nor U6989 (N_6989,N_6379,N_6596);
nand U6990 (N_6990,N_6536,N_6251);
xnor U6991 (N_6991,N_6063,N_6671);
or U6992 (N_6992,N_6248,N_6684);
and U6993 (N_6993,N_6475,N_6734);
nand U6994 (N_6994,N_6487,N_6522);
nand U6995 (N_6995,N_6548,N_6545);
nor U6996 (N_6996,N_6036,N_6089);
nor U6997 (N_6997,N_6267,N_6158);
nor U6998 (N_6998,N_6366,N_6182);
nand U6999 (N_6999,N_6002,N_6708);
nand U7000 (N_7000,N_6714,N_6406);
nand U7001 (N_7001,N_6673,N_6740);
nand U7002 (N_7002,N_6125,N_6032);
nor U7003 (N_7003,N_6461,N_6606);
or U7004 (N_7004,N_6350,N_6670);
xnor U7005 (N_7005,N_6640,N_6470);
xor U7006 (N_7006,N_6667,N_6354);
nor U7007 (N_7007,N_6749,N_6472);
nand U7008 (N_7008,N_6480,N_6009);
xnor U7009 (N_7009,N_6155,N_6339);
or U7010 (N_7010,N_6199,N_6250);
and U7011 (N_7011,N_6151,N_6072);
nor U7012 (N_7012,N_6326,N_6664);
or U7013 (N_7013,N_6167,N_6298);
nor U7014 (N_7014,N_6478,N_6380);
nor U7015 (N_7015,N_6415,N_6304);
or U7016 (N_7016,N_6620,N_6519);
nor U7017 (N_7017,N_6359,N_6621);
nand U7018 (N_7018,N_6688,N_6161);
and U7019 (N_7019,N_6318,N_6717);
nand U7020 (N_7020,N_6537,N_6186);
xor U7021 (N_7021,N_6501,N_6544);
or U7022 (N_7022,N_6403,N_6085);
or U7023 (N_7023,N_6506,N_6659);
nor U7024 (N_7024,N_6690,N_6686);
nor U7025 (N_7025,N_6373,N_6429);
and U7026 (N_7026,N_6613,N_6309);
and U7027 (N_7027,N_6024,N_6046);
nand U7028 (N_7028,N_6313,N_6393);
nand U7029 (N_7029,N_6517,N_6388);
nand U7030 (N_7030,N_6142,N_6296);
or U7031 (N_7031,N_6213,N_6689);
nor U7032 (N_7032,N_6082,N_6558);
nor U7033 (N_7033,N_6483,N_6102);
nor U7034 (N_7034,N_6727,N_6163);
nor U7035 (N_7035,N_6527,N_6600);
xor U7036 (N_7036,N_6652,N_6333);
or U7037 (N_7037,N_6568,N_6146);
nand U7038 (N_7038,N_6365,N_6594);
nor U7039 (N_7039,N_6426,N_6284);
or U7040 (N_7040,N_6361,N_6528);
nand U7041 (N_7041,N_6662,N_6398);
and U7042 (N_7042,N_6164,N_6553);
xor U7043 (N_7043,N_6630,N_6748);
and U7044 (N_7044,N_6090,N_6260);
nor U7045 (N_7045,N_6335,N_6421);
or U7046 (N_7046,N_6252,N_6491);
and U7047 (N_7047,N_6411,N_6264);
nor U7048 (N_7048,N_6567,N_6035);
and U7049 (N_7049,N_6049,N_6459);
or U7050 (N_7050,N_6327,N_6633);
nand U7051 (N_7051,N_6493,N_6739);
and U7052 (N_7052,N_6197,N_6012);
and U7053 (N_7053,N_6603,N_6399);
nand U7054 (N_7054,N_6114,N_6447);
xor U7055 (N_7055,N_6672,N_6585);
xor U7056 (N_7056,N_6683,N_6159);
nor U7057 (N_7057,N_6364,N_6243);
nor U7058 (N_7058,N_6485,N_6143);
and U7059 (N_7059,N_6057,N_6450);
nor U7060 (N_7060,N_6019,N_6360);
nand U7061 (N_7061,N_6462,N_6422);
nor U7062 (N_7062,N_6097,N_6392);
xnor U7063 (N_7063,N_6685,N_6410);
nor U7064 (N_7064,N_6694,N_6451);
and U7065 (N_7065,N_6303,N_6376);
xor U7066 (N_7066,N_6272,N_6691);
nor U7067 (N_7067,N_6214,N_6601);
xor U7068 (N_7068,N_6377,N_6120);
or U7069 (N_7069,N_6268,N_6658);
nand U7070 (N_7070,N_6427,N_6245);
nor U7071 (N_7071,N_6546,N_6017);
nor U7072 (N_7072,N_6221,N_6064);
xnor U7073 (N_7073,N_6572,N_6274);
nor U7074 (N_7074,N_6538,N_6565);
and U7075 (N_7075,N_6566,N_6521);
nor U7076 (N_7076,N_6492,N_6627);
or U7077 (N_7077,N_6160,N_6170);
nor U7078 (N_7078,N_6542,N_6004);
nand U7079 (N_7079,N_6275,N_6334);
and U7080 (N_7080,N_6011,N_6437);
nor U7081 (N_7081,N_6503,N_6322);
nand U7082 (N_7082,N_6041,N_6638);
nor U7083 (N_7083,N_6623,N_6108);
and U7084 (N_7084,N_6191,N_6310);
and U7085 (N_7085,N_6502,N_6166);
nand U7086 (N_7086,N_6512,N_6345);
and U7087 (N_7087,N_6632,N_6445);
nand U7088 (N_7088,N_6433,N_6467);
nand U7089 (N_7089,N_6374,N_6107);
nand U7090 (N_7090,N_6589,N_6368);
nor U7091 (N_7091,N_6173,N_6198);
nand U7092 (N_7092,N_6454,N_6455);
and U7093 (N_7093,N_6109,N_6058);
or U7094 (N_7094,N_6680,N_6137);
nand U7095 (N_7095,N_6128,N_6713);
nand U7096 (N_7096,N_6285,N_6059);
and U7097 (N_7097,N_6282,N_6203);
xnor U7098 (N_7098,N_6121,N_6560);
or U7099 (N_7099,N_6123,N_6730);
nand U7100 (N_7100,N_6323,N_6247);
nand U7101 (N_7101,N_6591,N_6188);
nor U7102 (N_7102,N_6249,N_6293);
and U7103 (N_7103,N_6220,N_6185);
and U7104 (N_7104,N_6413,N_6190);
xor U7105 (N_7105,N_6038,N_6469);
or U7106 (N_7106,N_6539,N_6408);
or U7107 (N_7107,N_6079,N_6276);
nor U7108 (N_7108,N_6205,N_6239);
nor U7109 (N_7109,N_6599,N_6162);
or U7110 (N_7110,N_6605,N_6745);
and U7111 (N_7111,N_6370,N_6397);
nand U7112 (N_7112,N_6314,N_6225);
and U7113 (N_7113,N_6529,N_6288);
nor U7114 (N_7114,N_6583,N_6656);
nor U7115 (N_7115,N_6552,N_6294);
and U7116 (N_7116,N_6172,N_6037);
nand U7117 (N_7117,N_6697,N_6523);
nor U7118 (N_7118,N_6610,N_6541);
xnor U7119 (N_7119,N_6201,N_6508);
nor U7120 (N_7120,N_6515,N_6226);
or U7121 (N_7121,N_6524,N_6712);
nand U7122 (N_7122,N_6095,N_6616);
nand U7123 (N_7123,N_6622,N_6253);
xor U7124 (N_7124,N_6614,N_6150);
nor U7125 (N_7125,N_6378,N_6077);
nor U7126 (N_7126,N_6651,N_6741);
nor U7127 (N_7127,N_6169,N_6532);
nand U7128 (N_7128,N_6299,N_6136);
nand U7129 (N_7129,N_6546,N_6040);
and U7130 (N_7130,N_6433,N_6420);
and U7131 (N_7131,N_6680,N_6545);
nor U7132 (N_7132,N_6165,N_6637);
or U7133 (N_7133,N_6744,N_6452);
xor U7134 (N_7134,N_6484,N_6238);
nor U7135 (N_7135,N_6747,N_6417);
or U7136 (N_7136,N_6162,N_6237);
xor U7137 (N_7137,N_6010,N_6092);
xnor U7138 (N_7138,N_6394,N_6280);
xor U7139 (N_7139,N_6329,N_6223);
nand U7140 (N_7140,N_6709,N_6170);
and U7141 (N_7141,N_6110,N_6327);
nor U7142 (N_7142,N_6117,N_6365);
and U7143 (N_7143,N_6260,N_6421);
nor U7144 (N_7144,N_6121,N_6529);
and U7145 (N_7145,N_6221,N_6236);
nor U7146 (N_7146,N_6643,N_6029);
and U7147 (N_7147,N_6276,N_6733);
and U7148 (N_7148,N_6219,N_6462);
or U7149 (N_7149,N_6672,N_6324);
nand U7150 (N_7150,N_6112,N_6623);
nor U7151 (N_7151,N_6195,N_6065);
nand U7152 (N_7152,N_6275,N_6128);
nor U7153 (N_7153,N_6520,N_6204);
nand U7154 (N_7154,N_6465,N_6478);
and U7155 (N_7155,N_6080,N_6472);
nand U7156 (N_7156,N_6147,N_6149);
nor U7157 (N_7157,N_6285,N_6393);
or U7158 (N_7158,N_6226,N_6661);
nor U7159 (N_7159,N_6237,N_6000);
xor U7160 (N_7160,N_6231,N_6472);
and U7161 (N_7161,N_6324,N_6703);
nor U7162 (N_7162,N_6579,N_6672);
and U7163 (N_7163,N_6485,N_6036);
nand U7164 (N_7164,N_6403,N_6446);
or U7165 (N_7165,N_6561,N_6608);
nand U7166 (N_7166,N_6526,N_6551);
nor U7167 (N_7167,N_6546,N_6054);
nor U7168 (N_7168,N_6155,N_6268);
xor U7169 (N_7169,N_6490,N_6485);
nor U7170 (N_7170,N_6532,N_6146);
nor U7171 (N_7171,N_6104,N_6030);
and U7172 (N_7172,N_6719,N_6532);
nor U7173 (N_7173,N_6567,N_6405);
and U7174 (N_7174,N_6284,N_6418);
and U7175 (N_7175,N_6473,N_6325);
nand U7176 (N_7176,N_6173,N_6600);
and U7177 (N_7177,N_6245,N_6635);
and U7178 (N_7178,N_6038,N_6425);
nor U7179 (N_7179,N_6501,N_6257);
and U7180 (N_7180,N_6588,N_6087);
nand U7181 (N_7181,N_6239,N_6287);
nand U7182 (N_7182,N_6469,N_6084);
nand U7183 (N_7183,N_6462,N_6356);
nand U7184 (N_7184,N_6388,N_6532);
nor U7185 (N_7185,N_6601,N_6518);
nor U7186 (N_7186,N_6387,N_6673);
or U7187 (N_7187,N_6085,N_6223);
nor U7188 (N_7188,N_6019,N_6492);
nand U7189 (N_7189,N_6439,N_6245);
nor U7190 (N_7190,N_6134,N_6453);
nor U7191 (N_7191,N_6017,N_6708);
nand U7192 (N_7192,N_6744,N_6087);
nor U7193 (N_7193,N_6308,N_6398);
and U7194 (N_7194,N_6288,N_6387);
xor U7195 (N_7195,N_6234,N_6424);
nor U7196 (N_7196,N_6680,N_6460);
nand U7197 (N_7197,N_6264,N_6407);
nand U7198 (N_7198,N_6158,N_6065);
or U7199 (N_7199,N_6728,N_6378);
or U7200 (N_7200,N_6677,N_6540);
xnor U7201 (N_7201,N_6370,N_6180);
nand U7202 (N_7202,N_6487,N_6157);
nand U7203 (N_7203,N_6616,N_6580);
xnor U7204 (N_7204,N_6100,N_6634);
nand U7205 (N_7205,N_6236,N_6699);
nor U7206 (N_7206,N_6000,N_6230);
nand U7207 (N_7207,N_6693,N_6384);
and U7208 (N_7208,N_6647,N_6344);
or U7209 (N_7209,N_6450,N_6430);
nor U7210 (N_7210,N_6480,N_6402);
nand U7211 (N_7211,N_6707,N_6367);
xor U7212 (N_7212,N_6541,N_6383);
nor U7213 (N_7213,N_6244,N_6030);
and U7214 (N_7214,N_6010,N_6573);
and U7215 (N_7215,N_6032,N_6441);
nor U7216 (N_7216,N_6567,N_6056);
and U7217 (N_7217,N_6526,N_6313);
and U7218 (N_7218,N_6070,N_6509);
or U7219 (N_7219,N_6531,N_6435);
nand U7220 (N_7220,N_6619,N_6219);
or U7221 (N_7221,N_6435,N_6205);
nand U7222 (N_7222,N_6359,N_6625);
nand U7223 (N_7223,N_6413,N_6688);
or U7224 (N_7224,N_6120,N_6169);
nor U7225 (N_7225,N_6205,N_6121);
nor U7226 (N_7226,N_6387,N_6441);
or U7227 (N_7227,N_6027,N_6443);
nand U7228 (N_7228,N_6254,N_6282);
or U7229 (N_7229,N_6088,N_6273);
or U7230 (N_7230,N_6646,N_6210);
nand U7231 (N_7231,N_6332,N_6260);
nor U7232 (N_7232,N_6697,N_6190);
or U7233 (N_7233,N_6008,N_6434);
nand U7234 (N_7234,N_6098,N_6280);
nor U7235 (N_7235,N_6053,N_6671);
nand U7236 (N_7236,N_6677,N_6516);
nor U7237 (N_7237,N_6143,N_6356);
nand U7238 (N_7238,N_6545,N_6691);
or U7239 (N_7239,N_6506,N_6499);
xnor U7240 (N_7240,N_6173,N_6452);
and U7241 (N_7241,N_6418,N_6247);
nand U7242 (N_7242,N_6617,N_6411);
xor U7243 (N_7243,N_6436,N_6653);
nor U7244 (N_7244,N_6162,N_6077);
nor U7245 (N_7245,N_6411,N_6514);
or U7246 (N_7246,N_6745,N_6308);
nand U7247 (N_7247,N_6698,N_6673);
nor U7248 (N_7248,N_6021,N_6022);
nand U7249 (N_7249,N_6564,N_6329);
or U7250 (N_7250,N_6292,N_6348);
and U7251 (N_7251,N_6162,N_6559);
nor U7252 (N_7252,N_6505,N_6327);
nand U7253 (N_7253,N_6661,N_6579);
nor U7254 (N_7254,N_6162,N_6002);
nand U7255 (N_7255,N_6599,N_6607);
nor U7256 (N_7256,N_6364,N_6446);
nor U7257 (N_7257,N_6555,N_6510);
nor U7258 (N_7258,N_6099,N_6683);
or U7259 (N_7259,N_6244,N_6591);
or U7260 (N_7260,N_6473,N_6653);
nor U7261 (N_7261,N_6005,N_6506);
nand U7262 (N_7262,N_6593,N_6743);
or U7263 (N_7263,N_6492,N_6092);
nor U7264 (N_7264,N_6297,N_6613);
and U7265 (N_7265,N_6531,N_6551);
xnor U7266 (N_7266,N_6048,N_6117);
and U7267 (N_7267,N_6477,N_6420);
and U7268 (N_7268,N_6413,N_6392);
nand U7269 (N_7269,N_6199,N_6420);
and U7270 (N_7270,N_6196,N_6097);
nor U7271 (N_7271,N_6080,N_6447);
or U7272 (N_7272,N_6070,N_6331);
and U7273 (N_7273,N_6427,N_6441);
xnor U7274 (N_7274,N_6472,N_6001);
nand U7275 (N_7275,N_6356,N_6467);
and U7276 (N_7276,N_6337,N_6550);
nand U7277 (N_7277,N_6406,N_6634);
and U7278 (N_7278,N_6576,N_6152);
nand U7279 (N_7279,N_6280,N_6251);
nor U7280 (N_7280,N_6673,N_6736);
xnor U7281 (N_7281,N_6159,N_6312);
or U7282 (N_7282,N_6153,N_6585);
or U7283 (N_7283,N_6145,N_6453);
xor U7284 (N_7284,N_6625,N_6276);
and U7285 (N_7285,N_6056,N_6693);
nor U7286 (N_7286,N_6647,N_6434);
and U7287 (N_7287,N_6671,N_6349);
or U7288 (N_7288,N_6311,N_6626);
nand U7289 (N_7289,N_6142,N_6708);
nor U7290 (N_7290,N_6694,N_6329);
or U7291 (N_7291,N_6316,N_6222);
or U7292 (N_7292,N_6399,N_6217);
nand U7293 (N_7293,N_6451,N_6003);
nand U7294 (N_7294,N_6491,N_6371);
nand U7295 (N_7295,N_6160,N_6730);
nand U7296 (N_7296,N_6590,N_6166);
or U7297 (N_7297,N_6339,N_6597);
nor U7298 (N_7298,N_6628,N_6279);
nor U7299 (N_7299,N_6483,N_6749);
and U7300 (N_7300,N_6108,N_6051);
nor U7301 (N_7301,N_6229,N_6625);
xnor U7302 (N_7302,N_6734,N_6599);
nand U7303 (N_7303,N_6020,N_6086);
xor U7304 (N_7304,N_6255,N_6360);
and U7305 (N_7305,N_6414,N_6535);
nand U7306 (N_7306,N_6264,N_6224);
and U7307 (N_7307,N_6570,N_6738);
and U7308 (N_7308,N_6059,N_6599);
nand U7309 (N_7309,N_6072,N_6023);
or U7310 (N_7310,N_6555,N_6117);
nand U7311 (N_7311,N_6157,N_6646);
or U7312 (N_7312,N_6204,N_6461);
or U7313 (N_7313,N_6160,N_6544);
and U7314 (N_7314,N_6315,N_6222);
nand U7315 (N_7315,N_6749,N_6655);
nor U7316 (N_7316,N_6067,N_6498);
nor U7317 (N_7317,N_6130,N_6017);
and U7318 (N_7318,N_6535,N_6079);
and U7319 (N_7319,N_6467,N_6330);
or U7320 (N_7320,N_6445,N_6200);
and U7321 (N_7321,N_6094,N_6458);
xor U7322 (N_7322,N_6011,N_6171);
nand U7323 (N_7323,N_6331,N_6315);
and U7324 (N_7324,N_6126,N_6251);
and U7325 (N_7325,N_6250,N_6493);
and U7326 (N_7326,N_6010,N_6413);
xnor U7327 (N_7327,N_6703,N_6677);
and U7328 (N_7328,N_6093,N_6222);
and U7329 (N_7329,N_6726,N_6565);
and U7330 (N_7330,N_6242,N_6645);
and U7331 (N_7331,N_6504,N_6160);
xor U7332 (N_7332,N_6261,N_6734);
or U7333 (N_7333,N_6638,N_6490);
and U7334 (N_7334,N_6509,N_6144);
and U7335 (N_7335,N_6069,N_6396);
nor U7336 (N_7336,N_6319,N_6357);
and U7337 (N_7337,N_6033,N_6732);
or U7338 (N_7338,N_6534,N_6467);
nand U7339 (N_7339,N_6368,N_6540);
or U7340 (N_7340,N_6101,N_6045);
nor U7341 (N_7341,N_6396,N_6400);
and U7342 (N_7342,N_6015,N_6321);
xor U7343 (N_7343,N_6417,N_6566);
nand U7344 (N_7344,N_6263,N_6090);
or U7345 (N_7345,N_6320,N_6735);
nand U7346 (N_7346,N_6410,N_6503);
nor U7347 (N_7347,N_6043,N_6128);
xnor U7348 (N_7348,N_6524,N_6452);
nand U7349 (N_7349,N_6197,N_6467);
or U7350 (N_7350,N_6534,N_6446);
or U7351 (N_7351,N_6137,N_6330);
nand U7352 (N_7352,N_6005,N_6669);
nor U7353 (N_7353,N_6253,N_6732);
nand U7354 (N_7354,N_6185,N_6524);
and U7355 (N_7355,N_6062,N_6047);
xnor U7356 (N_7356,N_6620,N_6184);
and U7357 (N_7357,N_6227,N_6511);
nand U7358 (N_7358,N_6607,N_6296);
and U7359 (N_7359,N_6378,N_6721);
nand U7360 (N_7360,N_6556,N_6240);
and U7361 (N_7361,N_6534,N_6189);
or U7362 (N_7362,N_6194,N_6359);
nor U7363 (N_7363,N_6252,N_6457);
or U7364 (N_7364,N_6149,N_6155);
and U7365 (N_7365,N_6264,N_6125);
and U7366 (N_7366,N_6592,N_6586);
or U7367 (N_7367,N_6236,N_6558);
nand U7368 (N_7368,N_6480,N_6712);
or U7369 (N_7369,N_6722,N_6169);
nand U7370 (N_7370,N_6254,N_6634);
and U7371 (N_7371,N_6087,N_6338);
nand U7372 (N_7372,N_6152,N_6252);
or U7373 (N_7373,N_6558,N_6245);
or U7374 (N_7374,N_6540,N_6338);
nand U7375 (N_7375,N_6716,N_6525);
nand U7376 (N_7376,N_6599,N_6365);
nand U7377 (N_7377,N_6361,N_6471);
xnor U7378 (N_7378,N_6370,N_6280);
and U7379 (N_7379,N_6499,N_6174);
and U7380 (N_7380,N_6349,N_6384);
xor U7381 (N_7381,N_6435,N_6546);
nor U7382 (N_7382,N_6563,N_6657);
or U7383 (N_7383,N_6095,N_6466);
xor U7384 (N_7384,N_6259,N_6099);
nor U7385 (N_7385,N_6234,N_6486);
nand U7386 (N_7386,N_6700,N_6202);
and U7387 (N_7387,N_6719,N_6419);
nand U7388 (N_7388,N_6380,N_6006);
and U7389 (N_7389,N_6281,N_6653);
xor U7390 (N_7390,N_6503,N_6412);
nor U7391 (N_7391,N_6595,N_6616);
and U7392 (N_7392,N_6632,N_6476);
and U7393 (N_7393,N_6122,N_6486);
and U7394 (N_7394,N_6554,N_6692);
nand U7395 (N_7395,N_6472,N_6136);
and U7396 (N_7396,N_6700,N_6401);
and U7397 (N_7397,N_6659,N_6608);
and U7398 (N_7398,N_6100,N_6243);
nor U7399 (N_7399,N_6517,N_6311);
xor U7400 (N_7400,N_6086,N_6639);
nor U7401 (N_7401,N_6017,N_6644);
nand U7402 (N_7402,N_6714,N_6094);
nor U7403 (N_7403,N_6259,N_6186);
and U7404 (N_7404,N_6452,N_6032);
nor U7405 (N_7405,N_6070,N_6313);
nor U7406 (N_7406,N_6014,N_6526);
nor U7407 (N_7407,N_6506,N_6009);
or U7408 (N_7408,N_6060,N_6543);
nor U7409 (N_7409,N_6182,N_6699);
and U7410 (N_7410,N_6748,N_6172);
or U7411 (N_7411,N_6484,N_6391);
and U7412 (N_7412,N_6587,N_6017);
or U7413 (N_7413,N_6682,N_6487);
xnor U7414 (N_7414,N_6456,N_6046);
xnor U7415 (N_7415,N_6639,N_6097);
nor U7416 (N_7416,N_6528,N_6184);
or U7417 (N_7417,N_6252,N_6718);
nor U7418 (N_7418,N_6234,N_6310);
nor U7419 (N_7419,N_6319,N_6342);
and U7420 (N_7420,N_6193,N_6066);
xor U7421 (N_7421,N_6586,N_6389);
nand U7422 (N_7422,N_6253,N_6546);
and U7423 (N_7423,N_6092,N_6545);
or U7424 (N_7424,N_6214,N_6097);
nand U7425 (N_7425,N_6631,N_6055);
nand U7426 (N_7426,N_6698,N_6058);
or U7427 (N_7427,N_6588,N_6635);
and U7428 (N_7428,N_6128,N_6358);
nand U7429 (N_7429,N_6070,N_6725);
or U7430 (N_7430,N_6385,N_6137);
or U7431 (N_7431,N_6305,N_6157);
nand U7432 (N_7432,N_6685,N_6072);
xnor U7433 (N_7433,N_6301,N_6715);
and U7434 (N_7434,N_6597,N_6674);
nand U7435 (N_7435,N_6136,N_6650);
nor U7436 (N_7436,N_6254,N_6132);
nand U7437 (N_7437,N_6005,N_6429);
and U7438 (N_7438,N_6321,N_6239);
or U7439 (N_7439,N_6694,N_6394);
nand U7440 (N_7440,N_6481,N_6121);
nor U7441 (N_7441,N_6542,N_6307);
nor U7442 (N_7442,N_6098,N_6293);
and U7443 (N_7443,N_6616,N_6476);
and U7444 (N_7444,N_6469,N_6143);
nand U7445 (N_7445,N_6034,N_6186);
nor U7446 (N_7446,N_6728,N_6543);
or U7447 (N_7447,N_6684,N_6445);
xor U7448 (N_7448,N_6599,N_6615);
nand U7449 (N_7449,N_6598,N_6345);
nor U7450 (N_7450,N_6395,N_6511);
nor U7451 (N_7451,N_6684,N_6444);
nand U7452 (N_7452,N_6022,N_6520);
nand U7453 (N_7453,N_6639,N_6022);
and U7454 (N_7454,N_6683,N_6594);
or U7455 (N_7455,N_6533,N_6276);
or U7456 (N_7456,N_6246,N_6008);
or U7457 (N_7457,N_6122,N_6666);
xnor U7458 (N_7458,N_6091,N_6307);
nand U7459 (N_7459,N_6361,N_6566);
or U7460 (N_7460,N_6210,N_6397);
nor U7461 (N_7461,N_6178,N_6404);
nand U7462 (N_7462,N_6164,N_6133);
nor U7463 (N_7463,N_6612,N_6494);
nand U7464 (N_7464,N_6322,N_6006);
or U7465 (N_7465,N_6456,N_6501);
and U7466 (N_7466,N_6199,N_6738);
nor U7467 (N_7467,N_6713,N_6365);
nand U7468 (N_7468,N_6600,N_6267);
nor U7469 (N_7469,N_6328,N_6617);
nand U7470 (N_7470,N_6543,N_6308);
nand U7471 (N_7471,N_6715,N_6640);
nor U7472 (N_7472,N_6281,N_6678);
xor U7473 (N_7473,N_6316,N_6370);
nor U7474 (N_7474,N_6190,N_6460);
xnor U7475 (N_7475,N_6340,N_6723);
nor U7476 (N_7476,N_6120,N_6511);
and U7477 (N_7477,N_6686,N_6458);
nand U7478 (N_7478,N_6079,N_6555);
nand U7479 (N_7479,N_6009,N_6223);
nand U7480 (N_7480,N_6356,N_6706);
or U7481 (N_7481,N_6433,N_6084);
nor U7482 (N_7482,N_6116,N_6719);
and U7483 (N_7483,N_6221,N_6350);
nor U7484 (N_7484,N_6394,N_6368);
nand U7485 (N_7485,N_6184,N_6456);
nand U7486 (N_7486,N_6413,N_6701);
or U7487 (N_7487,N_6634,N_6083);
nor U7488 (N_7488,N_6257,N_6637);
and U7489 (N_7489,N_6327,N_6212);
or U7490 (N_7490,N_6656,N_6275);
and U7491 (N_7491,N_6642,N_6425);
and U7492 (N_7492,N_6453,N_6657);
and U7493 (N_7493,N_6222,N_6188);
or U7494 (N_7494,N_6283,N_6055);
nand U7495 (N_7495,N_6444,N_6534);
nand U7496 (N_7496,N_6250,N_6129);
or U7497 (N_7497,N_6209,N_6543);
and U7498 (N_7498,N_6073,N_6521);
nor U7499 (N_7499,N_6018,N_6505);
and U7500 (N_7500,N_7287,N_7230);
xor U7501 (N_7501,N_7015,N_6937);
and U7502 (N_7502,N_7452,N_6980);
xnor U7503 (N_7503,N_7194,N_7434);
nand U7504 (N_7504,N_6966,N_7227);
nand U7505 (N_7505,N_7242,N_7326);
and U7506 (N_7506,N_6972,N_7276);
and U7507 (N_7507,N_6781,N_7265);
xor U7508 (N_7508,N_6885,N_7299);
or U7509 (N_7509,N_6750,N_6840);
nand U7510 (N_7510,N_6896,N_7302);
nand U7511 (N_7511,N_7125,N_6927);
and U7512 (N_7512,N_7359,N_6921);
and U7513 (N_7513,N_7049,N_6905);
nor U7514 (N_7514,N_7419,N_7007);
nand U7515 (N_7515,N_7033,N_7457);
nand U7516 (N_7516,N_7338,N_7271);
nand U7517 (N_7517,N_6890,N_6917);
nand U7518 (N_7518,N_7274,N_6982);
nand U7519 (N_7519,N_7108,N_7171);
xor U7520 (N_7520,N_7480,N_7013);
nand U7521 (N_7521,N_7121,N_7406);
nor U7522 (N_7522,N_6872,N_6929);
nand U7523 (N_7523,N_7346,N_7167);
or U7524 (N_7524,N_7428,N_6898);
nand U7525 (N_7525,N_7047,N_6847);
nor U7526 (N_7526,N_6884,N_6908);
nor U7527 (N_7527,N_7268,N_7247);
nand U7528 (N_7528,N_7120,N_7127);
nor U7529 (N_7529,N_7040,N_7239);
or U7530 (N_7530,N_6763,N_6958);
nand U7531 (N_7531,N_6957,N_7348);
or U7532 (N_7532,N_7106,N_7499);
nor U7533 (N_7533,N_7158,N_7012);
or U7534 (N_7534,N_7141,N_7357);
or U7535 (N_7535,N_7107,N_6837);
or U7536 (N_7536,N_7301,N_7386);
or U7537 (N_7537,N_6772,N_7124);
nor U7538 (N_7538,N_7298,N_7196);
and U7539 (N_7539,N_6904,N_7113);
nand U7540 (N_7540,N_6783,N_7062);
and U7541 (N_7541,N_7061,N_7427);
and U7542 (N_7542,N_7495,N_7005);
nand U7543 (N_7543,N_6989,N_7334);
or U7544 (N_7544,N_6955,N_7305);
nand U7545 (N_7545,N_6899,N_6756);
and U7546 (N_7546,N_7214,N_7039);
nand U7547 (N_7547,N_7168,N_7477);
xnor U7548 (N_7548,N_7447,N_7387);
or U7549 (N_7549,N_7414,N_6861);
nor U7550 (N_7550,N_6753,N_6997);
or U7551 (N_7551,N_7232,N_7486);
or U7552 (N_7552,N_7407,N_7281);
or U7553 (N_7553,N_7426,N_7014);
and U7554 (N_7554,N_6953,N_7489);
nand U7555 (N_7555,N_7116,N_6770);
and U7556 (N_7556,N_6968,N_7174);
nor U7557 (N_7557,N_7439,N_7019);
nand U7558 (N_7558,N_7320,N_6792);
nor U7559 (N_7559,N_7064,N_7077);
nor U7560 (N_7560,N_6876,N_7137);
or U7561 (N_7561,N_7494,N_7467);
and U7562 (N_7562,N_6823,N_7279);
xnor U7563 (N_7563,N_7004,N_7170);
and U7564 (N_7564,N_7068,N_6780);
nor U7565 (N_7565,N_6900,N_6888);
and U7566 (N_7566,N_7138,N_6999);
nand U7567 (N_7567,N_6799,N_7184);
and U7568 (N_7568,N_7311,N_7316);
or U7569 (N_7569,N_7011,N_7337);
nor U7570 (N_7570,N_6863,N_6962);
nand U7571 (N_7571,N_7104,N_6873);
nor U7572 (N_7572,N_7169,N_7295);
and U7573 (N_7573,N_7045,N_7403);
nand U7574 (N_7574,N_6846,N_7275);
xor U7575 (N_7575,N_7297,N_7092);
nor U7576 (N_7576,N_7384,N_7154);
nor U7577 (N_7577,N_6942,N_6752);
xnor U7578 (N_7578,N_6889,N_6887);
or U7579 (N_7579,N_6926,N_7074);
nor U7580 (N_7580,N_7289,N_7260);
and U7581 (N_7581,N_7048,N_7450);
nand U7582 (N_7582,N_7160,N_7270);
or U7583 (N_7583,N_7059,N_6786);
xnor U7584 (N_7584,N_7222,N_6848);
nand U7585 (N_7585,N_7296,N_7441);
xnor U7586 (N_7586,N_7416,N_7351);
nor U7587 (N_7587,N_6924,N_6893);
nand U7588 (N_7588,N_6931,N_7021);
xor U7589 (N_7589,N_6862,N_6869);
xor U7590 (N_7590,N_7038,N_6782);
nor U7591 (N_7591,N_7091,N_6995);
nand U7592 (N_7592,N_6932,N_7140);
nor U7593 (N_7593,N_7433,N_6762);
or U7594 (N_7594,N_7462,N_7231);
or U7595 (N_7595,N_7136,N_6883);
nor U7596 (N_7596,N_6916,N_7478);
nand U7597 (N_7597,N_7240,N_6991);
or U7598 (N_7598,N_7490,N_7037);
nand U7599 (N_7599,N_6813,N_6907);
nor U7600 (N_7600,N_7318,N_7129);
nor U7601 (N_7601,N_7304,N_7458);
and U7602 (N_7602,N_6842,N_7466);
nand U7603 (N_7603,N_6914,N_7056);
nor U7604 (N_7604,N_7029,N_7375);
and U7605 (N_7605,N_7044,N_7468);
nand U7606 (N_7606,N_7415,N_7492);
nor U7607 (N_7607,N_7109,N_7358);
or U7608 (N_7608,N_7204,N_7421);
or U7609 (N_7609,N_7224,N_6886);
nand U7610 (N_7610,N_7119,N_7321);
nand U7611 (N_7611,N_7202,N_6833);
or U7612 (N_7612,N_7130,N_7273);
or U7613 (N_7613,N_7382,N_6874);
nand U7614 (N_7614,N_7392,N_6766);
or U7615 (N_7615,N_7070,N_6860);
or U7616 (N_7616,N_6755,N_7461);
or U7617 (N_7617,N_7149,N_6771);
nand U7618 (N_7618,N_6858,N_7484);
nand U7619 (N_7619,N_6979,N_6785);
nand U7620 (N_7620,N_7391,N_7278);
nor U7621 (N_7621,N_6938,N_7464);
nand U7622 (N_7622,N_6910,N_7031);
nand U7623 (N_7623,N_6844,N_6764);
and U7624 (N_7624,N_6987,N_6796);
nor U7625 (N_7625,N_6943,N_7020);
and U7626 (N_7626,N_6951,N_7253);
or U7627 (N_7627,N_6952,N_7395);
nor U7628 (N_7628,N_6773,N_7185);
nand U7629 (N_7629,N_7042,N_7094);
nand U7630 (N_7630,N_7103,N_7465);
and U7631 (N_7631,N_6948,N_7442);
nor U7632 (N_7632,N_7422,N_7425);
and U7633 (N_7633,N_7379,N_7444);
nand U7634 (N_7634,N_6967,N_7207);
or U7635 (N_7635,N_7055,N_6903);
nand U7636 (N_7636,N_7206,N_7446);
and U7637 (N_7637,N_7163,N_7397);
xor U7638 (N_7638,N_6801,N_6841);
and U7639 (N_7639,N_7372,N_7235);
and U7640 (N_7640,N_7072,N_7388);
nor U7641 (N_7641,N_6870,N_7219);
and U7642 (N_7642,N_7215,N_7144);
nor U7643 (N_7643,N_7355,N_7132);
nand U7644 (N_7644,N_6923,N_7177);
nand U7645 (N_7645,N_7327,N_7365);
and U7646 (N_7646,N_7369,N_7436);
nand U7647 (N_7647,N_7491,N_6949);
nor U7648 (N_7648,N_6909,N_7420);
or U7649 (N_7649,N_7114,N_7079);
or U7650 (N_7650,N_7455,N_7225);
or U7651 (N_7651,N_7374,N_7394);
nor U7652 (N_7652,N_6965,N_7023);
nand U7653 (N_7653,N_6895,N_6864);
and U7654 (N_7654,N_6875,N_6960);
nand U7655 (N_7655,N_6919,N_7353);
or U7656 (N_7656,N_7306,N_6826);
or U7657 (N_7657,N_7449,N_7371);
and U7658 (N_7658,N_7146,N_7314);
nor U7659 (N_7659,N_7411,N_7498);
nor U7660 (N_7660,N_7463,N_7344);
and U7661 (N_7661,N_6757,N_7310);
nor U7662 (N_7662,N_7341,N_7319);
xnor U7663 (N_7663,N_6838,N_7035);
xor U7664 (N_7664,N_7487,N_7437);
or U7665 (N_7665,N_6839,N_6877);
or U7666 (N_7666,N_7071,N_7026);
xnor U7667 (N_7667,N_7046,N_6930);
xnor U7668 (N_7668,N_7131,N_7165);
xnor U7669 (N_7669,N_7368,N_6777);
nor U7670 (N_7670,N_7364,N_6808);
nor U7671 (N_7671,N_7256,N_7161);
and U7672 (N_7672,N_7145,N_6822);
nand U7673 (N_7673,N_7417,N_7356);
and U7674 (N_7674,N_7332,N_7361);
nand U7675 (N_7675,N_7376,N_6829);
nor U7676 (N_7676,N_6815,N_7402);
or U7677 (N_7677,N_6800,N_7085);
xor U7678 (N_7678,N_6998,N_7389);
or U7679 (N_7679,N_7259,N_7111);
or U7680 (N_7680,N_7248,N_7251);
or U7681 (N_7681,N_7135,N_7134);
nor U7682 (N_7682,N_7313,N_6956);
or U7683 (N_7683,N_7067,N_7234);
nor U7684 (N_7684,N_6939,N_6936);
nand U7685 (N_7685,N_6897,N_6810);
and U7686 (N_7686,N_6761,N_6825);
or U7687 (N_7687,N_7191,N_7432);
nand U7688 (N_7688,N_6767,N_7431);
xor U7689 (N_7689,N_6835,N_7459);
or U7690 (N_7690,N_7473,N_7350);
or U7691 (N_7691,N_7352,N_7093);
and U7692 (N_7692,N_7405,N_6986);
or U7693 (N_7693,N_6768,N_7244);
and U7694 (N_7694,N_7331,N_7166);
xnor U7695 (N_7695,N_7156,N_7159);
nor U7696 (N_7696,N_6769,N_6868);
or U7697 (N_7697,N_7126,N_7201);
nor U7698 (N_7698,N_6928,N_7367);
nand U7699 (N_7699,N_7142,N_6881);
nor U7700 (N_7700,N_7303,N_7220);
or U7701 (N_7701,N_7460,N_6775);
xnor U7702 (N_7702,N_7176,N_7211);
nor U7703 (N_7703,N_6880,N_7410);
and U7704 (N_7704,N_7399,N_6849);
and U7705 (N_7705,N_7323,N_7083);
and U7706 (N_7706,N_6831,N_7181);
nand U7707 (N_7707,N_7272,N_7285);
xor U7708 (N_7708,N_6854,N_6865);
nand U7709 (N_7709,N_6894,N_7485);
and U7710 (N_7710,N_6918,N_7451);
nand U7711 (N_7711,N_7221,N_7258);
nand U7712 (N_7712,N_7366,N_7254);
nand U7713 (N_7713,N_6959,N_7223);
nor U7714 (N_7714,N_7099,N_6915);
and U7715 (N_7715,N_7267,N_7117);
xor U7716 (N_7716,N_7342,N_7312);
or U7717 (N_7717,N_7470,N_7190);
nand U7718 (N_7718,N_7123,N_7363);
or U7719 (N_7719,N_6984,N_6845);
nor U7720 (N_7720,N_7218,N_7022);
nand U7721 (N_7721,N_7370,N_6790);
xnor U7722 (N_7722,N_6906,N_7000);
nor U7723 (N_7723,N_7180,N_7139);
xnor U7724 (N_7724,N_7241,N_6912);
nand U7725 (N_7725,N_6993,N_7330);
nor U7726 (N_7726,N_6954,N_7294);
nand U7727 (N_7727,N_6983,N_7153);
or U7728 (N_7728,N_6867,N_7243);
and U7729 (N_7729,N_6795,N_7252);
nand U7730 (N_7730,N_7418,N_7017);
or U7731 (N_7731,N_7122,N_7237);
and U7732 (N_7732,N_6811,N_7381);
or U7733 (N_7733,N_7378,N_6961);
nand U7734 (N_7734,N_7065,N_7233);
or U7735 (N_7735,N_7110,N_7148);
nand U7736 (N_7736,N_6827,N_7291);
or U7737 (N_7737,N_6940,N_7043);
xor U7738 (N_7738,N_7151,N_7288);
nor U7739 (N_7739,N_7347,N_7472);
nand U7740 (N_7740,N_7277,N_6812);
nor U7741 (N_7741,N_6882,N_6760);
or U7742 (N_7742,N_6765,N_6788);
nand U7743 (N_7743,N_7424,N_6797);
and U7744 (N_7744,N_7089,N_6922);
and U7745 (N_7745,N_7009,N_6935);
xnor U7746 (N_7746,N_7325,N_7335);
xor U7747 (N_7747,N_7456,N_7423);
or U7748 (N_7748,N_7345,N_7095);
or U7749 (N_7749,N_7333,N_6806);
nor U7750 (N_7750,N_7292,N_7102);
nand U7751 (N_7751,N_7096,N_7228);
and U7752 (N_7752,N_7157,N_7317);
nand U7753 (N_7753,N_6776,N_7474);
nand U7754 (N_7754,N_7250,N_6851);
nor U7755 (N_7755,N_6856,N_7112);
nand U7756 (N_7756,N_7283,N_7343);
and U7757 (N_7757,N_7380,N_7198);
and U7758 (N_7758,N_7401,N_7262);
nor U7759 (N_7759,N_6778,N_6804);
or U7760 (N_7760,N_7147,N_7360);
and U7761 (N_7761,N_7390,N_6824);
nor U7762 (N_7762,N_6866,N_7128);
nand U7763 (N_7763,N_7018,N_7229);
xnor U7764 (N_7764,N_6817,N_7078);
and U7765 (N_7765,N_7322,N_7186);
nand U7766 (N_7766,N_7377,N_7060);
nand U7767 (N_7767,N_7404,N_7249);
and U7768 (N_7768,N_6970,N_6941);
nor U7769 (N_7769,N_7027,N_7282);
or U7770 (N_7770,N_7188,N_6901);
nand U7771 (N_7771,N_7409,N_6859);
nand U7772 (N_7772,N_7084,N_7100);
nand U7773 (N_7773,N_6974,N_7440);
nand U7774 (N_7774,N_7238,N_6857);
nand U7775 (N_7775,N_7309,N_7082);
nor U7776 (N_7776,N_6946,N_7430);
xnor U7777 (N_7777,N_7398,N_6830);
nor U7778 (N_7778,N_7088,N_7090);
nand U7779 (N_7779,N_7408,N_7324);
or U7780 (N_7780,N_7193,N_6911);
or U7781 (N_7781,N_6794,N_7385);
nor U7782 (N_7782,N_7340,N_7143);
nand U7783 (N_7783,N_7483,N_7471);
and U7784 (N_7784,N_7179,N_7175);
nand U7785 (N_7785,N_7087,N_7307);
or U7786 (N_7786,N_7453,N_7028);
nand U7787 (N_7787,N_7263,N_7257);
nor U7788 (N_7788,N_7073,N_6981);
or U7789 (N_7789,N_7481,N_6934);
or U7790 (N_7790,N_6759,N_7066);
nor U7791 (N_7791,N_7032,N_6996);
xor U7792 (N_7792,N_7203,N_7209);
nor U7793 (N_7793,N_7349,N_6802);
nor U7794 (N_7794,N_6751,N_7226);
xnor U7795 (N_7795,N_7199,N_7172);
xor U7796 (N_7796,N_7069,N_7236);
or U7797 (N_7797,N_6994,N_7476);
nand U7798 (N_7798,N_7155,N_6879);
or U7799 (N_7799,N_7362,N_7445);
nand U7800 (N_7800,N_6969,N_6892);
xor U7801 (N_7801,N_6971,N_7150);
or U7802 (N_7802,N_6992,N_7086);
and U7803 (N_7803,N_7058,N_7438);
nor U7804 (N_7804,N_7400,N_7076);
nand U7805 (N_7805,N_7210,N_7162);
or U7806 (N_7806,N_7016,N_6843);
and U7807 (N_7807,N_7030,N_6990);
or U7808 (N_7808,N_7024,N_7200);
nand U7809 (N_7809,N_7006,N_7057);
or U7810 (N_7810,N_7469,N_6828);
xnor U7811 (N_7811,N_7189,N_6758);
or U7812 (N_7812,N_7001,N_7197);
nand U7813 (N_7813,N_6809,N_7255);
nand U7814 (N_7814,N_6976,N_6818);
or U7815 (N_7815,N_6933,N_7195);
nand U7816 (N_7816,N_7183,N_6853);
nor U7817 (N_7817,N_7493,N_7328);
and U7818 (N_7818,N_6836,N_7008);
and U7819 (N_7819,N_7264,N_6774);
and U7820 (N_7820,N_7010,N_6834);
nor U7821 (N_7821,N_6787,N_6871);
and U7822 (N_7822,N_7213,N_7383);
or U7823 (N_7823,N_7482,N_7290);
or U7824 (N_7824,N_6805,N_7329);
xnor U7825 (N_7825,N_6816,N_7097);
nand U7826 (N_7826,N_7053,N_6988);
nand U7827 (N_7827,N_7336,N_6793);
nor U7828 (N_7828,N_6950,N_6807);
nand U7829 (N_7829,N_7034,N_6789);
or U7830 (N_7830,N_7497,N_6820);
nand U7831 (N_7831,N_6791,N_7339);
and U7832 (N_7832,N_6975,N_6878);
and U7833 (N_7833,N_7105,N_7036);
or U7834 (N_7834,N_7479,N_7488);
and U7835 (N_7835,N_7269,N_7393);
and U7836 (N_7836,N_6784,N_7054);
or U7837 (N_7837,N_7075,N_7003);
nand U7838 (N_7838,N_6855,N_7152);
and U7839 (N_7839,N_6964,N_6891);
nand U7840 (N_7840,N_7261,N_6920);
nand U7841 (N_7841,N_7429,N_6779);
and U7842 (N_7842,N_7396,N_7293);
nor U7843 (N_7843,N_7212,N_7052);
nor U7844 (N_7844,N_7041,N_6947);
or U7845 (N_7845,N_6985,N_7308);
nor U7846 (N_7846,N_7205,N_7435);
xnor U7847 (N_7847,N_6814,N_7187);
or U7848 (N_7848,N_7412,N_6973);
nor U7849 (N_7849,N_7315,N_7354);
and U7850 (N_7850,N_7280,N_7373);
and U7851 (N_7851,N_6821,N_7475);
xnor U7852 (N_7852,N_7050,N_7081);
xor U7853 (N_7853,N_7133,N_7080);
and U7854 (N_7854,N_7178,N_6803);
and U7855 (N_7855,N_7246,N_7182);
xnor U7856 (N_7856,N_7300,N_7025);
or U7857 (N_7857,N_7164,N_7448);
and U7858 (N_7858,N_6798,N_6850);
nor U7859 (N_7859,N_7443,N_7063);
or U7860 (N_7860,N_7413,N_7454);
xnor U7861 (N_7861,N_6832,N_6978);
xnor U7862 (N_7862,N_7192,N_6925);
and U7863 (N_7863,N_7217,N_7266);
nand U7864 (N_7864,N_7101,N_7173);
xor U7865 (N_7865,N_7284,N_7118);
xor U7866 (N_7866,N_6944,N_6963);
nor U7867 (N_7867,N_6902,N_7216);
nor U7868 (N_7868,N_6913,N_7002);
xor U7869 (N_7869,N_7208,N_7245);
nor U7870 (N_7870,N_6852,N_6945);
nor U7871 (N_7871,N_7115,N_6754);
nand U7872 (N_7872,N_7496,N_6977);
and U7873 (N_7873,N_6819,N_7286);
or U7874 (N_7874,N_7051,N_7098);
or U7875 (N_7875,N_7413,N_7426);
nor U7876 (N_7876,N_7020,N_6900);
nand U7877 (N_7877,N_7343,N_7113);
or U7878 (N_7878,N_7465,N_6774);
nand U7879 (N_7879,N_7268,N_6751);
nor U7880 (N_7880,N_7041,N_7360);
or U7881 (N_7881,N_7004,N_6874);
and U7882 (N_7882,N_7132,N_7375);
nand U7883 (N_7883,N_6886,N_7120);
and U7884 (N_7884,N_6785,N_7469);
or U7885 (N_7885,N_7177,N_7277);
or U7886 (N_7886,N_7387,N_7494);
and U7887 (N_7887,N_6978,N_7029);
nor U7888 (N_7888,N_6889,N_7438);
and U7889 (N_7889,N_7295,N_7244);
and U7890 (N_7890,N_7147,N_7169);
and U7891 (N_7891,N_7328,N_7350);
or U7892 (N_7892,N_7046,N_7483);
or U7893 (N_7893,N_6789,N_7289);
nor U7894 (N_7894,N_7234,N_7116);
or U7895 (N_7895,N_7358,N_7027);
nor U7896 (N_7896,N_7089,N_7140);
nor U7897 (N_7897,N_6783,N_6810);
xor U7898 (N_7898,N_7464,N_7020);
or U7899 (N_7899,N_7034,N_6787);
and U7900 (N_7900,N_6951,N_7372);
nor U7901 (N_7901,N_7368,N_6934);
nand U7902 (N_7902,N_7311,N_6909);
nor U7903 (N_7903,N_7302,N_7272);
nor U7904 (N_7904,N_7326,N_7267);
nand U7905 (N_7905,N_7464,N_7410);
nand U7906 (N_7906,N_6786,N_7317);
nor U7907 (N_7907,N_6866,N_6814);
or U7908 (N_7908,N_6941,N_7310);
or U7909 (N_7909,N_7016,N_6926);
nor U7910 (N_7910,N_7457,N_6996);
nor U7911 (N_7911,N_7070,N_6834);
nor U7912 (N_7912,N_7147,N_7428);
or U7913 (N_7913,N_7059,N_7354);
or U7914 (N_7914,N_6937,N_7256);
xnor U7915 (N_7915,N_6815,N_7451);
or U7916 (N_7916,N_7367,N_7285);
nand U7917 (N_7917,N_7301,N_6890);
nor U7918 (N_7918,N_7209,N_6842);
nand U7919 (N_7919,N_7323,N_7221);
and U7920 (N_7920,N_7145,N_7278);
or U7921 (N_7921,N_7201,N_7436);
or U7922 (N_7922,N_7101,N_7035);
and U7923 (N_7923,N_7457,N_6842);
or U7924 (N_7924,N_7266,N_6916);
or U7925 (N_7925,N_6913,N_6847);
nand U7926 (N_7926,N_7360,N_7336);
and U7927 (N_7927,N_7100,N_7299);
or U7928 (N_7928,N_7182,N_6876);
or U7929 (N_7929,N_6808,N_7273);
or U7930 (N_7930,N_6750,N_7480);
and U7931 (N_7931,N_7069,N_7257);
or U7932 (N_7932,N_6947,N_6830);
nor U7933 (N_7933,N_6982,N_6801);
and U7934 (N_7934,N_7299,N_7318);
nor U7935 (N_7935,N_7033,N_6838);
nor U7936 (N_7936,N_7087,N_7089);
nand U7937 (N_7937,N_6891,N_7420);
nand U7938 (N_7938,N_7159,N_6891);
nor U7939 (N_7939,N_7283,N_7116);
nand U7940 (N_7940,N_7027,N_7175);
nand U7941 (N_7941,N_7291,N_7078);
and U7942 (N_7942,N_6886,N_6940);
and U7943 (N_7943,N_7399,N_7054);
nor U7944 (N_7944,N_7029,N_6991);
nor U7945 (N_7945,N_7128,N_7466);
or U7946 (N_7946,N_6856,N_7069);
nand U7947 (N_7947,N_7291,N_7225);
or U7948 (N_7948,N_6930,N_7370);
nor U7949 (N_7949,N_7017,N_6880);
xor U7950 (N_7950,N_7227,N_7130);
xnor U7951 (N_7951,N_7119,N_7443);
or U7952 (N_7952,N_6964,N_6920);
or U7953 (N_7953,N_7339,N_7411);
and U7954 (N_7954,N_7072,N_7341);
or U7955 (N_7955,N_7179,N_6969);
xor U7956 (N_7956,N_7020,N_7250);
and U7957 (N_7957,N_6990,N_7290);
or U7958 (N_7958,N_7151,N_7019);
nand U7959 (N_7959,N_7343,N_7340);
and U7960 (N_7960,N_7403,N_6849);
nand U7961 (N_7961,N_7297,N_6762);
xnor U7962 (N_7962,N_7117,N_7443);
or U7963 (N_7963,N_7481,N_6913);
or U7964 (N_7964,N_7150,N_7262);
nor U7965 (N_7965,N_7037,N_7069);
or U7966 (N_7966,N_6772,N_7463);
or U7967 (N_7967,N_7051,N_7332);
nor U7968 (N_7968,N_7069,N_7362);
or U7969 (N_7969,N_7366,N_7107);
nand U7970 (N_7970,N_7075,N_7053);
and U7971 (N_7971,N_7288,N_7141);
and U7972 (N_7972,N_6755,N_6899);
or U7973 (N_7973,N_7442,N_7456);
nor U7974 (N_7974,N_7448,N_7472);
nor U7975 (N_7975,N_7365,N_7182);
xor U7976 (N_7976,N_6925,N_7444);
or U7977 (N_7977,N_7436,N_6870);
nor U7978 (N_7978,N_7092,N_6783);
or U7979 (N_7979,N_6828,N_6842);
and U7980 (N_7980,N_7188,N_7228);
nor U7981 (N_7981,N_6779,N_7206);
nand U7982 (N_7982,N_7155,N_7135);
and U7983 (N_7983,N_7072,N_7125);
and U7984 (N_7984,N_6879,N_7114);
nor U7985 (N_7985,N_6821,N_7470);
and U7986 (N_7986,N_6854,N_7180);
or U7987 (N_7987,N_7261,N_7020);
nand U7988 (N_7988,N_7243,N_6870);
nor U7989 (N_7989,N_7283,N_7251);
and U7990 (N_7990,N_7409,N_7261);
and U7991 (N_7991,N_7080,N_7420);
nand U7992 (N_7992,N_7148,N_7480);
nand U7993 (N_7993,N_7470,N_7097);
or U7994 (N_7994,N_6761,N_7490);
xor U7995 (N_7995,N_7024,N_6797);
or U7996 (N_7996,N_7208,N_6898);
and U7997 (N_7997,N_7323,N_6937);
and U7998 (N_7998,N_7274,N_7387);
nand U7999 (N_7999,N_7230,N_7066);
or U8000 (N_8000,N_7378,N_6933);
nor U8001 (N_8001,N_6802,N_6759);
and U8002 (N_8002,N_6888,N_6980);
xnor U8003 (N_8003,N_7096,N_6957);
xnor U8004 (N_8004,N_7396,N_7440);
or U8005 (N_8005,N_7312,N_7462);
nor U8006 (N_8006,N_7481,N_7366);
nor U8007 (N_8007,N_7289,N_7276);
or U8008 (N_8008,N_7465,N_7120);
or U8009 (N_8009,N_6983,N_7109);
and U8010 (N_8010,N_7115,N_6885);
or U8011 (N_8011,N_6795,N_7108);
or U8012 (N_8012,N_7213,N_7140);
and U8013 (N_8013,N_6910,N_6792);
nand U8014 (N_8014,N_6753,N_6768);
or U8015 (N_8015,N_6966,N_6888);
or U8016 (N_8016,N_7467,N_6994);
nand U8017 (N_8017,N_6981,N_7209);
nor U8018 (N_8018,N_6983,N_7450);
nand U8019 (N_8019,N_7477,N_7112);
nand U8020 (N_8020,N_7079,N_7381);
and U8021 (N_8021,N_6839,N_7331);
nor U8022 (N_8022,N_7325,N_7109);
and U8023 (N_8023,N_7136,N_7282);
and U8024 (N_8024,N_7060,N_7149);
or U8025 (N_8025,N_7224,N_6994);
or U8026 (N_8026,N_6950,N_7190);
or U8027 (N_8027,N_6966,N_7391);
nor U8028 (N_8028,N_6849,N_7436);
xnor U8029 (N_8029,N_7205,N_7134);
and U8030 (N_8030,N_6834,N_7421);
nand U8031 (N_8031,N_7099,N_6963);
or U8032 (N_8032,N_7244,N_7466);
and U8033 (N_8033,N_7279,N_7070);
nand U8034 (N_8034,N_7160,N_7327);
xor U8035 (N_8035,N_7487,N_6899);
or U8036 (N_8036,N_7174,N_7146);
and U8037 (N_8037,N_7249,N_7442);
or U8038 (N_8038,N_7295,N_7362);
xnor U8039 (N_8039,N_6886,N_7059);
and U8040 (N_8040,N_7054,N_6912);
xor U8041 (N_8041,N_7015,N_6804);
and U8042 (N_8042,N_6865,N_7049);
nand U8043 (N_8043,N_7486,N_7298);
nand U8044 (N_8044,N_7284,N_7392);
or U8045 (N_8045,N_7302,N_7004);
or U8046 (N_8046,N_7364,N_6988);
nand U8047 (N_8047,N_6930,N_7253);
or U8048 (N_8048,N_7418,N_7071);
or U8049 (N_8049,N_6893,N_7220);
or U8050 (N_8050,N_7306,N_7090);
nor U8051 (N_8051,N_7268,N_7261);
nor U8052 (N_8052,N_7190,N_7097);
and U8053 (N_8053,N_7366,N_6938);
nor U8054 (N_8054,N_7219,N_7184);
xnor U8055 (N_8055,N_7011,N_7267);
and U8056 (N_8056,N_6878,N_7420);
nor U8057 (N_8057,N_7344,N_6822);
or U8058 (N_8058,N_6754,N_6860);
nor U8059 (N_8059,N_7150,N_7009);
nand U8060 (N_8060,N_6801,N_6825);
or U8061 (N_8061,N_6875,N_7215);
nor U8062 (N_8062,N_6790,N_7269);
or U8063 (N_8063,N_6755,N_6985);
and U8064 (N_8064,N_7011,N_7315);
nor U8065 (N_8065,N_7210,N_7456);
nand U8066 (N_8066,N_7344,N_7310);
xor U8067 (N_8067,N_6775,N_6779);
and U8068 (N_8068,N_7344,N_6776);
nor U8069 (N_8069,N_6835,N_7103);
nor U8070 (N_8070,N_6755,N_7048);
and U8071 (N_8071,N_7110,N_7378);
xor U8072 (N_8072,N_7298,N_7062);
nor U8073 (N_8073,N_6970,N_7094);
or U8074 (N_8074,N_7170,N_7338);
nor U8075 (N_8075,N_7080,N_7209);
or U8076 (N_8076,N_7079,N_7354);
and U8077 (N_8077,N_6896,N_7348);
and U8078 (N_8078,N_6768,N_7198);
and U8079 (N_8079,N_7276,N_7407);
and U8080 (N_8080,N_6807,N_7479);
or U8081 (N_8081,N_6770,N_6876);
nor U8082 (N_8082,N_7015,N_7207);
xor U8083 (N_8083,N_6969,N_7446);
nand U8084 (N_8084,N_7464,N_6774);
and U8085 (N_8085,N_7303,N_6779);
nor U8086 (N_8086,N_6950,N_7467);
xor U8087 (N_8087,N_7112,N_7324);
and U8088 (N_8088,N_7222,N_6972);
nand U8089 (N_8089,N_7146,N_7412);
nor U8090 (N_8090,N_6949,N_7264);
or U8091 (N_8091,N_7451,N_6785);
and U8092 (N_8092,N_6882,N_7093);
nand U8093 (N_8093,N_7008,N_7235);
nand U8094 (N_8094,N_7455,N_6785);
and U8095 (N_8095,N_6964,N_7373);
and U8096 (N_8096,N_6974,N_6895);
and U8097 (N_8097,N_7294,N_7093);
nor U8098 (N_8098,N_7145,N_7358);
and U8099 (N_8099,N_6755,N_6783);
and U8100 (N_8100,N_6973,N_6971);
xor U8101 (N_8101,N_7045,N_6868);
nor U8102 (N_8102,N_7221,N_7135);
or U8103 (N_8103,N_7108,N_7434);
nand U8104 (N_8104,N_7006,N_7449);
nor U8105 (N_8105,N_7433,N_7152);
nor U8106 (N_8106,N_7137,N_7291);
nand U8107 (N_8107,N_6815,N_7450);
or U8108 (N_8108,N_7406,N_7227);
and U8109 (N_8109,N_7355,N_7047);
nor U8110 (N_8110,N_7389,N_7416);
and U8111 (N_8111,N_6918,N_6880);
and U8112 (N_8112,N_6962,N_7115);
nor U8113 (N_8113,N_7071,N_7308);
or U8114 (N_8114,N_7136,N_7068);
nor U8115 (N_8115,N_7305,N_7487);
nand U8116 (N_8116,N_6774,N_6823);
xnor U8117 (N_8117,N_6993,N_6837);
and U8118 (N_8118,N_7088,N_7278);
nand U8119 (N_8119,N_7322,N_6922);
nor U8120 (N_8120,N_6831,N_6808);
or U8121 (N_8121,N_7065,N_7018);
nand U8122 (N_8122,N_7356,N_7484);
or U8123 (N_8123,N_7185,N_7224);
and U8124 (N_8124,N_7400,N_7372);
nor U8125 (N_8125,N_7084,N_6982);
or U8126 (N_8126,N_6869,N_7476);
xnor U8127 (N_8127,N_7452,N_6771);
nor U8128 (N_8128,N_7235,N_7100);
nor U8129 (N_8129,N_7431,N_6857);
and U8130 (N_8130,N_6781,N_7090);
nor U8131 (N_8131,N_7293,N_7327);
xnor U8132 (N_8132,N_7071,N_6983);
or U8133 (N_8133,N_6942,N_6990);
and U8134 (N_8134,N_7260,N_6905);
or U8135 (N_8135,N_7431,N_6837);
and U8136 (N_8136,N_6969,N_6987);
nor U8137 (N_8137,N_7127,N_7151);
and U8138 (N_8138,N_7294,N_7319);
nor U8139 (N_8139,N_7497,N_7019);
nor U8140 (N_8140,N_7043,N_6876);
or U8141 (N_8141,N_6919,N_7217);
xor U8142 (N_8142,N_6796,N_6809);
nor U8143 (N_8143,N_7092,N_7281);
nand U8144 (N_8144,N_6981,N_7406);
or U8145 (N_8145,N_7140,N_6944);
nand U8146 (N_8146,N_6989,N_6983);
nand U8147 (N_8147,N_6758,N_7252);
xnor U8148 (N_8148,N_7384,N_6945);
or U8149 (N_8149,N_6814,N_6819);
or U8150 (N_8150,N_6913,N_6935);
nand U8151 (N_8151,N_6763,N_6807);
nand U8152 (N_8152,N_7181,N_7031);
nand U8153 (N_8153,N_6772,N_7362);
nor U8154 (N_8154,N_7000,N_7312);
nand U8155 (N_8155,N_7028,N_7155);
xor U8156 (N_8156,N_6762,N_7000);
nor U8157 (N_8157,N_7234,N_7358);
and U8158 (N_8158,N_7373,N_7161);
nor U8159 (N_8159,N_7177,N_7239);
nor U8160 (N_8160,N_6954,N_7150);
nor U8161 (N_8161,N_6753,N_7377);
nand U8162 (N_8162,N_7353,N_7052);
and U8163 (N_8163,N_6898,N_6786);
xor U8164 (N_8164,N_7465,N_7490);
and U8165 (N_8165,N_7126,N_6865);
nand U8166 (N_8166,N_7075,N_7456);
and U8167 (N_8167,N_7441,N_6790);
or U8168 (N_8168,N_7398,N_7119);
and U8169 (N_8169,N_6954,N_6853);
nand U8170 (N_8170,N_6907,N_7063);
nor U8171 (N_8171,N_7417,N_6821);
and U8172 (N_8172,N_7211,N_7462);
or U8173 (N_8173,N_7297,N_7017);
nor U8174 (N_8174,N_7255,N_6951);
or U8175 (N_8175,N_7248,N_6972);
nand U8176 (N_8176,N_6992,N_6892);
or U8177 (N_8177,N_6990,N_7160);
nor U8178 (N_8178,N_7473,N_6773);
or U8179 (N_8179,N_7233,N_6915);
nand U8180 (N_8180,N_6979,N_7419);
xnor U8181 (N_8181,N_7410,N_6793);
and U8182 (N_8182,N_7474,N_7286);
nand U8183 (N_8183,N_7474,N_7193);
nand U8184 (N_8184,N_6949,N_7074);
or U8185 (N_8185,N_7044,N_7474);
or U8186 (N_8186,N_7360,N_6937);
xor U8187 (N_8187,N_7041,N_6820);
nor U8188 (N_8188,N_7324,N_6875);
and U8189 (N_8189,N_7006,N_7153);
nor U8190 (N_8190,N_6959,N_7074);
nor U8191 (N_8191,N_7364,N_6886);
or U8192 (N_8192,N_6812,N_7256);
nand U8193 (N_8193,N_7271,N_6884);
nand U8194 (N_8194,N_7145,N_7499);
and U8195 (N_8195,N_6967,N_7063);
or U8196 (N_8196,N_7047,N_7028);
or U8197 (N_8197,N_6802,N_6941);
and U8198 (N_8198,N_6868,N_6957);
and U8199 (N_8199,N_6804,N_6901);
or U8200 (N_8200,N_7412,N_7030);
nand U8201 (N_8201,N_7141,N_7172);
and U8202 (N_8202,N_6814,N_7440);
and U8203 (N_8203,N_7314,N_6790);
nand U8204 (N_8204,N_7046,N_6825);
or U8205 (N_8205,N_7378,N_7276);
nor U8206 (N_8206,N_6911,N_7160);
or U8207 (N_8207,N_6827,N_6834);
nand U8208 (N_8208,N_7197,N_6969);
nor U8209 (N_8209,N_7382,N_7104);
nor U8210 (N_8210,N_7114,N_7189);
or U8211 (N_8211,N_7449,N_6754);
nor U8212 (N_8212,N_7388,N_7317);
nand U8213 (N_8213,N_7057,N_7160);
nand U8214 (N_8214,N_7494,N_7306);
and U8215 (N_8215,N_7316,N_7040);
nor U8216 (N_8216,N_6950,N_6862);
nand U8217 (N_8217,N_7023,N_6818);
and U8218 (N_8218,N_6924,N_7469);
nand U8219 (N_8219,N_6880,N_6809);
nand U8220 (N_8220,N_6981,N_6966);
or U8221 (N_8221,N_7262,N_7318);
nor U8222 (N_8222,N_7387,N_6861);
or U8223 (N_8223,N_7357,N_7156);
or U8224 (N_8224,N_6986,N_7342);
nor U8225 (N_8225,N_7218,N_7149);
and U8226 (N_8226,N_7045,N_6799);
and U8227 (N_8227,N_7213,N_6937);
and U8228 (N_8228,N_6961,N_6807);
nand U8229 (N_8229,N_7086,N_6981);
nand U8230 (N_8230,N_7039,N_6840);
nand U8231 (N_8231,N_6922,N_7400);
xor U8232 (N_8232,N_6775,N_6984);
nand U8233 (N_8233,N_6903,N_7063);
xnor U8234 (N_8234,N_6857,N_7213);
and U8235 (N_8235,N_7490,N_6853);
and U8236 (N_8236,N_7167,N_7197);
or U8237 (N_8237,N_7405,N_6860);
xor U8238 (N_8238,N_7465,N_7209);
or U8239 (N_8239,N_7016,N_6832);
nand U8240 (N_8240,N_6792,N_7416);
or U8241 (N_8241,N_7423,N_7050);
and U8242 (N_8242,N_6831,N_6999);
xnor U8243 (N_8243,N_6867,N_6948);
xor U8244 (N_8244,N_6953,N_7270);
nor U8245 (N_8245,N_7487,N_7196);
and U8246 (N_8246,N_7310,N_6986);
xor U8247 (N_8247,N_6783,N_7007);
and U8248 (N_8248,N_7257,N_6855);
nand U8249 (N_8249,N_6785,N_7149);
nor U8250 (N_8250,N_8026,N_7830);
or U8251 (N_8251,N_8027,N_7732);
or U8252 (N_8252,N_8111,N_8007);
and U8253 (N_8253,N_7992,N_7780);
nor U8254 (N_8254,N_8132,N_7809);
nand U8255 (N_8255,N_7770,N_7647);
or U8256 (N_8256,N_7861,N_7827);
and U8257 (N_8257,N_7801,N_7936);
nor U8258 (N_8258,N_7738,N_8068);
and U8259 (N_8259,N_7857,N_8118);
xnor U8260 (N_8260,N_7989,N_7663);
and U8261 (N_8261,N_7950,N_8219);
nor U8262 (N_8262,N_8207,N_8012);
and U8263 (N_8263,N_8077,N_7561);
nor U8264 (N_8264,N_7674,N_7923);
or U8265 (N_8265,N_7626,N_7815);
nor U8266 (N_8266,N_7744,N_7838);
and U8267 (N_8267,N_7619,N_7650);
and U8268 (N_8268,N_7569,N_7695);
nand U8269 (N_8269,N_7781,N_7706);
xor U8270 (N_8270,N_8153,N_7922);
nand U8271 (N_8271,N_8208,N_8188);
or U8272 (N_8272,N_7716,N_7975);
nand U8273 (N_8273,N_7965,N_7935);
and U8274 (N_8274,N_8114,N_8190);
nand U8275 (N_8275,N_7517,N_8001);
nor U8276 (N_8276,N_7740,N_7798);
nor U8277 (N_8277,N_7546,N_7568);
or U8278 (N_8278,N_7671,N_8115);
nand U8279 (N_8279,N_8217,N_7721);
nor U8280 (N_8280,N_8195,N_7820);
and U8281 (N_8281,N_7636,N_8247);
or U8282 (N_8282,N_7694,N_7766);
nor U8283 (N_8283,N_7778,N_7967);
or U8284 (N_8284,N_7526,N_8122);
nor U8285 (N_8285,N_7842,N_7972);
and U8286 (N_8286,N_7964,N_7646);
nor U8287 (N_8287,N_8158,N_7955);
or U8288 (N_8288,N_7519,N_7714);
xnor U8289 (N_8289,N_8243,N_7513);
nand U8290 (N_8290,N_7587,N_8211);
and U8291 (N_8291,N_7712,N_7752);
or U8292 (N_8292,N_7944,N_7596);
and U8293 (N_8293,N_8245,N_7589);
and U8294 (N_8294,N_7533,N_8172);
and U8295 (N_8295,N_7993,N_7750);
and U8296 (N_8296,N_8226,N_7509);
and U8297 (N_8297,N_7786,N_8089);
and U8298 (N_8298,N_7635,N_8183);
and U8299 (N_8299,N_7860,N_7902);
nand U8300 (N_8300,N_7710,N_7537);
or U8301 (N_8301,N_8179,N_7954);
nand U8302 (N_8302,N_8167,N_8120);
nand U8303 (N_8303,N_7584,N_8006);
or U8304 (N_8304,N_8091,N_7855);
or U8305 (N_8305,N_7623,N_8055);
and U8306 (N_8306,N_7880,N_8127);
or U8307 (N_8307,N_7713,N_7545);
and U8308 (N_8308,N_7879,N_7831);
nor U8309 (N_8309,N_7631,N_8146);
or U8310 (N_8310,N_7934,N_7840);
or U8311 (N_8311,N_7620,N_7748);
xor U8312 (N_8312,N_7904,N_8223);
nand U8313 (N_8313,N_8009,N_7983);
and U8314 (N_8314,N_8229,N_8162);
nor U8315 (N_8315,N_7638,N_7867);
or U8316 (N_8316,N_7717,N_7961);
nor U8317 (N_8317,N_7814,N_7572);
or U8318 (N_8318,N_8075,N_7648);
or U8319 (N_8319,N_7667,N_7886);
nor U8320 (N_8320,N_7565,N_8192);
or U8321 (N_8321,N_7609,N_7743);
nor U8322 (N_8322,N_7624,N_7678);
nor U8323 (N_8323,N_7555,N_7615);
or U8324 (N_8324,N_7994,N_8071);
nand U8325 (N_8325,N_7977,N_7507);
nand U8326 (N_8326,N_8022,N_8094);
nand U8327 (N_8327,N_8169,N_7929);
xnor U8328 (N_8328,N_8129,N_7735);
or U8329 (N_8329,N_7554,N_8228);
or U8330 (N_8330,N_8051,N_7779);
or U8331 (N_8331,N_7919,N_7958);
or U8332 (N_8332,N_7805,N_7629);
and U8333 (N_8333,N_7693,N_8028);
or U8334 (N_8334,N_7604,N_7810);
and U8335 (N_8335,N_7811,N_7598);
or U8336 (N_8336,N_7749,N_8069);
or U8337 (N_8337,N_8239,N_7976);
nor U8338 (N_8338,N_7586,N_8103);
nor U8339 (N_8339,N_7821,N_7822);
or U8340 (N_8340,N_8102,N_8073);
nand U8341 (N_8341,N_7682,N_7816);
or U8342 (N_8342,N_8197,N_7728);
and U8343 (N_8343,N_7847,N_7567);
nor U8344 (N_8344,N_7829,N_8064);
nor U8345 (N_8345,N_7709,N_8076);
nor U8346 (N_8346,N_7872,N_7981);
xor U8347 (N_8347,N_7918,N_8106);
or U8348 (N_8348,N_7558,N_8086);
and U8349 (N_8349,N_8136,N_8005);
nor U8350 (N_8350,N_7907,N_8033);
nor U8351 (N_8351,N_7542,N_7874);
nor U8352 (N_8352,N_7696,N_8084);
and U8353 (N_8353,N_7697,N_7617);
and U8354 (N_8354,N_7762,N_8047);
nand U8355 (N_8355,N_8139,N_7530);
and U8356 (N_8356,N_7962,N_8154);
and U8357 (N_8357,N_7906,N_7737);
nand U8358 (N_8358,N_7873,N_7633);
and U8359 (N_8359,N_7689,N_7729);
nor U8360 (N_8360,N_8016,N_8175);
nor U8361 (N_8361,N_8096,N_7910);
nand U8362 (N_8362,N_7828,N_7684);
or U8363 (N_8363,N_8220,N_7951);
or U8364 (N_8364,N_7512,N_7772);
or U8365 (N_8365,N_7639,N_7601);
nand U8366 (N_8366,N_8019,N_8194);
and U8367 (N_8367,N_7621,N_7941);
and U8368 (N_8368,N_7754,N_8090);
nor U8369 (N_8369,N_7928,N_7869);
nor U8370 (N_8370,N_7597,N_7582);
nand U8371 (N_8371,N_8109,N_7571);
and U8372 (N_8372,N_8198,N_7850);
or U8373 (N_8373,N_7618,N_8024);
and U8374 (N_8374,N_7912,N_7503);
nor U8375 (N_8375,N_8107,N_7812);
xor U8376 (N_8376,N_7681,N_7726);
nand U8377 (N_8377,N_7819,N_7970);
nor U8378 (N_8378,N_8203,N_7607);
nand U8379 (N_8379,N_7769,N_8238);
and U8380 (N_8380,N_7871,N_7557);
or U8381 (N_8381,N_7913,N_7968);
nor U8382 (N_8382,N_7783,N_7903);
or U8383 (N_8383,N_7751,N_8215);
nand U8384 (N_8384,N_7818,N_7916);
and U8385 (N_8385,N_8044,N_8053);
nor U8386 (N_8386,N_7660,N_8140);
xor U8387 (N_8387,N_7654,N_7945);
nand U8388 (N_8388,N_7909,N_8065);
or U8389 (N_8389,N_7562,N_7643);
xor U8390 (N_8390,N_7984,N_7692);
or U8391 (N_8391,N_7501,N_7883);
or U8392 (N_8392,N_7771,N_8126);
or U8393 (N_8393,N_8248,N_7564);
or U8394 (N_8394,N_7759,N_7825);
nand U8395 (N_8395,N_7524,N_8095);
nand U8396 (N_8396,N_8130,N_7730);
and U8397 (N_8397,N_7698,N_7576);
nand U8398 (N_8398,N_7525,N_8039);
or U8399 (N_8399,N_7999,N_7959);
and U8400 (N_8400,N_7908,N_8209);
and U8401 (N_8401,N_8003,N_7747);
nor U8402 (N_8402,N_7785,N_8010);
nand U8403 (N_8403,N_7553,N_8184);
or U8404 (N_8404,N_7914,N_8020);
nor U8405 (N_8405,N_8119,N_7574);
or U8406 (N_8406,N_7843,N_7612);
nor U8407 (N_8407,N_8029,N_7892);
and U8408 (N_8408,N_7990,N_7588);
nand U8409 (N_8409,N_7532,N_7949);
xor U8410 (N_8410,N_7898,N_8214);
and U8411 (N_8411,N_7602,N_7960);
or U8412 (N_8412,N_7573,N_7520);
nand U8413 (N_8413,N_7947,N_7543);
nand U8414 (N_8414,N_7703,N_8133);
and U8415 (N_8415,N_7939,N_8110);
nor U8416 (N_8416,N_8151,N_8035);
and U8417 (N_8417,N_8100,N_7865);
or U8418 (N_8418,N_7998,N_8171);
nor U8419 (N_8419,N_7773,N_7931);
nor U8420 (N_8420,N_7651,N_8123);
xor U8421 (N_8421,N_8235,N_7683);
or U8422 (N_8422,N_8045,N_7600);
and U8423 (N_8423,N_7504,N_7884);
or U8424 (N_8424,N_7784,N_7536);
and U8425 (N_8425,N_7859,N_7722);
xnor U8426 (N_8426,N_7581,N_7645);
nor U8427 (N_8427,N_7836,N_7680);
nor U8428 (N_8428,N_8116,N_7637);
nor U8429 (N_8429,N_8186,N_7862);
or U8430 (N_8430,N_7523,N_8161);
nand U8431 (N_8431,N_7566,N_7579);
or U8432 (N_8432,N_8210,N_7725);
nand U8433 (N_8433,N_7644,N_7927);
nand U8434 (N_8434,N_8117,N_7905);
or U8435 (N_8435,N_7548,N_7807);
nor U8436 (N_8436,N_8178,N_7655);
or U8437 (N_8437,N_8227,N_7788);
nand U8438 (N_8438,N_7813,N_7736);
and U8439 (N_8439,N_7767,N_7677);
nor U8440 (N_8440,N_8034,N_8049);
or U8441 (N_8441,N_7616,N_8147);
nand U8442 (N_8442,N_7630,N_7516);
and U8443 (N_8443,N_8078,N_8234);
and U8444 (N_8444,N_7594,N_8166);
nand U8445 (N_8445,N_7940,N_7665);
or U8446 (N_8446,N_7510,N_7832);
xor U8447 (N_8447,N_8141,N_7622);
nand U8448 (N_8448,N_8206,N_7870);
xnor U8449 (N_8449,N_8205,N_8185);
and U8450 (N_8450,N_7711,N_8093);
or U8451 (N_8451,N_8191,N_7793);
xor U8452 (N_8452,N_7608,N_8164);
or U8453 (N_8453,N_7917,N_8159);
nand U8454 (N_8454,N_7837,N_7800);
and U8455 (N_8455,N_7764,N_7758);
or U8456 (N_8456,N_7658,N_8070);
and U8457 (N_8457,N_7757,N_7787);
or U8458 (N_8458,N_8128,N_7527);
or U8459 (N_8459,N_8231,N_7938);
or U8460 (N_8460,N_7895,N_8101);
xnor U8461 (N_8461,N_8112,N_7823);
or U8462 (N_8462,N_8213,N_7580);
or U8463 (N_8463,N_7844,N_7834);
or U8464 (N_8464,N_8092,N_8042);
and U8465 (N_8465,N_7763,N_7980);
and U8466 (N_8466,N_7911,N_7673);
nor U8467 (N_8467,N_7614,N_7782);
nor U8468 (N_8468,N_7518,N_7887);
nand U8469 (N_8469,N_7753,N_7672);
nor U8470 (N_8470,N_7888,N_7590);
nand U8471 (N_8471,N_7632,N_7666);
or U8472 (N_8472,N_7777,N_8142);
nand U8473 (N_8473,N_7560,N_7611);
and U8474 (N_8474,N_8050,N_7659);
nand U8475 (N_8475,N_7529,N_8031);
or U8476 (N_8476,N_8156,N_7760);
nand U8477 (N_8477,N_7641,N_7889);
and U8478 (N_8478,N_8021,N_7592);
nand U8479 (N_8479,N_8168,N_8113);
nor U8480 (N_8480,N_8187,N_7704);
nand U8481 (N_8481,N_7719,N_7505);
nor U8482 (N_8482,N_8018,N_7806);
xnor U8483 (N_8483,N_7851,N_8025);
nor U8484 (N_8484,N_8225,N_7701);
and U8485 (N_8485,N_7657,N_8040);
or U8486 (N_8486,N_7705,N_8131);
xor U8487 (N_8487,N_8163,N_7656);
or U8488 (N_8488,N_7853,N_7563);
nor U8489 (N_8489,N_8013,N_8056);
and U8490 (N_8490,N_7894,N_8081);
or U8491 (N_8491,N_8189,N_8082);
xor U8492 (N_8492,N_7627,N_7790);
and U8493 (N_8493,N_7978,N_7774);
or U8494 (N_8494,N_8058,N_7963);
nor U8495 (N_8495,N_7930,N_7556);
nand U8496 (N_8496,N_7846,N_7605);
or U8497 (N_8497,N_8000,N_7803);
nand U8498 (N_8498,N_8193,N_7733);
and U8499 (N_8499,N_8043,N_7603);
nor U8500 (N_8500,N_8204,N_8216);
xnor U8501 (N_8501,N_7549,N_7897);
nand U8502 (N_8502,N_8066,N_8170);
or U8503 (N_8503,N_7686,N_7915);
and U8504 (N_8504,N_7640,N_7599);
nand U8505 (N_8505,N_8036,N_8061);
and U8506 (N_8506,N_7761,N_8023);
nor U8507 (N_8507,N_7796,N_8222);
nand U8508 (N_8508,N_7799,N_7699);
xnor U8509 (N_8509,N_7987,N_7675);
nand U8510 (N_8510,N_7539,N_8182);
nor U8511 (N_8511,N_8083,N_7731);
or U8512 (N_8512,N_7690,N_8232);
nor U8513 (N_8513,N_8038,N_7577);
nand U8514 (N_8514,N_7552,N_8138);
and U8515 (N_8515,N_8157,N_7739);
xnor U8516 (N_8516,N_7966,N_7500);
nand U8517 (N_8517,N_8074,N_7741);
nor U8518 (N_8518,N_7804,N_8165);
nand U8519 (N_8519,N_8155,N_7792);
and U8520 (N_8520,N_8032,N_7583);
xnor U8521 (N_8521,N_7864,N_7541);
or U8522 (N_8522,N_8088,N_7765);
nor U8523 (N_8523,N_7676,N_7570);
nor U8524 (N_8524,N_8011,N_8149);
or U8525 (N_8525,N_7538,N_8236);
nor U8526 (N_8526,N_7891,N_8052);
and U8527 (N_8527,N_7925,N_7926);
xnor U8528 (N_8528,N_8041,N_7890);
and U8529 (N_8529,N_7547,N_7991);
nand U8530 (N_8530,N_7937,N_8137);
or U8531 (N_8531,N_8152,N_8224);
or U8532 (N_8532,N_7795,N_8199);
nand U8533 (N_8533,N_7610,N_7802);
or U8534 (N_8534,N_7756,N_7995);
or U8535 (N_8535,N_7595,N_7997);
xnor U8536 (N_8536,N_7863,N_7971);
nor U8537 (N_8537,N_8002,N_8063);
or U8538 (N_8538,N_7535,N_7585);
or U8539 (N_8539,N_8249,N_8060);
nor U8540 (N_8540,N_7882,N_8099);
nand U8541 (N_8541,N_7852,N_7559);
and U8542 (N_8542,N_7924,N_7669);
nor U8543 (N_8543,N_8059,N_7979);
nor U8544 (N_8544,N_7824,N_7901);
nor U8545 (N_8545,N_7856,N_7575);
nand U8546 (N_8546,N_7551,N_8054);
and U8547 (N_8547,N_8145,N_7508);
nor U8548 (N_8548,N_7946,N_8048);
and U8549 (N_8549,N_7839,N_8237);
or U8550 (N_8550,N_7953,N_7833);
nand U8551 (N_8551,N_7742,N_7982);
and U8552 (N_8552,N_8135,N_7920);
nand U8553 (N_8553,N_7877,N_8098);
or U8554 (N_8554,N_7727,N_8097);
nand U8555 (N_8555,N_7734,N_7723);
nor U8556 (N_8556,N_8201,N_7956);
or U8557 (N_8557,N_7593,N_7700);
or U8558 (N_8558,N_8202,N_8180);
and U8559 (N_8559,N_8244,N_8143);
nor U8560 (N_8560,N_8079,N_8014);
and U8561 (N_8561,N_7885,N_7745);
nor U8562 (N_8562,N_7652,N_7664);
nor U8563 (N_8563,N_8046,N_8108);
nor U8564 (N_8564,N_7625,N_8242);
or U8565 (N_8565,N_8057,N_7791);
nand U8566 (N_8566,N_7948,N_7514);
nor U8567 (N_8567,N_8181,N_8150);
or U8568 (N_8568,N_7670,N_7789);
or U8569 (N_8569,N_8067,N_8173);
nand U8570 (N_8570,N_7881,N_8212);
and U8571 (N_8571,N_7817,N_8072);
nand U8572 (N_8572,N_7591,N_7841);
or U8573 (N_8573,N_7942,N_7707);
and U8574 (N_8574,N_7679,N_7578);
nand U8575 (N_8575,N_7528,N_7985);
and U8576 (N_8576,N_7775,N_7797);
or U8577 (N_8577,N_7868,N_7540);
or U8578 (N_8578,N_8105,N_8200);
or U8579 (N_8579,N_7896,N_7613);
or U8580 (N_8580,N_8240,N_7996);
nand U8581 (N_8581,N_7845,N_7534);
nor U8582 (N_8582,N_7973,N_7718);
or U8583 (N_8583,N_7685,N_7986);
or U8584 (N_8584,N_7544,N_8062);
nand U8585 (N_8585,N_8144,N_7687);
and U8586 (N_8586,N_7988,N_8030);
and U8587 (N_8587,N_8246,N_7522);
or U8588 (N_8588,N_8177,N_7661);
nand U8589 (N_8589,N_7900,N_7849);
nand U8590 (N_8590,N_8221,N_7755);
nand U8591 (N_8591,N_7969,N_7933);
or U8592 (N_8592,N_8196,N_8176);
or U8593 (N_8593,N_8230,N_7708);
and U8594 (N_8594,N_8008,N_7974);
nand U8595 (N_8595,N_8087,N_7893);
nor U8596 (N_8596,N_7878,N_7688);
or U8597 (N_8597,N_7724,N_8080);
nand U8598 (N_8598,N_8037,N_8004);
or U8599 (N_8599,N_7776,N_8134);
or U8600 (N_8600,N_8233,N_7866);
nor U8601 (N_8601,N_7746,N_7848);
nand U8602 (N_8602,N_7858,N_7943);
nand U8603 (N_8603,N_7634,N_8160);
and U8604 (N_8604,N_7952,N_7662);
xnor U8605 (N_8605,N_7642,N_7521);
or U8606 (N_8606,N_8104,N_7768);
nand U8607 (N_8607,N_7876,N_8124);
or U8608 (N_8608,N_8015,N_7691);
or U8609 (N_8609,N_7794,N_7826);
or U8610 (N_8610,N_8148,N_7515);
or U8611 (N_8611,N_7875,N_8017);
nand U8612 (N_8612,N_7835,N_8241);
or U8613 (N_8613,N_7720,N_7511);
or U8614 (N_8614,N_7715,N_8218);
nand U8615 (N_8615,N_7702,N_8121);
or U8616 (N_8616,N_8085,N_7653);
xnor U8617 (N_8617,N_7957,N_7932);
xnor U8618 (N_8618,N_7531,N_7899);
and U8619 (N_8619,N_8174,N_8125);
or U8620 (N_8620,N_7506,N_7808);
or U8621 (N_8621,N_7668,N_7550);
or U8622 (N_8622,N_7628,N_7854);
nor U8623 (N_8623,N_7921,N_7502);
or U8624 (N_8624,N_7649,N_7606);
and U8625 (N_8625,N_8127,N_7603);
nand U8626 (N_8626,N_7782,N_7841);
or U8627 (N_8627,N_7772,N_7649);
or U8628 (N_8628,N_8227,N_7775);
xnor U8629 (N_8629,N_8083,N_7974);
or U8630 (N_8630,N_8020,N_7702);
or U8631 (N_8631,N_7999,N_8203);
nor U8632 (N_8632,N_8009,N_7604);
or U8633 (N_8633,N_7552,N_7789);
or U8634 (N_8634,N_7828,N_8020);
xnor U8635 (N_8635,N_7680,N_8034);
nor U8636 (N_8636,N_7563,N_7514);
nand U8637 (N_8637,N_7728,N_8081);
and U8638 (N_8638,N_7895,N_7746);
and U8639 (N_8639,N_7816,N_7771);
or U8640 (N_8640,N_7829,N_8106);
nand U8641 (N_8641,N_7716,N_7735);
nor U8642 (N_8642,N_8125,N_7639);
nor U8643 (N_8643,N_7783,N_7565);
and U8644 (N_8644,N_7952,N_8138);
nor U8645 (N_8645,N_7749,N_7519);
xor U8646 (N_8646,N_7922,N_8166);
nor U8647 (N_8647,N_7576,N_7794);
nor U8648 (N_8648,N_8224,N_7558);
and U8649 (N_8649,N_7507,N_7781);
nor U8650 (N_8650,N_7909,N_7673);
nor U8651 (N_8651,N_7714,N_7711);
or U8652 (N_8652,N_7851,N_8164);
or U8653 (N_8653,N_7521,N_7719);
or U8654 (N_8654,N_7952,N_8182);
nor U8655 (N_8655,N_7888,N_7917);
nor U8656 (N_8656,N_7603,N_8040);
nor U8657 (N_8657,N_8044,N_8194);
and U8658 (N_8658,N_7754,N_7857);
and U8659 (N_8659,N_8048,N_7719);
and U8660 (N_8660,N_7686,N_8241);
or U8661 (N_8661,N_7602,N_7864);
nor U8662 (N_8662,N_7967,N_7548);
and U8663 (N_8663,N_8074,N_8118);
and U8664 (N_8664,N_7917,N_7722);
or U8665 (N_8665,N_8192,N_7735);
xnor U8666 (N_8666,N_8073,N_7582);
or U8667 (N_8667,N_7575,N_7957);
and U8668 (N_8668,N_7690,N_8092);
nor U8669 (N_8669,N_7989,N_7616);
nand U8670 (N_8670,N_7523,N_7753);
and U8671 (N_8671,N_7553,N_7665);
nor U8672 (N_8672,N_7642,N_8123);
and U8673 (N_8673,N_7647,N_8180);
and U8674 (N_8674,N_7658,N_8177);
nand U8675 (N_8675,N_7781,N_8107);
or U8676 (N_8676,N_7835,N_8016);
nor U8677 (N_8677,N_8040,N_7985);
or U8678 (N_8678,N_7765,N_7724);
or U8679 (N_8679,N_7515,N_7902);
nor U8680 (N_8680,N_7742,N_7912);
and U8681 (N_8681,N_7983,N_8223);
nand U8682 (N_8682,N_8200,N_7864);
nand U8683 (N_8683,N_8078,N_7792);
or U8684 (N_8684,N_8233,N_8213);
and U8685 (N_8685,N_7933,N_7771);
and U8686 (N_8686,N_8233,N_7916);
or U8687 (N_8687,N_7550,N_7999);
nand U8688 (N_8688,N_7671,N_7521);
nand U8689 (N_8689,N_8008,N_7923);
and U8690 (N_8690,N_7926,N_7698);
nor U8691 (N_8691,N_8236,N_7882);
or U8692 (N_8692,N_8156,N_7809);
xor U8693 (N_8693,N_7561,N_7638);
and U8694 (N_8694,N_7524,N_7574);
or U8695 (N_8695,N_8084,N_7785);
or U8696 (N_8696,N_7685,N_8162);
or U8697 (N_8697,N_7646,N_7847);
xor U8698 (N_8698,N_7925,N_7727);
xnor U8699 (N_8699,N_7880,N_8114);
and U8700 (N_8700,N_8217,N_8165);
or U8701 (N_8701,N_7812,N_7749);
xnor U8702 (N_8702,N_7735,N_7787);
nand U8703 (N_8703,N_8048,N_7898);
nor U8704 (N_8704,N_7900,N_7593);
nor U8705 (N_8705,N_8030,N_8140);
and U8706 (N_8706,N_7660,N_7995);
nand U8707 (N_8707,N_8051,N_7958);
nor U8708 (N_8708,N_7792,N_8112);
nor U8709 (N_8709,N_7734,N_8080);
or U8710 (N_8710,N_7896,N_7603);
nand U8711 (N_8711,N_8055,N_8048);
nor U8712 (N_8712,N_8032,N_7620);
and U8713 (N_8713,N_7931,N_8189);
or U8714 (N_8714,N_7695,N_7997);
nor U8715 (N_8715,N_8247,N_7816);
nor U8716 (N_8716,N_7657,N_7589);
or U8717 (N_8717,N_7689,N_7815);
and U8718 (N_8718,N_7649,N_7731);
nor U8719 (N_8719,N_7630,N_7537);
and U8720 (N_8720,N_8060,N_7926);
nor U8721 (N_8721,N_7824,N_7647);
or U8722 (N_8722,N_8147,N_8099);
nand U8723 (N_8723,N_8051,N_7930);
and U8724 (N_8724,N_7730,N_7985);
or U8725 (N_8725,N_7651,N_7622);
nor U8726 (N_8726,N_7551,N_7856);
xnor U8727 (N_8727,N_7948,N_7806);
or U8728 (N_8728,N_7625,N_8146);
and U8729 (N_8729,N_7576,N_8156);
and U8730 (N_8730,N_8240,N_7774);
nand U8731 (N_8731,N_7514,N_7890);
and U8732 (N_8732,N_7696,N_7840);
nor U8733 (N_8733,N_7575,N_7512);
nor U8734 (N_8734,N_7814,N_7827);
nor U8735 (N_8735,N_7538,N_8033);
or U8736 (N_8736,N_7902,N_7801);
and U8737 (N_8737,N_7825,N_8078);
nor U8738 (N_8738,N_8185,N_7998);
nand U8739 (N_8739,N_7536,N_8076);
or U8740 (N_8740,N_8111,N_8214);
nor U8741 (N_8741,N_8030,N_8100);
nor U8742 (N_8742,N_8195,N_7798);
nand U8743 (N_8743,N_7526,N_7620);
nor U8744 (N_8744,N_7645,N_7702);
and U8745 (N_8745,N_7765,N_7587);
or U8746 (N_8746,N_7716,N_7509);
and U8747 (N_8747,N_7702,N_7590);
nor U8748 (N_8748,N_8136,N_8017);
nor U8749 (N_8749,N_7958,N_8112);
and U8750 (N_8750,N_8036,N_7693);
xor U8751 (N_8751,N_8159,N_7675);
nand U8752 (N_8752,N_7718,N_7937);
nand U8753 (N_8753,N_8179,N_7532);
and U8754 (N_8754,N_7934,N_7954);
and U8755 (N_8755,N_7937,N_7607);
and U8756 (N_8756,N_7799,N_8191);
nand U8757 (N_8757,N_7647,N_8200);
nand U8758 (N_8758,N_8155,N_8167);
and U8759 (N_8759,N_8231,N_8129);
nor U8760 (N_8760,N_7541,N_7563);
and U8761 (N_8761,N_7976,N_7990);
nor U8762 (N_8762,N_7995,N_7526);
and U8763 (N_8763,N_7737,N_8124);
nor U8764 (N_8764,N_7632,N_7622);
nand U8765 (N_8765,N_7965,N_8065);
or U8766 (N_8766,N_8030,N_7548);
nor U8767 (N_8767,N_7644,N_8049);
nand U8768 (N_8768,N_7706,N_8083);
nand U8769 (N_8769,N_7617,N_8210);
nor U8770 (N_8770,N_7540,N_8083);
nand U8771 (N_8771,N_8046,N_8001);
nand U8772 (N_8772,N_7767,N_8149);
nor U8773 (N_8773,N_8158,N_7780);
nand U8774 (N_8774,N_7877,N_8214);
xnor U8775 (N_8775,N_8215,N_8087);
and U8776 (N_8776,N_8117,N_7857);
nor U8777 (N_8777,N_8085,N_8190);
xor U8778 (N_8778,N_7652,N_7910);
and U8779 (N_8779,N_7500,N_7937);
nand U8780 (N_8780,N_7538,N_7609);
and U8781 (N_8781,N_7665,N_7593);
nor U8782 (N_8782,N_8041,N_8148);
or U8783 (N_8783,N_8091,N_7846);
nor U8784 (N_8784,N_7609,N_7823);
or U8785 (N_8785,N_7894,N_7779);
and U8786 (N_8786,N_8119,N_7807);
or U8787 (N_8787,N_7876,N_7645);
nor U8788 (N_8788,N_7759,N_7594);
nor U8789 (N_8789,N_7966,N_7515);
nor U8790 (N_8790,N_7840,N_7597);
and U8791 (N_8791,N_7502,N_7607);
nor U8792 (N_8792,N_7939,N_7962);
nor U8793 (N_8793,N_8223,N_8082);
nand U8794 (N_8794,N_8164,N_7615);
or U8795 (N_8795,N_8220,N_7830);
or U8796 (N_8796,N_7601,N_8165);
or U8797 (N_8797,N_7590,N_7925);
and U8798 (N_8798,N_7981,N_7842);
and U8799 (N_8799,N_8234,N_7875);
xor U8800 (N_8800,N_7986,N_7795);
nor U8801 (N_8801,N_8164,N_7683);
and U8802 (N_8802,N_8207,N_7786);
or U8803 (N_8803,N_7797,N_7532);
and U8804 (N_8804,N_7919,N_7648);
nor U8805 (N_8805,N_8087,N_8081);
or U8806 (N_8806,N_7712,N_8027);
nor U8807 (N_8807,N_8090,N_7552);
or U8808 (N_8808,N_7771,N_7620);
nor U8809 (N_8809,N_8047,N_7924);
nand U8810 (N_8810,N_7888,N_7709);
or U8811 (N_8811,N_7632,N_7755);
nand U8812 (N_8812,N_7895,N_7832);
or U8813 (N_8813,N_7692,N_7611);
nor U8814 (N_8814,N_7878,N_7991);
or U8815 (N_8815,N_7545,N_7850);
and U8816 (N_8816,N_8156,N_8147);
nor U8817 (N_8817,N_7583,N_7729);
or U8818 (N_8818,N_7880,N_8065);
and U8819 (N_8819,N_7619,N_8129);
xnor U8820 (N_8820,N_7583,N_8207);
nand U8821 (N_8821,N_8062,N_8219);
or U8822 (N_8822,N_7631,N_8184);
nor U8823 (N_8823,N_8247,N_7943);
nand U8824 (N_8824,N_8102,N_8113);
xor U8825 (N_8825,N_8018,N_8002);
or U8826 (N_8826,N_7650,N_7574);
and U8827 (N_8827,N_7902,N_8197);
and U8828 (N_8828,N_7994,N_7762);
or U8829 (N_8829,N_8216,N_7927);
nor U8830 (N_8830,N_8106,N_8088);
nand U8831 (N_8831,N_7868,N_7803);
and U8832 (N_8832,N_7819,N_7909);
nor U8833 (N_8833,N_8054,N_8167);
nor U8834 (N_8834,N_7746,N_7783);
and U8835 (N_8835,N_7656,N_7701);
nand U8836 (N_8836,N_7649,N_8033);
xnor U8837 (N_8837,N_8172,N_8236);
nor U8838 (N_8838,N_7599,N_7573);
nor U8839 (N_8839,N_7675,N_7714);
nand U8840 (N_8840,N_7623,N_8195);
or U8841 (N_8841,N_7924,N_7882);
and U8842 (N_8842,N_7822,N_8060);
and U8843 (N_8843,N_7909,N_7514);
and U8844 (N_8844,N_7617,N_8172);
nand U8845 (N_8845,N_7746,N_7575);
or U8846 (N_8846,N_7845,N_7753);
nor U8847 (N_8847,N_8095,N_8242);
nand U8848 (N_8848,N_7766,N_7997);
or U8849 (N_8849,N_8128,N_8173);
xor U8850 (N_8850,N_7780,N_8168);
and U8851 (N_8851,N_8208,N_7539);
xor U8852 (N_8852,N_8050,N_7706);
and U8853 (N_8853,N_8008,N_7715);
and U8854 (N_8854,N_8033,N_7826);
or U8855 (N_8855,N_7663,N_8019);
or U8856 (N_8856,N_7662,N_7545);
nor U8857 (N_8857,N_7621,N_7628);
or U8858 (N_8858,N_7851,N_7813);
nand U8859 (N_8859,N_8194,N_8159);
or U8860 (N_8860,N_7722,N_7599);
nand U8861 (N_8861,N_7543,N_8048);
and U8862 (N_8862,N_8014,N_8184);
nor U8863 (N_8863,N_7576,N_7976);
nor U8864 (N_8864,N_7642,N_7696);
or U8865 (N_8865,N_7669,N_7712);
and U8866 (N_8866,N_8144,N_7677);
and U8867 (N_8867,N_7851,N_8084);
and U8868 (N_8868,N_7531,N_7963);
and U8869 (N_8869,N_8123,N_7670);
and U8870 (N_8870,N_8070,N_7920);
and U8871 (N_8871,N_8198,N_7766);
nor U8872 (N_8872,N_7704,N_7994);
and U8873 (N_8873,N_8090,N_8233);
and U8874 (N_8874,N_8217,N_7943);
nor U8875 (N_8875,N_7814,N_7821);
xor U8876 (N_8876,N_8050,N_7586);
xor U8877 (N_8877,N_8155,N_7607);
nand U8878 (N_8878,N_7572,N_8073);
or U8879 (N_8879,N_7708,N_7922);
or U8880 (N_8880,N_7825,N_7814);
nand U8881 (N_8881,N_8011,N_7943);
or U8882 (N_8882,N_8103,N_8139);
or U8883 (N_8883,N_8209,N_8052);
nand U8884 (N_8884,N_7714,N_7826);
or U8885 (N_8885,N_7554,N_7778);
nor U8886 (N_8886,N_7687,N_8099);
nor U8887 (N_8887,N_8009,N_7547);
and U8888 (N_8888,N_7805,N_7627);
nor U8889 (N_8889,N_7613,N_7659);
or U8890 (N_8890,N_7839,N_7577);
or U8891 (N_8891,N_8130,N_7693);
nand U8892 (N_8892,N_7767,N_7944);
and U8893 (N_8893,N_8031,N_7518);
nor U8894 (N_8894,N_7936,N_7702);
nor U8895 (N_8895,N_8219,N_7536);
nor U8896 (N_8896,N_7907,N_8203);
or U8897 (N_8897,N_7846,N_8114);
nand U8898 (N_8898,N_7775,N_8185);
nor U8899 (N_8899,N_7541,N_7724);
nand U8900 (N_8900,N_7651,N_7710);
and U8901 (N_8901,N_8127,N_8113);
nor U8902 (N_8902,N_7953,N_7829);
nor U8903 (N_8903,N_8249,N_8079);
and U8904 (N_8904,N_7900,N_8231);
nor U8905 (N_8905,N_7522,N_8236);
and U8906 (N_8906,N_7697,N_8160);
nand U8907 (N_8907,N_7618,N_7876);
nor U8908 (N_8908,N_7513,N_7577);
and U8909 (N_8909,N_7727,N_7720);
nand U8910 (N_8910,N_8184,N_7741);
nand U8911 (N_8911,N_7859,N_8152);
nor U8912 (N_8912,N_7681,N_7779);
nor U8913 (N_8913,N_8173,N_7866);
and U8914 (N_8914,N_8187,N_8014);
nor U8915 (N_8915,N_7829,N_7974);
nor U8916 (N_8916,N_8060,N_7968);
and U8917 (N_8917,N_7651,N_7897);
xor U8918 (N_8918,N_8038,N_7910);
or U8919 (N_8919,N_8118,N_8003);
and U8920 (N_8920,N_7616,N_8059);
xnor U8921 (N_8921,N_8052,N_7522);
nor U8922 (N_8922,N_7668,N_7502);
xor U8923 (N_8923,N_8186,N_7642);
nor U8924 (N_8924,N_8052,N_7724);
nor U8925 (N_8925,N_8052,N_7892);
nor U8926 (N_8926,N_7932,N_8107);
nor U8927 (N_8927,N_7756,N_7975);
or U8928 (N_8928,N_7549,N_8236);
nand U8929 (N_8929,N_7531,N_7592);
or U8930 (N_8930,N_7832,N_7513);
nand U8931 (N_8931,N_7843,N_8029);
nor U8932 (N_8932,N_7620,N_7602);
and U8933 (N_8933,N_7755,N_7502);
nand U8934 (N_8934,N_7578,N_7899);
xnor U8935 (N_8935,N_7634,N_7772);
nor U8936 (N_8936,N_7942,N_7500);
and U8937 (N_8937,N_8140,N_7804);
xnor U8938 (N_8938,N_8094,N_8228);
nand U8939 (N_8939,N_7734,N_8139);
or U8940 (N_8940,N_7762,N_7551);
nor U8941 (N_8941,N_7875,N_7767);
and U8942 (N_8942,N_8097,N_7535);
nand U8943 (N_8943,N_8204,N_8040);
nor U8944 (N_8944,N_7537,N_8107);
nand U8945 (N_8945,N_7750,N_7820);
xor U8946 (N_8946,N_7639,N_7581);
and U8947 (N_8947,N_7964,N_8138);
and U8948 (N_8948,N_7555,N_8238);
or U8949 (N_8949,N_8028,N_8140);
nor U8950 (N_8950,N_8216,N_7808);
nor U8951 (N_8951,N_7832,N_8233);
nand U8952 (N_8952,N_7792,N_7841);
and U8953 (N_8953,N_7835,N_7840);
and U8954 (N_8954,N_7657,N_7731);
nand U8955 (N_8955,N_7585,N_7783);
nand U8956 (N_8956,N_8228,N_7836);
nor U8957 (N_8957,N_7887,N_7895);
or U8958 (N_8958,N_7872,N_7875);
or U8959 (N_8959,N_8220,N_8084);
nor U8960 (N_8960,N_7576,N_8224);
nor U8961 (N_8961,N_7574,N_7823);
and U8962 (N_8962,N_8049,N_8041);
or U8963 (N_8963,N_7769,N_7881);
and U8964 (N_8964,N_7552,N_8174);
nand U8965 (N_8965,N_7690,N_8108);
and U8966 (N_8966,N_7662,N_7644);
or U8967 (N_8967,N_7760,N_8105);
nor U8968 (N_8968,N_7996,N_7812);
nor U8969 (N_8969,N_8062,N_8071);
and U8970 (N_8970,N_7846,N_8062);
xor U8971 (N_8971,N_7949,N_7803);
xnor U8972 (N_8972,N_7721,N_8013);
or U8973 (N_8973,N_7519,N_7980);
nor U8974 (N_8974,N_7563,N_7803);
and U8975 (N_8975,N_7860,N_7717);
and U8976 (N_8976,N_7539,N_8049);
or U8977 (N_8977,N_7959,N_8140);
and U8978 (N_8978,N_7917,N_7952);
nor U8979 (N_8979,N_8096,N_7946);
nand U8980 (N_8980,N_7618,N_7660);
xor U8981 (N_8981,N_8074,N_8183);
nand U8982 (N_8982,N_7736,N_8106);
and U8983 (N_8983,N_7680,N_8193);
xnor U8984 (N_8984,N_8090,N_7965);
nand U8985 (N_8985,N_7966,N_7661);
or U8986 (N_8986,N_8188,N_8102);
or U8987 (N_8987,N_7869,N_8088);
nor U8988 (N_8988,N_7899,N_7906);
or U8989 (N_8989,N_7925,N_7688);
xnor U8990 (N_8990,N_7894,N_7881);
xor U8991 (N_8991,N_8139,N_8022);
xor U8992 (N_8992,N_8152,N_8200);
or U8993 (N_8993,N_7985,N_7694);
and U8994 (N_8994,N_7933,N_7524);
nand U8995 (N_8995,N_7982,N_7693);
and U8996 (N_8996,N_7849,N_8101);
and U8997 (N_8997,N_8031,N_7685);
nor U8998 (N_8998,N_7576,N_7731);
nand U8999 (N_8999,N_7575,N_7541);
or U9000 (N_9000,N_8958,N_8637);
and U9001 (N_9001,N_8257,N_8437);
nor U9002 (N_9002,N_8862,N_8779);
xnor U9003 (N_9003,N_8641,N_8802);
nand U9004 (N_9004,N_8457,N_8893);
nor U9005 (N_9005,N_8913,N_8730);
and U9006 (N_9006,N_8633,N_8382);
and U9007 (N_9007,N_8552,N_8657);
nor U9008 (N_9008,N_8423,N_8291);
xnor U9009 (N_9009,N_8817,N_8426);
nor U9010 (N_9010,N_8561,N_8911);
nor U9011 (N_9011,N_8790,N_8683);
xnor U9012 (N_9012,N_8290,N_8370);
xnor U9013 (N_9013,N_8313,N_8334);
nor U9014 (N_9014,N_8615,N_8727);
nor U9015 (N_9015,N_8937,N_8448);
nand U9016 (N_9016,N_8517,N_8999);
nand U9017 (N_9017,N_8472,N_8302);
and U9018 (N_9018,N_8551,N_8281);
or U9019 (N_9019,N_8521,N_8651);
and U9020 (N_9020,N_8411,N_8758);
nor U9021 (N_9021,N_8721,N_8665);
xnor U9022 (N_9022,N_8587,N_8420);
nor U9023 (N_9023,N_8687,N_8724);
nand U9024 (N_9024,N_8394,N_8498);
and U9025 (N_9025,N_8503,N_8546);
nand U9026 (N_9026,N_8908,N_8873);
nand U9027 (N_9027,N_8963,N_8629);
and U9028 (N_9028,N_8415,N_8664);
and U9029 (N_9029,N_8941,N_8754);
nand U9030 (N_9030,N_8703,N_8276);
nand U9031 (N_9031,N_8445,N_8306);
nor U9032 (N_9032,N_8593,N_8976);
xor U9033 (N_9033,N_8524,N_8901);
xor U9034 (N_9034,N_8384,N_8786);
xnor U9035 (N_9035,N_8607,N_8381);
nor U9036 (N_9036,N_8851,N_8856);
nand U9037 (N_9037,N_8975,N_8289);
or U9038 (N_9038,N_8295,N_8816);
nand U9039 (N_9039,N_8396,N_8293);
or U9040 (N_9040,N_8858,N_8461);
or U9041 (N_9041,N_8333,N_8272);
xor U9042 (N_9042,N_8386,N_8511);
or U9043 (N_9043,N_8948,N_8389);
or U9044 (N_9044,N_8667,N_8533);
or U9045 (N_9045,N_8788,N_8857);
nor U9046 (N_9046,N_8844,N_8717);
or U9047 (N_9047,N_8823,N_8564);
nor U9048 (N_9048,N_8403,N_8638);
or U9049 (N_9049,N_8861,N_8716);
and U9050 (N_9050,N_8864,N_8798);
xnor U9051 (N_9051,N_8617,N_8526);
and U9052 (N_9052,N_8782,N_8506);
nor U9053 (N_9053,N_8795,N_8902);
or U9054 (N_9054,N_8694,N_8635);
and U9055 (N_9055,N_8892,N_8537);
or U9056 (N_9056,N_8977,N_8375);
nor U9057 (N_9057,N_8297,N_8631);
xnor U9058 (N_9058,N_8841,N_8460);
nand U9059 (N_9059,N_8992,N_8956);
and U9060 (N_9060,N_8287,N_8601);
and U9061 (N_9061,N_8377,N_8895);
nand U9062 (N_9062,N_8422,N_8704);
xnor U9063 (N_9063,N_8510,N_8725);
nand U9064 (N_9064,N_8769,N_8990);
and U9065 (N_9065,N_8904,N_8489);
or U9066 (N_9066,N_8714,N_8345);
xnor U9067 (N_9067,N_8888,N_8357);
nor U9068 (N_9068,N_8602,N_8673);
and U9069 (N_9069,N_8924,N_8292);
nand U9070 (N_9070,N_8965,N_8989);
or U9071 (N_9071,N_8628,N_8718);
or U9072 (N_9072,N_8652,N_8960);
and U9073 (N_9073,N_8525,N_8926);
and U9074 (N_9074,N_8273,N_8860);
and U9075 (N_9075,N_8974,N_8402);
nand U9076 (N_9076,N_8656,N_8486);
xnor U9077 (N_9077,N_8449,N_8259);
nand U9078 (N_9078,N_8262,N_8418);
or U9079 (N_9079,N_8532,N_8740);
and U9080 (N_9080,N_8613,N_8496);
nand U9081 (N_9081,N_8907,N_8845);
nor U9082 (N_9082,N_8854,N_8722);
nor U9083 (N_9083,N_8658,N_8563);
xor U9084 (N_9084,N_8986,N_8996);
and U9085 (N_9085,N_8750,N_8550);
or U9086 (N_9086,N_8390,N_8995);
or U9087 (N_9087,N_8910,N_8570);
nand U9088 (N_9088,N_8916,N_8360);
xnor U9089 (N_9089,N_8475,N_8938);
nand U9090 (N_9090,N_8547,N_8485);
or U9091 (N_9091,N_8267,N_8930);
nor U9092 (N_9092,N_8378,N_8969);
nor U9093 (N_9093,N_8771,N_8369);
or U9094 (N_9094,N_8476,N_8367);
nor U9095 (N_9095,N_8534,N_8590);
xor U9096 (N_9096,N_8421,N_8441);
and U9097 (N_9097,N_8897,N_8275);
or U9098 (N_9098,N_8586,N_8775);
nand U9099 (N_9099,N_8604,N_8312);
and U9100 (N_9100,N_8591,N_8905);
xnor U9101 (N_9101,N_8654,N_8834);
nand U9102 (N_9102,N_8444,N_8899);
and U9103 (N_9103,N_8344,N_8253);
and U9104 (N_9104,N_8536,N_8516);
and U9105 (N_9105,N_8573,N_8686);
nor U9106 (N_9106,N_8791,N_8934);
nor U9107 (N_9107,N_8874,N_8745);
nor U9108 (N_9108,N_8349,N_8734);
xnor U9109 (N_9109,N_8464,N_8728);
or U9110 (N_9110,N_8364,N_8880);
nand U9111 (N_9111,N_8839,N_8626);
nand U9112 (N_9112,N_8338,N_8978);
xor U9113 (N_9113,N_8509,N_8413);
nand U9114 (N_9114,N_8630,N_8584);
nand U9115 (N_9115,N_8764,N_8599);
nor U9116 (N_9116,N_8720,N_8715);
or U9117 (N_9117,N_8685,N_8636);
nor U9118 (N_9118,N_8719,N_8330);
xnor U9119 (N_9119,N_8539,N_8871);
nor U9120 (N_9120,N_8768,N_8661);
or U9121 (N_9121,N_8575,N_8912);
xor U9122 (N_9122,N_8391,N_8723);
nor U9123 (N_9123,N_8774,N_8668);
nand U9124 (N_9124,N_8699,N_8530);
xnor U9125 (N_9125,N_8806,N_8675);
and U9126 (N_9126,N_8605,N_8314);
and U9127 (N_9127,N_8255,N_8821);
and U9128 (N_9128,N_8863,N_8434);
and U9129 (N_9129,N_8739,N_8680);
and U9130 (N_9130,N_8340,N_8596);
and U9131 (N_9131,N_8470,N_8726);
or U9132 (N_9132,N_8940,N_8918);
and U9133 (N_9133,N_8927,N_8603);
and U9134 (N_9134,N_8853,N_8608);
or U9135 (N_9135,N_8450,N_8358);
xnor U9136 (N_9136,N_8380,N_8909);
nand U9137 (N_9137,N_8556,N_8454);
or U9138 (N_9138,N_8371,N_8693);
nor U9139 (N_9139,N_8799,N_8884);
nor U9140 (N_9140,N_8811,N_8316);
xnor U9141 (N_9141,N_8438,N_8753);
and U9142 (N_9142,N_8640,N_8288);
nand U9143 (N_9143,N_8712,N_8757);
and U9144 (N_9144,N_8350,N_8898);
nor U9145 (N_9145,N_8512,N_8698);
nand U9146 (N_9146,N_8639,N_8416);
nand U9147 (N_9147,N_8588,N_8671);
or U9148 (N_9148,N_8343,N_8408);
or U9149 (N_9149,N_8317,N_8468);
nor U9150 (N_9150,N_8428,N_8818);
xnor U9151 (N_9151,N_8585,N_8677);
and U9152 (N_9152,N_8362,N_8881);
or U9153 (N_9153,N_8436,N_8875);
and U9154 (N_9154,N_8632,N_8906);
or U9155 (N_9155,N_8644,N_8501);
xor U9156 (N_9156,N_8766,N_8508);
or U9157 (N_9157,N_8886,N_8373);
and U9158 (N_9158,N_8756,N_8277);
nor U9159 (N_9159,N_8466,N_8385);
nand U9160 (N_9160,N_8323,N_8372);
xnor U9161 (N_9161,N_8932,N_8269);
or U9162 (N_9162,N_8462,N_8493);
nor U9163 (N_9163,N_8321,N_8700);
nor U9164 (N_9164,N_8335,N_8392);
and U9165 (N_9165,N_8645,N_8732);
or U9166 (N_9166,N_8773,N_8478);
and U9167 (N_9167,N_8882,N_8580);
nor U9168 (N_9168,N_8813,N_8548);
and U9169 (N_9169,N_8705,N_8947);
nor U9170 (N_9170,N_8847,N_8835);
nor U9171 (N_9171,N_8827,N_8304);
nand U9172 (N_9172,N_8964,N_8792);
and U9173 (N_9173,N_8830,N_8611);
nand U9174 (N_9174,N_8520,N_8824);
or U9175 (N_9175,N_8305,N_8810);
nand U9176 (N_9176,N_8252,N_8256);
xor U9177 (N_9177,N_8697,N_8443);
xnor U9178 (N_9178,N_8264,N_8737);
or U9179 (N_9179,N_8459,N_8622);
or U9180 (N_9180,N_8417,N_8527);
nor U9181 (N_9181,N_8981,N_8336);
nor U9182 (N_9182,N_8568,N_8574);
or U9183 (N_9183,N_8327,N_8936);
nand U9184 (N_9184,N_8351,N_8553);
and U9185 (N_9185,N_8455,N_8970);
and U9186 (N_9186,N_8966,N_8801);
or U9187 (N_9187,N_8746,N_8619);
or U9188 (N_9188,N_8943,N_8560);
and U9189 (N_9189,N_8832,N_8961);
or U9190 (N_9190,N_8933,N_8366);
and U9191 (N_9191,N_8274,N_8967);
and U9192 (N_9192,N_8915,N_8598);
or U9193 (N_9193,N_8263,N_8528);
nor U9194 (N_9194,N_8258,N_8777);
nand U9195 (N_9195,N_8648,N_8308);
or U9196 (N_9196,N_8365,N_8544);
and U9197 (N_9197,N_8543,N_8804);
or U9198 (N_9198,N_8618,N_8789);
or U9199 (N_9199,N_8278,N_8987);
and U9200 (N_9200,N_8922,N_8833);
nand U9201 (N_9201,N_8738,N_8713);
or U9202 (N_9202,N_8634,N_8866);
or U9203 (N_9203,N_8794,N_8407);
and U9204 (N_9204,N_8676,N_8749);
or U9205 (N_9205,N_8849,N_8928);
nand U9206 (N_9206,N_8925,N_8581);
or U9207 (N_9207,N_8250,N_8931);
nand U9208 (N_9208,N_8557,N_8567);
nor U9209 (N_9209,N_8812,N_8346);
and U9210 (N_9210,N_8623,N_8710);
xor U9211 (N_9211,N_8820,N_8848);
nand U9212 (N_9212,N_8807,N_8896);
nand U9213 (N_9213,N_8979,N_8435);
or U9214 (N_9214,N_8439,N_8660);
nor U9215 (N_9215,N_8747,N_8968);
or U9216 (N_9216,N_8577,N_8554);
nand U9217 (N_9217,N_8594,N_8669);
or U9218 (N_9218,N_8662,N_8299);
or U9219 (N_9219,N_8376,N_8867);
nand U9220 (N_9220,N_8379,N_8303);
nor U9221 (N_9221,N_8315,N_8878);
nand U9222 (N_9222,N_8569,N_8649);
or U9223 (N_9223,N_8784,N_8513);
or U9224 (N_9224,N_8555,N_8328);
xor U9225 (N_9225,N_8424,N_8920);
nand U9226 (N_9226,N_8751,N_8458);
and U9227 (N_9227,N_8514,N_8492);
or U9228 (N_9228,N_8760,N_8331);
nand U9229 (N_9229,N_8488,N_8405);
nor U9230 (N_9230,N_8280,N_8972);
nor U9231 (N_9231,N_8765,N_8497);
nor U9232 (N_9232,N_8393,N_8776);
or U9233 (N_9233,N_8842,N_8410);
nand U9234 (N_9234,N_8988,N_8284);
and U9235 (N_9235,N_8404,N_8374);
nor U9236 (N_9236,N_8770,N_8809);
xor U9237 (N_9237,N_8531,N_8610);
nor U9238 (N_9238,N_8491,N_8950);
and U9239 (N_9239,N_8761,N_8324);
nor U9240 (N_9240,N_8282,N_8625);
and U9241 (N_9241,N_8480,N_8692);
or U9242 (N_9242,N_8891,N_8877);
or U9243 (N_9243,N_8781,N_8887);
or U9244 (N_9244,N_8566,N_8953);
nor U9245 (N_9245,N_8744,N_8341);
or U9246 (N_9246,N_8592,N_8944);
and U9247 (N_9247,N_8653,N_8442);
or U9248 (N_9248,N_8843,N_8465);
or U9249 (N_9249,N_8535,N_8957);
and U9250 (N_9250,N_8432,N_8748);
nand U9251 (N_9251,N_8883,N_8778);
xor U9252 (N_9252,N_8310,N_8542);
or U9253 (N_9253,N_8627,N_8736);
nor U9254 (N_9254,N_8296,N_8828);
nand U9255 (N_9255,N_8419,N_8271);
nand U9256 (N_9256,N_8923,N_8733);
and U9257 (N_9257,N_8889,N_8939);
or U9258 (N_9258,N_8691,N_8954);
and U9259 (N_9259,N_8982,N_8935);
nand U9260 (N_9260,N_8595,N_8971);
or U9261 (N_9261,N_8870,N_8348);
xor U9262 (N_9262,N_8541,N_8279);
nand U9263 (N_9263,N_8518,N_8474);
or U9264 (N_9264,N_8285,N_8759);
and U9265 (N_9265,N_8919,N_8589);
and U9266 (N_9266,N_8325,N_8356);
nor U9267 (N_9267,N_8646,N_8479);
nor U9268 (N_9268,N_8872,N_8558);
and U9269 (N_9269,N_8650,N_8852);
or U9270 (N_9270,N_8743,N_8785);
nor U9271 (N_9271,N_8742,N_8682);
or U9272 (N_9272,N_8500,N_8412);
and U9273 (N_9273,N_8578,N_8406);
nand U9274 (N_9274,N_8672,N_8505);
nand U9275 (N_9275,N_8451,N_8300);
nand U9276 (N_9276,N_8565,N_8354);
nand U9277 (N_9277,N_8684,N_8819);
nor U9278 (N_9278,N_8890,N_8483);
nor U9279 (N_9279,N_8793,N_8855);
nor U9280 (N_9280,N_8355,N_8609);
nor U9281 (N_9281,N_8452,N_8398);
or U9282 (N_9282,N_8582,N_8741);
or U9283 (N_9283,N_8708,N_8689);
nand U9284 (N_9284,N_8467,N_8797);
or U9285 (N_9285,N_8701,N_8318);
and U9286 (N_9286,N_8709,N_8523);
and U9287 (N_9287,N_8850,N_8326);
and U9288 (N_9288,N_8984,N_8616);
and U9289 (N_9289,N_8767,N_8666);
and U9290 (N_9290,N_8456,N_8929);
xnor U9291 (N_9291,N_8755,N_8332);
or U9292 (N_9292,N_8283,N_8549);
xnor U9293 (N_9293,N_8307,N_8894);
xor U9294 (N_9294,N_8973,N_8729);
nor U9295 (N_9295,N_8495,N_8859);
nand U9296 (N_9296,N_8998,N_8337);
nor U9297 (N_9297,N_8469,N_8900);
nor U9298 (N_9298,N_8414,N_8397);
nand U9299 (N_9299,N_8903,N_8353);
or U9300 (N_9300,N_8363,N_8688);
and U9301 (N_9301,N_8731,N_8387);
or U9302 (N_9302,N_8361,N_8446);
nand U9303 (N_9303,N_8266,N_8286);
or U9304 (N_9304,N_8579,N_8829);
nor U9305 (N_9305,N_8805,N_8347);
nand U9306 (N_9306,N_8914,N_8803);
xnor U9307 (N_9307,N_8383,N_8846);
or U9308 (N_9308,N_8955,N_8427);
and U9309 (N_9309,N_8951,N_8942);
nand U9310 (N_9310,N_8440,N_8320);
nor U9311 (N_9311,N_8869,N_8559);
nand U9312 (N_9312,N_8695,N_8762);
xor U9313 (N_9313,N_8985,N_8322);
and U9314 (N_9314,N_8409,N_8808);
or U9315 (N_9315,N_8294,N_8752);
nand U9316 (N_9316,N_8368,N_8837);
or U9317 (N_9317,N_8572,N_8342);
or U9318 (N_9318,N_8621,N_8388);
and U9319 (N_9319,N_8983,N_8504);
or U9320 (N_9320,N_8494,N_8945);
nand U9321 (N_9321,N_8836,N_8484);
nor U9322 (N_9322,N_8879,N_8309);
nor U9323 (N_9323,N_8311,N_8576);
nand U9324 (N_9324,N_8401,N_8822);
and U9325 (N_9325,N_8433,N_8254);
nand U9326 (N_9326,N_8429,N_8329);
or U9327 (N_9327,N_8562,N_8921);
and U9328 (N_9328,N_8431,N_8959);
or U9329 (N_9329,N_8831,N_8826);
or U9330 (N_9330,N_8711,N_8814);
nor U9331 (N_9331,N_8670,N_8800);
nand U9332 (N_9332,N_8430,N_8359);
and U9333 (N_9333,N_8690,N_8519);
or U9334 (N_9334,N_8868,N_8647);
and U9335 (N_9335,N_8796,N_8696);
and U9336 (N_9336,N_8763,N_8477);
or U9337 (N_9337,N_8481,N_8991);
nand U9338 (N_9338,N_8735,N_8301);
or U9339 (N_9339,N_8490,N_8962);
nand U9340 (N_9340,N_8597,N_8298);
nor U9341 (N_9341,N_8499,N_8946);
and U9342 (N_9342,N_8917,N_8706);
or U9343 (N_9343,N_8952,N_8453);
nand U9344 (N_9344,N_8624,N_8463);
nand U9345 (N_9345,N_8702,N_8655);
xnor U9346 (N_9346,N_8674,N_8949);
or U9347 (N_9347,N_8659,N_8614);
nor U9348 (N_9348,N_8251,N_8339);
nand U9349 (N_9349,N_8612,N_8487);
nor U9350 (N_9350,N_8522,N_8352);
nor U9351 (N_9351,N_8681,N_8876);
and U9352 (N_9352,N_8482,N_8840);
or U9353 (N_9353,N_8865,N_8620);
or U9354 (N_9354,N_8471,N_8265);
and U9355 (N_9355,N_8260,N_8583);
nand U9356 (N_9356,N_8642,N_8606);
and U9357 (N_9357,N_8980,N_8507);
and U9358 (N_9358,N_8425,N_8825);
or U9359 (N_9359,N_8261,N_8571);
or U9360 (N_9360,N_8473,N_8783);
nor U9361 (N_9361,N_8997,N_8545);
xnor U9362 (N_9362,N_8707,N_8787);
nand U9363 (N_9363,N_8993,N_8815);
and U9364 (N_9364,N_8780,N_8502);
xor U9365 (N_9365,N_8678,N_8319);
nand U9366 (N_9366,N_8838,N_8395);
or U9367 (N_9367,N_8529,N_8643);
nand U9368 (N_9368,N_8268,N_8600);
nand U9369 (N_9369,N_8994,N_8538);
and U9370 (N_9370,N_8885,N_8270);
and U9371 (N_9371,N_8400,N_8399);
nor U9372 (N_9372,N_8679,N_8447);
nor U9373 (N_9373,N_8540,N_8772);
and U9374 (N_9374,N_8663,N_8515);
nor U9375 (N_9375,N_8618,N_8452);
and U9376 (N_9376,N_8322,N_8417);
nor U9377 (N_9377,N_8906,N_8388);
or U9378 (N_9378,N_8508,N_8372);
or U9379 (N_9379,N_8906,N_8796);
or U9380 (N_9380,N_8934,N_8673);
nand U9381 (N_9381,N_8738,N_8350);
nand U9382 (N_9382,N_8729,N_8322);
nor U9383 (N_9383,N_8419,N_8255);
or U9384 (N_9384,N_8726,N_8757);
nor U9385 (N_9385,N_8541,N_8658);
or U9386 (N_9386,N_8552,N_8386);
and U9387 (N_9387,N_8338,N_8259);
nor U9388 (N_9388,N_8775,N_8503);
or U9389 (N_9389,N_8822,N_8366);
and U9390 (N_9390,N_8299,N_8533);
or U9391 (N_9391,N_8952,N_8640);
or U9392 (N_9392,N_8279,N_8278);
or U9393 (N_9393,N_8380,N_8991);
nor U9394 (N_9394,N_8405,N_8719);
nor U9395 (N_9395,N_8842,N_8554);
nor U9396 (N_9396,N_8290,N_8592);
nand U9397 (N_9397,N_8373,N_8322);
nand U9398 (N_9398,N_8371,N_8721);
nor U9399 (N_9399,N_8261,N_8377);
nand U9400 (N_9400,N_8712,N_8792);
and U9401 (N_9401,N_8316,N_8928);
nand U9402 (N_9402,N_8923,N_8568);
nand U9403 (N_9403,N_8619,N_8892);
nand U9404 (N_9404,N_8475,N_8803);
nand U9405 (N_9405,N_8873,N_8802);
nand U9406 (N_9406,N_8272,N_8344);
xor U9407 (N_9407,N_8626,N_8742);
or U9408 (N_9408,N_8554,N_8303);
or U9409 (N_9409,N_8613,N_8835);
or U9410 (N_9410,N_8452,N_8523);
nor U9411 (N_9411,N_8883,N_8916);
xor U9412 (N_9412,N_8413,N_8999);
nand U9413 (N_9413,N_8991,N_8873);
xnor U9414 (N_9414,N_8507,N_8734);
nor U9415 (N_9415,N_8922,N_8510);
nor U9416 (N_9416,N_8938,N_8882);
nor U9417 (N_9417,N_8277,N_8681);
nand U9418 (N_9418,N_8738,N_8861);
nand U9419 (N_9419,N_8419,N_8314);
nor U9420 (N_9420,N_8730,N_8866);
and U9421 (N_9421,N_8311,N_8473);
and U9422 (N_9422,N_8911,N_8250);
nand U9423 (N_9423,N_8917,N_8985);
xor U9424 (N_9424,N_8796,N_8988);
nor U9425 (N_9425,N_8536,N_8720);
or U9426 (N_9426,N_8694,N_8697);
nand U9427 (N_9427,N_8562,N_8443);
and U9428 (N_9428,N_8713,N_8974);
or U9429 (N_9429,N_8602,N_8834);
and U9430 (N_9430,N_8582,N_8715);
nor U9431 (N_9431,N_8715,N_8514);
nand U9432 (N_9432,N_8802,N_8790);
nor U9433 (N_9433,N_8420,N_8264);
or U9434 (N_9434,N_8505,N_8438);
and U9435 (N_9435,N_8327,N_8335);
or U9436 (N_9436,N_8951,N_8670);
or U9437 (N_9437,N_8392,N_8484);
xor U9438 (N_9438,N_8745,N_8811);
nand U9439 (N_9439,N_8939,N_8953);
and U9440 (N_9440,N_8636,N_8648);
and U9441 (N_9441,N_8346,N_8702);
and U9442 (N_9442,N_8687,N_8606);
or U9443 (N_9443,N_8953,N_8276);
xnor U9444 (N_9444,N_8543,N_8338);
or U9445 (N_9445,N_8642,N_8699);
nor U9446 (N_9446,N_8330,N_8771);
nand U9447 (N_9447,N_8706,N_8379);
xnor U9448 (N_9448,N_8305,N_8312);
nor U9449 (N_9449,N_8384,N_8920);
nor U9450 (N_9450,N_8750,N_8736);
or U9451 (N_9451,N_8594,N_8753);
nand U9452 (N_9452,N_8410,N_8549);
or U9453 (N_9453,N_8751,N_8865);
nand U9454 (N_9454,N_8903,N_8604);
and U9455 (N_9455,N_8806,N_8616);
or U9456 (N_9456,N_8595,N_8323);
nand U9457 (N_9457,N_8460,N_8733);
and U9458 (N_9458,N_8384,N_8809);
or U9459 (N_9459,N_8371,N_8989);
nor U9460 (N_9460,N_8626,N_8275);
nand U9461 (N_9461,N_8607,N_8821);
and U9462 (N_9462,N_8587,N_8623);
nand U9463 (N_9463,N_8330,N_8890);
nand U9464 (N_9464,N_8476,N_8652);
nor U9465 (N_9465,N_8356,N_8874);
nor U9466 (N_9466,N_8654,N_8867);
nor U9467 (N_9467,N_8351,N_8799);
and U9468 (N_9468,N_8580,N_8983);
nand U9469 (N_9469,N_8275,N_8995);
nand U9470 (N_9470,N_8810,N_8369);
and U9471 (N_9471,N_8422,N_8533);
nor U9472 (N_9472,N_8291,N_8324);
and U9473 (N_9473,N_8928,N_8813);
nor U9474 (N_9474,N_8913,N_8309);
nand U9475 (N_9475,N_8599,N_8328);
nand U9476 (N_9476,N_8478,N_8493);
or U9477 (N_9477,N_8375,N_8665);
nand U9478 (N_9478,N_8615,N_8900);
nor U9479 (N_9479,N_8981,N_8980);
and U9480 (N_9480,N_8512,N_8961);
nand U9481 (N_9481,N_8810,N_8518);
xnor U9482 (N_9482,N_8472,N_8253);
nand U9483 (N_9483,N_8849,N_8810);
or U9484 (N_9484,N_8734,N_8590);
nand U9485 (N_9485,N_8643,N_8469);
xnor U9486 (N_9486,N_8426,N_8654);
or U9487 (N_9487,N_8979,N_8639);
or U9488 (N_9488,N_8562,N_8307);
and U9489 (N_9489,N_8590,N_8666);
nor U9490 (N_9490,N_8816,N_8868);
nand U9491 (N_9491,N_8724,N_8300);
nand U9492 (N_9492,N_8676,N_8833);
xnor U9493 (N_9493,N_8810,N_8659);
or U9494 (N_9494,N_8906,N_8496);
nor U9495 (N_9495,N_8596,N_8589);
and U9496 (N_9496,N_8827,N_8651);
and U9497 (N_9497,N_8992,N_8803);
and U9498 (N_9498,N_8856,N_8574);
nor U9499 (N_9499,N_8484,N_8728);
or U9500 (N_9500,N_8372,N_8919);
and U9501 (N_9501,N_8292,N_8658);
or U9502 (N_9502,N_8404,N_8692);
or U9503 (N_9503,N_8493,N_8630);
nor U9504 (N_9504,N_8541,N_8799);
nand U9505 (N_9505,N_8394,N_8767);
nor U9506 (N_9506,N_8952,N_8342);
nand U9507 (N_9507,N_8669,N_8804);
or U9508 (N_9508,N_8392,N_8687);
nor U9509 (N_9509,N_8648,N_8302);
nor U9510 (N_9510,N_8751,N_8774);
nand U9511 (N_9511,N_8681,N_8775);
or U9512 (N_9512,N_8728,N_8605);
or U9513 (N_9513,N_8480,N_8677);
nand U9514 (N_9514,N_8275,N_8321);
and U9515 (N_9515,N_8544,N_8528);
nand U9516 (N_9516,N_8900,N_8847);
nand U9517 (N_9517,N_8350,N_8352);
nand U9518 (N_9518,N_8810,N_8661);
xnor U9519 (N_9519,N_8632,N_8428);
and U9520 (N_9520,N_8827,N_8725);
xor U9521 (N_9521,N_8925,N_8544);
and U9522 (N_9522,N_8427,N_8883);
or U9523 (N_9523,N_8888,N_8859);
and U9524 (N_9524,N_8294,N_8289);
and U9525 (N_9525,N_8711,N_8844);
nand U9526 (N_9526,N_8549,N_8605);
nor U9527 (N_9527,N_8493,N_8731);
or U9528 (N_9528,N_8665,N_8493);
nor U9529 (N_9529,N_8421,N_8526);
nand U9530 (N_9530,N_8994,N_8649);
nor U9531 (N_9531,N_8911,N_8279);
nand U9532 (N_9532,N_8390,N_8760);
nand U9533 (N_9533,N_8419,N_8256);
nand U9534 (N_9534,N_8917,N_8500);
and U9535 (N_9535,N_8371,N_8666);
nor U9536 (N_9536,N_8838,N_8542);
and U9537 (N_9537,N_8476,N_8712);
nor U9538 (N_9538,N_8293,N_8360);
or U9539 (N_9539,N_8710,N_8854);
nand U9540 (N_9540,N_8992,N_8922);
nor U9541 (N_9541,N_8630,N_8398);
or U9542 (N_9542,N_8415,N_8328);
nand U9543 (N_9543,N_8921,N_8987);
and U9544 (N_9544,N_8455,N_8693);
nor U9545 (N_9545,N_8271,N_8343);
nand U9546 (N_9546,N_8413,N_8486);
and U9547 (N_9547,N_8717,N_8867);
or U9548 (N_9548,N_8610,N_8542);
and U9549 (N_9549,N_8896,N_8641);
or U9550 (N_9550,N_8490,N_8440);
nand U9551 (N_9551,N_8590,N_8826);
nand U9552 (N_9552,N_8476,N_8308);
or U9553 (N_9553,N_8323,N_8650);
and U9554 (N_9554,N_8742,N_8497);
nor U9555 (N_9555,N_8919,N_8313);
or U9556 (N_9556,N_8844,N_8825);
or U9557 (N_9557,N_8267,N_8945);
and U9558 (N_9558,N_8381,N_8921);
nor U9559 (N_9559,N_8870,N_8371);
or U9560 (N_9560,N_8669,N_8272);
or U9561 (N_9561,N_8485,N_8528);
and U9562 (N_9562,N_8650,N_8557);
and U9563 (N_9563,N_8964,N_8510);
nor U9564 (N_9564,N_8640,N_8833);
and U9565 (N_9565,N_8713,N_8819);
and U9566 (N_9566,N_8914,N_8693);
or U9567 (N_9567,N_8362,N_8416);
and U9568 (N_9568,N_8536,N_8873);
nand U9569 (N_9569,N_8680,N_8687);
and U9570 (N_9570,N_8691,N_8487);
and U9571 (N_9571,N_8754,N_8921);
and U9572 (N_9572,N_8381,N_8608);
or U9573 (N_9573,N_8871,N_8457);
nand U9574 (N_9574,N_8735,N_8354);
xnor U9575 (N_9575,N_8774,N_8933);
nand U9576 (N_9576,N_8737,N_8476);
nor U9577 (N_9577,N_8604,N_8940);
or U9578 (N_9578,N_8662,N_8754);
nor U9579 (N_9579,N_8920,N_8393);
or U9580 (N_9580,N_8278,N_8443);
or U9581 (N_9581,N_8955,N_8755);
and U9582 (N_9582,N_8396,N_8750);
and U9583 (N_9583,N_8256,N_8603);
nand U9584 (N_9584,N_8813,N_8880);
and U9585 (N_9585,N_8498,N_8527);
and U9586 (N_9586,N_8841,N_8466);
and U9587 (N_9587,N_8444,N_8901);
or U9588 (N_9588,N_8706,N_8664);
nand U9589 (N_9589,N_8721,N_8627);
xor U9590 (N_9590,N_8579,N_8417);
nand U9591 (N_9591,N_8434,N_8836);
nor U9592 (N_9592,N_8727,N_8795);
and U9593 (N_9593,N_8999,N_8377);
or U9594 (N_9594,N_8538,N_8612);
nor U9595 (N_9595,N_8771,N_8624);
or U9596 (N_9596,N_8461,N_8251);
nor U9597 (N_9597,N_8662,N_8518);
or U9598 (N_9598,N_8885,N_8333);
nor U9599 (N_9599,N_8303,N_8519);
nand U9600 (N_9600,N_8954,N_8969);
or U9601 (N_9601,N_8768,N_8779);
nor U9602 (N_9602,N_8892,N_8530);
nor U9603 (N_9603,N_8776,N_8589);
nand U9604 (N_9604,N_8707,N_8515);
or U9605 (N_9605,N_8370,N_8646);
nand U9606 (N_9606,N_8460,N_8657);
nor U9607 (N_9607,N_8929,N_8713);
or U9608 (N_9608,N_8351,N_8800);
nor U9609 (N_9609,N_8402,N_8429);
nand U9610 (N_9610,N_8824,N_8348);
or U9611 (N_9611,N_8297,N_8700);
nor U9612 (N_9612,N_8691,N_8679);
nand U9613 (N_9613,N_8793,N_8268);
and U9614 (N_9614,N_8412,N_8929);
and U9615 (N_9615,N_8744,N_8448);
xor U9616 (N_9616,N_8520,N_8736);
nor U9617 (N_9617,N_8482,N_8543);
nand U9618 (N_9618,N_8804,N_8321);
xnor U9619 (N_9619,N_8790,N_8654);
nor U9620 (N_9620,N_8818,N_8585);
nand U9621 (N_9621,N_8624,N_8493);
or U9622 (N_9622,N_8662,N_8549);
and U9623 (N_9623,N_8255,N_8862);
and U9624 (N_9624,N_8272,N_8828);
and U9625 (N_9625,N_8563,N_8429);
nand U9626 (N_9626,N_8364,N_8745);
or U9627 (N_9627,N_8703,N_8783);
xnor U9628 (N_9628,N_8752,N_8647);
or U9629 (N_9629,N_8447,N_8817);
or U9630 (N_9630,N_8972,N_8925);
and U9631 (N_9631,N_8866,N_8681);
nor U9632 (N_9632,N_8366,N_8865);
or U9633 (N_9633,N_8758,N_8879);
nand U9634 (N_9634,N_8762,N_8356);
xnor U9635 (N_9635,N_8491,N_8420);
and U9636 (N_9636,N_8768,N_8691);
or U9637 (N_9637,N_8445,N_8411);
nor U9638 (N_9638,N_8369,N_8263);
or U9639 (N_9639,N_8934,N_8527);
and U9640 (N_9640,N_8391,N_8379);
nor U9641 (N_9641,N_8428,N_8303);
or U9642 (N_9642,N_8369,N_8953);
xnor U9643 (N_9643,N_8420,N_8998);
and U9644 (N_9644,N_8678,N_8618);
or U9645 (N_9645,N_8279,N_8268);
nor U9646 (N_9646,N_8430,N_8959);
xnor U9647 (N_9647,N_8971,N_8660);
nor U9648 (N_9648,N_8258,N_8536);
and U9649 (N_9649,N_8823,N_8427);
nand U9650 (N_9650,N_8659,N_8615);
and U9651 (N_9651,N_8967,N_8835);
nand U9652 (N_9652,N_8857,N_8595);
or U9653 (N_9653,N_8862,N_8938);
or U9654 (N_9654,N_8944,N_8470);
nor U9655 (N_9655,N_8315,N_8289);
and U9656 (N_9656,N_8333,N_8478);
nand U9657 (N_9657,N_8946,N_8587);
or U9658 (N_9658,N_8913,N_8663);
xnor U9659 (N_9659,N_8287,N_8819);
nor U9660 (N_9660,N_8920,N_8970);
or U9661 (N_9661,N_8649,N_8664);
xor U9662 (N_9662,N_8554,N_8851);
nand U9663 (N_9663,N_8881,N_8288);
and U9664 (N_9664,N_8793,N_8878);
xnor U9665 (N_9665,N_8617,N_8628);
nor U9666 (N_9666,N_8803,N_8855);
and U9667 (N_9667,N_8795,N_8712);
nand U9668 (N_9668,N_8450,N_8770);
or U9669 (N_9669,N_8870,N_8949);
or U9670 (N_9670,N_8928,N_8680);
nand U9671 (N_9671,N_8760,N_8777);
xnor U9672 (N_9672,N_8290,N_8628);
and U9673 (N_9673,N_8399,N_8733);
or U9674 (N_9674,N_8643,N_8551);
and U9675 (N_9675,N_8270,N_8259);
nor U9676 (N_9676,N_8457,N_8579);
nor U9677 (N_9677,N_8296,N_8829);
nor U9678 (N_9678,N_8301,N_8456);
nor U9679 (N_9679,N_8830,N_8593);
nor U9680 (N_9680,N_8723,N_8573);
nor U9681 (N_9681,N_8760,N_8683);
nor U9682 (N_9682,N_8875,N_8998);
and U9683 (N_9683,N_8780,N_8352);
or U9684 (N_9684,N_8500,N_8604);
nor U9685 (N_9685,N_8473,N_8413);
xor U9686 (N_9686,N_8793,N_8836);
or U9687 (N_9687,N_8436,N_8489);
nand U9688 (N_9688,N_8882,N_8551);
nand U9689 (N_9689,N_8505,N_8627);
nor U9690 (N_9690,N_8440,N_8937);
and U9691 (N_9691,N_8975,N_8792);
nor U9692 (N_9692,N_8498,N_8974);
or U9693 (N_9693,N_8384,N_8893);
or U9694 (N_9694,N_8620,N_8967);
nor U9695 (N_9695,N_8901,N_8551);
or U9696 (N_9696,N_8807,N_8446);
xnor U9697 (N_9697,N_8377,N_8651);
nor U9698 (N_9698,N_8288,N_8393);
nand U9699 (N_9699,N_8669,N_8749);
nand U9700 (N_9700,N_8659,N_8686);
nor U9701 (N_9701,N_8858,N_8921);
or U9702 (N_9702,N_8883,N_8260);
or U9703 (N_9703,N_8549,N_8381);
nand U9704 (N_9704,N_8737,N_8758);
nor U9705 (N_9705,N_8746,N_8951);
and U9706 (N_9706,N_8301,N_8504);
nand U9707 (N_9707,N_8757,N_8728);
nor U9708 (N_9708,N_8636,N_8633);
nor U9709 (N_9709,N_8757,N_8714);
or U9710 (N_9710,N_8268,N_8721);
nand U9711 (N_9711,N_8846,N_8576);
nor U9712 (N_9712,N_8738,N_8419);
nand U9713 (N_9713,N_8822,N_8575);
nor U9714 (N_9714,N_8432,N_8485);
nor U9715 (N_9715,N_8317,N_8280);
nand U9716 (N_9716,N_8314,N_8554);
nand U9717 (N_9717,N_8774,N_8931);
nor U9718 (N_9718,N_8381,N_8981);
nand U9719 (N_9719,N_8972,N_8380);
nor U9720 (N_9720,N_8272,N_8452);
or U9721 (N_9721,N_8581,N_8483);
or U9722 (N_9722,N_8424,N_8519);
and U9723 (N_9723,N_8853,N_8711);
and U9724 (N_9724,N_8868,N_8322);
and U9725 (N_9725,N_8986,N_8335);
nor U9726 (N_9726,N_8341,N_8781);
and U9727 (N_9727,N_8925,N_8292);
nand U9728 (N_9728,N_8953,N_8887);
or U9729 (N_9729,N_8853,N_8945);
xnor U9730 (N_9730,N_8925,N_8662);
and U9731 (N_9731,N_8556,N_8575);
xor U9732 (N_9732,N_8829,N_8772);
xnor U9733 (N_9733,N_8474,N_8950);
nand U9734 (N_9734,N_8282,N_8551);
nor U9735 (N_9735,N_8836,N_8364);
and U9736 (N_9736,N_8283,N_8499);
nand U9737 (N_9737,N_8899,N_8567);
or U9738 (N_9738,N_8420,N_8301);
xor U9739 (N_9739,N_8483,N_8836);
and U9740 (N_9740,N_8298,N_8727);
and U9741 (N_9741,N_8323,N_8443);
nand U9742 (N_9742,N_8814,N_8345);
or U9743 (N_9743,N_8924,N_8718);
nor U9744 (N_9744,N_8669,N_8511);
or U9745 (N_9745,N_8260,N_8961);
and U9746 (N_9746,N_8391,N_8633);
nor U9747 (N_9747,N_8888,N_8597);
nor U9748 (N_9748,N_8950,N_8907);
or U9749 (N_9749,N_8346,N_8904);
or U9750 (N_9750,N_9173,N_9377);
nor U9751 (N_9751,N_9300,N_9220);
nand U9752 (N_9752,N_9000,N_9559);
nor U9753 (N_9753,N_9064,N_9349);
or U9754 (N_9754,N_9495,N_9638);
nor U9755 (N_9755,N_9091,N_9146);
nor U9756 (N_9756,N_9383,N_9303);
and U9757 (N_9757,N_9264,N_9746);
or U9758 (N_9758,N_9347,N_9435);
nor U9759 (N_9759,N_9253,N_9658);
or U9760 (N_9760,N_9351,N_9359);
nor U9761 (N_9761,N_9193,N_9293);
nand U9762 (N_9762,N_9339,N_9013);
nand U9763 (N_9763,N_9572,N_9677);
or U9764 (N_9764,N_9528,N_9421);
or U9765 (N_9765,N_9427,N_9222);
and U9766 (N_9766,N_9657,N_9499);
or U9767 (N_9767,N_9289,N_9231);
and U9768 (N_9768,N_9578,N_9602);
nor U9769 (N_9769,N_9471,N_9233);
nand U9770 (N_9770,N_9115,N_9162);
or U9771 (N_9771,N_9319,N_9729);
xnor U9772 (N_9772,N_9441,N_9726);
nor U9773 (N_9773,N_9371,N_9203);
nand U9774 (N_9774,N_9611,N_9036);
nand U9775 (N_9775,N_9154,N_9294);
and U9776 (N_9776,N_9413,N_9338);
nand U9777 (N_9777,N_9334,N_9095);
and U9778 (N_9778,N_9663,N_9044);
or U9779 (N_9779,N_9312,N_9191);
nor U9780 (N_9780,N_9344,N_9260);
or U9781 (N_9781,N_9695,N_9641);
nor U9782 (N_9782,N_9702,N_9135);
or U9783 (N_9783,N_9667,N_9336);
xor U9784 (N_9784,N_9144,N_9608);
or U9785 (N_9785,N_9448,N_9309);
and U9786 (N_9786,N_9538,N_9556);
and U9787 (N_9787,N_9614,N_9567);
or U9788 (N_9788,N_9683,N_9454);
and U9789 (N_9789,N_9600,N_9105);
nand U9790 (N_9790,N_9106,N_9092);
or U9791 (N_9791,N_9076,N_9698);
and U9792 (N_9792,N_9073,N_9432);
nor U9793 (N_9793,N_9691,N_9739);
and U9794 (N_9794,N_9420,N_9587);
nand U9795 (N_9795,N_9021,N_9205);
and U9796 (N_9796,N_9403,N_9425);
or U9797 (N_9797,N_9711,N_9131);
or U9798 (N_9798,N_9207,N_9439);
nor U9799 (N_9799,N_9047,N_9270);
or U9800 (N_9800,N_9062,N_9706);
or U9801 (N_9801,N_9554,N_9428);
nand U9802 (N_9802,N_9056,N_9626);
or U9803 (N_9803,N_9455,N_9615);
or U9804 (N_9804,N_9510,N_9089);
nor U9805 (N_9805,N_9249,N_9533);
and U9806 (N_9806,N_9248,N_9715);
or U9807 (N_9807,N_9335,N_9268);
and U9808 (N_9808,N_9027,N_9444);
nand U9809 (N_9809,N_9734,N_9265);
nand U9810 (N_9810,N_9684,N_9124);
nand U9811 (N_9811,N_9310,N_9450);
or U9812 (N_9812,N_9133,N_9058);
nor U9813 (N_9813,N_9186,N_9386);
and U9814 (N_9814,N_9185,N_9316);
nor U9815 (N_9815,N_9718,N_9355);
or U9816 (N_9816,N_9125,N_9071);
or U9817 (N_9817,N_9380,N_9748);
or U9818 (N_9818,N_9550,N_9093);
nor U9819 (N_9819,N_9422,N_9009);
nand U9820 (N_9820,N_9498,N_9308);
nand U9821 (N_9821,N_9030,N_9041);
and U9822 (N_9822,N_9070,N_9415);
and U9823 (N_9823,N_9512,N_9055);
nor U9824 (N_9824,N_9743,N_9668);
nand U9825 (N_9825,N_9731,N_9632);
xor U9826 (N_9826,N_9522,N_9273);
xnor U9827 (N_9827,N_9018,N_9118);
or U9828 (N_9828,N_9639,N_9674);
nor U9829 (N_9829,N_9470,N_9278);
and U9830 (N_9830,N_9145,N_9513);
nand U9831 (N_9831,N_9098,N_9024);
or U9832 (N_9832,N_9543,N_9122);
and U9833 (N_9833,N_9612,N_9040);
nor U9834 (N_9834,N_9490,N_9321);
nand U9835 (N_9835,N_9414,N_9214);
or U9836 (N_9836,N_9419,N_9655);
or U9837 (N_9837,N_9652,N_9127);
nor U9838 (N_9838,N_9103,N_9085);
xnor U9839 (N_9839,N_9688,N_9182);
nand U9840 (N_9840,N_9408,N_9477);
and U9841 (N_9841,N_9671,N_9116);
xor U9842 (N_9842,N_9317,N_9583);
or U9843 (N_9843,N_9094,N_9447);
xnor U9844 (N_9844,N_9057,N_9437);
and U9845 (N_9845,N_9476,N_9467);
or U9846 (N_9846,N_9560,N_9195);
or U9847 (N_9847,N_9694,N_9650);
or U9848 (N_9848,N_9519,N_9496);
and U9849 (N_9849,N_9117,N_9281);
nor U9850 (N_9850,N_9245,N_9722);
nor U9851 (N_9851,N_9177,N_9374);
nand U9852 (N_9852,N_9610,N_9465);
and U9853 (N_9853,N_9460,N_9217);
nand U9854 (N_9854,N_9163,N_9518);
and U9855 (N_9855,N_9553,N_9216);
nand U9856 (N_9856,N_9693,N_9251);
nor U9857 (N_9857,N_9372,N_9540);
and U9858 (N_9858,N_9341,N_9120);
nor U9859 (N_9859,N_9107,N_9311);
nand U9860 (N_9860,N_9628,N_9523);
nand U9861 (N_9861,N_9179,N_9088);
and U9862 (N_9862,N_9302,N_9576);
nand U9863 (N_9863,N_9114,N_9497);
nand U9864 (N_9864,N_9033,N_9174);
or U9865 (N_9865,N_9406,N_9430);
nor U9866 (N_9866,N_9016,N_9011);
and U9867 (N_9867,N_9581,N_9378);
xnor U9868 (N_9868,N_9325,N_9384);
or U9869 (N_9869,N_9619,N_9330);
or U9870 (N_9870,N_9015,N_9020);
xnor U9871 (N_9871,N_9599,N_9156);
and U9872 (N_9872,N_9633,N_9171);
or U9873 (N_9873,N_9346,N_9048);
nor U9874 (N_9874,N_9473,N_9049);
nor U9875 (N_9875,N_9043,N_9679);
nor U9876 (N_9876,N_9417,N_9243);
nor U9877 (N_9877,N_9622,N_9364);
and U9878 (N_9878,N_9666,N_9261);
nor U9879 (N_9879,N_9515,N_9449);
nor U9880 (N_9880,N_9431,N_9531);
nor U9881 (N_9881,N_9482,N_9200);
nand U9882 (N_9882,N_9597,N_9365);
nor U9883 (N_9883,N_9204,N_9451);
nand U9884 (N_9884,N_9389,N_9227);
nand U9885 (N_9885,N_9680,N_9104);
and U9886 (N_9886,N_9687,N_9485);
nor U9887 (N_9887,N_9291,N_9479);
nand U9888 (N_9888,N_9078,N_9022);
nor U9889 (N_9889,N_9646,N_9535);
and U9890 (N_9890,N_9290,N_9164);
nand U9891 (N_9891,N_9255,N_9254);
nand U9892 (N_9892,N_9516,N_9401);
xor U9893 (N_9893,N_9287,N_9388);
and U9894 (N_9894,N_9382,N_9053);
nor U9895 (N_9895,N_9202,N_9356);
xor U9896 (N_9896,N_9661,N_9409);
or U9897 (N_9897,N_9724,N_9052);
nand U9898 (N_9898,N_9669,N_9213);
or U9899 (N_9899,N_9352,N_9433);
xor U9900 (N_9900,N_9343,N_9462);
nor U9901 (N_9901,N_9398,N_9225);
nor U9902 (N_9902,N_9354,N_9461);
and U9903 (N_9903,N_9474,N_9358);
nand U9904 (N_9904,N_9604,N_9399);
nand U9905 (N_9905,N_9712,N_9244);
and U9906 (N_9906,N_9142,N_9566);
and U9907 (N_9907,N_9224,N_9525);
xnor U9908 (N_9908,N_9673,N_9703);
nor U9909 (N_9909,N_9579,N_9267);
nand U9910 (N_9910,N_9488,N_9670);
nor U9911 (N_9911,N_9035,N_9370);
or U9912 (N_9912,N_9453,N_9042);
nand U9913 (N_9913,N_9178,N_9545);
nor U9914 (N_9914,N_9002,N_9140);
and U9915 (N_9915,N_9304,N_9423);
nand U9916 (N_9916,N_9003,N_9594);
nor U9917 (N_9917,N_9521,N_9109);
nand U9918 (N_9918,N_9363,N_9621);
nor U9919 (N_9919,N_9169,N_9170);
xor U9920 (N_9920,N_9369,N_9494);
nor U9921 (N_9921,N_9740,N_9054);
xor U9922 (N_9922,N_9134,N_9315);
nor U9923 (N_9923,N_9649,N_9714);
and U9924 (N_9924,N_9299,N_9084);
or U9925 (N_9925,N_9440,N_9110);
xor U9926 (N_9926,N_9152,N_9457);
xor U9927 (N_9927,N_9590,N_9735);
nor U9928 (N_9928,N_9692,N_9544);
nor U9929 (N_9929,N_9723,N_9645);
and U9930 (N_9930,N_9180,N_9573);
and U9931 (N_9931,N_9329,N_9727);
or U9932 (N_9932,N_9716,N_9150);
nand U9933 (N_9933,N_9277,N_9353);
and U9934 (N_9934,N_9250,N_9198);
and U9935 (N_9935,N_9640,N_9491);
or U9936 (N_9936,N_9699,N_9407);
and U9937 (N_9937,N_9068,N_9357);
and U9938 (N_9938,N_9238,N_9029);
and U9939 (N_9939,N_9236,N_9242);
nor U9940 (N_9940,N_9630,N_9493);
and U9941 (N_9941,N_9627,N_9274);
and U9942 (N_9942,N_9552,N_9502);
nor U9943 (N_9943,N_9006,N_9379);
nand U9944 (N_9944,N_9527,N_9736);
nor U9945 (N_9945,N_9503,N_9588);
nand U9946 (N_9946,N_9537,N_9160);
and U9947 (N_9947,N_9279,N_9396);
nor U9948 (N_9948,N_9223,N_9445);
and U9949 (N_9949,N_9138,N_9209);
and U9950 (N_9950,N_9007,N_9241);
nor U9951 (N_9951,N_9368,N_9631);
xnor U9952 (N_9952,N_9136,N_9429);
and U9953 (N_9953,N_9411,N_9713);
xnor U9954 (N_9954,N_9466,N_9045);
or U9955 (N_9955,N_9201,N_9592);
or U9956 (N_9956,N_9732,N_9340);
xor U9957 (N_9957,N_9305,N_9288);
nand U9958 (N_9958,N_9475,N_9557);
nand U9959 (N_9959,N_9017,N_9524);
xnor U9960 (N_9960,N_9464,N_9327);
and U9961 (N_9961,N_9613,N_9511);
nor U9962 (N_9962,N_9656,N_9285);
nand U9963 (N_9963,N_9720,N_9326);
xnor U9964 (N_9964,N_9151,N_9301);
xor U9965 (N_9965,N_9585,N_9446);
nand U9966 (N_9966,N_9280,N_9155);
or U9967 (N_9967,N_9039,N_9292);
and U9968 (N_9968,N_9031,N_9741);
and U9969 (N_9969,N_9616,N_9589);
nand U9970 (N_9970,N_9595,N_9660);
and U9971 (N_9971,N_9549,N_9607);
or U9972 (N_9972,N_9617,N_9634);
nor U9973 (N_9973,N_9168,N_9458);
or U9974 (N_9974,N_9230,N_9418);
xnor U9975 (N_9975,N_9542,N_9012);
nor U9976 (N_9976,N_9059,N_9306);
or U9977 (N_9977,N_9086,N_9487);
or U9978 (N_9978,N_9728,N_9143);
or U9979 (N_9979,N_9392,N_9102);
and U9980 (N_9980,N_9130,N_9591);
or U9981 (N_9981,N_9077,N_9175);
xor U9982 (N_9982,N_9023,N_9412);
and U9983 (N_9983,N_9307,N_9097);
nand U9984 (N_9984,N_9189,N_9362);
nand U9985 (N_9985,N_9529,N_9436);
nand U9986 (N_9986,N_9026,N_9569);
or U9987 (N_9987,N_9108,N_9069);
nor U9988 (N_9988,N_9397,N_9025);
and U9989 (N_9989,N_9681,N_9580);
and U9990 (N_9990,N_9037,N_9424);
or U9991 (N_9991,N_9625,N_9212);
and U9992 (N_9992,N_9060,N_9258);
or U9993 (N_9993,N_9618,N_9119);
nor U9994 (N_9994,N_9096,N_9113);
nor U9995 (N_9995,N_9210,N_9153);
xnor U9996 (N_9996,N_9443,N_9367);
and U9997 (N_9997,N_9211,N_9416);
or U9998 (N_9998,N_9624,N_9456);
nand U9999 (N_9999,N_9452,N_9067);
and U10000 (N_10000,N_9080,N_9501);
nor U10001 (N_10001,N_9532,N_9232);
nor U10002 (N_10002,N_9161,N_9558);
nand U10003 (N_10003,N_9034,N_9066);
and U10004 (N_10004,N_9682,N_9514);
nand U10005 (N_10005,N_9707,N_9208);
or U10006 (N_10006,N_9390,N_9276);
or U10007 (N_10007,N_9239,N_9609);
nand U10008 (N_10008,N_9314,N_9324);
nand U10009 (N_10009,N_9313,N_9157);
or U10010 (N_10010,N_9745,N_9259);
nor U10011 (N_10011,N_9653,N_9730);
or U10012 (N_10012,N_9642,N_9165);
or U10013 (N_10013,N_9187,N_9263);
nand U10014 (N_10014,N_9075,N_9196);
nand U10015 (N_10015,N_9361,N_9697);
nand U10016 (N_10016,N_9240,N_9690);
xnor U10017 (N_10017,N_9530,N_9019);
nor U10018 (N_10018,N_9266,N_9584);
or U10019 (N_10019,N_9500,N_9749);
and U10020 (N_10020,N_9489,N_9298);
nand U10021 (N_10021,N_9717,N_9262);
nor U10022 (N_10022,N_9342,N_9644);
nor U10023 (N_10023,N_9541,N_9381);
nor U10024 (N_10024,N_9438,N_9664);
nor U10025 (N_10025,N_9742,N_9079);
and U10026 (N_10026,N_9141,N_9551);
or U10027 (N_10027,N_9637,N_9710);
nor U10028 (N_10028,N_9275,N_9725);
or U10029 (N_10029,N_9074,N_9562);
and U10030 (N_10030,N_9010,N_9662);
nand U10031 (N_10031,N_9139,N_9705);
and U10032 (N_10032,N_9520,N_9283);
nor U10033 (N_10033,N_9148,N_9629);
nor U10034 (N_10034,N_9555,N_9721);
xnor U10035 (N_10035,N_9719,N_9738);
nor U10036 (N_10036,N_9366,N_9028);
nand U10037 (N_10037,N_9385,N_9123);
or U10038 (N_10038,N_9546,N_9219);
or U10039 (N_10039,N_9272,N_9598);
and U10040 (N_10040,N_9159,N_9190);
nor U10041 (N_10041,N_9051,N_9484);
nand U10042 (N_10042,N_9506,N_9147);
nand U10043 (N_10043,N_9137,N_9747);
and U10044 (N_10044,N_9257,N_9676);
and U10045 (N_10045,N_9636,N_9271);
and U10046 (N_10046,N_9582,N_9647);
nor U10047 (N_10047,N_9623,N_9508);
and U10048 (N_10048,N_9686,N_9574);
or U10049 (N_10049,N_9606,N_9737);
xor U10050 (N_10050,N_9228,N_9593);
or U10051 (N_10051,N_9704,N_9548);
and U10052 (N_10052,N_9696,N_9038);
nor U10053 (N_10053,N_9247,N_9256);
nand U10054 (N_10054,N_9675,N_9348);
or U10055 (N_10055,N_9387,N_9149);
and U10056 (N_10056,N_9395,N_9082);
and U10057 (N_10057,N_9100,N_9376);
xor U10058 (N_10058,N_9481,N_9733);
xnor U10059 (N_10059,N_9472,N_9337);
and U10060 (N_10060,N_9001,N_9605);
or U10061 (N_10061,N_9563,N_9492);
or U10062 (N_10062,N_9375,N_9099);
nand U10063 (N_10063,N_9284,N_9601);
nand U10064 (N_10064,N_9183,N_9394);
or U10065 (N_10065,N_9121,N_9536);
nor U10066 (N_10066,N_9282,N_9286);
and U10067 (N_10067,N_9539,N_9570);
or U10068 (N_10068,N_9700,N_9126);
or U10069 (N_10069,N_9603,N_9206);
nand U10070 (N_10070,N_9129,N_9246);
nor U10071 (N_10071,N_9651,N_9320);
nand U10072 (N_10072,N_9547,N_9065);
or U10073 (N_10073,N_9237,N_9063);
nor U10074 (N_10074,N_9643,N_9654);
and U10075 (N_10075,N_9192,N_9295);
nand U10076 (N_10076,N_9504,N_9507);
or U10077 (N_10077,N_9072,N_9400);
and U10078 (N_10078,N_9410,N_9005);
nand U10079 (N_10079,N_9328,N_9360);
xor U10080 (N_10080,N_9032,N_9561);
and U10081 (N_10081,N_9486,N_9322);
nand U10082 (N_10082,N_9434,N_9061);
nor U10083 (N_10083,N_9402,N_9333);
nor U10084 (N_10084,N_9083,N_9226);
xor U10085 (N_10085,N_9564,N_9442);
nor U10086 (N_10086,N_9701,N_9483);
nor U10087 (N_10087,N_9744,N_9469);
xnor U10088 (N_10088,N_9586,N_9391);
nor U10089 (N_10089,N_9459,N_9112);
or U10090 (N_10090,N_9234,N_9081);
nand U10091 (N_10091,N_9111,N_9517);
and U10092 (N_10092,N_9405,N_9577);
or U10093 (N_10093,N_9331,N_9565);
or U10094 (N_10094,N_9158,N_9046);
nand U10095 (N_10095,N_9708,N_9393);
and U10096 (N_10096,N_9635,N_9087);
and U10097 (N_10097,N_9101,N_9184);
and U10098 (N_10098,N_9332,N_9199);
or U10099 (N_10099,N_9620,N_9176);
nor U10100 (N_10100,N_9181,N_9685);
nand U10101 (N_10101,N_9665,N_9345);
and U10102 (N_10102,N_9571,N_9128);
nand U10103 (N_10103,N_9188,N_9008);
xnor U10104 (N_10104,N_9004,N_9172);
and U10105 (N_10105,N_9672,N_9709);
nand U10106 (N_10106,N_9648,N_9166);
or U10107 (N_10107,N_9468,N_9132);
and U10108 (N_10108,N_9480,N_9050);
and U10109 (N_10109,N_9534,N_9318);
or U10110 (N_10110,N_9252,N_9194);
or U10111 (N_10111,N_9297,N_9463);
xnor U10112 (N_10112,N_9426,N_9090);
nor U10113 (N_10113,N_9678,N_9659);
and U10114 (N_10114,N_9215,N_9229);
nand U10115 (N_10115,N_9218,N_9596);
xor U10116 (N_10116,N_9323,N_9014);
nand U10117 (N_10117,N_9197,N_9373);
xor U10118 (N_10118,N_9296,N_9568);
nand U10119 (N_10119,N_9350,N_9509);
nor U10120 (N_10120,N_9505,N_9221);
nand U10121 (N_10121,N_9575,N_9526);
or U10122 (N_10122,N_9478,N_9404);
nor U10123 (N_10123,N_9167,N_9269);
and U10124 (N_10124,N_9689,N_9235);
or U10125 (N_10125,N_9607,N_9072);
nor U10126 (N_10126,N_9702,N_9082);
or U10127 (N_10127,N_9228,N_9710);
xor U10128 (N_10128,N_9415,N_9565);
xor U10129 (N_10129,N_9033,N_9426);
or U10130 (N_10130,N_9502,N_9205);
and U10131 (N_10131,N_9065,N_9219);
xor U10132 (N_10132,N_9271,N_9238);
or U10133 (N_10133,N_9342,N_9102);
xnor U10134 (N_10134,N_9265,N_9547);
xor U10135 (N_10135,N_9109,N_9185);
nor U10136 (N_10136,N_9296,N_9584);
xor U10137 (N_10137,N_9518,N_9070);
or U10138 (N_10138,N_9446,N_9619);
or U10139 (N_10139,N_9276,N_9039);
and U10140 (N_10140,N_9373,N_9417);
and U10141 (N_10141,N_9228,N_9655);
xor U10142 (N_10142,N_9545,N_9407);
and U10143 (N_10143,N_9274,N_9315);
and U10144 (N_10144,N_9654,N_9621);
and U10145 (N_10145,N_9642,N_9370);
nor U10146 (N_10146,N_9336,N_9483);
or U10147 (N_10147,N_9685,N_9275);
and U10148 (N_10148,N_9114,N_9300);
or U10149 (N_10149,N_9363,N_9216);
and U10150 (N_10150,N_9475,N_9053);
and U10151 (N_10151,N_9322,N_9733);
nor U10152 (N_10152,N_9721,N_9342);
or U10153 (N_10153,N_9498,N_9627);
xnor U10154 (N_10154,N_9713,N_9532);
nand U10155 (N_10155,N_9694,N_9209);
or U10156 (N_10156,N_9099,N_9482);
nand U10157 (N_10157,N_9141,N_9572);
or U10158 (N_10158,N_9599,N_9532);
and U10159 (N_10159,N_9195,N_9480);
nor U10160 (N_10160,N_9507,N_9595);
and U10161 (N_10161,N_9096,N_9014);
or U10162 (N_10162,N_9266,N_9657);
nand U10163 (N_10163,N_9096,N_9118);
nor U10164 (N_10164,N_9255,N_9113);
xnor U10165 (N_10165,N_9658,N_9323);
xor U10166 (N_10166,N_9108,N_9055);
nor U10167 (N_10167,N_9319,N_9746);
xnor U10168 (N_10168,N_9086,N_9174);
or U10169 (N_10169,N_9340,N_9611);
nor U10170 (N_10170,N_9125,N_9669);
and U10171 (N_10171,N_9745,N_9103);
and U10172 (N_10172,N_9524,N_9424);
nand U10173 (N_10173,N_9727,N_9280);
or U10174 (N_10174,N_9524,N_9729);
and U10175 (N_10175,N_9524,N_9364);
nor U10176 (N_10176,N_9214,N_9074);
nand U10177 (N_10177,N_9660,N_9540);
nor U10178 (N_10178,N_9454,N_9541);
nand U10179 (N_10179,N_9065,N_9236);
nor U10180 (N_10180,N_9369,N_9382);
or U10181 (N_10181,N_9334,N_9405);
nor U10182 (N_10182,N_9623,N_9090);
or U10183 (N_10183,N_9320,N_9359);
nor U10184 (N_10184,N_9380,N_9728);
nand U10185 (N_10185,N_9600,N_9610);
nor U10186 (N_10186,N_9310,N_9026);
xor U10187 (N_10187,N_9729,N_9666);
nor U10188 (N_10188,N_9314,N_9447);
or U10189 (N_10189,N_9685,N_9043);
nand U10190 (N_10190,N_9593,N_9743);
nand U10191 (N_10191,N_9372,N_9169);
nand U10192 (N_10192,N_9026,N_9614);
nand U10193 (N_10193,N_9321,N_9364);
nand U10194 (N_10194,N_9711,N_9283);
nor U10195 (N_10195,N_9747,N_9680);
or U10196 (N_10196,N_9096,N_9493);
xor U10197 (N_10197,N_9312,N_9109);
nor U10198 (N_10198,N_9243,N_9461);
or U10199 (N_10199,N_9472,N_9140);
or U10200 (N_10200,N_9499,N_9279);
nand U10201 (N_10201,N_9228,N_9459);
nand U10202 (N_10202,N_9038,N_9487);
nand U10203 (N_10203,N_9401,N_9378);
or U10204 (N_10204,N_9437,N_9386);
nand U10205 (N_10205,N_9445,N_9135);
nand U10206 (N_10206,N_9614,N_9113);
nor U10207 (N_10207,N_9574,N_9012);
and U10208 (N_10208,N_9682,N_9395);
nor U10209 (N_10209,N_9419,N_9718);
nand U10210 (N_10210,N_9646,N_9427);
nor U10211 (N_10211,N_9016,N_9667);
and U10212 (N_10212,N_9291,N_9091);
nand U10213 (N_10213,N_9624,N_9501);
nand U10214 (N_10214,N_9402,N_9583);
nand U10215 (N_10215,N_9436,N_9581);
or U10216 (N_10216,N_9325,N_9475);
nor U10217 (N_10217,N_9338,N_9309);
nand U10218 (N_10218,N_9175,N_9608);
nor U10219 (N_10219,N_9426,N_9427);
nand U10220 (N_10220,N_9029,N_9374);
or U10221 (N_10221,N_9339,N_9489);
and U10222 (N_10222,N_9521,N_9375);
and U10223 (N_10223,N_9048,N_9291);
nor U10224 (N_10224,N_9569,N_9642);
and U10225 (N_10225,N_9608,N_9294);
and U10226 (N_10226,N_9705,N_9723);
nor U10227 (N_10227,N_9477,N_9247);
or U10228 (N_10228,N_9311,N_9628);
nand U10229 (N_10229,N_9028,N_9614);
nand U10230 (N_10230,N_9669,N_9580);
and U10231 (N_10231,N_9517,N_9080);
or U10232 (N_10232,N_9396,N_9607);
or U10233 (N_10233,N_9314,N_9113);
nand U10234 (N_10234,N_9591,N_9104);
and U10235 (N_10235,N_9522,N_9064);
or U10236 (N_10236,N_9548,N_9226);
nor U10237 (N_10237,N_9208,N_9571);
nor U10238 (N_10238,N_9677,N_9280);
nand U10239 (N_10239,N_9007,N_9350);
and U10240 (N_10240,N_9159,N_9474);
and U10241 (N_10241,N_9211,N_9663);
nand U10242 (N_10242,N_9429,N_9300);
or U10243 (N_10243,N_9531,N_9080);
xnor U10244 (N_10244,N_9565,N_9156);
or U10245 (N_10245,N_9538,N_9537);
nand U10246 (N_10246,N_9300,N_9336);
and U10247 (N_10247,N_9659,N_9666);
nor U10248 (N_10248,N_9741,N_9076);
nand U10249 (N_10249,N_9663,N_9241);
xnor U10250 (N_10250,N_9536,N_9395);
or U10251 (N_10251,N_9010,N_9535);
nor U10252 (N_10252,N_9431,N_9258);
nor U10253 (N_10253,N_9238,N_9393);
or U10254 (N_10254,N_9336,N_9205);
nor U10255 (N_10255,N_9366,N_9141);
nor U10256 (N_10256,N_9510,N_9291);
nor U10257 (N_10257,N_9003,N_9547);
or U10258 (N_10258,N_9644,N_9119);
nor U10259 (N_10259,N_9231,N_9115);
xor U10260 (N_10260,N_9247,N_9677);
and U10261 (N_10261,N_9739,N_9280);
and U10262 (N_10262,N_9602,N_9049);
and U10263 (N_10263,N_9671,N_9060);
and U10264 (N_10264,N_9709,N_9682);
nand U10265 (N_10265,N_9383,N_9475);
nor U10266 (N_10266,N_9008,N_9127);
and U10267 (N_10267,N_9620,N_9069);
or U10268 (N_10268,N_9012,N_9733);
nor U10269 (N_10269,N_9006,N_9216);
nor U10270 (N_10270,N_9488,N_9565);
nand U10271 (N_10271,N_9015,N_9318);
nand U10272 (N_10272,N_9547,N_9397);
xnor U10273 (N_10273,N_9290,N_9025);
nand U10274 (N_10274,N_9534,N_9075);
nor U10275 (N_10275,N_9531,N_9538);
xor U10276 (N_10276,N_9623,N_9711);
nor U10277 (N_10277,N_9063,N_9143);
nand U10278 (N_10278,N_9065,N_9444);
nand U10279 (N_10279,N_9427,N_9304);
nor U10280 (N_10280,N_9036,N_9606);
nor U10281 (N_10281,N_9057,N_9544);
xor U10282 (N_10282,N_9530,N_9198);
xnor U10283 (N_10283,N_9510,N_9682);
nor U10284 (N_10284,N_9622,N_9659);
nand U10285 (N_10285,N_9570,N_9197);
or U10286 (N_10286,N_9291,N_9451);
or U10287 (N_10287,N_9322,N_9569);
xor U10288 (N_10288,N_9727,N_9300);
nand U10289 (N_10289,N_9565,N_9290);
and U10290 (N_10290,N_9081,N_9034);
nand U10291 (N_10291,N_9218,N_9524);
nor U10292 (N_10292,N_9409,N_9459);
nand U10293 (N_10293,N_9544,N_9732);
or U10294 (N_10294,N_9518,N_9724);
nor U10295 (N_10295,N_9136,N_9253);
xnor U10296 (N_10296,N_9430,N_9144);
or U10297 (N_10297,N_9093,N_9732);
nor U10298 (N_10298,N_9005,N_9154);
and U10299 (N_10299,N_9208,N_9393);
or U10300 (N_10300,N_9254,N_9113);
nor U10301 (N_10301,N_9349,N_9624);
or U10302 (N_10302,N_9153,N_9113);
or U10303 (N_10303,N_9467,N_9171);
nand U10304 (N_10304,N_9502,N_9134);
xor U10305 (N_10305,N_9161,N_9637);
and U10306 (N_10306,N_9688,N_9275);
and U10307 (N_10307,N_9092,N_9642);
or U10308 (N_10308,N_9608,N_9223);
nor U10309 (N_10309,N_9085,N_9691);
xor U10310 (N_10310,N_9479,N_9743);
nand U10311 (N_10311,N_9653,N_9395);
and U10312 (N_10312,N_9237,N_9394);
nand U10313 (N_10313,N_9317,N_9645);
nand U10314 (N_10314,N_9212,N_9165);
nor U10315 (N_10315,N_9576,N_9240);
or U10316 (N_10316,N_9283,N_9604);
nand U10317 (N_10317,N_9500,N_9684);
xnor U10318 (N_10318,N_9430,N_9215);
xnor U10319 (N_10319,N_9096,N_9144);
or U10320 (N_10320,N_9093,N_9746);
xnor U10321 (N_10321,N_9140,N_9662);
nand U10322 (N_10322,N_9264,N_9020);
and U10323 (N_10323,N_9040,N_9165);
and U10324 (N_10324,N_9484,N_9645);
and U10325 (N_10325,N_9529,N_9737);
and U10326 (N_10326,N_9400,N_9637);
or U10327 (N_10327,N_9072,N_9143);
nor U10328 (N_10328,N_9633,N_9477);
nor U10329 (N_10329,N_9078,N_9160);
nand U10330 (N_10330,N_9542,N_9690);
nand U10331 (N_10331,N_9716,N_9394);
or U10332 (N_10332,N_9130,N_9421);
nand U10333 (N_10333,N_9269,N_9172);
nand U10334 (N_10334,N_9025,N_9308);
nand U10335 (N_10335,N_9228,N_9579);
and U10336 (N_10336,N_9397,N_9537);
nand U10337 (N_10337,N_9159,N_9695);
nor U10338 (N_10338,N_9692,N_9435);
or U10339 (N_10339,N_9685,N_9530);
or U10340 (N_10340,N_9287,N_9746);
or U10341 (N_10341,N_9114,N_9320);
and U10342 (N_10342,N_9686,N_9337);
or U10343 (N_10343,N_9588,N_9494);
nor U10344 (N_10344,N_9088,N_9362);
nor U10345 (N_10345,N_9421,N_9397);
nor U10346 (N_10346,N_9462,N_9502);
and U10347 (N_10347,N_9226,N_9115);
and U10348 (N_10348,N_9231,N_9191);
nand U10349 (N_10349,N_9356,N_9190);
or U10350 (N_10350,N_9357,N_9225);
and U10351 (N_10351,N_9735,N_9047);
or U10352 (N_10352,N_9057,N_9281);
nand U10353 (N_10353,N_9480,N_9443);
nand U10354 (N_10354,N_9525,N_9316);
nand U10355 (N_10355,N_9530,N_9590);
nand U10356 (N_10356,N_9166,N_9127);
nand U10357 (N_10357,N_9431,N_9656);
and U10358 (N_10358,N_9310,N_9555);
nor U10359 (N_10359,N_9422,N_9488);
or U10360 (N_10360,N_9429,N_9590);
nand U10361 (N_10361,N_9656,N_9089);
nand U10362 (N_10362,N_9267,N_9291);
nor U10363 (N_10363,N_9228,N_9117);
and U10364 (N_10364,N_9227,N_9401);
or U10365 (N_10365,N_9527,N_9550);
nor U10366 (N_10366,N_9160,N_9450);
nand U10367 (N_10367,N_9241,N_9319);
xnor U10368 (N_10368,N_9257,N_9550);
and U10369 (N_10369,N_9274,N_9573);
or U10370 (N_10370,N_9537,N_9716);
and U10371 (N_10371,N_9078,N_9563);
nor U10372 (N_10372,N_9666,N_9016);
or U10373 (N_10373,N_9289,N_9542);
and U10374 (N_10374,N_9651,N_9422);
and U10375 (N_10375,N_9460,N_9504);
nand U10376 (N_10376,N_9029,N_9725);
or U10377 (N_10377,N_9288,N_9369);
nand U10378 (N_10378,N_9169,N_9158);
nor U10379 (N_10379,N_9469,N_9265);
and U10380 (N_10380,N_9174,N_9608);
or U10381 (N_10381,N_9268,N_9018);
nor U10382 (N_10382,N_9397,N_9566);
nand U10383 (N_10383,N_9195,N_9229);
or U10384 (N_10384,N_9208,N_9656);
and U10385 (N_10385,N_9525,N_9455);
nand U10386 (N_10386,N_9172,N_9564);
nor U10387 (N_10387,N_9179,N_9260);
or U10388 (N_10388,N_9732,N_9660);
nand U10389 (N_10389,N_9031,N_9444);
or U10390 (N_10390,N_9534,N_9684);
nor U10391 (N_10391,N_9120,N_9039);
nand U10392 (N_10392,N_9695,N_9208);
and U10393 (N_10393,N_9335,N_9395);
nor U10394 (N_10394,N_9546,N_9456);
nor U10395 (N_10395,N_9433,N_9718);
xnor U10396 (N_10396,N_9714,N_9664);
nand U10397 (N_10397,N_9139,N_9332);
and U10398 (N_10398,N_9669,N_9469);
xor U10399 (N_10399,N_9347,N_9728);
nor U10400 (N_10400,N_9013,N_9418);
xor U10401 (N_10401,N_9048,N_9388);
or U10402 (N_10402,N_9515,N_9075);
nor U10403 (N_10403,N_9598,N_9151);
nand U10404 (N_10404,N_9542,N_9137);
and U10405 (N_10405,N_9600,N_9061);
nand U10406 (N_10406,N_9318,N_9587);
nand U10407 (N_10407,N_9357,N_9595);
nor U10408 (N_10408,N_9727,N_9478);
nand U10409 (N_10409,N_9069,N_9115);
nand U10410 (N_10410,N_9481,N_9742);
or U10411 (N_10411,N_9747,N_9674);
xnor U10412 (N_10412,N_9655,N_9612);
nor U10413 (N_10413,N_9198,N_9696);
nor U10414 (N_10414,N_9446,N_9219);
nand U10415 (N_10415,N_9022,N_9065);
nor U10416 (N_10416,N_9146,N_9276);
xnor U10417 (N_10417,N_9266,N_9257);
nand U10418 (N_10418,N_9010,N_9334);
and U10419 (N_10419,N_9342,N_9251);
nor U10420 (N_10420,N_9226,N_9591);
nand U10421 (N_10421,N_9334,N_9557);
or U10422 (N_10422,N_9558,N_9426);
nand U10423 (N_10423,N_9465,N_9190);
and U10424 (N_10424,N_9552,N_9646);
nand U10425 (N_10425,N_9698,N_9532);
nand U10426 (N_10426,N_9311,N_9360);
and U10427 (N_10427,N_9487,N_9590);
nor U10428 (N_10428,N_9490,N_9477);
nor U10429 (N_10429,N_9422,N_9112);
and U10430 (N_10430,N_9118,N_9383);
nand U10431 (N_10431,N_9669,N_9077);
and U10432 (N_10432,N_9209,N_9143);
xor U10433 (N_10433,N_9106,N_9710);
and U10434 (N_10434,N_9324,N_9139);
nor U10435 (N_10435,N_9444,N_9311);
nor U10436 (N_10436,N_9473,N_9052);
xnor U10437 (N_10437,N_9549,N_9219);
or U10438 (N_10438,N_9055,N_9714);
and U10439 (N_10439,N_9443,N_9404);
nor U10440 (N_10440,N_9413,N_9554);
nand U10441 (N_10441,N_9661,N_9709);
or U10442 (N_10442,N_9436,N_9055);
and U10443 (N_10443,N_9415,N_9108);
and U10444 (N_10444,N_9103,N_9566);
and U10445 (N_10445,N_9030,N_9312);
nand U10446 (N_10446,N_9332,N_9295);
and U10447 (N_10447,N_9089,N_9212);
nor U10448 (N_10448,N_9445,N_9735);
or U10449 (N_10449,N_9437,N_9046);
nor U10450 (N_10450,N_9389,N_9477);
xnor U10451 (N_10451,N_9195,N_9381);
nand U10452 (N_10452,N_9448,N_9375);
nand U10453 (N_10453,N_9091,N_9190);
nand U10454 (N_10454,N_9543,N_9544);
nand U10455 (N_10455,N_9385,N_9715);
or U10456 (N_10456,N_9209,N_9225);
nand U10457 (N_10457,N_9566,N_9328);
nand U10458 (N_10458,N_9127,N_9225);
and U10459 (N_10459,N_9706,N_9287);
or U10460 (N_10460,N_9605,N_9405);
nor U10461 (N_10461,N_9501,N_9508);
nor U10462 (N_10462,N_9340,N_9728);
or U10463 (N_10463,N_9389,N_9671);
nor U10464 (N_10464,N_9155,N_9103);
or U10465 (N_10465,N_9073,N_9540);
xor U10466 (N_10466,N_9184,N_9289);
nand U10467 (N_10467,N_9272,N_9369);
or U10468 (N_10468,N_9339,N_9326);
or U10469 (N_10469,N_9102,N_9271);
and U10470 (N_10470,N_9720,N_9295);
xnor U10471 (N_10471,N_9557,N_9012);
or U10472 (N_10472,N_9057,N_9292);
xnor U10473 (N_10473,N_9086,N_9699);
nor U10474 (N_10474,N_9159,N_9193);
nor U10475 (N_10475,N_9223,N_9683);
nand U10476 (N_10476,N_9713,N_9312);
nor U10477 (N_10477,N_9050,N_9418);
nor U10478 (N_10478,N_9172,N_9622);
nor U10479 (N_10479,N_9521,N_9423);
and U10480 (N_10480,N_9201,N_9505);
nand U10481 (N_10481,N_9698,N_9120);
or U10482 (N_10482,N_9613,N_9133);
or U10483 (N_10483,N_9111,N_9327);
nor U10484 (N_10484,N_9458,N_9264);
or U10485 (N_10485,N_9178,N_9421);
or U10486 (N_10486,N_9303,N_9304);
nor U10487 (N_10487,N_9017,N_9364);
xnor U10488 (N_10488,N_9626,N_9010);
nor U10489 (N_10489,N_9231,N_9573);
nand U10490 (N_10490,N_9682,N_9036);
or U10491 (N_10491,N_9405,N_9576);
or U10492 (N_10492,N_9506,N_9290);
xor U10493 (N_10493,N_9473,N_9065);
and U10494 (N_10494,N_9743,N_9722);
nor U10495 (N_10495,N_9669,N_9262);
xor U10496 (N_10496,N_9083,N_9651);
or U10497 (N_10497,N_9420,N_9470);
nand U10498 (N_10498,N_9279,N_9293);
nor U10499 (N_10499,N_9547,N_9368);
and U10500 (N_10500,N_10317,N_9997);
and U10501 (N_10501,N_10224,N_10487);
xor U10502 (N_10502,N_9790,N_10477);
or U10503 (N_10503,N_10457,N_10361);
nand U10504 (N_10504,N_9852,N_10183);
nor U10505 (N_10505,N_9941,N_9774);
nand U10506 (N_10506,N_10357,N_9798);
nand U10507 (N_10507,N_10134,N_10377);
or U10508 (N_10508,N_9827,N_10354);
and U10509 (N_10509,N_9858,N_9815);
and U10510 (N_10510,N_9831,N_9856);
and U10511 (N_10511,N_10226,N_10182);
and U10512 (N_10512,N_10439,N_10077);
nor U10513 (N_10513,N_9800,N_10336);
nand U10514 (N_10514,N_10199,N_10192);
nor U10515 (N_10515,N_9962,N_10173);
or U10516 (N_10516,N_10236,N_9986);
or U10517 (N_10517,N_10310,N_10007);
or U10518 (N_10518,N_10018,N_9786);
nor U10519 (N_10519,N_10157,N_9878);
xor U10520 (N_10520,N_10086,N_10050);
and U10521 (N_10521,N_10290,N_10359);
nand U10522 (N_10522,N_10483,N_10385);
nor U10523 (N_10523,N_9785,N_9825);
and U10524 (N_10524,N_10459,N_10093);
and U10525 (N_10525,N_9796,N_10175);
xnor U10526 (N_10526,N_10446,N_9950);
xnor U10527 (N_10527,N_10325,N_10328);
and U10528 (N_10528,N_9801,N_10329);
and U10529 (N_10529,N_10153,N_9864);
or U10530 (N_10530,N_10131,N_10179);
nand U10531 (N_10531,N_10389,N_10168);
xor U10532 (N_10532,N_10479,N_10220);
xnor U10533 (N_10533,N_10291,N_10421);
and U10534 (N_10534,N_10424,N_10104);
nand U10535 (N_10535,N_9953,N_9799);
or U10536 (N_10536,N_10258,N_9853);
and U10537 (N_10537,N_9913,N_9837);
nand U10538 (N_10538,N_10367,N_10268);
nand U10539 (N_10539,N_10466,N_10478);
xor U10540 (N_10540,N_9984,N_10218);
nor U10541 (N_10541,N_10085,N_10038);
nor U10542 (N_10542,N_10090,N_10209);
or U10543 (N_10543,N_9813,N_10376);
nor U10544 (N_10544,N_9869,N_10072);
nor U10545 (N_10545,N_10193,N_9964);
nand U10546 (N_10546,N_10493,N_10341);
or U10547 (N_10547,N_10012,N_9781);
and U10548 (N_10548,N_10499,N_10396);
or U10549 (N_10549,N_10055,N_10471);
and U10550 (N_10550,N_10127,N_10075);
nand U10551 (N_10551,N_10304,N_10045);
xor U10552 (N_10552,N_10152,N_9940);
and U10553 (N_10553,N_10022,N_9885);
xor U10554 (N_10554,N_10383,N_10024);
nor U10555 (N_10555,N_9808,N_10240);
or U10556 (N_10556,N_10373,N_9814);
nand U10557 (N_10557,N_9752,N_10497);
nor U10558 (N_10558,N_10222,N_9886);
or U10559 (N_10559,N_10108,N_9865);
nor U10560 (N_10560,N_10340,N_9919);
and U10561 (N_10561,N_10350,N_9771);
and U10562 (N_10562,N_10032,N_10051);
or U10563 (N_10563,N_10380,N_10070);
nor U10564 (N_10564,N_10393,N_10261);
nand U10565 (N_10565,N_9947,N_10276);
nor U10566 (N_10566,N_10403,N_9860);
nor U10567 (N_10567,N_10027,N_10008);
nand U10568 (N_10568,N_10370,N_9980);
nor U10569 (N_10569,N_9904,N_10064);
or U10570 (N_10570,N_10492,N_10006);
nor U10571 (N_10571,N_10188,N_10144);
nand U10572 (N_10572,N_10302,N_9973);
nor U10573 (N_10573,N_9952,N_10481);
or U10574 (N_10574,N_10358,N_9916);
and U10575 (N_10575,N_10330,N_10475);
nand U10576 (N_10576,N_10409,N_10133);
and U10577 (N_10577,N_9863,N_9918);
and U10578 (N_10578,N_9944,N_9974);
and U10579 (N_10579,N_10023,N_10216);
or U10580 (N_10580,N_9993,N_10034);
and U10581 (N_10581,N_10000,N_10009);
xor U10582 (N_10582,N_9818,N_9971);
and U10583 (N_10583,N_10145,N_10252);
nand U10584 (N_10584,N_10489,N_10338);
nand U10585 (N_10585,N_9921,N_10476);
and U10586 (N_10586,N_10260,N_10337);
or U10587 (N_10587,N_9855,N_10442);
nand U10588 (N_10588,N_10427,N_10046);
or U10589 (N_10589,N_9914,N_10165);
nand U10590 (N_10590,N_10113,N_9767);
and U10591 (N_10591,N_9816,N_10114);
nor U10592 (N_10592,N_10102,N_9908);
nand U10593 (N_10593,N_10155,N_9893);
nand U10594 (N_10594,N_10109,N_9776);
nand U10595 (N_10595,N_10245,N_9835);
nor U10596 (N_10596,N_9762,N_10162);
xnor U10597 (N_10597,N_10399,N_10158);
or U10598 (N_10598,N_9938,N_10323);
and U10599 (N_10599,N_10130,N_10184);
or U10600 (N_10600,N_10456,N_10095);
or U10601 (N_10601,N_10147,N_9948);
and U10602 (N_10602,N_9846,N_10215);
or U10603 (N_10603,N_10124,N_9795);
nand U10604 (N_10604,N_9868,N_9793);
nor U10605 (N_10605,N_10266,N_10278);
and U10606 (N_10606,N_9770,N_10031);
nor U10607 (N_10607,N_9960,N_9757);
or U10608 (N_10608,N_10234,N_10042);
or U10609 (N_10609,N_10335,N_10029);
xor U10610 (N_10610,N_9876,N_9923);
and U10611 (N_10611,N_10472,N_9780);
or U10612 (N_10612,N_10422,N_10030);
nand U10613 (N_10613,N_10464,N_9990);
nand U10614 (N_10614,N_10288,N_9942);
nand U10615 (N_10615,N_9945,N_9961);
and U10616 (N_10616,N_10391,N_10308);
nand U10617 (N_10617,N_9955,N_9826);
and U10618 (N_10618,N_9978,N_10415);
and U10619 (N_10619,N_9873,N_10433);
or U10620 (N_10620,N_10300,N_9751);
or U10621 (N_10621,N_10397,N_9784);
xnor U10622 (N_10622,N_10198,N_9766);
nand U10623 (N_10623,N_10257,N_9843);
nor U10624 (N_10624,N_9934,N_10280);
and U10625 (N_10625,N_9807,N_9834);
xor U10626 (N_10626,N_9794,N_10004);
or U10627 (N_10627,N_10356,N_10473);
nand U10628 (N_10628,N_10021,N_10423);
nor U10629 (N_10629,N_9898,N_10071);
and U10630 (N_10630,N_9992,N_9922);
nand U10631 (N_10631,N_9805,N_10332);
or U10632 (N_10632,N_10149,N_10454);
xor U10633 (N_10633,N_9970,N_9870);
or U10634 (N_10634,N_9809,N_9845);
and U10635 (N_10635,N_9946,N_9896);
and U10636 (N_10636,N_10203,N_10307);
nor U10637 (N_10637,N_9832,N_10270);
nor U10638 (N_10638,N_10279,N_10106);
or U10639 (N_10639,N_9985,N_10141);
or U10640 (N_10640,N_10246,N_9877);
xnor U10641 (N_10641,N_9867,N_10043);
and U10642 (N_10642,N_9819,N_10387);
or U10643 (N_10643,N_10343,N_9811);
nor U10644 (N_10644,N_9967,N_10116);
nor U10645 (N_10645,N_9889,N_9912);
xnor U10646 (N_10646,N_10219,N_9951);
or U10647 (N_10647,N_10002,N_10296);
or U10648 (N_10648,N_10289,N_10191);
and U10649 (N_10649,N_10281,N_10394);
or U10650 (N_10650,N_9872,N_10255);
xor U10651 (N_10651,N_10154,N_10011);
or U10652 (N_10652,N_10275,N_10486);
xnor U10653 (N_10653,N_10405,N_10205);
or U10654 (N_10654,N_10416,N_9936);
nand U10655 (N_10655,N_9920,N_10259);
nand U10656 (N_10656,N_9803,N_10283);
and U10657 (N_10657,N_10419,N_10347);
and U10658 (N_10658,N_10312,N_10146);
or U10659 (N_10659,N_10441,N_10170);
or U10660 (N_10660,N_10488,N_10083);
or U10661 (N_10661,N_9958,N_10334);
and U10662 (N_10662,N_10440,N_10402);
and U10663 (N_10663,N_9829,N_9933);
nor U10664 (N_10664,N_10041,N_10292);
nand U10665 (N_10665,N_9847,N_10306);
nor U10666 (N_10666,N_10311,N_9894);
nor U10667 (N_10667,N_10429,N_10273);
nor U10668 (N_10668,N_10067,N_10298);
or U10669 (N_10669,N_9965,N_10431);
nor U10670 (N_10670,N_10408,N_10470);
and U10671 (N_10671,N_10436,N_10005);
and U10672 (N_10672,N_9966,N_10111);
xor U10673 (N_10673,N_10461,N_9778);
and U10674 (N_10674,N_9888,N_10189);
xor U10675 (N_10675,N_10434,N_10379);
nand U10676 (N_10676,N_10372,N_10204);
or U10677 (N_10677,N_10081,N_10301);
nand U10678 (N_10678,N_9791,N_10395);
nand U10679 (N_10679,N_10344,N_10003);
or U10680 (N_10680,N_10167,N_10212);
and U10681 (N_10681,N_9976,N_9817);
or U10682 (N_10682,N_10412,N_10069);
or U10683 (N_10683,N_10368,N_10314);
and U10684 (N_10684,N_10333,N_10411);
nor U10685 (N_10685,N_9820,N_9957);
and U10686 (N_10686,N_9972,N_10015);
or U10687 (N_10687,N_10062,N_10365);
xor U10688 (N_10688,N_9879,N_10139);
nand U10689 (N_10689,N_10094,N_10213);
nand U10690 (N_10690,N_10207,N_10232);
nor U10691 (N_10691,N_10404,N_10174);
nor U10692 (N_10692,N_9838,N_10088);
xor U10693 (N_10693,N_9821,N_9932);
and U10694 (N_10694,N_10110,N_9851);
nor U10695 (N_10695,N_10156,N_10371);
and U10696 (N_10696,N_10375,N_9979);
nor U10697 (N_10697,N_9887,N_10360);
nand U10698 (N_10698,N_10089,N_9789);
nand U10699 (N_10699,N_10233,N_9988);
nand U10700 (N_10700,N_10407,N_9849);
nor U10701 (N_10701,N_10313,N_10346);
and U10702 (N_10702,N_10120,N_10249);
and U10703 (N_10703,N_10128,N_10238);
and U10704 (N_10704,N_10010,N_10017);
and U10705 (N_10705,N_10248,N_10122);
or U10706 (N_10706,N_10166,N_9880);
xnor U10707 (N_10707,N_10037,N_10293);
nand U10708 (N_10708,N_10187,N_10498);
nor U10709 (N_10709,N_10227,N_10342);
nor U10710 (N_10710,N_9959,N_10348);
nor U10711 (N_10711,N_10103,N_10381);
nand U10712 (N_10712,N_10277,N_10214);
nor U10713 (N_10713,N_9759,N_10445);
and U10714 (N_10714,N_10345,N_10285);
or U10715 (N_10715,N_9975,N_10410);
nand U10716 (N_10716,N_10327,N_10105);
nor U10717 (N_10717,N_10016,N_9963);
and U10718 (N_10718,N_10449,N_10355);
and U10719 (N_10719,N_10142,N_10195);
nand U10720 (N_10720,N_9772,N_9968);
nand U10721 (N_10721,N_9859,N_10044);
or U10722 (N_10722,N_10417,N_10331);
nand U10723 (N_10723,N_9848,N_9833);
or U10724 (N_10724,N_10303,N_9861);
or U10725 (N_10725,N_10339,N_9930);
or U10726 (N_10726,N_10056,N_10469);
xor U10727 (N_10727,N_10353,N_10443);
or U10728 (N_10728,N_10190,N_9895);
nor U10729 (N_10729,N_9802,N_10181);
nand U10730 (N_10730,N_10140,N_9905);
or U10731 (N_10731,N_10091,N_10326);
nor U10732 (N_10732,N_10135,N_10161);
nand U10733 (N_10733,N_10059,N_10388);
xnor U10734 (N_10734,N_10467,N_9939);
nand U10735 (N_10735,N_9787,N_9812);
or U10736 (N_10736,N_10100,N_10305);
and U10737 (N_10737,N_10420,N_9983);
or U10738 (N_10738,N_9761,N_10036);
xor U10739 (N_10739,N_10262,N_10125);
and U10740 (N_10740,N_9989,N_9760);
xor U10741 (N_10741,N_10150,N_9931);
or U10742 (N_10742,N_9792,N_9764);
or U10743 (N_10743,N_9854,N_10014);
or U10744 (N_10744,N_10066,N_9937);
and U10745 (N_10745,N_10210,N_10185);
and U10746 (N_10746,N_10241,N_10495);
and U10747 (N_10747,N_10386,N_10484);
xnor U10748 (N_10748,N_10418,N_10269);
and U10749 (N_10749,N_10065,N_9755);
and U10750 (N_10750,N_10237,N_9783);
and U10751 (N_10751,N_9823,N_10052);
xnor U10752 (N_10752,N_10097,N_10164);
nand U10753 (N_10753,N_9765,N_9911);
nand U10754 (N_10754,N_10364,N_10132);
and U10755 (N_10755,N_10448,N_10073);
xnor U10756 (N_10756,N_10425,N_10490);
or U10757 (N_10757,N_9857,N_9871);
and U10758 (N_10758,N_9994,N_10148);
and U10759 (N_10759,N_10112,N_10206);
xnor U10760 (N_10760,N_9927,N_10398);
nor U10761 (N_10761,N_9754,N_10435);
nand U10762 (N_10762,N_10363,N_10460);
or U10763 (N_10763,N_10256,N_9901);
or U10764 (N_10764,N_10352,N_10137);
nand U10765 (N_10765,N_9999,N_10178);
or U10766 (N_10766,N_10078,N_10230);
xnor U10767 (N_10767,N_10171,N_9906);
and U10768 (N_10768,N_10201,N_10033);
or U10769 (N_10769,N_9756,N_10400);
and U10770 (N_10770,N_9915,N_10463);
and U10771 (N_10771,N_10229,N_10428);
nor U10772 (N_10772,N_10482,N_10468);
and U10773 (N_10773,N_10208,N_9758);
or U10774 (N_10774,N_9881,N_10079);
xnor U10775 (N_10775,N_9890,N_10076);
or U10776 (N_10776,N_9775,N_10284);
xnor U10777 (N_10777,N_10172,N_10058);
nand U10778 (N_10778,N_10319,N_10271);
xor U10779 (N_10779,N_10272,N_10063);
and U10780 (N_10780,N_9949,N_10251);
and U10781 (N_10781,N_9884,N_10294);
and U10782 (N_10782,N_9824,N_10082);
nor U10783 (N_10783,N_10239,N_9788);
or U10784 (N_10784,N_10013,N_10223);
nand U10785 (N_10785,N_9977,N_10384);
nand U10786 (N_10786,N_9830,N_10320);
nor U10787 (N_10787,N_10099,N_10480);
or U10788 (N_10788,N_10465,N_10321);
nor U10789 (N_10789,N_10322,N_9883);
nor U10790 (N_10790,N_9777,N_10426);
nor U10791 (N_10791,N_10282,N_10121);
and U10792 (N_10792,N_10366,N_10160);
and U10793 (N_10793,N_10228,N_10362);
xor U10794 (N_10794,N_10315,N_10485);
and U10795 (N_10795,N_10450,N_10453);
or U10796 (N_10796,N_10231,N_10039);
or U10797 (N_10797,N_10151,N_10458);
and U10798 (N_10798,N_10115,N_10068);
nand U10799 (N_10799,N_10474,N_9897);
nor U10800 (N_10800,N_10107,N_10318);
xor U10801 (N_10801,N_9902,N_9917);
nand U10802 (N_10802,N_9995,N_10020);
nor U10803 (N_10803,N_9996,N_9969);
or U10804 (N_10804,N_10451,N_10001);
nand U10805 (N_10805,N_10040,N_10123);
xor U10806 (N_10806,N_9822,N_10286);
nand U10807 (N_10807,N_10267,N_9875);
xor U10808 (N_10808,N_9782,N_10309);
xnor U10809 (N_10809,N_9768,N_10295);
and U10810 (N_10810,N_10047,N_10194);
or U10811 (N_10811,N_10126,N_10138);
or U10812 (N_10812,N_10287,N_9991);
or U10813 (N_10813,N_10054,N_10119);
nor U10814 (N_10814,N_9891,N_10049);
or U10815 (N_10815,N_10101,N_10378);
and U10816 (N_10816,N_10243,N_10143);
nand U10817 (N_10817,N_10176,N_9841);
and U10818 (N_10818,N_9935,N_9842);
nand U10819 (N_10819,N_9850,N_10196);
and U10820 (N_10820,N_9928,N_9804);
nor U10821 (N_10821,N_9866,N_10316);
nand U10822 (N_10822,N_10211,N_9874);
nand U10823 (N_10823,N_9779,N_10392);
nand U10824 (N_10824,N_10163,N_10035);
nor U10825 (N_10825,N_10274,N_10254);
xnor U10826 (N_10826,N_10096,N_9924);
nand U10827 (N_10827,N_10026,N_9954);
nand U10828 (N_10828,N_10351,N_10048);
or U10829 (N_10829,N_9806,N_9943);
and U10830 (N_10830,N_10430,N_9900);
nand U10831 (N_10831,N_10414,N_10080);
or U10832 (N_10832,N_10053,N_10061);
and U10833 (N_10833,N_10025,N_10202);
nand U10834 (N_10834,N_10217,N_10197);
nand U10835 (N_10835,N_10263,N_9840);
nor U10836 (N_10836,N_9763,N_10265);
xor U10837 (N_10837,N_9836,N_10117);
and U10838 (N_10838,N_10401,N_9753);
or U10839 (N_10839,N_10299,N_9828);
nand U10840 (N_10840,N_10136,N_9956);
nand U10841 (N_10841,N_10369,N_10159);
or U10842 (N_10842,N_9909,N_10247);
and U10843 (N_10843,N_10235,N_10250);
nand U10844 (N_10844,N_10225,N_9882);
nand U10845 (N_10845,N_10432,N_9982);
or U10846 (N_10846,N_9910,N_9899);
nor U10847 (N_10847,N_10242,N_10406);
xor U10848 (N_10848,N_10221,N_9926);
nand U10849 (N_10849,N_10390,N_9810);
nor U10850 (N_10850,N_10437,N_10324);
nor U10851 (N_10851,N_9929,N_10118);
and U10852 (N_10852,N_10177,N_9769);
nor U10853 (N_10853,N_9907,N_9998);
or U10854 (N_10854,N_10186,N_10084);
and U10855 (N_10855,N_9862,N_10180);
or U10856 (N_10856,N_10444,N_9844);
and U10857 (N_10857,N_10028,N_9903);
xnor U10858 (N_10858,N_9892,N_10382);
and U10859 (N_10859,N_9839,N_10253);
or U10860 (N_10860,N_9925,N_10413);
and U10861 (N_10861,N_10374,N_10129);
and U10862 (N_10862,N_10169,N_10019);
nand U10863 (N_10863,N_9987,N_10297);
nand U10864 (N_10864,N_10491,N_10060);
or U10865 (N_10865,N_10496,N_10057);
and U10866 (N_10866,N_10244,N_10494);
and U10867 (N_10867,N_10452,N_10087);
nor U10868 (N_10868,N_9750,N_10098);
nand U10869 (N_10869,N_9981,N_10200);
or U10870 (N_10870,N_10438,N_10447);
or U10871 (N_10871,N_10264,N_9797);
nor U10872 (N_10872,N_10074,N_10092);
xnor U10873 (N_10873,N_10349,N_9773);
nand U10874 (N_10874,N_10455,N_10462);
or U10875 (N_10875,N_10405,N_9793);
and U10876 (N_10876,N_10081,N_10027);
or U10877 (N_10877,N_10001,N_10191);
nor U10878 (N_10878,N_10437,N_10057);
nand U10879 (N_10879,N_10302,N_10355);
and U10880 (N_10880,N_9914,N_10039);
nor U10881 (N_10881,N_10115,N_10274);
or U10882 (N_10882,N_10361,N_10282);
xor U10883 (N_10883,N_10082,N_10057);
or U10884 (N_10884,N_9998,N_9798);
nand U10885 (N_10885,N_10322,N_10115);
nor U10886 (N_10886,N_10109,N_10203);
or U10887 (N_10887,N_10035,N_10488);
or U10888 (N_10888,N_10246,N_10260);
xor U10889 (N_10889,N_9905,N_10297);
nand U10890 (N_10890,N_10321,N_10128);
nand U10891 (N_10891,N_10187,N_10065);
nand U10892 (N_10892,N_10335,N_9970);
nor U10893 (N_10893,N_10242,N_9799);
or U10894 (N_10894,N_9884,N_9762);
nand U10895 (N_10895,N_10017,N_9966);
nand U10896 (N_10896,N_9828,N_10203);
or U10897 (N_10897,N_9843,N_10321);
and U10898 (N_10898,N_10097,N_9793);
or U10899 (N_10899,N_10373,N_10379);
or U10900 (N_10900,N_9914,N_10451);
and U10901 (N_10901,N_9832,N_10419);
nor U10902 (N_10902,N_9877,N_10232);
nand U10903 (N_10903,N_10110,N_10180);
or U10904 (N_10904,N_10121,N_10146);
nand U10905 (N_10905,N_10375,N_10067);
and U10906 (N_10906,N_10213,N_10260);
or U10907 (N_10907,N_10390,N_10396);
nor U10908 (N_10908,N_10077,N_10470);
nand U10909 (N_10909,N_10341,N_10317);
xor U10910 (N_10910,N_10353,N_9808);
nor U10911 (N_10911,N_10155,N_9926);
and U10912 (N_10912,N_10094,N_10429);
or U10913 (N_10913,N_10397,N_10170);
xor U10914 (N_10914,N_9873,N_10452);
or U10915 (N_10915,N_10266,N_10004);
and U10916 (N_10916,N_9900,N_10044);
or U10917 (N_10917,N_10261,N_9829);
nand U10918 (N_10918,N_9768,N_10231);
or U10919 (N_10919,N_10266,N_9898);
nand U10920 (N_10920,N_10077,N_9827);
nor U10921 (N_10921,N_9860,N_10448);
nand U10922 (N_10922,N_10025,N_9986);
nand U10923 (N_10923,N_10052,N_10231);
nor U10924 (N_10924,N_9980,N_10450);
xnor U10925 (N_10925,N_10425,N_9933);
nand U10926 (N_10926,N_10237,N_9857);
and U10927 (N_10927,N_10138,N_10283);
and U10928 (N_10928,N_10331,N_10023);
or U10929 (N_10929,N_10339,N_10376);
nand U10930 (N_10930,N_10149,N_10117);
nand U10931 (N_10931,N_10253,N_9996);
nand U10932 (N_10932,N_10208,N_9943);
xor U10933 (N_10933,N_10216,N_10127);
nor U10934 (N_10934,N_9981,N_9846);
nor U10935 (N_10935,N_9846,N_10069);
nand U10936 (N_10936,N_10132,N_10052);
nor U10937 (N_10937,N_9819,N_10072);
or U10938 (N_10938,N_10286,N_10496);
or U10939 (N_10939,N_10218,N_9814);
nand U10940 (N_10940,N_10334,N_9831);
and U10941 (N_10941,N_10284,N_10274);
nand U10942 (N_10942,N_9975,N_10157);
or U10943 (N_10943,N_10336,N_10315);
or U10944 (N_10944,N_10370,N_9828);
nor U10945 (N_10945,N_10144,N_9946);
or U10946 (N_10946,N_9889,N_10315);
and U10947 (N_10947,N_10141,N_10368);
nand U10948 (N_10948,N_9885,N_9864);
nand U10949 (N_10949,N_10056,N_10155);
or U10950 (N_10950,N_10445,N_10074);
or U10951 (N_10951,N_10346,N_10376);
nand U10952 (N_10952,N_9923,N_9750);
nor U10953 (N_10953,N_10061,N_10412);
nand U10954 (N_10954,N_10080,N_10423);
nor U10955 (N_10955,N_10196,N_9878);
nor U10956 (N_10956,N_10213,N_10275);
xor U10957 (N_10957,N_9946,N_10225);
or U10958 (N_10958,N_10313,N_10193);
and U10959 (N_10959,N_10295,N_9880);
nand U10960 (N_10960,N_9766,N_10392);
and U10961 (N_10961,N_10397,N_10469);
nor U10962 (N_10962,N_9996,N_10033);
nand U10963 (N_10963,N_10033,N_10290);
nor U10964 (N_10964,N_9812,N_9780);
xor U10965 (N_10965,N_10244,N_10045);
and U10966 (N_10966,N_9992,N_9966);
and U10967 (N_10967,N_10475,N_9769);
or U10968 (N_10968,N_10237,N_10397);
and U10969 (N_10969,N_10258,N_10212);
nor U10970 (N_10970,N_10306,N_9750);
nand U10971 (N_10971,N_10004,N_10453);
and U10972 (N_10972,N_10018,N_10393);
or U10973 (N_10973,N_9871,N_10493);
and U10974 (N_10974,N_10196,N_10049);
nand U10975 (N_10975,N_10231,N_9869);
nor U10976 (N_10976,N_10041,N_10148);
or U10977 (N_10977,N_10486,N_10432);
or U10978 (N_10978,N_10451,N_9829);
xnor U10979 (N_10979,N_9810,N_10281);
and U10980 (N_10980,N_10409,N_9953);
and U10981 (N_10981,N_9923,N_10073);
xnor U10982 (N_10982,N_10128,N_10299);
nor U10983 (N_10983,N_10198,N_9908);
nor U10984 (N_10984,N_10477,N_9841);
and U10985 (N_10985,N_10063,N_10444);
nor U10986 (N_10986,N_9997,N_9950);
or U10987 (N_10987,N_9874,N_10395);
nand U10988 (N_10988,N_10430,N_10491);
or U10989 (N_10989,N_10104,N_10278);
or U10990 (N_10990,N_10498,N_9754);
or U10991 (N_10991,N_9781,N_10263);
and U10992 (N_10992,N_10175,N_9824);
nand U10993 (N_10993,N_10222,N_10445);
nand U10994 (N_10994,N_9991,N_10057);
xnor U10995 (N_10995,N_10077,N_10209);
nand U10996 (N_10996,N_10498,N_10021);
nor U10997 (N_10997,N_10255,N_9966);
nor U10998 (N_10998,N_10238,N_10353);
or U10999 (N_10999,N_9890,N_10420);
nand U11000 (N_11000,N_10197,N_10116);
or U11001 (N_11001,N_10255,N_9805);
nor U11002 (N_11002,N_10140,N_10361);
nand U11003 (N_11003,N_9902,N_9932);
or U11004 (N_11004,N_9929,N_10348);
nor U11005 (N_11005,N_9759,N_9750);
or U11006 (N_11006,N_9962,N_10201);
nor U11007 (N_11007,N_10092,N_10380);
and U11008 (N_11008,N_9825,N_10460);
nor U11009 (N_11009,N_10241,N_10319);
nand U11010 (N_11010,N_9879,N_9752);
nand U11011 (N_11011,N_9768,N_10420);
xnor U11012 (N_11012,N_9783,N_10302);
nand U11013 (N_11013,N_10167,N_9854);
and U11014 (N_11014,N_9873,N_10380);
and U11015 (N_11015,N_9919,N_9834);
xor U11016 (N_11016,N_10298,N_10118);
and U11017 (N_11017,N_10271,N_10460);
nor U11018 (N_11018,N_9823,N_9902);
or U11019 (N_11019,N_10220,N_9890);
nor U11020 (N_11020,N_10299,N_10171);
nand U11021 (N_11021,N_9788,N_9848);
and U11022 (N_11022,N_10375,N_10219);
and U11023 (N_11023,N_9985,N_10316);
nor U11024 (N_11024,N_10313,N_9868);
and U11025 (N_11025,N_9778,N_10285);
xnor U11026 (N_11026,N_9869,N_9788);
nand U11027 (N_11027,N_10465,N_9858);
or U11028 (N_11028,N_10300,N_9951);
nor U11029 (N_11029,N_9907,N_10456);
or U11030 (N_11030,N_9955,N_10271);
nand U11031 (N_11031,N_10205,N_9942);
nor U11032 (N_11032,N_10420,N_10143);
nor U11033 (N_11033,N_10066,N_9787);
and U11034 (N_11034,N_9898,N_9924);
and U11035 (N_11035,N_10309,N_9939);
and U11036 (N_11036,N_10443,N_10471);
or U11037 (N_11037,N_10375,N_9860);
or U11038 (N_11038,N_10063,N_9816);
nand U11039 (N_11039,N_10102,N_10345);
or U11040 (N_11040,N_9945,N_10413);
and U11041 (N_11041,N_9924,N_10216);
nand U11042 (N_11042,N_10384,N_10419);
nor U11043 (N_11043,N_10272,N_10064);
xor U11044 (N_11044,N_10338,N_10289);
nor U11045 (N_11045,N_10461,N_9906);
nand U11046 (N_11046,N_10194,N_10167);
nor U11047 (N_11047,N_10027,N_9777);
nor U11048 (N_11048,N_10465,N_10298);
and U11049 (N_11049,N_9927,N_10197);
and U11050 (N_11050,N_10293,N_10430);
xor U11051 (N_11051,N_10036,N_10370);
and U11052 (N_11052,N_9876,N_9883);
and U11053 (N_11053,N_10357,N_10498);
and U11054 (N_11054,N_9922,N_10220);
xor U11055 (N_11055,N_9845,N_10391);
xnor U11056 (N_11056,N_10315,N_10025);
or U11057 (N_11057,N_10362,N_9908);
and U11058 (N_11058,N_10024,N_10282);
or U11059 (N_11059,N_9991,N_10383);
nand U11060 (N_11060,N_10087,N_10288);
nand U11061 (N_11061,N_9871,N_9903);
nor U11062 (N_11062,N_9832,N_9960);
and U11063 (N_11063,N_9945,N_9886);
xor U11064 (N_11064,N_10344,N_10411);
xor U11065 (N_11065,N_10057,N_9976);
and U11066 (N_11066,N_10179,N_10051);
nor U11067 (N_11067,N_9872,N_10475);
and U11068 (N_11068,N_9975,N_10040);
nand U11069 (N_11069,N_10151,N_10059);
and U11070 (N_11070,N_10112,N_9910);
nand U11071 (N_11071,N_10071,N_10234);
nor U11072 (N_11072,N_10270,N_9916);
nor U11073 (N_11073,N_10479,N_10026);
xor U11074 (N_11074,N_9925,N_9815);
nor U11075 (N_11075,N_10146,N_10475);
or U11076 (N_11076,N_9836,N_10493);
or U11077 (N_11077,N_10072,N_10283);
or U11078 (N_11078,N_10400,N_10349);
and U11079 (N_11079,N_9783,N_10016);
nor U11080 (N_11080,N_9844,N_10395);
and U11081 (N_11081,N_9833,N_10209);
or U11082 (N_11082,N_10251,N_10454);
nor U11083 (N_11083,N_10186,N_9754);
xnor U11084 (N_11084,N_9803,N_9867);
nand U11085 (N_11085,N_9753,N_9896);
or U11086 (N_11086,N_9857,N_10236);
nor U11087 (N_11087,N_10496,N_10251);
and U11088 (N_11088,N_10413,N_9992);
nand U11089 (N_11089,N_9911,N_10141);
nor U11090 (N_11090,N_10412,N_10214);
xnor U11091 (N_11091,N_9901,N_10415);
and U11092 (N_11092,N_9796,N_10146);
and U11093 (N_11093,N_10075,N_9795);
and U11094 (N_11094,N_10296,N_10033);
or U11095 (N_11095,N_9753,N_10246);
xor U11096 (N_11096,N_10145,N_10268);
nand U11097 (N_11097,N_10020,N_10384);
nor U11098 (N_11098,N_9868,N_9932);
or U11099 (N_11099,N_10124,N_10122);
nand U11100 (N_11100,N_9763,N_9818);
and U11101 (N_11101,N_9860,N_10290);
and U11102 (N_11102,N_9942,N_10482);
or U11103 (N_11103,N_9935,N_9800);
nand U11104 (N_11104,N_10231,N_10132);
nand U11105 (N_11105,N_10042,N_9965);
nand U11106 (N_11106,N_10124,N_10289);
nand U11107 (N_11107,N_9862,N_10489);
or U11108 (N_11108,N_9779,N_10272);
or U11109 (N_11109,N_10495,N_9928);
and U11110 (N_11110,N_10389,N_10083);
xor U11111 (N_11111,N_9916,N_10142);
nor U11112 (N_11112,N_9790,N_9926);
nor U11113 (N_11113,N_10073,N_10015);
nor U11114 (N_11114,N_10434,N_9816);
and U11115 (N_11115,N_10015,N_10025);
or U11116 (N_11116,N_10199,N_10449);
nor U11117 (N_11117,N_9802,N_10369);
nand U11118 (N_11118,N_10342,N_9997);
nor U11119 (N_11119,N_10420,N_9819);
nor U11120 (N_11120,N_10078,N_10083);
and U11121 (N_11121,N_10381,N_10464);
nand U11122 (N_11122,N_9867,N_9820);
nand U11123 (N_11123,N_10193,N_10153);
or U11124 (N_11124,N_10268,N_10242);
or U11125 (N_11125,N_10233,N_10387);
nor U11126 (N_11126,N_9976,N_10328);
nor U11127 (N_11127,N_10468,N_9982);
or U11128 (N_11128,N_10156,N_9889);
or U11129 (N_11129,N_10458,N_9950);
nor U11130 (N_11130,N_10148,N_9766);
xor U11131 (N_11131,N_10418,N_10165);
and U11132 (N_11132,N_10115,N_10242);
xnor U11133 (N_11133,N_10112,N_10355);
or U11134 (N_11134,N_9957,N_9885);
nor U11135 (N_11135,N_10068,N_9982);
and U11136 (N_11136,N_9997,N_10116);
nor U11137 (N_11137,N_10143,N_10426);
nor U11138 (N_11138,N_10053,N_10179);
and U11139 (N_11139,N_10453,N_10030);
nor U11140 (N_11140,N_9964,N_10317);
nand U11141 (N_11141,N_10207,N_9894);
or U11142 (N_11142,N_9884,N_10106);
or U11143 (N_11143,N_9998,N_10203);
and U11144 (N_11144,N_9879,N_10333);
xnor U11145 (N_11145,N_10405,N_10308);
or U11146 (N_11146,N_9824,N_9755);
nor U11147 (N_11147,N_10028,N_10090);
and U11148 (N_11148,N_10262,N_9823);
nor U11149 (N_11149,N_10091,N_10196);
or U11150 (N_11150,N_9963,N_9904);
or U11151 (N_11151,N_10099,N_10326);
or U11152 (N_11152,N_10427,N_10357);
or U11153 (N_11153,N_10187,N_10302);
or U11154 (N_11154,N_10315,N_9871);
nor U11155 (N_11155,N_9993,N_10096);
or U11156 (N_11156,N_10295,N_9945);
nand U11157 (N_11157,N_10009,N_9863);
xor U11158 (N_11158,N_10026,N_10082);
nand U11159 (N_11159,N_9883,N_9767);
nand U11160 (N_11160,N_10039,N_9849);
nand U11161 (N_11161,N_9910,N_10494);
nor U11162 (N_11162,N_10286,N_10488);
and U11163 (N_11163,N_9982,N_9786);
xnor U11164 (N_11164,N_10424,N_10142);
xor U11165 (N_11165,N_10165,N_9774);
and U11166 (N_11166,N_9895,N_10082);
or U11167 (N_11167,N_9828,N_10284);
nand U11168 (N_11168,N_10026,N_9968);
nor U11169 (N_11169,N_10428,N_10160);
nand U11170 (N_11170,N_10487,N_10174);
xor U11171 (N_11171,N_9845,N_10057);
or U11172 (N_11172,N_9877,N_10429);
or U11173 (N_11173,N_10460,N_9821);
or U11174 (N_11174,N_10198,N_10031);
xnor U11175 (N_11175,N_9873,N_10182);
nor U11176 (N_11176,N_9800,N_10155);
or U11177 (N_11177,N_10390,N_9877);
nand U11178 (N_11178,N_10031,N_9779);
nand U11179 (N_11179,N_10006,N_10451);
and U11180 (N_11180,N_10424,N_9978);
and U11181 (N_11181,N_10224,N_10164);
nand U11182 (N_11182,N_9791,N_10070);
or U11183 (N_11183,N_10385,N_9772);
nand U11184 (N_11184,N_10347,N_9941);
nand U11185 (N_11185,N_9918,N_10316);
nand U11186 (N_11186,N_10060,N_9793);
nand U11187 (N_11187,N_10072,N_10451);
nand U11188 (N_11188,N_10210,N_9754);
nand U11189 (N_11189,N_10425,N_10361);
nand U11190 (N_11190,N_10419,N_10372);
nor U11191 (N_11191,N_10291,N_9927);
nand U11192 (N_11192,N_9979,N_9957);
nor U11193 (N_11193,N_10472,N_9813);
nor U11194 (N_11194,N_10391,N_10045);
or U11195 (N_11195,N_10151,N_9922);
nand U11196 (N_11196,N_10497,N_9776);
and U11197 (N_11197,N_9785,N_10056);
and U11198 (N_11198,N_10432,N_10342);
xnor U11199 (N_11199,N_10453,N_10287);
nor U11200 (N_11200,N_9885,N_9801);
nor U11201 (N_11201,N_10242,N_10140);
nor U11202 (N_11202,N_9980,N_10465);
and U11203 (N_11203,N_10338,N_10043);
and U11204 (N_11204,N_9998,N_10252);
nor U11205 (N_11205,N_10325,N_10467);
nor U11206 (N_11206,N_9756,N_9934);
nand U11207 (N_11207,N_10496,N_9755);
xor U11208 (N_11208,N_10137,N_9992);
and U11209 (N_11209,N_10442,N_10388);
nor U11210 (N_11210,N_9800,N_10347);
nor U11211 (N_11211,N_9861,N_10211);
nand U11212 (N_11212,N_9798,N_9982);
or U11213 (N_11213,N_9817,N_10252);
nand U11214 (N_11214,N_9904,N_10063);
or U11215 (N_11215,N_9981,N_10003);
or U11216 (N_11216,N_9891,N_10367);
nand U11217 (N_11217,N_10374,N_10091);
nand U11218 (N_11218,N_9863,N_9761);
or U11219 (N_11219,N_10208,N_10455);
nor U11220 (N_11220,N_10159,N_9843);
nor U11221 (N_11221,N_9978,N_10081);
xor U11222 (N_11222,N_10287,N_10139);
and U11223 (N_11223,N_10354,N_9869);
and U11224 (N_11224,N_10040,N_10422);
xnor U11225 (N_11225,N_10174,N_10127);
nand U11226 (N_11226,N_10390,N_10119);
nor U11227 (N_11227,N_10075,N_10497);
nor U11228 (N_11228,N_9917,N_9933);
nor U11229 (N_11229,N_10168,N_10091);
and U11230 (N_11230,N_10402,N_10318);
or U11231 (N_11231,N_10296,N_10186);
and U11232 (N_11232,N_10457,N_10146);
nand U11233 (N_11233,N_10036,N_10280);
xnor U11234 (N_11234,N_10053,N_10404);
or U11235 (N_11235,N_10174,N_10323);
nor U11236 (N_11236,N_9846,N_9832);
or U11237 (N_11237,N_10158,N_10499);
nor U11238 (N_11238,N_10196,N_10463);
or U11239 (N_11239,N_10256,N_9969);
or U11240 (N_11240,N_10362,N_10249);
or U11241 (N_11241,N_10110,N_10266);
and U11242 (N_11242,N_10058,N_10247);
or U11243 (N_11243,N_9825,N_10007);
nor U11244 (N_11244,N_10013,N_10285);
nor U11245 (N_11245,N_10285,N_9827);
or U11246 (N_11246,N_10432,N_9869);
xnor U11247 (N_11247,N_10037,N_10255);
nand U11248 (N_11248,N_10238,N_9842);
and U11249 (N_11249,N_10010,N_10034);
xnor U11250 (N_11250,N_10706,N_11052);
and U11251 (N_11251,N_10520,N_10809);
nand U11252 (N_11252,N_10913,N_10892);
xor U11253 (N_11253,N_10941,N_10877);
and U11254 (N_11254,N_10678,N_11010);
and U11255 (N_11255,N_10810,N_11176);
or U11256 (N_11256,N_10690,N_11231);
or U11257 (N_11257,N_10987,N_10708);
or U11258 (N_11258,N_11186,N_11024);
and U11259 (N_11259,N_10766,N_10814);
and U11260 (N_11260,N_10560,N_10950);
or U11261 (N_11261,N_10540,N_11245);
nand U11262 (N_11262,N_10895,N_11153);
xor U11263 (N_11263,N_10837,N_11094);
nor U11264 (N_11264,N_11039,N_11148);
nand U11265 (N_11265,N_10923,N_10723);
and U11266 (N_11266,N_10805,N_10730);
or U11267 (N_11267,N_11003,N_10587);
nor U11268 (N_11268,N_10787,N_10506);
or U11269 (N_11269,N_10734,N_10769);
or U11270 (N_11270,N_10843,N_10953);
nor U11271 (N_11271,N_10544,N_10974);
and U11272 (N_11272,N_10686,N_10802);
xor U11273 (N_11273,N_10566,N_10516);
and U11274 (N_11274,N_11194,N_11184);
or U11275 (N_11275,N_10524,N_10561);
xor U11276 (N_11276,N_11041,N_11046);
and U11277 (N_11277,N_11142,N_11208);
and U11278 (N_11278,N_10590,N_11073);
or U11279 (N_11279,N_10732,N_11226);
nor U11280 (N_11280,N_10682,N_10920);
nor U11281 (N_11281,N_10806,N_11103);
xor U11282 (N_11282,N_11222,N_10530);
and U11283 (N_11283,N_11081,N_10937);
and U11284 (N_11284,N_11183,N_10922);
xnor U11285 (N_11285,N_10542,N_10977);
and U11286 (N_11286,N_11077,N_10967);
and U11287 (N_11287,N_10849,N_10755);
and U11288 (N_11288,N_11042,N_10826);
and U11289 (N_11289,N_11013,N_10729);
nor U11290 (N_11290,N_10654,N_11171);
nand U11291 (N_11291,N_10820,N_10903);
and U11292 (N_11292,N_10648,N_11174);
nor U11293 (N_11293,N_11150,N_11141);
nor U11294 (N_11294,N_10966,N_10889);
nand U11295 (N_11295,N_11197,N_10994);
and U11296 (N_11296,N_11137,N_10930);
nor U11297 (N_11297,N_10942,N_11213);
nand U11298 (N_11298,N_10633,N_11070);
xor U11299 (N_11299,N_11216,N_10675);
nor U11300 (N_11300,N_11240,N_10646);
xnor U11301 (N_11301,N_10608,N_10525);
nand U11302 (N_11302,N_10789,N_10502);
nand U11303 (N_11303,N_11045,N_10862);
nor U11304 (N_11304,N_11020,N_10927);
or U11305 (N_11305,N_10552,N_10905);
nor U11306 (N_11306,N_11212,N_10562);
and U11307 (N_11307,N_10881,N_10531);
and U11308 (N_11308,N_11018,N_11008);
and U11309 (N_11309,N_11078,N_11243);
nor U11310 (N_11310,N_10738,N_11029);
xnor U11311 (N_11311,N_11030,N_10796);
and U11312 (N_11312,N_11215,N_10649);
or U11313 (N_11313,N_10804,N_10836);
nand U11314 (N_11314,N_10722,N_10890);
xnor U11315 (N_11315,N_10572,N_11063);
nand U11316 (N_11316,N_11191,N_10824);
or U11317 (N_11317,N_11211,N_10639);
nor U11318 (N_11318,N_11207,N_11074);
and U11319 (N_11319,N_10749,N_10569);
and U11320 (N_11320,N_10545,N_10876);
and U11321 (N_11321,N_10832,N_10774);
nand U11322 (N_11322,N_10819,N_11056);
nor U11323 (N_11323,N_10564,N_10719);
nand U11324 (N_11324,N_10969,N_10860);
and U11325 (N_11325,N_10709,N_10598);
or U11326 (N_11326,N_10794,N_10713);
and U11327 (N_11327,N_10989,N_10674);
or U11328 (N_11328,N_11117,N_10586);
or U11329 (N_11329,N_11205,N_10912);
or U11330 (N_11330,N_10851,N_11085);
and U11331 (N_11331,N_10612,N_11169);
nor U11332 (N_11332,N_10760,N_11048);
xnor U11333 (N_11333,N_10632,N_10527);
nor U11334 (N_11334,N_10951,N_10956);
nand U11335 (N_11335,N_10500,N_10661);
nand U11336 (N_11336,N_10515,N_10813);
and U11337 (N_11337,N_10656,N_10743);
and U11338 (N_11338,N_10886,N_10720);
or U11339 (N_11339,N_10747,N_10899);
xor U11340 (N_11340,N_10990,N_11210);
and U11341 (N_11341,N_11120,N_11093);
and U11342 (N_11342,N_11027,N_10677);
and U11343 (N_11343,N_10961,N_11206);
nand U11344 (N_11344,N_10847,N_10750);
nand U11345 (N_11345,N_10915,N_11192);
or U11346 (N_11346,N_10988,N_10782);
nor U11347 (N_11347,N_10779,N_11004);
nand U11348 (N_11348,N_11170,N_10752);
or U11349 (N_11349,N_10935,N_10733);
and U11350 (N_11350,N_10635,N_10575);
or U11351 (N_11351,N_10807,N_10621);
nand U11352 (N_11352,N_11096,N_11097);
or U11353 (N_11353,N_10980,N_11202);
nor U11354 (N_11354,N_11116,N_10908);
nand U11355 (N_11355,N_10735,N_10762);
or U11356 (N_11356,N_11121,N_10916);
nor U11357 (N_11357,N_10968,N_11050);
and U11358 (N_11358,N_10725,N_11178);
nor U11359 (N_11359,N_11014,N_11007);
and U11360 (N_11360,N_10932,N_10781);
nor U11361 (N_11361,N_11083,N_10790);
nand U11362 (N_11362,N_10823,N_11036);
nor U11363 (N_11363,N_11165,N_10879);
and U11364 (N_11364,N_11034,N_10662);
nor U11365 (N_11365,N_10746,N_10551);
nor U11366 (N_11366,N_11238,N_10909);
and U11367 (N_11367,N_11055,N_10808);
and U11368 (N_11368,N_10817,N_11193);
nand U11369 (N_11369,N_10501,N_11017);
nor U11370 (N_11370,N_10775,N_10925);
nor U11371 (N_11371,N_10944,N_10883);
and U11372 (N_11372,N_10842,N_10865);
and U11373 (N_11373,N_11091,N_10534);
nand U11374 (N_11374,N_10548,N_10597);
xnor U11375 (N_11375,N_10803,N_10655);
nor U11376 (N_11376,N_11082,N_11175);
nand U11377 (N_11377,N_10900,N_10891);
or U11378 (N_11378,N_10670,N_10815);
nand U11379 (N_11379,N_10640,N_10873);
nor U11380 (N_11380,N_10882,N_11181);
and U11381 (N_11381,N_10739,N_11159);
nand U11382 (N_11382,N_10985,N_10791);
or U11383 (N_11383,N_10852,N_10767);
xor U11384 (N_11384,N_10504,N_11032);
nand U11385 (N_11385,N_10830,N_10973);
nand U11386 (N_11386,N_10991,N_10833);
nand U11387 (N_11387,N_10617,N_10550);
nand U11388 (N_11388,N_10519,N_10764);
nor U11389 (N_11389,N_10595,N_10602);
and U11390 (N_11390,N_11068,N_10904);
and U11391 (N_11391,N_10718,N_10650);
nor U11392 (N_11392,N_11227,N_10741);
nor U11393 (N_11393,N_11062,N_10695);
and U11394 (N_11394,N_10522,N_11025);
and U11395 (N_11395,N_11131,N_11187);
nand U11396 (N_11396,N_10858,N_10533);
and U11397 (N_11397,N_10600,N_10894);
nor U11398 (N_11398,N_11001,N_10939);
nand U11399 (N_11399,N_11233,N_11080);
or U11400 (N_11400,N_10982,N_10692);
nand U11401 (N_11401,N_11123,N_11006);
nor U11402 (N_11402,N_10714,N_10573);
or U11403 (N_11403,N_11016,N_11065);
or U11404 (N_11404,N_11180,N_11100);
nor U11405 (N_11405,N_10683,N_10924);
nand U11406 (N_11406,N_10971,N_10854);
or U11407 (N_11407,N_10710,N_10867);
and U11408 (N_11408,N_10715,N_11101);
or U11409 (N_11409,N_10517,N_10835);
xnor U11410 (N_11410,N_10963,N_10507);
nor U11411 (N_11411,N_10871,N_10954);
or U11412 (N_11412,N_10589,N_11000);
or U11413 (N_11413,N_10863,N_10699);
nor U11414 (N_11414,N_11110,N_10875);
xor U11415 (N_11415,N_10618,N_10556);
and U11416 (N_11416,N_10696,N_10606);
or U11417 (N_11417,N_10580,N_10671);
nand U11418 (N_11418,N_10605,N_10845);
or U11419 (N_11419,N_11196,N_10657);
nor U11420 (N_11420,N_10731,N_11067);
nor U11421 (N_11421,N_11071,N_11195);
nor U11422 (N_11422,N_11076,N_10770);
nand U11423 (N_11423,N_11015,N_11179);
nand U11424 (N_11424,N_10616,N_10869);
and U11425 (N_11425,N_10704,N_10840);
nand U11426 (N_11426,N_11095,N_10778);
and U11427 (N_11427,N_10570,N_11138);
xnor U11428 (N_11428,N_10740,N_10896);
and U11429 (N_11429,N_10970,N_10641);
nand U11430 (N_11430,N_11051,N_10513);
and U11431 (N_11431,N_11122,N_10693);
nand U11432 (N_11432,N_11220,N_10745);
nor U11433 (N_11433,N_10652,N_10582);
nor U11434 (N_11434,N_11209,N_10751);
and U11435 (N_11435,N_11249,N_10929);
nor U11436 (N_11436,N_10861,N_11054);
or U11437 (N_11437,N_10716,N_10559);
and U11438 (N_11438,N_10523,N_11201);
and U11439 (N_11439,N_10801,N_11158);
nand U11440 (N_11440,N_11133,N_10742);
xor U11441 (N_11441,N_10885,N_10567);
nand U11442 (N_11442,N_10642,N_10599);
nand U11443 (N_11443,N_11104,N_11084);
xor U11444 (N_11444,N_10689,N_10535);
and U11445 (N_11445,N_11087,N_10918);
or U11446 (N_11446,N_11102,N_11143);
or U11447 (N_11447,N_11037,N_11047);
nor U11448 (N_11448,N_10983,N_10630);
nand U11449 (N_11449,N_10888,N_10936);
nor U11450 (N_11450,N_10773,N_11185);
nor U11451 (N_11451,N_10962,N_10625);
nor U11452 (N_11452,N_11160,N_10651);
or U11453 (N_11453,N_10857,N_10958);
and U11454 (N_11454,N_10979,N_11058);
xnor U11455 (N_11455,N_10999,N_11075);
nand U11456 (N_11456,N_10822,N_10943);
or U11457 (N_11457,N_11228,N_10825);
nor U11458 (N_11458,N_10585,N_11011);
nor U11459 (N_11459,N_10995,N_10818);
nor U11460 (N_11460,N_10555,N_10947);
and U11461 (N_11461,N_10607,N_10754);
or U11462 (N_11462,N_10901,N_11188);
nand U11463 (N_11463,N_10549,N_11098);
and U11464 (N_11464,N_11089,N_10921);
or U11465 (N_11465,N_10902,N_10694);
nor U11466 (N_11466,N_10629,N_11200);
and U11467 (N_11467,N_10800,N_10672);
or U11468 (N_11468,N_10952,N_10557);
nor U11469 (N_11469,N_11079,N_11059);
and U11470 (N_11470,N_10705,N_11118);
nand U11471 (N_11471,N_11026,N_10978);
and U11472 (N_11472,N_10536,N_11247);
nand U11473 (N_11473,N_10872,N_10874);
nor U11474 (N_11474,N_10797,N_10508);
nand U11475 (N_11475,N_11119,N_11019);
nand U11476 (N_11476,N_10571,N_10634);
and U11477 (N_11477,N_11064,N_10996);
nor U11478 (N_11478,N_11111,N_11163);
nor U11479 (N_11479,N_10697,N_10702);
nand U11480 (N_11480,N_10631,N_10673);
nand U11481 (N_11481,N_10841,N_10821);
nand U11482 (N_11482,N_10509,N_10917);
nand U11483 (N_11483,N_10855,N_10563);
nand U11484 (N_11484,N_10931,N_10660);
nor U11485 (N_11485,N_11057,N_10676);
xnor U11486 (N_11486,N_10846,N_10853);
nand U11487 (N_11487,N_10898,N_10783);
nor U11488 (N_11488,N_11190,N_10510);
or U11489 (N_11489,N_10638,N_11198);
or U11490 (N_11490,N_10759,N_10761);
and U11491 (N_11491,N_11128,N_10701);
nor U11492 (N_11492,N_11232,N_10792);
nor U11493 (N_11493,N_11162,N_10757);
nand U11494 (N_11494,N_10707,N_10844);
nand U11495 (N_11495,N_10827,N_10763);
or U11496 (N_11496,N_10539,N_11225);
nand U11497 (N_11497,N_10780,N_10680);
or U11498 (N_11498,N_10583,N_11035);
nor U11499 (N_11499,N_11147,N_10964);
nand U11500 (N_11500,N_11132,N_11112);
and U11501 (N_11501,N_10647,N_10721);
nor U11502 (N_11502,N_10997,N_11236);
and U11503 (N_11503,N_10786,N_10645);
nor U11504 (N_11504,N_10604,N_11203);
nor U11505 (N_11505,N_10691,N_10665);
nor U11506 (N_11506,N_10960,N_10744);
nand U11507 (N_11507,N_11241,N_10636);
xor U11508 (N_11508,N_10518,N_10784);
nor U11509 (N_11509,N_10834,N_10793);
and U11510 (N_11510,N_10838,N_11224);
nor U11511 (N_11511,N_10788,N_11219);
and U11512 (N_11512,N_11105,N_10765);
and U11513 (N_11513,N_11152,N_10776);
nor U11514 (N_11514,N_10526,N_11234);
or U11515 (N_11515,N_10626,N_11099);
nand U11516 (N_11516,N_10588,N_10591);
nand U11517 (N_11517,N_10643,N_11177);
xnor U11518 (N_11518,N_10949,N_11139);
and U11519 (N_11519,N_10668,N_11109);
nand U11520 (N_11520,N_10965,N_10584);
and U11521 (N_11521,N_10868,N_11248);
nand U11522 (N_11522,N_11246,N_10611);
nand U11523 (N_11523,N_10541,N_10681);
or U11524 (N_11524,N_11135,N_10981);
and U11525 (N_11525,N_10798,N_11125);
nor U11526 (N_11526,N_10934,N_11028);
xor U11527 (N_11527,N_10957,N_11049);
xor U11528 (N_11528,N_10521,N_11217);
and U11529 (N_11529,N_10703,N_10603);
nand U11530 (N_11530,N_10887,N_11038);
nand U11531 (N_11531,N_11069,N_10712);
or U11532 (N_11532,N_10581,N_10659);
nor U11533 (N_11533,N_11229,N_11012);
nand U11534 (N_11534,N_10532,N_10622);
nand U11535 (N_11535,N_10687,N_10592);
or U11536 (N_11536,N_10717,N_10993);
and U11537 (N_11537,N_10593,N_10574);
and U11538 (N_11538,N_10777,N_10685);
nand U11539 (N_11539,N_11235,N_10679);
nor U11540 (N_11540,N_11072,N_10601);
xnor U11541 (N_11541,N_10620,N_10907);
nand U11542 (N_11542,N_10940,N_11140);
nor U11543 (N_11543,N_10812,N_10839);
xnor U11544 (N_11544,N_10724,N_11146);
or U11545 (N_11545,N_10623,N_10698);
nand U11546 (N_11546,N_11167,N_10537);
or U11547 (N_11547,N_11044,N_11066);
and U11548 (N_11548,N_10986,N_10768);
nor U11549 (N_11549,N_10528,N_11189);
nor U11550 (N_11550,N_11114,N_11033);
or U11551 (N_11551,N_10938,N_10554);
nand U11552 (N_11552,N_10700,N_10946);
and U11553 (N_11553,N_10848,N_10663);
and U11554 (N_11554,N_10864,N_10667);
nand U11555 (N_11555,N_10992,N_10906);
or U11556 (N_11556,N_10503,N_10831);
xnor U11557 (N_11557,N_10543,N_10850);
or U11558 (N_11558,N_10546,N_11136);
nand U11559 (N_11559,N_10911,N_10771);
xnor U11560 (N_11560,N_10558,N_10928);
xor U11561 (N_11561,N_11161,N_11134);
nand U11562 (N_11562,N_11144,N_10736);
nor U11563 (N_11563,N_10637,N_11124);
nand U11564 (N_11564,N_11221,N_10653);
or U11565 (N_11565,N_10547,N_11088);
nand U11566 (N_11566,N_10553,N_11155);
or U11567 (N_11567,N_10688,N_10785);
nand U11568 (N_11568,N_10975,N_11239);
and U11569 (N_11569,N_10666,N_10615);
or U11570 (N_11570,N_11108,N_10664);
and U11571 (N_11571,N_11151,N_11172);
nor U11572 (N_11572,N_11223,N_10933);
and U11573 (N_11573,N_10998,N_10511);
nand U11574 (N_11574,N_10758,N_10870);
or U11575 (N_11575,N_10514,N_11022);
nor U11576 (N_11576,N_10576,N_11053);
or U11577 (N_11577,N_10684,N_10737);
nor U11578 (N_11578,N_11145,N_10610);
or U11579 (N_11579,N_10945,N_11237);
xor U11580 (N_11580,N_10897,N_10753);
xnor U11581 (N_11581,N_11127,N_11061);
and U11582 (N_11582,N_10624,N_10972);
and U11583 (N_11583,N_10976,N_11090);
or U11584 (N_11584,N_10748,N_10578);
and U11585 (N_11585,N_10856,N_10596);
and U11586 (N_11586,N_11060,N_10505);
or U11587 (N_11587,N_10884,N_10594);
nor U11588 (N_11588,N_10538,N_10512);
nor U11589 (N_11589,N_11043,N_11157);
or U11590 (N_11590,N_10644,N_11002);
nor U11591 (N_11591,N_11021,N_11040);
or U11592 (N_11592,N_11107,N_10609);
xnor U11593 (N_11593,N_10955,N_10984);
nand U11594 (N_11594,N_11009,N_11115);
or U11595 (N_11595,N_11230,N_11204);
or U11596 (N_11596,N_10658,N_10628);
xnor U11597 (N_11597,N_10529,N_10959);
nand U11598 (N_11598,N_10568,N_10799);
or U11599 (N_11599,N_11156,N_10910);
and U11600 (N_11600,N_10811,N_10627);
nor U11601 (N_11601,N_10816,N_10795);
xnor U11602 (N_11602,N_10866,N_10613);
xnor U11603 (N_11603,N_11218,N_11130);
nor U11604 (N_11604,N_10893,N_11113);
or U11605 (N_11605,N_11106,N_11168);
nand U11606 (N_11606,N_11005,N_10711);
and U11607 (N_11607,N_11154,N_10914);
and U11608 (N_11608,N_10829,N_10919);
nand U11609 (N_11609,N_10577,N_11126);
nand U11610 (N_11610,N_11173,N_10828);
xor U11611 (N_11611,N_11166,N_10948);
nor U11612 (N_11612,N_10614,N_10727);
nand U11613 (N_11613,N_11031,N_11199);
nor U11614 (N_11614,N_11149,N_10726);
and U11615 (N_11615,N_10878,N_10669);
and U11616 (N_11616,N_10772,N_10579);
nand U11617 (N_11617,N_10565,N_11244);
nor U11618 (N_11618,N_11164,N_10859);
nor U11619 (N_11619,N_10619,N_10728);
and U11620 (N_11620,N_10926,N_11242);
nor U11621 (N_11621,N_10756,N_11092);
and U11622 (N_11622,N_11086,N_11129);
and U11623 (N_11623,N_10880,N_11182);
and U11624 (N_11624,N_11214,N_11023);
or U11625 (N_11625,N_10881,N_10723);
and U11626 (N_11626,N_10932,N_10884);
nor U11627 (N_11627,N_10812,N_10966);
or U11628 (N_11628,N_10663,N_10620);
nand U11629 (N_11629,N_11246,N_10721);
xnor U11630 (N_11630,N_10912,N_11196);
or U11631 (N_11631,N_11226,N_10716);
nor U11632 (N_11632,N_11034,N_10885);
or U11633 (N_11633,N_11221,N_10693);
xnor U11634 (N_11634,N_11062,N_10928);
nand U11635 (N_11635,N_10749,N_10975);
and U11636 (N_11636,N_11090,N_10917);
and U11637 (N_11637,N_10671,N_11022);
and U11638 (N_11638,N_11000,N_10671);
or U11639 (N_11639,N_10816,N_11177);
nand U11640 (N_11640,N_10722,N_10734);
nand U11641 (N_11641,N_10986,N_10822);
nand U11642 (N_11642,N_10725,N_10826);
nand U11643 (N_11643,N_10840,N_10712);
nor U11644 (N_11644,N_10717,N_10951);
and U11645 (N_11645,N_11035,N_11023);
or U11646 (N_11646,N_11124,N_10932);
nor U11647 (N_11647,N_10981,N_10524);
and U11648 (N_11648,N_11226,N_10557);
nand U11649 (N_11649,N_11220,N_10657);
and U11650 (N_11650,N_11051,N_11151);
and U11651 (N_11651,N_10765,N_11135);
nor U11652 (N_11652,N_10879,N_10839);
or U11653 (N_11653,N_11032,N_10625);
and U11654 (N_11654,N_11213,N_10558);
and U11655 (N_11655,N_11060,N_11151);
or U11656 (N_11656,N_11141,N_10647);
and U11657 (N_11657,N_10930,N_10850);
nor U11658 (N_11658,N_10728,N_10819);
and U11659 (N_11659,N_10702,N_11008);
nor U11660 (N_11660,N_11066,N_10975);
nand U11661 (N_11661,N_11183,N_10516);
xor U11662 (N_11662,N_10606,N_10632);
nand U11663 (N_11663,N_11223,N_10897);
or U11664 (N_11664,N_10710,N_11075);
or U11665 (N_11665,N_11083,N_10855);
or U11666 (N_11666,N_10555,N_11134);
and U11667 (N_11667,N_10584,N_11095);
nand U11668 (N_11668,N_11124,N_10602);
and U11669 (N_11669,N_11071,N_10831);
nor U11670 (N_11670,N_10651,N_11230);
nand U11671 (N_11671,N_11133,N_11241);
or U11672 (N_11672,N_11196,N_11219);
and U11673 (N_11673,N_10536,N_10516);
nand U11674 (N_11674,N_10811,N_11157);
nor U11675 (N_11675,N_10611,N_10761);
nor U11676 (N_11676,N_11015,N_10899);
nor U11677 (N_11677,N_11063,N_10647);
xor U11678 (N_11678,N_10614,N_10950);
nand U11679 (N_11679,N_10898,N_10841);
or U11680 (N_11680,N_10579,N_10789);
or U11681 (N_11681,N_10982,N_10807);
nand U11682 (N_11682,N_10748,N_10551);
and U11683 (N_11683,N_11141,N_10822);
or U11684 (N_11684,N_10512,N_10790);
or U11685 (N_11685,N_11145,N_10980);
and U11686 (N_11686,N_10742,N_11222);
nor U11687 (N_11687,N_10580,N_10573);
nor U11688 (N_11688,N_10616,N_10772);
or U11689 (N_11689,N_10741,N_10751);
or U11690 (N_11690,N_10589,N_10928);
and U11691 (N_11691,N_11107,N_10806);
xnor U11692 (N_11692,N_10595,N_10674);
nand U11693 (N_11693,N_11082,N_11081);
nand U11694 (N_11694,N_11035,N_10629);
and U11695 (N_11695,N_10559,N_10537);
xnor U11696 (N_11696,N_10795,N_11036);
or U11697 (N_11697,N_11207,N_10808);
or U11698 (N_11698,N_10996,N_10970);
nor U11699 (N_11699,N_10641,N_11038);
and U11700 (N_11700,N_10672,N_11092);
xor U11701 (N_11701,N_10855,N_10674);
nand U11702 (N_11702,N_10843,N_11179);
or U11703 (N_11703,N_11001,N_10689);
nand U11704 (N_11704,N_10901,N_10506);
or U11705 (N_11705,N_11125,N_10536);
nor U11706 (N_11706,N_10839,N_11221);
nor U11707 (N_11707,N_10731,N_11121);
nor U11708 (N_11708,N_10590,N_10513);
nand U11709 (N_11709,N_10726,N_11122);
nand U11710 (N_11710,N_11054,N_10528);
nor U11711 (N_11711,N_10663,N_11211);
or U11712 (N_11712,N_10660,N_10515);
or U11713 (N_11713,N_10955,N_10700);
nand U11714 (N_11714,N_10986,N_11024);
nand U11715 (N_11715,N_10785,N_11019);
nand U11716 (N_11716,N_10579,N_10982);
xnor U11717 (N_11717,N_10543,N_10548);
or U11718 (N_11718,N_10548,N_11235);
nand U11719 (N_11719,N_11138,N_10962);
or U11720 (N_11720,N_11156,N_11082);
and U11721 (N_11721,N_11227,N_11189);
and U11722 (N_11722,N_11220,N_10795);
nor U11723 (N_11723,N_10623,N_11244);
and U11724 (N_11724,N_10584,N_10591);
or U11725 (N_11725,N_10732,N_10595);
nand U11726 (N_11726,N_10883,N_10985);
and U11727 (N_11727,N_10566,N_11201);
and U11728 (N_11728,N_10701,N_10828);
and U11729 (N_11729,N_10712,N_10677);
or U11730 (N_11730,N_10606,N_10964);
or U11731 (N_11731,N_11219,N_10686);
nor U11732 (N_11732,N_10869,N_11134);
and U11733 (N_11733,N_10932,N_11141);
or U11734 (N_11734,N_10826,N_11051);
nor U11735 (N_11735,N_10561,N_10882);
nand U11736 (N_11736,N_10503,N_10825);
nand U11737 (N_11737,N_11110,N_10513);
or U11738 (N_11738,N_11027,N_10705);
or U11739 (N_11739,N_10934,N_10636);
xor U11740 (N_11740,N_10506,N_11244);
and U11741 (N_11741,N_10615,N_10604);
and U11742 (N_11742,N_10559,N_10915);
and U11743 (N_11743,N_10745,N_10916);
nor U11744 (N_11744,N_11114,N_11191);
nor U11745 (N_11745,N_10869,N_10626);
xor U11746 (N_11746,N_11156,N_10837);
and U11747 (N_11747,N_10967,N_10958);
nor U11748 (N_11748,N_10691,N_11114);
or U11749 (N_11749,N_10540,N_11111);
nor U11750 (N_11750,N_11070,N_11094);
or U11751 (N_11751,N_11175,N_11135);
and U11752 (N_11752,N_11228,N_10816);
and U11753 (N_11753,N_10615,N_11175);
or U11754 (N_11754,N_10569,N_10991);
nand U11755 (N_11755,N_11225,N_10918);
and U11756 (N_11756,N_10675,N_10915);
or U11757 (N_11757,N_10641,N_10567);
and U11758 (N_11758,N_10969,N_10832);
nor U11759 (N_11759,N_10700,N_11079);
nor U11760 (N_11760,N_10738,N_10761);
nor U11761 (N_11761,N_11145,N_10845);
xor U11762 (N_11762,N_10625,N_10830);
and U11763 (N_11763,N_10816,N_10932);
nand U11764 (N_11764,N_10561,N_11230);
and U11765 (N_11765,N_10533,N_10686);
and U11766 (N_11766,N_10609,N_10694);
nand U11767 (N_11767,N_11111,N_10619);
or U11768 (N_11768,N_11075,N_11008);
or U11769 (N_11769,N_11125,N_10793);
and U11770 (N_11770,N_10609,N_11014);
and U11771 (N_11771,N_10855,N_10870);
or U11772 (N_11772,N_11125,N_10585);
nor U11773 (N_11773,N_11091,N_11226);
xor U11774 (N_11774,N_10984,N_11152);
nor U11775 (N_11775,N_10711,N_11230);
and U11776 (N_11776,N_11202,N_10854);
nor U11777 (N_11777,N_10926,N_10875);
or U11778 (N_11778,N_11029,N_11023);
and U11779 (N_11779,N_10971,N_11193);
or U11780 (N_11780,N_10989,N_10942);
and U11781 (N_11781,N_10819,N_10778);
nor U11782 (N_11782,N_10515,N_11136);
nor U11783 (N_11783,N_10945,N_11179);
nand U11784 (N_11784,N_10689,N_11245);
nand U11785 (N_11785,N_11143,N_11089);
and U11786 (N_11786,N_10910,N_11221);
nand U11787 (N_11787,N_10556,N_10691);
nand U11788 (N_11788,N_10885,N_10804);
and U11789 (N_11789,N_11157,N_10603);
nand U11790 (N_11790,N_10963,N_10893);
or U11791 (N_11791,N_11197,N_10958);
nor U11792 (N_11792,N_11244,N_11223);
or U11793 (N_11793,N_11090,N_10860);
or U11794 (N_11794,N_10897,N_10540);
and U11795 (N_11795,N_10611,N_10618);
and U11796 (N_11796,N_11068,N_11234);
nor U11797 (N_11797,N_10981,N_10535);
nand U11798 (N_11798,N_10643,N_10750);
and U11799 (N_11799,N_11100,N_10793);
xor U11800 (N_11800,N_10563,N_10734);
and U11801 (N_11801,N_10812,N_10550);
nand U11802 (N_11802,N_10837,N_11121);
nor U11803 (N_11803,N_10919,N_10879);
xnor U11804 (N_11804,N_10840,N_10783);
or U11805 (N_11805,N_11083,N_10979);
or U11806 (N_11806,N_10895,N_10715);
or U11807 (N_11807,N_11186,N_10800);
or U11808 (N_11808,N_11009,N_10526);
or U11809 (N_11809,N_10614,N_11063);
and U11810 (N_11810,N_10851,N_10797);
nor U11811 (N_11811,N_11119,N_11018);
nand U11812 (N_11812,N_10795,N_10639);
or U11813 (N_11813,N_11021,N_10786);
nand U11814 (N_11814,N_11171,N_11164);
nand U11815 (N_11815,N_11158,N_10691);
nor U11816 (N_11816,N_11007,N_11214);
xor U11817 (N_11817,N_10931,N_10732);
or U11818 (N_11818,N_10896,N_10763);
or U11819 (N_11819,N_10530,N_10532);
nor U11820 (N_11820,N_10784,N_11096);
or U11821 (N_11821,N_10790,N_11087);
and U11822 (N_11822,N_11058,N_10640);
and U11823 (N_11823,N_10987,N_11037);
nand U11824 (N_11824,N_10922,N_10587);
nor U11825 (N_11825,N_11010,N_10624);
or U11826 (N_11826,N_11027,N_10862);
nand U11827 (N_11827,N_10724,N_10653);
and U11828 (N_11828,N_11207,N_10788);
nor U11829 (N_11829,N_10581,N_10744);
and U11830 (N_11830,N_10801,N_11174);
and U11831 (N_11831,N_10666,N_10715);
nand U11832 (N_11832,N_10993,N_11032);
or U11833 (N_11833,N_11201,N_10600);
or U11834 (N_11834,N_10526,N_11245);
and U11835 (N_11835,N_10613,N_10907);
and U11836 (N_11836,N_10736,N_10742);
and U11837 (N_11837,N_11016,N_10786);
and U11838 (N_11838,N_10799,N_11201);
or U11839 (N_11839,N_11128,N_10637);
xor U11840 (N_11840,N_10974,N_10731);
and U11841 (N_11841,N_10675,N_11174);
nand U11842 (N_11842,N_11155,N_10799);
or U11843 (N_11843,N_11016,N_10975);
and U11844 (N_11844,N_10773,N_10926);
nand U11845 (N_11845,N_11191,N_10592);
or U11846 (N_11846,N_11105,N_10796);
and U11847 (N_11847,N_10524,N_11011);
nor U11848 (N_11848,N_10608,N_11036);
or U11849 (N_11849,N_10566,N_11134);
or U11850 (N_11850,N_10644,N_10659);
or U11851 (N_11851,N_11180,N_10746);
nand U11852 (N_11852,N_10554,N_11095);
nand U11853 (N_11853,N_11192,N_11002);
or U11854 (N_11854,N_10938,N_10827);
nor U11855 (N_11855,N_10502,N_11238);
or U11856 (N_11856,N_10558,N_10961);
xor U11857 (N_11857,N_10788,N_10931);
xor U11858 (N_11858,N_10508,N_10620);
nor U11859 (N_11859,N_10937,N_10842);
or U11860 (N_11860,N_10528,N_10947);
nor U11861 (N_11861,N_11212,N_10904);
or U11862 (N_11862,N_10911,N_10999);
nor U11863 (N_11863,N_10581,N_11135);
xor U11864 (N_11864,N_10637,N_11040);
nor U11865 (N_11865,N_11148,N_10597);
or U11866 (N_11866,N_10980,N_10969);
or U11867 (N_11867,N_10695,N_10930);
nor U11868 (N_11868,N_10500,N_10572);
and U11869 (N_11869,N_10896,N_10578);
nor U11870 (N_11870,N_10678,N_10842);
or U11871 (N_11871,N_10513,N_10646);
nor U11872 (N_11872,N_10707,N_11194);
and U11873 (N_11873,N_10749,N_10523);
xnor U11874 (N_11874,N_10707,N_11015);
nand U11875 (N_11875,N_11229,N_11142);
and U11876 (N_11876,N_11052,N_10661);
and U11877 (N_11877,N_10526,N_11073);
or U11878 (N_11878,N_10951,N_10705);
nand U11879 (N_11879,N_11122,N_10751);
nand U11880 (N_11880,N_10922,N_11241);
xnor U11881 (N_11881,N_10528,N_11079);
nand U11882 (N_11882,N_10689,N_10691);
and U11883 (N_11883,N_10743,N_11166);
xor U11884 (N_11884,N_10511,N_10912);
xor U11885 (N_11885,N_10609,N_10935);
xnor U11886 (N_11886,N_11101,N_10938);
nand U11887 (N_11887,N_10570,N_10665);
or U11888 (N_11888,N_10620,N_10512);
nand U11889 (N_11889,N_11111,N_10609);
nor U11890 (N_11890,N_10921,N_10872);
or U11891 (N_11891,N_10626,N_10910);
nand U11892 (N_11892,N_11170,N_11223);
nand U11893 (N_11893,N_10877,N_10778);
and U11894 (N_11894,N_10809,N_11234);
and U11895 (N_11895,N_10622,N_10872);
xor U11896 (N_11896,N_10989,N_11016);
and U11897 (N_11897,N_11148,N_10829);
nor U11898 (N_11898,N_10767,N_11145);
nand U11899 (N_11899,N_11031,N_10723);
nor U11900 (N_11900,N_10788,N_11185);
or U11901 (N_11901,N_10627,N_11192);
and U11902 (N_11902,N_10669,N_10851);
or U11903 (N_11903,N_10927,N_10783);
nor U11904 (N_11904,N_11155,N_10838);
or U11905 (N_11905,N_11227,N_10884);
nor U11906 (N_11906,N_11136,N_10815);
nand U11907 (N_11907,N_10622,N_11165);
or U11908 (N_11908,N_11041,N_10789);
nand U11909 (N_11909,N_10940,N_11024);
nand U11910 (N_11910,N_10633,N_11098);
or U11911 (N_11911,N_10557,N_11180);
nor U11912 (N_11912,N_11030,N_10525);
and U11913 (N_11913,N_11137,N_11097);
nand U11914 (N_11914,N_11007,N_10751);
nor U11915 (N_11915,N_10977,N_10664);
or U11916 (N_11916,N_10643,N_10696);
nor U11917 (N_11917,N_10588,N_10521);
xor U11918 (N_11918,N_10821,N_10559);
and U11919 (N_11919,N_11070,N_10506);
and U11920 (N_11920,N_10716,N_10980);
and U11921 (N_11921,N_11168,N_10622);
xnor U11922 (N_11922,N_11173,N_10503);
or U11923 (N_11923,N_10870,N_10922);
nor U11924 (N_11924,N_10915,N_11238);
nand U11925 (N_11925,N_11115,N_10717);
xnor U11926 (N_11926,N_11033,N_10957);
or U11927 (N_11927,N_10658,N_11125);
and U11928 (N_11928,N_10549,N_10595);
xor U11929 (N_11929,N_11219,N_10786);
nor U11930 (N_11930,N_11091,N_11148);
and U11931 (N_11931,N_10997,N_10768);
and U11932 (N_11932,N_10749,N_11056);
nand U11933 (N_11933,N_11073,N_10620);
nor U11934 (N_11934,N_10636,N_10945);
and U11935 (N_11935,N_10707,N_10942);
nand U11936 (N_11936,N_10863,N_10644);
or U11937 (N_11937,N_10664,N_10817);
nand U11938 (N_11938,N_11155,N_11039);
nand U11939 (N_11939,N_10813,N_10666);
xnor U11940 (N_11940,N_10789,N_11000);
nor U11941 (N_11941,N_11139,N_10985);
xnor U11942 (N_11942,N_10873,N_10955);
and U11943 (N_11943,N_10579,N_10736);
and U11944 (N_11944,N_10822,N_10501);
xor U11945 (N_11945,N_10766,N_10784);
or U11946 (N_11946,N_10506,N_11204);
nor U11947 (N_11947,N_10559,N_11243);
nor U11948 (N_11948,N_10543,N_11002);
and U11949 (N_11949,N_10537,N_11092);
nand U11950 (N_11950,N_10805,N_10953);
nand U11951 (N_11951,N_10707,N_11133);
xor U11952 (N_11952,N_10961,N_10593);
nor U11953 (N_11953,N_10882,N_10610);
and U11954 (N_11954,N_10576,N_11008);
and U11955 (N_11955,N_10907,N_11192);
or U11956 (N_11956,N_10524,N_11034);
nor U11957 (N_11957,N_11239,N_10884);
and U11958 (N_11958,N_10918,N_10814);
nand U11959 (N_11959,N_11206,N_10855);
xor U11960 (N_11960,N_10916,N_10752);
xor U11961 (N_11961,N_10946,N_11084);
nand U11962 (N_11962,N_10865,N_10924);
and U11963 (N_11963,N_10599,N_10591);
nor U11964 (N_11964,N_10705,N_11147);
nand U11965 (N_11965,N_11238,N_11115);
and U11966 (N_11966,N_10698,N_11063);
xor U11967 (N_11967,N_11015,N_11120);
and U11968 (N_11968,N_10920,N_10864);
nor U11969 (N_11969,N_11166,N_10543);
and U11970 (N_11970,N_11164,N_11119);
and U11971 (N_11971,N_10729,N_10590);
nand U11972 (N_11972,N_10811,N_10582);
nor U11973 (N_11973,N_11150,N_11095);
xor U11974 (N_11974,N_11006,N_11130);
or U11975 (N_11975,N_11078,N_10810);
nand U11976 (N_11976,N_10871,N_11197);
nor U11977 (N_11977,N_10792,N_10772);
nor U11978 (N_11978,N_10707,N_10909);
nor U11979 (N_11979,N_10648,N_11041);
and U11980 (N_11980,N_10891,N_10507);
and U11981 (N_11981,N_10574,N_10921);
xnor U11982 (N_11982,N_10917,N_10582);
or U11983 (N_11983,N_10757,N_11012);
nand U11984 (N_11984,N_10959,N_10676);
and U11985 (N_11985,N_10764,N_10993);
and U11986 (N_11986,N_11112,N_10927);
or U11987 (N_11987,N_10583,N_10705);
nand U11988 (N_11988,N_10962,N_10612);
nor U11989 (N_11989,N_10677,N_10791);
nand U11990 (N_11990,N_10704,N_10527);
or U11991 (N_11991,N_11061,N_10920);
xor U11992 (N_11992,N_10775,N_10518);
nor U11993 (N_11993,N_10569,N_10523);
nand U11994 (N_11994,N_10917,N_10561);
nand U11995 (N_11995,N_11063,N_10660);
nor U11996 (N_11996,N_11208,N_10535);
or U11997 (N_11997,N_11206,N_11030);
and U11998 (N_11998,N_10561,N_11179);
or U11999 (N_11999,N_11165,N_10732);
xor U12000 (N_12000,N_11487,N_11281);
nor U12001 (N_12001,N_11714,N_11637);
and U12002 (N_12002,N_11944,N_11343);
nor U12003 (N_12003,N_11521,N_11638);
and U12004 (N_12004,N_11653,N_11333);
nor U12005 (N_12005,N_11518,N_11650);
and U12006 (N_12006,N_11728,N_11666);
nand U12007 (N_12007,N_11363,N_11270);
nand U12008 (N_12008,N_11615,N_11957);
nand U12009 (N_12009,N_11599,N_11265);
or U12010 (N_12010,N_11389,N_11764);
xor U12011 (N_12011,N_11842,N_11847);
and U12012 (N_12012,N_11353,N_11466);
or U12013 (N_12013,N_11706,N_11324);
nand U12014 (N_12014,N_11880,N_11507);
nor U12015 (N_12015,N_11545,N_11815);
nand U12016 (N_12016,N_11556,N_11554);
and U12017 (N_12017,N_11962,N_11705);
or U12018 (N_12018,N_11347,N_11330);
or U12019 (N_12019,N_11544,N_11422);
or U12020 (N_12020,N_11332,N_11374);
and U12021 (N_12021,N_11503,N_11611);
or U12022 (N_12022,N_11369,N_11617);
nor U12023 (N_12023,N_11255,N_11793);
nor U12024 (N_12024,N_11529,N_11651);
or U12025 (N_12025,N_11965,N_11497);
nor U12026 (N_12026,N_11568,N_11350);
nand U12027 (N_12027,N_11751,N_11375);
or U12028 (N_12028,N_11734,N_11627);
and U12029 (N_12029,N_11822,N_11912);
nor U12030 (N_12030,N_11681,N_11535);
nor U12031 (N_12031,N_11614,N_11571);
nor U12032 (N_12032,N_11893,N_11885);
nor U12033 (N_12033,N_11724,N_11876);
nor U12034 (N_12034,N_11258,N_11726);
nor U12035 (N_12035,N_11501,N_11426);
nor U12036 (N_12036,N_11383,N_11881);
and U12037 (N_12037,N_11536,N_11361);
and U12038 (N_12038,N_11538,N_11763);
or U12039 (N_12039,N_11262,N_11452);
or U12040 (N_12040,N_11486,N_11421);
xnor U12041 (N_12041,N_11618,N_11778);
nor U12042 (N_12042,N_11700,N_11622);
nand U12043 (N_12043,N_11686,N_11799);
nand U12044 (N_12044,N_11874,N_11780);
and U12045 (N_12045,N_11668,N_11745);
nand U12046 (N_12046,N_11587,N_11316);
or U12047 (N_12047,N_11604,N_11621);
and U12048 (N_12048,N_11581,N_11657);
nand U12049 (N_12049,N_11448,N_11307);
xnor U12050 (N_12050,N_11566,N_11288);
nor U12051 (N_12051,N_11929,N_11387);
or U12052 (N_12052,N_11643,N_11534);
or U12053 (N_12053,N_11349,N_11373);
nand U12054 (N_12054,N_11266,N_11377);
nor U12055 (N_12055,N_11738,N_11868);
and U12056 (N_12056,N_11319,N_11983);
and U12057 (N_12057,N_11510,N_11453);
xor U12058 (N_12058,N_11985,N_11355);
and U12059 (N_12059,N_11570,N_11256);
nand U12060 (N_12060,N_11574,N_11987);
and U12061 (N_12061,N_11539,N_11703);
and U12062 (N_12062,N_11612,N_11443);
and U12063 (N_12063,N_11998,N_11312);
nor U12064 (N_12064,N_11963,N_11419);
or U12065 (N_12065,N_11935,N_11743);
nand U12066 (N_12066,N_11855,N_11625);
or U12067 (N_12067,N_11903,N_11514);
nor U12068 (N_12068,N_11294,N_11829);
or U12069 (N_12069,N_11445,N_11372);
nor U12070 (N_12070,N_11284,N_11424);
or U12071 (N_12071,N_11508,N_11517);
xnor U12072 (N_12072,N_11459,N_11844);
xnor U12073 (N_12073,N_11827,N_11646);
and U12074 (N_12074,N_11435,N_11908);
and U12075 (N_12075,N_11687,N_11400);
and U12076 (N_12076,N_11674,N_11575);
and U12077 (N_12077,N_11818,N_11950);
nor U12078 (N_12078,N_11729,N_11490);
and U12079 (N_12079,N_11433,N_11794);
nor U12080 (N_12080,N_11557,N_11406);
nor U12081 (N_12081,N_11329,N_11562);
nand U12082 (N_12082,N_11933,N_11992);
nor U12083 (N_12083,N_11852,N_11592);
xor U12084 (N_12084,N_11783,N_11781);
nor U12085 (N_12085,N_11250,N_11341);
nor U12086 (N_12086,N_11327,N_11541);
xnor U12087 (N_12087,N_11840,N_11259);
or U12088 (N_12088,N_11528,N_11593);
and U12089 (N_12089,N_11600,N_11469);
and U12090 (N_12090,N_11252,N_11941);
or U12091 (N_12091,N_11440,N_11782);
nand U12092 (N_12092,N_11792,N_11302);
and U12093 (N_12093,N_11549,N_11836);
xnor U12094 (N_12094,N_11320,N_11475);
or U12095 (N_12095,N_11340,N_11770);
nand U12096 (N_12096,N_11923,N_11834);
nor U12097 (N_12097,N_11974,N_11429);
and U12098 (N_12098,N_11491,N_11506);
nand U12099 (N_12099,N_11613,N_11665);
nor U12100 (N_12100,N_11947,N_11851);
xor U12101 (N_12101,N_11482,N_11366);
and U12102 (N_12102,N_11537,N_11591);
and U12103 (N_12103,N_11584,N_11555);
or U12104 (N_12104,N_11640,N_11279);
nand U12105 (N_12105,N_11495,N_11552);
nand U12106 (N_12106,N_11848,N_11449);
nor U12107 (N_12107,N_11451,N_11427);
nand U12108 (N_12108,N_11344,N_11439);
and U12109 (N_12109,N_11411,N_11291);
and U12110 (N_12110,N_11919,N_11716);
nor U12111 (N_12111,N_11471,N_11454);
nand U12112 (N_12112,N_11282,N_11606);
xnor U12113 (N_12113,N_11395,N_11689);
nor U12114 (N_12114,N_11733,N_11649);
nand U12115 (N_12115,N_11582,N_11278);
nor U12116 (N_12116,N_11835,N_11367);
nor U12117 (N_12117,N_11602,N_11845);
and U12118 (N_12118,N_11945,N_11958);
nor U12119 (N_12119,N_11773,N_11772);
nand U12120 (N_12120,N_11317,N_11889);
nand U12121 (N_12121,N_11695,N_11629);
nor U12122 (N_12122,N_11523,N_11253);
nand U12123 (N_12123,N_11636,N_11870);
nand U12124 (N_12124,N_11678,N_11838);
xor U12125 (N_12125,N_11871,N_11386);
and U12126 (N_12126,N_11837,N_11295);
and U12127 (N_12127,N_11345,N_11989);
and U12128 (N_12128,N_11590,N_11318);
nor U12129 (N_12129,N_11438,N_11820);
xnor U12130 (N_12130,N_11644,N_11280);
nand U12131 (N_12131,N_11371,N_11902);
or U12132 (N_12132,N_11900,N_11548);
or U12133 (N_12133,N_11308,N_11381);
nand U12134 (N_12134,N_11789,N_11420);
nor U12135 (N_12135,N_11767,N_11458);
and U12136 (N_12136,N_11942,N_11964);
and U12137 (N_12137,N_11303,N_11786);
or U12138 (N_12138,N_11765,N_11718);
and U12139 (N_12139,N_11856,N_11342);
nor U12140 (N_12140,N_11825,N_11608);
nand U12141 (N_12141,N_11493,N_11533);
xnor U12142 (N_12142,N_11583,N_11785);
nor U12143 (N_12143,N_11735,N_11645);
and U12144 (N_12144,N_11939,N_11499);
or U12145 (N_12145,N_11354,N_11271);
nand U12146 (N_12146,N_11699,N_11661);
nand U12147 (N_12147,N_11547,N_11403);
nand U12148 (N_12148,N_11470,N_11955);
and U12149 (N_12149,N_11742,N_11525);
nand U12150 (N_12150,N_11833,N_11887);
or U12151 (N_12151,N_11810,N_11410);
nor U12152 (N_12152,N_11791,N_11727);
and U12153 (N_12153,N_11670,N_11702);
nor U12154 (N_12154,N_11531,N_11559);
and U12155 (N_12155,N_11346,N_11790);
nor U12156 (N_12156,N_11685,N_11601);
and U12157 (N_12157,N_11384,N_11623);
or U12158 (N_12158,N_11580,N_11257);
or U12159 (N_12159,N_11550,N_11981);
nand U12160 (N_12160,N_11652,N_11796);
or U12161 (N_12161,N_11988,N_11682);
nor U12162 (N_12162,N_11362,N_11512);
nor U12163 (N_12163,N_11949,N_11511);
xnor U12164 (N_12164,N_11722,N_11904);
or U12165 (N_12165,N_11694,N_11779);
and U12166 (N_12166,N_11832,N_11416);
nand U12167 (N_12167,N_11709,N_11717);
nand U12168 (N_12168,N_11866,N_11978);
or U12169 (N_12169,N_11680,N_11474);
and U12170 (N_12170,N_11816,N_11991);
nand U12171 (N_12171,N_11739,N_11274);
and U12172 (N_12172,N_11817,N_11428);
and U12173 (N_12173,N_11951,N_11489);
or U12174 (N_12174,N_11788,N_11920);
nor U12175 (N_12175,N_11806,N_11673);
or U12176 (N_12176,N_11313,N_11698);
xnor U12177 (N_12177,N_11500,N_11758);
and U12178 (N_12178,N_11732,N_11973);
nand U12179 (N_12179,N_11461,N_11276);
or U12180 (N_12180,N_11711,N_11522);
or U12181 (N_12181,N_11289,N_11701);
or U12182 (N_12182,N_11605,N_11563);
or U12183 (N_12183,N_11328,N_11922);
nand U12184 (N_12184,N_11692,N_11721);
or U12185 (N_12185,N_11567,N_11946);
nand U12186 (N_12186,N_11737,N_11543);
nand U12187 (N_12187,N_11392,N_11479);
nor U12188 (N_12188,N_11823,N_11578);
nor U12189 (N_12189,N_11663,N_11667);
and U12190 (N_12190,N_11476,N_11325);
nand U12191 (N_12191,N_11860,N_11331);
nor U12192 (N_12192,N_11713,N_11560);
nor U12193 (N_12193,N_11814,N_11664);
and U12194 (N_12194,N_11909,N_11824);
and U12195 (N_12195,N_11768,N_11296);
nor U12196 (N_12196,N_11924,N_11736);
and U12197 (N_12197,N_11975,N_11913);
nand U12198 (N_12198,N_11509,N_11251);
xnor U12199 (N_12199,N_11630,N_11805);
nor U12200 (N_12200,N_11391,N_11843);
or U12201 (N_12201,N_11378,N_11390);
or U12202 (N_12202,N_11432,N_11565);
and U12203 (N_12203,N_11821,N_11831);
or U12204 (N_12204,N_11969,N_11869);
and U12205 (N_12205,N_11937,N_11633);
and U12206 (N_12206,N_11393,N_11430);
nor U12207 (N_12207,N_11610,N_11936);
or U12208 (N_12208,N_11812,N_11408);
or U12209 (N_12209,N_11754,N_11967);
nor U12210 (N_12210,N_11468,N_11485);
nor U12211 (N_12211,N_11323,N_11305);
nand U12212 (N_12212,N_11994,N_11952);
nand U12213 (N_12213,N_11804,N_11660);
nand U12214 (N_12214,N_11360,N_11777);
or U12215 (N_12215,N_11997,N_11890);
and U12216 (N_12216,N_11561,N_11388);
or U12217 (N_12217,N_11865,N_11530);
and U12218 (N_12218,N_11596,N_11862);
and U12219 (N_12219,N_11572,N_11607);
nor U12220 (N_12220,N_11480,N_11684);
and U12221 (N_12221,N_11504,N_11588);
nand U12222 (N_12222,N_11888,N_11293);
xnor U12223 (N_12223,N_11899,N_11586);
nor U12224 (N_12224,N_11413,N_11409);
and U12225 (N_12225,N_11286,N_11376);
nand U12226 (N_12226,N_11897,N_11905);
xor U12227 (N_12227,N_11442,N_11656);
or U12228 (N_12228,N_11441,N_11697);
and U12229 (N_12229,N_11641,N_11415);
and U12230 (N_12230,N_11690,N_11287);
nor U12231 (N_12231,N_11766,N_11402);
nor U12232 (N_12232,N_11297,N_11423);
and U12233 (N_12233,N_11598,N_11960);
or U12234 (N_12234,N_11272,N_11401);
nor U12235 (N_12235,N_11339,N_11634);
or U12236 (N_12236,N_11999,N_11961);
xor U12237 (N_12237,N_11846,N_11589);
or U12238 (N_12238,N_11524,N_11996);
nand U12239 (N_12239,N_11731,N_11811);
and U12240 (N_12240,N_11879,N_11669);
nand U12241 (N_12241,N_11954,N_11917);
xor U12242 (N_12242,N_11655,N_11750);
or U12243 (N_12243,N_11801,N_11292);
nand U12244 (N_12244,N_11986,N_11380);
nand U12245 (N_12245,N_11407,N_11273);
xor U12246 (N_12246,N_11725,N_11425);
nand U12247 (N_12247,N_11826,N_11337);
nor U12248 (N_12248,N_11787,N_11465);
or U12249 (N_12249,N_11322,N_11382);
nor U12250 (N_12250,N_11857,N_11910);
and U12251 (N_12251,N_11762,N_11693);
nand U12252 (N_12252,N_11417,N_11784);
nand U12253 (N_12253,N_11966,N_11564);
nor U12254 (N_12254,N_11894,N_11677);
nor U12255 (N_12255,N_11456,N_11730);
and U12256 (N_12256,N_11595,N_11551);
or U12257 (N_12257,N_11311,N_11396);
or U12258 (N_12258,N_11746,N_11911);
nor U12259 (N_12259,N_11774,N_11603);
nor U12260 (N_12260,N_11467,N_11620);
or U12261 (N_12261,N_11414,N_11940);
nand U12262 (N_12262,N_11895,N_11352);
nor U12263 (N_12263,N_11853,N_11309);
nand U12264 (N_12264,N_11741,N_11267);
xor U12265 (N_12265,N_11654,N_11970);
and U12266 (N_12266,N_11723,N_11502);
nor U12267 (N_12267,N_11671,N_11505);
nor U12268 (N_12268,N_11368,N_11850);
and U12269 (N_12269,N_11385,N_11484);
nor U12270 (N_12270,N_11310,N_11577);
or U12271 (N_12271,N_11481,N_11304);
nor U12272 (N_12272,N_11397,N_11553);
nand U12273 (N_12273,N_11932,N_11800);
nor U12274 (N_12274,N_11631,N_11884);
or U12275 (N_12275,N_11283,N_11761);
nor U12276 (N_12276,N_11984,N_11807);
nor U12277 (N_12277,N_11968,N_11878);
or U12278 (N_12278,N_11464,N_11264);
or U12279 (N_12279,N_11624,N_11849);
nand U12280 (N_12280,N_11639,N_11976);
or U12281 (N_12281,N_11478,N_11956);
nor U12282 (N_12282,N_11915,N_11290);
nand U12283 (N_12283,N_11616,N_11628);
nor U12284 (N_12284,N_11990,N_11863);
or U12285 (N_12285,N_11841,N_11861);
nand U12286 (N_12286,N_11455,N_11626);
or U12287 (N_12287,N_11254,N_11472);
and U12288 (N_12288,N_11516,N_11594);
and U12289 (N_12289,N_11927,N_11883);
nor U12290 (N_12290,N_11275,N_11707);
and U12291 (N_12291,N_11527,N_11546);
xor U12292 (N_12292,N_11365,N_11398);
and U12293 (N_12293,N_11569,N_11914);
and U12294 (N_12294,N_11326,N_11519);
nand U12295 (N_12295,N_11370,N_11755);
or U12296 (N_12296,N_11712,N_11404);
or U12297 (N_12297,N_11938,N_11285);
nand U12298 (N_12298,N_11498,N_11399);
or U12299 (N_12299,N_11925,N_11875);
xnor U12300 (N_12300,N_11447,N_11691);
nand U12301 (N_12301,N_11338,N_11298);
or U12302 (N_12302,N_11993,N_11434);
nand U12303 (N_12303,N_11300,N_11431);
and U12304 (N_12304,N_11488,N_11926);
nor U12305 (N_12305,N_11306,N_11261);
nand U12306 (N_12306,N_11647,N_11642);
xnor U12307 (N_12307,N_11540,N_11858);
or U12308 (N_12308,N_11573,N_11959);
nor U12309 (N_12309,N_11704,N_11877);
and U12310 (N_12310,N_11418,N_11953);
or U12311 (N_12311,N_11776,N_11802);
and U12312 (N_12312,N_11526,N_11809);
or U12313 (N_12313,N_11675,N_11886);
and U12314 (N_12314,N_11972,N_11896);
and U12315 (N_12315,N_11585,N_11446);
xor U12316 (N_12316,N_11334,N_11819);
nor U12317 (N_12317,N_11916,N_11971);
nor U12318 (N_12318,N_11769,N_11662);
xnor U12319 (N_12319,N_11494,N_11797);
nand U12320 (N_12320,N_11364,N_11696);
and U12321 (N_12321,N_11979,N_11906);
or U12322 (N_12322,N_11457,N_11760);
xnor U12323 (N_12323,N_11719,N_11412);
xor U12324 (N_12324,N_11775,N_11934);
nand U12325 (N_12325,N_11263,N_11907);
and U12326 (N_12326,N_11379,N_11336);
and U12327 (N_12327,N_11748,N_11619);
nand U12328 (N_12328,N_11980,N_11394);
nand U12329 (N_12329,N_11859,N_11496);
nor U12330 (N_12330,N_11532,N_11928);
xor U12331 (N_12331,N_11520,N_11882);
nor U12332 (N_12332,N_11918,N_11688);
xor U12333 (N_12333,N_11752,N_11463);
nand U12334 (N_12334,N_11683,N_11740);
nor U12335 (N_12335,N_11357,N_11609);
nor U12336 (N_12336,N_11268,N_11813);
and U12337 (N_12337,N_11558,N_11720);
nor U12338 (N_12338,N_11260,N_11828);
or U12339 (N_12339,N_11672,N_11659);
nand U12340 (N_12340,N_11921,N_11808);
nor U12341 (N_12341,N_11715,N_11321);
or U12342 (N_12342,N_11437,N_11597);
nor U12343 (N_12343,N_11450,N_11873);
and U12344 (N_12344,N_11269,N_11348);
and U12345 (N_12345,N_11542,N_11436);
nor U12346 (N_12346,N_11632,N_11839);
or U12347 (N_12347,N_11749,N_11477);
nor U12348 (N_12348,N_11515,N_11795);
or U12349 (N_12349,N_11771,N_11930);
nor U12350 (N_12350,N_11658,N_11798);
nor U12351 (N_12351,N_11867,N_11854);
nor U12352 (N_12352,N_11492,N_11943);
or U12353 (N_12353,N_11473,N_11931);
or U12354 (N_12354,N_11462,N_11830);
or U12355 (N_12355,N_11460,N_11757);
nor U12356 (N_12356,N_11513,N_11892);
nand U12357 (N_12357,N_11872,N_11635);
nor U12358 (N_12358,N_11753,N_11444);
or U12359 (N_12359,N_11356,N_11483);
nand U12360 (N_12360,N_11891,N_11744);
nor U12361 (N_12361,N_11314,N_11299);
nand U12362 (N_12362,N_11864,N_11405);
xnor U12363 (N_12363,N_11901,N_11648);
or U12364 (N_12364,N_11710,N_11977);
nor U12365 (N_12365,N_11679,N_11579);
and U12366 (N_12366,N_11759,N_11576);
nor U12367 (N_12367,N_11948,N_11708);
and U12368 (N_12368,N_11803,N_11351);
or U12369 (N_12369,N_11335,N_11358);
nor U12370 (N_12370,N_11301,N_11995);
and U12371 (N_12371,N_11315,N_11676);
nand U12372 (N_12372,N_11982,N_11898);
nor U12373 (N_12373,N_11756,N_11747);
nor U12374 (N_12374,N_11359,N_11277);
or U12375 (N_12375,N_11734,N_11755);
or U12376 (N_12376,N_11569,N_11585);
nand U12377 (N_12377,N_11947,N_11985);
or U12378 (N_12378,N_11914,N_11876);
or U12379 (N_12379,N_11283,N_11649);
nor U12380 (N_12380,N_11283,N_11979);
nor U12381 (N_12381,N_11807,N_11866);
or U12382 (N_12382,N_11677,N_11748);
nand U12383 (N_12383,N_11631,N_11984);
nor U12384 (N_12384,N_11826,N_11476);
and U12385 (N_12385,N_11801,N_11453);
and U12386 (N_12386,N_11521,N_11847);
xor U12387 (N_12387,N_11591,N_11793);
and U12388 (N_12388,N_11719,N_11408);
nor U12389 (N_12389,N_11992,N_11263);
and U12390 (N_12390,N_11360,N_11343);
and U12391 (N_12391,N_11995,N_11459);
or U12392 (N_12392,N_11973,N_11798);
or U12393 (N_12393,N_11648,N_11283);
nor U12394 (N_12394,N_11557,N_11293);
and U12395 (N_12395,N_11399,N_11870);
nand U12396 (N_12396,N_11685,N_11585);
nand U12397 (N_12397,N_11769,N_11717);
nand U12398 (N_12398,N_11278,N_11765);
or U12399 (N_12399,N_11654,N_11850);
nor U12400 (N_12400,N_11681,N_11899);
and U12401 (N_12401,N_11681,N_11692);
or U12402 (N_12402,N_11770,N_11570);
and U12403 (N_12403,N_11488,N_11370);
nor U12404 (N_12404,N_11839,N_11790);
nor U12405 (N_12405,N_11928,N_11764);
nand U12406 (N_12406,N_11858,N_11498);
nor U12407 (N_12407,N_11274,N_11347);
nor U12408 (N_12408,N_11725,N_11319);
or U12409 (N_12409,N_11741,N_11292);
nor U12410 (N_12410,N_11817,N_11440);
nand U12411 (N_12411,N_11866,N_11320);
or U12412 (N_12412,N_11719,N_11497);
xor U12413 (N_12413,N_11833,N_11357);
nor U12414 (N_12414,N_11400,N_11758);
nand U12415 (N_12415,N_11694,N_11842);
or U12416 (N_12416,N_11349,N_11660);
nand U12417 (N_12417,N_11302,N_11352);
nand U12418 (N_12418,N_11692,N_11461);
and U12419 (N_12419,N_11976,N_11887);
and U12420 (N_12420,N_11430,N_11534);
and U12421 (N_12421,N_11787,N_11839);
and U12422 (N_12422,N_11546,N_11344);
xnor U12423 (N_12423,N_11703,N_11945);
or U12424 (N_12424,N_11577,N_11466);
or U12425 (N_12425,N_11780,N_11785);
or U12426 (N_12426,N_11525,N_11837);
nand U12427 (N_12427,N_11496,N_11477);
nor U12428 (N_12428,N_11253,N_11929);
or U12429 (N_12429,N_11898,N_11507);
nor U12430 (N_12430,N_11910,N_11569);
nor U12431 (N_12431,N_11838,N_11909);
and U12432 (N_12432,N_11610,N_11620);
nor U12433 (N_12433,N_11969,N_11261);
nor U12434 (N_12434,N_11376,N_11428);
nand U12435 (N_12435,N_11754,N_11915);
and U12436 (N_12436,N_11815,N_11614);
nor U12437 (N_12437,N_11939,N_11254);
or U12438 (N_12438,N_11322,N_11776);
nand U12439 (N_12439,N_11381,N_11409);
and U12440 (N_12440,N_11654,N_11971);
xor U12441 (N_12441,N_11815,N_11905);
or U12442 (N_12442,N_11397,N_11992);
nor U12443 (N_12443,N_11611,N_11933);
nand U12444 (N_12444,N_11678,N_11298);
or U12445 (N_12445,N_11292,N_11318);
xor U12446 (N_12446,N_11902,N_11556);
nand U12447 (N_12447,N_11557,N_11766);
nand U12448 (N_12448,N_11567,N_11950);
or U12449 (N_12449,N_11357,N_11898);
xnor U12450 (N_12450,N_11844,N_11827);
nor U12451 (N_12451,N_11439,N_11713);
nand U12452 (N_12452,N_11739,N_11480);
or U12453 (N_12453,N_11784,N_11769);
and U12454 (N_12454,N_11447,N_11623);
xor U12455 (N_12455,N_11535,N_11543);
nand U12456 (N_12456,N_11807,N_11505);
and U12457 (N_12457,N_11744,N_11558);
or U12458 (N_12458,N_11730,N_11458);
or U12459 (N_12459,N_11261,N_11324);
nor U12460 (N_12460,N_11386,N_11738);
nand U12461 (N_12461,N_11816,N_11713);
or U12462 (N_12462,N_11419,N_11635);
or U12463 (N_12463,N_11672,N_11751);
nand U12464 (N_12464,N_11469,N_11770);
nand U12465 (N_12465,N_11958,N_11734);
nand U12466 (N_12466,N_11744,N_11899);
and U12467 (N_12467,N_11573,N_11917);
nand U12468 (N_12468,N_11559,N_11717);
or U12469 (N_12469,N_11797,N_11969);
nor U12470 (N_12470,N_11257,N_11871);
or U12471 (N_12471,N_11423,N_11843);
nand U12472 (N_12472,N_11329,N_11622);
and U12473 (N_12473,N_11926,N_11652);
nand U12474 (N_12474,N_11455,N_11353);
xor U12475 (N_12475,N_11534,N_11423);
nand U12476 (N_12476,N_11483,N_11833);
or U12477 (N_12477,N_11903,N_11952);
nand U12478 (N_12478,N_11357,N_11691);
nand U12479 (N_12479,N_11799,N_11314);
nand U12480 (N_12480,N_11590,N_11459);
or U12481 (N_12481,N_11689,N_11773);
or U12482 (N_12482,N_11974,N_11639);
nor U12483 (N_12483,N_11829,N_11957);
nor U12484 (N_12484,N_11615,N_11897);
and U12485 (N_12485,N_11523,N_11600);
nor U12486 (N_12486,N_11267,N_11942);
xnor U12487 (N_12487,N_11544,N_11361);
nand U12488 (N_12488,N_11433,N_11545);
and U12489 (N_12489,N_11325,N_11785);
and U12490 (N_12490,N_11706,N_11513);
and U12491 (N_12491,N_11414,N_11796);
nand U12492 (N_12492,N_11486,N_11398);
nand U12493 (N_12493,N_11736,N_11284);
or U12494 (N_12494,N_11676,N_11827);
nor U12495 (N_12495,N_11347,N_11572);
and U12496 (N_12496,N_11964,N_11398);
nand U12497 (N_12497,N_11496,N_11870);
or U12498 (N_12498,N_11728,N_11460);
nor U12499 (N_12499,N_11713,N_11681);
or U12500 (N_12500,N_11750,N_11757);
xor U12501 (N_12501,N_11676,N_11433);
and U12502 (N_12502,N_11991,N_11371);
nand U12503 (N_12503,N_11751,N_11603);
nand U12504 (N_12504,N_11895,N_11470);
xnor U12505 (N_12505,N_11687,N_11597);
and U12506 (N_12506,N_11471,N_11709);
or U12507 (N_12507,N_11561,N_11458);
or U12508 (N_12508,N_11909,N_11343);
nand U12509 (N_12509,N_11286,N_11381);
and U12510 (N_12510,N_11539,N_11809);
and U12511 (N_12511,N_11589,N_11820);
nand U12512 (N_12512,N_11894,N_11701);
or U12513 (N_12513,N_11442,N_11556);
nor U12514 (N_12514,N_11799,N_11273);
and U12515 (N_12515,N_11810,N_11677);
nand U12516 (N_12516,N_11968,N_11410);
xor U12517 (N_12517,N_11584,N_11947);
xnor U12518 (N_12518,N_11717,N_11425);
xor U12519 (N_12519,N_11294,N_11419);
or U12520 (N_12520,N_11939,N_11930);
or U12521 (N_12521,N_11727,N_11255);
and U12522 (N_12522,N_11406,N_11639);
nand U12523 (N_12523,N_11720,N_11578);
nand U12524 (N_12524,N_11954,N_11435);
xor U12525 (N_12525,N_11253,N_11636);
xnor U12526 (N_12526,N_11292,N_11789);
and U12527 (N_12527,N_11560,N_11890);
and U12528 (N_12528,N_11995,N_11445);
and U12529 (N_12529,N_11441,N_11352);
nor U12530 (N_12530,N_11802,N_11418);
nor U12531 (N_12531,N_11555,N_11330);
nand U12532 (N_12532,N_11263,N_11289);
or U12533 (N_12533,N_11273,N_11710);
nor U12534 (N_12534,N_11537,N_11654);
or U12535 (N_12535,N_11598,N_11762);
and U12536 (N_12536,N_11973,N_11983);
or U12537 (N_12537,N_11793,N_11811);
nand U12538 (N_12538,N_11866,N_11361);
nor U12539 (N_12539,N_11266,N_11866);
nand U12540 (N_12540,N_11747,N_11372);
and U12541 (N_12541,N_11801,N_11482);
nor U12542 (N_12542,N_11607,N_11979);
nand U12543 (N_12543,N_11339,N_11809);
and U12544 (N_12544,N_11369,N_11514);
nor U12545 (N_12545,N_11977,N_11299);
or U12546 (N_12546,N_11500,N_11909);
and U12547 (N_12547,N_11518,N_11330);
nor U12548 (N_12548,N_11963,N_11986);
or U12549 (N_12549,N_11764,N_11942);
or U12550 (N_12550,N_11735,N_11287);
nor U12551 (N_12551,N_11734,N_11445);
nor U12552 (N_12552,N_11833,N_11256);
and U12553 (N_12553,N_11469,N_11251);
xnor U12554 (N_12554,N_11345,N_11574);
or U12555 (N_12555,N_11803,N_11812);
nor U12556 (N_12556,N_11331,N_11358);
and U12557 (N_12557,N_11576,N_11946);
and U12558 (N_12558,N_11839,N_11472);
and U12559 (N_12559,N_11315,N_11823);
and U12560 (N_12560,N_11621,N_11607);
nor U12561 (N_12561,N_11843,N_11727);
nand U12562 (N_12562,N_11411,N_11978);
xor U12563 (N_12563,N_11830,N_11684);
and U12564 (N_12564,N_11952,N_11398);
nor U12565 (N_12565,N_11442,N_11725);
and U12566 (N_12566,N_11854,N_11994);
and U12567 (N_12567,N_11830,N_11835);
nand U12568 (N_12568,N_11308,N_11797);
xnor U12569 (N_12569,N_11692,N_11527);
nor U12570 (N_12570,N_11931,N_11318);
xnor U12571 (N_12571,N_11300,N_11524);
xnor U12572 (N_12572,N_11744,N_11726);
and U12573 (N_12573,N_11263,N_11657);
nand U12574 (N_12574,N_11688,N_11521);
xor U12575 (N_12575,N_11408,N_11969);
nor U12576 (N_12576,N_11460,N_11298);
nand U12577 (N_12577,N_11271,N_11749);
nor U12578 (N_12578,N_11997,N_11697);
nor U12579 (N_12579,N_11873,N_11862);
or U12580 (N_12580,N_11459,N_11386);
and U12581 (N_12581,N_11650,N_11639);
nor U12582 (N_12582,N_11424,N_11809);
or U12583 (N_12583,N_11864,N_11472);
nand U12584 (N_12584,N_11768,N_11880);
and U12585 (N_12585,N_11770,N_11881);
and U12586 (N_12586,N_11320,N_11560);
or U12587 (N_12587,N_11409,N_11300);
and U12588 (N_12588,N_11499,N_11290);
and U12589 (N_12589,N_11620,N_11979);
or U12590 (N_12590,N_11537,N_11989);
or U12591 (N_12591,N_11803,N_11915);
or U12592 (N_12592,N_11365,N_11254);
and U12593 (N_12593,N_11413,N_11745);
nor U12594 (N_12594,N_11306,N_11288);
nor U12595 (N_12595,N_11758,N_11409);
nor U12596 (N_12596,N_11368,N_11736);
or U12597 (N_12597,N_11769,N_11478);
xnor U12598 (N_12598,N_11943,N_11946);
or U12599 (N_12599,N_11306,N_11683);
nand U12600 (N_12600,N_11370,N_11522);
xnor U12601 (N_12601,N_11453,N_11439);
nor U12602 (N_12602,N_11379,N_11581);
nand U12603 (N_12603,N_11698,N_11902);
nand U12604 (N_12604,N_11996,N_11439);
nand U12605 (N_12605,N_11849,N_11591);
or U12606 (N_12606,N_11801,N_11371);
nand U12607 (N_12607,N_11550,N_11903);
and U12608 (N_12608,N_11400,N_11272);
nor U12609 (N_12609,N_11791,N_11782);
nand U12610 (N_12610,N_11790,N_11332);
or U12611 (N_12611,N_11794,N_11786);
and U12612 (N_12612,N_11811,N_11364);
and U12613 (N_12613,N_11735,N_11847);
or U12614 (N_12614,N_11536,N_11298);
or U12615 (N_12615,N_11490,N_11745);
nand U12616 (N_12616,N_11575,N_11267);
and U12617 (N_12617,N_11445,N_11806);
nor U12618 (N_12618,N_11287,N_11879);
xor U12619 (N_12619,N_11441,N_11522);
nand U12620 (N_12620,N_11313,N_11539);
xnor U12621 (N_12621,N_11280,N_11583);
nor U12622 (N_12622,N_11425,N_11440);
and U12623 (N_12623,N_11270,N_11864);
or U12624 (N_12624,N_11300,N_11908);
and U12625 (N_12625,N_11722,N_11624);
xnor U12626 (N_12626,N_11265,N_11353);
or U12627 (N_12627,N_11689,N_11377);
and U12628 (N_12628,N_11887,N_11589);
nand U12629 (N_12629,N_11898,N_11524);
and U12630 (N_12630,N_11473,N_11541);
nor U12631 (N_12631,N_11730,N_11980);
or U12632 (N_12632,N_11476,N_11927);
nor U12633 (N_12633,N_11549,N_11699);
and U12634 (N_12634,N_11518,N_11836);
and U12635 (N_12635,N_11776,N_11386);
or U12636 (N_12636,N_11493,N_11297);
nor U12637 (N_12637,N_11926,N_11532);
xor U12638 (N_12638,N_11293,N_11752);
nand U12639 (N_12639,N_11945,N_11590);
nand U12640 (N_12640,N_11735,N_11683);
nor U12641 (N_12641,N_11523,N_11763);
nand U12642 (N_12642,N_11371,N_11255);
or U12643 (N_12643,N_11636,N_11713);
and U12644 (N_12644,N_11912,N_11288);
nor U12645 (N_12645,N_11365,N_11653);
and U12646 (N_12646,N_11561,N_11610);
or U12647 (N_12647,N_11272,N_11462);
and U12648 (N_12648,N_11996,N_11826);
nand U12649 (N_12649,N_11382,N_11778);
nor U12650 (N_12650,N_11422,N_11739);
xnor U12651 (N_12651,N_11285,N_11772);
and U12652 (N_12652,N_11740,N_11986);
nand U12653 (N_12653,N_11632,N_11920);
and U12654 (N_12654,N_11949,N_11409);
or U12655 (N_12655,N_11982,N_11688);
nand U12656 (N_12656,N_11426,N_11877);
and U12657 (N_12657,N_11638,N_11463);
nor U12658 (N_12658,N_11367,N_11924);
nor U12659 (N_12659,N_11319,N_11752);
nand U12660 (N_12660,N_11853,N_11928);
nor U12661 (N_12661,N_11375,N_11733);
xor U12662 (N_12662,N_11676,N_11614);
or U12663 (N_12663,N_11866,N_11971);
nand U12664 (N_12664,N_11398,N_11854);
and U12665 (N_12665,N_11424,N_11286);
xor U12666 (N_12666,N_11640,N_11303);
xor U12667 (N_12667,N_11267,N_11635);
nor U12668 (N_12668,N_11926,N_11555);
nand U12669 (N_12669,N_11926,N_11628);
and U12670 (N_12670,N_11741,N_11369);
and U12671 (N_12671,N_11332,N_11955);
xnor U12672 (N_12672,N_11634,N_11791);
xnor U12673 (N_12673,N_11360,N_11427);
nor U12674 (N_12674,N_11400,N_11569);
and U12675 (N_12675,N_11657,N_11642);
and U12676 (N_12676,N_11324,N_11714);
nand U12677 (N_12677,N_11447,N_11591);
nand U12678 (N_12678,N_11479,N_11385);
or U12679 (N_12679,N_11465,N_11267);
nor U12680 (N_12680,N_11750,N_11654);
xnor U12681 (N_12681,N_11365,N_11550);
nor U12682 (N_12682,N_11695,N_11495);
and U12683 (N_12683,N_11943,N_11253);
nand U12684 (N_12684,N_11636,N_11945);
or U12685 (N_12685,N_11945,N_11685);
nand U12686 (N_12686,N_11603,N_11987);
or U12687 (N_12687,N_11616,N_11524);
nor U12688 (N_12688,N_11315,N_11722);
nand U12689 (N_12689,N_11306,N_11480);
and U12690 (N_12690,N_11548,N_11918);
nand U12691 (N_12691,N_11947,N_11490);
and U12692 (N_12692,N_11818,N_11797);
nor U12693 (N_12693,N_11504,N_11757);
and U12694 (N_12694,N_11856,N_11667);
nand U12695 (N_12695,N_11685,N_11451);
and U12696 (N_12696,N_11403,N_11303);
nor U12697 (N_12697,N_11606,N_11426);
nor U12698 (N_12698,N_11443,N_11754);
nor U12699 (N_12699,N_11496,N_11250);
nand U12700 (N_12700,N_11595,N_11990);
and U12701 (N_12701,N_11517,N_11777);
nand U12702 (N_12702,N_11411,N_11523);
or U12703 (N_12703,N_11589,N_11679);
nor U12704 (N_12704,N_11311,N_11842);
and U12705 (N_12705,N_11651,N_11715);
nand U12706 (N_12706,N_11699,N_11795);
nor U12707 (N_12707,N_11415,N_11527);
nor U12708 (N_12708,N_11385,N_11426);
or U12709 (N_12709,N_11931,N_11587);
or U12710 (N_12710,N_11611,N_11968);
or U12711 (N_12711,N_11678,N_11290);
nand U12712 (N_12712,N_11996,N_11814);
or U12713 (N_12713,N_11886,N_11521);
and U12714 (N_12714,N_11394,N_11890);
xnor U12715 (N_12715,N_11300,N_11913);
or U12716 (N_12716,N_11995,N_11560);
and U12717 (N_12717,N_11900,N_11256);
and U12718 (N_12718,N_11863,N_11613);
nor U12719 (N_12719,N_11496,N_11610);
nand U12720 (N_12720,N_11579,N_11362);
xor U12721 (N_12721,N_11501,N_11332);
nor U12722 (N_12722,N_11887,N_11531);
and U12723 (N_12723,N_11359,N_11950);
nand U12724 (N_12724,N_11599,N_11422);
nand U12725 (N_12725,N_11840,N_11460);
nor U12726 (N_12726,N_11887,N_11628);
or U12727 (N_12727,N_11670,N_11309);
nor U12728 (N_12728,N_11591,N_11572);
nor U12729 (N_12729,N_11976,N_11305);
or U12730 (N_12730,N_11447,N_11924);
or U12731 (N_12731,N_11289,N_11697);
xnor U12732 (N_12732,N_11547,N_11410);
nand U12733 (N_12733,N_11492,N_11979);
nor U12734 (N_12734,N_11994,N_11263);
and U12735 (N_12735,N_11747,N_11928);
nor U12736 (N_12736,N_11367,N_11587);
nand U12737 (N_12737,N_11641,N_11620);
and U12738 (N_12738,N_11909,N_11868);
nor U12739 (N_12739,N_11598,N_11307);
or U12740 (N_12740,N_11676,N_11830);
or U12741 (N_12741,N_11426,N_11273);
nand U12742 (N_12742,N_11382,N_11302);
and U12743 (N_12743,N_11944,N_11637);
nand U12744 (N_12744,N_11838,N_11491);
or U12745 (N_12745,N_11956,N_11433);
nand U12746 (N_12746,N_11830,N_11651);
nor U12747 (N_12747,N_11477,N_11259);
and U12748 (N_12748,N_11328,N_11644);
xor U12749 (N_12749,N_11403,N_11682);
nand U12750 (N_12750,N_12604,N_12135);
and U12751 (N_12751,N_12409,N_12746);
or U12752 (N_12752,N_12251,N_12425);
or U12753 (N_12753,N_12556,N_12276);
nand U12754 (N_12754,N_12643,N_12025);
xor U12755 (N_12755,N_12460,N_12228);
nor U12756 (N_12756,N_12513,N_12118);
or U12757 (N_12757,N_12637,N_12654);
nand U12758 (N_12758,N_12588,N_12323);
and U12759 (N_12759,N_12043,N_12255);
nand U12760 (N_12760,N_12400,N_12231);
and U12761 (N_12761,N_12545,N_12666);
or U12762 (N_12762,N_12241,N_12442);
and U12763 (N_12763,N_12064,N_12395);
nor U12764 (N_12764,N_12273,N_12258);
nor U12765 (N_12765,N_12107,N_12480);
nand U12766 (N_12766,N_12670,N_12188);
nand U12767 (N_12767,N_12608,N_12354);
or U12768 (N_12768,N_12248,N_12557);
nand U12769 (N_12769,N_12221,N_12490);
or U12770 (N_12770,N_12578,N_12410);
nand U12771 (N_12771,N_12671,N_12407);
nand U12772 (N_12772,N_12408,N_12735);
nand U12773 (N_12773,N_12325,N_12472);
and U12774 (N_12774,N_12558,N_12309);
xnor U12775 (N_12775,N_12317,N_12101);
nand U12776 (N_12776,N_12374,N_12146);
nand U12777 (N_12777,N_12688,N_12530);
nor U12778 (N_12778,N_12290,N_12669);
xor U12779 (N_12779,N_12635,N_12569);
or U12780 (N_12780,N_12217,N_12040);
nor U12781 (N_12781,N_12443,N_12381);
nand U12782 (N_12782,N_12646,N_12121);
nand U12783 (N_12783,N_12029,N_12428);
or U12784 (N_12784,N_12544,N_12535);
xnor U12785 (N_12785,N_12445,N_12162);
and U12786 (N_12786,N_12726,N_12696);
and U12787 (N_12787,N_12300,N_12731);
nand U12788 (N_12788,N_12389,N_12277);
nor U12789 (N_12789,N_12385,N_12229);
nor U12790 (N_12790,N_12437,N_12620);
nand U12791 (N_12791,N_12542,N_12463);
nand U12792 (N_12792,N_12739,N_12705);
nand U12793 (N_12793,N_12244,N_12414);
and U12794 (N_12794,N_12479,N_12159);
and U12795 (N_12795,N_12194,N_12432);
nor U12796 (N_12796,N_12134,N_12176);
or U12797 (N_12797,N_12648,N_12239);
and U12798 (N_12798,N_12115,N_12464);
or U12799 (N_12799,N_12091,N_12185);
nand U12800 (N_12800,N_12059,N_12177);
nor U12801 (N_12801,N_12362,N_12289);
nand U12802 (N_12802,N_12291,N_12268);
nor U12803 (N_12803,N_12304,N_12266);
nor U12804 (N_12804,N_12543,N_12413);
or U12805 (N_12805,N_12677,N_12538);
nor U12806 (N_12806,N_12456,N_12070);
xnor U12807 (N_12807,N_12022,N_12250);
and U12808 (N_12808,N_12449,N_12576);
xnor U12809 (N_12809,N_12392,N_12675);
or U12810 (N_12810,N_12508,N_12020);
nand U12811 (N_12811,N_12729,N_12347);
or U12812 (N_12812,N_12516,N_12404);
and U12813 (N_12813,N_12361,N_12327);
and U12814 (N_12814,N_12458,N_12190);
nor U12815 (N_12815,N_12468,N_12682);
nand U12816 (N_12816,N_12519,N_12205);
and U12817 (N_12817,N_12088,N_12384);
and U12818 (N_12818,N_12685,N_12000);
and U12819 (N_12819,N_12707,N_12138);
nand U12820 (N_12820,N_12218,N_12322);
nor U12821 (N_12821,N_12537,N_12223);
or U12822 (N_12822,N_12096,N_12174);
nor U12823 (N_12823,N_12728,N_12242);
and U12824 (N_12824,N_12485,N_12524);
nor U12825 (N_12825,N_12306,N_12623);
nand U12826 (N_12826,N_12377,N_12252);
nor U12827 (N_12827,N_12582,N_12405);
nor U12828 (N_12828,N_12318,N_12717);
nand U12829 (N_12829,N_12099,N_12553);
nand U12830 (N_12830,N_12532,N_12390);
nand U12831 (N_12831,N_12411,N_12073);
nand U12832 (N_12832,N_12703,N_12527);
and U12833 (N_12833,N_12140,N_12195);
nand U12834 (N_12834,N_12048,N_12035);
and U12835 (N_12835,N_12511,N_12111);
and U12836 (N_12836,N_12216,N_12610);
nor U12837 (N_12837,N_12055,N_12619);
or U12838 (N_12838,N_12355,N_12271);
or U12839 (N_12839,N_12313,N_12534);
xor U12840 (N_12840,N_12503,N_12539);
xnor U12841 (N_12841,N_12267,N_12698);
nand U12842 (N_12842,N_12226,N_12279);
nand U12843 (N_12843,N_12398,N_12473);
or U12844 (N_12844,N_12531,N_12403);
xnor U12845 (N_12845,N_12214,N_12533);
nor U12846 (N_12846,N_12621,N_12585);
or U12847 (N_12847,N_12475,N_12122);
or U12848 (N_12848,N_12567,N_12393);
or U12849 (N_12849,N_12056,N_12343);
and U12850 (N_12850,N_12075,N_12492);
xor U12851 (N_12851,N_12329,N_12357);
nor U12852 (N_12852,N_12315,N_12388);
or U12853 (N_12853,N_12664,N_12548);
or U12854 (N_12854,N_12636,N_12676);
nand U12855 (N_12855,N_12068,N_12733);
or U12856 (N_12856,N_12320,N_12067);
nor U12857 (N_12857,N_12094,N_12353);
nor U12858 (N_12858,N_12642,N_12147);
or U12859 (N_12859,N_12287,N_12038);
nor U12860 (N_12860,N_12562,N_12382);
and U12861 (N_12861,N_12657,N_12074);
and U12862 (N_12862,N_12718,N_12697);
or U12863 (N_12863,N_12573,N_12219);
xor U12864 (N_12864,N_12150,N_12541);
nor U12865 (N_12865,N_12120,N_12574);
nor U12866 (N_12866,N_12615,N_12589);
or U12867 (N_12867,N_12256,N_12299);
or U12868 (N_12868,N_12607,N_12701);
nor U12869 (N_12869,N_12128,N_12166);
nand U12870 (N_12870,N_12416,N_12372);
nand U12871 (N_12871,N_12206,N_12584);
nor U12872 (N_12872,N_12618,N_12529);
and U12873 (N_12873,N_12233,N_12278);
and U12874 (N_12874,N_12023,N_12652);
xnor U12875 (N_12875,N_12011,N_12744);
nor U12876 (N_12876,N_12611,N_12502);
nor U12877 (N_12877,N_12518,N_12647);
or U12878 (N_12878,N_12366,N_12339);
xor U12879 (N_12879,N_12375,N_12336);
nand U12880 (N_12880,N_12429,N_12561);
nand U12881 (N_12881,N_12509,N_12139);
nor U12882 (N_12882,N_12046,N_12624);
or U12883 (N_12883,N_12178,N_12465);
xor U12884 (N_12884,N_12097,N_12655);
nor U12885 (N_12885,N_12148,N_12560);
and U12886 (N_12886,N_12047,N_12184);
nand U12887 (N_12887,N_12512,N_12462);
and U12888 (N_12888,N_12286,N_12272);
and U12889 (N_12889,N_12625,N_12100);
or U12890 (N_12890,N_12477,N_12732);
or U12891 (N_12891,N_12630,N_12716);
nor U12892 (N_12892,N_12015,N_12487);
or U12893 (N_12893,N_12238,N_12667);
xnor U12894 (N_12894,N_12161,N_12709);
nand U12895 (N_12895,N_12722,N_12734);
xnor U12896 (N_12896,N_12743,N_12123);
nand U12897 (N_12897,N_12145,N_12110);
or U12898 (N_12898,N_12672,N_12605);
or U12899 (N_12899,N_12358,N_12215);
nor U12900 (N_12900,N_12725,N_12466);
or U12901 (N_12901,N_12319,N_12476);
or U12902 (N_12902,N_12263,N_12684);
nand U12903 (N_12903,N_12702,N_12665);
or U12904 (N_12904,N_12474,N_12027);
and U12905 (N_12905,N_12564,N_12126);
nor U12906 (N_12906,N_12024,N_12658);
nand U12907 (N_12907,N_12417,N_12640);
or U12908 (N_12908,N_12663,N_12418);
or U12909 (N_12909,N_12203,N_12631);
and U12910 (N_12910,N_12246,N_12007);
nand U12911 (N_12911,N_12507,N_12438);
xor U12912 (N_12912,N_12453,N_12639);
nand U12913 (N_12913,N_12295,N_12280);
or U12914 (N_12914,N_12481,N_12435);
xnor U12915 (N_12915,N_12748,N_12613);
nand U12916 (N_12916,N_12211,N_12719);
or U12917 (N_12917,N_12371,N_12434);
or U12918 (N_12918,N_12152,N_12133);
nor U12919 (N_12919,N_12105,N_12365);
xnor U12920 (N_12920,N_12687,N_12247);
nor U12921 (N_12921,N_12198,N_12552);
nor U12922 (N_12922,N_12269,N_12540);
and U12923 (N_12923,N_12708,N_12264);
or U12924 (N_12924,N_12370,N_12634);
or U12925 (N_12925,N_12491,N_12420);
nand U12926 (N_12926,N_12285,N_12451);
nor U12927 (N_12927,N_12494,N_12575);
nand U12928 (N_12928,N_12419,N_12222);
nor U12929 (N_12929,N_12614,N_12501);
xnor U12930 (N_12930,N_12600,N_12436);
nand U12931 (N_12931,N_12338,N_12316);
and U12932 (N_12932,N_12302,N_12092);
nor U12933 (N_12933,N_12124,N_12712);
and U12934 (N_12934,N_12627,N_12660);
or U12935 (N_12935,N_12335,N_12207);
xor U12936 (N_12936,N_12373,N_12282);
nor U12937 (N_12937,N_12072,N_12587);
nor U12938 (N_12938,N_12412,N_12401);
and U12939 (N_12939,N_12051,N_12571);
nor U12940 (N_12940,N_12192,N_12061);
and U12941 (N_12941,N_12704,N_12397);
or U12942 (N_12942,N_12431,N_12379);
xor U12943 (N_12943,N_12077,N_12060);
nand U12944 (N_12944,N_12156,N_12334);
or U12945 (N_12945,N_12692,N_12199);
and U12946 (N_12946,N_12577,N_12583);
nand U12947 (N_12947,N_12202,N_12563);
and U12948 (N_12948,N_12549,N_12141);
xnor U12949 (N_12949,N_12522,N_12484);
nand U12950 (N_12950,N_12617,N_12193);
or U12951 (N_12951,N_12151,N_12298);
nand U12952 (N_12952,N_12525,N_12208);
nor U12953 (N_12953,N_12008,N_12296);
nor U12954 (N_12954,N_12209,N_12052);
nor U12955 (N_12955,N_12262,N_12283);
nand U12956 (N_12956,N_12363,N_12082);
nor U12957 (N_12957,N_12710,N_12127);
or U12958 (N_12958,N_12547,N_12235);
or U12959 (N_12959,N_12153,N_12259);
nand U12960 (N_12960,N_12210,N_12265);
or U12961 (N_12961,N_12175,N_12659);
nor U12962 (N_12962,N_12028,N_12130);
or U12963 (N_12963,N_12181,N_12695);
nand U12964 (N_12964,N_12715,N_12517);
nand U12965 (N_12965,N_12570,N_12469);
nor U12966 (N_12966,N_12565,N_12143);
nand U12967 (N_12967,N_12590,N_12650);
nand U12968 (N_12968,N_12036,N_12167);
xor U12969 (N_12969,N_12281,N_12505);
or U12970 (N_12970,N_12426,N_12312);
xor U12971 (N_12971,N_12224,N_12523);
or U12972 (N_12972,N_12144,N_12488);
and U12973 (N_12973,N_12087,N_12160);
and U12974 (N_12974,N_12661,N_12131);
and U12975 (N_12975,N_12689,N_12714);
nor U12976 (N_12976,N_12220,N_12737);
and U12977 (N_12977,N_12236,N_12173);
nor U12978 (N_12978,N_12076,N_12187);
xnor U12979 (N_12979,N_12616,N_12580);
nor U12980 (N_12980,N_12459,N_12747);
and U12981 (N_12981,N_12378,N_12498);
xnor U12982 (N_12982,N_12528,N_12171);
nor U12983 (N_12983,N_12430,N_12200);
nand U12984 (N_12984,N_12653,N_12245);
or U12985 (N_12985,N_12572,N_12034);
nand U12986 (N_12986,N_12489,N_12042);
or U12987 (N_12987,N_12172,N_12033);
nor U12988 (N_12988,N_12369,N_12341);
or U12989 (N_12989,N_12163,N_12196);
and U12990 (N_12990,N_12427,N_12448);
nand U12991 (N_12991,N_12439,N_12555);
xor U12992 (N_12992,N_12514,N_12031);
or U12993 (N_12993,N_12063,N_12597);
and U12994 (N_12994,N_12396,N_12201);
nand U12995 (N_12995,N_12711,N_12730);
nand U12996 (N_12996,N_12227,N_12510);
and U12997 (N_12997,N_12260,N_12310);
nand U12998 (N_12998,N_12331,N_12461);
nand U12999 (N_12999,N_12506,N_12603);
nand U13000 (N_13000,N_12204,N_12457);
nor U13001 (N_13001,N_12742,N_12149);
xnor U13002 (N_13002,N_12213,N_12332);
nor U13003 (N_13003,N_12307,N_12723);
or U13004 (N_13004,N_12612,N_12275);
nand U13005 (N_13005,N_12536,N_12521);
and U13006 (N_13006,N_12109,N_12380);
nor U13007 (N_13007,N_12526,N_12333);
nor U13008 (N_13008,N_12595,N_12674);
nor U13009 (N_13009,N_12550,N_12132);
nor U13010 (N_13010,N_12013,N_12649);
nor U13011 (N_13011,N_12119,N_12016);
nand U13012 (N_13012,N_12592,N_12157);
nor U13013 (N_13013,N_12344,N_12387);
nand U13014 (N_13014,N_12293,N_12467);
and U13015 (N_13015,N_12691,N_12738);
or U13016 (N_13016,N_12680,N_12057);
and U13017 (N_13017,N_12720,N_12500);
or U13018 (N_13018,N_12423,N_12212);
or U13019 (N_13019,N_12065,N_12638);
and U13020 (N_13020,N_12721,N_12305);
and U13021 (N_13021,N_12005,N_12651);
and U13022 (N_13022,N_12086,N_12261);
or U13023 (N_13023,N_12274,N_12125);
and U13024 (N_13024,N_12089,N_12058);
nand U13025 (N_13025,N_12154,N_12078);
nand U13026 (N_13026,N_12050,N_12232);
or U13027 (N_13027,N_12546,N_12191);
and U13028 (N_13028,N_12376,N_12006);
nand U13029 (N_13029,N_12444,N_12559);
xor U13030 (N_13030,N_12257,N_12054);
nand U13031 (N_13031,N_12049,N_12568);
and U13032 (N_13032,N_12402,N_12586);
nand U13033 (N_13033,N_12003,N_12359);
nand U13034 (N_13034,N_12520,N_12230);
nand U13035 (N_13035,N_12447,N_12345);
and U13036 (N_13036,N_12679,N_12069);
nand U13037 (N_13037,N_12504,N_12446);
nand U13038 (N_13038,N_12424,N_12019);
nand U13039 (N_13039,N_12083,N_12308);
nand U13040 (N_13040,N_12085,N_12495);
and U13041 (N_13041,N_12693,N_12662);
and U13042 (N_13042,N_12399,N_12137);
nand U13043 (N_13043,N_12002,N_12240);
nor U13044 (N_13044,N_12012,N_12724);
nor U13045 (N_13045,N_12324,N_12292);
nor U13046 (N_13046,N_12041,N_12001);
and U13047 (N_13047,N_12179,N_12515);
and U13048 (N_13048,N_12367,N_12297);
nor U13049 (N_13049,N_12116,N_12706);
or U13050 (N_13050,N_12673,N_12017);
nor U13051 (N_13051,N_12032,N_12591);
nand U13052 (N_13052,N_12346,N_12071);
nand U13053 (N_13053,N_12727,N_12197);
and U13054 (N_13054,N_12155,N_12062);
nor U13055 (N_13055,N_12243,N_12189);
and U13056 (N_13056,N_12303,N_12164);
nand U13057 (N_13057,N_12694,N_12601);
nand U13058 (N_13058,N_12606,N_12326);
nand U13059 (N_13059,N_12237,N_12018);
xor U13060 (N_13060,N_12579,N_12225);
or U13061 (N_13061,N_12004,N_12348);
nor U13062 (N_13062,N_12566,N_12644);
xor U13063 (N_13063,N_12483,N_12352);
nor U13064 (N_13064,N_12337,N_12478);
nor U13065 (N_13065,N_12632,N_12471);
nand U13066 (N_13066,N_12386,N_12112);
and U13067 (N_13067,N_12749,N_12598);
or U13068 (N_13068,N_12169,N_12093);
nand U13069 (N_13069,N_12328,N_12182);
nand U13070 (N_13070,N_12081,N_12368);
or U13071 (N_13071,N_12454,N_12356);
xor U13072 (N_13072,N_12641,N_12394);
and U13073 (N_13073,N_12079,N_12186);
nand U13074 (N_13074,N_12683,N_12106);
or U13075 (N_13075,N_12080,N_12441);
nor U13076 (N_13076,N_12009,N_12349);
nand U13077 (N_13077,N_12180,N_12014);
nand U13078 (N_13078,N_12098,N_12165);
nor U13079 (N_13079,N_12740,N_12690);
or U13080 (N_13080,N_12581,N_12628);
or U13081 (N_13081,N_12433,N_12095);
or U13082 (N_13082,N_12037,N_12351);
nand U13083 (N_13083,N_12391,N_12383);
or U13084 (N_13084,N_12629,N_12551);
nor U13085 (N_13085,N_12270,N_12168);
or U13086 (N_13086,N_12415,N_12450);
and U13087 (N_13087,N_12626,N_12599);
or U13088 (N_13088,N_12114,N_12045);
and U13089 (N_13089,N_12084,N_12103);
xnor U13090 (N_13090,N_12364,N_12311);
and U13091 (N_13091,N_12129,N_12596);
and U13092 (N_13092,N_12496,N_12645);
and U13093 (N_13093,N_12554,N_12736);
nor U13094 (N_13094,N_12142,N_12330);
or U13095 (N_13095,N_12158,N_12314);
xor U13096 (N_13096,N_12622,N_12609);
or U13097 (N_13097,N_12321,N_12486);
and U13098 (N_13098,N_12350,N_12288);
nor U13099 (N_13099,N_12421,N_12108);
and U13100 (N_13100,N_12010,N_12633);
and U13101 (N_13101,N_12342,N_12493);
nor U13102 (N_13102,N_12499,N_12497);
or U13103 (N_13103,N_12594,N_12681);
or U13104 (N_13104,N_12340,N_12090);
nor U13105 (N_13105,N_12452,N_12470);
nand U13106 (N_13106,N_12170,N_12284);
nor U13107 (N_13107,N_12482,N_12249);
xnor U13108 (N_13108,N_12253,N_12066);
and U13109 (N_13109,N_12668,N_12254);
nor U13110 (N_13110,N_12602,N_12301);
or U13111 (N_13111,N_12741,N_12656);
and U13112 (N_13112,N_12440,N_12360);
or U13113 (N_13113,N_12678,N_12713);
nand U13114 (N_13114,N_12117,N_12593);
nand U13115 (N_13115,N_12183,N_12021);
and U13116 (N_13116,N_12026,N_12102);
and U13117 (N_13117,N_12406,N_12422);
and U13118 (N_13118,N_12136,N_12455);
or U13119 (N_13119,N_12113,N_12039);
and U13120 (N_13120,N_12699,N_12745);
nand U13121 (N_13121,N_12030,N_12104);
or U13122 (N_13122,N_12700,N_12294);
and U13123 (N_13123,N_12234,N_12686);
or U13124 (N_13124,N_12044,N_12053);
xnor U13125 (N_13125,N_12190,N_12621);
nor U13126 (N_13126,N_12256,N_12245);
and U13127 (N_13127,N_12001,N_12163);
nor U13128 (N_13128,N_12311,N_12368);
nand U13129 (N_13129,N_12239,N_12555);
nand U13130 (N_13130,N_12478,N_12450);
and U13131 (N_13131,N_12717,N_12293);
and U13132 (N_13132,N_12333,N_12068);
nor U13133 (N_13133,N_12505,N_12640);
nor U13134 (N_13134,N_12020,N_12441);
nand U13135 (N_13135,N_12369,N_12311);
nor U13136 (N_13136,N_12383,N_12623);
xnor U13137 (N_13137,N_12043,N_12292);
nand U13138 (N_13138,N_12140,N_12244);
nor U13139 (N_13139,N_12557,N_12711);
or U13140 (N_13140,N_12123,N_12713);
or U13141 (N_13141,N_12280,N_12670);
nor U13142 (N_13142,N_12592,N_12250);
or U13143 (N_13143,N_12343,N_12002);
or U13144 (N_13144,N_12557,N_12738);
xnor U13145 (N_13145,N_12110,N_12358);
and U13146 (N_13146,N_12562,N_12551);
or U13147 (N_13147,N_12251,N_12467);
nand U13148 (N_13148,N_12693,N_12626);
xor U13149 (N_13149,N_12037,N_12365);
nor U13150 (N_13150,N_12602,N_12157);
nor U13151 (N_13151,N_12499,N_12355);
xnor U13152 (N_13152,N_12005,N_12368);
or U13153 (N_13153,N_12032,N_12494);
and U13154 (N_13154,N_12062,N_12088);
nor U13155 (N_13155,N_12191,N_12229);
or U13156 (N_13156,N_12181,N_12060);
or U13157 (N_13157,N_12268,N_12616);
nor U13158 (N_13158,N_12385,N_12460);
or U13159 (N_13159,N_12153,N_12636);
nand U13160 (N_13160,N_12213,N_12600);
nor U13161 (N_13161,N_12279,N_12557);
and U13162 (N_13162,N_12746,N_12538);
nand U13163 (N_13163,N_12429,N_12558);
and U13164 (N_13164,N_12564,N_12662);
nor U13165 (N_13165,N_12366,N_12030);
nor U13166 (N_13166,N_12268,N_12610);
or U13167 (N_13167,N_12635,N_12038);
nand U13168 (N_13168,N_12072,N_12169);
nor U13169 (N_13169,N_12480,N_12168);
and U13170 (N_13170,N_12342,N_12083);
xnor U13171 (N_13171,N_12479,N_12084);
nand U13172 (N_13172,N_12147,N_12649);
nor U13173 (N_13173,N_12296,N_12132);
nand U13174 (N_13174,N_12555,N_12342);
and U13175 (N_13175,N_12563,N_12272);
or U13176 (N_13176,N_12109,N_12034);
nor U13177 (N_13177,N_12665,N_12390);
nand U13178 (N_13178,N_12327,N_12557);
and U13179 (N_13179,N_12618,N_12307);
nor U13180 (N_13180,N_12697,N_12549);
nand U13181 (N_13181,N_12511,N_12525);
or U13182 (N_13182,N_12236,N_12744);
nor U13183 (N_13183,N_12104,N_12203);
nand U13184 (N_13184,N_12037,N_12086);
nor U13185 (N_13185,N_12115,N_12117);
or U13186 (N_13186,N_12189,N_12364);
or U13187 (N_13187,N_12157,N_12428);
xor U13188 (N_13188,N_12455,N_12076);
nor U13189 (N_13189,N_12470,N_12641);
nand U13190 (N_13190,N_12469,N_12490);
nand U13191 (N_13191,N_12238,N_12220);
nand U13192 (N_13192,N_12075,N_12126);
nor U13193 (N_13193,N_12477,N_12508);
and U13194 (N_13194,N_12679,N_12473);
and U13195 (N_13195,N_12162,N_12086);
or U13196 (N_13196,N_12176,N_12473);
nor U13197 (N_13197,N_12220,N_12316);
nor U13198 (N_13198,N_12098,N_12305);
nand U13199 (N_13199,N_12258,N_12479);
or U13200 (N_13200,N_12660,N_12568);
and U13201 (N_13201,N_12632,N_12583);
xor U13202 (N_13202,N_12105,N_12329);
nor U13203 (N_13203,N_12599,N_12596);
nor U13204 (N_13204,N_12459,N_12049);
nand U13205 (N_13205,N_12080,N_12165);
nor U13206 (N_13206,N_12119,N_12113);
nand U13207 (N_13207,N_12613,N_12203);
nand U13208 (N_13208,N_12171,N_12296);
and U13209 (N_13209,N_12019,N_12038);
nor U13210 (N_13210,N_12216,N_12692);
nor U13211 (N_13211,N_12121,N_12141);
nor U13212 (N_13212,N_12526,N_12031);
nand U13213 (N_13213,N_12086,N_12329);
or U13214 (N_13214,N_12356,N_12596);
xor U13215 (N_13215,N_12041,N_12525);
and U13216 (N_13216,N_12007,N_12632);
and U13217 (N_13217,N_12074,N_12559);
or U13218 (N_13218,N_12615,N_12704);
or U13219 (N_13219,N_12291,N_12701);
and U13220 (N_13220,N_12098,N_12423);
and U13221 (N_13221,N_12718,N_12059);
nand U13222 (N_13222,N_12093,N_12678);
and U13223 (N_13223,N_12410,N_12507);
and U13224 (N_13224,N_12656,N_12329);
and U13225 (N_13225,N_12385,N_12006);
or U13226 (N_13226,N_12178,N_12417);
nor U13227 (N_13227,N_12415,N_12545);
nand U13228 (N_13228,N_12051,N_12142);
nand U13229 (N_13229,N_12500,N_12323);
and U13230 (N_13230,N_12047,N_12707);
and U13231 (N_13231,N_12185,N_12194);
xnor U13232 (N_13232,N_12128,N_12676);
or U13233 (N_13233,N_12084,N_12418);
or U13234 (N_13234,N_12658,N_12442);
nand U13235 (N_13235,N_12576,N_12191);
or U13236 (N_13236,N_12745,N_12015);
or U13237 (N_13237,N_12068,N_12136);
or U13238 (N_13238,N_12273,N_12330);
nand U13239 (N_13239,N_12350,N_12411);
and U13240 (N_13240,N_12657,N_12216);
nor U13241 (N_13241,N_12654,N_12055);
nand U13242 (N_13242,N_12661,N_12432);
xor U13243 (N_13243,N_12258,N_12412);
nand U13244 (N_13244,N_12260,N_12133);
or U13245 (N_13245,N_12296,N_12142);
and U13246 (N_13246,N_12127,N_12040);
nand U13247 (N_13247,N_12214,N_12651);
nand U13248 (N_13248,N_12706,N_12578);
nor U13249 (N_13249,N_12081,N_12393);
or U13250 (N_13250,N_12126,N_12203);
nand U13251 (N_13251,N_12433,N_12435);
and U13252 (N_13252,N_12291,N_12290);
nor U13253 (N_13253,N_12355,N_12001);
nand U13254 (N_13254,N_12730,N_12082);
xnor U13255 (N_13255,N_12301,N_12327);
nor U13256 (N_13256,N_12590,N_12235);
nand U13257 (N_13257,N_12347,N_12416);
nor U13258 (N_13258,N_12167,N_12713);
or U13259 (N_13259,N_12102,N_12403);
nor U13260 (N_13260,N_12119,N_12243);
nand U13261 (N_13261,N_12371,N_12678);
and U13262 (N_13262,N_12482,N_12550);
and U13263 (N_13263,N_12289,N_12315);
nand U13264 (N_13264,N_12494,N_12022);
and U13265 (N_13265,N_12256,N_12698);
xor U13266 (N_13266,N_12647,N_12039);
and U13267 (N_13267,N_12211,N_12012);
or U13268 (N_13268,N_12111,N_12544);
or U13269 (N_13269,N_12474,N_12129);
and U13270 (N_13270,N_12164,N_12230);
nand U13271 (N_13271,N_12320,N_12152);
xnor U13272 (N_13272,N_12357,N_12268);
nand U13273 (N_13273,N_12323,N_12529);
nor U13274 (N_13274,N_12722,N_12235);
xnor U13275 (N_13275,N_12234,N_12336);
and U13276 (N_13276,N_12127,N_12012);
nand U13277 (N_13277,N_12279,N_12381);
xor U13278 (N_13278,N_12509,N_12151);
nand U13279 (N_13279,N_12227,N_12087);
xor U13280 (N_13280,N_12153,N_12123);
and U13281 (N_13281,N_12411,N_12573);
or U13282 (N_13282,N_12471,N_12124);
and U13283 (N_13283,N_12639,N_12081);
nor U13284 (N_13284,N_12653,N_12120);
nor U13285 (N_13285,N_12000,N_12118);
and U13286 (N_13286,N_12050,N_12122);
xor U13287 (N_13287,N_12445,N_12473);
and U13288 (N_13288,N_12673,N_12529);
nand U13289 (N_13289,N_12067,N_12598);
or U13290 (N_13290,N_12601,N_12656);
or U13291 (N_13291,N_12298,N_12133);
nor U13292 (N_13292,N_12243,N_12349);
or U13293 (N_13293,N_12639,N_12050);
nand U13294 (N_13294,N_12020,N_12632);
nor U13295 (N_13295,N_12665,N_12152);
nand U13296 (N_13296,N_12150,N_12705);
nand U13297 (N_13297,N_12172,N_12682);
and U13298 (N_13298,N_12129,N_12607);
xor U13299 (N_13299,N_12483,N_12422);
and U13300 (N_13300,N_12237,N_12495);
nand U13301 (N_13301,N_12254,N_12498);
or U13302 (N_13302,N_12182,N_12677);
and U13303 (N_13303,N_12323,N_12531);
nor U13304 (N_13304,N_12376,N_12123);
and U13305 (N_13305,N_12701,N_12599);
nand U13306 (N_13306,N_12429,N_12396);
and U13307 (N_13307,N_12740,N_12196);
nand U13308 (N_13308,N_12042,N_12093);
nor U13309 (N_13309,N_12716,N_12349);
or U13310 (N_13310,N_12401,N_12186);
xnor U13311 (N_13311,N_12158,N_12380);
xor U13312 (N_13312,N_12295,N_12381);
nor U13313 (N_13313,N_12013,N_12463);
nor U13314 (N_13314,N_12522,N_12460);
and U13315 (N_13315,N_12336,N_12022);
and U13316 (N_13316,N_12026,N_12251);
nand U13317 (N_13317,N_12429,N_12260);
nor U13318 (N_13318,N_12495,N_12561);
nor U13319 (N_13319,N_12300,N_12485);
or U13320 (N_13320,N_12670,N_12744);
or U13321 (N_13321,N_12078,N_12007);
and U13322 (N_13322,N_12294,N_12060);
nand U13323 (N_13323,N_12189,N_12619);
xor U13324 (N_13324,N_12601,N_12604);
and U13325 (N_13325,N_12301,N_12328);
and U13326 (N_13326,N_12667,N_12384);
nand U13327 (N_13327,N_12249,N_12132);
or U13328 (N_13328,N_12562,N_12117);
nor U13329 (N_13329,N_12522,N_12378);
nor U13330 (N_13330,N_12675,N_12499);
and U13331 (N_13331,N_12174,N_12544);
and U13332 (N_13332,N_12689,N_12502);
and U13333 (N_13333,N_12071,N_12477);
xnor U13334 (N_13334,N_12389,N_12009);
nand U13335 (N_13335,N_12600,N_12518);
xor U13336 (N_13336,N_12528,N_12376);
nand U13337 (N_13337,N_12550,N_12368);
nand U13338 (N_13338,N_12231,N_12567);
nor U13339 (N_13339,N_12477,N_12215);
nand U13340 (N_13340,N_12668,N_12726);
and U13341 (N_13341,N_12101,N_12649);
xnor U13342 (N_13342,N_12014,N_12430);
nor U13343 (N_13343,N_12666,N_12619);
nand U13344 (N_13344,N_12252,N_12646);
or U13345 (N_13345,N_12240,N_12744);
xnor U13346 (N_13346,N_12171,N_12161);
or U13347 (N_13347,N_12638,N_12293);
xnor U13348 (N_13348,N_12388,N_12071);
nor U13349 (N_13349,N_12542,N_12586);
or U13350 (N_13350,N_12109,N_12692);
or U13351 (N_13351,N_12490,N_12375);
nor U13352 (N_13352,N_12321,N_12416);
and U13353 (N_13353,N_12661,N_12619);
nor U13354 (N_13354,N_12644,N_12210);
nor U13355 (N_13355,N_12351,N_12053);
nand U13356 (N_13356,N_12610,N_12513);
nor U13357 (N_13357,N_12474,N_12526);
nor U13358 (N_13358,N_12272,N_12381);
xor U13359 (N_13359,N_12663,N_12395);
xnor U13360 (N_13360,N_12745,N_12020);
nand U13361 (N_13361,N_12352,N_12012);
or U13362 (N_13362,N_12471,N_12131);
nand U13363 (N_13363,N_12593,N_12496);
nor U13364 (N_13364,N_12476,N_12203);
or U13365 (N_13365,N_12202,N_12416);
nor U13366 (N_13366,N_12385,N_12729);
and U13367 (N_13367,N_12443,N_12093);
nor U13368 (N_13368,N_12552,N_12135);
nand U13369 (N_13369,N_12612,N_12484);
or U13370 (N_13370,N_12596,N_12717);
nand U13371 (N_13371,N_12132,N_12160);
and U13372 (N_13372,N_12214,N_12407);
or U13373 (N_13373,N_12740,N_12372);
nor U13374 (N_13374,N_12728,N_12057);
nand U13375 (N_13375,N_12464,N_12461);
nand U13376 (N_13376,N_12124,N_12694);
or U13377 (N_13377,N_12406,N_12236);
or U13378 (N_13378,N_12037,N_12589);
or U13379 (N_13379,N_12258,N_12015);
nor U13380 (N_13380,N_12206,N_12047);
nor U13381 (N_13381,N_12148,N_12680);
nand U13382 (N_13382,N_12488,N_12342);
and U13383 (N_13383,N_12605,N_12638);
or U13384 (N_13384,N_12087,N_12307);
or U13385 (N_13385,N_12141,N_12173);
or U13386 (N_13386,N_12622,N_12264);
or U13387 (N_13387,N_12010,N_12555);
xnor U13388 (N_13388,N_12031,N_12121);
xor U13389 (N_13389,N_12464,N_12093);
and U13390 (N_13390,N_12242,N_12098);
and U13391 (N_13391,N_12643,N_12236);
and U13392 (N_13392,N_12359,N_12286);
nand U13393 (N_13393,N_12170,N_12493);
and U13394 (N_13394,N_12743,N_12399);
xnor U13395 (N_13395,N_12692,N_12242);
nor U13396 (N_13396,N_12640,N_12406);
nor U13397 (N_13397,N_12618,N_12200);
or U13398 (N_13398,N_12583,N_12250);
and U13399 (N_13399,N_12492,N_12610);
and U13400 (N_13400,N_12699,N_12372);
and U13401 (N_13401,N_12634,N_12506);
and U13402 (N_13402,N_12419,N_12564);
nor U13403 (N_13403,N_12061,N_12398);
or U13404 (N_13404,N_12369,N_12346);
nand U13405 (N_13405,N_12216,N_12676);
and U13406 (N_13406,N_12037,N_12452);
xnor U13407 (N_13407,N_12346,N_12253);
nand U13408 (N_13408,N_12354,N_12444);
or U13409 (N_13409,N_12011,N_12662);
or U13410 (N_13410,N_12603,N_12056);
nand U13411 (N_13411,N_12106,N_12181);
nand U13412 (N_13412,N_12415,N_12556);
or U13413 (N_13413,N_12184,N_12110);
or U13414 (N_13414,N_12592,N_12433);
and U13415 (N_13415,N_12327,N_12253);
or U13416 (N_13416,N_12551,N_12484);
nand U13417 (N_13417,N_12133,N_12379);
nand U13418 (N_13418,N_12238,N_12235);
or U13419 (N_13419,N_12120,N_12420);
and U13420 (N_13420,N_12002,N_12450);
nand U13421 (N_13421,N_12540,N_12525);
nor U13422 (N_13422,N_12464,N_12457);
or U13423 (N_13423,N_12488,N_12468);
nor U13424 (N_13424,N_12000,N_12074);
nor U13425 (N_13425,N_12102,N_12625);
nor U13426 (N_13426,N_12063,N_12549);
nand U13427 (N_13427,N_12408,N_12434);
nor U13428 (N_13428,N_12606,N_12081);
and U13429 (N_13429,N_12348,N_12174);
nand U13430 (N_13430,N_12733,N_12727);
and U13431 (N_13431,N_12621,N_12453);
xnor U13432 (N_13432,N_12016,N_12705);
xor U13433 (N_13433,N_12028,N_12366);
and U13434 (N_13434,N_12259,N_12580);
or U13435 (N_13435,N_12335,N_12064);
and U13436 (N_13436,N_12707,N_12483);
nand U13437 (N_13437,N_12356,N_12290);
and U13438 (N_13438,N_12409,N_12032);
nor U13439 (N_13439,N_12302,N_12155);
and U13440 (N_13440,N_12021,N_12522);
xor U13441 (N_13441,N_12118,N_12138);
nor U13442 (N_13442,N_12384,N_12579);
and U13443 (N_13443,N_12405,N_12102);
or U13444 (N_13444,N_12662,N_12125);
and U13445 (N_13445,N_12361,N_12539);
nand U13446 (N_13446,N_12021,N_12739);
nand U13447 (N_13447,N_12014,N_12741);
nor U13448 (N_13448,N_12110,N_12450);
or U13449 (N_13449,N_12150,N_12374);
nor U13450 (N_13450,N_12242,N_12418);
nand U13451 (N_13451,N_12674,N_12356);
or U13452 (N_13452,N_12307,N_12264);
xnor U13453 (N_13453,N_12034,N_12036);
xnor U13454 (N_13454,N_12142,N_12647);
nor U13455 (N_13455,N_12640,N_12021);
xnor U13456 (N_13456,N_12376,N_12506);
and U13457 (N_13457,N_12575,N_12430);
nand U13458 (N_13458,N_12090,N_12305);
nand U13459 (N_13459,N_12161,N_12626);
or U13460 (N_13460,N_12686,N_12377);
or U13461 (N_13461,N_12434,N_12190);
and U13462 (N_13462,N_12290,N_12073);
nor U13463 (N_13463,N_12656,N_12339);
or U13464 (N_13464,N_12700,N_12026);
nand U13465 (N_13465,N_12262,N_12101);
nand U13466 (N_13466,N_12387,N_12053);
nand U13467 (N_13467,N_12581,N_12062);
nand U13468 (N_13468,N_12018,N_12618);
or U13469 (N_13469,N_12136,N_12273);
and U13470 (N_13470,N_12681,N_12530);
or U13471 (N_13471,N_12591,N_12337);
and U13472 (N_13472,N_12411,N_12556);
xnor U13473 (N_13473,N_12622,N_12017);
or U13474 (N_13474,N_12334,N_12443);
or U13475 (N_13475,N_12624,N_12211);
and U13476 (N_13476,N_12454,N_12684);
nand U13477 (N_13477,N_12142,N_12284);
and U13478 (N_13478,N_12215,N_12174);
or U13479 (N_13479,N_12401,N_12028);
and U13480 (N_13480,N_12274,N_12449);
and U13481 (N_13481,N_12040,N_12621);
nor U13482 (N_13482,N_12152,N_12587);
or U13483 (N_13483,N_12543,N_12368);
or U13484 (N_13484,N_12062,N_12299);
xnor U13485 (N_13485,N_12262,N_12113);
xor U13486 (N_13486,N_12028,N_12361);
xnor U13487 (N_13487,N_12571,N_12019);
nor U13488 (N_13488,N_12581,N_12468);
nor U13489 (N_13489,N_12645,N_12691);
xnor U13490 (N_13490,N_12659,N_12322);
nor U13491 (N_13491,N_12649,N_12735);
nor U13492 (N_13492,N_12254,N_12688);
nand U13493 (N_13493,N_12704,N_12505);
nor U13494 (N_13494,N_12030,N_12673);
nand U13495 (N_13495,N_12667,N_12573);
nand U13496 (N_13496,N_12530,N_12556);
or U13497 (N_13497,N_12375,N_12056);
nand U13498 (N_13498,N_12153,N_12029);
and U13499 (N_13499,N_12424,N_12736);
and U13500 (N_13500,N_13378,N_13002);
and U13501 (N_13501,N_12839,N_13177);
nor U13502 (N_13502,N_13014,N_12964);
nor U13503 (N_13503,N_12899,N_13405);
and U13504 (N_13504,N_13183,N_13376);
and U13505 (N_13505,N_12872,N_12883);
xnor U13506 (N_13506,N_13036,N_13171);
xor U13507 (N_13507,N_13164,N_13069);
or U13508 (N_13508,N_13366,N_12820);
and U13509 (N_13509,N_13367,N_12846);
nand U13510 (N_13510,N_13438,N_13220);
and U13511 (N_13511,N_13187,N_13157);
and U13512 (N_13512,N_13267,N_13426);
nand U13513 (N_13513,N_13296,N_12802);
xnor U13514 (N_13514,N_13265,N_12879);
nand U13515 (N_13515,N_13065,N_13450);
nor U13516 (N_13516,N_13478,N_13218);
and U13517 (N_13517,N_12998,N_13354);
and U13518 (N_13518,N_13015,N_12909);
and U13519 (N_13519,N_12885,N_13027);
and U13520 (N_13520,N_12760,N_12962);
nor U13521 (N_13521,N_12835,N_13243);
nor U13522 (N_13522,N_13113,N_12776);
nand U13523 (N_13523,N_13138,N_12854);
and U13524 (N_13524,N_12871,N_13095);
xor U13525 (N_13525,N_13222,N_12956);
xnor U13526 (N_13526,N_13320,N_12795);
nor U13527 (N_13527,N_12764,N_13104);
nor U13528 (N_13528,N_12766,N_12780);
and U13529 (N_13529,N_12882,N_13055);
nand U13530 (N_13530,N_13353,N_13482);
or U13531 (N_13531,N_12751,N_13050);
nand U13532 (N_13532,N_13030,N_13312);
xor U13533 (N_13533,N_13175,N_13230);
or U13534 (N_13534,N_13043,N_12755);
and U13535 (N_13535,N_13213,N_13136);
nor U13536 (N_13536,N_12801,N_13270);
xor U13537 (N_13537,N_12877,N_13060);
nand U13538 (N_13538,N_12831,N_13392);
nand U13539 (N_13539,N_13262,N_13274);
or U13540 (N_13540,N_13217,N_12916);
or U13541 (N_13541,N_13051,N_12827);
or U13542 (N_13542,N_13108,N_13295);
and U13543 (N_13543,N_13266,N_13040);
and U13544 (N_13544,N_12804,N_12958);
nor U13545 (N_13545,N_13067,N_13035);
nand U13546 (N_13546,N_13017,N_13384);
nor U13547 (N_13547,N_13470,N_13097);
and U13548 (N_13548,N_12887,N_13469);
nor U13549 (N_13549,N_13440,N_13082);
nor U13550 (N_13550,N_13374,N_13464);
or U13551 (N_13551,N_13143,N_12915);
nand U13552 (N_13552,N_12913,N_13241);
or U13553 (N_13553,N_12767,N_12758);
nor U13554 (N_13554,N_12851,N_12934);
nor U13555 (N_13555,N_12946,N_13324);
xor U13556 (N_13556,N_13172,N_13049);
nand U13557 (N_13557,N_12828,N_13141);
and U13558 (N_13558,N_13176,N_13173);
nor U13559 (N_13559,N_13351,N_13386);
or U13560 (N_13560,N_13100,N_13417);
nand U13561 (N_13561,N_13323,N_13225);
or U13562 (N_13562,N_13037,N_12873);
nand U13563 (N_13563,N_13340,N_12930);
nor U13564 (N_13564,N_12898,N_13352);
and U13565 (N_13565,N_13076,N_13291);
nand U13566 (N_13566,N_13306,N_13336);
nor U13567 (N_13567,N_12972,N_12761);
and U13568 (N_13568,N_12895,N_12834);
xor U13569 (N_13569,N_12955,N_13019);
xor U13570 (N_13570,N_13091,N_12845);
nor U13571 (N_13571,N_13223,N_13140);
nand U13572 (N_13572,N_13471,N_13190);
xnor U13573 (N_13573,N_13166,N_12939);
or U13574 (N_13574,N_13335,N_13429);
or U13575 (N_13575,N_12847,N_13337);
nand U13576 (N_13576,N_13347,N_13345);
and U13577 (N_13577,N_12932,N_12999);
nand U13578 (N_13578,N_13093,N_13278);
nand U13579 (N_13579,N_13328,N_12823);
nor U13580 (N_13580,N_13348,N_13299);
nor U13581 (N_13581,N_13131,N_13293);
xor U13582 (N_13582,N_13467,N_12929);
or U13583 (N_13583,N_13031,N_13486);
nand U13584 (N_13584,N_13499,N_13480);
and U13585 (N_13585,N_12908,N_13297);
and U13586 (N_13586,N_13439,N_12791);
xnor U13587 (N_13587,N_12979,N_13282);
xor U13588 (N_13588,N_13192,N_13089);
and U13589 (N_13589,N_12790,N_13443);
nor U13590 (N_13590,N_13178,N_12922);
nor U13591 (N_13591,N_13156,N_13410);
nor U13592 (N_13592,N_13124,N_12772);
xnor U13593 (N_13593,N_12920,N_13044);
nand U13594 (N_13594,N_13033,N_12897);
nand U13595 (N_13595,N_13142,N_13441);
or U13596 (N_13596,N_12757,N_12797);
nand U13597 (N_13597,N_13459,N_13349);
or U13598 (N_13598,N_13198,N_13012);
nor U13599 (N_13599,N_13163,N_13445);
nand U13600 (N_13600,N_13102,N_13240);
nand U13601 (N_13601,N_13029,N_13462);
xor U13602 (N_13602,N_13111,N_13253);
and U13603 (N_13603,N_13059,N_13453);
and U13604 (N_13604,N_12952,N_13281);
or U13605 (N_13605,N_12902,N_13399);
and U13606 (N_13606,N_12807,N_13318);
or U13607 (N_13607,N_13269,N_13316);
and U13608 (N_13608,N_13403,N_13001);
and U13609 (N_13609,N_13412,N_13120);
xnor U13610 (N_13610,N_13125,N_13046);
nor U13611 (N_13611,N_12843,N_13304);
and U13612 (N_13612,N_12949,N_12901);
xor U13613 (N_13613,N_13331,N_12857);
and U13614 (N_13614,N_13333,N_13170);
nand U13615 (N_13615,N_12756,N_13208);
nor U13616 (N_13616,N_12866,N_12859);
nor U13617 (N_13617,N_13212,N_13202);
xor U13618 (N_13618,N_13382,N_13215);
nor U13619 (N_13619,N_12765,N_13083);
nor U13620 (N_13620,N_12960,N_12778);
nor U13621 (N_13621,N_13314,N_13342);
or U13622 (N_13622,N_12982,N_12973);
or U13623 (N_13623,N_12985,N_12918);
nand U13624 (N_13624,N_12842,N_13105);
nor U13625 (N_13625,N_13099,N_13381);
nor U13626 (N_13626,N_13309,N_13455);
and U13627 (N_13627,N_13279,N_13461);
nor U13628 (N_13628,N_13234,N_13451);
or U13629 (N_13629,N_13161,N_12833);
or U13630 (N_13630,N_13437,N_13368);
or U13631 (N_13631,N_13180,N_13427);
nand U13632 (N_13632,N_12775,N_12850);
and U13633 (N_13633,N_12925,N_13460);
nor U13634 (N_13634,N_13285,N_13448);
and U13635 (N_13635,N_12886,N_13498);
and U13636 (N_13636,N_13165,N_12841);
nand U13637 (N_13637,N_13492,N_12825);
and U13638 (N_13638,N_13396,N_13475);
or U13639 (N_13639,N_12974,N_13088);
xor U13640 (N_13640,N_12894,N_13435);
nor U13641 (N_13641,N_13228,N_13332);
or U13642 (N_13642,N_13497,N_13458);
and U13643 (N_13643,N_13226,N_13096);
nand U13644 (N_13644,N_13092,N_13139);
or U13645 (N_13645,N_13305,N_13114);
nor U13646 (N_13646,N_12869,N_12966);
xor U13647 (N_13647,N_12994,N_13193);
and U13648 (N_13648,N_13365,N_13020);
nor U13649 (N_13649,N_12941,N_13201);
or U13650 (N_13650,N_13231,N_12855);
nand U13651 (N_13651,N_12988,N_12983);
or U13652 (N_13652,N_13276,N_12799);
nand U13653 (N_13653,N_13123,N_13203);
nand U13654 (N_13654,N_12959,N_12837);
and U13655 (N_13655,N_13013,N_13160);
and U13656 (N_13656,N_12944,N_13235);
and U13657 (N_13657,N_13360,N_13275);
nor U13658 (N_13658,N_12811,N_13398);
xnor U13659 (N_13659,N_12923,N_12926);
nand U13660 (N_13660,N_12863,N_12808);
nand U13661 (N_13661,N_13256,N_12968);
xnor U13662 (N_13662,N_13434,N_12953);
and U13663 (N_13663,N_12870,N_13414);
nand U13664 (N_13664,N_12789,N_12906);
nor U13665 (N_13665,N_13152,N_12809);
xnor U13666 (N_13666,N_13327,N_13074);
nor U13667 (N_13667,N_13232,N_13409);
nor U13668 (N_13668,N_13456,N_13329);
xor U13669 (N_13669,N_13288,N_13185);
and U13670 (N_13670,N_12798,N_12992);
nor U13671 (N_13671,N_12907,N_13424);
and U13672 (N_13672,N_13310,N_13024);
or U13673 (N_13673,N_12943,N_13107);
and U13674 (N_13674,N_12975,N_12940);
xor U13675 (N_13675,N_13199,N_13390);
nand U13676 (N_13676,N_12969,N_13224);
and U13677 (N_13677,N_13144,N_13137);
and U13678 (N_13678,N_13210,N_13477);
nand U13679 (N_13679,N_12981,N_12754);
nand U13680 (N_13680,N_13388,N_13248);
nor U13681 (N_13681,N_13494,N_12884);
and U13682 (N_13682,N_12824,N_13292);
or U13683 (N_13683,N_13115,N_12840);
nor U13684 (N_13684,N_13472,N_12830);
or U13685 (N_13685,N_13106,N_12881);
or U13686 (N_13686,N_13389,N_12903);
nor U13687 (N_13687,N_12793,N_12832);
or U13688 (N_13688,N_13385,N_13380);
and U13689 (N_13689,N_13326,N_13425);
nor U13690 (N_13690,N_13442,N_13407);
nand U13691 (N_13691,N_12977,N_13122);
nand U13692 (N_13692,N_12878,N_12784);
nand U13693 (N_13693,N_13200,N_13130);
nor U13694 (N_13694,N_13416,N_13168);
nand U13695 (N_13695,N_13422,N_12875);
nor U13696 (N_13696,N_13487,N_12861);
and U13697 (N_13697,N_12947,N_13290);
xor U13698 (N_13698,N_13186,N_13155);
xnor U13699 (N_13699,N_13496,N_13028);
or U13700 (N_13700,N_13356,N_12812);
and U13701 (N_13701,N_13153,N_12770);
and U13702 (N_13702,N_13247,N_13406);
nor U13703 (N_13703,N_13188,N_12777);
nor U13704 (N_13704,N_13209,N_12800);
nand U13705 (N_13705,N_13007,N_13394);
and U13706 (N_13706,N_12971,N_13479);
nand U13707 (N_13707,N_12961,N_13261);
nor U13708 (N_13708,N_13358,N_13039);
nor U13709 (N_13709,N_13058,N_13286);
nand U13710 (N_13710,N_12876,N_13148);
xor U13711 (N_13711,N_12867,N_13132);
nor U13712 (N_13712,N_13084,N_12914);
nand U13713 (N_13713,N_13255,N_13117);
xor U13714 (N_13714,N_13362,N_13071);
or U13715 (N_13715,N_13154,N_13334);
nor U13716 (N_13716,N_12786,N_13041);
and U13717 (N_13717,N_13483,N_13118);
or U13718 (N_13718,N_13465,N_13421);
nor U13719 (N_13719,N_13229,N_12888);
nor U13720 (N_13720,N_13109,N_13308);
nand U13721 (N_13721,N_12810,N_13449);
nand U13722 (N_13722,N_13116,N_13463);
nand U13723 (N_13723,N_13008,N_13061);
or U13724 (N_13724,N_12821,N_12905);
nor U13725 (N_13725,N_13404,N_13227);
or U13726 (N_13726,N_13273,N_13488);
or U13727 (N_13727,N_13271,N_13221);
nand U13728 (N_13728,N_13135,N_13101);
or U13729 (N_13729,N_13493,N_12788);
xor U13730 (N_13730,N_13194,N_13257);
nor U13731 (N_13731,N_12816,N_12917);
or U13732 (N_13732,N_13476,N_13303);
nand U13733 (N_13733,N_13211,N_12814);
nand U13734 (N_13734,N_12904,N_13025);
or U13735 (N_13735,N_13289,N_12792);
and U13736 (N_13736,N_12794,N_12750);
xor U13737 (N_13737,N_13436,N_13466);
nand U13738 (N_13738,N_12989,N_13119);
or U13739 (N_13739,N_13103,N_13151);
xor U13740 (N_13740,N_13233,N_13485);
and U13741 (N_13741,N_13249,N_12889);
nand U13742 (N_13742,N_13127,N_13204);
nand U13743 (N_13743,N_12782,N_13397);
nor U13744 (N_13744,N_12938,N_13149);
nand U13745 (N_13745,N_13189,N_13056);
or U13746 (N_13746,N_12951,N_13361);
and U13747 (N_13747,N_12819,N_13016);
or U13748 (N_13748,N_13245,N_13242);
nor U13749 (N_13749,N_13034,N_13315);
nor U13750 (N_13750,N_12954,N_13045);
or U13751 (N_13751,N_13359,N_13181);
or U13752 (N_13752,N_13018,N_13128);
or U13753 (N_13753,N_13073,N_13005);
nor U13754 (N_13754,N_12928,N_12817);
nand U13755 (N_13755,N_13010,N_13430);
nand U13756 (N_13756,N_13158,N_12900);
nor U13757 (N_13757,N_13263,N_12993);
and U13758 (N_13758,N_12924,N_12838);
nand U13759 (N_13759,N_12921,N_13004);
nand U13760 (N_13760,N_13495,N_13003);
nor U13761 (N_13761,N_13377,N_13444);
nand U13762 (N_13762,N_13419,N_13393);
nand U13763 (N_13763,N_12933,N_12984);
nor U13764 (N_13764,N_13064,N_13090);
and U13765 (N_13765,N_13167,N_13207);
nor U13766 (N_13766,N_12768,N_12779);
and U13767 (N_13767,N_13150,N_13277);
or U13768 (N_13768,N_13047,N_13077);
nand U13769 (N_13769,N_12759,N_13085);
or U13770 (N_13770,N_12848,N_13284);
nor U13771 (N_13771,N_13447,N_13283);
and U13772 (N_13772,N_13259,N_12781);
nor U13773 (N_13773,N_13490,N_13294);
nor U13774 (N_13774,N_13006,N_12976);
or U13775 (N_13775,N_13110,N_13147);
xor U13776 (N_13776,N_13317,N_12844);
and U13777 (N_13777,N_13428,N_12911);
and U13778 (N_13778,N_13216,N_12948);
and U13779 (N_13779,N_13344,N_13330);
nor U13780 (N_13780,N_13054,N_13489);
nand U13781 (N_13781,N_12815,N_12783);
xnor U13782 (N_13782,N_13357,N_12919);
nor U13783 (N_13783,N_13302,N_12860);
nor U13784 (N_13784,N_13338,N_12856);
and U13785 (N_13785,N_13134,N_13264);
xnor U13786 (N_13786,N_12796,N_12890);
nand U13787 (N_13787,N_13048,N_12997);
nor U13788 (N_13788,N_12785,N_13068);
nor U13789 (N_13789,N_12862,N_13280);
and U13790 (N_13790,N_13057,N_13179);
or U13791 (N_13791,N_13371,N_13042);
nand U13792 (N_13792,N_13395,N_12752);
and U13793 (N_13793,N_12963,N_13402);
and U13794 (N_13794,N_13238,N_13319);
xnor U13795 (N_13795,N_13184,N_12950);
nand U13796 (N_13796,N_12990,N_13370);
xnor U13797 (N_13797,N_13379,N_13053);
and U13798 (N_13798,N_13086,N_13237);
and U13799 (N_13799,N_12853,N_13411);
nor U13800 (N_13800,N_13433,N_13219);
xor U13801 (N_13801,N_12836,N_13011);
xor U13802 (N_13802,N_12806,N_13454);
nand U13803 (N_13803,N_13133,N_13321);
nand U13804 (N_13804,N_12822,N_13491);
xnor U13805 (N_13805,N_13174,N_12763);
or U13806 (N_13806,N_13474,N_13313);
or U13807 (N_13807,N_13457,N_13250);
nand U13808 (N_13808,N_13387,N_13126);
and U13809 (N_13809,N_13446,N_13206);
nand U13810 (N_13810,N_12864,N_13363);
nor U13811 (N_13811,N_12970,N_12892);
or U13812 (N_13812,N_13169,N_12927);
and U13813 (N_13813,N_13072,N_13159);
nor U13814 (N_13814,N_12868,N_13298);
nor U13815 (N_13815,N_13346,N_12935);
nor U13816 (N_13816,N_12995,N_13418);
nor U13817 (N_13817,N_13300,N_13239);
and U13818 (N_13818,N_12967,N_12880);
nand U13819 (N_13819,N_13272,N_12896);
nand U13820 (N_13820,N_13355,N_13009);
nand U13821 (N_13821,N_13078,N_12945);
nand U13822 (N_13822,N_13214,N_12891);
nor U13823 (N_13823,N_13162,N_12937);
nor U13824 (N_13824,N_13258,N_12978);
nor U13825 (N_13825,N_13066,N_13038);
nand U13826 (N_13826,N_13121,N_12813);
and U13827 (N_13827,N_13252,N_13484);
nor U13828 (N_13828,N_13023,N_13022);
nand U13829 (N_13829,N_12826,N_13400);
nor U13830 (N_13830,N_13431,N_13063);
or U13831 (N_13831,N_13081,N_12858);
nor U13832 (N_13832,N_12980,N_13000);
nor U13833 (N_13833,N_13191,N_13244);
or U13834 (N_13834,N_12986,N_12805);
xor U13835 (N_13835,N_13420,N_13468);
nor U13836 (N_13836,N_13205,N_12803);
and U13837 (N_13837,N_13146,N_12773);
nor U13838 (N_13838,N_13287,N_13254);
nand U13839 (N_13839,N_13375,N_13094);
or U13840 (N_13840,N_13087,N_13075);
nor U13841 (N_13841,N_13112,N_13021);
or U13842 (N_13842,N_13364,N_13341);
nand U13843 (N_13843,N_12849,N_13372);
nand U13844 (N_13844,N_12852,N_13423);
xnor U13845 (N_13845,N_12874,N_12829);
or U13846 (N_13846,N_13268,N_12942);
nand U13847 (N_13847,N_13401,N_13260);
and U13848 (N_13848,N_13413,N_12787);
or U13849 (N_13849,N_12912,N_12753);
and U13850 (N_13850,N_13473,N_12865);
or U13851 (N_13851,N_13481,N_13098);
nor U13852 (N_13852,N_13452,N_13236);
and U13853 (N_13853,N_13052,N_13343);
xor U13854 (N_13854,N_13246,N_13251);
xnor U13855 (N_13855,N_13026,N_12771);
and U13856 (N_13856,N_12987,N_13383);
nor U13857 (N_13857,N_13129,N_12818);
nor U13858 (N_13858,N_13391,N_13070);
nor U13859 (N_13859,N_12769,N_12762);
nand U13860 (N_13860,N_13432,N_12965);
and U13861 (N_13861,N_13325,N_13079);
and U13862 (N_13862,N_13350,N_13301);
nor U13863 (N_13863,N_12893,N_13062);
or U13864 (N_13864,N_13032,N_13373);
or U13865 (N_13865,N_12931,N_13408);
or U13866 (N_13866,N_13197,N_13415);
nand U13867 (N_13867,N_13182,N_13339);
nand U13868 (N_13868,N_13322,N_13195);
nand U13869 (N_13869,N_12957,N_13307);
xnor U13870 (N_13870,N_12910,N_13145);
or U13871 (N_13871,N_12774,N_13311);
nor U13872 (N_13872,N_13196,N_12991);
or U13873 (N_13873,N_12996,N_13369);
or U13874 (N_13874,N_13080,N_12936);
nand U13875 (N_13875,N_13344,N_12858);
nand U13876 (N_13876,N_13236,N_13042);
nor U13877 (N_13877,N_13323,N_13113);
nand U13878 (N_13878,N_13395,N_13041);
or U13879 (N_13879,N_13020,N_13206);
or U13880 (N_13880,N_13288,N_13418);
and U13881 (N_13881,N_12883,N_12800);
or U13882 (N_13882,N_12899,N_13457);
and U13883 (N_13883,N_12967,N_12988);
nand U13884 (N_13884,N_13345,N_13387);
and U13885 (N_13885,N_13122,N_13193);
nand U13886 (N_13886,N_12908,N_13393);
or U13887 (N_13887,N_13332,N_13401);
nand U13888 (N_13888,N_13310,N_13122);
nor U13889 (N_13889,N_12966,N_12763);
and U13890 (N_13890,N_12909,N_12906);
or U13891 (N_13891,N_13096,N_12991);
nand U13892 (N_13892,N_12787,N_12922);
or U13893 (N_13893,N_13480,N_13339);
nand U13894 (N_13894,N_12949,N_13368);
and U13895 (N_13895,N_13271,N_13462);
xnor U13896 (N_13896,N_12940,N_12777);
nand U13897 (N_13897,N_12764,N_13252);
or U13898 (N_13898,N_13147,N_13393);
and U13899 (N_13899,N_13002,N_12853);
nor U13900 (N_13900,N_13018,N_12789);
and U13901 (N_13901,N_12891,N_13323);
and U13902 (N_13902,N_13446,N_13372);
or U13903 (N_13903,N_13327,N_13356);
and U13904 (N_13904,N_12965,N_13105);
nand U13905 (N_13905,N_13300,N_13317);
and U13906 (N_13906,N_13252,N_12801);
nor U13907 (N_13907,N_13006,N_12848);
nor U13908 (N_13908,N_13207,N_13409);
nor U13909 (N_13909,N_12900,N_13357);
nand U13910 (N_13910,N_12978,N_12954);
nand U13911 (N_13911,N_13448,N_12905);
nor U13912 (N_13912,N_13206,N_13365);
or U13913 (N_13913,N_13471,N_13047);
nor U13914 (N_13914,N_13407,N_13444);
nor U13915 (N_13915,N_12791,N_13097);
xnor U13916 (N_13916,N_12844,N_13301);
nand U13917 (N_13917,N_13269,N_13480);
or U13918 (N_13918,N_12774,N_12924);
or U13919 (N_13919,N_13258,N_12827);
or U13920 (N_13920,N_12774,N_13305);
or U13921 (N_13921,N_12850,N_13398);
nor U13922 (N_13922,N_13033,N_13096);
nand U13923 (N_13923,N_12778,N_13350);
and U13924 (N_13924,N_13052,N_12947);
or U13925 (N_13925,N_13421,N_12759);
and U13926 (N_13926,N_13267,N_13285);
nor U13927 (N_13927,N_13311,N_13113);
nand U13928 (N_13928,N_13165,N_13331);
or U13929 (N_13929,N_13082,N_13305);
nor U13930 (N_13930,N_12989,N_12915);
or U13931 (N_13931,N_13126,N_12790);
or U13932 (N_13932,N_13257,N_13427);
nand U13933 (N_13933,N_13161,N_13076);
nor U13934 (N_13934,N_12943,N_13074);
nand U13935 (N_13935,N_12791,N_13054);
nor U13936 (N_13936,N_13424,N_13402);
nand U13937 (N_13937,N_12881,N_12909);
or U13938 (N_13938,N_13288,N_13001);
or U13939 (N_13939,N_13430,N_13117);
nand U13940 (N_13940,N_13363,N_12967);
nor U13941 (N_13941,N_13118,N_13392);
and U13942 (N_13942,N_12772,N_12969);
nand U13943 (N_13943,N_13447,N_13145);
nand U13944 (N_13944,N_13004,N_12965);
nor U13945 (N_13945,N_13080,N_12934);
or U13946 (N_13946,N_13084,N_12799);
and U13947 (N_13947,N_12909,N_13408);
or U13948 (N_13948,N_12932,N_13183);
and U13949 (N_13949,N_13029,N_13002);
and U13950 (N_13950,N_12971,N_12877);
or U13951 (N_13951,N_13099,N_13037);
or U13952 (N_13952,N_13347,N_13172);
or U13953 (N_13953,N_13365,N_13154);
and U13954 (N_13954,N_13488,N_13296);
and U13955 (N_13955,N_13352,N_12929);
or U13956 (N_13956,N_12803,N_13024);
or U13957 (N_13957,N_12788,N_12794);
and U13958 (N_13958,N_13054,N_12951);
nor U13959 (N_13959,N_13018,N_13169);
nor U13960 (N_13960,N_12773,N_12754);
and U13961 (N_13961,N_13050,N_13047);
or U13962 (N_13962,N_13181,N_13190);
and U13963 (N_13963,N_12785,N_13367);
xor U13964 (N_13964,N_13180,N_13033);
or U13965 (N_13965,N_13158,N_13062);
nor U13966 (N_13966,N_13374,N_12817);
xnor U13967 (N_13967,N_13432,N_12878);
nor U13968 (N_13968,N_13431,N_13041);
and U13969 (N_13969,N_13080,N_12928);
xor U13970 (N_13970,N_13253,N_12839);
xor U13971 (N_13971,N_13379,N_12810);
and U13972 (N_13972,N_13288,N_13038);
nand U13973 (N_13973,N_13138,N_13435);
nor U13974 (N_13974,N_13303,N_13077);
xor U13975 (N_13975,N_13139,N_12772);
or U13976 (N_13976,N_12921,N_12974);
nor U13977 (N_13977,N_13287,N_13059);
and U13978 (N_13978,N_13385,N_13172);
nor U13979 (N_13979,N_13139,N_13179);
and U13980 (N_13980,N_13470,N_12891);
nand U13981 (N_13981,N_13328,N_13019);
nand U13982 (N_13982,N_13127,N_12958);
or U13983 (N_13983,N_13161,N_13298);
or U13984 (N_13984,N_13114,N_13326);
or U13985 (N_13985,N_12982,N_13200);
and U13986 (N_13986,N_13307,N_13317);
and U13987 (N_13987,N_13106,N_13383);
or U13988 (N_13988,N_13359,N_13410);
xor U13989 (N_13989,N_12897,N_12806);
xor U13990 (N_13990,N_12815,N_12838);
and U13991 (N_13991,N_13338,N_12812);
or U13992 (N_13992,N_12822,N_12819);
nor U13993 (N_13993,N_13292,N_12967);
and U13994 (N_13994,N_13474,N_13260);
xnor U13995 (N_13995,N_12864,N_13271);
and U13996 (N_13996,N_12813,N_12791);
or U13997 (N_13997,N_12902,N_12945);
xnor U13998 (N_13998,N_13455,N_13295);
or U13999 (N_13999,N_12811,N_13421);
and U14000 (N_14000,N_12775,N_13282);
or U14001 (N_14001,N_13438,N_12909);
nor U14002 (N_14002,N_12957,N_13237);
nand U14003 (N_14003,N_13247,N_13091);
and U14004 (N_14004,N_13040,N_13405);
nor U14005 (N_14005,N_13120,N_13208);
or U14006 (N_14006,N_12833,N_13029);
and U14007 (N_14007,N_12849,N_13030);
nor U14008 (N_14008,N_13227,N_12912);
nand U14009 (N_14009,N_13217,N_13163);
or U14010 (N_14010,N_12985,N_12764);
xnor U14011 (N_14011,N_12898,N_13117);
and U14012 (N_14012,N_12915,N_13172);
nand U14013 (N_14013,N_12966,N_12947);
and U14014 (N_14014,N_13201,N_13446);
nor U14015 (N_14015,N_12821,N_13110);
or U14016 (N_14016,N_12864,N_13262);
or U14017 (N_14017,N_13486,N_12820);
or U14018 (N_14018,N_13328,N_13151);
or U14019 (N_14019,N_13178,N_13255);
nand U14020 (N_14020,N_13363,N_12752);
and U14021 (N_14021,N_12989,N_13338);
or U14022 (N_14022,N_13315,N_13466);
nor U14023 (N_14023,N_13499,N_13258);
or U14024 (N_14024,N_13491,N_13496);
and U14025 (N_14025,N_13069,N_13151);
or U14026 (N_14026,N_13272,N_13094);
nor U14027 (N_14027,N_13342,N_12771);
or U14028 (N_14028,N_13179,N_12901);
xor U14029 (N_14029,N_12928,N_12864);
and U14030 (N_14030,N_13087,N_13271);
nand U14031 (N_14031,N_13072,N_12982);
and U14032 (N_14032,N_13347,N_12779);
nor U14033 (N_14033,N_13097,N_13456);
or U14034 (N_14034,N_13363,N_13470);
or U14035 (N_14035,N_13417,N_13416);
nor U14036 (N_14036,N_13047,N_13245);
or U14037 (N_14037,N_13481,N_13061);
xor U14038 (N_14038,N_13215,N_13028);
nor U14039 (N_14039,N_12882,N_13420);
nand U14040 (N_14040,N_13116,N_13091);
nor U14041 (N_14041,N_12921,N_13476);
and U14042 (N_14042,N_12912,N_13426);
or U14043 (N_14043,N_13275,N_13254);
and U14044 (N_14044,N_13399,N_12892);
and U14045 (N_14045,N_12813,N_13166);
nand U14046 (N_14046,N_13126,N_13351);
nor U14047 (N_14047,N_12896,N_12822);
nor U14048 (N_14048,N_13324,N_13404);
and U14049 (N_14049,N_13197,N_13053);
or U14050 (N_14050,N_12972,N_13186);
nand U14051 (N_14051,N_13040,N_12850);
nand U14052 (N_14052,N_13314,N_12831);
nor U14053 (N_14053,N_12825,N_13423);
nor U14054 (N_14054,N_13048,N_12860);
nor U14055 (N_14055,N_13435,N_13264);
and U14056 (N_14056,N_13309,N_13034);
or U14057 (N_14057,N_13188,N_13201);
or U14058 (N_14058,N_13378,N_13326);
nor U14059 (N_14059,N_12897,N_13405);
or U14060 (N_14060,N_12816,N_12984);
nor U14061 (N_14061,N_13179,N_13040);
nor U14062 (N_14062,N_13071,N_13050);
nand U14063 (N_14063,N_12781,N_13055);
and U14064 (N_14064,N_13273,N_12902);
nor U14065 (N_14065,N_12980,N_13456);
or U14066 (N_14066,N_12894,N_12989);
nand U14067 (N_14067,N_13221,N_13091);
and U14068 (N_14068,N_13274,N_13064);
nand U14069 (N_14069,N_13177,N_13133);
xor U14070 (N_14070,N_12827,N_13010);
or U14071 (N_14071,N_13419,N_13228);
or U14072 (N_14072,N_12963,N_13372);
or U14073 (N_14073,N_13113,N_12840);
and U14074 (N_14074,N_13383,N_13184);
or U14075 (N_14075,N_13486,N_13408);
and U14076 (N_14076,N_13482,N_13472);
and U14077 (N_14077,N_13476,N_12862);
xnor U14078 (N_14078,N_13077,N_12754);
nand U14079 (N_14079,N_13191,N_13277);
and U14080 (N_14080,N_12762,N_13118);
and U14081 (N_14081,N_12846,N_13370);
nor U14082 (N_14082,N_12997,N_13434);
and U14083 (N_14083,N_13433,N_13205);
xnor U14084 (N_14084,N_13458,N_13171);
nor U14085 (N_14085,N_12983,N_13186);
or U14086 (N_14086,N_13134,N_13233);
and U14087 (N_14087,N_12879,N_13229);
nor U14088 (N_14088,N_13415,N_13221);
nor U14089 (N_14089,N_13141,N_13328);
and U14090 (N_14090,N_13396,N_12870);
and U14091 (N_14091,N_13278,N_13434);
and U14092 (N_14092,N_12882,N_13070);
and U14093 (N_14093,N_13371,N_13267);
and U14094 (N_14094,N_12856,N_13214);
and U14095 (N_14095,N_12846,N_13297);
xor U14096 (N_14096,N_12885,N_13132);
nor U14097 (N_14097,N_12753,N_12821);
and U14098 (N_14098,N_13056,N_12826);
and U14099 (N_14099,N_12899,N_13410);
nand U14100 (N_14100,N_12868,N_13078);
xor U14101 (N_14101,N_12965,N_13454);
xor U14102 (N_14102,N_13290,N_12994);
or U14103 (N_14103,N_12988,N_13040);
nand U14104 (N_14104,N_12772,N_13182);
or U14105 (N_14105,N_13430,N_13401);
and U14106 (N_14106,N_13411,N_13488);
and U14107 (N_14107,N_12955,N_13495);
and U14108 (N_14108,N_13389,N_12994);
and U14109 (N_14109,N_12935,N_12775);
or U14110 (N_14110,N_13307,N_13111);
or U14111 (N_14111,N_13449,N_13356);
and U14112 (N_14112,N_12762,N_13284);
nor U14113 (N_14113,N_12790,N_13287);
nor U14114 (N_14114,N_12823,N_13134);
and U14115 (N_14115,N_13219,N_13441);
nand U14116 (N_14116,N_12779,N_13427);
nor U14117 (N_14117,N_12985,N_12765);
nand U14118 (N_14118,N_12796,N_13267);
nor U14119 (N_14119,N_13474,N_13178);
nand U14120 (N_14120,N_13051,N_13207);
or U14121 (N_14121,N_12767,N_13261);
nand U14122 (N_14122,N_12991,N_13305);
nand U14123 (N_14123,N_13001,N_13134);
or U14124 (N_14124,N_13116,N_12957);
nand U14125 (N_14125,N_13278,N_13095);
nor U14126 (N_14126,N_12956,N_12752);
nor U14127 (N_14127,N_13022,N_12881);
and U14128 (N_14128,N_13178,N_13423);
nand U14129 (N_14129,N_13387,N_12892);
xnor U14130 (N_14130,N_13476,N_12926);
or U14131 (N_14131,N_12836,N_12826);
xor U14132 (N_14132,N_12865,N_13135);
and U14133 (N_14133,N_12907,N_13132);
nand U14134 (N_14134,N_13397,N_13179);
and U14135 (N_14135,N_13215,N_13173);
or U14136 (N_14136,N_12999,N_12986);
and U14137 (N_14137,N_12904,N_12770);
or U14138 (N_14138,N_13080,N_12954);
and U14139 (N_14139,N_13323,N_13132);
xnor U14140 (N_14140,N_12763,N_12908);
and U14141 (N_14141,N_13352,N_13148);
and U14142 (N_14142,N_13095,N_13450);
or U14143 (N_14143,N_13084,N_13447);
or U14144 (N_14144,N_12976,N_13467);
or U14145 (N_14145,N_13117,N_13195);
nand U14146 (N_14146,N_13179,N_13343);
nand U14147 (N_14147,N_13357,N_12836);
xnor U14148 (N_14148,N_12866,N_12858);
or U14149 (N_14149,N_13085,N_13232);
or U14150 (N_14150,N_13449,N_12798);
nand U14151 (N_14151,N_12760,N_12936);
nor U14152 (N_14152,N_12938,N_13328);
nor U14153 (N_14153,N_12899,N_13339);
nor U14154 (N_14154,N_12773,N_13347);
nand U14155 (N_14155,N_12905,N_13055);
and U14156 (N_14156,N_12917,N_13226);
or U14157 (N_14157,N_13078,N_13207);
nor U14158 (N_14158,N_13356,N_12921);
nor U14159 (N_14159,N_12803,N_12898);
or U14160 (N_14160,N_13051,N_13315);
or U14161 (N_14161,N_13186,N_13097);
xnor U14162 (N_14162,N_12897,N_12769);
nand U14163 (N_14163,N_12923,N_13170);
nand U14164 (N_14164,N_13416,N_13040);
nor U14165 (N_14165,N_12781,N_13091);
or U14166 (N_14166,N_13012,N_13245);
nand U14167 (N_14167,N_13439,N_12801);
xor U14168 (N_14168,N_13230,N_13083);
or U14169 (N_14169,N_13345,N_13149);
and U14170 (N_14170,N_13047,N_13021);
nor U14171 (N_14171,N_13181,N_12813);
nand U14172 (N_14172,N_12882,N_13186);
nor U14173 (N_14173,N_13275,N_12910);
nor U14174 (N_14174,N_13257,N_13386);
nor U14175 (N_14175,N_13154,N_13483);
nor U14176 (N_14176,N_13405,N_13381);
and U14177 (N_14177,N_13335,N_12841);
xor U14178 (N_14178,N_13137,N_13217);
and U14179 (N_14179,N_13320,N_12902);
and U14180 (N_14180,N_13205,N_12816);
nor U14181 (N_14181,N_13400,N_13135);
nand U14182 (N_14182,N_13134,N_13423);
nand U14183 (N_14183,N_13334,N_13280);
nand U14184 (N_14184,N_13286,N_13437);
or U14185 (N_14185,N_12859,N_13388);
and U14186 (N_14186,N_13351,N_13129);
nand U14187 (N_14187,N_13038,N_13439);
nor U14188 (N_14188,N_13202,N_13234);
or U14189 (N_14189,N_12969,N_12776);
nand U14190 (N_14190,N_12874,N_13312);
and U14191 (N_14191,N_13079,N_12943);
or U14192 (N_14192,N_12952,N_12753);
nand U14193 (N_14193,N_13468,N_13485);
nor U14194 (N_14194,N_12760,N_13394);
xor U14195 (N_14195,N_13025,N_13088);
nor U14196 (N_14196,N_13071,N_13465);
nor U14197 (N_14197,N_13358,N_13154);
or U14198 (N_14198,N_13074,N_13212);
nand U14199 (N_14199,N_12845,N_13327);
nor U14200 (N_14200,N_12784,N_12761);
nand U14201 (N_14201,N_12957,N_13071);
or U14202 (N_14202,N_13090,N_12908);
and U14203 (N_14203,N_13408,N_13384);
or U14204 (N_14204,N_12888,N_13166);
and U14205 (N_14205,N_12955,N_13485);
nor U14206 (N_14206,N_13227,N_13260);
nand U14207 (N_14207,N_13348,N_13235);
nand U14208 (N_14208,N_13411,N_12872);
nor U14209 (N_14209,N_12799,N_12774);
nand U14210 (N_14210,N_13268,N_13291);
nand U14211 (N_14211,N_13100,N_13342);
xor U14212 (N_14212,N_13333,N_12962);
and U14213 (N_14213,N_13454,N_12765);
nor U14214 (N_14214,N_13355,N_12996);
and U14215 (N_14215,N_13330,N_13283);
nand U14216 (N_14216,N_13475,N_13361);
or U14217 (N_14217,N_13099,N_12987);
and U14218 (N_14218,N_13285,N_13056);
and U14219 (N_14219,N_12832,N_12970);
nor U14220 (N_14220,N_13358,N_12895);
nor U14221 (N_14221,N_13006,N_13467);
and U14222 (N_14222,N_13201,N_12829);
or U14223 (N_14223,N_13317,N_13271);
or U14224 (N_14224,N_13251,N_12756);
nor U14225 (N_14225,N_12980,N_13286);
nor U14226 (N_14226,N_13229,N_13420);
and U14227 (N_14227,N_13457,N_13037);
nor U14228 (N_14228,N_13125,N_13355);
and U14229 (N_14229,N_13092,N_12836);
xor U14230 (N_14230,N_13370,N_13494);
nor U14231 (N_14231,N_13048,N_12930);
or U14232 (N_14232,N_13346,N_13135);
or U14233 (N_14233,N_13381,N_13352);
nor U14234 (N_14234,N_12871,N_13383);
nand U14235 (N_14235,N_13162,N_13382);
and U14236 (N_14236,N_13208,N_13181);
nor U14237 (N_14237,N_13027,N_13064);
and U14238 (N_14238,N_12927,N_13182);
nor U14239 (N_14239,N_13155,N_13220);
or U14240 (N_14240,N_12995,N_13327);
or U14241 (N_14241,N_13023,N_13365);
nor U14242 (N_14242,N_13204,N_12977);
nor U14243 (N_14243,N_13105,N_12922);
and U14244 (N_14244,N_13048,N_12918);
nor U14245 (N_14245,N_12960,N_13012);
or U14246 (N_14246,N_13385,N_13166);
or U14247 (N_14247,N_12924,N_12902);
xor U14248 (N_14248,N_13309,N_13490);
or U14249 (N_14249,N_12860,N_13106);
nand U14250 (N_14250,N_14081,N_14170);
and U14251 (N_14251,N_13827,N_14171);
nor U14252 (N_14252,N_13985,N_13734);
nand U14253 (N_14253,N_13737,N_14208);
or U14254 (N_14254,N_13910,N_13668);
nor U14255 (N_14255,N_13689,N_13508);
nor U14256 (N_14256,N_13535,N_14231);
xnor U14257 (N_14257,N_14247,N_13916);
nand U14258 (N_14258,N_14203,N_13748);
and U14259 (N_14259,N_14098,N_13659);
or U14260 (N_14260,N_13915,N_13775);
and U14261 (N_14261,N_13681,N_13701);
nor U14262 (N_14262,N_13988,N_13740);
nand U14263 (N_14263,N_14040,N_13601);
and U14264 (N_14264,N_13556,N_13928);
nand U14265 (N_14265,N_13519,N_14192);
nor U14266 (N_14266,N_13547,N_14046);
nor U14267 (N_14267,N_13699,N_13750);
or U14268 (N_14268,N_13595,N_13686);
or U14269 (N_14269,N_13691,N_13936);
and U14270 (N_14270,N_13784,N_14063);
nor U14271 (N_14271,N_13708,N_14165);
nor U14272 (N_14272,N_13912,N_13986);
or U14273 (N_14273,N_13887,N_14018);
nand U14274 (N_14274,N_14093,N_13884);
or U14275 (N_14275,N_14177,N_14058);
nand U14276 (N_14276,N_14119,N_13729);
nor U14277 (N_14277,N_13941,N_14014);
and U14278 (N_14278,N_13777,N_13837);
or U14279 (N_14279,N_13977,N_13832);
nand U14280 (N_14280,N_14054,N_13611);
and U14281 (N_14281,N_13579,N_14109);
or U14282 (N_14282,N_13888,N_14186);
or U14283 (N_14283,N_13581,N_13880);
nand U14284 (N_14284,N_13706,N_14175);
nand U14285 (N_14285,N_13931,N_14049);
and U14286 (N_14286,N_13656,N_14095);
or U14287 (N_14287,N_13692,N_13939);
or U14288 (N_14288,N_13690,N_13546);
or U14289 (N_14289,N_13603,N_13637);
nand U14290 (N_14290,N_13695,N_13548);
xnor U14291 (N_14291,N_14114,N_13920);
nor U14292 (N_14292,N_14075,N_13516);
and U14293 (N_14293,N_14073,N_14166);
nand U14294 (N_14294,N_13966,N_13505);
and U14295 (N_14295,N_13719,N_13904);
and U14296 (N_14296,N_14009,N_13746);
or U14297 (N_14297,N_13620,N_14090);
and U14298 (N_14298,N_14085,N_13964);
and U14299 (N_14299,N_13869,N_14199);
nor U14300 (N_14300,N_13864,N_14172);
nor U14301 (N_14301,N_14108,N_14005);
nor U14302 (N_14302,N_13545,N_14002);
and U14303 (N_14303,N_14178,N_13862);
or U14304 (N_14304,N_14047,N_13513);
nor U14305 (N_14305,N_13895,N_13510);
nand U14306 (N_14306,N_13707,N_13630);
nand U14307 (N_14307,N_14056,N_14068);
nand U14308 (N_14308,N_13634,N_14244);
or U14309 (N_14309,N_13532,N_13772);
xor U14310 (N_14310,N_13756,N_13974);
nand U14311 (N_14311,N_13802,N_13660);
xor U14312 (N_14312,N_14154,N_13696);
xor U14313 (N_14313,N_13543,N_13657);
nor U14314 (N_14314,N_13865,N_13716);
nor U14315 (N_14315,N_13918,N_13623);
xor U14316 (N_14316,N_13615,N_13585);
nand U14317 (N_14317,N_14230,N_13724);
nor U14318 (N_14318,N_14023,N_13945);
or U14319 (N_14319,N_14156,N_14245);
nand U14320 (N_14320,N_13676,N_13963);
nor U14321 (N_14321,N_13859,N_13504);
nand U14322 (N_14322,N_13886,N_13671);
nand U14323 (N_14323,N_14234,N_13577);
nand U14324 (N_14324,N_13744,N_13683);
xor U14325 (N_14325,N_13749,N_13572);
nor U14326 (N_14326,N_13952,N_13726);
nand U14327 (N_14327,N_13848,N_13534);
and U14328 (N_14328,N_13860,N_13942);
xnor U14329 (N_14329,N_13835,N_13600);
nor U14330 (N_14330,N_14238,N_14224);
nor U14331 (N_14331,N_14115,N_13815);
or U14332 (N_14332,N_13760,N_13927);
nand U14333 (N_14333,N_14039,N_13979);
nand U14334 (N_14334,N_13639,N_13751);
nor U14335 (N_14335,N_13998,N_13826);
xor U14336 (N_14336,N_14001,N_13560);
or U14337 (N_14337,N_13608,N_14248);
and U14338 (N_14338,N_13995,N_13822);
nor U14339 (N_14339,N_13563,N_14129);
nand U14340 (N_14340,N_13787,N_13654);
and U14341 (N_14341,N_14089,N_14028);
and U14342 (N_14342,N_13984,N_14216);
or U14343 (N_14343,N_14173,N_13541);
and U14344 (N_14344,N_14149,N_13538);
nor U14345 (N_14345,N_13664,N_13843);
nand U14346 (N_14346,N_14038,N_13967);
nand U14347 (N_14347,N_13885,N_13584);
or U14348 (N_14348,N_13901,N_13764);
nand U14349 (N_14349,N_13844,N_13622);
or U14350 (N_14350,N_13854,N_14083);
nand U14351 (N_14351,N_13809,N_13562);
and U14352 (N_14352,N_13644,N_14221);
xor U14353 (N_14353,N_13769,N_14176);
and U14354 (N_14354,N_13833,N_13721);
nand U14355 (N_14355,N_13900,N_13576);
and U14356 (N_14356,N_13774,N_13602);
xor U14357 (N_14357,N_14074,N_13632);
nor U14358 (N_14358,N_14196,N_13930);
nand U14359 (N_14359,N_13621,N_13828);
nand U14360 (N_14360,N_14008,N_13536);
nor U14361 (N_14361,N_14032,N_13793);
nand U14362 (N_14362,N_13643,N_13962);
nand U14363 (N_14363,N_13717,N_13728);
xor U14364 (N_14364,N_13530,N_13528);
nand U14365 (N_14365,N_13825,N_13551);
xor U14366 (N_14366,N_14194,N_13741);
and U14367 (N_14367,N_14134,N_13819);
and U14368 (N_14368,N_13669,N_13851);
or U14369 (N_14369,N_13824,N_14019);
nor U14370 (N_14370,N_13583,N_13976);
or U14371 (N_14371,N_13993,N_14117);
nor U14372 (N_14372,N_13882,N_13629);
nor U14373 (N_14373,N_13540,N_14213);
and U14374 (N_14374,N_13898,N_14107);
and U14375 (N_14375,N_13727,N_13514);
or U14376 (N_14376,N_13883,N_14029);
or U14377 (N_14377,N_14010,N_13703);
and U14378 (N_14378,N_13983,N_13752);
nand U14379 (N_14379,N_13868,N_13924);
xnor U14380 (N_14380,N_14144,N_13596);
nor U14381 (N_14381,N_13588,N_14239);
nand U14382 (N_14382,N_13926,N_13982);
and U14383 (N_14383,N_13732,N_13618);
nor U14384 (N_14384,N_14209,N_13817);
nor U14385 (N_14385,N_13960,N_13934);
and U14386 (N_14386,N_14204,N_13768);
nor U14387 (N_14387,N_13838,N_13839);
and U14388 (N_14388,N_13569,N_13881);
or U14389 (N_14389,N_13943,N_14103);
nor U14390 (N_14390,N_13627,N_13761);
nor U14391 (N_14391,N_13892,N_14214);
nand U14392 (N_14392,N_13914,N_13571);
nand U14393 (N_14393,N_14079,N_13821);
nand U14394 (N_14394,N_14077,N_13574);
or U14395 (N_14395,N_13994,N_14101);
nor U14396 (N_14396,N_13520,N_13872);
and U14397 (N_14397,N_13709,N_13972);
and U14398 (N_14398,N_13790,N_13922);
nand U14399 (N_14399,N_14207,N_13811);
nor U14400 (N_14400,N_13568,N_14059);
nand U14401 (N_14401,N_13720,N_13636);
or U14402 (N_14402,N_13804,N_13711);
or U14403 (N_14403,N_13559,N_13938);
nor U14404 (N_14404,N_14048,N_14035);
or U14405 (N_14405,N_13978,N_14210);
nor U14406 (N_14406,N_14030,N_14223);
nand U14407 (N_14407,N_13841,N_13929);
nor U14408 (N_14408,N_14243,N_13788);
nor U14409 (N_14409,N_13778,N_13905);
nand U14410 (N_14410,N_14169,N_14004);
and U14411 (N_14411,N_13682,N_14088);
or U14412 (N_14412,N_14227,N_13723);
xnor U14413 (N_14413,N_13614,N_13705);
nor U14414 (N_14414,N_14220,N_13968);
or U14415 (N_14415,N_14132,N_13628);
xnor U14416 (N_14416,N_13502,N_14128);
and U14417 (N_14417,N_14122,N_14064);
nand U14418 (N_14418,N_13797,N_13521);
nor U14419 (N_14419,N_13786,N_13800);
nor U14420 (N_14420,N_13799,N_13575);
nor U14421 (N_14421,N_14148,N_13511);
nand U14422 (N_14422,N_13919,N_13987);
or U14423 (N_14423,N_13680,N_13873);
nand U14424 (N_14424,N_13863,N_13955);
and U14425 (N_14425,N_13891,N_13996);
nor U14426 (N_14426,N_13758,N_14226);
xor U14427 (N_14427,N_14195,N_14218);
or U14428 (N_14428,N_13694,N_13566);
and U14429 (N_14429,N_14229,N_13911);
xor U14430 (N_14430,N_14102,N_14065);
or U14431 (N_14431,N_14147,N_13889);
nor U14432 (N_14432,N_13619,N_13874);
nor U14433 (N_14433,N_14016,N_14205);
and U14434 (N_14434,N_14110,N_14164);
nor U14435 (N_14435,N_13949,N_13606);
nand U14436 (N_14436,N_14161,N_13808);
nand U14437 (N_14437,N_13879,N_13806);
nand U14438 (N_14438,N_13655,N_14201);
and U14439 (N_14439,N_14105,N_13529);
and U14440 (N_14440,N_14111,N_13959);
or U14441 (N_14441,N_14136,N_13567);
and U14442 (N_14442,N_13624,N_13858);
or U14443 (N_14443,N_14120,N_14100);
nor U14444 (N_14444,N_13794,N_14168);
and U14445 (N_14445,N_13907,N_13507);
nor U14446 (N_14446,N_13923,N_14106);
nor U14447 (N_14447,N_13714,N_13743);
and U14448 (N_14448,N_14139,N_14055);
or U14449 (N_14449,N_13625,N_13965);
nor U14450 (N_14450,N_13524,N_14141);
xor U14451 (N_14451,N_14211,N_13702);
nand U14452 (N_14452,N_13876,N_13616);
nor U14453 (N_14453,N_14249,N_14027);
nand U14454 (N_14454,N_13957,N_13947);
or U14455 (N_14455,N_13853,N_14159);
nand U14456 (N_14456,N_14133,N_13552);
nand U14457 (N_14457,N_13757,N_13755);
nor U14458 (N_14458,N_13688,N_14037);
or U14459 (N_14459,N_13766,N_13666);
and U14460 (N_14460,N_13554,N_13836);
or U14461 (N_14461,N_13753,N_13733);
and U14462 (N_14462,N_13792,N_14190);
or U14463 (N_14463,N_14033,N_13807);
nor U14464 (N_14464,N_14062,N_13948);
and U14465 (N_14465,N_13813,N_14225);
or U14466 (N_14466,N_13593,N_14092);
nand U14467 (N_14467,N_13971,N_13570);
or U14468 (N_14468,N_13670,N_13877);
or U14469 (N_14469,N_14042,N_13674);
nand U14470 (N_14470,N_14096,N_14124);
nand U14471 (N_14471,N_13903,N_13932);
or U14472 (N_14472,N_13896,N_14069);
xor U14473 (N_14473,N_14003,N_13771);
xor U14474 (N_14474,N_13626,N_13767);
and U14475 (N_14475,N_14024,N_13649);
nand U14476 (N_14476,N_13801,N_13782);
nand U14477 (N_14477,N_13846,N_13565);
nand U14478 (N_14478,N_13635,N_13798);
xnor U14479 (N_14479,N_13899,N_13849);
nor U14480 (N_14480,N_14142,N_13871);
nor U14481 (N_14481,N_13515,N_13745);
nand U14482 (N_14482,N_13954,N_13875);
or U14483 (N_14483,N_13940,N_13999);
nor U14484 (N_14484,N_13679,N_13506);
or U14485 (N_14485,N_13677,N_13693);
nand U14486 (N_14486,N_13578,N_13557);
and U14487 (N_14487,N_13715,N_13830);
xor U14488 (N_14488,N_14097,N_13573);
and U14489 (N_14489,N_13867,N_14104);
nand U14490 (N_14490,N_14091,N_13989);
xnor U14491 (N_14491,N_14200,N_14246);
xnor U14492 (N_14492,N_14094,N_13975);
or U14493 (N_14493,N_13598,N_13653);
nand U14494 (N_14494,N_13725,N_14180);
and U14495 (N_14495,N_13834,N_13651);
or U14496 (N_14496,N_13731,N_14241);
nand U14497 (N_14497,N_13990,N_14015);
xnor U14498 (N_14498,N_14053,N_14181);
nand U14499 (N_14499,N_14183,N_13522);
nor U14500 (N_14500,N_13509,N_14125);
and U14501 (N_14501,N_13555,N_14121);
or U14502 (N_14502,N_14151,N_13564);
nand U14503 (N_14503,N_13890,N_14152);
or U14504 (N_14504,N_13527,N_13549);
and U14505 (N_14505,N_13878,N_14113);
nand U14506 (N_14506,N_13742,N_14212);
nor U14507 (N_14507,N_13662,N_13776);
nor U14508 (N_14508,N_14153,N_13908);
nand U14509 (N_14509,N_13542,N_13517);
nand U14510 (N_14510,N_14140,N_13533);
or U14511 (N_14511,N_13631,N_14137);
xnor U14512 (N_14512,N_14011,N_13779);
or U14513 (N_14513,N_13944,N_14017);
nand U14514 (N_14514,N_14116,N_13902);
nand U14515 (N_14515,N_14127,N_13870);
xnor U14516 (N_14516,N_13645,N_13638);
nand U14517 (N_14517,N_13582,N_13921);
and U14518 (N_14518,N_13970,N_13823);
nand U14519 (N_14519,N_13640,N_13780);
nor U14520 (N_14520,N_13847,N_13712);
nand U14521 (N_14521,N_13531,N_13933);
and U14522 (N_14522,N_14187,N_13605);
nand U14523 (N_14523,N_13909,N_14236);
or U14524 (N_14524,N_13526,N_13818);
nand U14525 (N_14525,N_13673,N_13935);
nor U14526 (N_14526,N_14143,N_14242);
nand U14527 (N_14527,N_14045,N_13857);
nand U14528 (N_14528,N_13658,N_13539);
nand U14529 (N_14529,N_14219,N_14232);
nor U14530 (N_14530,N_13675,N_13704);
xnor U14531 (N_14531,N_14007,N_14070);
nor U14532 (N_14532,N_14000,N_14162);
or U14533 (N_14533,N_14076,N_13893);
nor U14534 (N_14534,N_13597,N_13544);
nor U14535 (N_14535,N_13650,N_14157);
nand U14536 (N_14536,N_13866,N_13917);
or U14537 (N_14537,N_14179,N_13550);
nand U14538 (N_14538,N_13642,N_14036);
or U14539 (N_14539,N_13894,N_13558);
nand U14540 (N_14540,N_13759,N_14202);
nand U14541 (N_14541,N_13855,N_14051);
nor U14542 (N_14542,N_13861,N_13661);
nand U14543 (N_14543,N_13617,N_13961);
and U14544 (N_14544,N_14057,N_14044);
and U14545 (N_14545,N_13814,N_13805);
nor U14546 (N_14546,N_14158,N_13913);
and U14547 (N_14547,N_13652,N_13958);
xnor U14548 (N_14548,N_13796,N_14021);
and U14549 (N_14549,N_13803,N_13773);
and U14550 (N_14550,N_13586,N_13770);
and U14551 (N_14551,N_13648,N_14123);
or U14552 (N_14552,N_13840,N_13604);
or U14553 (N_14553,N_13633,N_14061);
nand U14554 (N_14554,N_13747,N_13845);
xnor U14555 (N_14555,N_14185,N_13980);
xnor U14556 (N_14556,N_13785,N_13946);
nand U14557 (N_14557,N_13810,N_13997);
nand U14558 (N_14558,N_14198,N_13981);
nor U14559 (N_14559,N_13697,N_13641);
xor U14560 (N_14560,N_13763,N_13500);
nand U14561 (N_14561,N_13525,N_14163);
and U14562 (N_14562,N_14084,N_13739);
nand U14563 (N_14563,N_13684,N_14174);
nor U14564 (N_14564,N_13523,N_14233);
and U14565 (N_14565,N_13783,N_13698);
nor U14566 (N_14566,N_13592,N_13850);
nand U14567 (N_14567,N_14167,N_14071);
nand U14568 (N_14568,N_14012,N_14067);
xnor U14569 (N_14569,N_13580,N_13816);
and U14570 (N_14570,N_14182,N_14222);
nor U14571 (N_14571,N_13587,N_13736);
xnor U14572 (N_14572,N_13937,N_13722);
nor U14573 (N_14573,N_14112,N_14034);
nand U14574 (N_14574,N_13735,N_13906);
xor U14575 (N_14575,N_14118,N_13594);
and U14576 (N_14576,N_14082,N_13607);
nand U14577 (N_14577,N_13647,N_13973);
and U14578 (N_14578,N_14066,N_13503);
xnor U14579 (N_14579,N_14240,N_14184);
or U14580 (N_14580,N_14193,N_14135);
and U14581 (N_14581,N_13561,N_13537);
or U14582 (N_14582,N_14197,N_14155);
or U14583 (N_14583,N_14189,N_13738);
nand U14584 (N_14584,N_14041,N_13512);
nand U14585 (N_14585,N_14080,N_13992);
nor U14586 (N_14586,N_14206,N_14099);
nor U14587 (N_14587,N_14217,N_13956);
nor U14588 (N_14588,N_14026,N_14022);
nand U14589 (N_14589,N_13820,N_13754);
or U14590 (N_14590,N_13609,N_13951);
xor U14591 (N_14591,N_13842,N_13665);
or U14592 (N_14592,N_14087,N_13646);
nor U14593 (N_14593,N_13700,N_13829);
and U14594 (N_14594,N_14126,N_13791);
and U14595 (N_14595,N_14145,N_14060);
nor U14596 (N_14596,N_13765,N_13518);
xor U14597 (N_14597,N_14235,N_13762);
xnor U14598 (N_14598,N_14160,N_13991);
nand U14599 (N_14599,N_14146,N_13667);
nor U14600 (N_14600,N_13856,N_13672);
and U14601 (N_14601,N_14086,N_14215);
and U14602 (N_14602,N_14078,N_13610);
or U14603 (N_14603,N_13599,N_13678);
and U14604 (N_14604,N_13795,N_13969);
nand U14605 (N_14605,N_14072,N_13501);
nand U14606 (N_14606,N_13925,N_13831);
nor U14607 (N_14607,N_14052,N_14228);
and U14608 (N_14608,N_13663,N_14050);
nand U14609 (N_14609,N_13950,N_14006);
and U14610 (N_14610,N_13812,N_13953);
or U14611 (N_14611,N_13589,N_14031);
nand U14612 (N_14612,N_13781,N_13553);
and U14613 (N_14613,N_13718,N_13590);
or U14614 (N_14614,N_13852,N_14130);
and U14615 (N_14615,N_13897,N_14020);
xnor U14616 (N_14616,N_13789,N_14150);
nor U14617 (N_14617,N_14191,N_13687);
or U14618 (N_14618,N_14013,N_13685);
and U14619 (N_14619,N_13713,N_14188);
xnor U14620 (N_14620,N_13591,N_13710);
and U14621 (N_14621,N_14131,N_13730);
nor U14622 (N_14622,N_14237,N_13612);
or U14623 (N_14623,N_13613,N_14138);
nand U14624 (N_14624,N_14025,N_14043);
nor U14625 (N_14625,N_13837,N_13901);
nor U14626 (N_14626,N_13905,N_13710);
or U14627 (N_14627,N_14074,N_13958);
nor U14628 (N_14628,N_13606,N_13722);
and U14629 (N_14629,N_13593,N_13834);
and U14630 (N_14630,N_14145,N_14083);
nor U14631 (N_14631,N_14141,N_13832);
nor U14632 (N_14632,N_13738,N_13716);
or U14633 (N_14633,N_14165,N_13538);
nand U14634 (N_14634,N_14167,N_13538);
nand U14635 (N_14635,N_14164,N_14090);
and U14636 (N_14636,N_13618,N_13980);
or U14637 (N_14637,N_14172,N_14082);
nor U14638 (N_14638,N_13912,N_13571);
nand U14639 (N_14639,N_13527,N_14148);
and U14640 (N_14640,N_14233,N_13741);
nor U14641 (N_14641,N_14150,N_14053);
and U14642 (N_14642,N_13806,N_13845);
or U14643 (N_14643,N_13863,N_13933);
nor U14644 (N_14644,N_13948,N_13666);
or U14645 (N_14645,N_13500,N_13580);
and U14646 (N_14646,N_13730,N_13726);
and U14647 (N_14647,N_13845,N_13542);
nor U14648 (N_14648,N_13923,N_14089);
nor U14649 (N_14649,N_14221,N_13857);
and U14650 (N_14650,N_13705,N_13728);
and U14651 (N_14651,N_13671,N_13948);
and U14652 (N_14652,N_14205,N_13510);
and U14653 (N_14653,N_14014,N_13537);
and U14654 (N_14654,N_13877,N_13921);
nand U14655 (N_14655,N_13722,N_14025);
or U14656 (N_14656,N_13938,N_13603);
nand U14657 (N_14657,N_13934,N_13810);
nand U14658 (N_14658,N_13652,N_14027);
or U14659 (N_14659,N_14205,N_13612);
or U14660 (N_14660,N_13758,N_14030);
nor U14661 (N_14661,N_13775,N_14220);
xnor U14662 (N_14662,N_13569,N_13756);
nor U14663 (N_14663,N_13743,N_13662);
and U14664 (N_14664,N_14056,N_13882);
nand U14665 (N_14665,N_13923,N_13954);
xor U14666 (N_14666,N_13565,N_13709);
and U14667 (N_14667,N_14090,N_13650);
or U14668 (N_14668,N_14112,N_13814);
nand U14669 (N_14669,N_14018,N_13513);
or U14670 (N_14670,N_13518,N_13677);
nand U14671 (N_14671,N_14230,N_13859);
and U14672 (N_14672,N_13748,N_13832);
and U14673 (N_14673,N_13710,N_13766);
and U14674 (N_14674,N_13779,N_13567);
or U14675 (N_14675,N_13955,N_13673);
nand U14676 (N_14676,N_14062,N_13907);
nor U14677 (N_14677,N_13712,N_14047);
and U14678 (N_14678,N_13878,N_13711);
or U14679 (N_14679,N_13723,N_14151);
and U14680 (N_14680,N_14146,N_14151);
nor U14681 (N_14681,N_13608,N_14207);
or U14682 (N_14682,N_14202,N_13970);
and U14683 (N_14683,N_14031,N_13674);
xor U14684 (N_14684,N_13759,N_13563);
nor U14685 (N_14685,N_13856,N_14221);
and U14686 (N_14686,N_13607,N_13568);
or U14687 (N_14687,N_14039,N_13892);
and U14688 (N_14688,N_13636,N_13794);
nand U14689 (N_14689,N_13530,N_14097);
and U14690 (N_14690,N_13800,N_14129);
or U14691 (N_14691,N_13957,N_13837);
xnor U14692 (N_14692,N_13735,N_13514);
xor U14693 (N_14693,N_14244,N_14023);
and U14694 (N_14694,N_14046,N_13663);
nand U14695 (N_14695,N_14005,N_14097);
and U14696 (N_14696,N_13780,N_13687);
nand U14697 (N_14697,N_13972,N_13595);
or U14698 (N_14698,N_14092,N_14112);
nor U14699 (N_14699,N_13613,N_13666);
xnor U14700 (N_14700,N_13906,N_13609);
and U14701 (N_14701,N_14206,N_14004);
and U14702 (N_14702,N_14145,N_13616);
or U14703 (N_14703,N_14003,N_13903);
nand U14704 (N_14704,N_14001,N_13678);
nand U14705 (N_14705,N_14152,N_14059);
and U14706 (N_14706,N_13844,N_13935);
nor U14707 (N_14707,N_13540,N_14161);
and U14708 (N_14708,N_13995,N_13839);
or U14709 (N_14709,N_13505,N_14160);
or U14710 (N_14710,N_13537,N_14088);
and U14711 (N_14711,N_13578,N_13994);
nor U14712 (N_14712,N_14112,N_13869);
and U14713 (N_14713,N_14079,N_13760);
nor U14714 (N_14714,N_13539,N_13762);
nand U14715 (N_14715,N_14169,N_13757);
nand U14716 (N_14716,N_13631,N_14106);
or U14717 (N_14717,N_14183,N_13718);
nand U14718 (N_14718,N_13871,N_13712);
nand U14719 (N_14719,N_13764,N_13800);
xnor U14720 (N_14720,N_13921,N_13938);
and U14721 (N_14721,N_14072,N_13737);
nor U14722 (N_14722,N_13542,N_13610);
or U14723 (N_14723,N_14085,N_13911);
and U14724 (N_14724,N_14005,N_13632);
nor U14725 (N_14725,N_13555,N_14074);
nand U14726 (N_14726,N_14088,N_13509);
xnor U14727 (N_14727,N_13935,N_13700);
and U14728 (N_14728,N_14116,N_14224);
nor U14729 (N_14729,N_14167,N_13837);
and U14730 (N_14730,N_13607,N_13644);
nor U14731 (N_14731,N_14102,N_13564);
or U14732 (N_14732,N_14176,N_13572);
and U14733 (N_14733,N_14141,N_13988);
and U14734 (N_14734,N_13542,N_13867);
or U14735 (N_14735,N_14005,N_13919);
nor U14736 (N_14736,N_13508,N_13616);
nand U14737 (N_14737,N_13887,N_13741);
and U14738 (N_14738,N_13583,N_14208);
nand U14739 (N_14739,N_14213,N_13736);
or U14740 (N_14740,N_13643,N_14192);
nand U14741 (N_14741,N_13520,N_13580);
or U14742 (N_14742,N_14178,N_13653);
and U14743 (N_14743,N_13673,N_14155);
or U14744 (N_14744,N_13563,N_13682);
or U14745 (N_14745,N_13545,N_13795);
xor U14746 (N_14746,N_13590,N_14028);
nor U14747 (N_14747,N_14077,N_14155);
nand U14748 (N_14748,N_13867,N_13892);
nor U14749 (N_14749,N_14231,N_14189);
and U14750 (N_14750,N_13723,N_13847);
and U14751 (N_14751,N_13582,N_13730);
nand U14752 (N_14752,N_13737,N_14199);
nor U14753 (N_14753,N_13787,N_14003);
nand U14754 (N_14754,N_13625,N_13929);
nor U14755 (N_14755,N_13700,N_14166);
nor U14756 (N_14756,N_14155,N_13657);
nand U14757 (N_14757,N_13700,N_14070);
and U14758 (N_14758,N_14200,N_13731);
nand U14759 (N_14759,N_13590,N_13631);
nand U14760 (N_14760,N_14217,N_14068);
nand U14761 (N_14761,N_14217,N_13990);
and U14762 (N_14762,N_14049,N_14244);
or U14763 (N_14763,N_14215,N_13596);
or U14764 (N_14764,N_13526,N_13953);
nand U14765 (N_14765,N_13726,N_14021);
nor U14766 (N_14766,N_14203,N_13554);
nand U14767 (N_14767,N_13813,N_13821);
xnor U14768 (N_14768,N_14142,N_14106);
nand U14769 (N_14769,N_13850,N_13664);
or U14770 (N_14770,N_14006,N_14170);
nor U14771 (N_14771,N_14192,N_14118);
nand U14772 (N_14772,N_14017,N_13843);
and U14773 (N_14773,N_14028,N_14241);
and U14774 (N_14774,N_13868,N_13738);
and U14775 (N_14775,N_14212,N_14006);
or U14776 (N_14776,N_13942,N_13670);
xnor U14777 (N_14777,N_13744,N_13591);
and U14778 (N_14778,N_13629,N_13919);
and U14779 (N_14779,N_13810,N_14162);
nor U14780 (N_14780,N_13926,N_14020);
nor U14781 (N_14781,N_13613,N_13960);
and U14782 (N_14782,N_13988,N_14013);
and U14783 (N_14783,N_13569,N_13791);
and U14784 (N_14784,N_13863,N_13575);
nor U14785 (N_14785,N_14029,N_14112);
and U14786 (N_14786,N_14050,N_13684);
nand U14787 (N_14787,N_13884,N_13594);
nor U14788 (N_14788,N_13708,N_13797);
nand U14789 (N_14789,N_14159,N_13609);
or U14790 (N_14790,N_13694,N_13526);
and U14791 (N_14791,N_14016,N_13652);
or U14792 (N_14792,N_14076,N_13541);
or U14793 (N_14793,N_13704,N_13906);
nor U14794 (N_14794,N_14059,N_13824);
or U14795 (N_14795,N_13840,N_14022);
nor U14796 (N_14796,N_14235,N_13675);
nand U14797 (N_14797,N_13957,N_13968);
nor U14798 (N_14798,N_13766,N_13873);
or U14799 (N_14799,N_13911,N_13862);
or U14800 (N_14800,N_13576,N_13557);
or U14801 (N_14801,N_14058,N_13665);
nor U14802 (N_14802,N_13635,N_13688);
nor U14803 (N_14803,N_13733,N_14209);
and U14804 (N_14804,N_13645,N_13800);
and U14805 (N_14805,N_14137,N_13816);
nor U14806 (N_14806,N_14125,N_13844);
and U14807 (N_14807,N_14168,N_13958);
and U14808 (N_14808,N_13624,N_14142);
nor U14809 (N_14809,N_13779,N_13916);
xnor U14810 (N_14810,N_13863,N_13851);
or U14811 (N_14811,N_13709,N_14070);
nor U14812 (N_14812,N_14184,N_14105);
nor U14813 (N_14813,N_14010,N_14055);
nor U14814 (N_14814,N_14190,N_13674);
and U14815 (N_14815,N_13740,N_13923);
nand U14816 (N_14816,N_13658,N_14086);
and U14817 (N_14817,N_14246,N_14026);
xnor U14818 (N_14818,N_14015,N_13865);
or U14819 (N_14819,N_13967,N_14062);
xnor U14820 (N_14820,N_14240,N_13990);
and U14821 (N_14821,N_13512,N_14225);
nand U14822 (N_14822,N_14076,N_13606);
or U14823 (N_14823,N_14155,N_13723);
nand U14824 (N_14824,N_13626,N_13578);
nor U14825 (N_14825,N_13883,N_14062);
and U14826 (N_14826,N_13587,N_13597);
nor U14827 (N_14827,N_13894,N_13718);
or U14828 (N_14828,N_13824,N_13599);
xnor U14829 (N_14829,N_13891,N_13692);
nand U14830 (N_14830,N_13951,N_13606);
and U14831 (N_14831,N_13786,N_13662);
and U14832 (N_14832,N_14092,N_14231);
and U14833 (N_14833,N_13715,N_13939);
nor U14834 (N_14834,N_13544,N_13532);
and U14835 (N_14835,N_13849,N_14012);
or U14836 (N_14836,N_13937,N_13799);
nor U14837 (N_14837,N_13674,N_14049);
nor U14838 (N_14838,N_14232,N_14200);
nor U14839 (N_14839,N_13609,N_14249);
nor U14840 (N_14840,N_13763,N_13691);
and U14841 (N_14841,N_13880,N_13803);
and U14842 (N_14842,N_13544,N_13746);
or U14843 (N_14843,N_14136,N_13532);
or U14844 (N_14844,N_14162,N_14224);
nor U14845 (N_14845,N_13667,N_13852);
or U14846 (N_14846,N_13686,N_13914);
nand U14847 (N_14847,N_13881,N_14146);
and U14848 (N_14848,N_13715,N_13951);
or U14849 (N_14849,N_13716,N_14127);
nor U14850 (N_14850,N_13859,N_13576);
and U14851 (N_14851,N_14245,N_13746);
xor U14852 (N_14852,N_14077,N_13605);
nor U14853 (N_14853,N_13605,N_13872);
nand U14854 (N_14854,N_13726,N_13650);
xnor U14855 (N_14855,N_14045,N_13814);
or U14856 (N_14856,N_13787,N_13730);
and U14857 (N_14857,N_13816,N_13629);
xnor U14858 (N_14858,N_13669,N_14237);
nor U14859 (N_14859,N_14071,N_14038);
or U14860 (N_14860,N_13882,N_13528);
xnor U14861 (N_14861,N_14195,N_13606);
and U14862 (N_14862,N_13915,N_14103);
nand U14863 (N_14863,N_13571,N_14247);
or U14864 (N_14864,N_14184,N_13612);
nand U14865 (N_14865,N_14139,N_13776);
and U14866 (N_14866,N_14216,N_13723);
or U14867 (N_14867,N_14169,N_13570);
and U14868 (N_14868,N_14045,N_13648);
xnor U14869 (N_14869,N_13634,N_13673);
and U14870 (N_14870,N_13892,N_14095);
xnor U14871 (N_14871,N_13900,N_14050);
xor U14872 (N_14872,N_14226,N_13737);
nor U14873 (N_14873,N_14233,N_13999);
nor U14874 (N_14874,N_13867,N_14091);
or U14875 (N_14875,N_13843,N_13637);
nor U14876 (N_14876,N_14100,N_13635);
nor U14877 (N_14877,N_14241,N_14230);
and U14878 (N_14878,N_14151,N_13544);
xnor U14879 (N_14879,N_13508,N_13646);
or U14880 (N_14880,N_14171,N_13739);
and U14881 (N_14881,N_13865,N_13997);
and U14882 (N_14882,N_14226,N_13766);
nand U14883 (N_14883,N_13685,N_13980);
or U14884 (N_14884,N_14148,N_14198);
or U14885 (N_14885,N_13952,N_13738);
nor U14886 (N_14886,N_13890,N_14140);
nand U14887 (N_14887,N_14229,N_14071);
xor U14888 (N_14888,N_14153,N_14061);
nand U14889 (N_14889,N_13580,N_13791);
or U14890 (N_14890,N_13680,N_14216);
nor U14891 (N_14891,N_13912,N_13715);
nor U14892 (N_14892,N_13654,N_13593);
or U14893 (N_14893,N_13831,N_14228);
xor U14894 (N_14894,N_13968,N_14224);
nor U14895 (N_14895,N_14191,N_13972);
or U14896 (N_14896,N_13827,N_14080);
nand U14897 (N_14897,N_13899,N_14066);
nand U14898 (N_14898,N_14089,N_14155);
and U14899 (N_14899,N_13606,N_13910);
nand U14900 (N_14900,N_13777,N_14120);
nand U14901 (N_14901,N_13882,N_13902);
nor U14902 (N_14902,N_13851,N_13760);
and U14903 (N_14903,N_14169,N_14044);
or U14904 (N_14904,N_13954,N_14101);
and U14905 (N_14905,N_13542,N_13741);
and U14906 (N_14906,N_13825,N_14010);
and U14907 (N_14907,N_14101,N_13970);
nand U14908 (N_14908,N_14247,N_14114);
nor U14909 (N_14909,N_13718,N_14096);
and U14910 (N_14910,N_13792,N_13930);
or U14911 (N_14911,N_13652,N_14146);
nor U14912 (N_14912,N_14172,N_13625);
and U14913 (N_14913,N_13586,N_13633);
and U14914 (N_14914,N_14222,N_13734);
nor U14915 (N_14915,N_13637,N_13905);
nand U14916 (N_14916,N_13885,N_13534);
nor U14917 (N_14917,N_13941,N_13667);
nand U14918 (N_14918,N_13502,N_13660);
or U14919 (N_14919,N_14220,N_13996);
or U14920 (N_14920,N_13508,N_13870);
or U14921 (N_14921,N_13663,N_14021);
nor U14922 (N_14922,N_13514,N_13833);
and U14923 (N_14923,N_13698,N_13824);
and U14924 (N_14924,N_13979,N_14007);
nand U14925 (N_14925,N_13858,N_14001);
and U14926 (N_14926,N_14004,N_14170);
xnor U14927 (N_14927,N_13651,N_14076);
nand U14928 (N_14928,N_14109,N_13799);
or U14929 (N_14929,N_13602,N_14101);
or U14930 (N_14930,N_13852,N_13884);
nor U14931 (N_14931,N_13546,N_13526);
nand U14932 (N_14932,N_14149,N_14246);
nand U14933 (N_14933,N_13686,N_13533);
nand U14934 (N_14934,N_14018,N_13707);
nand U14935 (N_14935,N_14117,N_14152);
nor U14936 (N_14936,N_13932,N_14113);
and U14937 (N_14937,N_14003,N_14212);
or U14938 (N_14938,N_13630,N_14167);
or U14939 (N_14939,N_14025,N_13828);
nor U14940 (N_14940,N_14213,N_14059);
nor U14941 (N_14941,N_13503,N_13564);
nand U14942 (N_14942,N_13717,N_14126);
or U14943 (N_14943,N_13564,N_13733);
xnor U14944 (N_14944,N_13508,N_14176);
nand U14945 (N_14945,N_14017,N_13898);
or U14946 (N_14946,N_14191,N_13706);
nor U14947 (N_14947,N_14132,N_14000);
or U14948 (N_14948,N_13790,N_14196);
and U14949 (N_14949,N_13780,N_13768);
nand U14950 (N_14950,N_14025,N_13580);
and U14951 (N_14951,N_13837,N_14171);
nor U14952 (N_14952,N_13553,N_14202);
and U14953 (N_14953,N_13504,N_13523);
or U14954 (N_14954,N_13525,N_13785);
or U14955 (N_14955,N_13757,N_13832);
and U14956 (N_14956,N_13898,N_14080);
nand U14957 (N_14957,N_13562,N_13669);
xor U14958 (N_14958,N_14150,N_14219);
nand U14959 (N_14959,N_13822,N_13955);
nand U14960 (N_14960,N_14063,N_14219);
nor U14961 (N_14961,N_13664,N_13527);
or U14962 (N_14962,N_13609,N_14154);
and U14963 (N_14963,N_13620,N_14095);
nand U14964 (N_14964,N_13798,N_13891);
nand U14965 (N_14965,N_13994,N_14030);
and U14966 (N_14966,N_13655,N_13922);
nand U14967 (N_14967,N_13818,N_14130);
nand U14968 (N_14968,N_13897,N_13847);
nand U14969 (N_14969,N_13769,N_13989);
nor U14970 (N_14970,N_14210,N_14065);
or U14971 (N_14971,N_13761,N_13932);
nor U14972 (N_14972,N_13719,N_14151);
or U14973 (N_14973,N_14021,N_14217);
nand U14974 (N_14974,N_13859,N_13789);
nor U14975 (N_14975,N_14003,N_13867);
nor U14976 (N_14976,N_13901,N_13739);
nand U14977 (N_14977,N_13822,N_13728);
nor U14978 (N_14978,N_13894,N_13792);
nand U14979 (N_14979,N_14102,N_14017);
or U14980 (N_14980,N_13814,N_13555);
and U14981 (N_14981,N_13854,N_13573);
xor U14982 (N_14982,N_13919,N_14240);
or U14983 (N_14983,N_13605,N_13639);
and U14984 (N_14984,N_14232,N_13545);
nand U14985 (N_14985,N_13741,N_13551);
and U14986 (N_14986,N_13835,N_13542);
or U14987 (N_14987,N_13543,N_13888);
or U14988 (N_14988,N_13958,N_14035);
or U14989 (N_14989,N_14033,N_13830);
nor U14990 (N_14990,N_13829,N_13626);
or U14991 (N_14991,N_13957,N_13793);
xor U14992 (N_14992,N_13591,N_13812);
nor U14993 (N_14993,N_13640,N_14226);
nand U14994 (N_14994,N_13733,N_13568);
nor U14995 (N_14995,N_13518,N_13982);
or U14996 (N_14996,N_13933,N_14217);
or U14997 (N_14997,N_14133,N_14022);
nor U14998 (N_14998,N_13790,N_14240);
and U14999 (N_14999,N_14055,N_13760);
or UO_0 (O_0,N_14965,N_14512);
or UO_1 (O_1,N_14383,N_14281);
or UO_2 (O_2,N_14523,N_14333);
nand UO_3 (O_3,N_14638,N_14838);
and UO_4 (O_4,N_14425,N_14624);
nand UO_5 (O_5,N_14556,N_14568);
and UO_6 (O_6,N_14521,N_14321);
nand UO_7 (O_7,N_14754,N_14348);
or UO_8 (O_8,N_14927,N_14776);
or UO_9 (O_9,N_14596,N_14466);
and UO_10 (O_10,N_14855,N_14361);
nand UO_11 (O_11,N_14816,N_14283);
and UO_12 (O_12,N_14574,N_14690);
and UO_13 (O_13,N_14478,N_14258);
and UO_14 (O_14,N_14431,N_14772);
nand UO_15 (O_15,N_14909,N_14504);
and UO_16 (O_16,N_14465,N_14675);
nor UO_17 (O_17,N_14547,N_14961);
or UO_18 (O_18,N_14765,N_14287);
or UO_19 (O_19,N_14609,N_14403);
and UO_20 (O_20,N_14317,N_14875);
or UO_21 (O_21,N_14810,N_14896);
nand UO_22 (O_22,N_14720,N_14856);
nand UO_23 (O_23,N_14994,N_14678);
or UO_24 (O_24,N_14885,N_14761);
and UO_25 (O_25,N_14549,N_14646);
nor UO_26 (O_26,N_14443,N_14968);
nor UO_27 (O_27,N_14584,N_14301);
xnor UO_28 (O_28,N_14682,N_14368);
or UO_29 (O_29,N_14878,N_14845);
nand UO_30 (O_30,N_14662,N_14589);
nand UO_31 (O_31,N_14435,N_14937);
or UO_32 (O_32,N_14851,N_14311);
nand UO_33 (O_33,N_14340,N_14446);
or UO_34 (O_34,N_14531,N_14917);
and UO_35 (O_35,N_14935,N_14977);
and UO_36 (O_36,N_14710,N_14603);
or UO_37 (O_37,N_14688,N_14873);
or UO_38 (O_38,N_14359,N_14586);
nor UO_39 (O_39,N_14483,N_14803);
nor UO_40 (O_40,N_14421,N_14929);
nand UO_41 (O_41,N_14762,N_14905);
or UO_42 (O_42,N_14413,N_14643);
nand UO_43 (O_43,N_14789,N_14899);
nand UO_44 (O_44,N_14460,N_14999);
and UO_45 (O_45,N_14319,N_14519);
nand UO_46 (O_46,N_14288,N_14402);
nand UO_47 (O_47,N_14978,N_14658);
nor UO_48 (O_48,N_14974,N_14818);
xnor UO_49 (O_49,N_14986,N_14707);
and UO_50 (O_50,N_14684,N_14472);
and UO_51 (O_51,N_14619,N_14698);
and UO_52 (O_52,N_14303,N_14382);
or UO_53 (O_53,N_14718,N_14256);
nand UO_54 (O_54,N_14820,N_14894);
nor UO_55 (O_55,N_14887,N_14979);
or UO_56 (O_56,N_14412,N_14262);
and UO_57 (O_57,N_14835,N_14976);
nor UO_58 (O_58,N_14757,N_14877);
or UO_59 (O_59,N_14396,N_14860);
and UO_60 (O_60,N_14514,N_14441);
and UO_61 (O_61,N_14781,N_14615);
nor UO_62 (O_62,N_14482,N_14993);
and UO_63 (O_63,N_14723,N_14585);
nor UO_64 (O_64,N_14387,N_14279);
and UO_65 (O_65,N_14526,N_14973);
nand UO_66 (O_66,N_14385,N_14278);
nor UO_67 (O_67,N_14839,N_14398);
nand UO_68 (O_68,N_14947,N_14959);
nand UO_69 (O_69,N_14798,N_14381);
nand UO_70 (O_70,N_14534,N_14951);
nor UO_71 (O_71,N_14270,N_14774);
nor UO_72 (O_72,N_14987,N_14492);
xnor UO_73 (O_73,N_14581,N_14632);
and UO_74 (O_74,N_14306,N_14452);
and UO_75 (O_75,N_14957,N_14604);
nand UO_76 (O_76,N_14966,N_14777);
nand UO_77 (O_77,N_14290,N_14712);
nand UO_78 (O_78,N_14980,N_14923);
nand UO_79 (O_79,N_14250,N_14797);
or UO_80 (O_80,N_14486,N_14814);
nor UO_81 (O_81,N_14631,N_14691);
nand UO_82 (O_82,N_14796,N_14499);
nor UO_83 (O_83,N_14367,N_14595);
and UO_84 (O_84,N_14889,N_14373);
and UO_85 (O_85,N_14756,N_14815);
nor UO_86 (O_86,N_14943,N_14576);
and UO_87 (O_87,N_14904,N_14656);
and UO_88 (O_88,N_14520,N_14990);
nor UO_89 (O_89,N_14299,N_14399);
nor UO_90 (O_90,N_14622,N_14846);
nor UO_91 (O_91,N_14956,N_14436);
nand UO_92 (O_92,N_14830,N_14612);
nor UO_93 (O_93,N_14423,N_14374);
nor UO_94 (O_94,N_14865,N_14420);
nand UO_95 (O_95,N_14379,N_14437);
and UO_96 (O_96,N_14580,N_14969);
xnor UO_97 (O_97,N_14392,N_14602);
nor UO_98 (O_98,N_14686,N_14694);
nand UO_99 (O_99,N_14608,N_14536);
or UO_100 (O_100,N_14828,N_14705);
or UO_101 (O_101,N_14992,N_14438);
and UO_102 (O_102,N_14975,N_14424);
or UO_103 (O_103,N_14357,N_14273);
and UO_104 (O_104,N_14310,N_14912);
or UO_105 (O_105,N_14958,N_14529);
nor UO_106 (O_106,N_14625,N_14759);
or UO_107 (O_107,N_14463,N_14430);
xor UO_108 (O_108,N_14857,N_14775);
xnor UO_109 (O_109,N_14308,N_14663);
and UO_110 (O_110,N_14351,N_14849);
nand UO_111 (O_111,N_14895,N_14884);
xnor UO_112 (O_112,N_14579,N_14479);
and UO_113 (O_113,N_14285,N_14605);
nand UO_114 (O_114,N_14664,N_14711);
and UO_115 (O_115,N_14347,N_14791);
and UO_116 (O_116,N_14352,N_14511);
nand UO_117 (O_117,N_14545,N_14669);
nand UO_118 (O_118,N_14747,N_14474);
nor UO_119 (O_119,N_14405,N_14764);
nand UO_120 (O_120,N_14569,N_14782);
and UO_121 (O_121,N_14869,N_14284);
nand UO_122 (O_122,N_14610,N_14661);
or UO_123 (O_123,N_14907,N_14445);
nand UO_124 (O_124,N_14832,N_14613);
xor UO_125 (O_125,N_14388,N_14307);
nor UO_126 (O_126,N_14433,N_14942);
xnor UO_127 (O_127,N_14670,N_14427);
xor UO_128 (O_128,N_14449,N_14516);
nor UO_129 (O_129,N_14847,N_14416);
nor UO_130 (O_130,N_14503,N_14349);
or UO_131 (O_131,N_14377,N_14600);
nand UO_132 (O_132,N_14844,N_14725);
nor UO_133 (O_133,N_14254,N_14471);
nor UO_134 (O_134,N_14537,N_14888);
and UO_135 (O_135,N_14751,N_14484);
nor UO_136 (O_136,N_14734,N_14949);
nor UO_137 (O_137,N_14954,N_14882);
and UO_138 (O_138,N_14840,N_14312);
nor UO_139 (O_139,N_14378,N_14591);
or UO_140 (O_140,N_14409,N_14850);
or UO_141 (O_141,N_14724,N_14448);
nor UO_142 (O_142,N_14414,N_14593);
or UO_143 (O_143,N_14962,N_14567);
or UO_144 (O_144,N_14495,N_14459);
nor UO_145 (O_145,N_14518,N_14527);
or UO_146 (O_146,N_14517,N_14298);
and UO_147 (O_147,N_14890,N_14647);
nor UO_148 (O_148,N_14326,N_14967);
and UO_149 (O_149,N_14716,N_14627);
nor UO_150 (O_150,N_14834,N_14852);
nor UO_151 (O_151,N_14771,N_14618);
nor UO_152 (O_152,N_14565,N_14826);
nor UO_153 (O_153,N_14410,N_14316);
or UO_154 (O_154,N_14350,N_14274);
or UO_155 (O_155,N_14322,N_14490);
nor UO_156 (O_156,N_14548,N_14265);
xor UO_157 (O_157,N_14336,N_14900);
nand UO_158 (O_158,N_14323,N_14864);
nand UO_159 (O_159,N_14394,N_14566);
and UO_160 (O_160,N_14741,N_14970);
or UO_161 (O_161,N_14522,N_14500);
xor UO_162 (O_162,N_14535,N_14344);
or UO_163 (O_163,N_14542,N_14269);
nor UO_164 (O_164,N_14442,N_14685);
and UO_165 (O_165,N_14641,N_14654);
nor UO_166 (O_166,N_14916,N_14315);
and UO_167 (O_167,N_14380,N_14588);
xor UO_168 (O_168,N_14788,N_14964);
nand UO_169 (O_169,N_14300,N_14778);
xnor UO_170 (O_170,N_14811,N_14473);
nand UO_171 (O_171,N_14628,N_14910);
nor UO_172 (O_172,N_14498,N_14680);
xor UO_173 (O_173,N_14808,N_14740);
nor UO_174 (O_174,N_14697,N_14925);
nand UO_175 (O_175,N_14502,N_14933);
and UO_176 (O_176,N_14749,N_14924);
and UO_177 (O_177,N_14945,N_14760);
nand UO_178 (O_178,N_14823,N_14389);
or UO_179 (O_179,N_14739,N_14748);
or UO_180 (O_180,N_14833,N_14713);
or UO_181 (O_181,N_14842,N_14914);
or UO_182 (O_182,N_14881,N_14475);
or UO_183 (O_183,N_14543,N_14932);
or UO_184 (O_184,N_14614,N_14305);
nor UO_185 (O_185,N_14984,N_14462);
and UO_186 (O_186,N_14393,N_14329);
and UO_187 (O_187,N_14458,N_14454);
nand UO_188 (O_188,N_14767,N_14773);
or UO_189 (O_189,N_14677,N_14444);
and UO_190 (O_190,N_14981,N_14507);
and UO_191 (O_191,N_14708,N_14768);
nor UO_192 (O_192,N_14268,N_14800);
nor UO_193 (O_193,N_14271,N_14544);
nand UO_194 (O_194,N_14313,N_14331);
nand UO_195 (O_195,N_14611,N_14450);
and UO_196 (O_196,N_14440,N_14871);
and UO_197 (O_197,N_14577,N_14750);
nor UO_198 (O_198,N_14702,N_14779);
xor UO_199 (O_199,N_14257,N_14730);
or UO_200 (O_200,N_14867,N_14919);
and UO_201 (O_201,N_14792,N_14858);
nand UO_202 (O_202,N_14699,N_14780);
or UO_203 (O_203,N_14571,N_14728);
nor UO_204 (O_204,N_14562,N_14453);
or UO_205 (O_205,N_14296,N_14709);
or UO_206 (O_206,N_14309,N_14515);
nand UO_207 (O_207,N_14971,N_14607);
and UO_208 (O_208,N_14883,N_14477);
and UO_209 (O_209,N_14679,N_14696);
nor UO_210 (O_210,N_14636,N_14601);
nand UO_211 (O_211,N_14572,N_14346);
and UO_212 (O_212,N_14341,N_14868);
and UO_213 (O_213,N_14369,N_14418);
nand UO_214 (O_214,N_14785,N_14489);
nand UO_215 (O_215,N_14415,N_14955);
nor UO_216 (O_216,N_14623,N_14872);
nand UO_217 (O_217,N_14982,N_14652);
and UO_218 (O_218,N_14640,N_14746);
or UO_219 (O_219,N_14722,N_14294);
or UO_220 (O_220,N_14695,N_14330);
nand UO_221 (O_221,N_14599,N_14906);
nand UO_222 (O_222,N_14375,N_14597);
or UO_223 (O_223,N_14338,N_14802);
or UO_224 (O_224,N_14752,N_14451);
xor UO_225 (O_225,N_14805,N_14952);
nand UO_226 (O_226,N_14386,N_14880);
and UO_227 (O_227,N_14715,N_14561);
and UO_228 (O_228,N_14550,N_14292);
or UO_229 (O_229,N_14532,N_14295);
nand UO_230 (O_230,N_14736,N_14496);
nor UO_231 (O_231,N_14264,N_14456);
or UO_232 (O_232,N_14991,N_14863);
and UO_233 (O_233,N_14738,N_14540);
xnor UO_234 (O_234,N_14841,N_14946);
nand UO_235 (O_235,N_14660,N_14583);
or UO_236 (O_236,N_14464,N_14795);
and UO_237 (O_237,N_14509,N_14719);
and UO_238 (O_238,N_14721,N_14275);
nor UO_239 (O_239,N_14928,N_14985);
and UO_240 (O_240,N_14617,N_14480);
or UO_241 (O_241,N_14806,N_14582);
nor UO_242 (O_242,N_14704,N_14908);
and UO_243 (O_243,N_14650,N_14541);
and UO_244 (O_244,N_14493,N_14575);
nor UO_245 (O_245,N_14457,N_14862);
xnor UO_246 (O_246,N_14960,N_14570);
or UO_247 (O_247,N_14941,N_14485);
nand UO_248 (O_248,N_14476,N_14513);
nand UO_249 (O_249,N_14280,N_14731);
nor UO_250 (O_250,N_14758,N_14786);
nor UO_251 (O_251,N_14983,N_14700);
nand UO_252 (O_252,N_14252,N_14481);
and UO_253 (O_253,N_14911,N_14809);
nor UO_254 (O_254,N_14384,N_14876);
nand UO_255 (O_255,N_14784,N_14787);
or UO_256 (O_256,N_14859,N_14689);
nor UO_257 (O_257,N_14897,N_14870);
nor UO_258 (O_258,N_14732,N_14996);
nor UO_259 (O_259,N_14419,N_14655);
or UO_260 (O_260,N_14372,N_14701);
or UO_261 (O_261,N_14854,N_14345);
nor UO_262 (O_262,N_14320,N_14649);
and UO_263 (O_263,N_14318,N_14726);
nor UO_264 (O_264,N_14745,N_14263);
nor UO_265 (O_265,N_14505,N_14633);
nor UO_266 (O_266,N_14592,N_14468);
or UO_267 (O_267,N_14717,N_14848);
or UO_268 (O_268,N_14439,N_14621);
and UO_269 (O_269,N_14934,N_14594);
nand UO_270 (O_270,N_14342,N_14671);
xor UO_271 (O_271,N_14343,N_14672);
nor UO_272 (O_272,N_14668,N_14902);
or UO_273 (O_273,N_14528,N_14755);
or UO_274 (O_274,N_14259,N_14302);
and UO_275 (O_275,N_14674,N_14395);
and UO_276 (O_276,N_14354,N_14735);
or UO_277 (O_277,N_14559,N_14822);
xor UO_278 (O_278,N_14948,N_14769);
nand UO_279 (O_279,N_14590,N_14365);
nor UO_280 (O_280,N_14467,N_14939);
nor UO_281 (O_281,N_14920,N_14819);
or UO_282 (O_282,N_14866,N_14564);
nor UO_283 (O_283,N_14358,N_14276);
xnor UO_284 (O_284,N_14598,N_14525);
and UO_285 (O_285,N_14277,N_14657);
nor UO_286 (O_286,N_14936,N_14325);
nor UO_287 (O_287,N_14553,N_14429);
or UO_288 (O_288,N_14799,N_14417);
nor UO_289 (O_289,N_14687,N_14998);
nor UO_290 (O_290,N_14364,N_14557);
nand UO_291 (O_291,N_14391,N_14953);
nand UO_292 (O_292,N_14606,N_14339);
nor UO_293 (O_293,N_14497,N_14703);
or UO_294 (O_294,N_14667,N_14644);
nand UO_295 (O_295,N_14332,N_14737);
and UO_296 (O_296,N_14578,N_14560);
or UO_297 (O_297,N_14404,N_14407);
and UO_298 (O_298,N_14861,N_14659);
nor UO_299 (O_299,N_14673,N_14573);
or UO_300 (O_300,N_14744,N_14563);
nand UO_301 (O_301,N_14807,N_14930);
and UO_302 (O_302,N_14639,N_14524);
and UO_303 (O_303,N_14693,N_14901);
nand UO_304 (O_304,N_14824,N_14918);
nand UO_305 (O_305,N_14530,N_14397);
nand UO_306 (O_306,N_14253,N_14813);
and UO_307 (O_307,N_14829,N_14558);
nand UO_308 (O_308,N_14626,N_14794);
xor UO_309 (O_309,N_14821,N_14455);
nand UO_310 (O_310,N_14616,N_14266);
and UO_311 (O_311,N_14790,N_14629);
nand UO_312 (O_312,N_14408,N_14293);
nor UO_313 (O_313,N_14825,N_14853);
or UO_314 (O_314,N_14676,N_14360);
and UO_315 (O_315,N_14488,N_14763);
nand UO_316 (O_316,N_14469,N_14337);
or UO_317 (O_317,N_14620,N_14411);
xor UO_318 (O_318,N_14366,N_14804);
or UO_319 (O_319,N_14304,N_14371);
or UO_320 (O_320,N_14554,N_14328);
nor UO_321 (O_321,N_14434,N_14487);
nor UO_322 (O_322,N_14827,N_14913);
nor UO_323 (O_323,N_14508,N_14362);
nor UO_324 (O_324,N_14692,N_14637);
nand UO_325 (O_325,N_14743,N_14255);
nand UO_326 (O_326,N_14491,N_14727);
nand UO_327 (O_327,N_14989,N_14766);
xnor UO_328 (O_328,N_14931,N_14356);
nand UO_329 (O_329,N_14260,N_14944);
or UO_330 (O_330,N_14447,N_14921);
and UO_331 (O_331,N_14915,N_14893);
and UO_332 (O_332,N_14665,N_14400);
nor UO_333 (O_333,N_14645,N_14297);
nor UO_334 (O_334,N_14376,N_14272);
nand UO_335 (O_335,N_14950,N_14494);
and UO_336 (O_336,N_14426,N_14363);
nand UO_337 (O_337,N_14886,N_14432);
and UO_338 (O_338,N_14891,N_14286);
and UO_339 (O_339,N_14422,N_14635);
nand UO_340 (O_340,N_14506,N_14706);
nand UO_341 (O_341,N_14898,N_14630);
nor UO_342 (O_342,N_14314,N_14267);
or UO_343 (O_343,N_14335,N_14892);
or UO_344 (O_344,N_14753,N_14995);
nor UO_345 (O_345,N_14831,N_14651);
and UO_346 (O_346,N_14903,N_14963);
or UO_347 (O_347,N_14533,N_14666);
xnor UO_348 (O_348,N_14538,N_14282);
or UO_349 (O_349,N_14683,N_14836);
and UO_350 (O_350,N_14642,N_14370);
nor UO_351 (O_351,N_14291,N_14355);
nand UO_352 (O_352,N_14261,N_14801);
nand UO_353 (O_353,N_14926,N_14988);
and UO_354 (O_354,N_14470,N_14539);
and UO_355 (O_355,N_14587,N_14461);
and UO_356 (O_356,N_14551,N_14812);
xnor UO_357 (O_357,N_14648,N_14555);
or UO_358 (O_358,N_14653,N_14634);
nand UO_359 (O_359,N_14334,N_14289);
nor UO_360 (O_360,N_14552,N_14327);
nand UO_361 (O_361,N_14251,N_14353);
or UO_362 (O_362,N_14770,N_14793);
nor UO_363 (O_363,N_14837,N_14874);
or UO_364 (O_364,N_14783,N_14733);
nand UO_365 (O_365,N_14406,N_14817);
nand UO_366 (O_366,N_14938,N_14972);
nand UO_367 (O_367,N_14390,N_14501);
nand UO_368 (O_368,N_14324,N_14997);
or UO_369 (O_369,N_14681,N_14843);
or UO_370 (O_370,N_14729,N_14940);
or UO_371 (O_371,N_14401,N_14742);
xnor UO_372 (O_372,N_14510,N_14879);
nor UO_373 (O_373,N_14428,N_14714);
nor UO_374 (O_374,N_14922,N_14546);
or UO_375 (O_375,N_14828,N_14358);
and UO_376 (O_376,N_14682,N_14471);
nor UO_377 (O_377,N_14464,N_14857);
nor UO_378 (O_378,N_14859,N_14760);
and UO_379 (O_379,N_14939,N_14769);
and UO_380 (O_380,N_14929,N_14325);
or UO_381 (O_381,N_14314,N_14768);
nand UO_382 (O_382,N_14557,N_14900);
and UO_383 (O_383,N_14750,N_14454);
and UO_384 (O_384,N_14535,N_14363);
or UO_385 (O_385,N_14747,N_14425);
and UO_386 (O_386,N_14481,N_14364);
xnor UO_387 (O_387,N_14671,N_14370);
and UO_388 (O_388,N_14958,N_14685);
nor UO_389 (O_389,N_14924,N_14269);
nor UO_390 (O_390,N_14681,N_14639);
or UO_391 (O_391,N_14805,N_14746);
or UO_392 (O_392,N_14745,N_14723);
nand UO_393 (O_393,N_14362,N_14308);
or UO_394 (O_394,N_14486,N_14629);
or UO_395 (O_395,N_14831,N_14273);
or UO_396 (O_396,N_14629,N_14989);
nor UO_397 (O_397,N_14669,N_14356);
or UO_398 (O_398,N_14807,N_14269);
nand UO_399 (O_399,N_14769,N_14431);
or UO_400 (O_400,N_14304,N_14252);
nor UO_401 (O_401,N_14842,N_14853);
nand UO_402 (O_402,N_14799,N_14562);
nand UO_403 (O_403,N_14885,N_14434);
nor UO_404 (O_404,N_14338,N_14741);
nor UO_405 (O_405,N_14613,N_14331);
and UO_406 (O_406,N_14865,N_14527);
nor UO_407 (O_407,N_14442,N_14875);
and UO_408 (O_408,N_14391,N_14261);
or UO_409 (O_409,N_14830,N_14273);
or UO_410 (O_410,N_14940,N_14316);
and UO_411 (O_411,N_14353,N_14647);
and UO_412 (O_412,N_14893,N_14870);
nand UO_413 (O_413,N_14961,N_14633);
or UO_414 (O_414,N_14330,N_14285);
nor UO_415 (O_415,N_14268,N_14275);
or UO_416 (O_416,N_14830,N_14341);
nand UO_417 (O_417,N_14890,N_14570);
nor UO_418 (O_418,N_14495,N_14254);
nand UO_419 (O_419,N_14875,N_14555);
nand UO_420 (O_420,N_14698,N_14821);
nor UO_421 (O_421,N_14318,N_14580);
or UO_422 (O_422,N_14505,N_14711);
and UO_423 (O_423,N_14998,N_14594);
and UO_424 (O_424,N_14481,N_14569);
nand UO_425 (O_425,N_14633,N_14503);
or UO_426 (O_426,N_14965,N_14880);
and UO_427 (O_427,N_14911,N_14280);
or UO_428 (O_428,N_14668,N_14489);
or UO_429 (O_429,N_14682,N_14342);
nand UO_430 (O_430,N_14521,N_14707);
or UO_431 (O_431,N_14830,N_14337);
and UO_432 (O_432,N_14549,N_14649);
or UO_433 (O_433,N_14797,N_14742);
and UO_434 (O_434,N_14281,N_14595);
nor UO_435 (O_435,N_14676,N_14875);
nor UO_436 (O_436,N_14713,N_14941);
nand UO_437 (O_437,N_14741,N_14909);
or UO_438 (O_438,N_14613,N_14265);
nor UO_439 (O_439,N_14962,N_14587);
or UO_440 (O_440,N_14379,N_14959);
and UO_441 (O_441,N_14336,N_14741);
or UO_442 (O_442,N_14696,N_14467);
xor UO_443 (O_443,N_14853,N_14973);
or UO_444 (O_444,N_14666,N_14992);
or UO_445 (O_445,N_14628,N_14484);
and UO_446 (O_446,N_14674,N_14726);
nor UO_447 (O_447,N_14386,N_14653);
or UO_448 (O_448,N_14747,N_14972);
and UO_449 (O_449,N_14267,N_14466);
nor UO_450 (O_450,N_14774,N_14284);
nor UO_451 (O_451,N_14944,N_14419);
or UO_452 (O_452,N_14720,N_14790);
xor UO_453 (O_453,N_14464,N_14834);
nor UO_454 (O_454,N_14894,N_14696);
or UO_455 (O_455,N_14332,N_14738);
or UO_456 (O_456,N_14947,N_14933);
xor UO_457 (O_457,N_14954,N_14466);
and UO_458 (O_458,N_14647,N_14598);
and UO_459 (O_459,N_14297,N_14509);
nand UO_460 (O_460,N_14902,N_14949);
nand UO_461 (O_461,N_14386,N_14748);
and UO_462 (O_462,N_14854,N_14861);
or UO_463 (O_463,N_14342,N_14452);
or UO_464 (O_464,N_14890,N_14879);
and UO_465 (O_465,N_14746,N_14914);
or UO_466 (O_466,N_14833,N_14295);
nor UO_467 (O_467,N_14516,N_14734);
or UO_468 (O_468,N_14351,N_14324);
xor UO_469 (O_469,N_14988,N_14623);
and UO_470 (O_470,N_14466,N_14826);
and UO_471 (O_471,N_14597,N_14948);
or UO_472 (O_472,N_14583,N_14516);
xnor UO_473 (O_473,N_14463,N_14281);
xnor UO_474 (O_474,N_14832,N_14511);
or UO_475 (O_475,N_14620,N_14612);
nor UO_476 (O_476,N_14818,N_14376);
and UO_477 (O_477,N_14477,N_14772);
xnor UO_478 (O_478,N_14527,N_14255);
nand UO_479 (O_479,N_14573,N_14785);
nor UO_480 (O_480,N_14791,N_14526);
and UO_481 (O_481,N_14257,N_14584);
nand UO_482 (O_482,N_14576,N_14410);
and UO_483 (O_483,N_14492,N_14709);
or UO_484 (O_484,N_14573,N_14814);
nand UO_485 (O_485,N_14694,N_14567);
and UO_486 (O_486,N_14543,N_14394);
nand UO_487 (O_487,N_14562,N_14538);
nor UO_488 (O_488,N_14769,N_14552);
nand UO_489 (O_489,N_14510,N_14507);
nand UO_490 (O_490,N_14963,N_14547);
and UO_491 (O_491,N_14886,N_14412);
or UO_492 (O_492,N_14851,N_14513);
xnor UO_493 (O_493,N_14385,N_14378);
nor UO_494 (O_494,N_14988,N_14556);
nor UO_495 (O_495,N_14846,N_14859);
xnor UO_496 (O_496,N_14938,N_14789);
nor UO_497 (O_497,N_14628,N_14952);
and UO_498 (O_498,N_14756,N_14821);
and UO_499 (O_499,N_14988,N_14950);
xnor UO_500 (O_500,N_14929,N_14276);
nand UO_501 (O_501,N_14743,N_14990);
xor UO_502 (O_502,N_14461,N_14278);
or UO_503 (O_503,N_14420,N_14862);
or UO_504 (O_504,N_14918,N_14258);
nor UO_505 (O_505,N_14869,N_14752);
nand UO_506 (O_506,N_14779,N_14740);
or UO_507 (O_507,N_14939,N_14290);
and UO_508 (O_508,N_14957,N_14806);
nand UO_509 (O_509,N_14448,N_14364);
and UO_510 (O_510,N_14831,N_14544);
nor UO_511 (O_511,N_14604,N_14450);
or UO_512 (O_512,N_14429,N_14715);
and UO_513 (O_513,N_14415,N_14819);
nor UO_514 (O_514,N_14463,N_14969);
and UO_515 (O_515,N_14856,N_14611);
nand UO_516 (O_516,N_14276,N_14489);
nand UO_517 (O_517,N_14329,N_14411);
and UO_518 (O_518,N_14601,N_14347);
nand UO_519 (O_519,N_14308,N_14578);
nor UO_520 (O_520,N_14314,N_14576);
or UO_521 (O_521,N_14719,N_14783);
nand UO_522 (O_522,N_14633,N_14906);
or UO_523 (O_523,N_14985,N_14453);
nand UO_524 (O_524,N_14551,N_14877);
and UO_525 (O_525,N_14627,N_14372);
nor UO_526 (O_526,N_14339,N_14503);
or UO_527 (O_527,N_14415,N_14312);
nor UO_528 (O_528,N_14737,N_14585);
nor UO_529 (O_529,N_14632,N_14983);
nor UO_530 (O_530,N_14818,N_14989);
nor UO_531 (O_531,N_14605,N_14448);
or UO_532 (O_532,N_14320,N_14307);
and UO_533 (O_533,N_14546,N_14748);
xor UO_534 (O_534,N_14904,N_14580);
xnor UO_535 (O_535,N_14927,N_14729);
xnor UO_536 (O_536,N_14450,N_14304);
and UO_537 (O_537,N_14254,N_14620);
nand UO_538 (O_538,N_14681,N_14418);
or UO_539 (O_539,N_14393,N_14377);
and UO_540 (O_540,N_14683,N_14454);
and UO_541 (O_541,N_14827,N_14569);
nor UO_542 (O_542,N_14440,N_14581);
nor UO_543 (O_543,N_14759,N_14360);
nand UO_544 (O_544,N_14714,N_14884);
and UO_545 (O_545,N_14777,N_14773);
nand UO_546 (O_546,N_14724,N_14906);
nand UO_547 (O_547,N_14934,N_14640);
nand UO_548 (O_548,N_14772,N_14820);
and UO_549 (O_549,N_14768,N_14645);
nor UO_550 (O_550,N_14838,N_14306);
nand UO_551 (O_551,N_14828,N_14438);
xor UO_552 (O_552,N_14271,N_14711);
and UO_553 (O_553,N_14262,N_14858);
nor UO_554 (O_554,N_14906,N_14563);
nor UO_555 (O_555,N_14936,N_14741);
or UO_556 (O_556,N_14995,N_14569);
nor UO_557 (O_557,N_14621,N_14481);
nand UO_558 (O_558,N_14362,N_14300);
xnor UO_559 (O_559,N_14852,N_14813);
nor UO_560 (O_560,N_14812,N_14600);
or UO_561 (O_561,N_14326,N_14451);
nor UO_562 (O_562,N_14725,N_14676);
nor UO_563 (O_563,N_14557,N_14471);
nand UO_564 (O_564,N_14446,N_14311);
nand UO_565 (O_565,N_14695,N_14420);
and UO_566 (O_566,N_14500,N_14519);
and UO_567 (O_567,N_14659,N_14269);
xnor UO_568 (O_568,N_14471,N_14407);
nand UO_569 (O_569,N_14730,N_14389);
nor UO_570 (O_570,N_14744,N_14416);
nand UO_571 (O_571,N_14631,N_14665);
nor UO_572 (O_572,N_14920,N_14270);
nand UO_573 (O_573,N_14548,N_14409);
or UO_574 (O_574,N_14993,N_14968);
xor UO_575 (O_575,N_14831,N_14481);
xnor UO_576 (O_576,N_14402,N_14481);
and UO_577 (O_577,N_14767,N_14487);
and UO_578 (O_578,N_14724,N_14774);
nor UO_579 (O_579,N_14646,N_14538);
xor UO_580 (O_580,N_14704,N_14801);
nand UO_581 (O_581,N_14833,N_14732);
or UO_582 (O_582,N_14336,N_14277);
nand UO_583 (O_583,N_14402,N_14669);
nor UO_584 (O_584,N_14859,N_14630);
or UO_585 (O_585,N_14550,N_14342);
nand UO_586 (O_586,N_14292,N_14660);
xor UO_587 (O_587,N_14363,N_14772);
nor UO_588 (O_588,N_14825,N_14565);
nand UO_589 (O_589,N_14521,N_14931);
or UO_590 (O_590,N_14912,N_14295);
nand UO_591 (O_591,N_14348,N_14599);
or UO_592 (O_592,N_14632,N_14481);
nand UO_593 (O_593,N_14617,N_14775);
or UO_594 (O_594,N_14988,N_14329);
and UO_595 (O_595,N_14314,N_14377);
nand UO_596 (O_596,N_14384,N_14267);
or UO_597 (O_597,N_14450,N_14815);
nor UO_598 (O_598,N_14893,N_14440);
xor UO_599 (O_599,N_14858,N_14546);
nand UO_600 (O_600,N_14260,N_14557);
nor UO_601 (O_601,N_14388,N_14251);
xnor UO_602 (O_602,N_14467,N_14485);
and UO_603 (O_603,N_14529,N_14940);
or UO_604 (O_604,N_14728,N_14403);
nor UO_605 (O_605,N_14407,N_14418);
nand UO_606 (O_606,N_14728,N_14692);
nor UO_607 (O_607,N_14253,N_14472);
nor UO_608 (O_608,N_14552,N_14314);
or UO_609 (O_609,N_14552,N_14595);
nor UO_610 (O_610,N_14252,N_14968);
and UO_611 (O_611,N_14597,N_14739);
xor UO_612 (O_612,N_14765,N_14545);
xnor UO_613 (O_613,N_14518,N_14277);
nand UO_614 (O_614,N_14453,N_14285);
or UO_615 (O_615,N_14623,N_14877);
nor UO_616 (O_616,N_14643,N_14943);
nor UO_617 (O_617,N_14482,N_14575);
nand UO_618 (O_618,N_14403,N_14288);
or UO_619 (O_619,N_14477,N_14389);
nor UO_620 (O_620,N_14877,N_14693);
or UO_621 (O_621,N_14891,N_14587);
and UO_622 (O_622,N_14589,N_14740);
xnor UO_623 (O_623,N_14633,N_14306);
and UO_624 (O_624,N_14313,N_14281);
and UO_625 (O_625,N_14906,N_14465);
and UO_626 (O_626,N_14254,N_14447);
and UO_627 (O_627,N_14870,N_14482);
and UO_628 (O_628,N_14367,N_14864);
nand UO_629 (O_629,N_14528,N_14598);
nand UO_630 (O_630,N_14784,N_14275);
and UO_631 (O_631,N_14397,N_14661);
or UO_632 (O_632,N_14800,N_14990);
and UO_633 (O_633,N_14691,N_14475);
nand UO_634 (O_634,N_14276,N_14899);
nand UO_635 (O_635,N_14545,N_14552);
nor UO_636 (O_636,N_14953,N_14923);
nor UO_637 (O_637,N_14688,N_14466);
nand UO_638 (O_638,N_14826,N_14996);
xor UO_639 (O_639,N_14476,N_14362);
nor UO_640 (O_640,N_14763,N_14739);
nor UO_641 (O_641,N_14567,N_14460);
nand UO_642 (O_642,N_14569,N_14580);
nor UO_643 (O_643,N_14727,N_14825);
or UO_644 (O_644,N_14621,N_14548);
or UO_645 (O_645,N_14468,N_14445);
and UO_646 (O_646,N_14294,N_14298);
or UO_647 (O_647,N_14265,N_14361);
or UO_648 (O_648,N_14484,N_14633);
nor UO_649 (O_649,N_14334,N_14284);
xor UO_650 (O_650,N_14925,N_14762);
and UO_651 (O_651,N_14940,N_14291);
and UO_652 (O_652,N_14491,N_14396);
nor UO_653 (O_653,N_14424,N_14547);
and UO_654 (O_654,N_14758,N_14903);
nor UO_655 (O_655,N_14316,N_14504);
xnor UO_656 (O_656,N_14846,N_14474);
or UO_657 (O_657,N_14732,N_14504);
and UO_658 (O_658,N_14740,N_14933);
nor UO_659 (O_659,N_14894,N_14997);
nand UO_660 (O_660,N_14904,N_14360);
and UO_661 (O_661,N_14474,N_14599);
nor UO_662 (O_662,N_14585,N_14943);
nor UO_663 (O_663,N_14253,N_14802);
or UO_664 (O_664,N_14894,N_14517);
or UO_665 (O_665,N_14412,N_14332);
nor UO_666 (O_666,N_14873,N_14893);
or UO_667 (O_667,N_14803,N_14513);
nand UO_668 (O_668,N_14430,N_14487);
nor UO_669 (O_669,N_14670,N_14517);
nand UO_670 (O_670,N_14323,N_14713);
and UO_671 (O_671,N_14955,N_14346);
nand UO_672 (O_672,N_14351,N_14965);
nand UO_673 (O_673,N_14965,N_14688);
nor UO_674 (O_674,N_14271,N_14744);
nor UO_675 (O_675,N_14979,N_14644);
nor UO_676 (O_676,N_14546,N_14463);
and UO_677 (O_677,N_14708,N_14252);
xor UO_678 (O_678,N_14263,N_14551);
or UO_679 (O_679,N_14991,N_14399);
nand UO_680 (O_680,N_14804,N_14559);
or UO_681 (O_681,N_14981,N_14436);
nor UO_682 (O_682,N_14456,N_14578);
nand UO_683 (O_683,N_14826,N_14654);
and UO_684 (O_684,N_14420,N_14834);
or UO_685 (O_685,N_14493,N_14984);
nand UO_686 (O_686,N_14541,N_14866);
nand UO_687 (O_687,N_14865,N_14781);
xnor UO_688 (O_688,N_14385,N_14579);
or UO_689 (O_689,N_14647,N_14571);
xor UO_690 (O_690,N_14696,N_14562);
nor UO_691 (O_691,N_14656,N_14685);
nor UO_692 (O_692,N_14582,N_14532);
nand UO_693 (O_693,N_14844,N_14777);
and UO_694 (O_694,N_14956,N_14796);
or UO_695 (O_695,N_14578,N_14790);
and UO_696 (O_696,N_14869,N_14544);
and UO_697 (O_697,N_14324,N_14361);
or UO_698 (O_698,N_14415,N_14965);
nand UO_699 (O_699,N_14406,N_14417);
nand UO_700 (O_700,N_14604,N_14404);
or UO_701 (O_701,N_14362,N_14622);
and UO_702 (O_702,N_14704,N_14920);
nor UO_703 (O_703,N_14927,N_14644);
or UO_704 (O_704,N_14554,N_14747);
and UO_705 (O_705,N_14564,N_14602);
nor UO_706 (O_706,N_14583,N_14548);
and UO_707 (O_707,N_14622,N_14524);
nor UO_708 (O_708,N_14688,N_14942);
or UO_709 (O_709,N_14592,N_14825);
xor UO_710 (O_710,N_14674,N_14634);
and UO_711 (O_711,N_14577,N_14841);
and UO_712 (O_712,N_14579,N_14880);
nor UO_713 (O_713,N_14760,N_14426);
nand UO_714 (O_714,N_14882,N_14944);
and UO_715 (O_715,N_14519,N_14376);
nand UO_716 (O_716,N_14579,N_14447);
nand UO_717 (O_717,N_14783,N_14964);
or UO_718 (O_718,N_14537,N_14912);
nand UO_719 (O_719,N_14729,N_14871);
nand UO_720 (O_720,N_14671,N_14350);
nand UO_721 (O_721,N_14496,N_14254);
nand UO_722 (O_722,N_14303,N_14878);
and UO_723 (O_723,N_14250,N_14299);
and UO_724 (O_724,N_14342,N_14969);
xnor UO_725 (O_725,N_14700,N_14978);
nand UO_726 (O_726,N_14673,N_14526);
xnor UO_727 (O_727,N_14785,N_14507);
nand UO_728 (O_728,N_14393,N_14655);
and UO_729 (O_729,N_14396,N_14536);
nor UO_730 (O_730,N_14806,N_14924);
nor UO_731 (O_731,N_14849,N_14292);
xor UO_732 (O_732,N_14266,N_14372);
xnor UO_733 (O_733,N_14682,N_14525);
or UO_734 (O_734,N_14714,N_14754);
nor UO_735 (O_735,N_14345,N_14344);
nand UO_736 (O_736,N_14506,N_14968);
and UO_737 (O_737,N_14897,N_14808);
and UO_738 (O_738,N_14877,N_14264);
and UO_739 (O_739,N_14825,N_14733);
or UO_740 (O_740,N_14317,N_14872);
or UO_741 (O_741,N_14409,N_14931);
or UO_742 (O_742,N_14250,N_14807);
or UO_743 (O_743,N_14307,N_14918);
or UO_744 (O_744,N_14524,N_14385);
nor UO_745 (O_745,N_14425,N_14864);
nand UO_746 (O_746,N_14784,N_14839);
xor UO_747 (O_747,N_14477,N_14680);
or UO_748 (O_748,N_14274,N_14565);
nand UO_749 (O_749,N_14858,N_14692);
or UO_750 (O_750,N_14644,N_14841);
nor UO_751 (O_751,N_14907,N_14376);
nor UO_752 (O_752,N_14496,N_14871);
nand UO_753 (O_753,N_14542,N_14845);
and UO_754 (O_754,N_14774,N_14816);
nand UO_755 (O_755,N_14368,N_14696);
and UO_756 (O_756,N_14617,N_14945);
nor UO_757 (O_757,N_14805,N_14598);
nand UO_758 (O_758,N_14658,N_14830);
nand UO_759 (O_759,N_14661,N_14574);
or UO_760 (O_760,N_14581,N_14544);
nor UO_761 (O_761,N_14513,N_14562);
and UO_762 (O_762,N_14539,N_14945);
or UO_763 (O_763,N_14330,N_14511);
nand UO_764 (O_764,N_14711,N_14577);
or UO_765 (O_765,N_14444,N_14620);
and UO_766 (O_766,N_14947,N_14580);
nand UO_767 (O_767,N_14440,N_14696);
nor UO_768 (O_768,N_14714,N_14991);
or UO_769 (O_769,N_14310,N_14676);
nor UO_770 (O_770,N_14655,N_14479);
nor UO_771 (O_771,N_14614,N_14431);
and UO_772 (O_772,N_14329,N_14614);
or UO_773 (O_773,N_14821,N_14806);
or UO_774 (O_774,N_14651,N_14877);
nand UO_775 (O_775,N_14874,N_14531);
nand UO_776 (O_776,N_14348,N_14597);
nand UO_777 (O_777,N_14712,N_14767);
nand UO_778 (O_778,N_14751,N_14416);
and UO_779 (O_779,N_14974,N_14258);
or UO_780 (O_780,N_14483,N_14771);
nand UO_781 (O_781,N_14495,N_14838);
or UO_782 (O_782,N_14974,N_14365);
or UO_783 (O_783,N_14391,N_14515);
nor UO_784 (O_784,N_14494,N_14980);
and UO_785 (O_785,N_14812,N_14336);
xnor UO_786 (O_786,N_14341,N_14592);
nor UO_787 (O_787,N_14795,N_14787);
and UO_788 (O_788,N_14626,N_14253);
and UO_789 (O_789,N_14330,N_14560);
xnor UO_790 (O_790,N_14876,N_14634);
or UO_791 (O_791,N_14450,N_14429);
or UO_792 (O_792,N_14646,N_14749);
or UO_793 (O_793,N_14320,N_14976);
xor UO_794 (O_794,N_14826,N_14371);
and UO_795 (O_795,N_14985,N_14872);
nand UO_796 (O_796,N_14293,N_14768);
nand UO_797 (O_797,N_14357,N_14738);
nand UO_798 (O_798,N_14951,N_14609);
xnor UO_799 (O_799,N_14707,N_14753);
or UO_800 (O_800,N_14459,N_14824);
nor UO_801 (O_801,N_14360,N_14603);
nor UO_802 (O_802,N_14718,N_14942);
and UO_803 (O_803,N_14822,N_14381);
and UO_804 (O_804,N_14620,N_14856);
and UO_805 (O_805,N_14815,N_14942);
and UO_806 (O_806,N_14389,N_14916);
nor UO_807 (O_807,N_14520,N_14840);
or UO_808 (O_808,N_14898,N_14552);
nand UO_809 (O_809,N_14275,N_14267);
xor UO_810 (O_810,N_14859,N_14552);
or UO_811 (O_811,N_14725,N_14608);
or UO_812 (O_812,N_14938,N_14794);
and UO_813 (O_813,N_14433,N_14531);
nor UO_814 (O_814,N_14763,N_14895);
nor UO_815 (O_815,N_14313,N_14441);
nor UO_816 (O_816,N_14468,N_14569);
xor UO_817 (O_817,N_14673,N_14888);
or UO_818 (O_818,N_14901,N_14384);
xor UO_819 (O_819,N_14293,N_14806);
nor UO_820 (O_820,N_14566,N_14885);
or UO_821 (O_821,N_14721,N_14258);
nor UO_822 (O_822,N_14445,N_14984);
nor UO_823 (O_823,N_14360,N_14291);
xor UO_824 (O_824,N_14260,N_14306);
xnor UO_825 (O_825,N_14438,N_14665);
nand UO_826 (O_826,N_14413,N_14429);
nor UO_827 (O_827,N_14333,N_14747);
nor UO_828 (O_828,N_14940,N_14902);
nand UO_829 (O_829,N_14436,N_14580);
nor UO_830 (O_830,N_14694,N_14630);
nand UO_831 (O_831,N_14339,N_14808);
nand UO_832 (O_832,N_14783,N_14540);
xor UO_833 (O_833,N_14762,N_14951);
nor UO_834 (O_834,N_14360,N_14401);
and UO_835 (O_835,N_14258,N_14961);
or UO_836 (O_836,N_14303,N_14717);
nand UO_837 (O_837,N_14869,N_14516);
nor UO_838 (O_838,N_14950,N_14627);
and UO_839 (O_839,N_14468,N_14302);
and UO_840 (O_840,N_14942,N_14503);
and UO_841 (O_841,N_14855,N_14264);
or UO_842 (O_842,N_14962,N_14687);
nand UO_843 (O_843,N_14498,N_14981);
nand UO_844 (O_844,N_14498,N_14493);
nor UO_845 (O_845,N_14543,N_14270);
nand UO_846 (O_846,N_14812,N_14830);
or UO_847 (O_847,N_14281,N_14345);
nor UO_848 (O_848,N_14345,N_14867);
and UO_849 (O_849,N_14958,N_14871);
nand UO_850 (O_850,N_14946,N_14848);
or UO_851 (O_851,N_14595,N_14861);
and UO_852 (O_852,N_14979,N_14347);
nand UO_853 (O_853,N_14764,N_14464);
and UO_854 (O_854,N_14436,N_14395);
nor UO_855 (O_855,N_14552,N_14848);
or UO_856 (O_856,N_14514,N_14843);
xor UO_857 (O_857,N_14579,N_14260);
xnor UO_858 (O_858,N_14937,N_14805);
xor UO_859 (O_859,N_14789,N_14687);
or UO_860 (O_860,N_14527,N_14367);
and UO_861 (O_861,N_14813,N_14296);
and UO_862 (O_862,N_14605,N_14407);
nor UO_863 (O_863,N_14319,N_14986);
nor UO_864 (O_864,N_14498,N_14706);
xnor UO_865 (O_865,N_14521,N_14732);
nor UO_866 (O_866,N_14692,N_14978);
nor UO_867 (O_867,N_14383,N_14963);
nor UO_868 (O_868,N_14694,N_14855);
and UO_869 (O_869,N_14592,N_14507);
nor UO_870 (O_870,N_14800,N_14880);
xor UO_871 (O_871,N_14736,N_14989);
nand UO_872 (O_872,N_14547,N_14411);
and UO_873 (O_873,N_14281,N_14710);
nor UO_874 (O_874,N_14900,N_14762);
nand UO_875 (O_875,N_14376,N_14511);
and UO_876 (O_876,N_14962,N_14452);
and UO_877 (O_877,N_14880,N_14484);
xor UO_878 (O_878,N_14312,N_14501);
or UO_879 (O_879,N_14767,N_14748);
or UO_880 (O_880,N_14491,N_14627);
nand UO_881 (O_881,N_14921,N_14742);
nor UO_882 (O_882,N_14594,N_14282);
and UO_883 (O_883,N_14717,N_14681);
nor UO_884 (O_884,N_14478,N_14338);
nand UO_885 (O_885,N_14556,N_14784);
or UO_886 (O_886,N_14410,N_14366);
nor UO_887 (O_887,N_14453,N_14933);
nand UO_888 (O_888,N_14299,N_14546);
and UO_889 (O_889,N_14877,N_14280);
xor UO_890 (O_890,N_14806,N_14807);
or UO_891 (O_891,N_14429,N_14558);
nor UO_892 (O_892,N_14429,N_14345);
and UO_893 (O_893,N_14317,N_14904);
nor UO_894 (O_894,N_14378,N_14722);
or UO_895 (O_895,N_14984,N_14983);
nor UO_896 (O_896,N_14953,N_14669);
or UO_897 (O_897,N_14484,N_14554);
or UO_898 (O_898,N_14954,N_14269);
nor UO_899 (O_899,N_14587,N_14850);
or UO_900 (O_900,N_14376,N_14454);
nand UO_901 (O_901,N_14823,N_14950);
and UO_902 (O_902,N_14594,N_14313);
nand UO_903 (O_903,N_14587,N_14314);
or UO_904 (O_904,N_14880,N_14778);
nand UO_905 (O_905,N_14675,N_14960);
or UO_906 (O_906,N_14757,N_14475);
and UO_907 (O_907,N_14973,N_14355);
nor UO_908 (O_908,N_14924,N_14576);
nor UO_909 (O_909,N_14808,N_14639);
or UO_910 (O_910,N_14988,N_14857);
or UO_911 (O_911,N_14597,N_14989);
nor UO_912 (O_912,N_14535,N_14993);
nand UO_913 (O_913,N_14410,N_14511);
nor UO_914 (O_914,N_14352,N_14503);
or UO_915 (O_915,N_14346,N_14281);
or UO_916 (O_916,N_14806,N_14707);
nor UO_917 (O_917,N_14483,N_14311);
and UO_918 (O_918,N_14819,N_14405);
nor UO_919 (O_919,N_14647,N_14745);
nor UO_920 (O_920,N_14813,N_14767);
nand UO_921 (O_921,N_14997,N_14898);
nand UO_922 (O_922,N_14806,N_14390);
or UO_923 (O_923,N_14878,N_14783);
and UO_924 (O_924,N_14722,N_14970);
xor UO_925 (O_925,N_14763,N_14438);
nor UO_926 (O_926,N_14568,N_14822);
or UO_927 (O_927,N_14589,N_14867);
nand UO_928 (O_928,N_14922,N_14992);
or UO_929 (O_929,N_14714,N_14338);
nor UO_930 (O_930,N_14963,N_14797);
nor UO_931 (O_931,N_14882,N_14813);
nor UO_932 (O_932,N_14608,N_14440);
and UO_933 (O_933,N_14763,N_14697);
and UO_934 (O_934,N_14544,N_14699);
nor UO_935 (O_935,N_14559,N_14750);
nor UO_936 (O_936,N_14857,N_14415);
nor UO_937 (O_937,N_14418,N_14917);
or UO_938 (O_938,N_14957,N_14346);
or UO_939 (O_939,N_14572,N_14271);
or UO_940 (O_940,N_14467,N_14606);
or UO_941 (O_941,N_14421,N_14452);
nor UO_942 (O_942,N_14476,N_14393);
and UO_943 (O_943,N_14369,N_14480);
or UO_944 (O_944,N_14836,N_14611);
and UO_945 (O_945,N_14547,N_14687);
nor UO_946 (O_946,N_14859,N_14855);
or UO_947 (O_947,N_14401,N_14560);
xnor UO_948 (O_948,N_14656,N_14450);
nor UO_949 (O_949,N_14597,N_14467);
and UO_950 (O_950,N_14678,N_14571);
nand UO_951 (O_951,N_14422,N_14748);
nor UO_952 (O_952,N_14530,N_14551);
and UO_953 (O_953,N_14698,N_14409);
nand UO_954 (O_954,N_14353,N_14996);
nor UO_955 (O_955,N_14511,N_14841);
nand UO_956 (O_956,N_14275,N_14728);
xor UO_957 (O_957,N_14775,N_14538);
or UO_958 (O_958,N_14986,N_14276);
or UO_959 (O_959,N_14548,N_14751);
and UO_960 (O_960,N_14387,N_14924);
nand UO_961 (O_961,N_14309,N_14826);
and UO_962 (O_962,N_14921,N_14975);
nand UO_963 (O_963,N_14813,N_14535);
and UO_964 (O_964,N_14661,N_14800);
or UO_965 (O_965,N_14823,N_14418);
nand UO_966 (O_966,N_14275,N_14841);
nand UO_967 (O_967,N_14462,N_14576);
and UO_968 (O_968,N_14563,N_14933);
nor UO_969 (O_969,N_14625,N_14342);
nand UO_970 (O_970,N_14761,N_14417);
nor UO_971 (O_971,N_14759,N_14291);
nor UO_972 (O_972,N_14318,N_14383);
nand UO_973 (O_973,N_14622,N_14640);
and UO_974 (O_974,N_14467,N_14360);
or UO_975 (O_975,N_14937,N_14362);
and UO_976 (O_976,N_14759,N_14460);
nor UO_977 (O_977,N_14411,N_14260);
nand UO_978 (O_978,N_14782,N_14723);
nand UO_979 (O_979,N_14364,N_14415);
nor UO_980 (O_980,N_14781,N_14411);
and UO_981 (O_981,N_14954,N_14756);
or UO_982 (O_982,N_14638,N_14679);
nand UO_983 (O_983,N_14558,N_14610);
and UO_984 (O_984,N_14954,N_14774);
and UO_985 (O_985,N_14949,N_14971);
nor UO_986 (O_986,N_14793,N_14959);
nor UO_987 (O_987,N_14297,N_14589);
nand UO_988 (O_988,N_14859,N_14823);
or UO_989 (O_989,N_14531,N_14727);
or UO_990 (O_990,N_14367,N_14887);
and UO_991 (O_991,N_14860,N_14312);
nor UO_992 (O_992,N_14417,N_14700);
or UO_993 (O_993,N_14942,N_14817);
or UO_994 (O_994,N_14737,N_14484);
nor UO_995 (O_995,N_14259,N_14869);
xnor UO_996 (O_996,N_14462,N_14582);
xnor UO_997 (O_997,N_14930,N_14506);
nand UO_998 (O_998,N_14896,N_14573);
and UO_999 (O_999,N_14482,N_14337);
nor UO_1000 (O_1000,N_14894,N_14808);
nor UO_1001 (O_1001,N_14921,N_14328);
or UO_1002 (O_1002,N_14566,N_14989);
nor UO_1003 (O_1003,N_14290,N_14685);
or UO_1004 (O_1004,N_14584,N_14443);
or UO_1005 (O_1005,N_14391,N_14492);
nand UO_1006 (O_1006,N_14847,N_14869);
or UO_1007 (O_1007,N_14894,N_14489);
nand UO_1008 (O_1008,N_14505,N_14809);
or UO_1009 (O_1009,N_14489,N_14857);
nand UO_1010 (O_1010,N_14589,N_14663);
nand UO_1011 (O_1011,N_14561,N_14527);
or UO_1012 (O_1012,N_14553,N_14480);
nand UO_1013 (O_1013,N_14624,N_14361);
nor UO_1014 (O_1014,N_14954,N_14845);
nor UO_1015 (O_1015,N_14936,N_14753);
xor UO_1016 (O_1016,N_14687,N_14496);
and UO_1017 (O_1017,N_14465,N_14700);
or UO_1018 (O_1018,N_14600,N_14792);
and UO_1019 (O_1019,N_14905,N_14988);
and UO_1020 (O_1020,N_14655,N_14928);
nor UO_1021 (O_1021,N_14784,N_14672);
and UO_1022 (O_1022,N_14551,N_14466);
nor UO_1023 (O_1023,N_14843,N_14496);
nor UO_1024 (O_1024,N_14433,N_14411);
and UO_1025 (O_1025,N_14910,N_14867);
and UO_1026 (O_1026,N_14735,N_14286);
xnor UO_1027 (O_1027,N_14586,N_14378);
nor UO_1028 (O_1028,N_14706,N_14460);
xor UO_1029 (O_1029,N_14797,N_14477);
nor UO_1030 (O_1030,N_14661,N_14342);
nor UO_1031 (O_1031,N_14980,N_14821);
and UO_1032 (O_1032,N_14711,N_14563);
or UO_1033 (O_1033,N_14282,N_14584);
and UO_1034 (O_1034,N_14847,N_14770);
nand UO_1035 (O_1035,N_14977,N_14263);
nor UO_1036 (O_1036,N_14578,N_14383);
xnor UO_1037 (O_1037,N_14764,N_14795);
nor UO_1038 (O_1038,N_14895,N_14952);
xnor UO_1039 (O_1039,N_14801,N_14815);
or UO_1040 (O_1040,N_14338,N_14262);
nand UO_1041 (O_1041,N_14622,N_14279);
and UO_1042 (O_1042,N_14422,N_14993);
nor UO_1043 (O_1043,N_14436,N_14388);
nor UO_1044 (O_1044,N_14845,N_14696);
nand UO_1045 (O_1045,N_14724,N_14767);
and UO_1046 (O_1046,N_14266,N_14362);
nor UO_1047 (O_1047,N_14548,N_14283);
and UO_1048 (O_1048,N_14274,N_14774);
nor UO_1049 (O_1049,N_14291,N_14290);
xor UO_1050 (O_1050,N_14809,N_14971);
or UO_1051 (O_1051,N_14487,N_14946);
nor UO_1052 (O_1052,N_14546,N_14605);
or UO_1053 (O_1053,N_14737,N_14322);
and UO_1054 (O_1054,N_14523,N_14271);
and UO_1055 (O_1055,N_14720,N_14662);
nand UO_1056 (O_1056,N_14595,N_14503);
or UO_1057 (O_1057,N_14798,N_14389);
nand UO_1058 (O_1058,N_14560,N_14573);
nand UO_1059 (O_1059,N_14913,N_14768);
and UO_1060 (O_1060,N_14856,N_14654);
or UO_1061 (O_1061,N_14697,N_14922);
and UO_1062 (O_1062,N_14370,N_14494);
nor UO_1063 (O_1063,N_14439,N_14564);
nor UO_1064 (O_1064,N_14975,N_14843);
nand UO_1065 (O_1065,N_14713,N_14581);
and UO_1066 (O_1066,N_14577,N_14712);
or UO_1067 (O_1067,N_14817,N_14969);
nand UO_1068 (O_1068,N_14567,N_14518);
nor UO_1069 (O_1069,N_14348,N_14495);
nor UO_1070 (O_1070,N_14938,N_14377);
nor UO_1071 (O_1071,N_14822,N_14948);
nor UO_1072 (O_1072,N_14358,N_14638);
xnor UO_1073 (O_1073,N_14460,N_14888);
xor UO_1074 (O_1074,N_14631,N_14635);
and UO_1075 (O_1075,N_14508,N_14711);
nand UO_1076 (O_1076,N_14677,N_14480);
and UO_1077 (O_1077,N_14546,N_14457);
and UO_1078 (O_1078,N_14856,N_14364);
and UO_1079 (O_1079,N_14686,N_14499);
and UO_1080 (O_1080,N_14802,N_14920);
and UO_1081 (O_1081,N_14938,N_14529);
nand UO_1082 (O_1082,N_14851,N_14892);
nor UO_1083 (O_1083,N_14450,N_14411);
nand UO_1084 (O_1084,N_14547,N_14490);
and UO_1085 (O_1085,N_14562,N_14876);
or UO_1086 (O_1086,N_14302,N_14995);
nand UO_1087 (O_1087,N_14277,N_14292);
nand UO_1088 (O_1088,N_14738,N_14289);
or UO_1089 (O_1089,N_14688,N_14337);
or UO_1090 (O_1090,N_14837,N_14845);
nor UO_1091 (O_1091,N_14260,N_14362);
nand UO_1092 (O_1092,N_14367,N_14729);
or UO_1093 (O_1093,N_14669,N_14587);
or UO_1094 (O_1094,N_14713,N_14398);
nand UO_1095 (O_1095,N_14930,N_14379);
or UO_1096 (O_1096,N_14893,N_14707);
xor UO_1097 (O_1097,N_14485,N_14877);
nor UO_1098 (O_1098,N_14915,N_14372);
nand UO_1099 (O_1099,N_14501,N_14346);
nand UO_1100 (O_1100,N_14387,N_14559);
nor UO_1101 (O_1101,N_14422,N_14843);
xor UO_1102 (O_1102,N_14536,N_14565);
and UO_1103 (O_1103,N_14537,N_14293);
nand UO_1104 (O_1104,N_14515,N_14671);
and UO_1105 (O_1105,N_14528,N_14277);
nor UO_1106 (O_1106,N_14671,N_14640);
nor UO_1107 (O_1107,N_14271,N_14660);
and UO_1108 (O_1108,N_14621,N_14753);
xnor UO_1109 (O_1109,N_14593,N_14607);
nor UO_1110 (O_1110,N_14490,N_14992);
nand UO_1111 (O_1111,N_14475,N_14729);
nor UO_1112 (O_1112,N_14735,N_14826);
xor UO_1113 (O_1113,N_14862,N_14831);
and UO_1114 (O_1114,N_14787,N_14973);
nand UO_1115 (O_1115,N_14302,N_14692);
nor UO_1116 (O_1116,N_14342,N_14838);
nor UO_1117 (O_1117,N_14446,N_14496);
nor UO_1118 (O_1118,N_14295,N_14842);
nand UO_1119 (O_1119,N_14333,N_14847);
nand UO_1120 (O_1120,N_14798,N_14343);
and UO_1121 (O_1121,N_14968,N_14643);
xor UO_1122 (O_1122,N_14347,N_14492);
or UO_1123 (O_1123,N_14254,N_14709);
or UO_1124 (O_1124,N_14832,N_14917);
nand UO_1125 (O_1125,N_14489,N_14440);
and UO_1126 (O_1126,N_14811,N_14611);
nand UO_1127 (O_1127,N_14745,N_14770);
nor UO_1128 (O_1128,N_14999,N_14389);
and UO_1129 (O_1129,N_14747,N_14314);
and UO_1130 (O_1130,N_14688,N_14951);
and UO_1131 (O_1131,N_14294,N_14549);
nor UO_1132 (O_1132,N_14654,N_14352);
or UO_1133 (O_1133,N_14784,N_14906);
nor UO_1134 (O_1134,N_14558,N_14750);
and UO_1135 (O_1135,N_14545,N_14824);
nand UO_1136 (O_1136,N_14415,N_14398);
nor UO_1137 (O_1137,N_14630,N_14942);
and UO_1138 (O_1138,N_14316,N_14466);
nor UO_1139 (O_1139,N_14784,N_14352);
nand UO_1140 (O_1140,N_14961,N_14524);
or UO_1141 (O_1141,N_14789,N_14978);
or UO_1142 (O_1142,N_14409,N_14272);
nor UO_1143 (O_1143,N_14371,N_14604);
or UO_1144 (O_1144,N_14432,N_14557);
nor UO_1145 (O_1145,N_14340,N_14283);
or UO_1146 (O_1146,N_14694,N_14342);
nor UO_1147 (O_1147,N_14649,N_14290);
xor UO_1148 (O_1148,N_14373,N_14388);
or UO_1149 (O_1149,N_14666,N_14722);
xnor UO_1150 (O_1150,N_14645,N_14459);
nand UO_1151 (O_1151,N_14326,N_14421);
nor UO_1152 (O_1152,N_14525,N_14859);
nor UO_1153 (O_1153,N_14978,N_14449);
xnor UO_1154 (O_1154,N_14933,N_14281);
nor UO_1155 (O_1155,N_14468,N_14710);
or UO_1156 (O_1156,N_14346,N_14711);
nor UO_1157 (O_1157,N_14723,N_14594);
or UO_1158 (O_1158,N_14311,N_14841);
nor UO_1159 (O_1159,N_14931,N_14328);
and UO_1160 (O_1160,N_14876,N_14811);
or UO_1161 (O_1161,N_14739,N_14665);
nand UO_1162 (O_1162,N_14933,N_14961);
or UO_1163 (O_1163,N_14428,N_14291);
nand UO_1164 (O_1164,N_14613,N_14518);
nand UO_1165 (O_1165,N_14334,N_14512);
and UO_1166 (O_1166,N_14806,N_14862);
or UO_1167 (O_1167,N_14769,N_14469);
xnor UO_1168 (O_1168,N_14824,N_14371);
nor UO_1169 (O_1169,N_14331,N_14330);
nor UO_1170 (O_1170,N_14845,N_14506);
and UO_1171 (O_1171,N_14461,N_14340);
nand UO_1172 (O_1172,N_14640,N_14752);
nand UO_1173 (O_1173,N_14257,N_14720);
nand UO_1174 (O_1174,N_14819,N_14815);
nor UO_1175 (O_1175,N_14541,N_14463);
or UO_1176 (O_1176,N_14655,N_14990);
or UO_1177 (O_1177,N_14393,N_14787);
and UO_1178 (O_1178,N_14455,N_14323);
nand UO_1179 (O_1179,N_14908,N_14303);
and UO_1180 (O_1180,N_14572,N_14511);
and UO_1181 (O_1181,N_14832,N_14895);
and UO_1182 (O_1182,N_14815,N_14473);
nor UO_1183 (O_1183,N_14929,N_14821);
or UO_1184 (O_1184,N_14766,N_14686);
and UO_1185 (O_1185,N_14698,N_14622);
nor UO_1186 (O_1186,N_14956,N_14891);
or UO_1187 (O_1187,N_14990,N_14457);
nand UO_1188 (O_1188,N_14711,N_14357);
and UO_1189 (O_1189,N_14312,N_14959);
nor UO_1190 (O_1190,N_14770,N_14346);
and UO_1191 (O_1191,N_14641,N_14315);
and UO_1192 (O_1192,N_14593,N_14878);
or UO_1193 (O_1193,N_14617,N_14579);
xor UO_1194 (O_1194,N_14675,N_14662);
or UO_1195 (O_1195,N_14433,N_14809);
or UO_1196 (O_1196,N_14308,N_14699);
or UO_1197 (O_1197,N_14904,N_14405);
and UO_1198 (O_1198,N_14765,N_14620);
or UO_1199 (O_1199,N_14816,N_14528);
nor UO_1200 (O_1200,N_14983,N_14466);
nand UO_1201 (O_1201,N_14460,N_14814);
or UO_1202 (O_1202,N_14880,N_14796);
or UO_1203 (O_1203,N_14924,N_14993);
and UO_1204 (O_1204,N_14584,N_14747);
and UO_1205 (O_1205,N_14768,N_14736);
and UO_1206 (O_1206,N_14488,N_14448);
nand UO_1207 (O_1207,N_14827,N_14971);
nor UO_1208 (O_1208,N_14372,N_14920);
or UO_1209 (O_1209,N_14268,N_14327);
nand UO_1210 (O_1210,N_14330,N_14265);
xnor UO_1211 (O_1211,N_14766,N_14342);
xor UO_1212 (O_1212,N_14612,N_14503);
or UO_1213 (O_1213,N_14641,N_14772);
or UO_1214 (O_1214,N_14514,N_14586);
or UO_1215 (O_1215,N_14886,N_14991);
nand UO_1216 (O_1216,N_14492,N_14897);
or UO_1217 (O_1217,N_14627,N_14715);
nor UO_1218 (O_1218,N_14701,N_14326);
nand UO_1219 (O_1219,N_14891,N_14660);
nor UO_1220 (O_1220,N_14347,N_14447);
nor UO_1221 (O_1221,N_14407,N_14504);
nand UO_1222 (O_1222,N_14327,N_14640);
nand UO_1223 (O_1223,N_14821,N_14534);
nand UO_1224 (O_1224,N_14947,N_14497);
and UO_1225 (O_1225,N_14715,N_14420);
nand UO_1226 (O_1226,N_14484,N_14343);
xor UO_1227 (O_1227,N_14861,N_14497);
or UO_1228 (O_1228,N_14432,N_14742);
or UO_1229 (O_1229,N_14338,N_14622);
xnor UO_1230 (O_1230,N_14337,N_14622);
or UO_1231 (O_1231,N_14465,N_14305);
nand UO_1232 (O_1232,N_14940,N_14574);
nand UO_1233 (O_1233,N_14274,N_14847);
or UO_1234 (O_1234,N_14507,N_14320);
or UO_1235 (O_1235,N_14367,N_14807);
nor UO_1236 (O_1236,N_14474,N_14831);
and UO_1237 (O_1237,N_14720,N_14353);
and UO_1238 (O_1238,N_14633,N_14611);
nand UO_1239 (O_1239,N_14995,N_14743);
nand UO_1240 (O_1240,N_14479,N_14938);
nand UO_1241 (O_1241,N_14283,N_14613);
nor UO_1242 (O_1242,N_14291,N_14380);
nand UO_1243 (O_1243,N_14993,N_14910);
or UO_1244 (O_1244,N_14933,N_14644);
nor UO_1245 (O_1245,N_14585,N_14261);
or UO_1246 (O_1246,N_14735,N_14495);
and UO_1247 (O_1247,N_14302,N_14861);
or UO_1248 (O_1248,N_14313,N_14661);
nand UO_1249 (O_1249,N_14973,N_14705);
nor UO_1250 (O_1250,N_14940,N_14850);
or UO_1251 (O_1251,N_14953,N_14295);
or UO_1252 (O_1252,N_14719,N_14971);
nor UO_1253 (O_1253,N_14710,N_14601);
or UO_1254 (O_1254,N_14311,N_14605);
and UO_1255 (O_1255,N_14915,N_14570);
and UO_1256 (O_1256,N_14914,N_14455);
nor UO_1257 (O_1257,N_14814,N_14762);
nor UO_1258 (O_1258,N_14453,N_14624);
nand UO_1259 (O_1259,N_14309,N_14310);
nand UO_1260 (O_1260,N_14649,N_14634);
nand UO_1261 (O_1261,N_14700,N_14399);
xnor UO_1262 (O_1262,N_14508,N_14611);
and UO_1263 (O_1263,N_14978,N_14973);
or UO_1264 (O_1264,N_14962,N_14837);
nand UO_1265 (O_1265,N_14412,N_14491);
xnor UO_1266 (O_1266,N_14640,N_14331);
nor UO_1267 (O_1267,N_14915,N_14482);
and UO_1268 (O_1268,N_14615,N_14679);
xnor UO_1269 (O_1269,N_14766,N_14284);
and UO_1270 (O_1270,N_14864,N_14806);
xor UO_1271 (O_1271,N_14355,N_14674);
nor UO_1272 (O_1272,N_14528,N_14455);
and UO_1273 (O_1273,N_14522,N_14476);
or UO_1274 (O_1274,N_14690,N_14529);
xnor UO_1275 (O_1275,N_14795,N_14801);
and UO_1276 (O_1276,N_14565,N_14878);
and UO_1277 (O_1277,N_14480,N_14889);
nand UO_1278 (O_1278,N_14636,N_14454);
nand UO_1279 (O_1279,N_14434,N_14469);
or UO_1280 (O_1280,N_14724,N_14590);
nand UO_1281 (O_1281,N_14362,N_14830);
and UO_1282 (O_1282,N_14419,N_14913);
nand UO_1283 (O_1283,N_14971,N_14816);
nand UO_1284 (O_1284,N_14256,N_14656);
xor UO_1285 (O_1285,N_14483,N_14430);
or UO_1286 (O_1286,N_14439,N_14716);
and UO_1287 (O_1287,N_14605,N_14451);
and UO_1288 (O_1288,N_14979,N_14563);
and UO_1289 (O_1289,N_14854,N_14277);
or UO_1290 (O_1290,N_14917,N_14854);
and UO_1291 (O_1291,N_14647,N_14830);
or UO_1292 (O_1292,N_14814,N_14348);
xnor UO_1293 (O_1293,N_14942,N_14896);
nor UO_1294 (O_1294,N_14728,N_14365);
nand UO_1295 (O_1295,N_14615,N_14920);
and UO_1296 (O_1296,N_14785,N_14633);
xnor UO_1297 (O_1297,N_14754,N_14271);
nand UO_1298 (O_1298,N_14431,N_14348);
xor UO_1299 (O_1299,N_14339,N_14900);
nand UO_1300 (O_1300,N_14825,N_14900);
xnor UO_1301 (O_1301,N_14950,N_14312);
nor UO_1302 (O_1302,N_14618,N_14335);
or UO_1303 (O_1303,N_14928,N_14802);
and UO_1304 (O_1304,N_14425,N_14736);
nand UO_1305 (O_1305,N_14915,N_14807);
or UO_1306 (O_1306,N_14652,N_14883);
nand UO_1307 (O_1307,N_14299,N_14317);
or UO_1308 (O_1308,N_14303,N_14481);
and UO_1309 (O_1309,N_14297,N_14912);
xnor UO_1310 (O_1310,N_14683,N_14477);
and UO_1311 (O_1311,N_14800,N_14687);
and UO_1312 (O_1312,N_14494,N_14408);
and UO_1313 (O_1313,N_14533,N_14978);
xor UO_1314 (O_1314,N_14647,N_14258);
nor UO_1315 (O_1315,N_14364,N_14421);
xor UO_1316 (O_1316,N_14823,N_14691);
or UO_1317 (O_1317,N_14670,N_14363);
nand UO_1318 (O_1318,N_14534,N_14813);
nor UO_1319 (O_1319,N_14938,N_14420);
nor UO_1320 (O_1320,N_14552,N_14269);
nor UO_1321 (O_1321,N_14974,N_14895);
and UO_1322 (O_1322,N_14910,N_14780);
or UO_1323 (O_1323,N_14763,N_14998);
nor UO_1324 (O_1324,N_14316,N_14915);
xnor UO_1325 (O_1325,N_14736,N_14757);
nor UO_1326 (O_1326,N_14534,N_14501);
nor UO_1327 (O_1327,N_14600,N_14737);
nor UO_1328 (O_1328,N_14290,N_14896);
nor UO_1329 (O_1329,N_14736,N_14432);
and UO_1330 (O_1330,N_14573,N_14867);
nand UO_1331 (O_1331,N_14587,N_14279);
nor UO_1332 (O_1332,N_14954,N_14321);
and UO_1333 (O_1333,N_14870,N_14635);
nand UO_1334 (O_1334,N_14700,N_14480);
nand UO_1335 (O_1335,N_14333,N_14622);
or UO_1336 (O_1336,N_14852,N_14348);
nand UO_1337 (O_1337,N_14808,N_14387);
and UO_1338 (O_1338,N_14717,N_14807);
nor UO_1339 (O_1339,N_14291,N_14455);
nand UO_1340 (O_1340,N_14952,N_14415);
and UO_1341 (O_1341,N_14298,N_14411);
nand UO_1342 (O_1342,N_14887,N_14780);
and UO_1343 (O_1343,N_14813,N_14872);
nor UO_1344 (O_1344,N_14636,N_14642);
or UO_1345 (O_1345,N_14505,N_14949);
nor UO_1346 (O_1346,N_14597,N_14414);
or UO_1347 (O_1347,N_14520,N_14598);
or UO_1348 (O_1348,N_14623,N_14359);
nor UO_1349 (O_1349,N_14890,N_14441);
or UO_1350 (O_1350,N_14289,N_14910);
xor UO_1351 (O_1351,N_14654,N_14467);
or UO_1352 (O_1352,N_14664,N_14416);
and UO_1353 (O_1353,N_14550,N_14391);
nand UO_1354 (O_1354,N_14640,N_14918);
nor UO_1355 (O_1355,N_14738,N_14733);
and UO_1356 (O_1356,N_14455,N_14788);
and UO_1357 (O_1357,N_14878,N_14281);
and UO_1358 (O_1358,N_14798,N_14356);
nand UO_1359 (O_1359,N_14690,N_14369);
nor UO_1360 (O_1360,N_14415,N_14589);
nor UO_1361 (O_1361,N_14287,N_14648);
or UO_1362 (O_1362,N_14875,N_14373);
nor UO_1363 (O_1363,N_14436,N_14511);
or UO_1364 (O_1364,N_14444,N_14681);
nand UO_1365 (O_1365,N_14557,N_14383);
xnor UO_1366 (O_1366,N_14707,N_14349);
nand UO_1367 (O_1367,N_14609,N_14982);
nand UO_1368 (O_1368,N_14872,N_14628);
nor UO_1369 (O_1369,N_14353,N_14921);
and UO_1370 (O_1370,N_14279,N_14673);
or UO_1371 (O_1371,N_14431,N_14511);
xnor UO_1372 (O_1372,N_14865,N_14923);
nor UO_1373 (O_1373,N_14643,N_14471);
nor UO_1374 (O_1374,N_14712,N_14623);
nand UO_1375 (O_1375,N_14353,N_14261);
nor UO_1376 (O_1376,N_14629,N_14416);
nor UO_1377 (O_1377,N_14363,N_14976);
or UO_1378 (O_1378,N_14992,N_14967);
or UO_1379 (O_1379,N_14382,N_14410);
xor UO_1380 (O_1380,N_14522,N_14773);
nand UO_1381 (O_1381,N_14672,N_14967);
or UO_1382 (O_1382,N_14357,N_14697);
nand UO_1383 (O_1383,N_14846,N_14553);
or UO_1384 (O_1384,N_14614,N_14281);
xnor UO_1385 (O_1385,N_14959,N_14710);
or UO_1386 (O_1386,N_14785,N_14699);
xor UO_1387 (O_1387,N_14330,N_14811);
or UO_1388 (O_1388,N_14678,N_14849);
and UO_1389 (O_1389,N_14509,N_14486);
nand UO_1390 (O_1390,N_14450,N_14483);
nand UO_1391 (O_1391,N_14680,N_14579);
nand UO_1392 (O_1392,N_14510,N_14344);
or UO_1393 (O_1393,N_14824,N_14568);
nor UO_1394 (O_1394,N_14282,N_14432);
and UO_1395 (O_1395,N_14283,N_14941);
and UO_1396 (O_1396,N_14876,N_14750);
or UO_1397 (O_1397,N_14719,N_14941);
or UO_1398 (O_1398,N_14416,N_14572);
nand UO_1399 (O_1399,N_14949,N_14594);
nand UO_1400 (O_1400,N_14815,N_14875);
nand UO_1401 (O_1401,N_14624,N_14696);
and UO_1402 (O_1402,N_14381,N_14278);
or UO_1403 (O_1403,N_14877,N_14809);
and UO_1404 (O_1404,N_14321,N_14412);
nand UO_1405 (O_1405,N_14513,N_14915);
nand UO_1406 (O_1406,N_14733,N_14456);
and UO_1407 (O_1407,N_14270,N_14860);
nand UO_1408 (O_1408,N_14477,N_14287);
and UO_1409 (O_1409,N_14801,N_14285);
and UO_1410 (O_1410,N_14399,N_14599);
nor UO_1411 (O_1411,N_14838,N_14753);
and UO_1412 (O_1412,N_14887,N_14810);
nor UO_1413 (O_1413,N_14401,N_14367);
nand UO_1414 (O_1414,N_14838,N_14483);
nor UO_1415 (O_1415,N_14435,N_14687);
or UO_1416 (O_1416,N_14951,N_14992);
nand UO_1417 (O_1417,N_14872,N_14574);
and UO_1418 (O_1418,N_14366,N_14688);
nand UO_1419 (O_1419,N_14311,N_14900);
and UO_1420 (O_1420,N_14953,N_14331);
nand UO_1421 (O_1421,N_14281,N_14647);
nand UO_1422 (O_1422,N_14508,N_14885);
nor UO_1423 (O_1423,N_14327,N_14719);
nand UO_1424 (O_1424,N_14732,N_14451);
or UO_1425 (O_1425,N_14488,N_14320);
nor UO_1426 (O_1426,N_14418,N_14705);
and UO_1427 (O_1427,N_14883,N_14990);
nand UO_1428 (O_1428,N_14803,N_14618);
nand UO_1429 (O_1429,N_14774,N_14351);
nand UO_1430 (O_1430,N_14345,N_14363);
nand UO_1431 (O_1431,N_14517,N_14831);
or UO_1432 (O_1432,N_14822,N_14375);
and UO_1433 (O_1433,N_14314,N_14764);
nor UO_1434 (O_1434,N_14265,N_14349);
and UO_1435 (O_1435,N_14624,N_14597);
nor UO_1436 (O_1436,N_14558,N_14975);
and UO_1437 (O_1437,N_14399,N_14685);
nand UO_1438 (O_1438,N_14317,N_14919);
nor UO_1439 (O_1439,N_14562,N_14309);
nand UO_1440 (O_1440,N_14812,N_14965);
or UO_1441 (O_1441,N_14620,N_14938);
nor UO_1442 (O_1442,N_14413,N_14503);
nor UO_1443 (O_1443,N_14314,N_14350);
or UO_1444 (O_1444,N_14607,N_14544);
nor UO_1445 (O_1445,N_14387,N_14463);
nand UO_1446 (O_1446,N_14277,N_14326);
nor UO_1447 (O_1447,N_14943,N_14484);
or UO_1448 (O_1448,N_14938,N_14623);
and UO_1449 (O_1449,N_14637,N_14499);
and UO_1450 (O_1450,N_14462,N_14850);
or UO_1451 (O_1451,N_14658,N_14902);
or UO_1452 (O_1452,N_14417,N_14566);
xnor UO_1453 (O_1453,N_14750,N_14695);
nor UO_1454 (O_1454,N_14898,N_14331);
and UO_1455 (O_1455,N_14467,N_14873);
xnor UO_1456 (O_1456,N_14926,N_14700);
nand UO_1457 (O_1457,N_14447,N_14800);
nor UO_1458 (O_1458,N_14470,N_14824);
and UO_1459 (O_1459,N_14559,N_14597);
nand UO_1460 (O_1460,N_14443,N_14505);
nand UO_1461 (O_1461,N_14328,N_14780);
nor UO_1462 (O_1462,N_14763,N_14633);
and UO_1463 (O_1463,N_14395,N_14473);
nand UO_1464 (O_1464,N_14886,N_14686);
and UO_1465 (O_1465,N_14944,N_14513);
and UO_1466 (O_1466,N_14824,N_14961);
nor UO_1467 (O_1467,N_14347,N_14739);
xor UO_1468 (O_1468,N_14833,N_14902);
and UO_1469 (O_1469,N_14956,N_14353);
nor UO_1470 (O_1470,N_14835,N_14625);
or UO_1471 (O_1471,N_14728,N_14510);
nand UO_1472 (O_1472,N_14443,N_14955);
and UO_1473 (O_1473,N_14512,N_14320);
nor UO_1474 (O_1474,N_14354,N_14884);
and UO_1475 (O_1475,N_14400,N_14561);
or UO_1476 (O_1476,N_14941,N_14361);
or UO_1477 (O_1477,N_14390,N_14888);
and UO_1478 (O_1478,N_14565,N_14371);
xnor UO_1479 (O_1479,N_14866,N_14371);
nor UO_1480 (O_1480,N_14521,N_14544);
nand UO_1481 (O_1481,N_14528,N_14266);
nor UO_1482 (O_1482,N_14937,N_14337);
and UO_1483 (O_1483,N_14725,N_14761);
and UO_1484 (O_1484,N_14671,N_14874);
and UO_1485 (O_1485,N_14979,N_14273);
and UO_1486 (O_1486,N_14579,N_14914);
xnor UO_1487 (O_1487,N_14629,N_14498);
nor UO_1488 (O_1488,N_14442,N_14712);
nor UO_1489 (O_1489,N_14577,N_14672);
nor UO_1490 (O_1490,N_14853,N_14954);
xnor UO_1491 (O_1491,N_14685,N_14546);
nand UO_1492 (O_1492,N_14981,N_14486);
xor UO_1493 (O_1493,N_14494,N_14566);
nand UO_1494 (O_1494,N_14653,N_14290);
nand UO_1495 (O_1495,N_14522,N_14928);
or UO_1496 (O_1496,N_14993,N_14460);
nand UO_1497 (O_1497,N_14775,N_14867);
and UO_1498 (O_1498,N_14592,N_14519);
or UO_1499 (O_1499,N_14521,N_14632);
or UO_1500 (O_1500,N_14881,N_14682);
nor UO_1501 (O_1501,N_14931,N_14781);
nor UO_1502 (O_1502,N_14784,N_14426);
or UO_1503 (O_1503,N_14444,N_14314);
nor UO_1504 (O_1504,N_14642,N_14664);
nor UO_1505 (O_1505,N_14400,N_14662);
nor UO_1506 (O_1506,N_14447,N_14292);
nor UO_1507 (O_1507,N_14275,N_14289);
nand UO_1508 (O_1508,N_14893,N_14689);
nor UO_1509 (O_1509,N_14688,N_14756);
or UO_1510 (O_1510,N_14968,N_14727);
and UO_1511 (O_1511,N_14324,N_14971);
nand UO_1512 (O_1512,N_14906,N_14593);
nand UO_1513 (O_1513,N_14982,N_14579);
nand UO_1514 (O_1514,N_14931,N_14684);
nand UO_1515 (O_1515,N_14269,N_14673);
and UO_1516 (O_1516,N_14519,N_14700);
nand UO_1517 (O_1517,N_14983,N_14680);
nand UO_1518 (O_1518,N_14768,N_14847);
or UO_1519 (O_1519,N_14895,N_14603);
or UO_1520 (O_1520,N_14339,N_14657);
or UO_1521 (O_1521,N_14481,N_14290);
nand UO_1522 (O_1522,N_14889,N_14996);
or UO_1523 (O_1523,N_14311,N_14490);
nand UO_1524 (O_1524,N_14374,N_14722);
xor UO_1525 (O_1525,N_14601,N_14426);
or UO_1526 (O_1526,N_14413,N_14269);
and UO_1527 (O_1527,N_14351,N_14613);
or UO_1528 (O_1528,N_14781,N_14611);
and UO_1529 (O_1529,N_14766,N_14781);
nand UO_1530 (O_1530,N_14255,N_14700);
xnor UO_1531 (O_1531,N_14683,N_14960);
and UO_1532 (O_1532,N_14299,N_14458);
nand UO_1533 (O_1533,N_14557,N_14462);
and UO_1534 (O_1534,N_14385,N_14655);
nor UO_1535 (O_1535,N_14537,N_14573);
nor UO_1536 (O_1536,N_14620,N_14257);
or UO_1537 (O_1537,N_14253,N_14949);
or UO_1538 (O_1538,N_14524,N_14750);
xnor UO_1539 (O_1539,N_14430,N_14952);
and UO_1540 (O_1540,N_14728,N_14916);
xor UO_1541 (O_1541,N_14524,N_14292);
and UO_1542 (O_1542,N_14532,N_14903);
or UO_1543 (O_1543,N_14323,N_14685);
or UO_1544 (O_1544,N_14598,N_14706);
nand UO_1545 (O_1545,N_14556,N_14769);
or UO_1546 (O_1546,N_14514,N_14671);
or UO_1547 (O_1547,N_14659,N_14652);
or UO_1548 (O_1548,N_14894,N_14781);
nand UO_1549 (O_1549,N_14665,N_14637);
nor UO_1550 (O_1550,N_14920,N_14720);
or UO_1551 (O_1551,N_14463,N_14483);
nor UO_1552 (O_1552,N_14880,N_14832);
nand UO_1553 (O_1553,N_14304,N_14761);
nor UO_1554 (O_1554,N_14919,N_14548);
nand UO_1555 (O_1555,N_14540,N_14260);
and UO_1556 (O_1556,N_14439,N_14657);
nor UO_1557 (O_1557,N_14952,N_14905);
xnor UO_1558 (O_1558,N_14288,N_14334);
nand UO_1559 (O_1559,N_14939,N_14993);
or UO_1560 (O_1560,N_14908,N_14984);
or UO_1561 (O_1561,N_14454,N_14507);
or UO_1562 (O_1562,N_14835,N_14986);
and UO_1563 (O_1563,N_14870,N_14306);
nand UO_1564 (O_1564,N_14350,N_14604);
nor UO_1565 (O_1565,N_14309,N_14454);
nand UO_1566 (O_1566,N_14617,N_14544);
and UO_1567 (O_1567,N_14750,N_14421);
nand UO_1568 (O_1568,N_14887,N_14494);
nand UO_1569 (O_1569,N_14354,N_14924);
nand UO_1570 (O_1570,N_14915,N_14730);
nand UO_1571 (O_1571,N_14583,N_14985);
or UO_1572 (O_1572,N_14563,N_14480);
nor UO_1573 (O_1573,N_14918,N_14932);
nand UO_1574 (O_1574,N_14758,N_14322);
and UO_1575 (O_1575,N_14919,N_14363);
nor UO_1576 (O_1576,N_14533,N_14857);
nand UO_1577 (O_1577,N_14337,N_14936);
or UO_1578 (O_1578,N_14339,N_14627);
nand UO_1579 (O_1579,N_14910,N_14846);
xnor UO_1580 (O_1580,N_14656,N_14854);
and UO_1581 (O_1581,N_14256,N_14623);
nor UO_1582 (O_1582,N_14994,N_14421);
nor UO_1583 (O_1583,N_14332,N_14597);
nor UO_1584 (O_1584,N_14884,N_14410);
nor UO_1585 (O_1585,N_14845,N_14281);
and UO_1586 (O_1586,N_14445,N_14446);
xnor UO_1587 (O_1587,N_14501,N_14872);
nand UO_1588 (O_1588,N_14401,N_14893);
or UO_1589 (O_1589,N_14542,N_14807);
or UO_1590 (O_1590,N_14957,N_14468);
or UO_1591 (O_1591,N_14991,N_14732);
or UO_1592 (O_1592,N_14963,N_14855);
xnor UO_1593 (O_1593,N_14358,N_14678);
nor UO_1594 (O_1594,N_14790,N_14756);
or UO_1595 (O_1595,N_14448,N_14603);
xor UO_1596 (O_1596,N_14926,N_14643);
nor UO_1597 (O_1597,N_14267,N_14871);
nand UO_1598 (O_1598,N_14779,N_14354);
and UO_1599 (O_1599,N_14292,N_14580);
nand UO_1600 (O_1600,N_14277,N_14836);
or UO_1601 (O_1601,N_14788,N_14479);
nor UO_1602 (O_1602,N_14970,N_14491);
and UO_1603 (O_1603,N_14406,N_14484);
or UO_1604 (O_1604,N_14472,N_14731);
and UO_1605 (O_1605,N_14915,N_14383);
nor UO_1606 (O_1606,N_14994,N_14655);
and UO_1607 (O_1607,N_14255,N_14728);
nand UO_1608 (O_1608,N_14313,N_14272);
nor UO_1609 (O_1609,N_14619,N_14615);
or UO_1610 (O_1610,N_14557,N_14770);
nand UO_1611 (O_1611,N_14798,N_14284);
or UO_1612 (O_1612,N_14908,N_14682);
nand UO_1613 (O_1613,N_14986,N_14709);
and UO_1614 (O_1614,N_14453,N_14536);
and UO_1615 (O_1615,N_14388,N_14390);
or UO_1616 (O_1616,N_14676,N_14617);
nand UO_1617 (O_1617,N_14328,N_14858);
and UO_1618 (O_1618,N_14704,N_14352);
and UO_1619 (O_1619,N_14652,N_14971);
or UO_1620 (O_1620,N_14641,N_14437);
nand UO_1621 (O_1621,N_14887,N_14647);
nand UO_1622 (O_1622,N_14926,N_14756);
nand UO_1623 (O_1623,N_14908,N_14833);
or UO_1624 (O_1624,N_14743,N_14647);
or UO_1625 (O_1625,N_14916,N_14850);
nand UO_1626 (O_1626,N_14480,N_14896);
or UO_1627 (O_1627,N_14967,N_14763);
or UO_1628 (O_1628,N_14762,N_14958);
nand UO_1629 (O_1629,N_14702,N_14921);
nor UO_1630 (O_1630,N_14379,N_14609);
nand UO_1631 (O_1631,N_14894,N_14480);
nor UO_1632 (O_1632,N_14970,N_14633);
and UO_1633 (O_1633,N_14719,N_14259);
xnor UO_1634 (O_1634,N_14584,N_14524);
and UO_1635 (O_1635,N_14966,N_14575);
and UO_1636 (O_1636,N_14691,N_14258);
nor UO_1637 (O_1637,N_14659,N_14461);
nor UO_1638 (O_1638,N_14471,N_14677);
and UO_1639 (O_1639,N_14649,N_14417);
xor UO_1640 (O_1640,N_14870,N_14924);
xnor UO_1641 (O_1641,N_14618,N_14633);
nor UO_1642 (O_1642,N_14529,N_14801);
or UO_1643 (O_1643,N_14547,N_14373);
or UO_1644 (O_1644,N_14496,N_14447);
nor UO_1645 (O_1645,N_14453,N_14427);
and UO_1646 (O_1646,N_14386,N_14289);
nor UO_1647 (O_1647,N_14772,N_14665);
and UO_1648 (O_1648,N_14653,N_14645);
nand UO_1649 (O_1649,N_14631,N_14512);
and UO_1650 (O_1650,N_14391,N_14681);
nand UO_1651 (O_1651,N_14397,N_14579);
nor UO_1652 (O_1652,N_14264,N_14270);
or UO_1653 (O_1653,N_14491,N_14972);
and UO_1654 (O_1654,N_14321,N_14475);
xnor UO_1655 (O_1655,N_14327,N_14742);
and UO_1656 (O_1656,N_14453,N_14785);
or UO_1657 (O_1657,N_14706,N_14423);
and UO_1658 (O_1658,N_14985,N_14791);
and UO_1659 (O_1659,N_14510,N_14596);
or UO_1660 (O_1660,N_14733,N_14353);
and UO_1661 (O_1661,N_14723,N_14754);
or UO_1662 (O_1662,N_14498,N_14403);
nor UO_1663 (O_1663,N_14392,N_14519);
nand UO_1664 (O_1664,N_14419,N_14820);
xor UO_1665 (O_1665,N_14277,N_14970);
and UO_1666 (O_1666,N_14295,N_14584);
or UO_1667 (O_1667,N_14514,N_14716);
nand UO_1668 (O_1668,N_14916,N_14843);
nor UO_1669 (O_1669,N_14619,N_14956);
or UO_1670 (O_1670,N_14754,N_14900);
nor UO_1671 (O_1671,N_14385,N_14803);
nand UO_1672 (O_1672,N_14564,N_14939);
nand UO_1673 (O_1673,N_14880,N_14693);
nand UO_1674 (O_1674,N_14303,N_14335);
nor UO_1675 (O_1675,N_14314,N_14665);
nor UO_1676 (O_1676,N_14257,N_14508);
nand UO_1677 (O_1677,N_14346,N_14904);
or UO_1678 (O_1678,N_14921,N_14436);
and UO_1679 (O_1679,N_14949,N_14424);
or UO_1680 (O_1680,N_14365,N_14504);
nor UO_1681 (O_1681,N_14798,N_14374);
nand UO_1682 (O_1682,N_14423,N_14616);
and UO_1683 (O_1683,N_14776,N_14631);
nor UO_1684 (O_1684,N_14334,N_14707);
and UO_1685 (O_1685,N_14491,N_14688);
nand UO_1686 (O_1686,N_14895,N_14877);
xor UO_1687 (O_1687,N_14701,N_14796);
xor UO_1688 (O_1688,N_14402,N_14507);
or UO_1689 (O_1689,N_14550,N_14692);
nand UO_1690 (O_1690,N_14373,N_14979);
or UO_1691 (O_1691,N_14953,N_14672);
nor UO_1692 (O_1692,N_14282,N_14276);
nor UO_1693 (O_1693,N_14477,N_14635);
nand UO_1694 (O_1694,N_14685,N_14332);
and UO_1695 (O_1695,N_14795,N_14912);
or UO_1696 (O_1696,N_14686,N_14835);
nand UO_1697 (O_1697,N_14705,N_14771);
xor UO_1698 (O_1698,N_14311,N_14786);
or UO_1699 (O_1699,N_14635,N_14279);
or UO_1700 (O_1700,N_14622,N_14491);
nand UO_1701 (O_1701,N_14892,N_14359);
nor UO_1702 (O_1702,N_14848,N_14415);
or UO_1703 (O_1703,N_14544,N_14293);
nor UO_1704 (O_1704,N_14989,N_14688);
nor UO_1705 (O_1705,N_14421,N_14829);
nand UO_1706 (O_1706,N_14578,N_14326);
or UO_1707 (O_1707,N_14449,N_14365);
or UO_1708 (O_1708,N_14546,N_14791);
nor UO_1709 (O_1709,N_14879,N_14585);
nor UO_1710 (O_1710,N_14261,N_14315);
and UO_1711 (O_1711,N_14417,N_14298);
xor UO_1712 (O_1712,N_14343,N_14490);
nor UO_1713 (O_1713,N_14580,N_14258);
nand UO_1714 (O_1714,N_14340,N_14345);
nor UO_1715 (O_1715,N_14548,N_14530);
or UO_1716 (O_1716,N_14419,N_14310);
nor UO_1717 (O_1717,N_14825,N_14819);
nor UO_1718 (O_1718,N_14293,N_14867);
nand UO_1719 (O_1719,N_14330,N_14310);
and UO_1720 (O_1720,N_14889,N_14520);
or UO_1721 (O_1721,N_14605,N_14784);
or UO_1722 (O_1722,N_14584,N_14899);
or UO_1723 (O_1723,N_14776,N_14806);
nor UO_1724 (O_1724,N_14960,N_14419);
or UO_1725 (O_1725,N_14762,N_14702);
or UO_1726 (O_1726,N_14843,N_14654);
and UO_1727 (O_1727,N_14383,N_14505);
and UO_1728 (O_1728,N_14346,N_14450);
or UO_1729 (O_1729,N_14880,N_14604);
or UO_1730 (O_1730,N_14963,N_14885);
or UO_1731 (O_1731,N_14471,N_14922);
and UO_1732 (O_1732,N_14835,N_14864);
and UO_1733 (O_1733,N_14743,N_14940);
nor UO_1734 (O_1734,N_14937,N_14346);
xor UO_1735 (O_1735,N_14666,N_14367);
or UO_1736 (O_1736,N_14907,N_14382);
nor UO_1737 (O_1737,N_14305,N_14952);
xor UO_1738 (O_1738,N_14259,N_14971);
nand UO_1739 (O_1739,N_14424,N_14940);
nand UO_1740 (O_1740,N_14845,N_14559);
nand UO_1741 (O_1741,N_14705,N_14303);
nand UO_1742 (O_1742,N_14807,N_14898);
or UO_1743 (O_1743,N_14378,N_14694);
nand UO_1744 (O_1744,N_14482,N_14643);
xnor UO_1745 (O_1745,N_14505,N_14419);
xor UO_1746 (O_1746,N_14493,N_14562);
nand UO_1747 (O_1747,N_14829,N_14361);
or UO_1748 (O_1748,N_14764,N_14495);
nand UO_1749 (O_1749,N_14782,N_14541);
or UO_1750 (O_1750,N_14290,N_14457);
nor UO_1751 (O_1751,N_14594,N_14516);
or UO_1752 (O_1752,N_14267,N_14482);
nor UO_1753 (O_1753,N_14599,N_14390);
and UO_1754 (O_1754,N_14834,N_14457);
nor UO_1755 (O_1755,N_14738,N_14383);
and UO_1756 (O_1756,N_14964,N_14275);
nand UO_1757 (O_1757,N_14368,N_14855);
nand UO_1758 (O_1758,N_14485,N_14591);
or UO_1759 (O_1759,N_14616,N_14758);
and UO_1760 (O_1760,N_14392,N_14741);
and UO_1761 (O_1761,N_14265,N_14893);
or UO_1762 (O_1762,N_14418,N_14548);
nor UO_1763 (O_1763,N_14832,N_14305);
nand UO_1764 (O_1764,N_14885,N_14416);
or UO_1765 (O_1765,N_14809,N_14815);
nor UO_1766 (O_1766,N_14393,N_14300);
nand UO_1767 (O_1767,N_14434,N_14641);
and UO_1768 (O_1768,N_14641,N_14862);
and UO_1769 (O_1769,N_14991,N_14777);
or UO_1770 (O_1770,N_14738,N_14330);
or UO_1771 (O_1771,N_14992,N_14794);
or UO_1772 (O_1772,N_14383,N_14885);
or UO_1773 (O_1773,N_14773,N_14902);
and UO_1774 (O_1774,N_14558,N_14308);
nand UO_1775 (O_1775,N_14736,N_14784);
nand UO_1776 (O_1776,N_14571,N_14281);
and UO_1777 (O_1777,N_14651,N_14920);
nand UO_1778 (O_1778,N_14960,N_14912);
and UO_1779 (O_1779,N_14895,N_14947);
xor UO_1780 (O_1780,N_14613,N_14602);
xor UO_1781 (O_1781,N_14910,N_14351);
and UO_1782 (O_1782,N_14340,N_14298);
or UO_1783 (O_1783,N_14873,N_14663);
and UO_1784 (O_1784,N_14949,N_14369);
or UO_1785 (O_1785,N_14612,N_14727);
or UO_1786 (O_1786,N_14956,N_14639);
nor UO_1787 (O_1787,N_14932,N_14285);
nand UO_1788 (O_1788,N_14605,N_14468);
nor UO_1789 (O_1789,N_14655,N_14496);
nor UO_1790 (O_1790,N_14993,N_14846);
xnor UO_1791 (O_1791,N_14348,N_14842);
and UO_1792 (O_1792,N_14592,N_14697);
and UO_1793 (O_1793,N_14902,N_14507);
or UO_1794 (O_1794,N_14984,N_14613);
nor UO_1795 (O_1795,N_14503,N_14814);
and UO_1796 (O_1796,N_14401,N_14416);
nor UO_1797 (O_1797,N_14283,N_14312);
nor UO_1798 (O_1798,N_14777,N_14302);
nor UO_1799 (O_1799,N_14296,N_14692);
and UO_1800 (O_1800,N_14509,N_14826);
and UO_1801 (O_1801,N_14403,N_14678);
xnor UO_1802 (O_1802,N_14541,N_14486);
and UO_1803 (O_1803,N_14991,N_14344);
or UO_1804 (O_1804,N_14702,N_14763);
or UO_1805 (O_1805,N_14614,N_14535);
or UO_1806 (O_1806,N_14775,N_14997);
xnor UO_1807 (O_1807,N_14429,N_14670);
or UO_1808 (O_1808,N_14772,N_14438);
nand UO_1809 (O_1809,N_14394,N_14324);
and UO_1810 (O_1810,N_14440,N_14330);
nor UO_1811 (O_1811,N_14765,N_14413);
nor UO_1812 (O_1812,N_14842,N_14582);
or UO_1813 (O_1813,N_14691,N_14968);
and UO_1814 (O_1814,N_14272,N_14836);
and UO_1815 (O_1815,N_14819,N_14694);
xor UO_1816 (O_1816,N_14556,N_14311);
nand UO_1817 (O_1817,N_14742,N_14860);
or UO_1818 (O_1818,N_14473,N_14334);
nand UO_1819 (O_1819,N_14374,N_14967);
or UO_1820 (O_1820,N_14409,N_14577);
nor UO_1821 (O_1821,N_14879,N_14670);
and UO_1822 (O_1822,N_14749,N_14267);
or UO_1823 (O_1823,N_14554,N_14540);
nand UO_1824 (O_1824,N_14912,N_14993);
nand UO_1825 (O_1825,N_14278,N_14744);
nor UO_1826 (O_1826,N_14958,N_14869);
or UO_1827 (O_1827,N_14629,N_14519);
nand UO_1828 (O_1828,N_14454,N_14734);
and UO_1829 (O_1829,N_14659,N_14905);
nor UO_1830 (O_1830,N_14969,N_14911);
and UO_1831 (O_1831,N_14713,N_14720);
and UO_1832 (O_1832,N_14268,N_14601);
and UO_1833 (O_1833,N_14965,N_14375);
nand UO_1834 (O_1834,N_14483,N_14389);
nand UO_1835 (O_1835,N_14280,N_14459);
nor UO_1836 (O_1836,N_14260,N_14891);
and UO_1837 (O_1837,N_14539,N_14933);
and UO_1838 (O_1838,N_14798,N_14726);
and UO_1839 (O_1839,N_14292,N_14627);
xor UO_1840 (O_1840,N_14695,N_14479);
nor UO_1841 (O_1841,N_14566,N_14298);
or UO_1842 (O_1842,N_14894,N_14591);
nand UO_1843 (O_1843,N_14916,N_14399);
nand UO_1844 (O_1844,N_14511,N_14409);
xnor UO_1845 (O_1845,N_14438,N_14925);
or UO_1846 (O_1846,N_14472,N_14340);
nor UO_1847 (O_1847,N_14871,N_14572);
or UO_1848 (O_1848,N_14776,N_14434);
and UO_1849 (O_1849,N_14672,N_14304);
or UO_1850 (O_1850,N_14863,N_14848);
nand UO_1851 (O_1851,N_14535,N_14601);
or UO_1852 (O_1852,N_14353,N_14959);
nor UO_1853 (O_1853,N_14280,N_14654);
nor UO_1854 (O_1854,N_14715,N_14489);
nand UO_1855 (O_1855,N_14687,N_14596);
nor UO_1856 (O_1856,N_14873,N_14509);
nand UO_1857 (O_1857,N_14852,N_14511);
nor UO_1858 (O_1858,N_14597,N_14460);
or UO_1859 (O_1859,N_14837,N_14909);
nor UO_1860 (O_1860,N_14961,N_14692);
or UO_1861 (O_1861,N_14510,N_14313);
or UO_1862 (O_1862,N_14618,N_14646);
nand UO_1863 (O_1863,N_14387,N_14954);
nand UO_1864 (O_1864,N_14645,N_14789);
nand UO_1865 (O_1865,N_14364,N_14735);
nand UO_1866 (O_1866,N_14744,N_14444);
nand UO_1867 (O_1867,N_14537,N_14447);
nor UO_1868 (O_1868,N_14810,N_14608);
xor UO_1869 (O_1869,N_14716,N_14728);
or UO_1870 (O_1870,N_14882,N_14796);
or UO_1871 (O_1871,N_14647,N_14717);
nor UO_1872 (O_1872,N_14940,N_14294);
xnor UO_1873 (O_1873,N_14761,N_14986);
and UO_1874 (O_1874,N_14674,N_14768);
xor UO_1875 (O_1875,N_14322,N_14413);
or UO_1876 (O_1876,N_14664,N_14926);
and UO_1877 (O_1877,N_14688,N_14857);
or UO_1878 (O_1878,N_14587,N_14551);
nand UO_1879 (O_1879,N_14891,N_14777);
and UO_1880 (O_1880,N_14285,N_14271);
nand UO_1881 (O_1881,N_14317,N_14517);
nand UO_1882 (O_1882,N_14922,N_14404);
nand UO_1883 (O_1883,N_14450,N_14978);
xor UO_1884 (O_1884,N_14801,N_14541);
nand UO_1885 (O_1885,N_14724,N_14829);
or UO_1886 (O_1886,N_14431,N_14304);
or UO_1887 (O_1887,N_14654,N_14591);
and UO_1888 (O_1888,N_14608,N_14495);
and UO_1889 (O_1889,N_14303,N_14910);
nor UO_1890 (O_1890,N_14659,N_14520);
nand UO_1891 (O_1891,N_14732,N_14454);
xor UO_1892 (O_1892,N_14503,N_14429);
and UO_1893 (O_1893,N_14257,N_14711);
nand UO_1894 (O_1894,N_14824,N_14399);
or UO_1895 (O_1895,N_14266,N_14513);
xor UO_1896 (O_1896,N_14766,N_14294);
or UO_1897 (O_1897,N_14873,N_14917);
and UO_1898 (O_1898,N_14922,N_14840);
nor UO_1899 (O_1899,N_14502,N_14349);
nand UO_1900 (O_1900,N_14656,N_14551);
nand UO_1901 (O_1901,N_14323,N_14597);
xor UO_1902 (O_1902,N_14776,N_14976);
nand UO_1903 (O_1903,N_14555,N_14363);
and UO_1904 (O_1904,N_14710,N_14589);
nor UO_1905 (O_1905,N_14862,N_14955);
nor UO_1906 (O_1906,N_14781,N_14658);
nand UO_1907 (O_1907,N_14274,N_14451);
or UO_1908 (O_1908,N_14951,N_14258);
xor UO_1909 (O_1909,N_14342,N_14601);
nor UO_1910 (O_1910,N_14987,N_14378);
nor UO_1911 (O_1911,N_14489,N_14984);
and UO_1912 (O_1912,N_14607,N_14446);
and UO_1913 (O_1913,N_14744,N_14823);
or UO_1914 (O_1914,N_14678,N_14527);
nand UO_1915 (O_1915,N_14498,N_14624);
nor UO_1916 (O_1916,N_14767,N_14352);
or UO_1917 (O_1917,N_14399,N_14695);
or UO_1918 (O_1918,N_14429,N_14533);
and UO_1919 (O_1919,N_14670,N_14350);
or UO_1920 (O_1920,N_14561,N_14848);
and UO_1921 (O_1921,N_14572,N_14821);
or UO_1922 (O_1922,N_14597,N_14962);
or UO_1923 (O_1923,N_14524,N_14415);
or UO_1924 (O_1924,N_14962,N_14510);
and UO_1925 (O_1925,N_14430,N_14559);
and UO_1926 (O_1926,N_14796,N_14731);
nand UO_1927 (O_1927,N_14780,N_14962);
nor UO_1928 (O_1928,N_14378,N_14862);
nor UO_1929 (O_1929,N_14412,N_14282);
and UO_1930 (O_1930,N_14496,N_14568);
or UO_1931 (O_1931,N_14742,N_14625);
nand UO_1932 (O_1932,N_14556,N_14722);
nand UO_1933 (O_1933,N_14445,N_14269);
and UO_1934 (O_1934,N_14893,N_14822);
and UO_1935 (O_1935,N_14572,N_14540);
and UO_1936 (O_1936,N_14664,N_14813);
nor UO_1937 (O_1937,N_14774,N_14491);
nand UO_1938 (O_1938,N_14739,N_14664);
nand UO_1939 (O_1939,N_14756,N_14902);
nand UO_1940 (O_1940,N_14698,N_14705);
xor UO_1941 (O_1941,N_14972,N_14814);
or UO_1942 (O_1942,N_14508,N_14265);
or UO_1943 (O_1943,N_14454,N_14463);
nor UO_1944 (O_1944,N_14468,N_14517);
nor UO_1945 (O_1945,N_14530,N_14372);
nand UO_1946 (O_1946,N_14991,N_14696);
or UO_1947 (O_1947,N_14371,N_14768);
or UO_1948 (O_1948,N_14474,N_14303);
nand UO_1949 (O_1949,N_14562,N_14350);
or UO_1950 (O_1950,N_14617,N_14439);
and UO_1951 (O_1951,N_14374,N_14667);
nor UO_1952 (O_1952,N_14322,N_14271);
nand UO_1953 (O_1953,N_14848,N_14619);
and UO_1954 (O_1954,N_14350,N_14281);
and UO_1955 (O_1955,N_14500,N_14595);
or UO_1956 (O_1956,N_14937,N_14262);
and UO_1957 (O_1957,N_14853,N_14532);
nor UO_1958 (O_1958,N_14342,N_14709);
and UO_1959 (O_1959,N_14767,N_14863);
nand UO_1960 (O_1960,N_14792,N_14559);
and UO_1961 (O_1961,N_14924,N_14603);
nor UO_1962 (O_1962,N_14285,N_14593);
xor UO_1963 (O_1963,N_14781,N_14629);
or UO_1964 (O_1964,N_14813,N_14963);
nand UO_1965 (O_1965,N_14376,N_14595);
or UO_1966 (O_1966,N_14442,N_14784);
or UO_1967 (O_1967,N_14626,N_14505);
nor UO_1968 (O_1968,N_14326,N_14737);
and UO_1969 (O_1969,N_14692,N_14355);
and UO_1970 (O_1970,N_14423,N_14321);
and UO_1971 (O_1971,N_14723,N_14388);
nor UO_1972 (O_1972,N_14343,N_14405);
or UO_1973 (O_1973,N_14598,N_14377);
and UO_1974 (O_1974,N_14791,N_14316);
or UO_1975 (O_1975,N_14336,N_14649);
or UO_1976 (O_1976,N_14315,N_14846);
xor UO_1977 (O_1977,N_14869,N_14402);
or UO_1978 (O_1978,N_14295,N_14880);
nor UO_1979 (O_1979,N_14896,N_14571);
and UO_1980 (O_1980,N_14880,N_14313);
or UO_1981 (O_1981,N_14874,N_14600);
nor UO_1982 (O_1982,N_14409,N_14618);
or UO_1983 (O_1983,N_14316,N_14327);
or UO_1984 (O_1984,N_14269,N_14964);
and UO_1985 (O_1985,N_14371,N_14765);
nand UO_1986 (O_1986,N_14322,N_14919);
nor UO_1987 (O_1987,N_14953,N_14366);
or UO_1988 (O_1988,N_14655,N_14273);
nor UO_1989 (O_1989,N_14439,N_14278);
or UO_1990 (O_1990,N_14477,N_14929);
and UO_1991 (O_1991,N_14678,N_14436);
nor UO_1992 (O_1992,N_14736,N_14397);
nand UO_1993 (O_1993,N_14536,N_14838);
or UO_1994 (O_1994,N_14636,N_14716);
or UO_1995 (O_1995,N_14595,N_14279);
or UO_1996 (O_1996,N_14993,N_14883);
or UO_1997 (O_1997,N_14730,N_14457);
and UO_1998 (O_1998,N_14884,N_14649);
nand UO_1999 (O_1999,N_14259,N_14587);
endmodule