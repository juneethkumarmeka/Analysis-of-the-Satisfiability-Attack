module basic_1000_10000_1500_2_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5001,N_5004,N_5005,N_5006,N_5008,N_5009,N_5010,N_5014,N_5015,N_5016,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5026,N_5028,N_5029,N_5033,N_5034,N_5036,N_5037,N_5039,N_5041,N_5042,N_5043,N_5044,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5057,N_5059,N_5060,N_5061,N_5063,N_5067,N_5068,N_5070,N_5073,N_5075,N_5076,N_5078,N_5079,N_5080,N_5081,N_5084,N_5085,N_5088,N_5089,N_5093,N_5094,N_5095,N_5098,N_5099,N_5101,N_5102,N_5103,N_5105,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5123,N_5124,N_5125,N_5126,N_5128,N_5129,N_5130,N_5131,N_5133,N_5134,N_5136,N_5137,N_5140,N_5141,N_5143,N_5144,N_5146,N_5147,N_5152,N_5154,N_5155,N_5157,N_5161,N_5162,N_5165,N_5166,N_5167,N_5169,N_5171,N_5172,N_5174,N_5175,N_5176,N_5178,N_5180,N_5181,N_5183,N_5184,N_5186,N_5187,N_5189,N_5190,N_5191,N_5192,N_5195,N_5196,N_5198,N_5200,N_5201,N_5202,N_5203,N_5204,N_5206,N_5211,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5222,N_5226,N_5227,N_5230,N_5232,N_5233,N_5235,N_5239,N_5242,N_5244,N_5245,N_5246,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5259,N_5260,N_5262,N_5264,N_5265,N_5267,N_5268,N_5269,N_5270,N_5272,N_5274,N_5276,N_5277,N_5281,N_5282,N_5283,N_5285,N_5289,N_5293,N_5294,N_5295,N_5299,N_5300,N_5305,N_5307,N_5308,N_5309,N_5310,N_5311,N_5313,N_5314,N_5316,N_5317,N_5319,N_5320,N_5321,N_5322,N_5323,N_5326,N_5328,N_5329,N_5330,N_5332,N_5333,N_5334,N_5335,N_5336,N_5342,N_5343,N_5344,N_5346,N_5347,N_5349,N_5352,N_5353,N_5357,N_5359,N_5360,N_5361,N_5363,N_5364,N_5365,N_5366,N_5367,N_5369,N_5370,N_5371,N_5373,N_5375,N_5376,N_5379,N_5380,N_5381,N_5382,N_5384,N_5385,N_5388,N_5395,N_5396,N_5397,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5413,N_5414,N_5417,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5429,N_5430,N_5431,N_5432,N_5433,N_5436,N_5437,N_5439,N_5440,N_5441,N_5442,N_5444,N_5446,N_5447,N_5448,N_5449,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5459,N_5461,N_5464,N_5465,N_5467,N_5468,N_5470,N_5472,N_5474,N_5475,N_5476,N_5479,N_5480,N_5481,N_5484,N_5487,N_5488,N_5490,N_5491,N_5492,N_5493,N_5494,N_5497,N_5498,N_5499,N_5501,N_5504,N_5506,N_5508,N_5509,N_5512,N_5513,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5523,N_5524,N_5529,N_5530,N_5531,N_5532,N_5533,N_5536,N_5537,N_5538,N_5539,N_5544,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5559,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5570,N_5573,N_5574,N_5576,N_5577,N_5578,N_5581,N_5582,N_5583,N_5584,N_5585,N_5587,N_5589,N_5591,N_5592,N_5593,N_5594,N_5597,N_5598,N_5599,N_5600,N_5602,N_5603,N_5604,N_5606,N_5608,N_5609,N_5612,N_5613,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5627,N_5629,N_5630,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5646,N_5647,N_5650,N_5651,N_5652,N_5653,N_5654,N_5656,N_5658,N_5659,N_5661,N_5662,N_5663,N_5667,N_5668,N_5669,N_5671,N_5673,N_5675,N_5677,N_5678,N_5682,N_5684,N_5686,N_5687,N_5688,N_5691,N_5692,N_5694,N_5696,N_5697,N_5699,N_5700,N_5701,N_5703,N_5704,N_5705,N_5706,N_5709,N_5711,N_5712,N_5715,N_5719,N_5722,N_5723,N_5728,N_5729,N_5730,N_5732,N_5733,N_5734,N_5735,N_5737,N_5739,N_5741,N_5742,N_5743,N_5748,N_5749,N_5750,N_5751,N_5752,N_5755,N_5758,N_5759,N_5762,N_5764,N_5765,N_5767,N_5768,N_5769,N_5771,N_5772,N_5774,N_5778,N_5779,N_5781,N_5783,N_5786,N_5787,N_5789,N_5790,N_5792,N_5793,N_5795,N_5796,N_5798,N_5799,N_5801,N_5802,N_5804,N_5805,N_5808,N_5811,N_5813,N_5815,N_5816,N_5817,N_5818,N_5820,N_5821,N_5823,N_5826,N_5828,N_5833,N_5834,N_5835,N_5836,N_5840,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5858,N_5859,N_5862,N_5865,N_5866,N_5869,N_5871,N_5872,N_5875,N_5876,N_5877,N_5878,N_5880,N_5883,N_5885,N_5886,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5895,N_5896,N_5898,N_5899,N_5902,N_5903,N_5906,N_5908,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5922,N_5923,N_5924,N_5925,N_5926,N_5928,N_5929,N_5930,N_5931,N_5933,N_5934,N_5938,N_5939,N_5944,N_5945,N_5946,N_5948,N_5950,N_5951,N_5953,N_5954,N_5956,N_5957,N_5960,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5980,N_5981,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5992,N_5993,N_5995,N_5996,N_5998,N_5999,N_6002,N_6005,N_6006,N_6008,N_6009,N_6010,N_6012,N_6015,N_6019,N_6020,N_6021,N_6022,N_6023,N_6025,N_6026,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6039,N_6040,N_6041,N_6042,N_6044,N_6045,N_6046,N_6047,N_6048,N_6052,N_6054,N_6056,N_6057,N_6058,N_6061,N_6062,N_6064,N_6065,N_6066,N_6068,N_6072,N_6080,N_6081,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6092,N_6094,N_6095,N_6096,N_6097,N_6099,N_6100,N_6101,N_6102,N_6106,N_6110,N_6111,N_6112,N_6114,N_6115,N_6117,N_6118,N_6119,N_6120,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6129,N_6132,N_6136,N_6137,N_6142,N_6143,N_6145,N_6147,N_6148,N_6150,N_6151,N_6152,N_6153,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6163,N_6164,N_6168,N_6169,N_6170,N_6173,N_6174,N_6175,N_6176,N_6177,N_6182,N_6183,N_6184,N_6185,N_6186,N_6188,N_6190,N_6191,N_6192,N_6193,N_6198,N_6201,N_6202,N_6204,N_6205,N_6206,N_6208,N_6209,N_6213,N_6214,N_6217,N_6219,N_6220,N_6222,N_6223,N_6224,N_6225,N_6230,N_6232,N_6233,N_6234,N_6238,N_6242,N_6243,N_6244,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6255,N_6261,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6272,N_6276,N_6281,N_6282,N_6285,N_6286,N_6288,N_6289,N_6293,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6305,N_6306,N_6308,N_6311,N_6312,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6325,N_6326,N_6327,N_6330,N_6331,N_6332,N_6333,N_6335,N_6337,N_6338,N_6341,N_6342,N_6346,N_6350,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6361,N_6362,N_6363,N_6365,N_6366,N_6367,N_6371,N_6372,N_6375,N_6376,N_6377,N_6380,N_6381,N_6382,N_6383,N_6384,N_6389,N_6392,N_6393,N_6395,N_6396,N_6397,N_6398,N_6400,N_6402,N_6404,N_6407,N_6409,N_6410,N_6411,N_6412,N_6414,N_6415,N_6416,N_6417,N_6419,N_6420,N_6421,N_6423,N_6425,N_6428,N_6429,N_6430,N_6431,N_6433,N_6434,N_6436,N_6438,N_6442,N_6444,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6459,N_6460,N_6462,N_6463,N_6466,N_6468,N_6471,N_6472,N_6473,N_6475,N_6477,N_6478,N_6479,N_6481,N_6482,N_6484,N_6485,N_6487,N_6489,N_6490,N_6492,N_6496,N_6498,N_6500,N_6501,N_6502,N_6503,N_6505,N_6507,N_6508,N_6511,N_6512,N_6513,N_6514,N_6515,N_6517,N_6518,N_6520,N_6521,N_6529,N_6530,N_6531,N_6532,N_6534,N_6535,N_6536,N_6537,N_6539,N_6540,N_6542,N_6543,N_6547,N_6548,N_6549,N_6551,N_6557,N_6558,N_6559,N_6562,N_6563,N_6565,N_6567,N_6568,N_6569,N_6570,N_6571,N_6573,N_6575,N_6576,N_6579,N_6581,N_6584,N_6589,N_6590,N_6591,N_6596,N_6597,N_6598,N_6599,N_6600,N_6603,N_6604,N_6606,N_6608,N_6612,N_6613,N_6614,N_6616,N_6619,N_6623,N_6624,N_6625,N_6626,N_6627,N_6630,N_6631,N_6633,N_6635,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6644,N_6645,N_6646,N_6649,N_6650,N_6653,N_6654,N_6656,N_6657,N_6658,N_6659,N_6660,N_6663,N_6665,N_6666,N_6670,N_6671,N_6672,N_6673,N_6675,N_6678,N_6680,N_6681,N_6683,N_6684,N_6686,N_6687,N_6688,N_6690,N_6691,N_6692,N_6694,N_6695,N_6700,N_6702,N_6704,N_6708,N_6709,N_6711,N_6715,N_6716,N_6717,N_6718,N_6721,N_6722,N_6723,N_6724,N_6726,N_6728,N_6729,N_6731,N_6732,N_6733,N_6741,N_6743,N_6744,N_6745,N_6750,N_6751,N_6753,N_6755,N_6756,N_6757,N_6760,N_6762,N_6763,N_6767,N_6769,N_6771,N_6772,N_6774,N_6775,N_6776,N_6777,N_6779,N_6780,N_6783,N_6784,N_6785,N_6788,N_6790,N_6791,N_6792,N_6797,N_6798,N_6800,N_6802,N_6803,N_6805,N_6806,N_6808,N_6811,N_6812,N_6813,N_6814,N_6815,N_6817,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6828,N_6829,N_6830,N_6831,N_6832,N_6834,N_6835,N_6836,N_6839,N_6840,N_6841,N_6842,N_6845,N_6847,N_6848,N_6850,N_6851,N_6852,N_6853,N_6854,N_6856,N_6857,N_6861,N_6862,N_6863,N_6866,N_6867,N_6869,N_6873,N_6874,N_6875,N_6877,N_6878,N_6879,N_6883,N_6885,N_6888,N_6891,N_6892,N_6893,N_6894,N_6896,N_6897,N_6899,N_6900,N_6903,N_6904,N_6908,N_6910,N_6912,N_6913,N_6915,N_6917,N_6921,N_6922,N_6925,N_6927,N_6935,N_6937,N_6940,N_6941,N_6942,N_6943,N_6944,N_6946,N_6947,N_6949,N_6950,N_6953,N_6954,N_6955,N_6956,N_6957,N_6959,N_6960,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6979,N_6980,N_6984,N_6985,N_6986,N_6989,N_6992,N_6996,N_6998,N_6999,N_7000,N_7001,N_7003,N_7006,N_7007,N_7008,N_7010,N_7011,N_7012,N_7014,N_7018,N_7019,N_7020,N_7021,N_7022,N_7024,N_7025,N_7027,N_7028,N_7031,N_7032,N_7033,N_7035,N_7036,N_7037,N_7038,N_7041,N_7042,N_7045,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7068,N_7071,N_7075,N_7076,N_7078,N_7080,N_7081,N_7082,N_7083,N_7085,N_7086,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7098,N_7099,N_7102,N_7106,N_7108,N_7109,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7119,N_7120,N_7121,N_7122,N_7125,N_7126,N_7127,N_7128,N_7132,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7151,N_7153,N_7155,N_7156,N_7158,N_7159,N_7160,N_7164,N_7165,N_7166,N_7167,N_7172,N_7173,N_7176,N_7177,N_7178,N_7179,N_7180,N_7182,N_7183,N_7185,N_7186,N_7188,N_7189,N_7193,N_7194,N_7196,N_7197,N_7199,N_7200,N_7202,N_7203,N_7205,N_7206,N_7211,N_7213,N_7215,N_7216,N_7219,N_7221,N_7225,N_7226,N_7227,N_7228,N_7229,N_7231,N_7232,N_7233,N_7234,N_7236,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7246,N_7248,N_7249,N_7251,N_7252,N_7253,N_7254,N_7255,N_7260,N_7261,N_7262,N_7264,N_7265,N_7272,N_7273,N_7274,N_7277,N_7279,N_7280,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7291,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7302,N_7306,N_7307,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7324,N_7325,N_7326,N_7327,N_7328,N_7330,N_7332,N_7333,N_7334,N_7335,N_7336,N_7338,N_7339,N_7340,N_7343,N_7344,N_7345,N_7347,N_7348,N_7349,N_7350,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7360,N_7361,N_7363,N_7366,N_7367,N_7368,N_7369,N_7371,N_7373,N_7375,N_7376,N_7378,N_7380,N_7381,N_7384,N_7386,N_7391,N_7392,N_7394,N_7395,N_7396,N_7397,N_7398,N_7400,N_7403,N_7404,N_7405,N_7409,N_7410,N_7411,N_7415,N_7416,N_7419,N_7421,N_7423,N_7424,N_7425,N_7426,N_7428,N_7430,N_7431,N_7432,N_7433,N_7434,N_7437,N_7438,N_7440,N_7443,N_7444,N_7446,N_7447,N_7448,N_7452,N_7453,N_7455,N_7458,N_7459,N_7460,N_7462,N_7463,N_7465,N_7466,N_7467,N_7468,N_7469,N_7472,N_7473,N_7474,N_7475,N_7476,N_7479,N_7480,N_7483,N_7484,N_7487,N_7490,N_7491,N_7493,N_7494,N_7496,N_7497,N_7498,N_7499,N_7502,N_7503,N_7505,N_7506,N_7507,N_7508,N_7510,N_7512,N_7515,N_7516,N_7518,N_7520,N_7521,N_7523,N_7524,N_7526,N_7527,N_7529,N_7530,N_7531,N_7534,N_7535,N_7536,N_7538,N_7539,N_7540,N_7541,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7554,N_7559,N_7560,N_7562,N_7564,N_7565,N_7566,N_7567,N_7569,N_7571,N_7575,N_7576,N_7578,N_7579,N_7580,N_7586,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7596,N_7598,N_7600,N_7601,N_7602,N_7603,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7612,N_7613,N_7615,N_7616,N_7618,N_7620,N_7622,N_7623,N_7624,N_7628,N_7629,N_7632,N_7633,N_7634,N_7637,N_7638,N_7639,N_7640,N_7641,N_7644,N_7647,N_7648,N_7649,N_7652,N_7656,N_7657,N_7658,N_7660,N_7662,N_7663,N_7666,N_7667,N_7668,N_7670,N_7671,N_7673,N_7674,N_7675,N_7676,N_7678,N_7680,N_7682,N_7683,N_7684,N_7685,N_7687,N_7689,N_7690,N_7693,N_7697,N_7699,N_7700,N_7701,N_7702,N_7704,N_7708,N_7710,N_7711,N_7712,N_7714,N_7716,N_7720,N_7722,N_7723,N_7724,N_7725,N_7726,N_7729,N_7730,N_7731,N_7732,N_7734,N_7735,N_7736,N_7737,N_7739,N_7742,N_7746,N_7747,N_7751,N_7752,N_7753,N_7756,N_7757,N_7758,N_7759,N_7761,N_7762,N_7763,N_7764,N_7766,N_7767,N_7769,N_7771,N_7773,N_7774,N_7778,N_7780,N_7781,N_7782,N_7784,N_7788,N_7790,N_7792,N_7793,N_7794,N_7795,N_7796,N_7799,N_7800,N_7801,N_7802,N_7805,N_7806,N_7809,N_7810,N_7813,N_7814,N_7815,N_7816,N_7819,N_7823,N_7825,N_7826,N_7829,N_7831,N_7834,N_7835,N_7838,N_7839,N_7841,N_7843,N_7847,N_7848,N_7849,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7860,N_7863,N_7864,N_7866,N_7870,N_7871,N_7872,N_7874,N_7875,N_7877,N_7879,N_7880,N_7881,N_7883,N_7885,N_7886,N_7887,N_7889,N_7891,N_7892,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7904,N_7906,N_7907,N_7908,N_7909,N_7910,N_7913,N_7915,N_7916,N_7917,N_7918,N_7919,N_7921,N_7923,N_7924,N_7927,N_7929,N_7930,N_7937,N_7942,N_7944,N_7946,N_7947,N_7948,N_7949,N_7955,N_7959,N_7960,N_7961,N_7964,N_7965,N_7967,N_7968,N_7969,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7978,N_7980,N_7982,N_7985,N_7987,N_7988,N_7991,N_7997,N_7998,N_7999,N_8000,N_8001,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8013,N_8014,N_8015,N_8017,N_8018,N_8019,N_8023,N_8024,N_8025,N_8026,N_8027,N_8029,N_8030,N_8031,N_8032,N_8034,N_8035,N_8036,N_8037,N_8039,N_8040,N_8042,N_8043,N_8044,N_8045,N_8046,N_8048,N_8050,N_8054,N_8055,N_8057,N_8058,N_8061,N_8062,N_8065,N_8066,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8078,N_8081,N_8082,N_8085,N_8086,N_8088,N_8089,N_8090,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8104,N_8108,N_8109,N_8110,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8123,N_8124,N_8126,N_8127,N_8128,N_8130,N_8133,N_8134,N_8136,N_8140,N_8141,N_8142,N_8145,N_8147,N_8148,N_8150,N_8154,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8165,N_8166,N_8168,N_8171,N_8172,N_8174,N_8175,N_8176,N_8177,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8196,N_8197,N_8198,N_8199,N_8200,N_8202,N_8204,N_8205,N_8206,N_8207,N_8208,N_8213,N_8217,N_8218,N_8219,N_8220,N_8222,N_8223,N_8224,N_8226,N_8227,N_8229,N_8230,N_8233,N_8235,N_8236,N_8237,N_8238,N_8241,N_8242,N_8244,N_8245,N_8246,N_8248,N_8249,N_8250,N_8252,N_8253,N_8254,N_8261,N_8264,N_8265,N_8269,N_8271,N_8273,N_8274,N_8275,N_8276,N_8277,N_8279,N_8283,N_8284,N_8288,N_8289,N_8290,N_8294,N_8295,N_8296,N_8297,N_8299,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8309,N_8312,N_8315,N_8316,N_8318,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8330,N_8331,N_8333,N_8334,N_8335,N_8336,N_8337,N_8339,N_8340,N_8341,N_8342,N_8343,N_8345,N_8346,N_8348,N_8349,N_8350,N_8352,N_8355,N_8357,N_8358,N_8359,N_8360,N_8362,N_8363,N_8365,N_8366,N_8369,N_8370,N_8373,N_8376,N_8378,N_8380,N_8382,N_8384,N_8386,N_8387,N_8388,N_8391,N_8393,N_8394,N_8395,N_8396,N_8400,N_8401,N_8402,N_8404,N_8406,N_8407,N_8410,N_8413,N_8414,N_8415,N_8416,N_8417,N_8419,N_8420,N_8424,N_8425,N_8428,N_8430,N_8431,N_8432,N_8434,N_8435,N_8436,N_8438,N_8439,N_8442,N_8445,N_8446,N_8447,N_8449,N_8451,N_8452,N_8457,N_8460,N_8461,N_8463,N_8464,N_8467,N_8469,N_8470,N_8471,N_8472,N_8475,N_8476,N_8477,N_8480,N_8481,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8502,N_8503,N_8505,N_8506,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8519,N_8520,N_8521,N_8524,N_8525,N_8527,N_8528,N_8531,N_8533,N_8535,N_8536,N_8537,N_8539,N_8541,N_8543,N_8546,N_8547,N_8549,N_8550,N_8551,N_8553,N_8554,N_8555,N_8560,N_8562,N_8564,N_8567,N_8568,N_8569,N_8570,N_8573,N_8580,N_8582,N_8583,N_8587,N_8588,N_8590,N_8592,N_8593,N_8595,N_8598,N_8601,N_8602,N_8603,N_8606,N_8608,N_8610,N_8611,N_8615,N_8616,N_8619,N_8620,N_8621,N_8622,N_8627,N_8630,N_8632,N_8634,N_8636,N_8637,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8647,N_8648,N_8649,N_8650,N_8653,N_8655,N_8656,N_8660,N_8663,N_8665,N_8666,N_8669,N_8670,N_8671,N_8673,N_8675,N_8676,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8689,N_8692,N_8694,N_8695,N_8696,N_8698,N_8699,N_8700,N_8702,N_8704,N_8705,N_8706,N_8709,N_8710,N_8711,N_8715,N_8719,N_8720,N_8722,N_8723,N_8724,N_8725,N_8727,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8742,N_8743,N_8744,N_8745,N_8747,N_8748,N_8749,N_8753,N_8754,N_8757,N_8759,N_8764,N_8766,N_8767,N_8771,N_8774,N_8777,N_8780,N_8783,N_8785,N_8787,N_8788,N_8792,N_8793,N_8796,N_8797,N_8799,N_8800,N_8802,N_8807,N_8808,N_8814,N_8815,N_8816,N_8817,N_8819,N_8820,N_8822,N_8823,N_8824,N_8825,N_8826,N_8828,N_8829,N_8831,N_8832,N_8836,N_8838,N_8839,N_8841,N_8842,N_8845,N_8846,N_8847,N_8848,N_8850,N_8851,N_8855,N_8857,N_8859,N_8860,N_8862,N_8863,N_8866,N_8867,N_8868,N_8871,N_8873,N_8875,N_8876,N_8878,N_8883,N_8884,N_8885,N_8886,N_8887,N_8889,N_8890,N_8892,N_8893,N_8894,N_8895,N_8897,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8930,N_8932,N_8933,N_8936,N_8937,N_8938,N_8940,N_8941,N_8943,N_8944,N_8945,N_8949,N_8952,N_8953,N_8955,N_8956,N_8957,N_8958,N_8960,N_8962,N_8964,N_8965,N_8967,N_8968,N_8969,N_8971,N_8972,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8999,N_9000,N_9001,N_9004,N_9005,N_9006,N_9008,N_9009,N_9010,N_9013,N_9019,N_9020,N_9021,N_9023,N_9024,N_9025,N_9026,N_9029,N_9031,N_9032,N_9035,N_9036,N_9039,N_9040,N_9041,N_9044,N_9048,N_9050,N_9051,N_9052,N_9054,N_9056,N_9058,N_9060,N_9062,N_9063,N_9066,N_9068,N_9070,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9080,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9098,N_9099,N_9100,N_9101,N_9105,N_9106,N_9107,N_9110,N_9112,N_9113,N_9115,N_9118,N_9120,N_9121,N_9122,N_9123,N_9124,N_9127,N_9128,N_9129,N_9131,N_9132,N_9135,N_9137,N_9138,N_9139,N_9141,N_9144,N_9145,N_9147,N_9149,N_9150,N_9151,N_9152,N_9153,N_9158,N_9159,N_9161,N_9162,N_9163,N_9164,N_9165,N_9167,N_9168,N_9169,N_9170,N_9172,N_9174,N_9175,N_9176,N_9177,N_9178,N_9181,N_9183,N_9185,N_9190,N_9192,N_9195,N_9196,N_9198,N_9199,N_9200,N_9201,N_9203,N_9204,N_9205,N_9207,N_9209,N_9210,N_9211,N_9214,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9241,N_9242,N_9245,N_9247,N_9248,N_9249,N_9251,N_9252,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9262,N_9263,N_9265,N_9267,N_9270,N_9272,N_9273,N_9274,N_9275,N_9276,N_9278,N_9279,N_9280,N_9282,N_9283,N_9284,N_9285,N_9287,N_9289,N_9290,N_9292,N_9296,N_9297,N_9298,N_9299,N_9300,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9319,N_9324,N_9327,N_9330,N_9331,N_9333,N_9334,N_9339,N_9340,N_9341,N_9343,N_9344,N_9345,N_9346,N_9348,N_9354,N_9355,N_9358,N_9360,N_9361,N_9362,N_9364,N_9365,N_9369,N_9371,N_9372,N_9373,N_9374,N_9376,N_9377,N_9379,N_9380,N_9382,N_9383,N_9384,N_9385,N_9387,N_9389,N_9391,N_9392,N_9393,N_9394,N_9397,N_9398,N_9399,N_9400,N_9403,N_9405,N_9407,N_9409,N_9411,N_9412,N_9416,N_9418,N_9421,N_9422,N_9423,N_9424,N_9426,N_9427,N_9429,N_9431,N_9433,N_9434,N_9437,N_9439,N_9440,N_9441,N_9442,N_9443,N_9447,N_9448,N_9450,N_9451,N_9456,N_9457,N_9458,N_9460,N_9461,N_9463,N_9469,N_9471,N_9473,N_9475,N_9478,N_9479,N_9480,N_9482,N_9485,N_9488,N_9489,N_9490,N_9493,N_9494,N_9496,N_9497,N_9498,N_9500,N_9502,N_9503,N_9505,N_9506,N_9507,N_9509,N_9511,N_9513,N_9515,N_9516,N_9517,N_9518,N_9519,N_9521,N_9522,N_9523,N_9525,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9539,N_9540,N_9542,N_9543,N_9544,N_9545,N_9547,N_9548,N_9549,N_9550,N_9554,N_9557,N_9558,N_9559,N_9560,N_9561,N_9564,N_9565,N_9567,N_9568,N_9571,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9587,N_9590,N_9591,N_9593,N_9594,N_9595,N_9597,N_9598,N_9599,N_9603,N_9604,N_9605,N_9607,N_9609,N_9611,N_9612,N_9613,N_9614,N_9615,N_9618,N_9619,N_9621,N_9622,N_9625,N_9627,N_9631,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9640,N_9641,N_9642,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9653,N_9658,N_9659,N_9660,N_9662,N_9665,N_9667,N_9670,N_9671,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9681,N_9682,N_9683,N_9684,N_9689,N_9691,N_9693,N_9694,N_9697,N_9698,N_9699,N_9703,N_9705,N_9706,N_9710,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9721,N_9723,N_9725,N_9727,N_9728,N_9729,N_9730,N_9733,N_9735,N_9738,N_9739,N_9740,N_9743,N_9749,N_9753,N_9754,N_9755,N_9756,N_9757,N_9760,N_9761,N_9762,N_9765,N_9766,N_9767,N_9769,N_9770,N_9771,N_9773,N_9774,N_9775,N_9779,N_9780,N_9781,N_9784,N_9786,N_9788,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9801,N_9803,N_9804,N_9805,N_9807,N_9808,N_9810,N_9813,N_9814,N_9815,N_9816,N_9818,N_9819,N_9821,N_9822,N_9823,N_9826,N_9827,N_9828,N_9832,N_9833,N_9834,N_9835,N_9836,N_9839,N_9841,N_9842,N_9843,N_9844,N_9850,N_9851,N_9854,N_9855,N_9856,N_9858,N_9859,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9874,N_9876,N_9878,N_9882,N_9883,N_9884,N_9886,N_9887,N_9891,N_9892,N_9893,N_9896,N_9898,N_9900,N_9902,N_9903,N_9904,N_9905,N_9907,N_9908,N_9909,N_9911,N_9912,N_9913,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9924,N_9925,N_9927,N_9929,N_9935,N_9936,N_9937,N_9938,N_9942,N_9943,N_9945,N_9947,N_9951,N_9954,N_9955,N_9959,N_9961,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9971,N_9974,N_9975,N_9977,N_9978,N_9984,N_9985,N_9987,N_9988,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9999;
and U0 (N_0,In_715,In_862);
or U1 (N_1,In_204,In_172);
and U2 (N_2,In_410,In_173);
and U3 (N_3,In_148,In_470);
nor U4 (N_4,In_850,In_647);
or U5 (N_5,In_94,In_434);
or U6 (N_6,In_448,In_664);
and U7 (N_7,In_444,In_32);
or U8 (N_8,In_467,In_269);
or U9 (N_9,In_258,In_814);
and U10 (N_10,In_157,In_372);
nor U11 (N_11,In_104,In_183);
nand U12 (N_12,In_868,In_68);
or U13 (N_13,In_507,In_412);
or U14 (N_14,In_76,In_777);
or U15 (N_15,In_220,In_120);
nor U16 (N_16,In_798,In_234);
nand U17 (N_17,In_841,In_768);
nor U18 (N_18,In_922,In_266);
or U19 (N_19,In_252,In_766);
nand U20 (N_20,In_761,In_665);
or U21 (N_21,In_392,In_597);
and U22 (N_22,In_592,In_573);
and U23 (N_23,In_683,In_442);
nand U24 (N_24,In_343,In_737);
and U25 (N_25,In_318,In_539);
and U26 (N_26,In_880,In_418);
nand U27 (N_27,In_72,In_799);
nor U28 (N_28,In_322,In_793);
or U29 (N_29,In_757,In_602);
nor U30 (N_30,In_424,In_188);
nand U31 (N_31,In_363,In_297);
or U32 (N_32,In_888,In_180);
and U33 (N_33,In_670,In_274);
or U34 (N_34,In_519,In_505);
nor U35 (N_35,In_371,In_785);
nand U36 (N_36,In_83,In_631);
nand U37 (N_37,In_253,In_451);
and U38 (N_38,In_884,In_200);
and U39 (N_39,In_503,In_560);
and U40 (N_40,In_205,In_810);
nor U41 (N_41,In_201,In_36);
or U42 (N_42,In_358,In_991);
nor U43 (N_43,In_469,In_527);
nor U44 (N_44,In_136,In_751);
nor U45 (N_45,In_7,In_844);
and U46 (N_46,In_355,In_14);
nor U47 (N_47,In_818,In_228);
and U48 (N_48,In_895,In_796);
and U49 (N_49,In_826,In_979);
nand U50 (N_50,In_992,In_168);
or U51 (N_51,In_778,In_154);
and U52 (N_52,In_216,In_459);
and U53 (N_53,In_816,In_93);
nand U54 (N_54,In_845,In_864);
and U55 (N_55,In_137,In_189);
or U56 (N_56,In_73,In_755);
nand U57 (N_57,In_135,In_566);
nand U58 (N_58,In_501,In_985);
and U59 (N_59,In_33,In_346);
nor U60 (N_60,In_280,In_240);
or U61 (N_61,In_226,In_484);
and U62 (N_62,In_866,In_417);
nand U63 (N_63,In_194,In_693);
and U64 (N_64,In_341,In_208);
nand U65 (N_65,In_657,In_942);
or U66 (N_66,In_732,In_974);
xnor U67 (N_67,In_184,In_323);
or U68 (N_68,In_374,In_537);
nand U69 (N_69,In_476,In_313);
or U70 (N_70,In_382,In_70);
and U71 (N_71,In_175,In_572);
nor U72 (N_72,In_67,In_704);
nand U73 (N_73,In_820,In_49);
or U74 (N_74,In_497,In_262);
nor U75 (N_75,In_301,In_261);
nand U76 (N_76,In_995,In_753);
nand U77 (N_77,In_381,In_509);
or U78 (N_78,In_99,In_405);
nor U79 (N_79,In_164,In_743);
and U80 (N_80,In_831,In_975);
or U81 (N_81,In_515,In_292);
or U82 (N_82,In_911,In_812);
or U83 (N_83,In_697,In_764);
or U84 (N_84,In_186,In_538);
nand U85 (N_85,In_217,In_558);
and U86 (N_86,In_541,In_703);
nand U87 (N_87,In_998,In_615);
and U88 (N_88,In_177,In_811);
and U89 (N_89,In_516,In_265);
nand U90 (N_90,In_643,In_413);
nand U91 (N_91,In_859,In_399);
or U92 (N_92,In_807,In_999);
or U93 (N_93,In_147,In_257);
nand U94 (N_94,In_846,In_432);
nor U95 (N_95,In_155,In_856);
nor U96 (N_96,In_908,In_134);
or U97 (N_97,In_513,In_993);
and U98 (N_98,In_124,In_976);
nand U99 (N_99,In_359,In_806);
nor U100 (N_100,In_797,In_948);
and U101 (N_101,In_89,In_913);
nand U102 (N_102,In_331,In_421);
nor U103 (N_103,In_914,In_910);
and U104 (N_104,In_673,In_171);
nor U105 (N_105,In_722,In_851);
nor U106 (N_106,In_277,In_239);
or U107 (N_107,In_306,In_316);
or U108 (N_108,In_726,In_518);
nor U109 (N_109,In_493,In_475);
nand U110 (N_110,In_708,In_511);
nand U111 (N_111,In_229,In_928);
nor U112 (N_112,In_970,In_642);
and U113 (N_113,In_639,In_867);
nand U114 (N_114,In_494,In_464);
or U115 (N_115,In_508,In_984);
nand U116 (N_116,In_881,In_370);
nand U117 (N_117,In_391,In_746);
or U118 (N_118,In_953,In_563);
and U119 (N_119,In_672,In_242);
nand U120 (N_120,In_267,In_273);
or U121 (N_121,In_738,In_303);
nand U122 (N_122,In_601,In_871);
and U123 (N_123,In_907,In_312);
xor U124 (N_124,In_106,In_994);
and U125 (N_125,In_238,In_441);
and U126 (N_126,In_428,In_139);
nor U127 (N_127,In_546,In_415);
nand U128 (N_128,In_236,In_460);
nor U129 (N_129,In_619,In_794);
nand U130 (N_130,In_44,In_748);
nor U131 (N_131,In_455,In_533);
nand U132 (N_132,In_326,In_325);
and U133 (N_133,In_191,In_917);
nor U134 (N_134,In_271,In_309);
and U135 (N_135,In_608,In_512);
nor U136 (N_136,In_98,In_514);
and U137 (N_137,In_224,In_495);
and U138 (N_138,In_332,In_34);
or U139 (N_139,In_623,In_401);
and U140 (N_140,In_131,In_964);
or U141 (N_141,In_92,In_452);
or U142 (N_142,In_376,In_349);
and U143 (N_143,In_268,In_29);
and U144 (N_144,In_24,In_645);
or U145 (N_145,In_30,In_270);
and U146 (N_146,In_659,In_128);
nand U147 (N_147,In_122,In_365);
nand U148 (N_148,In_640,In_0);
and U149 (N_149,In_570,In_540);
nor U150 (N_150,In_287,In_237);
and U151 (N_151,In_354,In_815);
or U152 (N_152,In_660,In_2);
nor U153 (N_153,In_404,In_996);
and U154 (N_154,In_833,In_350);
nor U155 (N_155,In_65,In_574);
or U156 (N_156,In_641,In_593);
xnor U157 (N_157,In_259,In_912);
and U158 (N_158,In_586,In_825);
nor U159 (N_159,In_712,In_153);
and U160 (N_160,In_407,In_486);
nor U161 (N_161,In_959,In_677);
and U162 (N_162,In_838,In_161);
or U163 (N_163,In_179,In_159);
or U164 (N_164,In_101,In_808);
or U165 (N_165,In_174,In_754);
or U166 (N_166,In_215,In_938);
nor U167 (N_167,In_81,In_528);
or U168 (N_168,In_679,In_57);
and U169 (N_169,In_983,In_646);
nor U170 (N_170,In_3,In_957);
nand U171 (N_171,In_731,In_395);
or U172 (N_172,In_479,In_612);
nor U173 (N_173,In_710,In_906);
nor U174 (N_174,In_875,In_145);
xnor U175 (N_175,In_614,In_278);
nor U176 (N_176,In_130,In_351);
or U177 (N_177,In_698,In_225);
and U178 (N_178,In_109,In_377);
nand U179 (N_179,In_489,In_931);
and U180 (N_180,In_689,In_110);
and U181 (N_181,In_22,In_561);
nand U182 (N_182,In_185,In_899);
and U183 (N_183,In_324,In_709);
nand U184 (N_184,In_9,In_190);
nor U185 (N_185,In_305,In_655);
nor U186 (N_186,In_716,In_676);
nor U187 (N_187,In_396,In_891);
nor U188 (N_188,In_43,In_594);
and U189 (N_189,In_883,In_954);
xnor U190 (N_190,In_763,In_687);
or U191 (N_191,In_209,In_232);
and U192 (N_192,In_750,In_565);
or U193 (N_193,In_213,In_842);
nand U194 (N_194,In_613,In_781);
nand U195 (N_195,In_15,In_218);
nand U196 (N_196,In_182,In_207);
or U197 (N_197,In_767,In_304);
or U198 (N_198,In_66,In_827);
and U199 (N_199,In_530,In_1);
and U200 (N_200,In_133,In_830);
and U201 (N_201,In_384,In_411);
nor U202 (N_202,In_10,In_936);
nor U203 (N_203,In_552,In_564);
nand U204 (N_204,In_127,In_345);
nor U205 (N_205,In_474,In_946);
nor U206 (N_206,In_387,In_658);
and U207 (N_207,In_490,In_456);
and U208 (N_208,In_553,In_809);
or U209 (N_209,In_74,In_690);
nor U210 (N_210,In_531,In_802);
nor U211 (N_211,In_621,In_944);
nor U212 (N_212,In_963,In_12);
or U213 (N_213,In_952,In_822);
nand U214 (N_214,In_924,In_571);
or U215 (N_215,In_939,In_836);
nor U216 (N_216,In_523,In_863);
or U217 (N_217,In_656,In_422);
and U218 (N_218,In_247,In_115);
and U219 (N_219,In_562,In_918);
and U220 (N_220,In_400,In_477);
or U221 (N_221,In_91,In_95);
or U222 (N_222,In_885,In_583);
or U223 (N_223,In_638,In_357);
nand U224 (N_224,In_940,In_554);
or U225 (N_225,In_299,In_744);
and U226 (N_226,In_887,In_196);
nor U227 (N_227,In_40,In_107);
nand U228 (N_228,In_680,In_719);
nand U229 (N_229,In_307,In_6);
and U230 (N_230,In_852,In_532);
or U231 (N_231,In_694,In_627);
nand U232 (N_232,In_745,In_786);
or U233 (N_233,In_702,In_667);
and U234 (N_234,In_803,In_958);
or U235 (N_235,In_315,In_51);
or U236 (N_236,In_26,In_500);
nand U237 (N_237,In_791,In_425);
or U238 (N_238,In_480,In_142);
nand U239 (N_239,In_792,In_662);
or U240 (N_240,In_718,In_861);
nor U241 (N_241,In_466,In_210);
nand U242 (N_242,In_853,In_282);
nand U243 (N_243,In_443,In_149);
and U244 (N_244,In_364,In_348);
and U245 (N_245,In_705,In_166);
and U246 (N_246,In_295,In_978);
nor U247 (N_247,In_310,In_813);
nand U248 (N_248,In_577,In_882);
nand U249 (N_249,In_787,In_281);
or U250 (N_250,In_111,In_943);
nor U251 (N_251,In_765,In_916);
nor U252 (N_252,In_96,In_473);
or U253 (N_253,In_223,In_622);
and U254 (N_254,In_692,In_669);
nand U255 (N_255,In_966,In_340);
or U256 (N_256,In_839,In_487);
xor U257 (N_257,In_260,In_522);
nand U258 (N_258,In_626,In_872);
or U259 (N_259,In_937,In_45);
nor U260 (N_260,In_661,In_535);
nand U261 (N_261,In_961,In_596);
and U262 (N_262,In_595,In_870);
and U263 (N_263,In_502,In_835);
nor U264 (N_264,In_905,In_485);
nand U265 (N_265,In_776,In_431);
and U266 (N_266,In_321,In_114);
and U267 (N_267,In_248,In_187);
or U268 (N_268,In_847,In_178);
nand U269 (N_269,In_103,In_52);
nor U270 (N_270,In_255,In_385);
nand U271 (N_271,In_610,In_821);
or U272 (N_272,In_653,In_279);
nand U273 (N_273,In_86,In_333);
or U274 (N_274,In_982,In_921);
and U275 (N_275,In_580,In_534);
or U276 (N_276,In_169,In_526);
and U277 (N_277,In_393,In_688);
or U278 (N_278,In_206,In_618);
or U279 (N_279,In_64,In_249);
nand U280 (N_280,In_181,In_909);
or U281 (N_281,In_8,In_633);
xnor U282 (N_282,In_13,In_648);
or U283 (N_283,In_857,In_457);
and U284 (N_284,In_50,In_233);
xor U285 (N_285,In_138,In_294);
nor U286 (N_286,In_406,In_699);
nand U287 (N_287,In_80,In_890);
nand U288 (N_288,In_150,In_873);
nand U289 (N_289,In_987,In_288);
nor U290 (N_290,In_293,In_214);
or U291 (N_291,In_625,In_706);
nand U292 (N_292,In_569,In_197);
or U293 (N_293,In_230,In_789);
and U294 (N_294,In_617,In_607);
and U295 (N_295,In_654,In_747);
nand U296 (N_296,In_21,In_823);
nor U297 (N_297,In_876,In_504);
or U298 (N_298,In_369,In_430);
nand U299 (N_299,In_678,In_499);
nor U300 (N_300,In_723,In_129);
and U301 (N_301,In_721,In_90);
nor U302 (N_302,In_624,In_419);
nand U303 (N_303,In_988,In_433);
nor U304 (N_304,In_893,In_837);
or U305 (N_305,In_492,In_828);
nor U306 (N_306,In_491,In_462);
nor U307 (N_307,In_256,In_285);
nand U308 (N_308,In_311,In_517);
or U309 (N_309,In_276,In_557);
nand U310 (N_310,In_900,In_632);
nand U311 (N_311,In_663,In_222);
or U312 (N_312,In_123,In_79);
xnor U313 (N_313,In_770,In_152);
and U314 (N_314,In_735,In_556);
nor U315 (N_315,In_46,In_356);
nand U316 (N_316,In_934,In_611);
and U317 (N_317,In_758,In_858);
and U318 (N_318,In_529,In_652);
nand U319 (N_319,In_840,In_675);
xor U320 (N_320,In_771,In_724);
nor U321 (N_321,In_132,In_481);
nand U322 (N_322,In_956,In_775);
and U323 (N_323,In_17,In_446);
nand U324 (N_324,In_930,In_31);
or U325 (N_325,In_77,In_437);
or U326 (N_326,In_227,In_100);
nor U327 (N_327,In_752,In_686);
nor U328 (N_328,In_666,In_423);
or U329 (N_329,In_160,In_892);
nand U330 (N_330,In_585,In_965);
or U331 (N_331,In_843,In_860);
or U332 (N_332,In_482,In_420);
nor U333 (N_333,In_603,In_590);
and U334 (N_334,In_458,In_714);
nand U335 (N_335,In_926,In_877);
nor U336 (N_336,In_591,In_11);
or U337 (N_337,In_496,In_829);
nand U338 (N_338,In_849,In_498);
or U339 (N_339,In_5,In_362);
nor U340 (N_340,In_336,In_383);
and U341 (N_341,In_616,In_25);
or U342 (N_342,In_366,In_163);
nor U343 (N_343,In_337,In_547);
and U344 (N_344,In_329,In_582);
xor U345 (N_345,In_733,In_390);
or U346 (N_346,In_973,In_932);
nor U347 (N_347,In_636,In_55);
nor U348 (N_348,In_193,In_449);
nand U349 (N_349,In_435,In_720);
nor U350 (N_350,In_426,In_804);
and U351 (N_351,In_241,In_375);
or U352 (N_352,In_69,In_955);
nand U353 (N_353,In_854,In_581);
nor U354 (N_354,In_730,In_682);
nor U355 (N_355,In_819,In_634);
and U356 (N_356,In_61,In_865);
nand U357 (N_357,In_403,In_711);
nor U358 (N_358,In_118,In_472);
nand U359 (N_359,In_598,In_378);
and U360 (N_360,In_298,In_971);
nor U361 (N_361,In_684,In_219);
and U362 (N_362,In_170,In_725);
or U363 (N_363,In_707,In_695);
or U364 (N_364,In_167,In_674);
nor U365 (N_365,In_254,In_398);
nor U366 (N_366,In_780,In_729);
nor U367 (N_367,In_445,In_935);
or U368 (N_368,In_54,In_379);
and U369 (N_369,In_87,In_454);
or U370 (N_370,In_555,In_923);
nand U371 (N_371,In_402,In_19);
nor U372 (N_372,In_668,In_203);
nand U373 (N_373,In_88,In_869);
or U374 (N_374,In_314,In_981);
or U375 (N_375,In_328,In_126);
nand U376 (N_376,In_782,In_896);
and U377 (N_377,In_728,In_408);
nand U378 (N_378,In_394,In_388);
and U379 (N_379,In_915,In_251);
and U380 (N_380,In_713,In_296);
nor U381 (N_381,In_524,In_635);
or U382 (N_382,In_342,In_628);
nand U383 (N_383,In_198,In_20);
nor U384 (N_384,In_438,In_264);
or U385 (N_385,In_416,In_542);
nor U386 (N_386,In_604,In_62);
or U387 (N_387,In_801,In_549);
or U388 (N_388,In_536,In_283);
nor U389 (N_389,In_760,In_904);
and U390 (N_390,In_275,In_60);
nand U391 (N_391,In_568,In_4);
nand U392 (N_392,In_461,In_327);
nand U393 (N_393,In_263,In_788);
and U394 (N_394,In_947,In_483);
or U395 (N_395,In_949,In_116);
nor U396 (N_396,In_18,In_739);
and U397 (N_397,In_567,In_986);
and U398 (N_398,In_784,In_620);
and U399 (N_399,In_587,In_951);
nand U400 (N_400,In_286,In_38);
or U401 (N_401,In_889,In_834);
nor U402 (N_402,In_78,In_37);
nand U403 (N_403,In_990,In_800);
nor U404 (N_404,In_246,In_344);
or U405 (N_405,In_550,In_589);
or U406 (N_406,In_629,In_28);
and U407 (N_407,In_980,In_158);
nand U408 (N_408,In_644,In_151);
or U409 (N_409,In_681,In_972);
and U410 (N_410,In_832,In_649);
nor U411 (N_411,In_386,In_960);
nor U412 (N_412,In_544,In_339);
nand U413 (N_413,In_997,In_736);
and U414 (N_414,In_521,In_691);
nor U415 (N_415,In_927,In_48);
nor U416 (N_416,In_319,In_898);
or U417 (N_417,In_16,In_63);
nand U418 (N_418,In_27,In_244);
nor U419 (N_419,In_579,In_609);
nor U420 (N_420,In_272,In_548);
or U421 (N_421,In_289,In_925);
or U422 (N_422,In_671,In_463);
and U423 (N_423,In_165,In_685);
nor U424 (N_424,In_41,In_117);
nand U425 (N_425,In_968,In_941);
nor U426 (N_426,In_734,In_762);
nand U427 (N_427,In_105,In_637);
nor U428 (N_428,In_284,In_773);
nand U429 (N_429,In_429,In_75);
nand U430 (N_430,In_605,In_969);
and U431 (N_431,In_855,In_933);
or U432 (N_432,In_520,In_334);
xnor U433 (N_433,In_878,In_967);
nor U434 (N_434,In_478,In_606);
and U435 (N_435,In_848,In_397);
and U436 (N_436,In_510,In_450);
nor U437 (N_437,In_389,In_414);
or U438 (N_438,In_59,In_156);
and U439 (N_439,In_112,In_950);
nand U440 (N_440,In_361,In_929);
nor U441 (N_441,In_874,In_779);
nor U442 (N_442,In_805,In_584);
and U443 (N_443,In_576,In_290);
and U444 (N_444,In_600,In_85);
or U445 (N_445,In_551,In_250);
or U446 (N_446,In_919,In_195);
nor U447 (N_447,In_47,In_108);
nand U448 (N_448,In_212,In_920);
nand U449 (N_449,In_360,In_465);
nor U450 (N_450,In_774,In_901);
nor U451 (N_451,In_488,In_427);
and U452 (N_452,In_58,In_367);
and U453 (N_453,In_373,In_347);
and U454 (N_454,In_468,In_176);
nand U455 (N_455,In_338,In_989);
nor U456 (N_456,In_352,In_97);
and U457 (N_457,In_409,In_144);
and U458 (N_458,In_742,In_795);
and U459 (N_459,In_440,In_300);
or U460 (N_460,In_439,In_783);
and U461 (N_461,In_545,In_353);
nor U462 (N_462,In_113,In_543);
nor U463 (N_463,In_650,In_962);
or U464 (N_464,In_141,In_102);
nor U465 (N_465,In_772,In_817);
nor U466 (N_466,In_790,In_243);
or U467 (N_467,In_42,In_245);
nor U468 (N_468,In_879,In_894);
or U469 (N_469,In_308,In_902);
and U470 (N_470,In_23,In_977);
nand U471 (N_471,In_125,In_302);
nand U472 (N_472,In_559,In_903);
nand U473 (N_473,In_727,In_471);
and U474 (N_474,In_769,In_506);
and U475 (N_475,In_121,In_291);
and U476 (N_476,In_740,In_886);
nand U477 (N_477,In_436,In_330);
nand U478 (N_478,In_897,In_320);
nand U479 (N_479,In_35,In_317);
or U480 (N_480,In_717,In_146);
nor U481 (N_481,In_82,In_235);
nor U482 (N_482,In_578,In_696);
nand U483 (N_483,In_162,In_231);
nor U484 (N_484,In_756,In_824);
nor U485 (N_485,In_701,In_630);
or U486 (N_486,In_39,In_945);
or U487 (N_487,In_759,In_199);
nand U488 (N_488,In_192,In_84);
nor U489 (N_489,In_143,In_453);
nand U490 (N_490,In_749,In_651);
nand U491 (N_491,In_56,In_335);
nor U492 (N_492,In_221,In_447);
or U493 (N_493,In_588,In_368);
nand U494 (N_494,In_575,In_53);
or U495 (N_495,In_380,In_599);
nor U496 (N_496,In_741,In_71);
nor U497 (N_497,In_202,In_700);
nor U498 (N_498,In_140,In_211);
nand U499 (N_499,In_119,In_525);
or U500 (N_500,In_64,In_849);
and U501 (N_501,In_298,In_772);
nand U502 (N_502,In_67,In_965);
nand U503 (N_503,In_502,In_23);
or U504 (N_504,In_683,In_728);
or U505 (N_505,In_35,In_47);
nor U506 (N_506,In_113,In_442);
nor U507 (N_507,In_683,In_505);
and U508 (N_508,In_504,In_372);
and U509 (N_509,In_369,In_341);
nand U510 (N_510,In_189,In_547);
nor U511 (N_511,In_184,In_377);
nand U512 (N_512,In_708,In_197);
nor U513 (N_513,In_726,In_779);
nand U514 (N_514,In_326,In_205);
nor U515 (N_515,In_38,In_34);
and U516 (N_516,In_751,In_934);
and U517 (N_517,In_271,In_916);
xor U518 (N_518,In_877,In_965);
or U519 (N_519,In_603,In_278);
and U520 (N_520,In_82,In_366);
xnor U521 (N_521,In_196,In_464);
nand U522 (N_522,In_622,In_724);
or U523 (N_523,In_437,In_115);
and U524 (N_524,In_705,In_524);
nand U525 (N_525,In_130,In_874);
nand U526 (N_526,In_794,In_219);
and U527 (N_527,In_780,In_22);
or U528 (N_528,In_586,In_564);
and U529 (N_529,In_185,In_747);
or U530 (N_530,In_138,In_924);
xor U531 (N_531,In_419,In_423);
or U532 (N_532,In_928,In_933);
or U533 (N_533,In_743,In_57);
and U534 (N_534,In_152,In_704);
or U535 (N_535,In_872,In_6);
and U536 (N_536,In_621,In_414);
nand U537 (N_537,In_698,In_274);
nor U538 (N_538,In_885,In_404);
or U539 (N_539,In_661,In_879);
and U540 (N_540,In_274,In_555);
nor U541 (N_541,In_580,In_711);
nand U542 (N_542,In_883,In_501);
or U543 (N_543,In_976,In_945);
nand U544 (N_544,In_758,In_971);
or U545 (N_545,In_929,In_285);
and U546 (N_546,In_655,In_911);
nand U547 (N_547,In_500,In_483);
or U548 (N_548,In_831,In_644);
nor U549 (N_549,In_853,In_608);
or U550 (N_550,In_275,In_222);
and U551 (N_551,In_841,In_147);
or U552 (N_552,In_755,In_959);
xor U553 (N_553,In_838,In_687);
nor U554 (N_554,In_741,In_718);
and U555 (N_555,In_303,In_591);
or U556 (N_556,In_686,In_277);
nand U557 (N_557,In_468,In_221);
or U558 (N_558,In_431,In_313);
nor U559 (N_559,In_947,In_361);
or U560 (N_560,In_604,In_974);
nand U561 (N_561,In_694,In_771);
and U562 (N_562,In_695,In_255);
nor U563 (N_563,In_796,In_570);
nor U564 (N_564,In_667,In_670);
or U565 (N_565,In_619,In_539);
and U566 (N_566,In_629,In_234);
or U567 (N_567,In_42,In_741);
or U568 (N_568,In_999,In_307);
nand U569 (N_569,In_972,In_218);
and U570 (N_570,In_686,In_875);
or U571 (N_571,In_59,In_944);
nand U572 (N_572,In_632,In_444);
nor U573 (N_573,In_651,In_95);
and U574 (N_574,In_856,In_878);
nand U575 (N_575,In_434,In_497);
nand U576 (N_576,In_248,In_286);
and U577 (N_577,In_963,In_71);
nand U578 (N_578,In_22,In_424);
nor U579 (N_579,In_322,In_71);
and U580 (N_580,In_111,In_5);
nand U581 (N_581,In_149,In_172);
or U582 (N_582,In_230,In_627);
and U583 (N_583,In_231,In_446);
and U584 (N_584,In_161,In_910);
or U585 (N_585,In_254,In_692);
nor U586 (N_586,In_600,In_292);
nand U587 (N_587,In_267,In_810);
nor U588 (N_588,In_64,In_926);
or U589 (N_589,In_320,In_9);
or U590 (N_590,In_691,In_533);
and U591 (N_591,In_56,In_728);
nor U592 (N_592,In_938,In_895);
nand U593 (N_593,In_870,In_136);
nor U594 (N_594,In_187,In_554);
nand U595 (N_595,In_884,In_312);
nand U596 (N_596,In_837,In_983);
nor U597 (N_597,In_540,In_714);
nand U598 (N_598,In_751,In_25);
and U599 (N_599,In_749,In_446);
nor U600 (N_600,In_161,In_152);
and U601 (N_601,In_762,In_344);
nand U602 (N_602,In_459,In_498);
or U603 (N_603,In_819,In_157);
nor U604 (N_604,In_675,In_587);
nor U605 (N_605,In_311,In_451);
nand U606 (N_606,In_493,In_702);
xor U607 (N_607,In_989,In_670);
nor U608 (N_608,In_603,In_949);
or U609 (N_609,In_164,In_819);
or U610 (N_610,In_526,In_802);
nor U611 (N_611,In_14,In_91);
and U612 (N_612,In_972,In_350);
and U613 (N_613,In_620,In_758);
nor U614 (N_614,In_979,In_124);
nor U615 (N_615,In_401,In_246);
and U616 (N_616,In_647,In_410);
nand U617 (N_617,In_211,In_772);
nor U618 (N_618,In_729,In_311);
and U619 (N_619,In_976,In_735);
nor U620 (N_620,In_510,In_277);
and U621 (N_621,In_916,In_933);
and U622 (N_622,In_878,In_759);
nor U623 (N_623,In_625,In_988);
xor U624 (N_624,In_483,In_325);
or U625 (N_625,In_583,In_876);
or U626 (N_626,In_317,In_672);
and U627 (N_627,In_649,In_671);
or U628 (N_628,In_824,In_650);
or U629 (N_629,In_304,In_835);
nand U630 (N_630,In_21,In_426);
or U631 (N_631,In_896,In_406);
or U632 (N_632,In_454,In_761);
nand U633 (N_633,In_554,In_930);
xor U634 (N_634,In_368,In_359);
nor U635 (N_635,In_367,In_403);
or U636 (N_636,In_948,In_904);
nor U637 (N_637,In_345,In_392);
nand U638 (N_638,In_930,In_8);
nor U639 (N_639,In_554,In_715);
nand U640 (N_640,In_551,In_920);
nand U641 (N_641,In_517,In_920);
nor U642 (N_642,In_802,In_659);
nand U643 (N_643,In_52,In_604);
nand U644 (N_644,In_716,In_660);
and U645 (N_645,In_326,In_858);
nor U646 (N_646,In_493,In_383);
nor U647 (N_647,In_495,In_710);
nand U648 (N_648,In_538,In_828);
nor U649 (N_649,In_490,In_109);
or U650 (N_650,In_710,In_392);
nand U651 (N_651,In_880,In_744);
or U652 (N_652,In_531,In_381);
and U653 (N_653,In_13,In_34);
and U654 (N_654,In_707,In_733);
nor U655 (N_655,In_639,In_125);
or U656 (N_656,In_804,In_945);
or U657 (N_657,In_640,In_611);
nor U658 (N_658,In_459,In_397);
and U659 (N_659,In_974,In_173);
nor U660 (N_660,In_460,In_688);
and U661 (N_661,In_93,In_732);
or U662 (N_662,In_853,In_91);
nor U663 (N_663,In_108,In_498);
nor U664 (N_664,In_955,In_368);
nand U665 (N_665,In_23,In_405);
and U666 (N_666,In_843,In_99);
and U667 (N_667,In_743,In_770);
and U668 (N_668,In_55,In_487);
or U669 (N_669,In_521,In_353);
and U670 (N_670,In_292,In_928);
nand U671 (N_671,In_310,In_870);
nor U672 (N_672,In_202,In_290);
or U673 (N_673,In_208,In_990);
and U674 (N_674,In_884,In_823);
nand U675 (N_675,In_692,In_40);
nand U676 (N_676,In_792,In_111);
nand U677 (N_677,In_73,In_698);
or U678 (N_678,In_205,In_690);
or U679 (N_679,In_985,In_493);
and U680 (N_680,In_823,In_802);
nor U681 (N_681,In_950,In_25);
nor U682 (N_682,In_636,In_601);
nand U683 (N_683,In_287,In_857);
nand U684 (N_684,In_295,In_329);
or U685 (N_685,In_958,In_582);
and U686 (N_686,In_394,In_751);
nand U687 (N_687,In_491,In_418);
nand U688 (N_688,In_528,In_682);
and U689 (N_689,In_88,In_662);
or U690 (N_690,In_832,In_28);
and U691 (N_691,In_897,In_248);
or U692 (N_692,In_644,In_501);
nor U693 (N_693,In_249,In_882);
and U694 (N_694,In_422,In_640);
or U695 (N_695,In_573,In_44);
or U696 (N_696,In_807,In_723);
nand U697 (N_697,In_600,In_804);
nor U698 (N_698,In_292,In_65);
nor U699 (N_699,In_670,In_440);
nor U700 (N_700,In_290,In_523);
or U701 (N_701,In_410,In_332);
nor U702 (N_702,In_756,In_894);
or U703 (N_703,In_553,In_288);
and U704 (N_704,In_498,In_191);
nand U705 (N_705,In_737,In_266);
nor U706 (N_706,In_28,In_874);
or U707 (N_707,In_882,In_83);
nand U708 (N_708,In_863,In_746);
nand U709 (N_709,In_778,In_107);
nor U710 (N_710,In_777,In_868);
nand U711 (N_711,In_755,In_198);
and U712 (N_712,In_132,In_109);
nand U713 (N_713,In_488,In_329);
or U714 (N_714,In_922,In_131);
nand U715 (N_715,In_829,In_208);
or U716 (N_716,In_326,In_227);
nor U717 (N_717,In_93,In_644);
nor U718 (N_718,In_975,In_564);
or U719 (N_719,In_75,In_844);
and U720 (N_720,In_592,In_42);
or U721 (N_721,In_397,In_212);
nor U722 (N_722,In_254,In_341);
nor U723 (N_723,In_926,In_39);
nand U724 (N_724,In_328,In_594);
and U725 (N_725,In_964,In_379);
and U726 (N_726,In_115,In_218);
and U727 (N_727,In_983,In_917);
nor U728 (N_728,In_723,In_999);
nand U729 (N_729,In_520,In_272);
or U730 (N_730,In_337,In_635);
or U731 (N_731,In_747,In_564);
and U732 (N_732,In_305,In_441);
or U733 (N_733,In_424,In_897);
or U734 (N_734,In_643,In_370);
or U735 (N_735,In_288,In_446);
nand U736 (N_736,In_144,In_143);
nand U737 (N_737,In_333,In_971);
nor U738 (N_738,In_751,In_646);
and U739 (N_739,In_29,In_273);
or U740 (N_740,In_207,In_356);
nor U741 (N_741,In_731,In_319);
nand U742 (N_742,In_844,In_177);
nand U743 (N_743,In_726,In_579);
nand U744 (N_744,In_621,In_966);
or U745 (N_745,In_988,In_770);
nand U746 (N_746,In_493,In_684);
nor U747 (N_747,In_41,In_330);
or U748 (N_748,In_506,In_846);
nor U749 (N_749,In_681,In_534);
nand U750 (N_750,In_358,In_244);
nand U751 (N_751,In_734,In_185);
and U752 (N_752,In_815,In_726);
nor U753 (N_753,In_825,In_593);
nor U754 (N_754,In_878,In_322);
or U755 (N_755,In_644,In_379);
nand U756 (N_756,In_391,In_448);
nand U757 (N_757,In_57,In_636);
or U758 (N_758,In_938,In_841);
nand U759 (N_759,In_730,In_339);
nor U760 (N_760,In_36,In_967);
nor U761 (N_761,In_750,In_46);
nand U762 (N_762,In_556,In_23);
nand U763 (N_763,In_231,In_35);
or U764 (N_764,In_580,In_751);
or U765 (N_765,In_190,In_482);
nand U766 (N_766,In_937,In_443);
nand U767 (N_767,In_845,In_417);
nand U768 (N_768,In_25,In_326);
and U769 (N_769,In_333,In_669);
nand U770 (N_770,In_808,In_932);
nor U771 (N_771,In_751,In_489);
or U772 (N_772,In_994,In_888);
and U773 (N_773,In_579,In_818);
nor U774 (N_774,In_951,In_564);
nor U775 (N_775,In_693,In_441);
or U776 (N_776,In_512,In_869);
nand U777 (N_777,In_28,In_938);
nor U778 (N_778,In_225,In_66);
or U779 (N_779,In_315,In_933);
nand U780 (N_780,In_871,In_243);
nor U781 (N_781,In_755,In_756);
or U782 (N_782,In_517,In_717);
or U783 (N_783,In_693,In_349);
nand U784 (N_784,In_48,In_833);
and U785 (N_785,In_311,In_186);
nand U786 (N_786,In_316,In_765);
nor U787 (N_787,In_384,In_651);
nor U788 (N_788,In_538,In_700);
nand U789 (N_789,In_73,In_785);
nor U790 (N_790,In_248,In_490);
and U791 (N_791,In_100,In_748);
and U792 (N_792,In_744,In_468);
and U793 (N_793,In_401,In_67);
nand U794 (N_794,In_588,In_999);
or U795 (N_795,In_231,In_208);
nand U796 (N_796,In_81,In_801);
or U797 (N_797,In_852,In_584);
or U798 (N_798,In_5,In_489);
or U799 (N_799,In_531,In_334);
or U800 (N_800,In_707,In_223);
or U801 (N_801,In_775,In_486);
and U802 (N_802,In_755,In_884);
nor U803 (N_803,In_465,In_843);
and U804 (N_804,In_343,In_851);
nand U805 (N_805,In_293,In_871);
nand U806 (N_806,In_430,In_977);
nand U807 (N_807,In_649,In_572);
nor U808 (N_808,In_203,In_557);
or U809 (N_809,In_476,In_50);
nand U810 (N_810,In_93,In_160);
or U811 (N_811,In_268,In_410);
nand U812 (N_812,In_672,In_636);
or U813 (N_813,In_66,In_30);
xnor U814 (N_814,In_976,In_636);
and U815 (N_815,In_102,In_982);
and U816 (N_816,In_212,In_596);
and U817 (N_817,In_355,In_907);
or U818 (N_818,In_188,In_124);
nand U819 (N_819,In_900,In_262);
nor U820 (N_820,In_988,In_165);
nand U821 (N_821,In_538,In_999);
and U822 (N_822,In_177,In_143);
or U823 (N_823,In_149,In_732);
and U824 (N_824,In_896,In_875);
nor U825 (N_825,In_912,In_565);
or U826 (N_826,In_592,In_829);
nand U827 (N_827,In_807,In_286);
or U828 (N_828,In_248,In_358);
or U829 (N_829,In_227,In_331);
and U830 (N_830,In_565,In_403);
nor U831 (N_831,In_109,In_46);
nor U832 (N_832,In_73,In_672);
or U833 (N_833,In_637,In_268);
nand U834 (N_834,In_209,In_516);
nand U835 (N_835,In_488,In_392);
or U836 (N_836,In_186,In_572);
or U837 (N_837,In_989,In_795);
nor U838 (N_838,In_736,In_91);
or U839 (N_839,In_211,In_160);
or U840 (N_840,In_377,In_887);
and U841 (N_841,In_609,In_320);
and U842 (N_842,In_236,In_900);
nand U843 (N_843,In_156,In_970);
and U844 (N_844,In_66,In_73);
and U845 (N_845,In_221,In_866);
nand U846 (N_846,In_458,In_895);
and U847 (N_847,In_467,In_349);
nand U848 (N_848,In_778,In_506);
or U849 (N_849,In_481,In_286);
and U850 (N_850,In_839,In_666);
or U851 (N_851,In_190,In_805);
or U852 (N_852,In_806,In_317);
nor U853 (N_853,In_438,In_241);
and U854 (N_854,In_474,In_546);
nor U855 (N_855,In_42,In_124);
and U856 (N_856,In_839,In_425);
or U857 (N_857,In_774,In_70);
nor U858 (N_858,In_881,In_987);
or U859 (N_859,In_854,In_185);
and U860 (N_860,In_374,In_418);
nand U861 (N_861,In_209,In_335);
or U862 (N_862,In_424,In_550);
nor U863 (N_863,In_956,In_471);
or U864 (N_864,In_796,In_342);
xnor U865 (N_865,In_773,In_954);
nand U866 (N_866,In_195,In_358);
nor U867 (N_867,In_975,In_917);
and U868 (N_868,In_355,In_473);
nor U869 (N_869,In_345,In_869);
nor U870 (N_870,In_884,In_467);
and U871 (N_871,In_0,In_699);
nor U872 (N_872,In_818,In_208);
nor U873 (N_873,In_404,In_217);
and U874 (N_874,In_99,In_812);
or U875 (N_875,In_82,In_442);
nand U876 (N_876,In_784,In_218);
nand U877 (N_877,In_957,In_438);
and U878 (N_878,In_322,In_867);
nand U879 (N_879,In_320,In_17);
nand U880 (N_880,In_794,In_488);
or U881 (N_881,In_352,In_559);
or U882 (N_882,In_879,In_666);
and U883 (N_883,In_829,In_547);
nand U884 (N_884,In_834,In_576);
nor U885 (N_885,In_149,In_645);
and U886 (N_886,In_94,In_703);
and U887 (N_887,In_267,In_925);
nor U888 (N_888,In_372,In_64);
nand U889 (N_889,In_961,In_320);
nand U890 (N_890,In_439,In_972);
nand U891 (N_891,In_968,In_827);
or U892 (N_892,In_494,In_286);
nand U893 (N_893,In_589,In_646);
or U894 (N_894,In_544,In_471);
nor U895 (N_895,In_172,In_133);
nor U896 (N_896,In_61,In_743);
and U897 (N_897,In_531,In_687);
or U898 (N_898,In_121,In_977);
nor U899 (N_899,In_804,In_108);
nand U900 (N_900,In_370,In_299);
or U901 (N_901,In_325,In_805);
nand U902 (N_902,In_789,In_794);
nand U903 (N_903,In_989,In_420);
or U904 (N_904,In_837,In_926);
and U905 (N_905,In_259,In_671);
or U906 (N_906,In_979,In_566);
or U907 (N_907,In_342,In_249);
or U908 (N_908,In_133,In_436);
and U909 (N_909,In_538,In_324);
nand U910 (N_910,In_64,In_702);
nor U911 (N_911,In_311,In_509);
and U912 (N_912,In_390,In_520);
or U913 (N_913,In_408,In_450);
nand U914 (N_914,In_976,In_173);
nand U915 (N_915,In_329,In_519);
and U916 (N_916,In_294,In_388);
and U917 (N_917,In_807,In_3);
and U918 (N_918,In_296,In_946);
nor U919 (N_919,In_662,In_891);
nand U920 (N_920,In_88,In_249);
or U921 (N_921,In_170,In_377);
or U922 (N_922,In_68,In_388);
nor U923 (N_923,In_399,In_898);
or U924 (N_924,In_89,In_416);
nor U925 (N_925,In_171,In_34);
nor U926 (N_926,In_783,In_219);
or U927 (N_927,In_383,In_598);
nand U928 (N_928,In_312,In_1);
nor U929 (N_929,In_125,In_45);
nor U930 (N_930,In_456,In_373);
or U931 (N_931,In_461,In_933);
nand U932 (N_932,In_380,In_543);
or U933 (N_933,In_465,In_256);
nand U934 (N_934,In_485,In_163);
nor U935 (N_935,In_146,In_598);
nand U936 (N_936,In_474,In_642);
nor U937 (N_937,In_778,In_981);
and U938 (N_938,In_456,In_87);
nand U939 (N_939,In_799,In_195);
nand U940 (N_940,In_309,In_24);
and U941 (N_941,In_593,In_487);
and U942 (N_942,In_599,In_96);
or U943 (N_943,In_838,In_323);
or U944 (N_944,In_759,In_625);
or U945 (N_945,In_967,In_364);
or U946 (N_946,In_706,In_396);
nor U947 (N_947,In_569,In_661);
or U948 (N_948,In_762,In_851);
or U949 (N_949,In_198,In_203);
nand U950 (N_950,In_10,In_330);
nor U951 (N_951,In_794,In_332);
nor U952 (N_952,In_974,In_616);
and U953 (N_953,In_609,In_577);
nand U954 (N_954,In_268,In_69);
and U955 (N_955,In_228,In_181);
and U956 (N_956,In_211,In_591);
nand U957 (N_957,In_350,In_611);
and U958 (N_958,In_633,In_943);
or U959 (N_959,In_700,In_479);
nand U960 (N_960,In_353,In_102);
nand U961 (N_961,In_391,In_499);
nand U962 (N_962,In_130,In_936);
nor U963 (N_963,In_64,In_963);
nand U964 (N_964,In_518,In_663);
and U965 (N_965,In_12,In_183);
or U966 (N_966,In_64,In_1);
nor U967 (N_967,In_242,In_911);
nand U968 (N_968,In_928,In_744);
nand U969 (N_969,In_22,In_188);
nand U970 (N_970,In_181,In_85);
nor U971 (N_971,In_850,In_102);
nand U972 (N_972,In_963,In_128);
nand U973 (N_973,In_607,In_170);
or U974 (N_974,In_224,In_634);
or U975 (N_975,In_525,In_776);
or U976 (N_976,In_441,In_623);
nor U977 (N_977,In_396,In_303);
or U978 (N_978,In_623,In_127);
nand U979 (N_979,In_67,In_855);
nor U980 (N_980,In_268,In_668);
or U981 (N_981,In_726,In_191);
or U982 (N_982,In_970,In_599);
or U983 (N_983,In_223,In_502);
nand U984 (N_984,In_688,In_234);
and U985 (N_985,In_569,In_715);
and U986 (N_986,In_556,In_277);
and U987 (N_987,In_511,In_873);
or U988 (N_988,In_281,In_603);
nand U989 (N_989,In_394,In_495);
nor U990 (N_990,In_891,In_4);
or U991 (N_991,In_901,In_16);
and U992 (N_992,In_828,In_972);
nor U993 (N_993,In_635,In_582);
and U994 (N_994,In_199,In_319);
nor U995 (N_995,In_352,In_176);
or U996 (N_996,In_370,In_957);
nand U997 (N_997,In_580,In_914);
nor U998 (N_998,In_240,In_440);
nand U999 (N_999,In_942,In_257);
or U1000 (N_1000,In_687,In_833);
and U1001 (N_1001,In_29,In_898);
or U1002 (N_1002,In_863,In_178);
or U1003 (N_1003,In_250,In_98);
nand U1004 (N_1004,In_322,In_317);
and U1005 (N_1005,In_115,In_710);
nor U1006 (N_1006,In_551,In_422);
and U1007 (N_1007,In_715,In_14);
nand U1008 (N_1008,In_940,In_451);
and U1009 (N_1009,In_433,In_602);
and U1010 (N_1010,In_61,In_518);
or U1011 (N_1011,In_433,In_100);
and U1012 (N_1012,In_764,In_538);
or U1013 (N_1013,In_9,In_706);
or U1014 (N_1014,In_936,In_351);
nand U1015 (N_1015,In_904,In_138);
and U1016 (N_1016,In_570,In_137);
or U1017 (N_1017,In_916,In_1);
nand U1018 (N_1018,In_490,In_13);
or U1019 (N_1019,In_997,In_48);
or U1020 (N_1020,In_286,In_833);
nor U1021 (N_1021,In_710,In_489);
nor U1022 (N_1022,In_438,In_830);
and U1023 (N_1023,In_723,In_534);
and U1024 (N_1024,In_73,In_57);
and U1025 (N_1025,In_525,In_378);
or U1026 (N_1026,In_475,In_448);
and U1027 (N_1027,In_281,In_466);
and U1028 (N_1028,In_432,In_813);
and U1029 (N_1029,In_549,In_740);
and U1030 (N_1030,In_206,In_528);
and U1031 (N_1031,In_573,In_463);
or U1032 (N_1032,In_808,In_675);
nand U1033 (N_1033,In_61,In_886);
or U1034 (N_1034,In_816,In_9);
nand U1035 (N_1035,In_85,In_827);
nand U1036 (N_1036,In_574,In_781);
nor U1037 (N_1037,In_964,In_729);
nor U1038 (N_1038,In_186,In_383);
and U1039 (N_1039,In_196,In_122);
or U1040 (N_1040,In_178,In_461);
nand U1041 (N_1041,In_524,In_708);
nand U1042 (N_1042,In_198,In_991);
nor U1043 (N_1043,In_831,In_826);
or U1044 (N_1044,In_109,In_425);
nand U1045 (N_1045,In_91,In_389);
or U1046 (N_1046,In_593,In_995);
or U1047 (N_1047,In_43,In_742);
xnor U1048 (N_1048,In_39,In_796);
and U1049 (N_1049,In_607,In_599);
nor U1050 (N_1050,In_29,In_688);
or U1051 (N_1051,In_233,In_386);
nor U1052 (N_1052,In_900,In_921);
nand U1053 (N_1053,In_880,In_682);
nor U1054 (N_1054,In_798,In_519);
nand U1055 (N_1055,In_221,In_929);
nand U1056 (N_1056,In_194,In_469);
and U1057 (N_1057,In_323,In_557);
nor U1058 (N_1058,In_19,In_192);
and U1059 (N_1059,In_812,In_798);
or U1060 (N_1060,In_667,In_712);
or U1061 (N_1061,In_808,In_879);
or U1062 (N_1062,In_544,In_641);
nand U1063 (N_1063,In_877,In_8);
nand U1064 (N_1064,In_264,In_903);
and U1065 (N_1065,In_13,In_284);
nor U1066 (N_1066,In_410,In_620);
or U1067 (N_1067,In_496,In_735);
nor U1068 (N_1068,In_125,In_1);
or U1069 (N_1069,In_837,In_264);
nor U1070 (N_1070,In_867,In_930);
nand U1071 (N_1071,In_761,In_831);
or U1072 (N_1072,In_607,In_156);
nor U1073 (N_1073,In_551,In_478);
or U1074 (N_1074,In_656,In_744);
nor U1075 (N_1075,In_263,In_343);
and U1076 (N_1076,In_184,In_47);
or U1077 (N_1077,In_297,In_531);
nand U1078 (N_1078,In_799,In_795);
or U1079 (N_1079,In_63,In_544);
nand U1080 (N_1080,In_315,In_217);
and U1081 (N_1081,In_819,In_869);
nor U1082 (N_1082,In_545,In_172);
or U1083 (N_1083,In_668,In_492);
or U1084 (N_1084,In_457,In_966);
nor U1085 (N_1085,In_390,In_10);
and U1086 (N_1086,In_272,In_160);
nor U1087 (N_1087,In_629,In_231);
and U1088 (N_1088,In_233,In_554);
or U1089 (N_1089,In_856,In_909);
nand U1090 (N_1090,In_255,In_553);
or U1091 (N_1091,In_616,In_443);
xor U1092 (N_1092,In_618,In_96);
nand U1093 (N_1093,In_349,In_546);
and U1094 (N_1094,In_360,In_93);
and U1095 (N_1095,In_1,In_667);
or U1096 (N_1096,In_459,In_592);
or U1097 (N_1097,In_450,In_657);
and U1098 (N_1098,In_584,In_10);
and U1099 (N_1099,In_756,In_482);
nand U1100 (N_1100,In_595,In_904);
or U1101 (N_1101,In_396,In_865);
nand U1102 (N_1102,In_436,In_968);
or U1103 (N_1103,In_918,In_875);
nor U1104 (N_1104,In_202,In_212);
and U1105 (N_1105,In_117,In_160);
nand U1106 (N_1106,In_948,In_183);
or U1107 (N_1107,In_269,In_431);
or U1108 (N_1108,In_307,In_585);
or U1109 (N_1109,In_115,In_405);
nand U1110 (N_1110,In_707,In_387);
or U1111 (N_1111,In_956,In_362);
nor U1112 (N_1112,In_115,In_983);
nand U1113 (N_1113,In_188,In_79);
or U1114 (N_1114,In_911,In_626);
or U1115 (N_1115,In_240,In_811);
nand U1116 (N_1116,In_469,In_792);
nand U1117 (N_1117,In_224,In_245);
nand U1118 (N_1118,In_712,In_948);
nor U1119 (N_1119,In_252,In_681);
nand U1120 (N_1120,In_341,In_820);
and U1121 (N_1121,In_750,In_903);
and U1122 (N_1122,In_189,In_253);
nor U1123 (N_1123,In_646,In_197);
nand U1124 (N_1124,In_541,In_613);
xnor U1125 (N_1125,In_800,In_493);
nand U1126 (N_1126,In_264,In_295);
or U1127 (N_1127,In_864,In_42);
nand U1128 (N_1128,In_503,In_183);
nand U1129 (N_1129,In_173,In_905);
nand U1130 (N_1130,In_63,In_563);
nor U1131 (N_1131,In_192,In_276);
and U1132 (N_1132,In_830,In_18);
nand U1133 (N_1133,In_770,In_108);
nand U1134 (N_1134,In_604,In_293);
or U1135 (N_1135,In_933,In_483);
nand U1136 (N_1136,In_868,In_877);
nor U1137 (N_1137,In_509,In_337);
nor U1138 (N_1138,In_222,In_907);
or U1139 (N_1139,In_537,In_554);
nor U1140 (N_1140,In_473,In_495);
nor U1141 (N_1141,In_319,In_607);
and U1142 (N_1142,In_134,In_302);
and U1143 (N_1143,In_927,In_9);
nand U1144 (N_1144,In_675,In_408);
nor U1145 (N_1145,In_578,In_61);
nand U1146 (N_1146,In_6,In_414);
and U1147 (N_1147,In_702,In_378);
or U1148 (N_1148,In_807,In_385);
nor U1149 (N_1149,In_303,In_946);
or U1150 (N_1150,In_112,In_388);
nand U1151 (N_1151,In_721,In_64);
nand U1152 (N_1152,In_782,In_449);
nand U1153 (N_1153,In_5,In_241);
or U1154 (N_1154,In_351,In_492);
or U1155 (N_1155,In_854,In_88);
nand U1156 (N_1156,In_296,In_623);
and U1157 (N_1157,In_923,In_800);
nor U1158 (N_1158,In_761,In_346);
xnor U1159 (N_1159,In_436,In_558);
or U1160 (N_1160,In_430,In_360);
and U1161 (N_1161,In_204,In_211);
nand U1162 (N_1162,In_732,In_570);
nor U1163 (N_1163,In_560,In_977);
nand U1164 (N_1164,In_796,In_136);
or U1165 (N_1165,In_853,In_814);
or U1166 (N_1166,In_250,In_440);
or U1167 (N_1167,In_420,In_822);
nand U1168 (N_1168,In_483,In_959);
nand U1169 (N_1169,In_891,In_309);
nand U1170 (N_1170,In_116,In_135);
nand U1171 (N_1171,In_999,In_409);
nand U1172 (N_1172,In_916,In_658);
nand U1173 (N_1173,In_960,In_288);
nor U1174 (N_1174,In_585,In_394);
nor U1175 (N_1175,In_995,In_304);
nor U1176 (N_1176,In_331,In_498);
nor U1177 (N_1177,In_368,In_936);
and U1178 (N_1178,In_390,In_16);
and U1179 (N_1179,In_232,In_175);
nand U1180 (N_1180,In_916,In_535);
nand U1181 (N_1181,In_59,In_162);
nand U1182 (N_1182,In_417,In_556);
or U1183 (N_1183,In_515,In_617);
and U1184 (N_1184,In_627,In_565);
or U1185 (N_1185,In_551,In_483);
nor U1186 (N_1186,In_91,In_437);
nand U1187 (N_1187,In_380,In_851);
nand U1188 (N_1188,In_142,In_610);
or U1189 (N_1189,In_601,In_788);
or U1190 (N_1190,In_573,In_745);
nand U1191 (N_1191,In_469,In_192);
and U1192 (N_1192,In_853,In_706);
and U1193 (N_1193,In_22,In_182);
nand U1194 (N_1194,In_704,In_268);
nor U1195 (N_1195,In_970,In_903);
and U1196 (N_1196,In_237,In_898);
nand U1197 (N_1197,In_589,In_955);
and U1198 (N_1198,In_643,In_591);
and U1199 (N_1199,In_121,In_797);
nand U1200 (N_1200,In_915,In_525);
nand U1201 (N_1201,In_944,In_295);
nor U1202 (N_1202,In_986,In_284);
nor U1203 (N_1203,In_788,In_896);
and U1204 (N_1204,In_841,In_518);
nand U1205 (N_1205,In_172,In_732);
or U1206 (N_1206,In_937,In_292);
or U1207 (N_1207,In_213,In_304);
nor U1208 (N_1208,In_122,In_329);
and U1209 (N_1209,In_820,In_633);
nor U1210 (N_1210,In_678,In_691);
nor U1211 (N_1211,In_795,In_760);
nor U1212 (N_1212,In_420,In_824);
nor U1213 (N_1213,In_23,In_836);
nand U1214 (N_1214,In_414,In_823);
nor U1215 (N_1215,In_589,In_516);
nor U1216 (N_1216,In_637,In_301);
and U1217 (N_1217,In_618,In_482);
nand U1218 (N_1218,In_711,In_71);
nand U1219 (N_1219,In_667,In_312);
or U1220 (N_1220,In_107,In_101);
or U1221 (N_1221,In_213,In_273);
and U1222 (N_1222,In_406,In_156);
nand U1223 (N_1223,In_894,In_671);
nor U1224 (N_1224,In_648,In_460);
nand U1225 (N_1225,In_188,In_752);
nor U1226 (N_1226,In_83,In_302);
nor U1227 (N_1227,In_511,In_964);
or U1228 (N_1228,In_983,In_938);
or U1229 (N_1229,In_991,In_24);
nand U1230 (N_1230,In_374,In_574);
nor U1231 (N_1231,In_912,In_545);
nor U1232 (N_1232,In_856,In_532);
nor U1233 (N_1233,In_278,In_988);
or U1234 (N_1234,In_342,In_22);
xor U1235 (N_1235,In_293,In_372);
or U1236 (N_1236,In_880,In_100);
nand U1237 (N_1237,In_668,In_199);
nand U1238 (N_1238,In_4,In_112);
nand U1239 (N_1239,In_30,In_7);
and U1240 (N_1240,In_253,In_615);
and U1241 (N_1241,In_299,In_846);
and U1242 (N_1242,In_244,In_769);
or U1243 (N_1243,In_778,In_356);
nor U1244 (N_1244,In_841,In_898);
nand U1245 (N_1245,In_607,In_450);
nor U1246 (N_1246,In_365,In_711);
nor U1247 (N_1247,In_131,In_130);
or U1248 (N_1248,In_782,In_443);
nor U1249 (N_1249,In_218,In_265);
nand U1250 (N_1250,In_394,In_251);
xor U1251 (N_1251,In_188,In_442);
and U1252 (N_1252,In_306,In_28);
and U1253 (N_1253,In_260,In_50);
or U1254 (N_1254,In_562,In_68);
or U1255 (N_1255,In_657,In_302);
nand U1256 (N_1256,In_21,In_753);
nand U1257 (N_1257,In_294,In_703);
or U1258 (N_1258,In_965,In_621);
nand U1259 (N_1259,In_130,In_682);
or U1260 (N_1260,In_907,In_852);
or U1261 (N_1261,In_413,In_919);
and U1262 (N_1262,In_696,In_185);
nor U1263 (N_1263,In_408,In_363);
nor U1264 (N_1264,In_352,In_968);
nor U1265 (N_1265,In_274,In_288);
or U1266 (N_1266,In_167,In_606);
and U1267 (N_1267,In_796,In_212);
nand U1268 (N_1268,In_43,In_123);
or U1269 (N_1269,In_502,In_960);
nor U1270 (N_1270,In_600,In_295);
and U1271 (N_1271,In_876,In_471);
and U1272 (N_1272,In_981,In_185);
and U1273 (N_1273,In_514,In_595);
nor U1274 (N_1274,In_483,In_634);
and U1275 (N_1275,In_247,In_392);
nor U1276 (N_1276,In_232,In_234);
nand U1277 (N_1277,In_947,In_584);
or U1278 (N_1278,In_52,In_427);
nor U1279 (N_1279,In_741,In_346);
or U1280 (N_1280,In_918,In_213);
and U1281 (N_1281,In_125,In_117);
and U1282 (N_1282,In_282,In_734);
and U1283 (N_1283,In_288,In_53);
or U1284 (N_1284,In_421,In_422);
or U1285 (N_1285,In_87,In_635);
and U1286 (N_1286,In_573,In_32);
nand U1287 (N_1287,In_13,In_955);
or U1288 (N_1288,In_714,In_710);
nor U1289 (N_1289,In_599,In_592);
nor U1290 (N_1290,In_886,In_415);
nand U1291 (N_1291,In_815,In_3);
nand U1292 (N_1292,In_416,In_298);
nor U1293 (N_1293,In_536,In_151);
or U1294 (N_1294,In_746,In_739);
nand U1295 (N_1295,In_934,In_172);
or U1296 (N_1296,In_565,In_360);
and U1297 (N_1297,In_896,In_466);
nand U1298 (N_1298,In_760,In_583);
nor U1299 (N_1299,In_77,In_560);
nor U1300 (N_1300,In_930,In_234);
nor U1301 (N_1301,In_822,In_34);
nor U1302 (N_1302,In_302,In_242);
and U1303 (N_1303,In_563,In_327);
nor U1304 (N_1304,In_910,In_974);
nand U1305 (N_1305,In_257,In_575);
or U1306 (N_1306,In_89,In_264);
nor U1307 (N_1307,In_683,In_386);
nor U1308 (N_1308,In_714,In_566);
and U1309 (N_1309,In_683,In_595);
nand U1310 (N_1310,In_490,In_52);
and U1311 (N_1311,In_219,In_55);
nor U1312 (N_1312,In_828,In_689);
nor U1313 (N_1313,In_81,In_98);
and U1314 (N_1314,In_267,In_136);
or U1315 (N_1315,In_12,In_127);
and U1316 (N_1316,In_439,In_665);
nand U1317 (N_1317,In_27,In_532);
or U1318 (N_1318,In_835,In_162);
or U1319 (N_1319,In_361,In_772);
xnor U1320 (N_1320,In_362,In_367);
nand U1321 (N_1321,In_917,In_204);
and U1322 (N_1322,In_990,In_679);
or U1323 (N_1323,In_809,In_784);
and U1324 (N_1324,In_816,In_428);
or U1325 (N_1325,In_921,In_824);
nand U1326 (N_1326,In_88,In_471);
nand U1327 (N_1327,In_839,In_473);
nor U1328 (N_1328,In_57,In_831);
and U1329 (N_1329,In_753,In_655);
nand U1330 (N_1330,In_43,In_319);
and U1331 (N_1331,In_177,In_705);
xnor U1332 (N_1332,In_849,In_20);
nand U1333 (N_1333,In_180,In_797);
nor U1334 (N_1334,In_803,In_595);
nand U1335 (N_1335,In_411,In_602);
nand U1336 (N_1336,In_572,In_656);
or U1337 (N_1337,In_381,In_493);
nand U1338 (N_1338,In_197,In_61);
nor U1339 (N_1339,In_572,In_647);
and U1340 (N_1340,In_131,In_793);
nor U1341 (N_1341,In_653,In_275);
nand U1342 (N_1342,In_234,In_483);
nor U1343 (N_1343,In_541,In_800);
or U1344 (N_1344,In_151,In_496);
nand U1345 (N_1345,In_376,In_250);
or U1346 (N_1346,In_406,In_976);
nor U1347 (N_1347,In_915,In_766);
and U1348 (N_1348,In_193,In_397);
or U1349 (N_1349,In_513,In_808);
or U1350 (N_1350,In_795,In_875);
or U1351 (N_1351,In_79,In_602);
and U1352 (N_1352,In_79,In_252);
and U1353 (N_1353,In_880,In_937);
and U1354 (N_1354,In_322,In_202);
or U1355 (N_1355,In_530,In_423);
nand U1356 (N_1356,In_290,In_261);
nor U1357 (N_1357,In_924,In_665);
and U1358 (N_1358,In_146,In_485);
nor U1359 (N_1359,In_937,In_129);
or U1360 (N_1360,In_178,In_115);
and U1361 (N_1361,In_762,In_804);
and U1362 (N_1362,In_793,In_557);
nor U1363 (N_1363,In_217,In_584);
and U1364 (N_1364,In_469,In_979);
or U1365 (N_1365,In_281,In_114);
and U1366 (N_1366,In_369,In_692);
nor U1367 (N_1367,In_126,In_46);
and U1368 (N_1368,In_182,In_647);
and U1369 (N_1369,In_789,In_143);
nor U1370 (N_1370,In_191,In_603);
nand U1371 (N_1371,In_51,In_632);
nand U1372 (N_1372,In_735,In_838);
nand U1373 (N_1373,In_66,In_488);
or U1374 (N_1374,In_371,In_39);
nand U1375 (N_1375,In_888,In_988);
and U1376 (N_1376,In_550,In_799);
and U1377 (N_1377,In_135,In_992);
or U1378 (N_1378,In_237,In_416);
and U1379 (N_1379,In_5,In_410);
or U1380 (N_1380,In_431,In_295);
and U1381 (N_1381,In_512,In_147);
nand U1382 (N_1382,In_651,In_54);
nand U1383 (N_1383,In_688,In_541);
nor U1384 (N_1384,In_11,In_466);
nand U1385 (N_1385,In_467,In_460);
nand U1386 (N_1386,In_524,In_281);
nand U1387 (N_1387,In_492,In_684);
nor U1388 (N_1388,In_204,In_602);
nand U1389 (N_1389,In_896,In_464);
or U1390 (N_1390,In_12,In_478);
nand U1391 (N_1391,In_415,In_813);
nand U1392 (N_1392,In_819,In_199);
nor U1393 (N_1393,In_630,In_159);
nand U1394 (N_1394,In_545,In_737);
nand U1395 (N_1395,In_478,In_864);
and U1396 (N_1396,In_808,In_141);
or U1397 (N_1397,In_687,In_427);
nor U1398 (N_1398,In_444,In_840);
nand U1399 (N_1399,In_722,In_729);
nand U1400 (N_1400,In_481,In_789);
and U1401 (N_1401,In_194,In_375);
or U1402 (N_1402,In_752,In_910);
and U1403 (N_1403,In_466,In_606);
or U1404 (N_1404,In_789,In_872);
and U1405 (N_1405,In_520,In_62);
nand U1406 (N_1406,In_408,In_32);
nand U1407 (N_1407,In_282,In_847);
nand U1408 (N_1408,In_273,In_707);
and U1409 (N_1409,In_692,In_539);
and U1410 (N_1410,In_285,In_402);
and U1411 (N_1411,In_163,In_7);
and U1412 (N_1412,In_959,In_663);
and U1413 (N_1413,In_555,In_895);
nand U1414 (N_1414,In_542,In_613);
nand U1415 (N_1415,In_812,In_166);
and U1416 (N_1416,In_194,In_537);
or U1417 (N_1417,In_361,In_826);
nand U1418 (N_1418,In_786,In_942);
nor U1419 (N_1419,In_919,In_448);
nor U1420 (N_1420,In_759,In_815);
or U1421 (N_1421,In_722,In_513);
nor U1422 (N_1422,In_974,In_52);
nand U1423 (N_1423,In_708,In_96);
nor U1424 (N_1424,In_810,In_76);
nor U1425 (N_1425,In_651,In_241);
and U1426 (N_1426,In_999,In_150);
nand U1427 (N_1427,In_725,In_578);
or U1428 (N_1428,In_718,In_767);
or U1429 (N_1429,In_974,In_939);
and U1430 (N_1430,In_329,In_774);
nor U1431 (N_1431,In_600,In_604);
and U1432 (N_1432,In_771,In_233);
nand U1433 (N_1433,In_157,In_674);
and U1434 (N_1434,In_184,In_853);
and U1435 (N_1435,In_190,In_97);
nand U1436 (N_1436,In_116,In_527);
or U1437 (N_1437,In_925,In_997);
and U1438 (N_1438,In_305,In_284);
nand U1439 (N_1439,In_98,In_877);
nor U1440 (N_1440,In_755,In_65);
nor U1441 (N_1441,In_357,In_282);
or U1442 (N_1442,In_258,In_240);
nand U1443 (N_1443,In_99,In_602);
nand U1444 (N_1444,In_649,In_610);
and U1445 (N_1445,In_26,In_207);
nand U1446 (N_1446,In_577,In_869);
nor U1447 (N_1447,In_73,In_860);
nand U1448 (N_1448,In_873,In_173);
or U1449 (N_1449,In_857,In_179);
or U1450 (N_1450,In_671,In_365);
nand U1451 (N_1451,In_337,In_911);
nand U1452 (N_1452,In_586,In_897);
nor U1453 (N_1453,In_928,In_191);
nor U1454 (N_1454,In_934,In_569);
or U1455 (N_1455,In_361,In_217);
nor U1456 (N_1456,In_179,In_538);
and U1457 (N_1457,In_604,In_668);
or U1458 (N_1458,In_193,In_970);
nor U1459 (N_1459,In_28,In_417);
and U1460 (N_1460,In_900,In_569);
nand U1461 (N_1461,In_101,In_451);
nor U1462 (N_1462,In_461,In_384);
or U1463 (N_1463,In_233,In_986);
nor U1464 (N_1464,In_723,In_748);
or U1465 (N_1465,In_35,In_120);
or U1466 (N_1466,In_648,In_332);
nand U1467 (N_1467,In_836,In_357);
and U1468 (N_1468,In_549,In_4);
nor U1469 (N_1469,In_749,In_603);
nand U1470 (N_1470,In_283,In_330);
and U1471 (N_1471,In_16,In_557);
nand U1472 (N_1472,In_357,In_661);
nand U1473 (N_1473,In_825,In_931);
nand U1474 (N_1474,In_43,In_135);
nor U1475 (N_1475,In_939,In_850);
nand U1476 (N_1476,In_877,In_594);
or U1477 (N_1477,In_607,In_103);
or U1478 (N_1478,In_636,In_286);
nand U1479 (N_1479,In_36,In_30);
nor U1480 (N_1480,In_390,In_481);
nor U1481 (N_1481,In_869,In_699);
and U1482 (N_1482,In_107,In_159);
or U1483 (N_1483,In_462,In_94);
and U1484 (N_1484,In_636,In_897);
and U1485 (N_1485,In_247,In_832);
and U1486 (N_1486,In_767,In_220);
and U1487 (N_1487,In_208,In_682);
nand U1488 (N_1488,In_825,In_612);
and U1489 (N_1489,In_530,In_350);
nor U1490 (N_1490,In_641,In_686);
or U1491 (N_1491,In_960,In_605);
nand U1492 (N_1492,In_445,In_683);
nor U1493 (N_1493,In_756,In_626);
or U1494 (N_1494,In_936,In_815);
and U1495 (N_1495,In_969,In_764);
nand U1496 (N_1496,In_490,In_6);
or U1497 (N_1497,In_902,In_398);
and U1498 (N_1498,In_745,In_845);
nor U1499 (N_1499,In_619,In_525);
nor U1500 (N_1500,In_541,In_525);
or U1501 (N_1501,In_102,In_942);
nand U1502 (N_1502,In_386,In_505);
or U1503 (N_1503,In_190,In_654);
and U1504 (N_1504,In_835,In_530);
or U1505 (N_1505,In_458,In_192);
nor U1506 (N_1506,In_759,In_764);
or U1507 (N_1507,In_69,In_173);
and U1508 (N_1508,In_469,In_429);
or U1509 (N_1509,In_124,In_119);
and U1510 (N_1510,In_839,In_221);
nand U1511 (N_1511,In_164,In_317);
and U1512 (N_1512,In_402,In_843);
nor U1513 (N_1513,In_732,In_760);
or U1514 (N_1514,In_136,In_186);
nand U1515 (N_1515,In_933,In_418);
nor U1516 (N_1516,In_970,In_786);
and U1517 (N_1517,In_554,In_672);
xor U1518 (N_1518,In_500,In_603);
nor U1519 (N_1519,In_15,In_275);
nand U1520 (N_1520,In_532,In_599);
or U1521 (N_1521,In_308,In_725);
nand U1522 (N_1522,In_14,In_382);
and U1523 (N_1523,In_210,In_176);
nand U1524 (N_1524,In_822,In_51);
and U1525 (N_1525,In_990,In_611);
nand U1526 (N_1526,In_171,In_133);
nor U1527 (N_1527,In_474,In_632);
and U1528 (N_1528,In_37,In_210);
and U1529 (N_1529,In_214,In_27);
or U1530 (N_1530,In_588,In_858);
and U1531 (N_1531,In_835,In_245);
nand U1532 (N_1532,In_337,In_831);
and U1533 (N_1533,In_288,In_591);
or U1534 (N_1534,In_738,In_914);
nor U1535 (N_1535,In_591,In_395);
nor U1536 (N_1536,In_267,In_765);
or U1537 (N_1537,In_126,In_26);
and U1538 (N_1538,In_573,In_358);
or U1539 (N_1539,In_884,In_998);
or U1540 (N_1540,In_47,In_517);
and U1541 (N_1541,In_81,In_188);
or U1542 (N_1542,In_860,In_163);
nand U1543 (N_1543,In_444,In_233);
or U1544 (N_1544,In_573,In_101);
nor U1545 (N_1545,In_582,In_197);
nor U1546 (N_1546,In_946,In_206);
or U1547 (N_1547,In_437,In_970);
nand U1548 (N_1548,In_620,In_865);
or U1549 (N_1549,In_338,In_508);
nor U1550 (N_1550,In_234,In_271);
or U1551 (N_1551,In_297,In_701);
and U1552 (N_1552,In_30,In_671);
or U1553 (N_1553,In_148,In_413);
and U1554 (N_1554,In_729,In_239);
nor U1555 (N_1555,In_246,In_996);
nor U1556 (N_1556,In_848,In_605);
nor U1557 (N_1557,In_676,In_503);
nand U1558 (N_1558,In_4,In_865);
or U1559 (N_1559,In_741,In_127);
or U1560 (N_1560,In_317,In_74);
nand U1561 (N_1561,In_137,In_794);
or U1562 (N_1562,In_175,In_52);
nand U1563 (N_1563,In_422,In_711);
nor U1564 (N_1564,In_95,In_143);
nand U1565 (N_1565,In_361,In_878);
or U1566 (N_1566,In_684,In_848);
nor U1567 (N_1567,In_970,In_164);
nand U1568 (N_1568,In_198,In_606);
nand U1569 (N_1569,In_889,In_259);
or U1570 (N_1570,In_908,In_400);
nand U1571 (N_1571,In_315,In_459);
nor U1572 (N_1572,In_313,In_414);
nand U1573 (N_1573,In_407,In_280);
and U1574 (N_1574,In_479,In_278);
or U1575 (N_1575,In_504,In_35);
nand U1576 (N_1576,In_494,In_233);
or U1577 (N_1577,In_350,In_51);
nor U1578 (N_1578,In_96,In_496);
nand U1579 (N_1579,In_633,In_631);
nor U1580 (N_1580,In_223,In_980);
or U1581 (N_1581,In_773,In_248);
nor U1582 (N_1582,In_971,In_294);
and U1583 (N_1583,In_371,In_719);
and U1584 (N_1584,In_857,In_81);
or U1585 (N_1585,In_303,In_433);
or U1586 (N_1586,In_531,In_126);
and U1587 (N_1587,In_929,In_398);
nand U1588 (N_1588,In_518,In_146);
and U1589 (N_1589,In_197,In_319);
or U1590 (N_1590,In_652,In_430);
or U1591 (N_1591,In_909,In_592);
nand U1592 (N_1592,In_56,In_684);
nand U1593 (N_1593,In_330,In_781);
or U1594 (N_1594,In_553,In_589);
and U1595 (N_1595,In_780,In_540);
and U1596 (N_1596,In_380,In_207);
or U1597 (N_1597,In_827,In_191);
nand U1598 (N_1598,In_801,In_614);
nand U1599 (N_1599,In_583,In_40);
nand U1600 (N_1600,In_682,In_367);
or U1601 (N_1601,In_279,In_494);
and U1602 (N_1602,In_141,In_136);
or U1603 (N_1603,In_961,In_165);
or U1604 (N_1604,In_155,In_721);
nor U1605 (N_1605,In_985,In_464);
and U1606 (N_1606,In_882,In_613);
or U1607 (N_1607,In_989,In_617);
or U1608 (N_1608,In_131,In_984);
nor U1609 (N_1609,In_0,In_788);
and U1610 (N_1610,In_407,In_118);
nor U1611 (N_1611,In_896,In_909);
nand U1612 (N_1612,In_902,In_756);
nor U1613 (N_1613,In_356,In_386);
nor U1614 (N_1614,In_331,In_773);
and U1615 (N_1615,In_764,In_913);
or U1616 (N_1616,In_534,In_703);
and U1617 (N_1617,In_998,In_951);
nand U1618 (N_1618,In_731,In_849);
nor U1619 (N_1619,In_424,In_126);
nand U1620 (N_1620,In_552,In_857);
nand U1621 (N_1621,In_886,In_970);
nor U1622 (N_1622,In_475,In_559);
and U1623 (N_1623,In_151,In_825);
nand U1624 (N_1624,In_524,In_707);
nor U1625 (N_1625,In_208,In_252);
nor U1626 (N_1626,In_743,In_774);
nand U1627 (N_1627,In_716,In_629);
nand U1628 (N_1628,In_700,In_878);
nand U1629 (N_1629,In_159,In_725);
nor U1630 (N_1630,In_235,In_307);
nand U1631 (N_1631,In_316,In_883);
and U1632 (N_1632,In_659,In_277);
nand U1633 (N_1633,In_479,In_305);
nand U1634 (N_1634,In_421,In_625);
and U1635 (N_1635,In_776,In_664);
nor U1636 (N_1636,In_352,In_330);
or U1637 (N_1637,In_377,In_964);
nand U1638 (N_1638,In_993,In_856);
or U1639 (N_1639,In_444,In_388);
nand U1640 (N_1640,In_659,In_750);
or U1641 (N_1641,In_261,In_505);
nand U1642 (N_1642,In_526,In_48);
or U1643 (N_1643,In_745,In_973);
or U1644 (N_1644,In_296,In_631);
and U1645 (N_1645,In_812,In_389);
or U1646 (N_1646,In_569,In_996);
nand U1647 (N_1647,In_706,In_820);
nor U1648 (N_1648,In_511,In_419);
or U1649 (N_1649,In_672,In_1);
or U1650 (N_1650,In_176,In_292);
and U1651 (N_1651,In_519,In_408);
and U1652 (N_1652,In_307,In_601);
or U1653 (N_1653,In_192,In_788);
nor U1654 (N_1654,In_694,In_727);
and U1655 (N_1655,In_853,In_985);
xor U1656 (N_1656,In_22,In_978);
and U1657 (N_1657,In_275,In_600);
and U1658 (N_1658,In_629,In_555);
nand U1659 (N_1659,In_443,In_359);
nor U1660 (N_1660,In_271,In_42);
or U1661 (N_1661,In_570,In_637);
nor U1662 (N_1662,In_812,In_813);
nand U1663 (N_1663,In_612,In_655);
and U1664 (N_1664,In_516,In_464);
nand U1665 (N_1665,In_392,In_630);
or U1666 (N_1666,In_265,In_128);
or U1667 (N_1667,In_689,In_698);
or U1668 (N_1668,In_606,In_827);
nor U1669 (N_1669,In_884,In_851);
xor U1670 (N_1670,In_60,In_690);
nor U1671 (N_1671,In_513,In_889);
or U1672 (N_1672,In_914,In_276);
xnor U1673 (N_1673,In_43,In_124);
and U1674 (N_1674,In_966,In_373);
and U1675 (N_1675,In_617,In_110);
and U1676 (N_1676,In_307,In_336);
and U1677 (N_1677,In_639,In_314);
or U1678 (N_1678,In_636,In_402);
nor U1679 (N_1679,In_90,In_671);
nor U1680 (N_1680,In_744,In_497);
nand U1681 (N_1681,In_760,In_445);
nand U1682 (N_1682,In_990,In_517);
and U1683 (N_1683,In_233,In_369);
or U1684 (N_1684,In_990,In_540);
and U1685 (N_1685,In_68,In_347);
nand U1686 (N_1686,In_892,In_268);
nand U1687 (N_1687,In_979,In_472);
nor U1688 (N_1688,In_884,In_109);
and U1689 (N_1689,In_183,In_317);
or U1690 (N_1690,In_834,In_527);
nor U1691 (N_1691,In_268,In_12);
or U1692 (N_1692,In_537,In_730);
nand U1693 (N_1693,In_106,In_797);
and U1694 (N_1694,In_363,In_355);
nor U1695 (N_1695,In_36,In_534);
or U1696 (N_1696,In_369,In_640);
and U1697 (N_1697,In_113,In_511);
or U1698 (N_1698,In_821,In_673);
and U1699 (N_1699,In_171,In_261);
nor U1700 (N_1700,In_566,In_771);
and U1701 (N_1701,In_63,In_156);
nand U1702 (N_1702,In_873,In_351);
nor U1703 (N_1703,In_108,In_806);
nor U1704 (N_1704,In_141,In_348);
and U1705 (N_1705,In_323,In_836);
and U1706 (N_1706,In_695,In_51);
or U1707 (N_1707,In_481,In_238);
nand U1708 (N_1708,In_909,In_681);
and U1709 (N_1709,In_120,In_411);
and U1710 (N_1710,In_868,In_126);
nand U1711 (N_1711,In_562,In_812);
or U1712 (N_1712,In_307,In_846);
nor U1713 (N_1713,In_14,In_966);
and U1714 (N_1714,In_575,In_14);
nand U1715 (N_1715,In_454,In_39);
or U1716 (N_1716,In_392,In_939);
nand U1717 (N_1717,In_110,In_587);
nor U1718 (N_1718,In_458,In_556);
and U1719 (N_1719,In_788,In_759);
nand U1720 (N_1720,In_836,In_2);
nand U1721 (N_1721,In_966,In_290);
and U1722 (N_1722,In_848,In_246);
or U1723 (N_1723,In_441,In_266);
nor U1724 (N_1724,In_291,In_288);
or U1725 (N_1725,In_735,In_102);
or U1726 (N_1726,In_276,In_560);
and U1727 (N_1727,In_349,In_797);
or U1728 (N_1728,In_704,In_791);
and U1729 (N_1729,In_100,In_667);
or U1730 (N_1730,In_579,In_240);
nor U1731 (N_1731,In_294,In_694);
nor U1732 (N_1732,In_525,In_544);
nand U1733 (N_1733,In_476,In_282);
and U1734 (N_1734,In_922,In_635);
or U1735 (N_1735,In_187,In_93);
xnor U1736 (N_1736,In_446,In_784);
nand U1737 (N_1737,In_703,In_347);
and U1738 (N_1738,In_213,In_951);
and U1739 (N_1739,In_504,In_32);
nand U1740 (N_1740,In_668,In_846);
nand U1741 (N_1741,In_407,In_675);
nor U1742 (N_1742,In_266,In_912);
nor U1743 (N_1743,In_754,In_529);
or U1744 (N_1744,In_335,In_817);
nand U1745 (N_1745,In_3,In_602);
or U1746 (N_1746,In_420,In_108);
and U1747 (N_1747,In_390,In_274);
or U1748 (N_1748,In_906,In_186);
nand U1749 (N_1749,In_438,In_615);
nand U1750 (N_1750,In_837,In_842);
nor U1751 (N_1751,In_306,In_938);
nor U1752 (N_1752,In_690,In_733);
nand U1753 (N_1753,In_48,In_967);
nand U1754 (N_1754,In_986,In_854);
nand U1755 (N_1755,In_685,In_339);
nand U1756 (N_1756,In_784,In_609);
nand U1757 (N_1757,In_601,In_450);
nor U1758 (N_1758,In_167,In_481);
or U1759 (N_1759,In_819,In_58);
or U1760 (N_1760,In_608,In_31);
and U1761 (N_1761,In_715,In_642);
and U1762 (N_1762,In_132,In_226);
and U1763 (N_1763,In_283,In_647);
nor U1764 (N_1764,In_221,In_838);
and U1765 (N_1765,In_212,In_160);
or U1766 (N_1766,In_225,In_311);
nand U1767 (N_1767,In_840,In_438);
nand U1768 (N_1768,In_219,In_966);
nor U1769 (N_1769,In_702,In_81);
or U1770 (N_1770,In_351,In_484);
and U1771 (N_1771,In_75,In_875);
nand U1772 (N_1772,In_624,In_804);
nor U1773 (N_1773,In_441,In_200);
and U1774 (N_1774,In_153,In_405);
nand U1775 (N_1775,In_785,In_932);
nor U1776 (N_1776,In_159,In_763);
and U1777 (N_1777,In_477,In_33);
and U1778 (N_1778,In_564,In_808);
or U1779 (N_1779,In_887,In_769);
and U1780 (N_1780,In_86,In_883);
and U1781 (N_1781,In_832,In_825);
nor U1782 (N_1782,In_976,In_657);
or U1783 (N_1783,In_734,In_310);
nor U1784 (N_1784,In_129,In_811);
and U1785 (N_1785,In_278,In_643);
and U1786 (N_1786,In_43,In_355);
or U1787 (N_1787,In_394,In_756);
or U1788 (N_1788,In_955,In_370);
nand U1789 (N_1789,In_853,In_710);
nor U1790 (N_1790,In_340,In_961);
and U1791 (N_1791,In_658,In_239);
or U1792 (N_1792,In_222,In_60);
and U1793 (N_1793,In_592,In_966);
and U1794 (N_1794,In_358,In_987);
or U1795 (N_1795,In_193,In_111);
or U1796 (N_1796,In_584,In_158);
nor U1797 (N_1797,In_720,In_876);
and U1798 (N_1798,In_858,In_641);
nor U1799 (N_1799,In_773,In_226);
xor U1800 (N_1800,In_278,In_813);
xor U1801 (N_1801,In_120,In_732);
nand U1802 (N_1802,In_609,In_854);
nand U1803 (N_1803,In_763,In_971);
nand U1804 (N_1804,In_8,In_924);
or U1805 (N_1805,In_260,In_244);
or U1806 (N_1806,In_587,In_987);
nor U1807 (N_1807,In_835,In_800);
nor U1808 (N_1808,In_421,In_636);
nand U1809 (N_1809,In_16,In_78);
nor U1810 (N_1810,In_695,In_371);
nor U1811 (N_1811,In_134,In_18);
nand U1812 (N_1812,In_539,In_725);
and U1813 (N_1813,In_986,In_832);
or U1814 (N_1814,In_555,In_259);
nor U1815 (N_1815,In_843,In_405);
xor U1816 (N_1816,In_111,In_130);
and U1817 (N_1817,In_686,In_79);
nor U1818 (N_1818,In_440,In_146);
nand U1819 (N_1819,In_636,In_68);
nor U1820 (N_1820,In_574,In_854);
or U1821 (N_1821,In_411,In_264);
nor U1822 (N_1822,In_649,In_163);
nor U1823 (N_1823,In_715,In_613);
nand U1824 (N_1824,In_961,In_150);
nand U1825 (N_1825,In_538,In_401);
nand U1826 (N_1826,In_701,In_393);
nor U1827 (N_1827,In_39,In_198);
and U1828 (N_1828,In_279,In_954);
and U1829 (N_1829,In_665,In_605);
nor U1830 (N_1830,In_335,In_488);
nor U1831 (N_1831,In_764,In_287);
nor U1832 (N_1832,In_919,In_488);
nor U1833 (N_1833,In_194,In_458);
and U1834 (N_1834,In_365,In_72);
and U1835 (N_1835,In_828,In_152);
and U1836 (N_1836,In_473,In_92);
and U1837 (N_1837,In_477,In_947);
nor U1838 (N_1838,In_396,In_211);
and U1839 (N_1839,In_275,In_389);
or U1840 (N_1840,In_68,In_696);
or U1841 (N_1841,In_702,In_642);
or U1842 (N_1842,In_145,In_572);
nand U1843 (N_1843,In_695,In_937);
nand U1844 (N_1844,In_302,In_606);
nand U1845 (N_1845,In_582,In_471);
or U1846 (N_1846,In_771,In_523);
nand U1847 (N_1847,In_494,In_820);
and U1848 (N_1848,In_860,In_883);
or U1849 (N_1849,In_164,In_582);
nand U1850 (N_1850,In_241,In_883);
nand U1851 (N_1851,In_998,In_217);
and U1852 (N_1852,In_278,In_704);
nor U1853 (N_1853,In_537,In_772);
and U1854 (N_1854,In_849,In_500);
or U1855 (N_1855,In_181,In_192);
nor U1856 (N_1856,In_44,In_239);
and U1857 (N_1857,In_365,In_381);
or U1858 (N_1858,In_1,In_33);
nand U1859 (N_1859,In_876,In_590);
and U1860 (N_1860,In_117,In_394);
nor U1861 (N_1861,In_449,In_304);
and U1862 (N_1862,In_920,In_717);
and U1863 (N_1863,In_814,In_548);
or U1864 (N_1864,In_908,In_615);
nor U1865 (N_1865,In_784,In_751);
nor U1866 (N_1866,In_710,In_961);
nand U1867 (N_1867,In_414,In_830);
or U1868 (N_1868,In_734,In_399);
and U1869 (N_1869,In_101,In_18);
nor U1870 (N_1870,In_28,In_725);
or U1871 (N_1871,In_395,In_797);
and U1872 (N_1872,In_450,In_445);
or U1873 (N_1873,In_511,In_711);
nor U1874 (N_1874,In_924,In_257);
or U1875 (N_1875,In_473,In_22);
nand U1876 (N_1876,In_646,In_880);
or U1877 (N_1877,In_711,In_391);
and U1878 (N_1878,In_640,In_777);
and U1879 (N_1879,In_905,In_682);
nor U1880 (N_1880,In_9,In_803);
nor U1881 (N_1881,In_793,In_341);
or U1882 (N_1882,In_95,In_483);
and U1883 (N_1883,In_567,In_614);
and U1884 (N_1884,In_234,In_633);
or U1885 (N_1885,In_745,In_358);
nand U1886 (N_1886,In_635,In_279);
nand U1887 (N_1887,In_330,In_567);
or U1888 (N_1888,In_44,In_64);
and U1889 (N_1889,In_122,In_15);
nand U1890 (N_1890,In_750,In_332);
nor U1891 (N_1891,In_374,In_31);
nand U1892 (N_1892,In_309,In_991);
or U1893 (N_1893,In_923,In_489);
nor U1894 (N_1894,In_430,In_697);
nor U1895 (N_1895,In_338,In_128);
nor U1896 (N_1896,In_957,In_406);
nor U1897 (N_1897,In_646,In_244);
nor U1898 (N_1898,In_449,In_485);
or U1899 (N_1899,In_621,In_112);
and U1900 (N_1900,In_455,In_37);
and U1901 (N_1901,In_915,In_483);
or U1902 (N_1902,In_886,In_494);
or U1903 (N_1903,In_794,In_660);
nor U1904 (N_1904,In_981,In_783);
nand U1905 (N_1905,In_88,In_695);
and U1906 (N_1906,In_771,In_398);
and U1907 (N_1907,In_993,In_466);
and U1908 (N_1908,In_289,In_614);
and U1909 (N_1909,In_745,In_105);
and U1910 (N_1910,In_292,In_915);
nor U1911 (N_1911,In_505,In_319);
or U1912 (N_1912,In_158,In_732);
nor U1913 (N_1913,In_424,In_482);
nand U1914 (N_1914,In_816,In_963);
nand U1915 (N_1915,In_428,In_732);
nand U1916 (N_1916,In_789,In_920);
nor U1917 (N_1917,In_986,In_595);
nand U1918 (N_1918,In_874,In_582);
nor U1919 (N_1919,In_638,In_137);
nor U1920 (N_1920,In_497,In_54);
nand U1921 (N_1921,In_139,In_163);
or U1922 (N_1922,In_892,In_117);
and U1923 (N_1923,In_956,In_811);
or U1924 (N_1924,In_897,In_130);
or U1925 (N_1925,In_710,In_361);
nand U1926 (N_1926,In_935,In_508);
nand U1927 (N_1927,In_100,In_422);
nand U1928 (N_1928,In_397,In_872);
nor U1929 (N_1929,In_356,In_518);
and U1930 (N_1930,In_455,In_459);
and U1931 (N_1931,In_642,In_927);
or U1932 (N_1932,In_22,In_325);
nand U1933 (N_1933,In_934,In_161);
or U1934 (N_1934,In_730,In_331);
nor U1935 (N_1935,In_682,In_971);
nor U1936 (N_1936,In_114,In_713);
nor U1937 (N_1937,In_93,In_515);
or U1938 (N_1938,In_321,In_170);
or U1939 (N_1939,In_835,In_684);
nand U1940 (N_1940,In_159,In_973);
and U1941 (N_1941,In_1,In_591);
or U1942 (N_1942,In_167,In_349);
or U1943 (N_1943,In_526,In_490);
and U1944 (N_1944,In_752,In_574);
and U1945 (N_1945,In_901,In_458);
and U1946 (N_1946,In_372,In_73);
and U1947 (N_1947,In_219,In_673);
nor U1948 (N_1948,In_526,In_703);
or U1949 (N_1949,In_526,In_843);
nor U1950 (N_1950,In_988,In_417);
or U1951 (N_1951,In_385,In_73);
nand U1952 (N_1952,In_319,In_764);
nor U1953 (N_1953,In_399,In_659);
nand U1954 (N_1954,In_855,In_171);
nor U1955 (N_1955,In_384,In_767);
xor U1956 (N_1956,In_233,In_701);
and U1957 (N_1957,In_99,In_806);
nor U1958 (N_1958,In_138,In_982);
nand U1959 (N_1959,In_931,In_102);
nand U1960 (N_1960,In_511,In_968);
nand U1961 (N_1961,In_985,In_163);
nor U1962 (N_1962,In_637,In_776);
or U1963 (N_1963,In_980,In_5);
or U1964 (N_1964,In_100,In_747);
or U1965 (N_1965,In_176,In_402);
nor U1966 (N_1966,In_766,In_155);
or U1967 (N_1967,In_909,In_472);
or U1968 (N_1968,In_811,In_607);
and U1969 (N_1969,In_283,In_474);
and U1970 (N_1970,In_230,In_463);
or U1971 (N_1971,In_548,In_936);
or U1972 (N_1972,In_128,In_48);
and U1973 (N_1973,In_30,In_837);
or U1974 (N_1974,In_752,In_502);
and U1975 (N_1975,In_725,In_635);
nor U1976 (N_1976,In_799,In_692);
and U1977 (N_1977,In_945,In_782);
nor U1978 (N_1978,In_322,In_653);
nor U1979 (N_1979,In_50,In_425);
and U1980 (N_1980,In_385,In_357);
nor U1981 (N_1981,In_709,In_673);
nand U1982 (N_1982,In_805,In_134);
nor U1983 (N_1983,In_734,In_107);
or U1984 (N_1984,In_442,In_5);
nand U1985 (N_1985,In_175,In_177);
and U1986 (N_1986,In_454,In_940);
nor U1987 (N_1987,In_49,In_162);
nor U1988 (N_1988,In_125,In_176);
nand U1989 (N_1989,In_543,In_316);
and U1990 (N_1990,In_68,In_71);
and U1991 (N_1991,In_15,In_786);
and U1992 (N_1992,In_958,In_779);
and U1993 (N_1993,In_768,In_332);
or U1994 (N_1994,In_333,In_974);
nor U1995 (N_1995,In_372,In_507);
or U1996 (N_1996,In_508,In_977);
or U1997 (N_1997,In_457,In_563);
nor U1998 (N_1998,In_735,In_633);
and U1999 (N_1999,In_722,In_288);
and U2000 (N_2000,In_861,In_433);
nand U2001 (N_2001,In_716,In_78);
and U2002 (N_2002,In_269,In_52);
nand U2003 (N_2003,In_610,In_592);
and U2004 (N_2004,In_63,In_938);
nand U2005 (N_2005,In_151,In_398);
nor U2006 (N_2006,In_327,In_366);
or U2007 (N_2007,In_962,In_509);
or U2008 (N_2008,In_683,In_724);
nand U2009 (N_2009,In_905,In_404);
or U2010 (N_2010,In_179,In_739);
nand U2011 (N_2011,In_695,In_933);
nand U2012 (N_2012,In_818,In_124);
nor U2013 (N_2013,In_712,In_242);
nor U2014 (N_2014,In_405,In_462);
or U2015 (N_2015,In_825,In_707);
or U2016 (N_2016,In_802,In_529);
nor U2017 (N_2017,In_760,In_352);
nor U2018 (N_2018,In_299,In_581);
nand U2019 (N_2019,In_139,In_729);
or U2020 (N_2020,In_748,In_216);
nand U2021 (N_2021,In_781,In_191);
nand U2022 (N_2022,In_705,In_763);
and U2023 (N_2023,In_934,In_128);
nand U2024 (N_2024,In_154,In_353);
and U2025 (N_2025,In_779,In_928);
or U2026 (N_2026,In_518,In_670);
nor U2027 (N_2027,In_266,In_91);
nor U2028 (N_2028,In_99,In_152);
or U2029 (N_2029,In_215,In_286);
or U2030 (N_2030,In_990,In_715);
and U2031 (N_2031,In_362,In_129);
nand U2032 (N_2032,In_975,In_484);
or U2033 (N_2033,In_307,In_613);
nor U2034 (N_2034,In_523,In_401);
and U2035 (N_2035,In_664,In_761);
or U2036 (N_2036,In_900,In_701);
nor U2037 (N_2037,In_102,In_637);
and U2038 (N_2038,In_639,In_606);
nor U2039 (N_2039,In_182,In_272);
nand U2040 (N_2040,In_905,In_20);
nand U2041 (N_2041,In_710,In_769);
nor U2042 (N_2042,In_556,In_524);
or U2043 (N_2043,In_82,In_604);
or U2044 (N_2044,In_350,In_785);
nor U2045 (N_2045,In_720,In_841);
or U2046 (N_2046,In_207,In_402);
or U2047 (N_2047,In_436,In_585);
nor U2048 (N_2048,In_46,In_311);
nand U2049 (N_2049,In_998,In_790);
and U2050 (N_2050,In_397,In_451);
and U2051 (N_2051,In_345,In_685);
nand U2052 (N_2052,In_147,In_591);
nand U2053 (N_2053,In_775,In_838);
nand U2054 (N_2054,In_482,In_656);
nand U2055 (N_2055,In_145,In_917);
nand U2056 (N_2056,In_404,In_259);
and U2057 (N_2057,In_114,In_412);
nand U2058 (N_2058,In_477,In_508);
and U2059 (N_2059,In_489,In_239);
and U2060 (N_2060,In_172,In_38);
and U2061 (N_2061,In_46,In_919);
nor U2062 (N_2062,In_783,In_211);
nand U2063 (N_2063,In_271,In_649);
or U2064 (N_2064,In_981,In_796);
and U2065 (N_2065,In_339,In_492);
or U2066 (N_2066,In_195,In_554);
or U2067 (N_2067,In_211,In_697);
nor U2068 (N_2068,In_215,In_218);
or U2069 (N_2069,In_601,In_725);
nand U2070 (N_2070,In_718,In_729);
and U2071 (N_2071,In_890,In_509);
nand U2072 (N_2072,In_426,In_894);
and U2073 (N_2073,In_271,In_525);
nor U2074 (N_2074,In_225,In_959);
nor U2075 (N_2075,In_950,In_398);
and U2076 (N_2076,In_626,In_604);
or U2077 (N_2077,In_339,In_245);
or U2078 (N_2078,In_737,In_948);
xnor U2079 (N_2079,In_286,In_811);
nand U2080 (N_2080,In_714,In_954);
and U2081 (N_2081,In_684,In_754);
or U2082 (N_2082,In_10,In_161);
and U2083 (N_2083,In_43,In_454);
nand U2084 (N_2084,In_251,In_226);
nand U2085 (N_2085,In_222,In_670);
or U2086 (N_2086,In_630,In_900);
nor U2087 (N_2087,In_924,In_972);
and U2088 (N_2088,In_305,In_383);
nand U2089 (N_2089,In_910,In_573);
nor U2090 (N_2090,In_991,In_54);
or U2091 (N_2091,In_791,In_786);
nand U2092 (N_2092,In_303,In_249);
or U2093 (N_2093,In_216,In_349);
nor U2094 (N_2094,In_653,In_433);
nor U2095 (N_2095,In_557,In_636);
nand U2096 (N_2096,In_378,In_913);
nand U2097 (N_2097,In_117,In_389);
and U2098 (N_2098,In_374,In_44);
and U2099 (N_2099,In_767,In_178);
nand U2100 (N_2100,In_375,In_25);
and U2101 (N_2101,In_693,In_296);
nand U2102 (N_2102,In_779,In_878);
or U2103 (N_2103,In_471,In_882);
nand U2104 (N_2104,In_466,In_432);
nor U2105 (N_2105,In_576,In_709);
nand U2106 (N_2106,In_990,In_166);
or U2107 (N_2107,In_273,In_580);
and U2108 (N_2108,In_99,In_667);
or U2109 (N_2109,In_688,In_967);
nor U2110 (N_2110,In_615,In_229);
or U2111 (N_2111,In_184,In_695);
and U2112 (N_2112,In_673,In_774);
or U2113 (N_2113,In_944,In_64);
nor U2114 (N_2114,In_997,In_400);
or U2115 (N_2115,In_438,In_512);
and U2116 (N_2116,In_559,In_361);
nor U2117 (N_2117,In_473,In_273);
and U2118 (N_2118,In_301,In_579);
or U2119 (N_2119,In_517,In_946);
or U2120 (N_2120,In_236,In_425);
and U2121 (N_2121,In_254,In_38);
and U2122 (N_2122,In_551,In_304);
nand U2123 (N_2123,In_1,In_261);
nand U2124 (N_2124,In_790,In_641);
nand U2125 (N_2125,In_721,In_810);
and U2126 (N_2126,In_829,In_721);
and U2127 (N_2127,In_961,In_822);
or U2128 (N_2128,In_771,In_494);
or U2129 (N_2129,In_256,In_998);
or U2130 (N_2130,In_225,In_452);
nor U2131 (N_2131,In_715,In_386);
nor U2132 (N_2132,In_545,In_130);
or U2133 (N_2133,In_560,In_102);
or U2134 (N_2134,In_92,In_878);
and U2135 (N_2135,In_563,In_170);
or U2136 (N_2136,In_383,In_980);
nor U2137 (N_2137,In_534,In_743);
nor U2138 (N_2138,In_109,In_765);
and U2139 (N_2139,In_577,In_364);
and U2140 (N_2140,In_601,In_425);
and U2141 (N_2141,In_306,In_174);
or U2142 (N_2142,In_414,In_634);
nor U2143 (N_2143,In_970,In_488);
and U2144 (N_2144,In_815,In_99);
nor U2145 (N_2145,In_187,In_99);
nand U2146 (N_2146,In_319,In_585);
or U2147 (N_2147,In_16,In_843);
nand U2148 (N_2148,In_576,In_961);
or U2149 (N_2149,In_536,In_67);
nand U2150 (N_2150,In_861,In_338);
and U2151 (N_2151,In_294,In_510);
nand U2152 (N_2152,In_601,In_924);
nor U2153 (N_2153,In_933,In_833);
or U2154 (N_2154,In_722,In_480);
nand U2155 (N_2155,In_89,In_728);
nand U2156 (N_2156,In_771,In_439);
nand U2157 (N_2157,In_351,In_648);
nor U2158 (N_2158,In_313,In_282);
or U2159 (N_2159,In_945,In_890);
or U2160 (N_2160,In_690,In_948);
nand U2161 (N_2161,In_103,In_560);
and U2162 (N_2162,In_741,In_227);
nand U2163 (N_2163,In_253,In_221);
nor U2164 (N_2164,In_621,In_536);
nand U2165 (N_2165,In_803,In_415);
nor U2166 (N_2166,In_525,In_494);
nand U2167 (N_2167,In_409,In_644);
or U2168 (N_2168,In_655,In_800);
or U2169 (N_2169,In_55,In_795);
or U2170 (N_2170,In_300,In_775);
nor U2171 (N_2171,In_99,In_496);
nor U2172 (N_2172,In_112,In_93);
xnor U2173 (N_2173,In_793,In_572);
and U2174 (N_2174,In_5,In_742);
and U2175 (N_2175,In_962,In_715);
and U2176 (N_2176,In_350,In_159);
or U2177 (N_2177,In_640,In_265);
and U2178 (N_2178,In_285,In_305);
nor U2179 (N_2179,In_799,In_774);
nor U2180 (N_2180,In_502,In_945);
and U2181 (N_2181,In_837,In_908);
or U2182 (N_2182,In_998,In_15);
or U2183 (N_2183,In_353,In_397);
nand U2184 (N_2184,In_49,In_143);
and U2185 (N_2185,In_976,In_199);
nor U2186 (N_2186,In_805,In_84);
or U2187 (N_2187,In_929,In_617);
nand U2188 (N_2188,In_889,In_543);
or U2189 (N_2189,In_631,In_95);
and U2190 (N_2190,In_601,In_548);
or U2191 (N_2191,In_829,In_697);
nand U2192 (N_2192,In_416,In_422);
and U2193 (N_2193,In_239,In_798);
nand U2194 (N_2194,In_134,In_825);
and U2195 (N_2195,In_950,In_446);
nand U2196 (N_2196,In_935,In_105);
nor U2197 (N_2197,In_23,In_715);
nor U2198 (N_2198,In_543,In_13);
and U2199 (N_2199,In_69,In_975);
xnor U2200 (N_2200,In_437,In_228);
or U2201 (N_2201,In_472,In_693);
or U2202 (N_2202,In_230,In_668);
nand U2203 (N_2203,In_730,In_644);
nor U2204 (N_2204,In_888,In_567);
nand U2205 (N_2205,In_303,In_302);
and U2206 (N_2206,In_232,In_403);
and U2207 (N_2207,In_11,In_106);
and U2208 (N_2208,In_554,In_241);
nor U2209 (N_2209,In_704,In_596);
nor U2210 (N_2210,In_634,In_992);
or U2211 (N_2211,In_410,In_326);
or U2212 (N_2212,In_95,In_61);
nor U2213 (N_2213,In_685,In_492);
or U2214 (N_2214,In_400,In_999);
and U2215 (N_2215,In_792,In_56);
or U2216 (N_2216,In_472,In_708);
or U2217 (N_2217,In_896,In_685);
nand U2218 (N_2218,In_232,In_531);
nor U2219 (N_2219,In_127,In_406);
nand U2220 (N_2220,In_756,In_930);
nor U2221 (N_2221,In_478,In_600);
and U2222 (N_2222,In_834,In_584);
nor U2223 (N_2223,In_494,In_920);
nand U2224 (N_2224,In_162,In_96);
or U2225 (N_2225,In_109,In_441);
nand U2226 (N_2226,In_212,In_362);
and U2227 (N_2227,In_149,In_186);
nand U2228 (N_2228,In_864,In_692);
or U2229 (N_2229,In_345,In_630);
or U2230 (N_2230,In_340,In_815);
nor U2231 (N_2231,In_639,In_856);
or U2232 (N_2232,In_858,In_31);
and U2233 (N_2233,In_966,In_496);
and U2234 (N_2234,In_576,In_981);
or U2235 (N_2235,In_338,In_1);
or U2236 (N_2236,In_547,In_370);
and U2237 (N_2237,In_811,In_430);
nand U2238 (N_2238,In_53,In_826);
nand U2239 (N_2239,In_916,In_223);
and U2240 (N_2240,In_888,In_580);
or U2241 (N_2241,In_749,In_628);
nand U2242 (N_2242,In_373,In_938);
nor U2243 (N_2243,In_128,In_792);
and U2244 (N_2244,In_470,In_927);
nand U2245 (N_2245,In_213,In_251);
nor U2246 (N_2246,In_9,In_938);
and U2247 (N_2247,In_587,In_864);
and U2248 (N_2248,In_278,In_912);
and U2249 (N_2249,In_2,In_597);
nand U2250 (N_2250,In_124,In_496);
nor U2251 (N_2251,In_31,In_188);
nor U2252 (N_2252,In_400,In_407);
or U2253 (N_2253,In_362,In_763);
or U2254 (N_2254,In_774,In_718);
nand U2255 (N_2255,In_731,In_19);
nor U2256 (N_2256,In_640,In_378);
nor U2257 (N_2257,In_759,In_478);
or U2258 (N_2258,In_954,In_965);
or U2259 (N_2259,In_432,In_892);
nand U2260 (N_2260,In_771,In_80);
and U2261 (N_2261,In_106,In_214);
or U2262 (N_2262,In_438,In_415);
nor U2263 (N_2263,In_852,In_516);
nor U2264 (N_2264,In_138,In_190);
and U2265 (N_2265,In_112,In_464);
and U2266 (N_2266,In_855,In_588);
and U2267 (N_2267,In_79,In_776);
or U2268 (N_2268,In_481,In_275);
or U2269 (N_2269,In_1,In_803);
nor U2270 (N_2270,In_513,In_237);
nand U2271 (N_2271,In_784,In_415);
or U2272 (N_2272,In_582,In_725);
and U2273 (N_2273,In_744,In_146);
nand U2274 (N_2274,In_270,In_812);
xnor U2275 (N_2275,In_197,In_919);
nor U2276 (N_2276,In_667,In_498);
and U2277 (N_2277,In_174,In_147);
nor U2278 (N_2278,In_819,In_718);
and U2279 (N_2279,In_211,In_843);
or U2280 (N_2280,In_724,In_200);
and U2281 (N_2281,In_162,In_338);
nor U2282 (N_2282,In_437,In_456);
and U2283 (N_2283,In_924,In_819);
nor U2284 (N_2284,In_40,In_263);
and U2285 (N_2285,In_297,In_667);
nor U2286 (N_2286,In_846,In_170);
and U2287 (N_2287,In_91,In_581);
and U2288 (N_2288,In_7,In_440);
nand U2289 (N_2289,In_764,In_485);
and U2290 (N_2290,In_514,In_868);
nor U2291 (N_2291,In_613,In_870);
nand U2292 (N_2292,In_670,In_332);
or U2293 (N_2293,In_856,In_214);
nand U2294 (N_2294,In_842,In_841);
and U2295 (N_2295,In_231,In_961);
and U2296 (N_2296,In_538,In_938);
nand U2297 (N_2297,In_223,In_114);
nand U2298 (N_2298,In_796,In_637);
nand U2299 (N_2299,In_716,In_27);
nand U2300 (N_2300,In_681,In_840);
nor U2301 (N_2301,In_933,In_320);
and U2302 (N_2302,In_228,In_708);
nor U2303 (N_2303,In_467,In_600);
or U2304 (N_2304,In_293,In_328);
nor U2305 (N_2305,In_114,In_697);
nor U2306 (N_2306,In_183,In_157);
or U2307 (N_2307,In_888,In_550);
and U2308 (N_2308,In_918,In_157);
and U2309 (N_2309,In_395,In_413);
or U2310 (N_2310,In_855,In_743);
and U2311 (N_2311,In_336,In_135);
nor U2312 (N_2312,In_300,In_247);
or U2313 (N_2313,In_748,In_161);
or U2314 (N_2314,In_949,In_362);
nand U2315 (N_2315,In_739,In_736);
or U2316 (N_2316,In_385,In_834);
nor U2317 (N_2317,In_641,In_171);
and U2318 (N_2318,In_698,In_799);
and U2319 (N_2319,In_906,In_180);
nand U2320 (N_2320,In_335,In_130);
or U2321 (N_2321,In_337,In_850);
or U2322 (N_2322,In_523,In_364);
nand U2323 (N_2323,In_122,In_467);
nor U2324 (N_2324,In_397,In_384);
nand U2325 (N_2325,In_427,In_411);
nand U2326 (N_2326,In_121,In_331);
or U2327 (N_2327,In_559,In_922);
and U2328 (N_2328,In_339,In_273);
and U2329 (N_2329,In_375,In_347);
nand U2330 (N_2330,In_685,In_213);
or U2331 (N_2331,In_752,In_126);
nor U2332 (N_2332,In_651,In_697);
and U2333 (N_2333,In_973,In_401);
nor U2334 (N_2334,In_940,In_664);
and U2335 (N_2335,In_543,In_770);
nor U2336 (N_2336,In_593,In_196);
nand U2337 (N_2337,In_670,In_622);
nor U2338 (N_2338,In_638,In_316);
or U2339 (N_2339,In_200,In_436);
and U2340 (N_2340,In_291,In_394);
nor U2341 (N_2341,In_735,In_745);
or U2342 (N_2342,In_884,In_551);
and U2343 (N_2343,In_959,In_517);
nor U2344 (N_2344,In_752,In_858);
nor U2345 (N_2345,In_821,In_221);
nand U2346 (N_2346,In_973,In_273);
nor U2347 (N_2347,In_332,In_405);
nand U2348 (N_2348,In_603,In_562);
and U2349 (N_2349,In_930,In_0);
and U2350 (N_2350,In_295,In_943);
nor U2351 (N_2351,In_676,In_208);
and U2352 (N_2352,In_704,In_283);
nor U2353 (N_2353,In_648,In_672);
and U2354 (N_2354,In_453,In_820);
nand U2355 (N_2355,In_331,In_363);
nor U2356 (N_2356,In_473,In_378);
nor U2357 (N_2357,In_787,In_517);
or U2358 (N_2358,In_863,In_524);
nor U2359 (N_2359,In_670,In_652);
nand U2360 (N_2360,In_855,In_238);
nor U2361 (N_2361,In_472,In_989);
and U2362 (N_2362,In_30,In_901);
nand U2363 (N_2363,In_94,In_81);
or U2364 (N_2364,In_195,In_603);
or U2365 (N_2365,In_550,In_708);
nor U2366 (N_2366,In_80,In_483);
nor U2367 (N_2367,In_906,In_557);
nor U2368 (N_2368,In_725,In_390);
nor U2369 (N_2369,In_443,In_577);
and U2370 (N_2370,In_438,In_917);
and U2371 (N_2371,In_3,In_530);
or U2372 (N_2372,In_329,In_161);
nand U2373 (N_2373,In_255,In_282);
nor U2374 (N_2374,In_110,In_708);
nor U2375 (N_2375,In_640,In_483);
nor U2376 (N_2376,In_915,In_883);
nor U2377 (N_2377,In_989,In_800);
and U2378 (N_2378,In_906,In_292);
nor U2379 (N_2379,In_229,In_658);
or U2380 (N_2380,In_484,In_76);
nand U2381 (N_2381,In_138,In_861);
nand U2382 (N_2382,In_718,In_940);
nor U2383 (N_2383,In_171,In_570);
nand U2384 (N_2384,In_216,In_303);
nor U2385 (N_2385,In_427,In_629);
or U2386 (N_2386,In_313,In_352);
and U2387 (N_2387,In_223,In_362);
nand U2388 (N_2388,In_807,In_340);
nand U2389 (N_2389,In_950,In_980);
nor U2390 (N_2390,In_452,In_472);
or U2391 (N_2391,In_611,In_848);
or U2392 (N_2392,In_63,In_768);
and U2393 (N_2393,In_149,In_718);
nand U2394 (N_2394,In_597,In_438);
or U2395 (N_2395,In_668,In_108);
nor U2396 (N_2396,In_404,In_670);
nor U2397 (N_2397,In_505,In_835);
nor U2398 (N_2398,In_957,In_206);
nor U2399 (N_2399,In_167,In_791);
nor U2400 (N_2400,In_12,In_136);
and U2401 (N_2401,In_679,In_745);
nor U2402 (N_2402,In_48,In_242);
nand U2403 (N_2403,In_878,In_349);
and U2404 (N_2404,In_75,In_902);
and U2405 (N_2405,In_682,In_351);
nand U2406 (N_2406,In_759,In_49);
and U2407 (N_2407,In_239,In_785);
nor U2408 (N_2408,In_633,In_967);
or U2409 (N_2409,In_60,In_594);
nor U2410 (N_2410,In_833,In_80);
nor U2411 (N_2411,In_610,In_709);
nand U2412 (N_2412,In_34,In_640);
and U2413 (N_2413,In_596,In_143);
nor U2414 (N_2414,In_67,In_618);
nand U2415 (N_2415,In_21,In_722);
and U2416 (N_2416,In_413,In_132);
and U2417 (N_2417,In_400,In_138);
and U2418 (N_2418,In_757,In_640);
or U2419 (N_2419,In_291,In_837);
nand U2420 (N_2420,In_750,In_144);
nand U2421 (N_2421,In_808,In_604);
nor U2422 (N_2422,In_348,In_239);
nand U2423 (N_2423,In_283,In_50);
or U2424 (N_2424,In_411,In_841);
and U2425 (N_2425,In_602,In_389);
nand U2426 (N_2426,In_458,In_627);
or U2427 (N_2427,In_247,In_470);
or U2428 (N_2428,In_982,In_652);
nor U2429 (N_2429,In_503,In_946);
and U2430 (N_2430,In_46,In_387);
nand U2431 (N_2431,In_128,In_754);
or U2432 (N_2432,In_974,In_648);
or U2433 (N_2433,In_463,In_438);
or U2434 (N_2434,In_443,In_744);
or U2435 (N_2435,In_653,In_534);
nand U2436 (N_2436,In_34,In_318);
and U2437 (N_2437,In_688,In_659);
or U2438 (N_2438,In_966,In_200);
nor U2439 (N_2439,In_899,In_238);
and U2440 (N_2440,In_373,In_488);
and U2441 (N_2441,In_814,In_292);
and U2442 (N_2442,In_81,In_49);
nor U2443 (N_2443,In_934,In_944);
and U2444 (N_2444,In_455,In_214);
nor U2445 (N_2445,In_457,In_556);
nand U2446 (N_2446,In_632,In_590);
nor U2447 (N_2447,In_921,In_257);
or U2448 (N_2448,In_930,In_641);
or U2449 (N_2449,In_941,In_127);
and U2450 (N_2450,In_820,In_999);
nor U2451 (N_2451,In_174,In_21);
or U2452 (N_2452,In_418,In_524);
or U2453 (N_2453,In_54,In_645);
nor U2454 (N_2454,In_436,In_843);
and U2455 (N_2455,In_275,In_169);
or U2456 (N_2456,In_602,In_554);
or U2457 (N_2457,In_653,In_217);
nor U2458 (N_2458,In_407,In_301);
nand U2459 (N_2459,In_967,In_150);
nand U2460 (N_2460,In_936,In_6);
nor U2461 (N_2461,In_452,In_213);
nand U2462 (N_2462,In_419,In_413);
and U2463 (N_2463,In_341,In_661);
and U2464 (N_2464,In_175,In_492);
or U2465 (N_2465,In_322,In_501);
or U2466 (N_2466,In_858,In_280);
and U2467 (N_2467,In_313,In_536);
and U2468 (N_2468,In_939,In_61);
and U2469 (N_2469,In_68,In_961);
nor U2470 (N_2470,In_153,In_243);
or U2471 (N_2471,In_909,In_384);
or U2472 (N_2472,In_889,In_294);
nand U2473 (N_2473,In_666,In_646);
and U2474 (N_2474,In_866,In_434);
and U2475 (N_2475,In_673,In_822);
or U2476 (N_2476,In_98,In_549);
nor U2477 (N_2477,In_696,In_975);
nand U2478 (N_2478,In_825,In_359);
nand U2479 (N_2479,In_625,In_244);
nand U2480 (N_2480,In_50,In_620);
nor U2481 (N_2481,In_655,In_361);
nand U2482 (N_2482,In_623,In_816);
nand U2483 (N_2483,In_284,In_446);
or U2484 (N_2484,In_680,In_937);
and U2485 (N_2485,In_731,In_966);
nor U2486 (N_2486,In_497,In_854);
and U2487 (N_2487,In_851,In_588);
and U2488 (N_2488,In_400,In_388);
or U2489 (N_2489,In_579,In_82);
and U2490 (N_2490,In_817,In_860);
and U2491 (N_2491,In_220,In_82);
xor U2492 (N_2492,In_339,In_344);
or U2493 (N_2493,In_716,In_206);
or U2494 (N_2494,In_298,In_297);
or U2495 (N_2495,In_710,In_119);
nor U2496 (N_2496,In_296,In_459);
or U2497 (N_2497,In_212,In_115);
or U2498 (N_2498,In_643,In_892);
nor U2499 (N_2499,In_776,In_228);
nand U2500 (N_2500,In_615,In_421);
or U2501 (N_2501,In_184,In_872);
nor U2502 (N_2502,In_648,In_547);
nor U2503 (N_2503,In_561,In_181);
or U2504 (N_2504,In_52,In_338);
nor U2505 (N_2505,In_295,In_868);
nor U2506 (N_2506,In_215,In_389);
and U2507 (N_2507,In_494,In_235);
or U2508 (N_2508,In_420,In_288);
and U2509 (N_2509,In_884,In_65);
nand U2510 (N_2510,In_49,In_199);
and U2511 (N_2511,In_94,In_213);
or U2512 (N_2512,In_998,In_941);
or U2513 (N_2513,In_825,In_328);
nor U2514 (N_2514,In_279,In_461);
or U2515 (N_2515,In_419,In_549);
or U2516 (N_2516,In_320,In_668);
or U2517 (N_2517,In_380,In_503);
and U2518 (N_2518,In_367,In_602);
and U2519 (N_2519,In_167,In_490);
or U2520 (N_2520,In_81,In_749);
nor U2521 (N_2521,In_966,In_956);
nand U2522 (N_2522,In_295,In_704);
nand U2523 (N_2523,In_592,In_995);
and U2524 (N_2524,In_96,In_672);
or U2525 (N_2525,In_27,In_938);
nor U2526 (N_2526,In_7,In_120);
nand U2527 (N_2527,In_861,In_937);
or U2528 (N_2528,In_301,In_401);
nand U2529 (N_2529,In_897,In_297);
or U2530 (N_2530,In_178,In_720);
or U2531 (N_2531,In_648,In_628);
and U2532 (N_2532,In_675,In_824);
nor U2533 (N_2533,In_619,In_241);
or U2534 (N_2534,In_548,In_845);
xnor U2535 (N_2535,In_118,In_120);
nor U2536 (N_2536,In_433,In_716);
nor U2537 (N_2537,In_418,In_94);
nand U2538 (N_2538,In_252,In_447);
nor U2539 (N_2539,In_663,In_346);
and U2540 (N_2540,In_686,In_824);
nand U2541 (N_2541,In_218,In_591);
and U2542 (N_2542,In_34,In_424);
and U2543 (N_2543,In_382,In_714);
nand U2544 (N_2544,In_228,In_727);
nor U2545 (N_2545,In_849,In_670);
nor U2546 (N_2546,In_403,In_194);
and U2547 (N_2547,In_683,In_969);
nand U2548 (N_2548,In_956,In_834);
or U2549 (N_2549,In_66,In_515);
nor U2550 (N_2550,In_10,In_97);
and U2551 (N_2551,In_830,In_611);
nor U2552 (N_2552,In_437,In_653);
and U2553 (N_2553,In_242,In_90);
nand U2554 (N_2554,In_43,In_30);
and U2555 (N_2555,In_190,In_230);
nor U2556 (N_2556,In_468,In_939);
nand U2557 (N_2557,In_486,In_749);
or U2558 (N_2558,In_543,In_50);
nand U2559 (N_2559,In_275,In_29);
and U2560 (N_2560,In_1,In_136);
nor U2561 (N_2561,In_252,In_633);
and U2562 (N_2562,In_957,In_358);
or U2563 (N_2563,In_96,In_511);
nand U2564 (N_2564,In_139,In_738);
and U2565 (N_2565,In_641,In_657);
nor U2566 (N_2566,In_202,In_242);
or U2567 (N_2567,In_839,In_892);
and U2568 (N_2568,In_173,In_8);
nor U2569 (N_2569,In_263,In_11);
or U2570 (N_2570,In_241,In_807);
nor U2571 (N_2571,In_810,In_320);
or U2572 (N_2572,In_582,In_625);
and U2573 (N_2573,In_325,In_355);
nor U2574 (N_2574,In_766,In_744);
nor U2575 (N_2575,In_650,In_495);
or U2576 (N_2576,In_879,In_862);
nor U2577 (N_2577,In_491,In_57);
nand U2578 (N_2578,In_179,In_407);
nor U2579 (N_2579,In_137,In_21);
and U2580 (N_2580,In_559,In_5);
or U2581 (N_2581,In_323,In_414);
nand U2582 (N_2582,In_287,In_456);
or U2583 (N_2583,In_75,In_568);
and U2584 (N_2584,In_198,In_666);
nor U2585 (N_2585,In_44,In_35);
nor U2586 (N_2586,In_997,In_689);
and U2587 (N_2587,In_747,In_106);
nor U2588 (N_2588,In_662,In_677);
nor U2589 (N_2589,In_617,In_184);
nand U2590 (N_2590,In_261,In_974);
nor U2591 (N_2591,In_299,In_498);
or U2592 (N_2592,In_743,In_812);
or U2593 (N_2593,In_16,In_662);
nand U2594 (N_2594,In_145,In_550);
nand U2595 (N_2595,In_387,In_715);
or U2596 (N_2596,In_555,In_733);
nand U2597 (N_2597,In_347,In_497);
nand U2598 (N_2598,In_610,In_124);
and U2599 (N_2599,In_185,In_742);
nor U2600 (N_2600,In_525,In_228);
and U2601 (N_2601,In_121,In_346);
nand U2602 (N_2602,In_643,In_914);
nor U2603 (N_2603,In_487,In_762);
and U2604 (N_2604,In_96,In_880);
and U2605 (N_2605,In_95,In_395);
nor U2606 (N_2606,In_496,In_30);
and U2607 (N_2607,In_390,In_84);
and U2608 (N_2608,In_338,In_295);
and U2609 (N_2609,In_191,In_887);
or U2610 (N_2610,In_639,In_918);
nand U2611 (N_2611,In_468,In_335);
nand U2612 (N_2612,In_402,In_844);
nor U2613 (N_2613,In_836,In_430);
or U2614 (N_2614,In_912,In_354);
and U2615 (N_2615,In_71,In_173);
and U2616 (N_2616,In_17,In_584);
nor U2617 (N_2617,In_432,In_204);
or U2618 (N_2618,In_777,In_806);
and U2619 (N_2619,In_465,In_235);
nor U2620 (N_2620,In_691,In_516);
nand U2621 (N_2621,In_361,In_791);
and U2622 (N_2622,In_547,In_155);
nand U2623 (N_2623,In_667,In_431);
or U2624 (N_2624,In_253,In_934);
or U2625 (N_2625,In_918,In_230);
and U2626 (N_2626,In_563,In_236);
or U2627 (N_2627,In_96,In_93);
xnor U2628 (N_2628,In_883,In_841);
nand U2629 (N_2629,In_132,In_992);
nor U2630 (N_2630,In_414,In_450);
nand U2631 (N_2631,In_794,In_496);
nor U2632 (N_2632,In_679,In_201);
nand U2633 (N_2633,In_883,In_28);
and U2634 (N_2634,In_220,In_191);
nand U2635 (N_2635,In_973,In_853);
nor U2636 (N_2636,In_64,In_619);
nand U2637 (N_2637,In_267,In_313);
and U2638 (N_2638,In_641,In_846);
nor U2639 (N_2639,In_169,In_260);
or U2640 (N_2640,In_852,In_599);
xnor U2641 (N_2641,In_896,In_445);
nand U2642 (N_2642,In_658,In_786);
or U2643 (N_2643,In_238,In_927);
nand U2644 (N_2644,In_91,In_565);
nand U2645 (N_2645,In_380,In_781);
nor U2646 (N_2646,In_543,In_447);
nand U2647 (N_2647,In_791,In_49);
nor U2648 (N_2648,In_608,In_762);
or U2649 (N_2649,In_164,In_721);
and U2650 (N_2650,In_419,In_916);
nand U2651 (N_2651,In_858,In_99);
and U2652 (N_2652,In_23,In_500);
nor U2653 (N_2653,In_984,In_712);
and U2654 (N_2654,In_757,In_441);
and U2655 (N_2655,In_842,In_871);
nor U2656 (N_2656,In_39,In_304);
and U2657 (N_2657,In_240,In_524);
and U2658 (N_2658,In_320,In_48);
nand U2659 (N_2659,In_191,In_677);
and U2660 (N_2660,In_205,In_523);
nor U2661 (N_2661,In_945,In_986);
or U2662 (N_2662,In_509,In_196);
nor U2663 (N_2663,In_629,In_568);
or U2664 (N_2664,In_61,In_673);
and U2665 (N_2665,In_715,In_196);
nor U2666 (N_2666,In_600,In_44);
or U2667 (N_2667,In_59,In_38);
or U2668 (N_2668,In_718,In_192);
nand U2669 (N_2669,In_126,In_249);
or U2670 (N_2670,In_785,In_43);
xnor U2671 (N_2671,In_582,In_357);
or U2672 (N_2672,In_407,In_91);
or U2673 (N_2673,In_558,In_227);
nor U2674 (N_2674,In_84,In_664);
nand U2675 (N_2675,In_445,In_623);
nor U2676 (N_2676,In_50,In_834);
and U2677 (N_2677,In_926,In_416);
and U2678 (N_2678,In_657,In_491);
or U2679 (N_2679,In_22,In_43);
and U2680 (N_2680,In_956,In_1);
and U2681 (N_2681,In_889,In_850);
nor U2682 (N_2682,In_712,In_969);
and U2683 (N_2683,In_19,In_710);
nor U2684 (N_2684,In_452,In_12);
or U2685 (N_2685,In_229,In_43);
xor U2686 (N_2686,In_980,In_988);
nand U2687 (N_2687,In_272,In_847);
or U2688 (N_2688,In_307,In_587);
nor U2689 (N_2689,In_940,In_315);
nand U2690 (N_2690,In_442,In_659);
and U2691 (N_2691,In_55,In_336);
nand U2692 (N_2692,In_62,In_497);
and U2693 (N_2693,In_598,In_525);
nand U2694 (N_2694,In_347,In_189);
and U2695 (N_2695,In_979,In_387);
and U2696 (N_2696,In_988,In_825);
and U2697 (N_2697,In_729,In_776);
nor U2698 (N_2698,In_370,In_726);
nand U2699 (N_2699,In_229,In_805);
and U2700 (N_2700,In_757,In_553);
or U2701 (N_2701,In_235,In_873);
nor U2702 (N_2702,In_111,In_815);
and U2703 (N_2703,In_395,In_918);
or U2704 (N_2704,In_160,In_477);
and U2705 (N_2705,In_191,In_13);
and U2706 (N_2706,In_609,In_347);
and U2707 (N_2707,In_702,In_734);
nand U2708 (N_2708,In_780,In_460);
nand U2709 (N_2709,In_744,In_51);
nor U2710 (N_2710,In_704,In_698);
nor U2711 (N_2711,In_469,In_169);
or U2712 (N_2712,In_498,In_653);
nor U2713 (N_2713,In_487,In_748);
xnor U2714 (N_2714,In_256,In_615);
or U2715 (N_2715,In_318,In_194);
nand U2716 (N_2716,In_253,In_513);
or U2717 (N_2717,In_604,In_143);
and U2718 (N_2718,In_959,In_393);
nor U2719 (N_2719,In_297,In_370);
nor U2720 (N_2720,In_350,In_43);
nor U2721 (N_2721,In_778,In_49);
nor U2722 (N_2722,In_573,In_969);
or U2723 (N_2723,In_385,In_308);
or U2724 (N_2724,In_813,In_500);
and U2725 (N_2725,In_31,In_956);
nor U2726 (N_2726,In_719,In_106);
or U2727 (N_2727,In_816,In_651);
or U2728 (N_2728,In_623,In_874);
and U2729 (N_2729,In_791,In_778);
nand U2730 (N_2730,In_79,In_313);
or U2731 (N_2731,In_400,In_254);
nand U2732 (N_2732,In_197,In_776);
and U2733 (N_2733,In_228,In_690);
nand U2734 (N_2734,In_834,In_693);
or U2735 (N_2735,In_260,In_648);
nor U2736 (N_2736,In_364,In_262);
nor U2737 (N_2737,In_350,In_547);
and U2738 (N_2738,In_839,In_848);
or U2739 (N_2739,In_457,In_503);
nor U2740 (N_2740,In_652,In_388);
or U2741 (N_2741,In_972,In_67);
or U2742 (N_2742,In_227,In_162);
or U2743 (N_2743,In_436,In_586);
and U2744 (N_2744,In_380,In_49);
nand U2745 (N_2745,In_731,In_428);
nor U2746 (N_2746,In_329,In_395);
or U2747 (N_2747,In_846,In_280);
or U2748 (N_2748,In_697,In_613);
nand U2749 (N_2749,In_961,In_77);
or U2750 (N_2750,In_567,In_349);
and U2751 (N_2751,In_873,In_736);
nand U2752 (N_2752,In_24,In_546);
nor U2753 (N_2753,In_797,In_61);
nand U2754 (N_2754,In_861,In_37);
nor U2755 (N_2755,In_770,In_746);
or U2756 (N_2756,In_694,In_85);
nand U2757 (N_2757,In_437,In_357);
nand U2758 (N_2758,In_487,In_459);
nor U2759 (N_2759,In_868,In_860);
nand U2760 (N_2760,In_927,In_453);
nand U2761 (N_2761,In_303,In_390);
and U2762 (N_2762,In_311,In_866);
and U2763 (N_2763,In_798,In_198);
and U2764 (N_2764,In_10,In_669);
or U2765 (N_2765,In_277,In_216);
and U2766 (N_2766,In_203,In_266);
and U2767 (N_2767,In_44,In_644);
nor U2768 (N_2768,In_760,In_52);
and U2769 (N_2769,In_369,In_860);
or U2770 (N_2770,In_128,In_389);
or U2771 (N_2771,In_157,In_977);
and U2772 (N_2772,In_349,In_159);
and U2773 (N_2773,In_14,In_735);
nand U2774 (N_2774,In_904,In_538);
or U2775 (N_2775,In_583,In_981);
nand U2776 (N_2776,In_187,In_672);
or U2777 (N_2777,In_307,In_700);
nor U2778 (N_2778,In_646,In_458);
and U2779 (N_2779,In_467,In_912);
or U2780 (N_2780,In_774,In_256);
nand U2781 (N_2781,In_916,In_865);
nand U2782 (N_2782,In_734,In_550);
and U2783 (N_2783,In_923,In_869);
nand U2784 (N_2784,In_96,In_896);
or U2785 (N_2785,In_679,In_343);
and U2786 (N_2786,In_319,In_355);
nand U2787 (N_2787,In_315,In_378);
nor U2788 (N_2788,In_277,In_688);
nand U2789 (N_2789,In_188,In_980);
or U2790 (N_2790,In_467,In_715);
and U2791 (N_2791,In_130,In_199);
nand U2792 (N_2792,In_832,In_472);
or U2793 (N_2793,In_912,In_996);
and U2794 (N_2794,In_149,In_89);
or U2795 (N_2795,In_191,In_575);
and U2796 (N_2796,In_250,In_510);
nand U2797 (N_2797,In_493,In_746);
and U2798 (N_2798,In_306,In_99);
nand U2799 (N_2799,In_528,In_39);
and U2800 (N_2800,In_841,In_162);
and U2801 (N_2801,In_743,In_874);
or U2802 (N_2802,In_235,In_612);
nor U2803 (N_2803,In_286,In_505);
or U2804 (N_2804,In_881,In_648);
or U2805 (N_2805,In_408,In_304);
nand U2806 (N_2806,In_231,In_20);
nor U2807 (N_2807,In_723,In_566);
or U2808 (N_2808,In_717,In_31);
nor U2809 (N_2809,In_63,In_652);
or U2810 (N_2810,In_24,In_11);
nand U2811 (N_2811,In_569,In_101);
nand U2812 (N_2812,In_896,In_51);
and U2813 (N_2813,In_797,In_294);
and U2814 (N_2814,In_272,In_365);
nor U2815 (N_2815,In_374,In_927);
nor U2816 (N_2816,In_464,In_417);
nor U2817 (N_2817,In_649,In_726);
nand U2818 (N_2818,In_477,In_18);
nand U2819 (N_2819,In_696,In_689);
or U2820 (N_2820,In_864,In_206);
or U2821 (N_2821,In_841,In_987);
nand U2822 (N_2822,In_453,In_525);
nand U2823 (N_2823,In_996,In_261);
or U2824 (N_2824,In_917,In_544);
nor U2825 (N_2825,In_437,In_268);
nor U2826 (N_2826,In_427,In_636);
nor U2827 (N_2827,In_448,In_35);
nand U2828 (N_2828,In_280,In_90);
and U2829 (N_2829,In_608,In_226);
nor U2830 (N_2830,In_924,In_67);
nor U2831 (N_2831,In_338,In_184);
or U2832 (N_2832,In_397,In_808);
and U2833 (N_2833,In_849,In_873);
nand U2834 (N_2834,In_919,In_773);
or U2835 (N_2835,In_929,In_636);
or U2836 (N_2836,In_331,In_747);
nor U2837 (N_2837,In_654,In_91);
nand U2838 (N_2838,In_938,In_876);
and U2839 (N_2839,In_398,In_887);
xnor U2840 (N_2840,In_791,In_972);
and U2841 (N_2841,In_635,In_910);
or U2842 (N_2842,In_942,In_462);
nor U2843 (N_2843,In_277,In_809);
nand U2844 (N_2844,In_911,In_186);
and U2845 (N_2845,In_498,In_737);
nand U2846 (N_2846,In_411,In_627);
or U2847 (N_2847,In_705,In_528);
nand U2848 (N_2848,In_375,In_368);
nand U2849 (N_2849,In_459,In_433);
or U2850 (N_2850,In_669,In_227);
nor U2851 (N_2851,In_646,In_600);
or U2852 (N_2852,In_976,In_886);
nor U2853 (N_2853,In_522,In_251);
nor U2854 (N_2854,In_529,In_450);
nor U2855 (N_2855,In_628,In_987);
or U2856 (N_2856,In_134,In_677);
nand U2857 (N_2857,In_73,In_643);
xnor U2858 (N_2858,In_846,In_273);
and U2859 (N_2859,In_527,In_41);
nand U2860 (N_2860,In_361,In_259);
or U2861 (N_2861,In_24,In_900);
nor U2862 (N_2862,In_475,In_30);
or U2863 (N_2863,In_289,In_856);
nor U2864 (N_2864,In_442,In_526);
nor U2865 (N_2865,In_842,In_539);
or U2866 (N_2866,In_219,In_511);
nand U2867 (N_2867,In_47,In_329);
and U2868 (N_2868,In_147,In_668);
nand U2869 (N_2869,In_463,In_140);
and U2870 (N_2870,In_932,In_121);
nor U2871 (N_2871,In_846,In_755);
and U2872 (N_2872,In_237,In_176);
and U2873 (N_2873,In_93,In_236);
nand U2874 (N_2874,In_789,In_803);
nor U2875 (N_2875,In_219,In_32);
nand U2876 (N_2876,In_898,In_7);
nor U2877 (N_2877,In_479,In_190);
nor U2878 (N_2878,In_385,In_489);
nand U2879 (N_2879,In_97,In_421);
nor U2880 (N_2880,In_827,In_559);
nand U2881 (N_2881,In_993,In_586);
nand U2882 (N_2882,In_560,In_628);
nor U2883 (N_2883,In_812,In_608);
nor U2884 (N_2884,In_69,In_370);
nor U2885 (N_2885,In_956,In_28);
nand U2886 (N_2886,In_555,In_695);
or U2887 (N_2887,In_962,In_556);
nand U2888 (N_2888,In_702,In_863);
nor U2889 (N_2889,In_436,In_885);
or U2890 (N_2890,In_72,In_851);
nand U2891 (N_2891,In_61,In_149);
and U2892 (N_2892,In_645,In_344);
nor U2893 (N_2893,In_850,In_822);
nor U2894 (N_2894,In_123,In_60);
nor U2895 (N_2895,In_302,In_738);
or U2896 (N_2896,In_532,In_248);
and U2897 (N_2897,In_761,In_296);
nor U2898 (N_2898,In_696,In_114);
nand U2899 (N_2899,In_354,In_758);
nor U2900 (N_2900,In_299,In_137);
or U2901 (N_2901,In_761,In_403);
or U2902 (N_2902,In_794,In_213);
and U2903 (N_2903,In_330,In_177);
or U2904 (N_2904,In_63,In_829);
or U2905 (N_2905,In_221,In_348);
nor U2906 (N_2906,In_307,In_439);
nor U2907 (N_2907,In_630,In_356);
nor U2908 (N_2908,In_874,In_729);
nand U2909 (N_2909,In_228,In_17);
xor U2910 (N_2910,In_495,In_105);
and U2911 (N_2911,In_274,In_92);
nand U2912 (N_2912,In_602,In_705);
or U2913 (N_2913,In_92,In_270);
and U2914 (N_2914,In_39,In_864);
and U2915 (N_2915,In_873,In_826);
nand U2916 (N_2916,In_383,In_29);
nand U2917 (N_2917,In_320,In_751);
or U2918 (N_2918,In_832,In_83);
xnor U2919 (N_2919,In_859,In_11);
or U2920 (N_2920,In_537,In_499);
nor U2921 (N_2921,In_818,In_374);
nand U2922 (N_2922,In_612,In_597);
or U2923 (N_2923,In_358,In_282);
or U2924 (N_2924,In_725,In_866);
nor U2925 (N_2925,In_17,In_112);
and U2926 (N_2926,In_321,In_391);
nand U2927 (N_2927,In_371,In_34);
nand U2928 (N_2928,In_23,In_358);
nand U2929 (N_2929,In_762,In_867);
nor U2930 (N_2930,In_134,In_552);
nor U2931 (N_2931,In_35,In_990);
or U2932 (N_2932,In_450,In_2);
and U2933 (N_2933,In_806,In_998);
or U2934 (N_2934,In_914,In_900);
nand U2935 (N_2935,In_615,In_219);
and U2936 (N_2936,In_692,In_32);
nor U2937 (N_2937,In_185,In_780);
or U2938 (N_2938,In_315,In_488);
or U2939 (N_2939,In_715,In_977);
or U2940 (N_2940,In_240,In_796);
nor U2941 (N_2941,In_291,In_975);
nand U2942 (N_2942,In_730,In_919);
or U2943 (N_2943,In_229,In_965);
or U2944 (N_2944,In_737,In_899);
and U2945 (N_2945,In_190,In_439);
or U2946 (N_2946,In_763,In_549);
and U2947 (N_2947,In_778,In_507);
and U2948 (N_2948,In_481,In_662);
and U2949 (N_2949,In_121,In_431);
nor U2950 (N_2950,In_282,In_95);
or U2951 (N_2951,In_843,In_151);
nand U2952 (N_2952,In_721,In_961);
or U2953 (N_2953,In_151,In_376);
nand U2954 (N_2954,In_733,In_65);
or U2955 (N_2955,In_723,In_992);
and U2956 (N_2956,In_302,In_460);
or U2957 (N_2957,In_951,In_609);
or U2958 (N_2958,In_321,In_999);
or U2959 (N_2959,In_408,In_317);
nand U2960 (N_2960,In_906,In_860);
nand U2961 (N_2961,In_69,In_315);
nor U2962 (N_2962,In_431,In_342);
and U2963 (N_2963,In_422,In_569);
and U2964 (N_2964,In_887,In_554);
nor U2965 (N_2965,In_531,In_971);
or U2966 (N_2966,In_788,In_842);
or U2967 (N_2967,In_381,In_465);
or U2968 (N_2968,In_514,In_712);
and U2969 (N_2969,In_666,In_724);
or U2970 (N_2970,In_194,In_578);
nand U2971 (N_2971,In_891,In_404);
nand U2972 (N_2972,In_516,In_617);
nand U2973 (N_2973,In_781,In_796);
and U2974 (N_2974,In_181,In_260);
and U2975 (N_2975,In_136,In_675);
and U2976 (N_2976,In_754,In_678);
xnor U2977 (N_2977,In_723,In_557);
or U2978 (N_2978,In_461,In_93);
nor U2979 (N_2979,In_217,In_232);
nand U2980 (N_2980,In_624,In_486);
nor U2981 (N_2981,In_440,In_625);
and U2982 (N_2982,In_875,In_401);
nor U2983 (N_2983,In_487,In_654);
and U2984 (N_2984,In_401,In_440);
nand U2985 (N_2985,In_93,In_270);
and U2986 (N_2986,In_285,In_347);
or U2987 (N_2987,In_40,In_77);
nand U2988 (N_2988,In_286,In_511);
nand U2989 (N_2989,In_408,In_314);
and U2990 (N_2990,In_348,In_214);
and U2991 (N_2991,In_183,In_549);
nand U2992 (N_2992,In_847,In_715);
and U2993 (N_2993,In_936,In_655);
or U2994 (N_2994,In_866,In_57);
and U2995 (N_2995,In_423,In_900);
and U2996 (N_2996,In_242,In_266);
and U2997 (N_2997,In_66,In_326);
nor U2998 (N_2998,In_555,In_744);
or U2999 (N_2999,In_444,In_901);
nor U3000 (N_3000,In_551,In_135);
nor U3001 (N_3001,In_141,In_775);
or U3002 (N_3002,In_257,In_312);
and U3003 (N_3003,In_798,In_176);
and U3004 (N_3004,In_891,In_201);
nand U3005 (N_3005,In_582,In_829);
nand U3006 (N_3006,In_912,In_926);
and U3007 (N_3007,In_76,In_628);
or U3008 (N_3008,In_92,In_327);
nand U3009 (N_3009,In_166,In_7);
nand U3010 (N_3010,In_482,In_0);
nand U3011 (N_3011,In_962,In_523);
nor U3012 (N_3012,In_397,In_295);
and U3013 (N_3013,In_711,In_877);
nor U3014 (N_3014,In_963,In_456);
or U3015 (N_3015,In_415,In_452);
nand U3016 (N_3016,In_240,In_880);
nor U3017 (N_3017,In_696,In_102);
nor U3018 (N_3018,In_792,In_654);
nand U3019 (N_3019,In_722,In_620);
nand U3020 (N_3020,In_913,In_49);
nor U3021 (N_3021,In_825,In_279);
nand U3022 (N_3022,In_37,In_112);
and U3023 (N_3023,In_801,In_11);
nor U3024 (N_3024,In_668,In_422);
or U3025 (N_3025,In_420,In_758);
and U3026 (N_3026,In_11,In_409);
and U3027 (N_3027,In_432,In_131);
and U3028 (N_3028,In_545,In_206);
nor U3029 (N_3029,In_947,In_405);
and U3030 (N_3030,In_887,In_853);
nor U3031 (N_3031,In_158,In_557);
or U3032 (N_3032,In_56,In_580);
nor U3033 (N_3033,In_631,In_212);
and U3034 (N_3034,In_663,In_660);
and U3035 (N_3035,In_656,In_528);
nand U3036 (N_3036,In_498,In_976);
or U3037 (N_3037,In_883,In_458);
nor U3038 (N_3038,In_760,In_772);
nand U3039 (N_3039,In_965,In_973);
nor U3040 (N_3040,In_201,In_831);
and U3041 (N_3041,In_889,In_389);
xor U3042 (N_3042,In_793,In_409);
and U3043 (N_3043,In_80,In_989);
or U3044 (N_3044,In_451,In_982);
or U3045 (N_3045,In_178,In_891);
and U3046 (N_3046,In_128,In_385);
or U3047 (N_3047,In_722,In_274);
and U3048 (N_3048,In_442,In_370);
and U3049 (N_3049,In_809,In_858);
or U3050 (N_3050,In_986,In_805);
nor U3051 (N_3051,In_332,In_740);
nand U3052 (N_3052,In_677,In_920);
nand U3053 (N_3053,In_926,In_222);
nor U3054 (N_3054,In_844,In_687);
nor U3055 (N_3055,In_796,In_162);
and U3056 (N_3056,In_208,In_768);
nor U3057 (N_3057,In_411,In_888);
nand U3058 (N_3058,In_930,In_614);
or U3059 (N_3059,In_995,In_490);
nand U3060 (N_3060,In_955,In_228);
or U3061 (N_3061,In_198,In_702);
and U3062 (N_3062,In_757,In_604);
nand U3063 (N_3063,In_244,In_781);
or U3064 (N_3064,In_223,In_873);
nor U3065 (N_3065,In_700,In_79);
and U3066 (N_3066,In_45,In_769);
nand U3067 (N_3067,In_995,In_666);
nand U3068 (N_3068,In_690,In_124);
and U3069 (N_3069,In_943,In_95);
or U3070 (N_3070,In_632,In_975);
nor U3071 (N_3071,In_428,In_985);
nand U3072 (N_3072,In_595,In_657);
xnor U3073 (N_3073,In_333,In_182);
and U3074 (N_3074,In_935,In_519);
and U3075 (N_3075,In_466,In_709);
and U3076 (N_3076,In_854,In_167);
nand U3077 (N_3077,In_803,In_708);
xor U3078 (N_3078,In_497,In_27);
and U3079 (N_3079,In_25,In_82);
or U3080 (N_3080,In_686,In_295);
nor U3081 (N_3081,In_707,In_283);
or U3082 (N_3082,In_811,In_926);
nor U3083 (N_3083,In_956,In_698);
and U3084 (N_3084,In_106,In_319);
nor U3085 (N_3085,In_575,In_740);
nand U3086 (N_3086,In_107,In_619);
and U3087 (N_3087,In_705,In_833);
nor U3088 (N_3088,In_128,In_348);
nor U3089 (N_3089,In_482,In_301);
and U3090 (N_3090,In_963,In_66);
and U3091 (N_3091,In_824,In_589);
nor U3092 (N_3092,In_486,In_717);
nor U3093 (N_3093,In_48,In_728);
or U3094 (N_3094,In_150,In_149);
or U3095 (N_3095,In_82,In_411);
xor U3096 (N_3096,In_242,In_858);
nor U3097 (N_3097,In_867,In_848);
or U3098 (N_3098,In_83,In_255);
nand U3099 (N_3099,In_779,In_862);
nor U3100 (N_3100,In_455,In_530);
or U3101 (N_3101,In_342,In_309);
nand U3102 (N_3102,In_295,In_961);
or U3103 (N_3103,In_425,In_325);
and U3104 (N_3104,In_690,In_628);
nand U3105 (N_3105,In_920,In_502);
nor U3106 (N_3106,In_593,In_961);
and U3107 (N_3107,In_639,In_952);
nor U3108 (N_3108,In_262,In_304);
nor U3109 (N_3109,In_600,In_166);
or U3110 (N_3110,In_917,In_769);
or U3111 (N_3111,In_475,In_394);
nand U3112 (N_3112,In_565,In_563);
or U3113 (N_3113,In_578,In_67);
nand U3114 (N_3114,In_194,In_441);
and U3115 (N_3115,In_343,In_509);
or U3116 (N_3116,In_326,In_122);
or U3117 (N_3117,In_743,In_896);
nand U3118 (N_3118,In_231,In_311);
and U3119 (N_3119,In_248,In_835);
and U3120 (N_3120,In_71,In_688);
nor U3121 (N_3121,In_824,In_778);
or U3122 (N_3122,In_608,In_922);
nand U3123 (N_3123,In_658,In_748);
nor U3124 (N_3124,In_192,In_449);
nor U3125 (N_3125,In_913,In_812);
or U3126 (N_3126,In_646,In_927);
or U3127 (N_3127,In_695,In_794);
or U3128 (N_3128,In_216,In_148);
and U3129 (N_3129,In_569,In_579);
and U3130 (N_3130,In_306,In_221);
nor U3131 (N_3131,In_722,In_527);
nand U3132 (N_3132,In_810,In_204);
or U3133 (N_3133,In_784,In_761);
nor U3134 (N_3134,In_111,In_134);
and U3135 (N_3135,In_150,In_524);
nand U3136 (N_3136,In_760,In_683);
and U3137 (N_3137,In_741,In_897);
or U3138 (N_3138,In_523,In_302);
nor U3139 (N_3139,In_237,In_538);
nand U3140 (N_3140,In_263,In_633);
and U3141 (N_3141,In_466,In_25);
nand U3142 (N_3142,In_899,In_549);
nor U3143 (N_3143,In_224,In_678);
or U3144 (N_3144,In_182,In_772);
nand U3145 (N_3145,In_805,In_75);
nor U3146 (N_3146,In_140,In_277);
nor U3147 (N_3147,In_147,In_454);
and U3148 (N_3148,In_351,In_771);
nor U3149 (N_3149,In_118,In_80);
or U3150 (N_3150,In_354,In_141);
or U3151 (N_3151,In_352,In_238);
nand U3152 (N_3152,In_616,In_218);
or U3153 (N_3153,In_915,In_423);
or U3154 (N_3154,In_800,In_610);
nand U3155 (N_3155,In_217,In_780);
and U3156 (N_3156,In_552,In_320);
and U3157 (N_3157,In_805,In_208);
and U3158 (N_3158,In_692,In_59);
and U3159 (N_3159,In_864,In_648);
or U3160 (N_3160,In_690,In_345);
nand U3161 (N_3161,In_314,In_317);
and U3162 (N_3162,In_752,In_122);
or U3163 (N_3163,In_161,In_806);
nand U3164 (N_3164,In_720,In_447);
and U3165 (N_3165,In_315,In_401);
and U3166 (N_3166,In_836,In_993);
or U3167 (N_3167,In_610,In_652);
and U3168 (N_3168,In_606,In_61);
or U3169 (N_3169,In_267,In_423);
or U3170 (N_3170,In_655,In_519);
or U3171 (N_3171,In_655,In_237);
and U3172 (N_3172,In_622,In_736);
nand U3173 (N_3173,In_330,In_897);
nor U3174 (N_3174,In_640,In_336);
nand U3175 (N_3175,In_713,In_396);
or U3176 (N_3176,In_560,In_865);
and U3177 (N_3177,In_970,In_737);
nand U3178 (N_3178,In_923,In_251);
nor U3179 (N_3179,In_499,In_6);
and U3180 (N_3180,In_482,In_163);
or U3181 (N_3181,In_263,In_112);
or U3182 (N_3182,In_712,In_524);
nor U3183 (N_3183,In_48,In_926);
or U3184 (N_3184,In_535,In_722);
and U3185 (N_3185,In_207,In_533);
nand U3186 (N_3186,In_247,In_917);
and U3187 (N_3187,In_926,In_273);
nor U3188 (N_3188,In_717,In_993);
nand U3189 (N_3189,In_504,In_660);
or U3190 (N_3190,In_307,In_311);
nor U3191 (N_3191,In_572,In_249);
nand U3192 (N_3192,In_656,In_371);
or U3193 (N_3193,In_285,In_103);
and U3194 (N_3194,In_701,In_150);
or U3195 (N_3195,In_589,In_322);
nor U3196 (N_3196,In_168,In_558);
nand U3197 (N_3197,In_866,In_387);
or U3198 (N_3198,In_414,In_251);
nand U3199 (N_3199,In_913,In_445);
and U3200 (N_3200,In_688,In_1);
and U3201 (N_3201,In_395,In_828);
or U3202 (N_3202,In_472,In_509);
nor U3203 (N_3203,In_371,In_417);
and U3204 (N_3204,In_656,In_36);
nor U3205 (N_3205,In_618,In_179);
nor U3206 (N_3206,In_312,In_21);
or U3207 (N_3207,In_48,In_809);
nor U3208 (N_3208,In_852,In_136);
nand U3209 (N_3209,In_62,In_491);
and U3210 (N_3210,In_882,In_867);
nor U3211 (N_3211,In_58,In_43);
xor U3212 (N_3212,In_104,In_817);
and U3213 (N_3213,In_633,In_970);
and U3214 (N_3214,In_497,In_784);
or U3215 (N_3215,In_881,In_869);
nor U3216 (N_3216,In_878,In_237);
or U3217 (N_3217,In_596,In_154);
and U3218 (N_3218,In_284,In_432);
nand U3219 (N_3219,In_356,In_522);
nor U3220 (N_3220,In_619,In_593);
nor U3221 (N_3221,In_299,In_6);
and U3222 (N_3222,In_560,In_713);
nor U3223 (N_3223,In_356,In_306);
or U3224 (N_3224,In_907,In_786);
or U3225 (N_3225,In_155,In_567);
and U3226 (N_3226,In_39,In_212);
nand U3227 (N_3227,In_314,In_55);
nand U3228 (N_3228,In_81,In_701);
and U3229 (N_3229,In_176,In_106);
nand U3230 (N_3230,In_887,In_936);
and U3231 (N_3231,In_721,In_572);
nand U3232 (N_3232,In_290,In_188);
nor U3233 (N_3233,In_289,In_829);
or U3234 (N_3234,In_515,In_897);
or U3235 (N_3235,In_309,In_109);
nand U3236 (N_3236,In_168,In_84);
nor U3237 (N_3237,In_819,In_363);
nor U3238 (N_3238,In_983,In_850);
nor U3239 (N_3239,In_525,In_888);
or U3240 (N_3240,In_568,In_414);
nor U3241 (N_3241,In_845,In_775);
nand U3242 (N_3242,In_19,In_450);
or U3243 (N_3243,In_116,In_186);
nand U3244 (N_3244,In_152,In_449);
and U3245 (N_3245,In_322,In_454);
or U3246 (N_3246,In_616,In_899);
and U3247 (N_3247,In_670,In_659);
nor U3248 (N_3248,In_785,In_190);
nand U3249 (N_3249,In_407,In_144);
nor U3250 (N_3250,In_880,In_332);
or U3251 (N_3251,In_223,In_586);
nand U3252 (N_3252,In_851,In_652);
and U3253 (N_3253,In_741,In_701);
nand U3254 (N_3254,In_447,In_353);
nor U3255 (N_3255,In_736,In_838);
nand U3256 (N_3256,In_647,In_447);
nor U3257 (N_3257,In_104,In_970);
and U3258 (N_3258,In_592,In_370);
and U3259 (N_3259,In_719,In_483);
and U3260 (N_3260,In_446,In_840);
nor U3261 (N_3261,In_650,In_98);
and U3262 (N_3262,In_433,In_153);
nand U3263 (N_3263,In_690,In_476);
nor U3264 (N_3264,In_790,In_521);
or U3265 (N_3265,In_210,In_894);
or U3266 (N_3266,In_986,In_176);
nor U3267 (N_3267,In_247,In_736);
and U3268 (N_3268,In_355,In_543);
or U3269 (N_3269,In_281,In_856);
and U3270 (N_3270,In_805,In_938);
nor U3271 (N_3271,In_489,In_844);
or U3272 (N_3272,In_133,In_256);
and U3273 (N_3273,In_893,In_120);
or U3274 (N_3274,In_571,In_573);
nor U3275 (N_3275,In_292,In_872);
nand U3276 (N_3276,In_645,In_566);
or U3277 (N_3277,In_523,In_912);
and U3278 (N_3278,In_312,In_968);
and U3279 (N_3279,In_562,In_518);
nand U3280 (N_3280,In_365,In_803);
nor U3281 (N_3281,In_105,In_162);
and U3282 (N_3282,In_495,In_892);
nand U3283 (N_3283,In_631,In_602);
and U3284 (N_3284,In_925,In_507);
and U3285 (N_3285,In_949,In_659);
nor U3286 (N_3286,In_654,In_409);
nand U3287 (N_3287,In_528,In_734);
or U3288 (N_3288,In_156,In_514);
and U3289 (N_3289,In_824,In_357);
nand U3290 (N_3290,In_312,In_747);
nor U3291 (N_3291,In_745,In_841);
or U3292 (N_3292,In_358,In_342);
and U3293 (N_3293,In_349,In_479);
nor U3294 (N_3294,In_285,In_676);
nor U3295 (N_3295,In_850,In_609);
or U3296 (N_3296,In_783,In_534);
nand U3297 (N_3297,In_442,In_462);
nor U3298 (N_3298,In_809,In_217);
nor U3299 (N_3299,In_916,In_156);
or U3300 (N_3300,In_40,In_401);
or U3301 (N_3301,In_69,In_636);
or U3302 (N_3302,In_458,In_893);
or U3303 (N_3303,In_752,In_607);
nand U3304 (N_3304,In_62,In_40);
nor U3305 (N_3305,In_739,In_113);
or U3306 (N_3306,In_360,In_619);
nor U3307 (N_3307,In_855,In_536);
nand U3308 (N_3308,In_523,In_712);
nand U3309 (N_3309,In_699,In_567);
nand U3310 (N_3310,In_656,In_562);
nand U3311 (N_3311,In_388,In_731);
nor U3312 (N_3312,In_89,In_991);
nor U3313 (N_3313,In_664,In_839);
or U3314 (N_3314,In_556,In_308);
nor U3315 (N_3315,In_957,In_378);
nand U3316 (N_3316,In_862,In_523);
and U3317 (N_3317,In_835,In_807);
nor U3318 (N_3318,In_645,In_820);
or U3319 (N_3319,In_380,In_450);
nand U3320 (N_3320,In_892,In_315);
or U3321 (N_3321,In_547,In_72);
or U3322 (N_3322,In_564,In_476);
and U3323 (N_3323,In_68,In_667);
and U3324 (N_3324,In_600,In_805);
nor U3325 (N_3325,In_171,In_386);
or U3326 (N_3326,In_144,In_203);
nand U3327 (N_3327,In_697,In_490);
and U3328 (N_3328,In_430,In_492);
and U3329 (N_3329,In_210,In_648);
or U3330 (N_3330,In_536,In_742);
or U3331 (N_3331,In_351,In_428);
and U3332 (N_3332,In_821,In_38);
and U3333 (N_3333,In_989,In_11);
and U3334 (N_3334,In_666,In_753);
or U3335 (N_3335,In_97,In_759);
and U3336 (N_3336,In_386,In_150);
or U3337 (N_3337,In_136,In_731);
nand U3338 (N_3338,In_595,In_847);
or U3339 (N_3339,In_973,In_872);
or U3340 (N_3340,In_3,In_824);
and U3341 (N_3341,In_526,In_487);
nor U3342 (N_3342,In_785,In_561);
nand U3343 (N_3343,In_210,In_861);
nor U3344 (N_3344,In_703,In_417);
or U3345 (N_3345,In_955,In_558);
or U3346 (N_3346,In_643,In_191);
nor U3347 (N_3347,In_726,In_997);
nor U3348 (N_3348,In_592,In_128);
nand U3349 (N_3349,In_892,In_76);
and U3350 (N_3350,In_345,In_913);
and U3351 (N_3351,In_805,In_12);
and U3352 (N_3352,In_565,In_757);
nand U3353 (N_3353,In_217,In_603);
and U3354 (N_3354,In_378,In_619);
or U3355 (N_3355,In_12,In_367);
nor U3356 (N_3356,In_411,In_201);
nor U3357 (N_3357,In_147,In_540);
nor U3358 (N_3358,In_361,In_147);
or U3359 (N_3359,In_721,In_129);
nor U3360 (N_3360,In_459,In_540);
nor U3361 (N_3361,In_180,In_181);
nand U3362 (N_3362,In_827,In_283);
nor U3363 (N_3363,In_298,In_8);
nand U3364 (N_3364,In_348,In_474);
nor U3365 (N_3365,In_54,In_142);
nand U3366 (N_3366,In_367,In_504);
nand U3367 (N_3367,In_504,In_653);
or U3368 (N_3368,In_482,In_17);
and U3369 (N_3369,In_674,In_949);
and U3370 (N_3370,In_57,In_585);
and U3371 (N_3371,In_706,In_100);
nor U3372 (N_3372,In_987,In_821);
nand U3373 (N_3373,In_416,In_742);
nor U3374 (N_3374,In_87,In_942);
or U3375 (N_3375,In_578,In_930);
or U3376 (N_3376,In_740,In_557);
and U3377 (N_3377,In_34,In_230);
nand U3378 (N_3378,In_421,In_198);
or U3379 (N_3379,In_868,In_402);
or U3380 (N_3380,In_730,In_970);
nor U3381 (N_3381,In_247,In_933);
and U3382 (N_3382,In_318,In_770);
nor U3383 (N_3383,In_498,In_58);
nand U3384 (N_3384,In_936,In_89);
and U3385 (N_3385,In_212,In_641);
and U3386 (N_3386,In_308,In_133);
or U3387 (N_3387,In_887,In_840);
and U3388 (N_3388,In_613,In_181);
nand U3389 (N_3389,In_924,In_6);
or U3390 (N_3390,In_813,In_283);
nor U3391 (N_3391,In_959,In_282);
nand U3392 (N_3392,In_336,In_833);
and U3393 (N_3393,In_567,In_29);
and U3394 (N_3394,In_953,In_346);
nand U3395 (N_3395,In_80,In_946);
nand U3396 (N_3396,In_641,In_365);
or U3397 (N_3397,In_735,In_871);
or U3398 (N_3398,In_765,In_30);
and U3399 (N_3399,In_722,In_765);
or U3400 (N_3400,In_188,In_356);
nor U3401 (N_3401,In_251,In_808);
nand U3402 (N_3402,In_987,In_126);
or U3403 (N_3403,In_197,In_604);
nand U3404 (N_3404,In_170,In_612);
nor U3405 (N_3405,In_664,In_5);
and U3406 (N_3406,In_601,In_935);
nor U3407 (N_3407,In_542,In_678);
nand U3408 (N_3408,In_305,In_330);
nor U3409 (N_3409,In_733,In_146);
and U3410 (N_3410,In_330,In_288);
nand U3411 (N_3411,In_322,In_39);
nor U3412 (N_3412,In_986,In_305);
nand U3413 (N_3413,In_550,In_656);
nor U3414 (N_3414,In_717,In_213);
or U3415 (N_3415,In_540,In_40);
nand U3416 (N_3416,In_233,In_392);
nor U3417 (N_3417,In_72,In_514);
nor U3418 (N_3418,In_270,In_172);
or U3419 (N_3419,In_327,In_866);
nor U3420 (N_3420,In_487,In_645);
and U3421 (N_3421,In_701,In_896);
and U3422 (N_3422,In_16,In_879);
or U3423 (N_3423,In_987,In_919);
or U3424 (N_3424,In_166,In_304);
nor U3425 (N_3425,In_36,In_580);
nand U3426 (N_3426,In_911,In_174);
and U3427 (N_3427,In_265,In_548);
or U3428 (N_3428,In_658,In_542);
nand U3429 (N_3429,In_860,In_111);
nor U3430 (N_3430,In_291,In_634);
and U3431 (N_3431,In_854,In_699);
or U3432 (N_3432,In_117,In_862);
and U3433 (N_3433,In_34,In_42);
nand U3434 (N_3434,In_514,In_154);
nor U3435 (N_3435,In_617,In_343);
nor U3436 (N_3436,In_620,In_601);
or U3437 (N_3437,In_414,In_361);
or U3438 (N_3438,In_814,In_244);
nand U3439 (N_3439,In_259,In_358);
nor U3440 (N_3440,In_933,In_670);
nand U3441 (N_3441,In_966,In_61);
nand U3442 (N_3442,In_815,In_463);
nand U3443 (N_3443,In_624,In_393);
nand U3444 (N_3444,In_632,In_772);
or U3445 (N_3445,In_721,In_703);
and U3446 (N_3446,In_846,In_682);
nor U3447 (N_3447,In_505,In_245);
xnor U3448 (N_3448,In_764,In_813);
or U3449 (N_3449,In_904,In_90);
nand U3450 (N_3450,In_484,In_269);
or U3451 (N_3451,In_606,In_523);
and U3452 (N_3452,In_187,In_129);
or U3453 (N_3453,In_107,In_941);
nor U3454 (N_3454,In_124,In_648);
nand U3455 (N_3455,In_219,In_444);
nand U3456 (N_3456,In_648,In_638);
nor U3457 (N_3457,In_808,In_285);
nand U3458 (N_3458,In_502,In_199);
nand U3459 (N_3459,In_80,In_122);
nor U3460 (N_3460,In_798,In_686);
xnor U3461 (N_3461,In_8,In_819);
nand U3462 (N_3462,In_481,In_413);
nand U3463 (N_3463,In_690,In_238);
nor U3464 (N_3464,In_326,In_295);
nor U3465 (N_3465,In_625,In_485);
nor U3466 (N_3466,In_916,In_22);
and U3467 (N_3467,In_249,In_283);
or U3468 (N_3468,In_785,In_906);
or U3469 (N_3469,In_464,In_375);
nand U3470 (N_3470,In_29,In_832);
and U3471 (N_3471,In_271,In_140);
nor U3472 (N_3472,In_117,In_711);
or U3473 (N_3473,In_667,In_688);
nor U3474 (N_3474,In_778,In_829);
and U3475 (N_3475,In_4,In_108);
or U3476 (N_3476,In_143,In_241);
nand U3477 (N_3477,In_437,In_526);
or U3478 (N_3478,In_257,In_671);
and U3479 (N_3479,In_810,In_702);
nand U3480 (N_3480,In_523,In_636);
nor U3481 (N_3481,In_367,In_97);
nand U3482 (N_3482,In_314,In_750);
and U3483 (N_3483,In_797,In_893);
nand U3484 (N_3484,In_71,In_92);
nor U3485 (N_3485,In_254,In_258);
nor U3486 (N_3486,In_534,In_432);
nor U3487 (N_3487,In_393,In_159);
or U3488 (N_3488,In_429,In_738);
and U3489 (N_3489,In_9,In_545);
and U3490 (N_3490,In_238,In_970);
nand U3491 (N_3491,In_781,In_930);
nand U3492 (N_3492,In_472,In_716);
and U3493 (N_3493,In_37,In_879);
nand U3494 (N_3494,In_445,In_948);
nand U3495 (N_3495,In_678,In_8);
or U3496 (N_3496,In_305,In_363);
nor U3497 (N_3497,In_469,In_538);
or U3498 (N_3498,In_252,In_440);
nand U3499 (N_3499,In_438,In_19);
nand U3500 (N_3500,In_634,In_279);
and U3501 (N_3501,In_987,In_373);
and U3502 (N_3502,In_247,In_623);
and U3503 (N_3503,In_60,In_876);
nor U3504 (N_3504,In_880,In_498);
nor U3505 (N_3505,In_253,In_784);
or U3506 (N_3506,In_427,In_5);
or U3507 (N_3507,In_746,In_376);
nand U3508 (N_3508,In_967,In_370);
or U3509 (N_3509,In_423,In_12);
nor U3510 (N_3510,In_632,In_364);
nor U3511 (N_3511,In_894,In_18);
nand U3512 (N_3512,In_401,In_932);
and U3513 (N_3513,In_141,In_228);
nand U3514 (N_3514,In_520,In_277);
and U3515 (N_3515,In_661,In_474);
nand U3516 (N_3516,In_382,In_308);
nand U3517 (N_3517,In_938,In_424);
nand U3518 (N_3518,In_148,In_582);
and U3519 (N_3519,In_788,In_416);
nor U3520 (N_3520,In_460,In_143);
and U3521 (N_3521,In_110,In_616);
and U3522 (N_3522,In_846,In_427);
xnor U3523 (N_3523,In_980,In_824);
or U3524 (N_3524,In_983,In_895);
nand U3525 (N_3525,In_600,In_620);
or U3526 (N_3526,In_390,In_386);
and U3527 (N_3527,In_0,In_73);
and U3528 (N_3528,In_840,In_730);
nor U3529 (N_3529,In_334,In_594);
or U3530 (N_3530,In_959,In_468);
and U3531 (N_3531,In_724,In_378);
and U3532 (N_3532,In_77,In_775);
nor U3533 (N_3533,In_743,In_300);
or U3534 (N_3534,In_916,In_561);
nand U3535 (N_3535,In_394,In_624);
nor U3536 (N_3536,In_451,In_551);
nand U3537 (N_3537,In_863,In_569);
nor U3538 (N_3538,In_454,In_142);
nand U3539 (N_3539,In_582,In_174);
nor U3540 (N_3540,In_754,In_62);
nor U3541 (N_3541,In_795,In_878);
and U3542 (N_3542,In_190,In_234);
nor U3543 (N_3543,In_485,In_904);
or U3544 (N_3544,In_146,In_110);
nor U3545 (N_3545,In_492,In_187);
or U3546 (N_3546,In_786,In_555);
and U3547 (N_3547,In_195,In_202);
or U3548 (N_3548,In_574,In_660);
or U3549 (N_3549,In_50,In_152);
nor U3550 (N_3550,In_414,In_855);
nor U3551 (N_3551,In_27,In_159);
and U3552 (N_3552,In_970,In_265);
nor U3553 (N_3553,In_925,In_299);
nand U3554 (N_3554,In_600,In_490);
nand U3555 (N_3555,In_53,In_727);
or U3556 (N_3556,In_35,In_521);
nand U3557 (N_3557,In_130,In_255);
nor U3558 (N_3558,In_598,In_503);
or U3559 (N_3559,In_593,In_977);
nor U3560 (N_3560,In_425,In_725);
nand U3561 (N_3561,In_715,In_0);
and U3562 (N_3562,In_93,In_822);
or U3563 (N_3563,In_754,In_173);
or U3564 (N_3564,In_488,In_941);
nand U3565 (N_3565,In_842,In_224);
and U3566 (N_3566,In_352,In_146);
or U3567 (N_3567,In_357,In_939);
and U3568 (N_3568,In_869,In_880);
nor U3569 (N_3569,In_355,In_861);
nor U3570 (N_3570,In_556,In_26);
nand U3571 (N_3571,In_95,In_253);
nor U3572 (N_3572,In_138,In_163);
nor U3573 (N_3573,In_972,In_319);
or U3574 (N_3574,In_79,In_193);
nand U3575 (N_3575,In_626,In_780);
and U3576 (N_3576,In_646,In_868);
and U3577 (N_3577,In_812,In_48);
nand U3578 (N_3578,In_29,In_137);
or U3579 (N_3579,In_43,In_376);
nand U3580 (N_3580,In_813,In_429);
nand U3581 (N_3581,In_422,In_413);
nand U3582 (N_3582,In_292,In_870);
nand U3583 (N_3583,In_893,In_868);
nor U3584 (N_3584,In_182,In_119);
nand U3585 (N_3585,In_858,In_731);
nor U3586 (N_3586,In_558,In_237);
nor U3587 (N_3587,In_237,In_276);
nand U3588 (N_3588,In_430,In_7);
nor U3589 (N_3589,In_778,In_688);
nand U3590 (N_3590,In_245,In_560);
nand U3591 (N_3591,In_129,In_196);
or U3592 (N_3592,In_489,In_122);
nand U3593 (N_3593,In_534,In_180);
and U3594 (N_3594,In_970,In_402);
nand U3595 (N_3595,In_99,In_776);
nand U3596 (N_3596,In_173,In_801);
nor U3597 (N_3597,In_176,In_307);
or U3598 (N_3598,In_732,In_912);
nand U3599 (N_3599,In_949,In_481);
or U3600 (N_3600,In_471,In_75);
or U3601 (N_3601,In_15,In_413);
and U3602 (N_3602,In_419,In_278);
and U3603 (N_3603,In_708,In_356);
or U3604 (N_3604,In_348,In_366);
nor U3605 (N_3605,In_618,In_754);
nor U3606 (N_3606,In_482,In_743);
nor U3607 (N_3607,In_675,In_569);
and U3608 (N_3608,In_952,In_245);
or U3609 (N_3609,In_211,In_153);
or U3610 (N_3610,In_621,In_360);
and U3611 (N_3611,In_669,In_986);
and U3612 (N_3612,In_423,In_101);
nor U3613 (N_3613,In_331,In_771);
nand U3614 (N_3614,In_197,In_800);
or U3615 (N_3615,In_505,In_238);
and U3616 (N_3616,In_717,In_433);
nand U3617 (N_3617,In_920,In_597);
and U3618 (N_3618,In_891,In_63);
or U3619 (N_3619,In_493,In_167);
nor U3620 (N_3620,In_329,In_332);
nand U3621 (N_3621,In_960,In_950);
nor U3622 (N_3622,In_974,In_862);
nor U3623 (N_3623,In_703,In_723);
nor U3624 (N_3624,In_481,In_24);
nand U3625 (N_3625,In_395,In_32);
nand U3626 (N_3626,In_478,In_514);
or U3627 (N_3627,In_588,In_668);
nor U3628 (N_3628,In_792,In_842);
and U3629 (N_3629,In_912,In_139);
and U3630 (N_3630,In_371,In_960);
nor U3631 (N_3631,In_328,In_708);
nor U3632 (N_3632,In_751,In_966);
or U3633 (N_3633,In_523,In_778);
nand U3634 (N_3634,In_274,In_730);
nor U3635 (N_3635,In_757,In_711);
nand U3636 (N_3636,In_360,In_831);
nand U3637 (N_3637,In_806,In_546);
nand U3638 (N_3638,In_791,In_950);
nor U3639 (N_3639,In_433,In_338);
and U3640 (N_3640,In_880,In_45);
nand U3641 (N_3641,In_380,In_829);
nor U3642 (N_3642,In_927,In_318);
nand U3643 (N_3643,In_743,In_498);
or U3644 (N_3644,In_119,In_269);
and U3645 (N_3645,In_94,In_245);
or U3646 (N_3646,In_159,In_318);
and U3647 (N_3647,In_366,In_326);
nand U3648 (N_3648,In_77,In_981);
nor U3649 (N_3649,In_271,In_236);
nand U3650 (N_3650,In_28,In_942);
nand U3651 (N_3651,In_364,In_723);
or U3652 (N_3652,In_471,In_696);
nand U3653 (N_3653,In_908,In_233);
nor U3654 (N_3654,In_461,In_759);
or U3655 (N_3655,In_966,In_182);
nor U3656 (N_3656,In_642,In_145);
or U3657 (N_3657,In_603,In_985);
or U3658 (N_3658,In_350,In_539);
or U3659 (N_3659,In_938,In_512);
nand U3660 (N_3660,In_147,In_534);
or U3661 (N_3661,In_155,In_16);
nand U3662 (N_3662,In_586,In_997);
and U3663 (N_3663,In_263,In_694);
nor U3664 (N_3664,In_313,In_330);
or U3665 (N_3665,In_692,In_955);
or U3666 (N_3666,In_85,In_380);
nor U3667 (N_3667,In_741,In_871);
nor U3668 (N_3668,In_282,In_859);
nor U3669 (N_3669,In_370,In_368);
or U3670 (N_3670,In_603,In_348);
nor U3671 (N_3671,In_990,In_165);
nor U3672 (N_3672,In_909,In_272);
xor U3673 (N_3673,In_858,In_386);
nand U3674 (N_3674,In_700,In_659);
xor U3675 (N_3675,In_213,In_659);
nand U3676 (N_3676,In_524,In_408);
nor U3677 (N_3677,In_969,In_779);
nand U3678 (N_3678,In_674,In_708);
nand U3679 (N_3679,In_878,In_964);
nand U3680 (N_3680,In_304,In_210);
nor U3681 (N_3681,In_149,In_442);
or U3682 (N_3682,In_508,In_136);
nand U3683 (N_3683,In_832,In_374);
and U3684 (N_3684,In_417,In_707);
nor U3685 (N_3685,In_775,In_360);
and U3686 (N_3686,In_474,In_846);
nand U3687 (N_3687,In_372,In_197);
nand U3688 (N_3688,In_511,In_793);
and U3689 (N_3689,In_352,In_376);
or U3690 (N_3690,In_461,In_838);
nand U3691 (N_3691,In_787,In_452);
nand U3692 (N_3692,In_966,In_127);
and U3693 (N_3693,In_415,In_966);
or U3694 (N_3694,In_250,In_163);
or U3695 (N_3695,In_662,In_43);
nand U3696 (N_3696,In_881,In_835);
or U3697 (N_3697,In_228,In_48);
xnor U3698 (N_3698,In_100,In_195);
nand U3699 (N_3699,In_257,In_383);
nor U3700 (N_3700,In_473,In_432);
and U3701 (N_3701,In_676,In_715);
nor U3702 (N_3702,In_677,In_91);
and U3703 (N_3703,In_180,In_722);
and U3704 (N_3704,In_531,In_862);
nand U3705 (N_3705,In_430,In_864);
or U3706 (N_3706,In_585,In_326);
nor U3707 (N_3707,In_169,In_450);
and U3708 (N_3708,In_707,In_755);
and U3709 (N_3709,In_5,In_487);
nand U3710 (N_3710,In_18,In_800);
xnor U3711 (N_3711,In_785,In_334);
and U3712 (N_3712,In_330,In_810);
or U3713 (N_3713,In_283,In_973);
or U3714 (N_3714,In_787,In_181);
or U3715 (N_3715,In_265,In_921);
and U3716 (N_3716,In_384,In_932);
nand U3717 (N_3717,In_517,In_86);
nand U3718 (N_3718,In_56,In_430);
xor U3719 (N_3719,In_884,In_714);
nor U3720 (N_3720,In_660,In_416);
and U3721 (N_3721,In_564,In_704);
or U3722 (N_3722,In_187,In_132);
or U3723 (N_3723,In_429,In_660);
nor U3724 (N_3724,In_342,In_940);
or U3725 (N_3725,In_921,In_107);
and U3726 (N_3726,In_582,In_75);
nor U3727 (N_3727,In_872,In_837);
nand U3728 (N_3728,In_75,In_836);
and U3729 (N_3729,In_499,In_198);
and U3730 (N_3730,In_131,In_795);
nand U3731 (N_3731,In_42,In_127);
or U3732 (N_3732,In_330,In_503);
nor U3733 (N_3733,In_405,In_397);
and U3734 (N_3734,In_785,In_683);
and U3735 (N_3735,In_737,In_574);
nand U3736 (N_3736,In_857,In_320);
and U3737 (N_3737,In_598,In_41);
and U3738 (N_3738,In_969,In_676);
or U3739 (N_3739,In_638,In_668);
nand U3740 (N_3740,In_76,In_69);
and U3741 (N_3741,In_54,In_630);
nand U3742 (N_3742,In_14,In_432);
nor U3743 (N_3743,In_947,In_809);
or U3744 (N_3744,In_115,In_135);
nand U3745 (N_3745,In_580,In_577);
and U3746 (N_3746,In_550,In_674);
and U3747 (N_3747,In_492,In_635);
and U3748 (N_3748,In_184,In_356);
or U3749 (N_3749,In_988,In_408);
or U3750 (N_3750,In_452,In_610);
or U3751 (N_3751,In_904,In_459);
nand U3752 (N_3752,In_185,In_720);
nor U3753 (N_3753,In_83,In_434);
nand U3754 (N_3754,In_776,In_862);
and U3755 (N_3755,In_266,In_667);
nand U3756 (N_3756,In_964,In_936);
and U3757 (N_3757,In_420,In_838);
or U3758 (N_3758,In_985,In_924);
or U3759 (N_3759,In_324,In_402);
and U3760 (N_3760,In_975,In_341);
nor U3761 (N_3761,In_28,In_914);
or U3762 (N_3762,In_636,In_780);
nand U3763 (N_3763,In_823,In_348);
nor U3764 (N_3764,In_858,In_369);
and U3765 (N_3765,In_90,In_309);
nor U3766 (N_3766,In_78,In_444);
and U3767 (N_3767,In_4,In_499);
nor U3768 (N_3768,In_709,In_166);
and U3769 (N_3769,In_39,In_149);
nand U3770 (N_3770,In_614,In_891);
nor U3771 (N_3771,In_630,In_106);
nand U3772 (N_3772,In_621,In_441);
or U3773 (N_3773,In_667,In_452);
and U3774 (N_3774,In_87,In_928);
or U3775 (N_3775,In_183,In_127);
or U3776 (N_3776,In_172,In_996);
nor U3777 (N_3777,In_116,In_249);
nor U3778 (N_3778,In_536,In_37);
or U3779 (N_3779,In_342,In_165);
nor U3780 (N_3780,In_354,In_279);
nor U3781 (N_3781,In_406,In_479);
nor U3782 (N_3782,In_216,In_761);
nand U3783 (N_3783,In_939,In_511);
nand U3784 (N_3784,In_760,In_710);
and U3785 (N_3785,In_980,In_234);
and U3786 (N_3786,In_438,In_644);
and U3787 (N_3787,In_997,In_989);
or U3788 (N_3788,In_944,In_622);
or U3789 (N_3789,In_444,In_863);
or U3790 (N_3790,In_35,In_69);
nand U3791 (N_3791,In_59,In_108);
and U3792 (N_3792,In_213,In_468);
nor U3793 (N_3793,In_800,In_567);
nand U3794 (N_3794,In_888,In_458);
and U3795 (N_3795,In_723,In_289);
nand U3796 (N_3796,In_356,In_813);
and U3797 (N_3797,In_476,In_285);
or U3798 (N_3798,In_866,In_82);
or U3799 (N_3799,In_563,In_160);
and U3800 (N_3800,In_941,In_891);
nor U3801 (N_3801,In_403,In_343);
and U3802 (N_3802,In_987,In_391);
nand U3803 (N_3803,In_485,In_769);
and U3804 (N_3804,In_873,In_375);
and U3805 (N_3805,In_429,In_377);
or U3806 (N_3806,In_472,In_782);
or U3807 (N_3807,In_460,In_366);
nor U3808 (N_3808,In_440,In_818);
nor U3809 (N_3809,In_998,In_812);
nand U3810 (N_3810,In_391,In_115);
or U3811 (N_3811,In_590,In_199);
nand U3812 (N_3812,In_256,In_161);
nand U3813 (N_3813,In_599,In_617);
nand U3814 (N_3814,In_293,In_644);
nor U3815 (N_3815,In_388,In_970);
nand U3816 (N_3816,In_992,In_521);
and U3817 (N_3817,In_989,In_936);
and U3818 (N_3818,In_329,In_159);
xor U3819 (N_3819,In_303,In_447);
and U3820 (N_3820,In_735,In_847);
or U3821 (N_3821,In_888,In_755);
or U3822 (N_3822,In_311,In_157);
xor U3823 (N_3823,In_727,In_263);
or U3824 (N_3824,In_77,In_466);
nand U3825 (N_3825,In_174,In_124);
nand U3826 (N_3826,In_687,In_905);
and U3827 (N_3827,In_81,In_108);
nand U3828 (N_3828,In_348,In_323);
and U3829 (N_3829,In_353,In_212);
and U3830 (N_3830,In_647,In_563);
nand U3831 (N_3831,In_49,In_72);
nand U3832 (N_3832,In_134,In_339);
or U3833 (N_3833,In_50,In_262);
and U3834 (N_3834,In_379,In_272);
or U3835 (N_3835,In_720,In_543);
nor U3836 (N_3836,In_12,In_847);
nand U3837 (N_3837,In_972,In_854);
xnor U3838 (N_3838,In_856,In_814);
or U3839 (N_3839,In_579,In_132);
nand U3840 (N_3840,In_142,In_176);
nor U3841 (N_3841,In_351,In_446);
and U3842 (N_3842,In_291,In_391);
or U3843 (N_3843,In_438,In_122);
nor U3844 (N_3844,In_332,In_180);
nand U3845 (N_3845,In_43,In_978);
and U3846 (N_3846,In_541,In_24);
nor U3847 (N_3847,In_257,In_941);
nand U3848 (N_3848,In_606,In_790);
nor U3849 (N_3849,In_734,In_655);
or U3850 (N_3850,In_514,In_341);
or U3851 (N_3851,In_645,In_615);
and U3852 (N_3852,In_289,In_561);
and U3853 (N_3853,In_149,In_239);
nor U3854 (N_3854,In_871,In_317);
nand U3855 (N_3855,In_279,In_228);
nor U3856 (N_3856,In_700,In_615);
nand U3857 (N_3857,In_450,In_88);
nor U3858 (N_3858,In_975,In_181);
nor U3859 (N_3859,In_80,In_184);
nand U3860 (N_3860,In_309,In_830);
or U3861 (N_3861,In_900,In_257);
or U3862 (N_3862,In_394,In_683);
nor U3863 (N_3863,In_891,In_763);
nand U3864 (N_3864,In_63,In_933);
or U3865 (N_3865,In_504,In_95);
nand U3866 (N_3866,In_317,In_481);
or U3867 (N_3867,In_111,In_682);
nor U3868 (N_3868,In_225,In_831);
or U3869 (N_3869,In_386,In_847);
nor U3870 (N_3870,In_217,In_564);
and U3871 (N_3871,In_887,In_92);
and U3872 (N_3872,In_355,In_914);
and U3873 (N_3873,In_362,In_597);
and U3874 (N_3874,In_719,In_440);
nand U3875 (N_3875,In_828,In_998);
nand U3876 (N_3876,In_655,In_458);
or U3877 (N_3877,In_883,In_760);
nor U3878 (N_3878,In_367,In_297);
and U3879 (N_3879,In_626,In_300);
nand U3880 (N_3880,In_989,In_649);
or U3881 (N_3881,In_661,In_221);
or U3882 (N_3882,In_242,In_825);
and U3883 (N_3883,In_674,In_945);
or U3884 (N_3884,In_308,In_964);
nand U3885 (N_3885,In_302,In_960);
or U3886 (N_3886,In_709,In_867);
or U3887 (N_3887,In_194,In_131);
and U3888 (N_3888,In_431,In_285);
and U3889 (N_3889,In_317,In_733);
and U3890 (N_3890,In_208,In_772);
or U3891 (N_3891,In_362,In_153);
nand U3892 (N_3892,In_861,In_408);
and U3893 (N_3893,In_580,In_790);
and U3894 (N_3894,In_816,In_250);
nor U3895 (N_3895,In_195,In_812);
nor U3896 (N_3896,In_857,In_817);
and U3897 (N_3897,In_160,In_555);
nor U3898 (N_3898,In_237,In_927);
and U3899 (N_3899,In_601,In_610);
nor U3900 (N_3900,In_419,In_559);
nand U3901 (N_3901,In_186,In_139);
nand U3902 (N_3902,In_717,In_852);
and U3903 (N_3903,In_552,In_936);
and U3904 (N_3904,In_715,In_148);
and U3905 (N_3905,In_22,In_133);
nand U3906 (N_3906,In_23,In_883);
nand U3907 (N_3907,In_501,In_780);
nand U3908 (N_3908,In_36,In_811);
nand U3909 (N_3909,In_226,In_707);
or U3910 (N_3910,In_821,In_191);
or U3911 (N_3911,In_73,In_620);
or U3912 (N_3912,In_6,In_145);
or U3913 (N_3913,In_763,In_342);
and U3914 (N_3914,In_621,In_708);
and U3915 (N_3915,In_452,In_32);
nand U3916 (N_3916,In_828,In_258);
nand U3917 (N_3917,In_336,In_511);
xor U3918 (N_3918,In_953,In_525);
or U3919 (N_3919,In_321,In_776);
nand U3920 (N_3920,In_644,In_359);
and U3921 (N_3921,In_241,In_25);
and U3922 (N_3922,In_541,In_744);
xnor U3923 (N_3923,In_880,In_141);
nand U3924 (N_3924,In_845,In_871);
or U3925 (N_3925,In_189,In_395);
and U3926 (N_3926,In_433,In_226);
and U3927 (N_3927,In_783,In_720);
or U3928 (N_3928,In_816,In_169);
nand U3929 (N_3929,In_882,In_583);
nor U3930 (N_3930,In_813,In_387);
and U3931 (N_3931,In_898,In_937);
nand U3932 (N_3932,In_535,In_448);
and U3933 (N_3933,In_79,In_782);
and U3934 (N_3934,In_132,In_352);
or U3935 (N_3935,In_605,In_185);
nand U3936 (N_3936,In_554,In_392);
or U3937 (N_3937,In_451,In_10);
and U3938 (N_3938,In_55,In_120);
and U3939 (N_3939,In_485,In_856);
or U3940 (N_3940,In_988,In_254);
nand U3941 (N_3941,In_410,In_175);
or U3942 (N_3942,In_930,In_125);
nor U3943 (N_3943,In_426,In_640);
nand U3944 (N_3944,In_666,In_66);
nand U3945 (N_3945,In_478,In_34);
or U3946 (N_3946,In_152,In_634);
and U3947 (N_3947,In_595,In_248);
nand U3948 (N_3948,In_809,In_369);
and U3949 (N_3949,In_608,In_880);
nand U3950 (N_3950,In_86,In_964);
or U3951 (N_3951,In_307,In_72);
nor U3952 (N_3952,In_79,In_311);
nand U3953 (N_3953,In_380,In_396);
and U3954 (N_3954,In_138,In_222);
or U3955 (N_3955,In_173,In_185);
and U3956 (N_3956,In_8,In_57);
or U3957 (N_3957,In_969,In_688);
and U3958 (N_3958,In_32,In_342);
and U3959 (N_3959,In_272,In_697);
and U3960 (N_3960,In_318,In_759);
nand U3961 (N_3961,In_463,In_958);
nor U3962 (N_3962,In_743,In_775);
or U3963 (N_3963,In_469,In_24);
or U3964 (N_3964,In_797,In_110);
nor U3965 (N_3965,In_703,In_678);
or U3966 (N_3966,In_682,In_276);
nand U3967 (N_3967,In_304,In_735);
or U3968 (N_3968,In_995,In_451);
nor U3969 (N_3969,In_774,In_157);
and U3970 (N_3970,In_0,In_182);
nor U3971 (N_3971,In_754,In_725);
nand U3972 (N_3972,In_376,In_291);
nor U3973 (N_3973,In_346,In_690);
and U3974 (N_3974,In_256,In_616);
nand U3975 (N_3975,In_699,In_847);
nand U3976 (N_3976,In_638,In_33);
nor U3977 (N_3977,In_862,In_979);
nand U3978 (N_3978,In_202,In_735);
or U3979 (N_3979,In_255,In_727);
nor U3980 (N_3980,In_457,In_601);
or U3981 (N_3981,In_225,In_722);
or U3982 (N_3982,In_454,In_498);
and U3983 (N_3983,In_54,In_654);
nor U3984 (N_3984,In_838,In_478);
and U3985 (N_3985,In_560,In_42);
nor U3986 (N_3986,In_625,In_161);
nand U3987 (N_3987,In_282,In_205);
or U3988 (N_3988,In_805,In_305);
nor U3989 (N_3989,In_360,In_642);
and U3990 (N_3990,In_370,In_682);
nor U3991 (N_3991,In_688,In_998);
and U3992 (N_3992,In_803,In_278);
nor U3993 (N_3993,In_93,In_258);
or U3994 (N_3994,In_683,In_520);
nor U3995 (N_3995,In_257,In_197);
nand U3996 (N_3996,In_101,In_940);
nor U3997 (N_3997,In_399,In_274);
or U3998 (N_3998,In_322,In_295);
nand U3999 (N_3999,In_154,In_424);
and U4000 (N_4000,In_237,In_194);
and U4001 (N_4001,In_467,In_682);
and U4002 (N_4002,In_335,In_521);
and U4003 (N_4003,In_382,In_823);
or U4004 (N_4004,In_990,In_388);
nand U4005 (N_4005,In_601,In_729);
nand U4006 (N_4006,In_714,In_296);
and U4007 (N_4007,In_138,In_459);
nor U4008 (N_4008,In_430,In_635);
and U4009 (N_4009,In_178,In_243);
or U4010 (N_4010,In_250,In_246);
nor U4011 (N_4011,In_279,In_373);
or U4012 (N_4012,In_275,In_833);
and U4013 (N_4013,In_508,In_423);
and U4014 (N_4014,In_188,In_590);
and U4015 (N_4015,In_24,In_589);
nor U4016 (N_4016,In_226,In_497);
nor U4017 (N_4017,In_275,In_939);
or U4018 (N_4018,In_621,In_775);
nand U4019 (N_4019,In_57,In_127);
nand U4020 (N_4020,In_704,In_148);
nor U4021 (N_4021,In_721,In_958);
nor U4022 (N_4022,In_85,In_864);
nand U4023 (N_4023,In_59,In_145);
and U4024 (N_4024,In_93,In_194);
nand U4025 (N_4025,In_583,In_236);
nor U4026 (N_4026,In_716,In_409);
and U4027 (N_4027,In_132,In_315);
nand U4028 (N_4028,In_283,In_892);
and U4029 (N_4029,In_392,In_898);
nor U4030 (N_4030,In_332,In_88);
nor U4031 (N_4031,In_209,In_728);
or U4032 (N_4032,In_627,In_491);
nand U4033 (N_4033,In_890,In_622);
nor U4034 (N_4034,In_28,In_982);
or U4035 (N_4035,In_310,In_605);
or U4036 (N_4036,In_611,In_253);
nor U4037 (N_4037,In_224,In_984);
or U4038 (N_4038,In_848,In_761);
and U4039 (N_4039,In_331,In_931);
and U4040 (N_4040,In_622,In_683);
nand U4041 (N_4041,In_120,In_557);
nand U4042 (N_4042,In_432,In_868);
and U4043 (N_4043,In_526,In_957);
nand U4044 (N_4044,In_77,In_991);
nor U4045 (N_4045,In_673,In_868);
nor U4046 (N_4046,In_863,In_220);
and U4047 (N_4047,In_930,In_770);
and U4048 (N_4048,In_670,In_203);
and U4049 (N_4049,In_33,In_830);
nand U4050 (N_4050,In_375,In_619);
nor U4051 (N_4051,In_987,In_763);
nor U4052 (N_4052,In_483,In_364);
nand U4053 (N_4053,In_729,In_939);
or U4054 (N_4054,In_371,In_145);
or U4055 (N_4055,In_248,In_806);
nor U4056 (N_4056,In_845,In_29);
and U4057 (N_4057,In_67,In_129);
and U4058 (N_4058,In_906,In_0);
nor U4059 (N_4059,In_582,In_697);
and U4060 (N_4060,In_574,In_661);
nand U4061 (N_4061,In_798,In_534);
nor U4062 (N_4062,In_519,In_996);
or U4063 (N_4063,In_8,In_820);
and U4064 (N_4064,In_735,In_846);
nor U4065 (N_4065,In_546,In_705);
nor U4066 (N_4066,In_802,In_902);
or U4067 (N_4067,In_62,In_454);
or U4068 (N_4068,In_924,In_879);
and U4069 (N_4069,In_494,In_171);
nor U4070 (N_4070,In_453,In_779);
nor U4071 (N_4071,In_626,In_576);
nand U4072 (N_4072,In_534,In_46);
nand U4073 (N_4073,In_59,In_678);
nor U4074 (N_4074,In_545,In_778);
or U4075 (N_4075,In_633,In_726);
or U4076 (N_4076,In_494,In_292);
nor U4077 (N_4077,In_551,In_100);
nor U4078 (N_4078,In_326,In_582);
nor U4079 (N_4079,In_391,In_904);
nand U4080 (N_4080,In_842,In_763);
and U4081 (N_4081,In_964,In_889);
and U4082 (N_4082,In_461,In_400);
or U4083 (N_4083,In_21,In_697);
nand U4084 (N_4084,In_475,In_535);
and U4085 (N_4085,In_708,In_103);
xor U4086 (N_4086,In_303,In_410);
or U4087 (N_4087,In_280,In_918);
nand U4088 (N_4088,In_828,In_179);
or U4089 (N_4089,In_214,In_699);
nand U4090 (N_4090,In_678,In_98);
nor U4091 (N_4091,In_397,In_418);
nor U4092 (N_4092,In_308,In_552);
nand U4093 (N_4093,In_584,In_194);
nand U4094 (N_4094,In_143,In_565);
and U4095 (N_4095,In_584,In_271);
or U4096 (N_4096,In_487,In_732);
nand U4097 (N_4097,In_287,In_515);
or U4098 (N_4098,In_660,In_513);
nor U4099 (N_4099,In_138,In_504);
and U4100 (N_4100,In_812,In_554);
nand U4101 (N_4101,In_317,In_283);
or U4102 (N_4102,In_997,In_330);
or U4103 (N_4103,In_832,In_194);
or U4104 (N_4104,In_639,In_763);
nor U4105 (N_4105,In_484,In_348);
and U4106 (N_4106,In_449,In_34);
nand U4107 (N_4107,In_954,In_235);
and U4108 (N_4108,In_761,In_173);
nor U4109 (N_4109,In_960,In_223);
nand U4110 (N_4110,In_358,In_196);
and U4111 (N_4111,In_212,In_855);
or U4112 (N_4112,In_330,In_774);
and U4113 (N_4113,In_301,In_148);
and U4114 (N_4114,In_885,In_558);
and U4115 (N_4115,In_588,In_871);
nand U4116 (N_4116,In_143,In_409);
nor U4117 (N_4117,In_763,In_552);
and U4118 (N_4118,In_350,In_965);
and U4119 (N_4119,In_831,In_182);
and U4120 (N_4120,In_924,In_42);
and U4121 (N_4121,In_369,In_520);
nor U4122 (N_4122,In_595,In_578);
nor U4123 (N_4123,In_189,In_771);
nand U4124 (N_4124,In_959,In_389);
nand U4125 (N_4125,In_134,In_179);
xnor U4126 (N_4126,In_178,In_729);
nand U4127 (N_4127,In_302,In_854);
or U4128 (N_4128,In_7,In_206);
nor U4129 (N_4129,In_800,In_883);
nor U4130 (N_4130,In_526,In_371);
nand U4131 (N_4131,In_630,In_513);
and U4132 (N_4132,In_302,In_278);
nand U4133 (N_4133,In_39,In_358);
xnor U4134 (N_4134,In_910,In_526);
and U4135 (N_4135,In_331,In_981);
nand U4136 (N_4136,In_418,In_730);
or U4137 (N_4137,In_495,In_319);
and U4138 (N_4138,In_295,In_344);
and U4139 (N_4139,In_617,In_157);
and U4140 (N_4140,In_846,In_245);
nand U4141 (N_4141,In_268,In_736);
nand U4142 (N_4142,In_35,In_470);
or U4143 (N_4143,In_859,In_588);
nand U4144 (N_4144,In_251,In_998);
or U4145 (N_4145,In_451,In_337);
and U4146 (N_4146,In_96,In_726);
and U4147 (N_4147,In_270,In_935);
or U4148 (N_4148,In_795,In_619);
or U4149 (N_4149,In_302,In_939);
nor U4150 (N_4150,In_916,In_207);
or U4151 (N_4151,In_73,In_281);
nand U4152 (N_4152,In_267,In_337);
nand U4153 (N_4153,In_192,In_250);
and U4154 (N_4154,In_459,In_999);
and U4155 (N_4155,In_926,In_272);
or U4156 (N_4156,In_405,In_360);
nand U4157 (N_4157,In_398,In_126);
and U4158 (N_4158,In_265,In_954);
or U4159 (N_4159,In_822,In_893);
nand U4160 (N_4160,In_558,In_380);
nand U4161 (N_4161,In_667,In_108);
nand U4162 (N_4162,In_91,In_648);
and U4163 (N_4163,In_63,In_984);
and U4164 (N_4164,In_430,In_54);
and U4165 (N_4165,In_883,In_753);
and U4166 (N_4166,In_353,In_217);
nand U4167 (N_4167,In_68,In_193);
nor U4168 (N_4168,In_408,In_420);
and U4169 (N_4169,In_58,In_942);
and U4170 (N_4170,In_408,In_564);
nand U4171 (N_4171,In_263,In_713);
or U4172 (N_4172,In_890,In_9);
and U4173 (N_4173,In_739,In_968);
or U4174 (N_4174,In_764,In_448);
or U4175 (N_4175,In_273,In_71);
or U4176 (N_4176,In_431,In_443);
and U4177 (N_4177,In_775,In_427);
nand U4178 (N_4178,In_729,In_146);
and U4179 (N_4179,In_111,In_410);
nor U4180 (N_4180,In_643,In_980);
or U4181 (N_4181,In_958,In_315);
and U4182 (N_4182,In_707,In_444);
and U4183 (N_4183,In_16,In_697);
nor U4184 (N_4184,In_176,In_919);
nor U4185 (N_4185,In_983,In_529);
and U4186 (N_4186,In_935,In_763);
xor U4187 (N_4187,In_737,In_326);
or U4188 (N_4188,In_566,In_802);
or U4189 (N_4189,In_513,In_385);
and U4190 (N_4190,In_586,In_555);
or U4191 (N_4191,In_809,In_387);
or U4192 (N_4192,In_965,In_751);
nor U4193 (N_4193,In_263,In_970);
and U4194 (N_4194,In_526,In_462);
or U4195 (N_4195,In_628,In_444);
nor U4196 (N_4196,In_758,In_414);
and U4197 (N_4197,In_589,In_471);
or U4198 (N_4198,In_296,In_742);
nor U4199 (N_4199,In_195,In_610);
and U4200 (N_4200,In_436,In_529);
nand U4201 (N_4201,In_723,In_725);
and U4202 (N_4202,In_37,In_251);
or U4203 (N_4203,In_617,In_702);
nor U4204 (N_4204,In_380,In_304);
nor U4205 (N_4205,In_76,In_5);
or U4206 (N_4206,In_215,In_272);
nand U4207 (N_4207,In_855,In_105);
or U4208 (N_4208,In_351,In_966);
or U4209 (N_4209,In_493,In_471);
nor U4210 (N_4210,In_181,In_504);
and U4211 (N_4211,In_631,In_320);
nor U4212 (N_4212,In_279,In_323);
and U4213 (N_4213,In_70,In_529);
or U4214 (N_4214,In_96,In_240);
or U4215 (N_4215,In_566,In_529);
and U4216 (N_4216,In_910,In_34);
or U4217 (N_4217,In_172,In_866);
nor U4218 (N_4218,In_877,In_190);
or U4219 (N_4219,In_760,In_173);
or U4220 (N_4220,In_475,In_739);
nand U4221 (N_4221,In_994,In_523);
and U4222 (N_4222,In_759,In_748);
and U4223 (N_4223,In_117,In_413);
nand U4224 (N_4224,In_766,In_254);
and U4225 (N_4225,In_261,In_213);
and U4226 (N_4226,In_679,In_833);
or U4227 (N_4227,In_633,In_471);
nor U4228 (N_4228,In_320,In_646);
nand U4229 (N_4229,In_973,In_449);
and U4230 (N_4230,In_992,In_143);
nor U4231 (N_4231,In_146,In_542);
or U4232 (N_4232,In_319,In_500);
nor U4233 (N_4233,In_385,In_830);
or U4234 (N_4234,In_981,In_61);
nand U4235 (N_4235,In_944,In_401);
or U4236 (N_4236,In_780,In_634);
and U4237 (N_4237,In_906,In_409);
and U4238 (N_4238,In_363,In_490);
nand U4239 (N_4239,In_854,In_11);
or U4240 (N_4240,In_566,In_20);
nand U4241 (N_4241,In_106,In_920);
nor U4242 (N_4242,In_85,In_157);
nor U4243 (N_4243,In_30,In_550);
nor U4244 (N_4244,In_430,In_601);
nand U4245 (N_4245,In_672,In_103);
nand U4246 (N_4246,In_741,In_75);
or U4247 (N_4247,In_761,In_726);
or U4248 (N_4248,In_862,In_912);
nand U4249 (N_4249,In_406,In_819);
nand U4250 (N_4250,In_991,In_600);
nor U4251 (N_4251,In_34,In_968);
nand U4252 (N_4252,In_862,In_709);
or U4253 (N_4253,In_783,In_115);
nand U4254 (N_4254,In_119,In_260);
nand U4255 (N_4255,In_574,In_373);
nor U4256 (N_4256,In_580,In_214);
or U4257 (N_4257,In_616,In_352);
nor U4258 (N_4258,In_410,In_825);
nor U4259 (N_4259,In_725,In_843);
nand U4260 (N_4260,In_243,In_128);
or U4261 (N_4261,In_81,In_545);
and U4262 (N_4262,In_700,In_111);
nand U4263 (N_4263,In_251,In_517);
or U4264 (N_4264,In_572,In_483);
nor U4265 (N_4265,In_196,In_642);
or U4266 (N_4266,In_176,In_694);
nand U4267 (N_4267,In_844,In_218);
or U4268 (N_4268,In_242,In_540);
and U4269 (N_4269,In_504,In_543);
nand U4270 (N_4270,In_68,In_101);
nor U4271 (N_4271,In_715,In_235);
nor U4272 (N_4272,In_50,In_782);
nand U4273 (N_4273,In_85,In_736);
and U4274 (N_4274,In_761,In_343);
or U4275 (N_4275,In_141,In_694);
nor U4276 (N_4276,In_607,In_205);
nand U4277 (N_4277,In_293,In_931);
nor U4278 (N_4278,In_48,In_879);
or U4279 (N_4279,In_136,In_696);
nand U4280 (N_4280,In_888,In_848);
and U4281 (N_4281,In_754,In_949);
nor U4282 (N_4282,In_131,In_377);
and U4283 (N_4283,In_126,In_713);
and U4284 (N_4284,In_994,In_534);
nand U4285 (N_4285,In_17,In_252);
or U4286 (N_4286,In_579,In_857);
and U4287 (N_4287,In_502,In_887);
nor U4288 (N_4288,In_274,In_926);
and U4289 (N_4289,In_996,In_130);
nor U4290 (N_4290,In_824,In_322);
or U4291 (N_4291,In_912,In_691);
and U4292 (N_4292,In_270,In_856);
nand U4293 (N_4293,In_364,In_311);
nor U4294 (N_4294,In_75,In_206);
nand U4295 (N_4295,In_543,In_929);
or U4296 (N_4296,In_684,In_759);
and U4297 (N_4297,In_842,In_719);
nand U4298 (N_4298,In_489,In_136);
and U4299 (N_4299,In_946,In_884);
or U4300 (N_4300,In_387,In_895);
nor U4301 (N_4301,In_336,In_498);
or U4302 (N_4302,In_876,In_152);
and U4303 (N_4303,In_272,In_689);
nand U4304 (N_4304,In_712,In_539);
and U4305 (N_4305,In_922,In_54);
or U4306 (N_4306,In_379,In_188);
nand U4307 (N_4307,In_464,In_378);
nor U4308 (N_4308,In_105,In_403);
nor U4309 (N_4309,In_692,In_350);
or U4310 (N_4310,In_828,In_996);
or U4311 (N_4311,In_633,In_679);
or U4312 (N_4312,In_368,In_671);
and U4313 (N_4313,In_616,In_143);
nand U4314 (N_4314,In_919,In_142);
and U4315 (N_4315,In_671,In_848);
xor U4316 (N_4316,In_857,In_384);
nor U4317 (N_4317,In_768,In_411);
nand U4318 (N_4318,In_530,In_379);
or U4319 (N_4319,In_845,In_19);
and U4320 (N_4320,In_273,In_955);
nor U4321 (N_4321,In_754,In_218);
or U4322 (N_4322,In_204,In_520);
or U4323 (N_4323,In_382,In_50);
or U4324 (N_4324,In_167,In_289);
nand U4325 (N_4325,In_191,In_90);
and U4326 (N_4326,In_373,In_0);
and U4327 (N_4327,In_16,In_56);
nor U4328 (N_4328,In_995,In_498);
or U4329 (N_4329,In_385,In_556);
and U4330 (N_4330,In_599,In_328);
nand U4331 (N_4331,In_799,In_699);
and U4332 (N_4332,In_373,In_964);
nor U4333 (N_4333,In_600,In_625);
and U4334 (N_4334,In_68,In_210);
nor U4335 (N_4335,In_606,In_467);
nand U4336 (N_4336,In_151,In_364);
nand U4337 (N_4337,In_822,In_874);
and U4338 (N_4338,In_672,In_178);
or U4339 (N_4339,In_439,In_61);
or U4340 (N_4340,In_225,In_955);
or U4341 (N_4341,In_986,In_247);
or U4342 (N_4342,In_596,In_482);
nor U4343 (N_4343,In_537,In_505);
nor U4344 (N_4344,In_388,In_245);
and U4345 (N_4345,In_796,In_123);
nand U4346 (N_4346,In_787,In_328);
or U4347 (N_4347,In_263,In_761);
or U4348 (N_4348,In_93,In_848);
nand U4349 (N_4349,In_571,In_21);
nor U4350 (N_4350,In_489,In_440);
nand U4351 (N_4351,In_101,In_380);
nor U4352 (N_4352,In_873,In_962);
nor U4353 (N_4353,In_345,In_243);
nor U4354 (N_4354,In_518,In_901);
or U4355 (N_4355,In_656,In_968);
nor U4356 (N_4356,In_299,In_525);
or U4357 (N_4357,In_686,In_370);
or U4358 (N_4358,In_830,In_933);
nand U4359 (N_4359,In_157,In_79);
and U4360 (N_4360,In_521,In_309);
or U4361 (N_4361,In_743,In_163);
nand U4362 (N_4362,In_256,In_471);
nand U4363 (N_4363,In_509,In_352);
nand U4364 (N_4364,In_879,In_903);
or U4365 (N_4365,In_258,In_634);
nand U4366 (N_4366,In_262,In_976);
and U4367 (N_4367,In_310,In_481);
nand U4368 (N_4368,In_119,In_675);
and U4369 (N_4369,In_895,In_763);
nand U4370 (N_4370,In_258,In_260);
nand U4371 (N_4371,In_194,In_874);
and U4372 (N_4372,In_697,In_158);
and U4373 (N_4373,In_888,In_775);
or U4374 (N_4374,In_86,In_991);
or U4375 (N_4375,In_514,In_876);
nand U4376 (N_4376,In_224,In_924);
nor U4377 (N_4377,In_845,In_427);
and U4378 (N_4378,In_51,In_197);
and U4379 (N_4379,In_625,In_322);
nand U4380 (N_4380,In_95,In_755);
nand U4381 (N_4381,In_503,In_808);
nand U4382 (N_4382,In_894,In_938);
or U4383 (N_4383,In_941,In_905);
and U4384 (N_4384,In_217,In_36);
nor U4385 (N_4385,In_367,In_138);
nor U4386 (N_4386,In_725,In_80);
nor U4387 (N_4387,In_80,In_993);
nand U4388 (N_4388,In_704,In_526);
nor U4389 (N_4389,In_180,In_695);
or U4390 (N_4390,In_712,In_307);
nor U4391 (N_4391,In_928,In_973);
and U4392 (N_4392,In_266,In_547);
nor U4393 (N_4393,In_543,In_893);
or U4394 (N_4394,In_320,In_812);
nand U4395 (N_4395,In_451,In_433);
nor U4396 (N_4396,In_802,In_851);
and U4397 (N_4397,In_779,In_772);
nor U4398 (N_4398,In_321,In_129);
or U4399 (N_4399,In_800,In_729);
nor U4400 (N_4400,In_575,In_164);
and U4401 (N_4401,In_426,In_551);
and U4402 (N_4402,In_232,In_923);
or U4403 (N_4403,In_910,In_917);
or U4404 (N_4404,In_676,In_144);
and U4405 (N_4405,In_182,In_104);
nand U4406 (N_4406,In_683,In_21);
and U4407 (N_4407,In_563,In_498);
nand U4408 (N_4408,In_348,In_958);
nor U4409 (N_4409,In_347,In_191);
nor U4410 (N_4410,In_150,In_894);
nor U4411 (N_4411,In_549,In_234);
nor U4412 (N_4412,In_696,In_629);
or U4413 (N_4413,In_489,In_212);
nand U4414 (N_4414,In_853,In_733);
and U4415 (N_4415,In_445,In_206);
or U4416 (N_4416,In_774,In_756);
or U4417 (N_4417,In_475,In_904);
nand U4418 (N_4418,In_359,In_652);
and U4419 (N_4419,In_542,In_297);
nand U4420 (N_4420,In_594,In_106);
nand U4421 (N_4421,In_639,In_183);
and U4422 (N_4422,In_180,In_88);
and U4423 (N_4423,In_256,In_830);
nand U4424 (N_4424,In_353,In_554);
xnor U4425 (N_4425,In_205,In_678);
or U4426 (N_4426,In_644,In_586);
nor U4427 (N_4427,In_70,In_489);
and U4428 (N_4428,In_794,In_70);
nand U4429 (N_4429,In_845,In_640);
nor U4430 (N_4430,In_651,In_647);
or U4431 (N_4431,In_904,In_281);
and U4432 (N_4432,In_346,In_308);
or U4433 (N_4433,In_171,In_367);
nand U4434 (N_4434,In_661,In_261);
or U4435 (N_4435,In_361,In_835);
nand U4436 (N_4436,In_802,In_738);
nor U4437 (N_4437,In_483,In_969);
nor U4438 (N_4438,In_757,In_198);
and U4439 (N_4439,In_251,In_159);
nor U4440 (N_4440,In_674,In_543);
and U4441 (N_4441,In_551,In_982);
or U4442 (N_4442,In_108,In_9);
and U4443 (N_4443,In_804,In_736);
nor U4444 (N_4444,In_37,In_371);
nor U4445 (N_4445,In_936,In_234);
or U4446 (N_4446,In_649,In_905);
nor U4447 (N_4447,In_497,In_22);
and U4448 (N_4448,In_302,In_824);
and U4449 (N_4449,In_107,In_315);
or U4450 (N_4450,In_181,In_338);
nand U4451 (N_4451,In_244,In_560);
or U4452 (N_4452,In_998,In_429);
nor U4453 (N_4453,In_839,In_731);
nand U4454 (N_4454,In_563,In_662);
nor U4455 (N_4455,In_699,In_980);
nor U4456 (N_4456,In_807,In_625);
xor U4457 (N_4457,In_938,In_362);
nor U4458 (N_4458,In_442,In_163);
and U4459 (N_4459,In_457,In_272);
or U4460 (N_4460,In_991,In_134);
or U4461 (N_4461,In_810,In_394);
nor U4462 (N_4462,In_390,In_556);
nand U4463 (N_4463,In_709,In_690);
nor U4464 (N_4464,In_989,In_808);
or U4465 (N_4465,In_800,In_826);
or U4466 (N_4466,In_676,In_337);
or U4467 (N_4467,In_308,In_74);
or U4468 (N_4468,In_221,In_581);
nand U4469 (N_4469,In_315,In_194);
nand U4470 (N_4470,In_706,In_683);
nor U4471 (N_4471,In_661,In_365);
nor U4472 (N_4472,In_982,In_285);
and U4473 (N_4473,In_719,In_912);
nand U4474 (N_4474,In_749,In_611);
or U4475 (N_4475,In_505,In_413);
and U4476 (N_4476,In_171,In_897);
or U4477 (N_4477,In_732,In_505);
or U4478 (N_4478,In_200,In_160);
xor U4479 (N_4479,In_458,In_455);
or U4480 (N_4480,In_889,In_87);
and U4481 (N_4481,In_600,In_135);
nand U4482 (N_4482,In_281,In_991);
nor U4483 (N_4483,In_66,In_145);
and U4484 (N_4484,In_224,In_37);
nor U4485 (N_4485,In_764,In_693);
nor U4486 (N_4486,In_471,In_899);
nor U4487 (N_4487,In_561,In_252);
and U4488 (N_4488,In_701,In_528);
or U4489 (N_4489,In_967,In_617);
and U4490 (N_4490,In_757,In_975);
and U4491 (N_4491,In_378,In_309);
xor U4492 (N_4492,In_166,In_124);
or U4493 (N_4493,In_146,In_932);
xnor U4494 (N_4494,In_331,In_881);
nand U4495 (N_4495,In_932,In_861);
nand U4496 (N_4496,In_240,In_475);
and U4497 (N_4497,In_911,In_928);
nand U4498 (N_4498,In_58,In_417);
or U4499 (N_4499,In_549,In_222);
nand U4500 (N_4500,In_763,In_96);
nor U4501 (N_4501,In_743,In_304);
nor U4502 (N_4502,In_146,In_136);
xnor U4503 (N_4503,In_607,In_2);
or U4504 (N_4504,In_198,In_827);
or U4505 (N_4505,In_368,In_429);
nor U4506 (N_4506,In_433,In_816);
nand U4507 (N_4507,In_395,In_231);
nand U4508 (N_4508,In_770,In_810);
nor U4509 (N_4509,In_159,In_712);
nor U4510 (N_4510,In_38,In_303);
nand U4511 (N_4511,In_986,In_838);
nor U4512 (N_4512,In_743,In_479);
or U4513 (N_4513,In_249,In_22);
nor U4514 (N_4514,In_124,In_41);
nor U4515 (N_4515,In_143,In_982);
and U4516 (N_4516,In_88,In_702);
or U4517 (N_4517,In_781,In_661);
and U4518 (N_4518,In_885,In_669);
and U4519 (N_4519,In_966,In_370);
and U4520 (N_4520,In_30,In_254);
nand U4521 (N_4521,In_525,In_197);
or U4522 (N_4522,In_687,In_342);
nor U4523 (N_4523,In_495,In_678);
nand U4524 (N_4524,In_53,In_336);
nor U4525 (N_4525,In_980,In_781);
nand U4526 (N_4526,In_556,In_754);
or U4527 (N_4527,In_172,In_414);
and U4528 (N_4528,In_411,In_702);
or U4529 (N_4529,In_390,In_660);
nor U4530 (N_4530,In_993,In_243);
and U4531 (N_4531,In_11,In_710);
nor U4532 (N_4532,In_121,In_568);
nor U4533 (N_4533,In_64,In_704);
or U4534 (N_4534,In_546,In_996);
nor U4535 (N_4535,In_53,In_132);
and U4536 (N_4536,In_434,In_886);
and U4537 (N_4537,In_509,In_371);
nor U4538 (N_4538,In_305,In_887);
nand U4539 (N_4539,In_834,In_981);
nand U4540 (N_4540,In_613,In_330);
and U4541 (N_4541,In_459,In_392);
or U4542 (N_4542,In_448,In_813);
or U4543 (N_4543,In_98,In_991);
nand U4544 (N_4544,In_472,In_281);
or U4545 (N_4545,In_797,In_7);
and U4546 (N_4546,In_308,In_609);
nor U4547 (N_4547,In_794,In_181);
nand U4548 (N_4548,In_891,In_40);
or U4549 (N_4549,In_700,In_781);
or U4550 (N_4550,In_820,In_379);
nand U4551 (N_4551,In_920,In_236);
and U4552 (N_4552,In_917,In_610);
nand U4553 (N_4553,In_616,In_683);
nand U4554 (N_4554,In_737,In_555);
nand U4555 (N_4555,In_768,In_1);
and U4556 (N_4556,In_359,In_239);
nand U4557 (N_4557,In_959,In_630);
nand U4558 (N_4558,In_901,In_762);
and U4559 (N_4559,In_878,In_321);
nor U4560 (N_4560,In_822,In_261);
nand U4561 (N_4561,In_920,In_105);
and U4562 (N_4562,In_727,In_639);
or U4563 (N_4563,In_486,In_110);
or U4564 (N_4564,In_865,In_33);
nor U4565 (N_4565,In_242,In_797);
or U4566 (N_4566,In_607,In_942);
and U4567 (N_4567,In_909,In_692);
or U4568 (N_4568,In_533,In_867);
or U4569 (N_4569,In_991,In_998);
nand U4570 (N_4570,In_470,In_487);
or U4571 (N_4571,In_334,In_650);
nand U4572 (N_4572,In_454,In_919);
and U4573 (N_4573,In_257,In_558);
and U4574 (N_4574,In_119,In_604);
nor U4575 (N_4575,In_837,In_322);
nand U4576 (N_4576,In_100,In_228);
or U4577 (N_4577,In_616,In_706);
nor U4578 (N_4578,In_655,In_733);
and U4579 (N_4579,In_647,In_574);
or U4580 (N_4580,In_837,In_547);
nand U4581 (N_4581,In_272,In_222);
and U4582 (N_4582,In_190,In_104);
nor U4583 (N_4583,In_362,In_968);
nor U4584 (N_4584,In_899,In_9);
nand U4585 (N_4585,In_167,In_6);
or U4586 (N_4586,In_642,In_155);
nand U4587 (N_4587,In_45,In_968);
nand U4588 (N_4588,In_204,In_718);
nor U4589 (N_4589,In_259,In_115);
and U4590 (N_4590,In_167,In_637);
or U4591 (N_4591,In_852,In_785);
nand U4592 (N_4592,In_426,In_902);
and U4593 (N_4593,In_680,In_336);
or U4594 (N_4594,In_369,In_656);
nor U4595 (N_4595,In_246,In_160);
nor U4596 (N_4596,In_63,In_9);
and U4597 (N_4597,In_600,In_364);
or U4598 (N_4598,In_282,In_695);
nor U4599 (N_4599,In_710,In_852);
and U4600 (N_4600,In_92,In_838);
nor U4601 (N_4601,In_685,In_207);
or U4602 (N_4602,In_12,In_673);
nor U4603 (N_4603,In_771,In_729);
nor U4604 (N_4604,In_579,In_770);
or U4605 (N_4605,In_944,In_527);
nor U4606 (N_4606,In_115,In_311);
or U4607 (N_4607,In_720,In_524);
nor U4608 (N_4608,In_330,In_875);
nand U4609 (N_4609,In_47,In_234);
or U4610 (N_4610,In_141,In_993);
or U4611 (N_4611,In_66,In_895);
or U4612 (N_4612,In_74,In_44);
nor U4613 (N_4613,In_685,In_35);
nand U4614 (N_4614,In_45,In_374);
nand U4615 (N_4615,In_837,In_898);
nand U4616 (N_4616,In_11,In_319);
or U4617 (N_4617,In_950,In_602);
nand U4618 (N_4618,In_107,In_575);
xor U4619 (N_4619,In_571,In_250);
or U4620 (N_4620,In_568,In_66);
nand U4621 (N_4621,In_754,In_169);
nand U4622 (N_4622,In_585,In_637);
or U4623 (N_4623,In_643,In_628);
or U4624 (N_4624,In_442,In_666);
or U4625 (N_4625,In_256,In_294);
nand U4626 (N_4626,In_698,In_841);
nand U4627 (N_4627,In_734,In_923);
and U4628 (N_4628,In_691,In_344);
nand U4629 (N_4629,In_152,In_739);
and U4630 (N_4630,In_779,In_295);
and U4631 (N_4631,In_531,In_24);
xor U4632 (N_4632,In_874,In_869);
or U4633 (N_4633,In_870,In_385);
and U4634 (N_4634,In_989,In_252);
nor U4635 (N_4635,In_328,In_486);
and U4636 (N_4636,In_153,In_198);
nand U4637 (N_4637,In_329,In_761);
nor U4638 (N_4638,In_857,In_302);
nor U4639 (N_4639,In_511,In_609);
and U4640 (N_4640,In_664,In_181);
or U4641 (N_4641,In_506,In_26);
nor U4642 (N_4642,In_465,In_287);
nand U4643 (N_4643,In_492,In_910);
nor U4644 (N_4644,In_389,In_932);
nand U4645 (N_4645,In_54,In_744);
or U4646 (N_4646,In_76,In_2);
and U4647 (N_4647,In_30,In_965);
and U4648 (N_4648,In_323,In_481);
nor U4649 (N_4649,In_75,In_781);
and U4650 (N_4650,In_483,In_10);
nand U4651 (N_4651,In_914,In_654);
and U4652 (N_4652,In_444,In_970);
nor U4653 (N_4653,In_610,In_329);
nand U4654 (N_4654,In_454,In_585);
nand U4655 (N_4655,In_72,In_361);
or U4656 (N_4656,In_697,In_148);
nand U4657 (N_4657,In_760,In_624);
and U4658 (N_4658,In_502,In_637);
and U4659 (N_4659,In_458,In_878);
and U4660 (N_4660,In_163,In_870);
nor U4661 (N_4661,In_341,In_611);
or U4662 (N_4662,In_310,In_913);
nor U4663 (N_4663,In_633,In_982);
and U4664 (N_4664,In_42,In_24);
nand U4665 (N_4665,In_817,In_217);
or U4666 (N_4666,In_985,In_217);
and U4667 (N_4667,In_652,In_693);
or U4668 (N_4668,In_798,In_126);
or U4669 (N_4669,In_593,In_570);
nand U4670 (N_4670,In_672,In_909);
nor U4671 (N_4671,In_231,In_249);
or U4672 (N_4672,In_287,In_330);
or U4673 (N_4673,In_148,In_456);
and U4674 (N_4674,In_244,In_579);
or U4675 (N_4675,In_599,In_527);
or U4676 (N_4676,In_939,In_327);
nor U4677 (N_4677,In_934,In_127);
and U4678 (N_4678,In_996,In_602);
or U4679 (N_4679,In_276,In_199);
nor U4680 (N_4680,In_862,In_432);
and U4681 (N_4681,In_324,In_308);
or U4682 (N_4682,In_732,In_827);
nand U4683 (N_4683,In_725,In_384);
nor U4684 (N_4684,In_623,In_615);
or U4685 (N_4685,In_327,In_128);
or U4686 (N_4686,In_609,In_359);
nand U4687 (N_4687,In_826,In_740);
nor U4688 (N_4688,In_439,In_758);
and U4689 (N_4689,In_218,In_155);
or U4690 (N_4690,In_887,In_706);
nand U4691 (N_4691,In_252,In_602);
nor U4692 (N_4692,In_343,In_85);
and U4693 (N_4693,In_664,In_519);
and U4694 (N_4694,In_361,In_413);
or U4695 (N_4695,In_228,In_126);
nor U4696 (N_4696,In_371,In_807);
or U4697 (N_4697,In_453,In_580);
nor U4698 (N_4698,In_477,In_599);
nor U4699 (N_4699,In_173,In_184);
and U4700 (N_4700,In_70,In_343);
or U4701 (N_4701,In_467,In_901);
and U4702 (N_4702,In_941,In_500);
and U4703 (N_4703,In_380,In_64);
and U4704 (N_4704,In_453,In_282);
and U4705 (N_4705,In_821,In_463);
or U4706 (N_4706,In_130,In_998);
xor U4707 (N_4707,In_578,In_588);
nor U4708 (N_4708,In_768,In_711);
or U4709 (N_4709,In_502,In_956);
and U4710 (N_4710,In_144,In_996);
or U4711 (N_4711,In_648,In_236);
and U4712 (N_4712,In_999,In_452);
nor U4713 (N_4713,In_119,In_444);
and U4714 (N_4714,In_700,In_439);
or U4715 (N_4715,In_467,In_79);
and U4716 (N_4716,In_189,In_173);
nor U4717 (N_4717,In_43,In_830);
and U4718 (N_4718,In_463,In_71);
nor U4719 (N_4719,In_8,In_649);
nor U4720 (N_4720,In_269,In_633);
nand U4721 (N_4721,In_918,In_365);
or U4722 (N_4722,In_945,In_218);
or U4723 (N_4723,In_227,In_447);
nand U4724 (N_4724,In_798,In_65);
or U4725 (N_4725,In_671,In_450);
or U4726 (N_4726,In_439,In_772);
or U4727 (N_4727,In_499,In_304);
nor U4728 (N_4728,In_509,In_350);
or U4729 (N_4729,In_608,In_770);
nand U4730 (N_4730,In_664,In_239);
nand U4731 (N_4731,In_952,In_993);
and U4732 (N_4732,In_120,In_251);
and U4733 (N_4733,In_179,In_86);
nand U4734 (N_4734,In_584,In_109);
and U4735 (N_4735,In_36,In_273);
or U4736 (N_4736,In_726,In_190);
or U4737 (N_4737,In_135,In_769);
nand U4738 (N_4738,In_967,In_288);
nand U4739 (N_4739,In_827,In_125);
or U4740 (N_4740,In_377,In_471);
and U4741 (N_4741,In_642,In_269);
or U4742 (N_4742,In_901,In_658);
or U4743 (N_4743,In_728,In_417);
or U4744 (N_4744,In_416,In_53);
nor U4745 (N_4745,In_269,In_224);
nor U4746 (N_4746,In_54,In_899);
nand U4747 (N_4747,In_795,In_123);
or U4748 (N_4748,In_880,In_383);
or U4749 (N_4749,In_315,In_189);
nand U4750 (N_4750,In_132,In_913);
and U4751 (N_4751,In_758,In_656);
nor U4752 (N_4752,In_268,In_587);
and U4753 (N_4753,In_741,In_699);
nand U4754 (N_4754,In_142,In_946);
nand U4755 (N_4755,In_385,In_516);
and U4756 (N_4756,In_573,In_717);
nand U4757 (N_4757,In_805,In_479);
nand U4758 (N_4758,In_660,In_843);
or U4759 (N_4759,In_301,In_536);
or U4760 (N_4760,In_676,In_288);
and U4761 (N_4761,In_688,In_769);
xor U4762 (N_4762,In_415,In_878);
nor U4763 (N_4763,In_829,In_512);
nor U4764 (N_4764,In_139,In_848);
nor U4765 (N_4765,In_71,In_999);
or U4766 (N_4766,In_69,In_468);
nand U4767 (N_4767,In_35,In_957);
nor U4768 (N_4768,In_613,In_687);
or U4769 (N_4769,In_94,In_540);
and U4770 (N_4770,In_307,In_814);
nand U4771 (N_4771,In_374,In_518);
nand U4772 (N_4772,In_882,In_744);
nor U4773 (N_4773,In_597,In_834);
and U4774 (N_4774,In_784,In_202);
nand U4775 (N_4775,In_802,In_353);
nor U4776 (N_4776,In_280,In_736);
nor U4777 (N_4777,In_868,In_982);
nand U4778 (N_4778,In_333,In_192);
and U4779 (N_4779,In_709,In_574);
and U4780 (N_4780,In_972,In_225);
or U4781 (N_4781,In_588,In_682);
nand U4782 (N_4782,In_478,In_263);
nor U4783 (N_4783,In_847,In_287);
nand U4784 (N_4784,In_732,In_395);
and U4785 (N_4785,In_340,In_332);
nand U4786 (N_4786,In_51,In_848);
nor U4787 (N_4787,In_597,In_117);
nand U4788 (N_4788,In_658,In_223);
nor U4789 (N_4789,In_876,In_494);
or U4790 (N_4790,In_947,In_897);
and U4791 (N_4791,In_125,In_298);
and U4792 (N_4792,In_31,In_46);
or U4793 (N_4793,In_497,In_493);
nand U4794 (N_4794,In_944,In_42);
nor U4795 (N_4795,In_215,In_297);
nor U4796 (N_4796,In_843,In_666);
nor U4797 (N_4797,In_212,In_75);
nor U4798 (N_4798,In_285,In_549);
and U4799 (N_4799,In_636,In_696);
nor U4800 (N_4800,In_775,In_852);
nor U4801 (N_4801,In_542,In_818);
nand U4802 (N_4802,In_992,In_186);
nor U4803 (N_4803,In_760,In_176);
or U4804 (N_4804,In_133,In_947);
nor U4805 (N_4805,In_206,In_125);
nor U4806 (N_4806,In_40,In_947);
nor U4807 (N_4807,In_304,In_629);
and U4808 (N_4808,In_740,In_580);
nand U4809 (N_4809,In_352,In_594);
nor U4810 (N_4810,In_718,In_373);
or U4811 (N_4811,In_891,In_164);
nand U4812 (N_4812,In_408,In_953);
or U4813 (N_4813,In_38,In_877);
nand U4814 (N_4814,In_577,In_674);
or U4815 (N_4815,In_179,In_599);
nor U4816 (N_4816,In_884,In_524);
nand U4817 (N_4817,In_188,In_281);
or U4818 (N_4818,In_145,In_763);
and U4819 (N_4819,In_412,In_964);
nand U4820 (N_4820,In_814,In_448);
nand U4821 (N_4821,In_945,In_978);
nor U4822 (N_4822,In_125,In_829);
or U4823 (N_4823,In_684,In_60);
nor U4824 (N_4824,In_628,In_896);
or U4825 (N_4825,In_947,In_723);
or U4826 (N_4826,In_495,In_209);
and U4827 (N_4827,In_294,In_53);
and U4828 (N_4828,In_119,In_798);
xnor U4829 (N_4829,In_646,In_801);
nor U4830 (N_4830,In_730,In_587);
nand U4831 (N_4831,In_86,In_132);
or U4832 (N_4832,In_130,In_577);
and U4833 (N_4833,In_706,In_908);
nor U4834 (N_4834,In_874,In_747);
nor U4835 (N_4835,In_975,In_883);
nand U4836 (N_4836,In_420,In_212);
and U4837 (N_4837,In_276,In_553);
nand U4838 (N_4838,In_138,In_572);
and U4839 (N_4839,In_594,In_221);
nand U4840 (N_4840,In_119,In_456);
nor U4841 (N_4841,In_442,In_726);
nor U4842 (N_4842,In_194,In_867);
and U4843 (N_4843,In_624,In_258);
or U4844 (N_4844,In_100,In_187);
and U4845 (N_4845,In_110,In_246);
nand U4846 (N_4846,In_857,In_896);
nor U4847 (N_4847,In_80,In_374);
nand U4848 (N_4848,In_390,In_632);
or U4849 (N_4849,In_674,In_634);
nand U4850 (N_4850,In_571,In_768);
and U4851 (N_4851,In_872,In_617);
and U4852 (N_4852,In_444,In_779);
nand U4853 (N_4853,In_670,In_259);
nor U4854 (N_4854,In_492,In_726);
nor U4855 (N_4855,In_894,In_754);
nand U4856 (N_4856,In_545,In_803);
or U4857 (N_4857,In_879,In_233);
and U4858 (N_4858,In_734,In_422);
nor U4859 (N_4859,In_820,In_238);
or U4860 (N_4860,In_964,In_233);
nand U4861 (N_4861,In_207,In_197);
and U4862 (N_4862,In_844,In_112);
and U4863 (N_4863,In_204,In_850);
or U4864 (N_4864,In_990,In_343);
nor U4865 (N_4865,In_849,In_790);
or U4866 (N_4866,In_643,In_409);
or U4867 (N_4867,In_778,In_385);
or U4868 (N_4868,In_690,In_31);
nand U4869 (N_4869,In_152,In_727);
nand U4870 (N_4870,In_114,In_365);
nor U4871 (N_4871,In_769,In_60);
and U4872 (N_4872,In_810,In_321);
or U4873 (N_4873,In_228,In_592);
nand U4874 (N_4874,In_977,In_219);
nor U4875 (N_4875,In_189,In_68);
nor U4876 (N_4876,In_324,In_139);
or U4877 (N_4877,In_457,In_183);
and U4878 (N_4878,In_479,In_214);
nor U4879 (N_4879,In_809,In_902);
and U4880 (N_4880,In_344,In_376);
nand U4881 (N_4881,In_453,In_21);
nand U4882 (N_4882,In_113,In_723);
or U4883 (N_4883,In_150,In_101);
nor U4884 (N_4884,In_167,In_262);
and U4885 (N_4885,In_564,In_602);
nand U4886 (N_4886,In_145,In_64);
and U4887 (N_4887,In_227,In_295);
and U4888 (N_4888,In_707,In_89);
and U4889 (N_4889,In_644,In_63);
and U4890 (N_4890,In_469,In_106);
and U4891 (N_4891,In_625,In_81);
and U4892 (N_4892,In_773,In_999);
and U4893 (N_4893,In_755,In_170);
nand U4894 (N_4894,In_933,In_491);
and U4895 (N_4895,In_355,In_844);
nor U4896 (N_4896,In_509,In_816);
or U4897 (N_4897,In_842,In_652);
nand U4898 (N_4898,In_969,In_928);
or U4899 (N_4899,In_181,In_688);
or U4900 (N_4900,In_357,In_469);
nor U4901 (N_4901,In_565,In_584);
or U4902 (N_4902,In_262,In_649);
nor U4903 (N_4903,In_532,In_567);
or U4904 (N_4904,In_311,In_641);
or U4905 (N_4905,In_556,In_54);
nand U4906 (N_4906,In_149,In_818);
nor U4907 (N_4907,In_197,In_77);
and U4908 (N_4908,In_366,In_213);
nand U4909 (N_4909,In_866,In_904);
and U4910 (N_4910,In_603,In_437);
or U4911 (N_4911,In_108,In_939);
and U4912 (N_4912,In_986,In_952);
nor U4913 (N_4913,In_788,In_87);
nand U4914 (N_4914,In_552,In_272);
and U4915 (N_4915,In_488,In_148);
or U4916 (N_4916,In_666,In_708);
and U4917 (N_4917,In_562,In_614);
nor U4918 (N_4918,In_376,In_515);
nand U4919 (N_4919,In_624,In_718);
and U4920 (N_4920,In_548,In_359);
nor U4921 (N_4921,In_122,In_632);
and U4922 (N_4922,In_963,In_367);
nand U4923 (N_4923,In_44,In_898);
or U4924 (N_4924,In_667,In_977);
nand U4925 (N_4925,In_726,In_283);
nor U4926 (N_4926,In_563,In_93);
nor U4927 (N_4927,In_129,In_638);
nor U4928 (N_4928,In_682,In_997);
or U4929 (N_4929,In_54,In_381);
or U4930 (N_4930,In_20,In_1);
nor U4931 (N_4931,In_120,In_193);
nand U4932 (N_4932,In_858,In_595);
nor U4933 (N_4933,In_940,In_397);
nand U4934 (N_4934,In_489,In_585);
and U4935 (N_4935,In_657,In_100);
nor U4936 (N_4936,In_927,In_98);
nor U4937 (N_4937,In_693,In_270);
nor U4938 (N_4938,In_337,In_222);
and U4939 (N_4939,In_0,In_762);
nor U4940 (N_4940,In_794,In_446);
or U4941 (N_4941,In_958,In_965);
and U4942 (N_4942,In_314,In_356);
or U4943 (N_4943,In_91,In_295);
nor U4944 (N_4944,In_427,In_232);
nor U4945 (N_4945,In_811,In_433);
and U4946 (N_4946,In_920,In_189);
or U4947 (N_4947,In_844,In_724);
nand U4948 (N_4948,In_204,In_72);
and U4949 (N_4949,In_810,In_881);
or U4950 (N_4950,In_148,In_955);
xnor U4951 (N_4951,In_939,In_958);
nor U4952 (N_4952,In_804,In_226);
nor U4953 (N_4953,In_91,In_576);
nand U4954 (N_4954,In_407,In_607);
and U4955 (N_4955,In_521,In_80);
and U4956 (N_4956,In_408,In_66);
and U4957 (N_4957,In_677,In_748);
and U4958 (N_4958,In_479,In_632);
nor U4959 (N_4959,In_407,In_44);
nor U4960 (N_4960,In_442,In_349);
nor U4961 (N_4961,In_858,In_725);
or U4962 (N_4962,In_512,In_346);
and U4963 (N_4963,In_270,In_241);
nand U4964 (N_4964,In_922,In_253);
nor U4965 (N_4965,In_892,In_713);
nor U4966 (N_4966,In_676,In_642);
nand U4967 (N_4967,In_547,In_916);
nor U4968 (N_4968,In_585,In_617);
or U4969 (N_4969,In_268,In_993);
nand U4970 (N_4970,In_35,In_890);
nor U4971 (N_4971,In_286,In_909);
or U4972 (N_4972,In_458,In_20);
and U4973 (N_4973,In_361,In_457);
nand U4974 (N_4974,In_419,In_828);
or U4975 (N_4975,In_801,In_995);
nand U4976 (N_4976,In_665,In_912);
and U4977 (N_4977,In_31,In_679);
and U4978 (N_4978,In_279,In_793);
and U4979 (N_4979,In_537,In_80);
nand U4980 (N_4980,In_840,In_550);
nor U4981 (N_4981,In_114,In_706);
nor U4982 (N_4982,In_823,In_799);
nand U4983 (N_4983,In_474,In_257);
and U4984 (N_4984,In_37,In_471);
or U4985 (N_4985,In_90,In_463);
nor U4986 (N_4986,In_292,In_653);
and U4987 (N_4987,In_640,In_54);
and U4988 (N_4988,In_678,In_650);
xnor U4989 (N_4989,In_773,In_143);
nor U4990 (N_4990,In_575,In_936);
nor U4991 (N_4991,In_101,In_826);
and U4992 (N_4992,In_229,In_155);
nor U4993 (N_4993,In_375,In_61);
or U4994 (N_4994,In_79,In_122);
nand U4995 (N_4995,In_554,In_641);
and U4996 (N_4996,In_901,In_81);
and U4997 (N_4997,In_894,In_270);
and U4998 (N_4998,In_14,In_417);
nor U4999 (N_4999,In_409,In_890);
nor U5000 (N_5000,N_947,N_1210);
nand U5001 (N_5001,N_4855,N_4911);
nor U5002 (N_5002,N_1261,N_2517);
or U5003 (N_5003,N_1147,N_975);
and U5004 (N_5004,N_794,N_2812);
xor U5005 (N_5005,N_4641,N_978);
nand U5006 (N_5006,N_3959,N_4785);
or U5007 (N_5007,N_4833,N_744);
nand U5008 (N_5008,N_2154,N_4440);
nor U5009 (N_5009,N_3910,N_3075);
nand U5010 (N_5010,N_871,N_4350);
nor U5011 (N_5011,N_3104,N_1958);
nor U5012 (N_5012,N_4314,N_3393);
and U5013 (N_5013,N_2087,N_3941);
or U5014 (N_5014,N_4149,N_1111);
and U5015 (N_5015,N_1616,N_3994);
or U5016 (N_5016,N_2222,N_184);
nand U5017 (N_5017,N_452,N_3659);
nor U5018 (N_5018,N_1380,N_3302);
and U5019 (N_5019,N_639,N_3477);
nor U5020 (N_5020,N_2740,N_4625);
or U5021 (N_5021,N_4604,N_2617);
or U5022 (N_5022,N_1513,N_3406);
or U5023 (N_5023,N_938,N_1893);
and U5024 (N_5024,N_4530,N_1570);
nand U5025 (N_5025,N_4005,N_4474);
nor U5026 (N_5026,N_2485,N_3399);
and U5027 (N_5027,N_3449,N_2065);
nor U5028 (N_5028,N_278,N_4402);
nor U5029 (N_5029,N_2986,N_4082);
nand U5030 (N_5030,N_795,N_3587);
nand U5031 (N_5031,N_3598,N_2990);
nor U5032 (N_5032,N_2304,N_2531);
nand U5033 (N_5033,N_126,N_842);
nor U5034 (N_5034,N_333,N_757);
or U5035 (N_5035,N_4268,N_3632);
nor U5036 (N_5036,N_1586,N_2596);
nor U5037 (N_5037,N_2206,N_4171);
nor U5038 (N_5038,N_1449,N_3433);
and U5039 (N_5039,N_3546,N_1177);
nor U5040 (N_5040,N_1233,N_738);
and U5041 (N_5041,N_1443,N_2476);
nand U5042 (N_5042,N_3432,N_1678);
or U5043 (N_5043,N_3019,N_4122);
and U5044 (N_5044,N_432,N_2980);
or U5045 (N_5045,N_3968,N_3863);
nor U5046 (N_5046,N_3115,N_4098);
nand U5047 (N_5047,N_3760,N_53);
and U5048 (N_5048,N_2686,N_2984);
or U5049 (N_5049,N_2816,N_2032);
or U5050 (N_5050,N_125,N_1218);
nand U5051 (N_5051,N_1707,N_260);
nor U5052 (N_5052,N_1734,N_4483);
and U5053 (N_5053,N_1219,N_2766);
or U5054 (N_5054,N_4512,N_4009);
nor U5055 (N_5055,N_1230,N_2139);
nand U5056 (N_5056,N_1687,N_1390);
or U5057 (N_5057,N_73,N_2633);
nand U5058 (N_5058,N_1000,N_1247);
or U5059 (N_5059,N_4730,N_3146);
nor U5060 (N_5060,N_4822,N_1151);
nand U5061 (N_5061,N_711,N_571);
or U5062 (N_5062,N_4576,N_2512);
and U5063 (N_5063,N_4112,N_3502);
and U5064 (N_5064,N_1714,N_3699);
nor U5065 (N_5065,N_1669,N_1292);
nand U5066 (N_5066,N_1942,N_4254);
or U5067 (N_5067,N_2684,N_1325);
or U5068 (N_5068,N_3703,N_820);
and U5069 (N_5069,N_2580,N_941);
nor U5070 (N_5070,N_1319,N_547);
or U5071 (N_5071,N_1766,N_564);
nand U5072 (N_5072,N_2395,N_3772);
and U5073 (N_5073,N_4482,N_3023);
or U5074 (N_5074,N_1432,N_3386);
nor U5075 (N_5075,N_2142,N_81);
or U5076 (N_5076,N_1618,N_2760);
nand U5077 (N_5077,N_2377,N_2870);
nor U5078 (N_5078,N_4523,N_4374);
nand U5079 (N_5079,N_2040,N_2286);
or U5080 (N_5080,N_2762,N_3780);
and U5081 (N_5081,N_1485,N_4176);
or U5082 (N_5082,N_4917,N_387);
or U5083 (N_5083,N_4330,N_3591);
nand U5084 (N_5084,N_3882,N_3912);
and U5085 (N_5085,N_2358,N_4167);
and U5086 (N_5086,N_3915,N_2179);
nand U5087 (N_5087,N_2058,N_4362);
nand U5088 (N_5088,N_289,N_4748);
or U5089 (N_5089,N_455,N_2481);
nand U5090 (N_5090,N_4449,N_1953);
and U5091 (N_5091,N_1551,N_4277);
nand U5092 (N_5092,N_2938,N_1100);
nor U5093 (N_5093,N_2078,N_1662);
nor U5094 (N_5094,N_3745,N_1491);
or U5095 (N_5095,N_238,N_4749);
nand U5096 (N_5096,N_1280,N_745);
nand U5097 (N_5097,N_1540,N_3131);
and U5098 (N_5098,N_4629,N_3499);
and U5099 (N_5099,N_4455,N_695);
or U5100 (N_5100,N_106,N_4670);
or U5101 (N_5101,N_4237,N_1289);
or U5102 (N_5102,N_228,N_2759);
and U5103 (N_5103,N_3400,N_4695);
nor U5104 (N_5104,N_2153,N_2814);
and U5105 (N_5105,N_678,N_191);
and U5106 (N_5106,N_3479,N_594);
and U5107 (N_5107,N_2082,N_358);
or U5108 (N_5108,N_4764,N_2627);
or U5109 (N_5109,N_1308,N_1153);
or U5110 (N_5110,N_194,N_3308);
nand U5111 (N_5111,N_2002,N_1342);
and U5112 (N_5112,N_3349,N_1822);
nand U5113 (N_5113,N_138,N_850);
and U5114 (N_5114,N_2346,N_171);
and U5115 (N_5115,N_800,N_120);
or U5116 (N_5116,N_3181,N_1691);
nand U5117 (N_5117,N_3648,N_4049);
or U5118 (N_5118,N_4377,N_2510);
and U5119 (N_5119,N_2347,N_857);
nor U5120 (N_5120,N_837,N_62);
or U5121 (N_5121,N_3306,N_4983);
nand U5122 (N_5122,N_3036,N_4419);
nand U5123 (N_5123,N_4241,N_3493);
nand U5124 (N_5124,N_1157,N_1811);
and U5125 (N_5125,N_1050,N_4635);
nor U5126 (N_5126,N_2190,N_3113);
nor U5127 (N_5127,N_270,N_3784);
or U5128 (N_5128,N_2080,N_1413);
or U5129 (N_5129,N_4216,N_2325);
or U5130 (N_5130,N_1383,N_3260);
nand U5131 (N_5131,N_4899,N_3750);
and U5132 (N_5132,N_4376,N_99);
or U5133 (N_5133,N_4024,N_2429);
nor U5134 (N_5134,N_4729,N_3582);
nor U5135 (N_5135,N_1988,N_3685);
nor U5136 (N_5136,N_1915,N_3478);
nand U5137 (N_5137,N_763,N_1730);
nand U5138 (N_5138,N_1974,N_4008);
nand U5139 (N_5139,N_2319,N_4527);
or U5140 (N_5140,N_1658,N_974);
nand U5141 (N_5141,N_3663,N_2635);
nor U5142 (N_5142,N_1259,N_4018);
nand U5143 (N_5143,N_3342,N_2436);
nor U5144 (N_5144,N_1828,N_4838);
nand U5145 (N_5145,N_1183,N_2782);
nand U5146 (N_5146,N_685,N_1436);
and U5147 (N_5147,N_2774,N_1220);
nor U5148 (N_5148,N_3518,N_3027);
nor U5149 (N_5149,N_2342,N_4579);
and U5150 (N_5150,N_488,N_288);
or U5151 (N_5151,N_2114,N_10);
and U5152 (N_5152,N_2932,N_2267);
or U5153 (N_5153,N_4524,N_652);
nand U5154 (N_5154,N_254,N_3535);
xor U5155 (N_5155,N_665,N_3641);
or U5156 (N_5156,N_2212,N_1320);
nand U5157 (N_5157,N_2471,N_244);
nand U5158 (N_5158,N_1339,N_2334);
nor U5159 (N_5159,N_1706,N_2937);
or U5160 (N_5160,N_926,N_4674);
nand U5161 (N_5161,N_3021,N_1655);
nor U5162 (N_5162,N_863,N_4133);
nor U5163 (N_5163,N_2605,N_3822);
nand U5164 (N_5164,N_3491,N_1411);
and U5165 (N_5165,N_2900,N_3076);
nand U5166 (N_5166,N_876,N_2350);
nand U5167 (N_5167,N_3025,N_1267);
and U5168 (N_5168,N_1047,N_4708);
or U5169 (N_5169,N_4487,N_1978);
nand U5170 (N_5170,N_2732,N_4079);
xor U5171 (N_5171,N_2493,N_672);
nor U5172 (N_5172,N_2682,N_3480);
nor U5173 (N_5173,N_508,N_3683);
or U5174 (N_5174,N_2243,N_1797);
nor U5175 (N_5175,N_1381,N_4484);
or U5176 (N_5176,N_2752,N_2768);
and U5177 (N_5177,N_1187,N_1429);
or U5178 (N_5178,N_4568,N_4584);
nand U5179 (N_5179,N_3544,N_4728);
or U5180 (N_5180,N_243,N_4818);
nand U5181 (N_5181,N_4824,N_1639);
nand U5182 (N_5182,N_168,N_3837);
nor U5183 (N_5183,N_345,N_1060);
nor U5184 (N_5184,N_1067,N_3788);
nor U5185 (N_5185,N_764,N_761);
nor U5186 (N_5186,N_1084,N_1989);
or U5187 (N_5187,N_3394,N_3294);
nand U5188 (N_5188,N_4348,N_3531);
nand U5189 (N_5189,N_4551,N_4780);
nand U5190 (N_5190,N_1331,N_1577);
or U5191 (N_5191,N_155,N_2841);
nor U5192 (N_5192,N_537,N_2291);
nand U5193 (N_5193,N_1468,N_439);
and U5194 (N_5194,N_4373,N_50);
or U5195 (N_5195,N_1727,N_220);
nor U5196 (N_5196,N_1832,N_186);
and U5197 (N_5197,N_3093,N_4944);
and U5198 (N_5198,N_4634,N_1200);
nor U5199 (N_5199,N_881,N_3442);
or U5200 (N_5200,N_1037,N_825);
or U5201 (N_5201,N_1098,N_2166);
nand U5202 (N_5202,N_4364,N_715);
nand U5203 (N_5203,N_914,N_485);
or U5204 (N_5204,N_4581,N_1911);
or U5205 (N_5205,N_2445,N_1216);
and U5206 (N_5206,N_3127,N_2897);
or U5207 (N_5207,N_3921,N_4801);
nor U5208 (N_5208,N_35,N_3561);
or U5209 (N_5209,N_4520,N_3527);
and U5210 (N_5210,N_2951,N_2138);
or U5211 (N_5211,N_3835,N_72);
nand U5212 (N_5212,N_3424,N_4074);
or U5213 (N_5213,N_2117,N_1025);
and U5214 (N_5214,N_4195,N_4808);
nor U5215 (N_5215,N_1640,N_2950);
or U5216 (N_5216,N_4918,N_4055);
nor U5217 (N_5217,N_4382,N_1791);
nand U5218 (N_5218,N_1099,N_1940);
and U5219 (N_5219,N_352,N_4211);
and U5220 (N_5220,N_1193,N_2368);
or U5221 (N_5221,N_421,N_573);
nand U5222 (N_5222,N_4323,N_4477);
nand U5223 (N_5223,N_1574,N_3376);
nand U5224 (N_5224,N_2503,N_2136);
and U5225 (N_5225,N_3147,N_2896);
or U5226 (N_5226,N_3483,N_2210);
or U5227 (N_5227,N_1161,N_897);
and U5228 (N_5228,N_15,N_1999);
nand U5229 (N_5229,N_4701,N_465);
and U5230 (N_5230,N_983,N_3734);
nor U5231 (N_5231,N_1124,N_1802);
and U5232 (N_5232,N_263,N_1189);
and U5233 (N_5233,N_1591,N_2149);
and U5234 (N_5234,N_1115,N_3830);
or U5235 (N_5235,N_3861,N_2533);
or U5236 (N_5236,N_1737,N_420);
or U5237 (N_5237,N_1985,N_4789);
nor U5238 (N_5238,N_686,N_1757);
or U5239 (N_5239,N_2828,N_3754);
nand U5240 (N_5240,N_2218,N_483);
xor U5241 (N_5241,N_4212,N_1938);
nor U5242 (N_5242,N_3794,N_287);
or U5243 (N_5243,N_3853,N_4718);
nand U5244 (N_5244,N_1769,N_3223);
or U5245 (N_5245,N_1906,N_3790);
nand U5246 (N_5246,N_1199,N_4933);
and U5247 (N_5247,N_2538,N_965);
nor U5248 (N_5248,N_3774,N_4193);
nor U5249 (N_5249,N_327,N_2246);
nor U5250 (N_5250,N_3049,N_1531);
nand U5251 (N_5251,N_2013,N_3680);
and U5252 (N_5252,N_2653,N_3571);
nor U5253 (N_5253,N_4346,N_645);
and U5254 (N_5254,N_1745,N_2671);
nor U5255 (N_5255,N_4452,N_480);
and U5256 (N_5256,N_4352,N_870);
nand U5257 (N_5257,N_1435,N_3566);
or U5258 (N_5258,N_1417,N_3196);
and U5259 (N_5259,N_179,N_153);
or U5260 (N_5260,N_606,N_4113);
nand U5261 (N_5261,N_2299,N_190);
nor U5262 (N_5262,N_4002,N_454);
nand U5263 (N_5263,N_1719,N_2922);
or U5264 (N_5264,N_4327,N_4578);
or U5265 (N_5265,N_739,N_621);
or U5266 (N_5266,N_3463,N_4906);
or U5267 (N_5267,N_4162,N_2844);
nand U5268 (N_5268,N_3567,N_2885);
and U5269 (N_5269,N_1993,N_3579);
nor U5270 (N_5270,N_641,N_2432);
and U5271 (N_5271,N_1445,N_4255);
or U5272 (N_5272,N_3966,N_2366);
nand U5273 (N_5273,N_4058,N_950);
nor U5274 (N_5274,N_796,N_2262);
or U5275 (N_5275,N_4329,N_3281);
nand U5276 (N_5276,N_616,N_1937);
and U5277 (N_5277,N_2796,N_2620);
nand U5278 (N_5278,N_4210,N_2124);
and U5279 (N_5279,N_22,N_2838);
nand U5280 (N_5280,N_2257,N_961);
nand U5281 (N_5281,N_3460,N_4588);
and U5282 (N_5282,N_4281,N_2854);
nor U5283 (N_5283,N_2738,N_3520);
nand U5284 (N_5284,N_538,N_2354);
or U5285 (N_5285,N_4639,N_4020);
and U5286 (N_5286,N_1345,N_4782);
nand U5287 (N_5287,N_4692,N_649);
or U5288 (N_5288,N_192,N_4138);
and U5289 (N_5289,N_3589,N_3005);
and U5290 (N_5290,N_1610,N_1130);
nor U5291 (N_5291,N_290,N_499);
nand U5292 (N_5292,N_3991,N_4083);
or U5293 (N_5293,N_3939,N_4198);
or U5294 (N_5294,N_75,N_3380);
and U5295 (N_5295,N_3954,N_3833);
nand U5296 (N_5296,N_3771,N_2526);
or U5297 (N_5297,N_3604,N_1856);
or U5298 (N_5298,N_2042,N_2193);
nor U5299 (N_5299,N_2349,N_3725);
or U5300 (N_5300,N_550,N_3961);
and U5301 (N_5301,N_4795,N_1555);
and U5302 (N_5302,N_2910,N_4868);
and U5303 (N_5303,N_1785,N_925);
xnor U5304 (N_5304,N_159,N_4820);
nor U5305 (N_5305,N_1410,N_316);
or U5306 (N_5306,N_446,N_3046);
nand U5307 (N_5307,N_1295,N_4644);
nand U5308 (N_5308,N_3585,N_1234);
or U5309 (N_5309,N_6,N_2359);
or U5310 (N_5310,N_3859,N_3462);
and U5311 (N_5311,N_2033,N_1677);
nand U5312 (N_5312,N_4598,N_3600);
nor U5313 (N_5313,N_580,N_2636);
and U5314 (N_5314,N_2448,N_3307);
nand U5315 (N_5315,N_4339,N_2601);
or U5316 (N_5316,N_4236,N_344);
and U5317 (N_5317,N_4776,N_3109);
and U5318 (N_5318,N_646,N_4228);
or U5319 (N_5319,N_2886,N_1431);
nand U5320 (N_5320,N_3201,N_1851);
nor U5321 (N_5321,N_1642,N_4128);
and U5322 (N_5322,N_3143,N_3576);
or U5323 (N_5323,N_2324,N_2869);
and U5324 (N_5324,N_2137,N_1321);
and U5325 (N_5325,N_617,N_1232);
nor U5326 (N_5326,N_4783,N_3423);
and U5327 (N_5327,N_2469,N_3695);
and U5328 (N_5328,N_2,N_2726);
or U5329 (N_5329,N_2789,N_2929);
nand U5330 (N_5330,N_4383,N_919);
and U5331 (N_5331,N_3679,N_4717);
nand U5332 (N_5332,N_2890,N_1996);
nor U5333 (N_5333,N_2985,N_4980);
and U5334 (N_5334,N_404,N_1961);
nor U5335 (N_5335,N_2098,N_3364);
and U5336 (N_5336,N_362,N_759);
nand U5337 (N_5337,N_375,N_4740);
and U5338 (N_5338,N_4586,N_4790);
or U5339 (N_5339,N_2808,N_2340);
nor U5340 (N_5340,N_3274,N_2848);
nor U5341 (N_5341,N_3615,N_567);
nor U5342 (N_5342,N_3940,N_2070);
nand U5343 (N_5343,N_2957,N_1090);
and U5344 (N_5344,N_648,N_110);
nor U5345 (N_5345,N_403,N_376);
and U5346 (N_5346,N_4769,N_964);
nor U5347 (N_5347,N_3316,N_4233);
and U5348 (N_5348,N_2468,N_2433);
nand U5349 (N_5349,N_883,N_3883);
nor U5350 (N_5350,N_2112,N_602);
nor U5351 (N_5351,N_2573,N_1945);
or U5352 (N_5352,N_1487,N_1708);
nor U5353 (N_5353,N_4461,N_3123);
and U5354 (N_5354,N_3461,N_2451);
nand U5355 (N_5355,N_3253,N_1164);
nor U5356 (N_5356,N_855,N_4556);
and U5357 (N_5357,N_4473,N_3536);
and U5358 (N_5358,N_3170,N_44);
nor U5359 (N_5359,N_2637,N_4539);
and U5360 (N_5360,N_3368,N_4444);
and U5361 (N_5361,N_109,N_4654);
or U5362 (N_5362,N_1501,N_2832);
nand U5363 (N_5363,N_3009,N_3978);
nand U5364 (N_5364,N_4156,N_3034);
nand U5365 (N_5365,N_2645,N_2045);
or U5366 (N_5366,N_3996,N_1516);
nor U5367 (N_5367,N_3211,N_4261);
nand U5368 (N_5368,N_4743,N_4939);
and U5369 (N_5369,N_748,N_2833);
nor U5370 (N_5370,N_1351,N_4612);
and U5371 (N_5371,N_1266,N_49);
or U5372 (N_5372,N_2083,N_4860);
and U5373 (N_5373,N_3373,N_497);
and U5374 (N_5374,N_4761,N_1182);
or U5375 (N_5375,N_4157,N_1593);
and U5376 (N_5376,N_4736,N_2908);
and U5377 (N_5377,N_777,N_4321);
nand U5378 (N_5378,N_4406,N_1076);
nor U5379 (N_5379,N_4033,N_3943);
nand U5380 (N_5380,N_3165,N_1524);
or U5381 (N_5381,N_1529,N_3669);
nand U5382 (N_5382,N_3168,N_980);
and U5383 (N_5383,N_3383,N_3033);
nand U5384 (N_5384,N_4519,N_3238);
and U5385 (N_5385,N_4945,N_3476);
or U5386 (N_5386,N_4777,N_3510);
or U5387 (N_5387,N_487,N_388);
or U5388 (N_5388,N_3574,N_1553);
or U5389 (N_5389,N_2550,N_1509);
or U5390 (N_5390,N_511,N_4132);
or U5391 (N_5391,N_1612,N_1348);
nand U5392 (N_5392,N_1852,N_4656);
and U5393 (N_5393,N_43,N_2113);
and U5394 (N_5394,N_956,N_304);
nor U5395 (N_5395,N_3155,N_3958);
or U5396 (N_5396,N_1519,N_4573);
and U5397 (N_5397,N_1235,N_4544);
nand U5398 (N_5398,N_4124,N_1256);
nand U5399 (N_5399,N_4472,N_1622);
or U5400 (N_5400,N_2464,N_1674);
and U5401 (N_5401,N_4505,N_4415);
or U5402 (N_5402,N_1672,N_654);
and U5403 (N_5403,N_4480,N_637);
and U5404 (N_5404,N_3649,N_1370);
or U5405 (N_5405,N_3178,N_4869);
and U5406 (N_5406,N_1855,N_312);
nand U5407 (N_5407,N_1185,N_285);
nand U5408 (N_5408,N_1843,N_907);
and U5409 (N_5409,N_4878,N_257);
or U5410 (N_5410,N_3800,N_3);
nor U5411 (N_5411,N_698,N_2919);
nand U5412 (N_5412,N_3272,N_127);
nand U5413 (N_5413,N_4199,N_2029);
and U5414 (N_5414,N_4711,N_3124);
and U5415 (N_5415,N_4290,N_1440);
nor U5416 (N_5416,N_4518,N_2453);
nand U5417 (N_5417,N_3553,N_3284);
nand U5418 (N_5418,N_4657,N_2125);
and U5419 (N_5419,N_2077,N_1777);
and U5420 (N_5420,N_2722,N_3533);
nand U5421 (N_5421,N_3638,N_137);
or U5422 (N_5422,N_3409,N_3095);
nor U5423 (N_5423,N_4072,N_3436);
or U5424 (N_5424,N_26,N_4227);
nand U5425 (N_5425,N_2827,N_4916);
nand U5426 (N_5426,N_2997,N_104);
and U5427 (N_5427,N_2901,N_866);
nor U5428 (N_5428,N_2442,N_1975);
nor U5429 (N_5429,N_4252,N_4197);
nand U5430 (N_5430,N_5,N_3041);
nand U5431 (N_5431,N_3700,N_408);
and U5432 (N_5432,N_979,N_3712);
nand U5433 (N_5433,N_1659,N_2096);
and U5434 (N_5434,N_4887,N_1633);
and U5435 (N_5435,N_4832,N_1213);
or U5436 (N_5436,N_681,N_1150);
nor U5437 (N_5437,N_3819,N_4204);
nor U5438 (N_5438,N_2912,N_47);
or U5439 (N_5439,N_3623,N_2184);
nor U5440 (N_5440,N_3551,N_4497);
or U5441 (N_5441,N_1464,N_1720);
nor U5442 (N_5442,N_4436,N_527);
or U5443 (N_5443,N_1631,N_3194);
or U5444 (N_5444,N_4226,N_1272);
nand U5445 (N_5445,N_48,N_4147);
nor U5446 (N_5446,N_526,N_4636);
or U5447 (N_5447,N_386,N_1916);
nor U5448 (N_5448,N_2805,N_2561);
and U5449 (N_5449,N_1424,N_3743);
or U5450 (N_5450,N_4966,N_3554);
and U5451 (N_5451,N_2066,N_4835);
nand U5452 (N_5452,N_108,N_2552);
nor U5453 (N_5453,N_4326,N_2398);
and U5454 (N_5454,N_3401,N_3643);
nor U5455 (N_5455,N_4248,N_613);
or U5456 (N_5456,N_4873,N_4224);
and U5457 (N_5457,N_593,N_595);
nor U5458 (N_5458,N_3603,N_444);
and U5459 (N_5459,N_2883,N_3840);
and U5460 (N_5460,N_2056,N_1057);
nand U5461 (N_5461,N_1303,N_3766);
or U5462 (N_5462,N_2679,N_4686);
nor U5463 (N_5463,N_493,N_1052);
or U5464 (N_5464,N_4811,N_2409);
and U5465 (N_5465,N_4660,N_4411);
and U5466 (N_5466,N_322,N_418);
nor U5467 (N_5467,N_3217,N_4607);
or U5468 (N_5468,N_231,N_4796);
nor U5469 (N_5469,N_4235,N_3248);
nor U5470 (N_5470,N_4309,N_482);
nand U5471 (N_5471,N_2015,N_2779);
nor U5472 (N_5472,N_2666,N_1176);
nand U5473 (N_5473,N_4349,N_167);
nor U5474 (N_5474,N_4146,N_4086);
and U5475 (N_5475,N_4279,N_1004);
nand U5476 (N_5476,N_610,N_861);
and U5477 (N_5477,N_1427,N_1334);
and U5478 (N_5478,N_2059,N_2506);
and U5479 (N_5479,N_4425,N_790);
and U5480 (N_5480,N_4456,N_632);
and U5481 (N_5481,N_2331,N_320);
or U5482 (N_5482,N_2092,N_135);
nand U5483 (N_5483,N_2967,N_773);
xor U5484 (N_5484,N_1683,N_3793);
nor U5485 (N_5485,N_1480,N_4475);
nor U5486 (N_5486,N_2280,N_3426);
and U5487 (N_5487,N_4902,N_3494);
and U5488 (N_5488,N_4390,N_402);
or U5489 (N_5489,N_612,N_2427);
nand U5490 (N_5490,N_1028,N_1136);
and U5491 (N_5491,N_3257,N_1081);
and U5492 (N_5492,N_1904,N_2693);
nand U5493 (N_5493,N_1188,N_4685);
nand U5494 (N_5494,N_984,N_3767);
or U5495 (N_5495,N_3132,N_88);
and U5496 (N_5496,N_1168,N_575);
or U5497 (N_5497,N_3408,N_3960);
xnor U5498 (N_5498,N_3644,N_1254);
nand U5499 (N_5499,N_2790,N_2351);
or U5500 (N_5500,N_812,N_4294);
nand U5501 (N_5501,N_3816,N_3042);
or U5502 (N_5502,N_3549,N_4935);
nand U5503 (N_5503,N_2522,N_2905);
nor U5504 (N_5504,N_2852,N_3485);
nand U5505 (N_5505,N_3250,N_94);
nor U5506 (N_5506,N_258,N_620);
or U5507 (N_5507,N_4208,N_2380);
or U5508 (N_5508,N_3378,N_1718);
nor U5509 (N_5509,N_1787,N_2876);
nor U5510 (N_5510,N_3278,N_3841);
or U5511 (N_5511,N_36,N_182);
nor U5512 (N_5512,N_1392,N_1954);
xor U5513 (N_5513,N_1173,N_3923);
nand U5514 (N_5514,N_1378,N_647);
nand U5515 (N_5515,N_1850,N_675);
nor U5516 (N_5516,N_2392,N_2703);
nand U5517 (N_5517,N_532,N_2130);
or U5518 (N_5518,N_1543,N_4784);
or U5519 (N_5519,N_4194,N_336);
nand U5520 (N_5520,N_2192,N_4912);
nand U5521 (N_5521,N_4810,N_4057);
or U5522 (N_5522,N_2423,N_82);
nand U5523 (N_5523,N_326,N_3183);
nand U5524 (N_5524,N_912,N_1457);
nor U5525 (N_5525,N_392,N_2081);
or U5526 (N_5526,N_1684,N_1728);
nand U5527 (N_5527,N_1583,N_4021);
or U5528 (N_5528,N_2053,N_3578);
or U5529 (N_5529,N_1952,N_3936);
nor U5530 (N_5530,N_4041,N_1371);
and U5531 (N_5531,N_2450,N_1842);
and U5532 (N_5532,N_3735,N_4609);
nand U5533 (N_5533,N_447,N_3665);
nor U5534 (N_5534,N_2498,N_4242);
nor U5535 (N_5535,N_1770,N_242);
or U5536 (N_5536,N_442,N_3255);
nand U5537 (N_5537,N_1327,N_1946);
or U5538 (N_5538,N_1030,N_635);
and U5539 (N_5539,N_4438,N_3366);
and U5540 (N_5540,N_3739,N_2882);
nor U5541 (N_5541,N_1595,N_4569);
or U5542 (N_5542,N_3592,N_4938);
and U5543 (N_5543,N_4863,N_3782);
nor U5544 (N_5544,N_2616,N_887);
and U5545 (N_5545,N_3110,N_2298);
and U5546 (N_5546,N_2757,N_4700);
or U5547 (N_5547,N_2401,N_3528);
and U5548 (N_5548,N_517,N_2723);
nand U5549 (N_5549,N_3525,N_4786);
or U5550 (N_5550,N_551,N_2019);
and U5551 (N_5551,N_3625,N_1552);
and U5552 (N_5552,N_2236,N_294);
nor U5553 (N_5553,N_3708,N_525);
or U5554 (N_5554,N_4239,N_3810);
and U5555 (N_5555,N_2648,N_1005);
nand U5556 (N_5556,N_4052,N_1355);
nor U5557 (N_5557,N_3271,N_1158);
nor U5558 (N_5558,N_1103,N_1887);
nor U5559 (N_5559,N_3503,N_557);
or U5560 (N_5560,N_2602,N_2025);
nor U5561 (N_5561,N_1845,N_331);
nand U5562 (N_5562,N_671,N_3509);
nor U5563 (N_5563,N_4763,N_4849);
nand U5564 (N_5564,N_2609,N_1763);
or U5565 (N_5565,N_2629,N_998);
nand U5566 (N_5566,N_1074,N_1338);
nand U5567 (N_5567,N_2615,N_3098);
or U5568 (N_5568,N_4244,N_1407);
or U5569 (N_5569,N_3370,N_1512);
nand U5570 (N_5570,N_2675,N_1118);
nor U5571 (N_5571,N_1615,N_3166);
or U5572 (N_5572,N_1414,N_2930);
nor U5573 (N_5573,N_3672,N_4303);
and U5574 (N_5574,N_3507,N_298);
and U5575 (N_5575,N_4613,N_1771);
nor U5576 (N_5576,N_951,N_4460);
and U5577 (N_5577,N_2229,N_4668);
or U5578 (N_5578,N_2164,N_4857);
nand U5579 (N_5579,N_625,N_2577);
or U5580 (N_5580,N_1892,N_2194);
nand U5581 (N_5581,N_805,N_2385);
or U5582 (N_5582,N_4471,N_3639);
and U5583 (N_5583,N_3851,N_4571);
and U5584 (N_5584,N_3114,N_198);
nand U5585 (N_5585,N_3225,N_3144);
and U5586 (N_5586,N_949,N_3619);
nor U5587 (N_5587,N_1806,N_1986);
nand U5588 (N_5588,N_1091,N_3929);
and U5589 (N_5589,N_3577,N_4567);
nor U5590 (N_5590,N_3301,N_4328);
or U5591 (N_5591,N_3411,N_124);
nand U5592 (N_5592,N_1105,N_3454);
and U5593 (N_5593,N_4683,N_3045);
nor U5594 (N_5594,N_3320,N_4974);
or U5595 (N_5595,N_3671,N_1347);
or U5596 (N_5596,N_4663,N_727);
nor U5597 (N_5597,N_1357,N_239);
xnor U5598 (N_5598,N_2316,N_3249);
and U5599 (N_5599,N_3989,N_1711);
or U5600 (N_5600,N_4883,N_1296);
nand U5601 (N_5601,N_3674,N_2147);
or U5602 (N_5602,N_2422,N_1333);
nor U5603 (N_5603,N_1944,N_2674);
nand U5604 (N_5604,N_498,N_489);
nor U5605 (N_5605,N_2692,N_1019);
or U5606 (N_5606,N_2562,N_2715);
nand U5607 (N_5607,N_2122,N_4557);
nor U5608 (N_5608,N_1567,N_1853);
or U5609 (N_5609,N_4549,N_338);
and U5610 (N_5610,N_3054,N_2793);
nand U5611 (N_5611,N_3328,N_4192);
xor U5612 (N_5612,N_3246,N_1661);
and U5613 (N_5613,N_2582,N_1697);
and U5614 (N_5614,N_1031,N_3067);
nor U5615 (N_5615,N_4225,N_3336);
nor U5616 (N_5616,N_150,N_2009);
nand U5617 (N_5617,N_3416,N_1948);
or U5618 (N_5618,N_2800,N_1315);
and U5619 (N_5619,N_2374,N_4953);
and U5620 (N_5620,N_399,N_2963);
nand U5621 (N_5621,N_4698,N_4675);
or U5622 (N_5622,N_3451,N_490);
nand U5623 (N_5623,N_4036,N_2372);
nand U5624 (N_5624,N_4061,N_768);
or U5625 (N_5625,N_4735,N_3992);
or U5626 (N_5626,N_1015,N_1497);
and U5627 (N_5627,N_2914,N_708);
nand U5628 (N_5628,N_832,N_720);
or U5629 (N_5629,N_4665,N_4069);
nand U5630 (N_5630,N_2443,N_4928);
nor U5631 (N_5631,N_709,N_1453);
or U5632 (N_5632,N_2983,N_4332);
nand U5633 (N_5633,N_4940,N_3039);
nor U5634 (N_5634,N_1796,N_3471);
and U5635 (N_5635,N_4864,N_2746);
or U5636 (N_5636,N_4495,N_3806);
or U5637 (N_5637,N_3897,N_1603);
or U5638 (N_5638,N_2360,N_831);
nand U5639 (N_5639,N_592,N_121);
and U5640 (N_5640,N_1939,N_1362);
or U5641 (N_5641,N_1346,N_12);
and U5642 (N_5642,N_622,N_4885);
nor U5643 (N_5643,N_2311,N_2539);
or U5644 (N_5644,N_3823,N_2831);
nand U5645 (N_5645,N_66,N_1224);
or U5646 (N_5646,N_4485,N_4905);
and U5647 (N_5647,N_1743,N_208);
nand U5648 (N_5648,N_4839,N_1859);
or U5649 (N_5649,N_2565,N_3296);
or U5650 (N_5650,N_2461,N_3082);
or U5651 (N_5651,N_2094,N_1533);
or U5652 (N_5652,N_1505,N_3065);
nor U5653 (N_5653,N_1608,N_2010);
or U5654 (N_5654,N_2564,N_585);
xnor U5655 (N_5655,N_3444,N_4408);
and U5656 (N_5656,N_560,N_273);
nor U5657 (N_5657,N_1307,N_1765);
and U5658 (N_5658,N_4032,N_4181);
nand U5659 (N_5659,N_3263,N_3831);
nand U5660 (N_5660,N_2003,N_3186);
nor U5661 (N_5661,N_247,N_2660);
and U5662 (N_5662,N_4011,N_2126);
nor U5663 (N_5663,N_4102,N_4845);
nand U5664 (N_5664,N_2297,N_3858);
or U5665 (N_5665,N_427,N_4854);
nand U5666 (N_5666,N_2949,N_2672);
nor U5667 (N_5667,N_4664,N_3473);
or U5668 (N_5668,N_55,N_4405);
nor U5669 (N_5669,N_1647,N_4993);
nor U5670 (N_5670,N_13,N_4391);
and U5671 (N_5671,N_205,N_817);
xor U5672 (N_5672,N_1192,N_1035);
or U5673 (N_5673,N_1242,N_4101);
nand U5674 (N_5674,N_3259,N_2127);
nand U5675 (N_5675,N_3581,N_995);
nand U5676 (N_5676,N_1799,N_4071);
nand U5677 (N_5677,N_3177,N_2570);
or U5678 (N_5678,N_2458,N_581);
or U5679 (N_5679,N_3369,N_1818);
and U5680 (N_5680,N_3707,N_1481);
nand U5681 (N_5681,N_2559,N_1258);
or U5682 (N_5682,N_1660,N_4222);
nor U5683 (N_5683,N_2600,N_3305);
nor U5684 (N_5684,N_1092,N_3037);
nor U5685 (N_5685,N_603,N_4770);
nor U5686 (N_5686,N_854,N_4398);
or U5687 (N_5687,N_1717,N_3570);
nor U5688 (N_5688,N_828,N_4443);
nand U5689 (N_5689,N_4590,N_2008);
nor U5690 (N_5690,N_3898,N_867);
nand U5691 (N_5691,N_3206,N_319);
nand U5692 (N_5692,N_200,N_3829);
or U5693 (N_5693,N_865,N_4798);
nand U5694 (N_5694,N_3231,N_4751);
nand U5695 (N_5695,N_1521,N_4805);
and U5696 (N_5696,N_619,N_4431);
xnor U5697 (N_5697,N_3628,N_3894);
nand U5698 (N_5698,N_3015,N_2467);
and U5699 (N_5699,N_521,N_4467);
nor U5700 (N_5700,N_274,N_2284);
or U5701 (N_5701,N_2505,N_638);
nor U5702 (N_5702,N_1596,N_3440);
nand U5703 (N_5703,N_1026,N_1373);
and U5704 (N_5704,N_3595,N_372);
nor U5705 (N_5705,N_4829,N_1879);
nor U5706 (N_5706,N_2634,N_1726);
nand U5707 (N_5707,N_4642,N_607);
and U5708 (N_5708,N_1379,N_1356);
or U5709 (N_5709,N_3254,N_1844);
nor U5710 (N_5710,N_3681,N_2798);
nor U5711 (N_5711,N_2478,N_3849);
nor U5712 (N_5712,N_4982,N_1498);
or U5713 (N_5713,N_437,N_4022);
nand U5714 (N_5714,N_310,N_3826);
or U5715 (N_5715,N_3497,N_3321);
and U5716 (N_5716,N_4213,N_3496);
nand U5717 (N_5717,N_1712,N_2778);
or U5718 (N_5718,N_3997,N_3151);
or U5719 (N_5719,N_1375,N_2927);
nand U5720 (N_5720,N_113,N_2174);
or U5721 (N_5721,N_351,N_2628);
and U5722 (N_5722,N_4272,N_3293);
or U5723 (N_5723,N_1651,N_1257);
nor U5724 (N_5724,N_2737,N_3003);
or U5725 (N_5725,N_3637,N_419);
or U5726 (N_5726,N_501,N_558);
xnor U5727 (N_5727,N_3572,N_553);
or U5728 (N_5728,N_4559,N_2370);
nand U5729 (N_5729,N_2680,N_428);
nor U5730 (N_5730,N_241,N_1686);
xnor U5731 (N_5731,N_640,N_213);
or U5732 (N_5732,N_1349,N_2851);
and U5733 (N_5733,N_3030,N_4954);
nor U5734 (N_5734,N_227,N_3645);
nor U5735 (N_5735,N_3756,N_3984);
or U5736 (N_5736,N_1329,N_1458);
nor U5737 (N_5737,N_4418,N_3781);
nand U5738 (N_5738,N_3908,N_3977);
nand U5739 (N_5739,N_3618,N_95);
and U5740 (N_5740,N_1814,N_2165);
nand U5741 (N_5741,N_2486,N_3565);
and U5742 (N_5742,N_2470,N_1260);
or U5743 (N_5743,N_1504,N_3657);
xor U5744 (N_5744,N_2397,N_1696);
nor U5745 (N_5745,N_1703,N_3724);
nand U5746 (N_5746,N_1096,N_2772);
or U5747 (N_5747,N_1395,N_275);
and U5748 (N_5748,N_118,N_2750);
and U5749 (N_5749,N_3523,N_3314);
nor U5750 (N_5750,N_397,N_4757);
or U5751 (N_5751,N_3063,N_577);
nand U5752 (N_5752,N_3993,N_2589);
nor U5753 (N_5753,N_1511,N_1389);
nor U5754 (N_5754,N_2610,N_2741);
or U5755 (N_5755,N_3617,N_2781);
nor U5756 (N_5756,N_3635,N_211);
and U5757 (N_5757,N_2488,N_1862);
and U5758 (N_5758,N_2054,N_833);
nor U5759 (N_5759,N_4732,N_4134);
or U5760 (N_5760,N_1628,N_2632);
nand U5761 (N_5761,N_3425,N_1838);
nand U5762 (N_5762,N_1072,N_2753);
nor U5763 (N_5763,N_4690,N_4767);
or U5764 (N_5764,N_2705,N_2525);
nand U5765 (N_5765,N_4221,N_4793);
nor U5766 (N_5766,N_2592,N_1310);
and U5767 (N_5767,N_3475,N_1069);
or U5768 (N_5768,N_2022,N_1048);
or U5769 (N_5769,N_3976,N_4872);
or U5770 (N_5770,N_1965,N_3060);
or U5771 (N_5771,N_3190,N_3627);
nand U5772 (N_5772,N_2644,N_2535);
or U5773 (N_5773,N_2318,N_4831);
or U5774 (N_5774,N_1835,N_3472);
or U5775 (N_5775,N_3538,N_4109);
or U5776 (N_5776,N_4317,N_2224);
nand U5777 (N_5777,N_3267,N_2274);
nand U5778 (N_5778,N_2038,N_3235);
nand U5779 (N_5779,N_4338,N_4442);
nand U5780 (N_5780,N_4476,N_1788);
or U5781 (N_5781,N_4010,N_4672);
or U5782 (N_5782,N_3983,N_3847);
and U5783 (N_5783,N_1146,N_512);
nand U5784 (N_5784,N_2244,N_844);
or U5785 (N_5785,N_1121,N_1592);
or U5786 (N_5786,N_803,N_2294);
or U5787 (N_5787,N_1698,N_4127);
nand U5788 (N_5788,N_4907,N_3506);
nand U5789 (N_5789,N_4126,N_400);
nand U5790 (N_5790,N_303,N_282);
or U5791 (N_5791,N_4647,N_141);
or U5792 (N_5792,N_2205,N_4363);
nor U5793 (N_5793,N_54,N_3287);
nor U5794 (N_5794,N_4014,N_4920);
and U5795 (N_5795,N_279,N_3785);
nor U5796 (N_5796,N_3952,N_4105);
nor U5797 (N_5797,N_1359,N_3758);
and U5798 (N_5798,N_3704,N_4392);
or U5799 (N_5799,N_798,N_4738);
nand U5800 (N_5800,N_1169,N_3050);
and U5801 (N_5801,N_4116,N_229);
nand U5802 (N_5802,N_4599,N_4429);
nand U5803 (N_5803,N_3876,N_3159);
or U5804 (N_5804,N_348,N_4503);
nand U5805 (N_5805,N_1558,N_2439);
nor U5806 (N_5806,N_4428,N_2994);
nand U5807 (N_5807,N_2649,N_3787);
nand U5808 (N_5808,N_1399,N_4468);
nand U5809 (N_5809,N_1995,N_329);
or U5810 (N_5810,N_4787,N_3214);
and U5811 (N_5811,N_1694,N_3903);
nor U5812 (N_5812,N_2731,N_475);
nand U5813 (N_5813,N_3139,N_391);
nor U5814 (N_5814,N_1547,N_2934);
xor U5815 (N_5815,N_206,N_3842);
or U5816 (N_5816,N_1682,N_4043);
nor U5817 (N_5817,N_819,N_4068);
and U5818 (N_5818,N_1826,N_1520);
nand U5819 (N_5819,N_441,N_3624);
nor U5820 (N_5820,N_1222,N_207);
nand U5821 (N_5821,N_4492,N_3926);
nand U5822 (N_5822,N_467,N_2959);
nor U5823 (N_5823,N_28,N_1964);
nand U5824 (N_5824,N_2144,N_149);
nor U5825 (N_5825,N_4843,N_4044);
or U5826 (N_5826,N_3431,N_1473);
nand U5827 (N_5827,N_2247,N_3256);
and U5828 (N_5828,N_1680,N_4500);
or U5829 (N_5829,N_1109,N_173);
nand U5830 (N_5830,N_3878,N_245);
nor U5831 (N_5831,N_2921,N_2940);
or U5832 (N_5832,N_1488,N_3405);
xor U5833 (N_5833,N_1131,N_1670);
or U5834 (N_5834,N_248,N_4550);
and U5835 (N_5835,N_4802,N_4096);
nand U5836 (N_5836,N_1798,N_3804);
or U5837 (N_5837,N_3714,N_3653);
nor U5838 (N_5838,N_4533,N_2681);
and U5839 (N_5839,N_4858,N_2399);
nand U5840 (N_5840,N_4889,N_3631);
nor U5841 (N_5841,N_3962,N_4646);
nor U5842 (N_5842,N_3004,N_1565);
and U5843 (N_5843,N_4358,N_545);
nor U5844 (N_5844,N_4291,N_4552);
nand U5845 (N_5845,N_4856,N_890);
nor U5846 (N_5846,N_2804,N_2654);
or U5847 (N_5847,N_986,N_3560);
or U5848 (N_5848,N_4929,N_4416);
and U5849 (N_5849,N_657,N_2260);
nand U5850 (N_5850,N_3942,N_3412);
nand U5851 (N_5851,N_4384,N_2006);
or U5852 (N_5852,N_219,N_7);
and U5853 (N_5853,N_536,N_4342);
or U5854 (N_5854,N_1085,N_3286);
or U5855 (N_5855,N_4006,N_3359);
or U5856 (N_5856,N_1619,N_856);
nor U5857 (N_5857,N_3134,N_2074);
nor U5858 (N_5858,N_4977,N_2785);
and U5859 (N_5859,N_4545,N_4565);
nor U5860 (N_5860,N_235,N_3698);
nand U5861 (N_5861,N_3360,N_4876);
nor U5862 (N_5862,N_383,N_659);
nand U5863 (N_5863,N_2642,N_3322);
nand U5864 (N_5864,N_893,N_1452);
nor U5865 (N_5865,N_4491,N_4274);
nor U5866 (N_5866,N_1022,N_3228);
nor U5867 (N_5867,N_4336,N_4713);
and U5868 (N_5868,N_533,N_1525);
nor U5869 (N_5869,N_2797,N_67);
nor U5870 (N_5870,N_3813,N_518);
nor U5871 (N_5871,N_3489,N_2749);
nor U5872 (N_5872,N_3309,N_1913);
and U5873 (N_5873,N_3808,N_2611);
or U5874 (N_5874,N_2877,N_4961);
nor U5875 (N_5875,N_2742,N_3453);
nor U5876 (N_5876,N_1779,N_1125);
nand U5877 (N_5877,N_2282,N_3119);
nand U5878 (N_5878,N_2902,N_1625);
nor U5879 (N_5879,N_4553,N_752);
and U5880 (N_5880,N_1575,N_4238);
and U5881 (N_5881,N_3227,N_3728);
nand U5882 (N_5882,N_86,N_3495);
nand U5883 (N_5883,N_1063,N_1336);
and U5884 (N_5884,N_1038,N_3338);
and U5885 (N_5885,N_4959,N_2103);
or U5886 (N_5886,N_478,N_1313);
xnor U5887 (N_5887,N_2962,N_3071);
nand U5888 (N_5888,N_128,N_1133);
nand U5889 (N_5889,N_2894,N_78);
nand U5890 (N_5890,N_3118,N_3055);
nand U5891 (N_5891,N_2036,N_2463);
or U5892 (N_5892,N_1710,N_1144);
and U5893 (N_5893,N_76,N_163);
nor U5894 (N_5894,N_4602,N_2253);
nand U5895 (N_5895,N_4110,N_730);
nand U5896 (N_5896,N_1700,N_4689);
or U5897 (N_5897,N_2773,N_3356);
nand U5898 (N_5898,N_1557,N_2585);
nand U5899 (N_5899,N_2756,N_4025);
nor U5900 (N_5900,N_1820,N_1009);
nand U5901 (N_5901,N_2892,N_423);
or U5902 (N_5902,N_1201,N_4600);
nand U5903 (N_5903,N_3701,N_3348);
or U5904 (N_5904,N_930,N_2387);
nand U5905 (N_5905,N_3283,N_3946);
and U5906 (N_5906,N_2460,N_4975);
nor U5907 (N_5907,N_1465,N_462);
and U5908 (N_5908,N_1108,N_3607);
nor U5909 (N_5909,N_1129,N_3291);
nor U5910 (N_5910,N_3064,N_115);
nor U5911 (N_5911,N_1865,N_4304);
or U5912 (N_5912,N_4278,N_2704);
nor U5913 (N_5913,N_2004,N_3988);
and U5914 (N_5914,N_3530,N_340);
or U5915 (N_5915,N_2647,N_3948);
or U5916 (N_5916,N_2613,N_4201);
or U5917 (N_5917,N_3737,N_928);
nand U5918 (N_5918,N_246,N_2606);
nand U5919 (N_5919,N_3824,N_2575);
xor U5920 (N_5920,N_2554,N_4794);
or U5921 (N_5921,N_2578,N_374);
nor U5922 (N_5922,N_1054,N_1636);
and U5923 (N_5923,N_215,N_3029);
or U5924 (N_5924,N_2903,N_1848);
nand U5925 (N_5925,N_4427,N_3856);
nand U5926 (N_5926,N_3072,N_484);
nor U5927 (N_5927,N_2515,N_2135);
or U5928 (N_5928,N_1,N_693);
and U5929 (N_5929,N_4637,N_1977);
nand U5930 (N_5930,N_4315,N_2946);
or U5931 (N_5931,N_2250,N_1097);
nand U5932 (N_5932,N_3995,N_1194);
nand U5933 (N_5933,N_1484,N_2285);
and U5934 (N_5934,N_2075,N_2860);
and U5935 (N_5935,N_4270,N_4608);
nor U5936 (N_5936,N_3130,N_1196);
nor U5937 (N_5937,N_1180,N_1704);
and U5938 (N_5938,N_4063,N_2817);
nor U5939 (N_5939,N_960,N_2393);
nor U5940 (N_5940,N_2425,N_2712);
nand U5941 (N_5941,N_299,N_2061);
nor U5942 (N_5942,N_862,N_4531);
nor U5943 (N_5943,N_3594,N_157);
nand U5944 (N_5944,N_4687,N_4202);
and U5945 (N_5945,N_4834,N_2330);
nand U5946 (N_5946,N_4814,N_1899);
nor U5947 (N_5947,N_4163,N_2830);
nor U5948 (N_5948,N_1175,N_1002);
nand U5949 (N_5949,N_590,N_2764);
or U5950 (N_5950,N_4087,N_1386);
nor U5951 (N_5951,N_4054,N_3696);
or U5952 (N_5952,N_3532,N_3580);
nor U5953 (N_5953,N_2404,N_4830);
or U5954 (N_5954,N_3415,N_1871);
nor U5955 (N_5955,N_2657,N_31);
nor U5956 (N_5956,N_424,N_102);
and U5957 (N_5957,N_4280,N_908);
or U5958 (N_5958,N_3332,N_1437);
nand U5959 (N_5959,N_2496,N_1556);
xor U5960 (N_5960,N_4030,N_2223);
or U5961 (N_5961,N_3500,N_1634);
and U5962 (N_5962,N_4186,N_4155);
nand U5963 (N_5963,N_1029,N_1723);
or U5964 (N_5964,N_1819,N_3070);
nor U5965 (N_5965,N_3455,N_4926);
nand U5966 (N_5966,N_677,N_1482);
xor U5967 (N_5967,N_2150,N_716);
nand U5968 (N_5968,N_3797,N_2663);
nand U5969 (N_5969,N_2225,N_2251);
or U5970 (N_5970,N_2698,N_1447);
and U5971 (N_5971,N_1679,N_2276);
nor U5972 (N_5972,N_1493,N_4893);
and U5973 (N_5973,N_2926,N_1532);
or U5974 (N_5974,N_2920,N_1376);
nand U5975 (N_5975,N_201,N_2079);
nor U5976 (N_5976,N_3769,N_767);
nor U5977 (N_5977,N_56,N_684);
nor U5978 (N_5978,N_4908,N_2031);
and U5979 (N_5979,N_4409,N_233);
nand U5980 (N_5980,N_4847,N_996);
or U5981 (N_5981,N_1905,N_2241);
or U5982 (N_5982,N_3562,N_3967);
nand U5983 (N_5983,N_3172,N_742);
nor U5984 (N_5984,N_4394,N_2279);
nand U5985 (N_5985,N_725,N_2803);
nor U5986 (N_5986,N_3160,N_2109);
or U5987 (N_5987,N_3417,N_197);
and U5988 (N_5988,N_4502,N_3410);
nand U5989 (N_5989,N_898,N_3512);
and U5990 (N_5990,N_2072,N_4215);
nor U5991 (N_5991,N_2159,N_2809);
or U5992 (N_5992,N_3656,N_707);
nand U5993 (N_5993,N_311,N_45);
or U5994 (N_5994,N_988,N_1195);
and U5995 (N_5995,N_4190,N_1701);
and U5996 (N_5996,N_608,N_4837);
and U5997 (N_5997,N_4874,N_1514);
nand U5998 (N_5998,N_3930,N_2482);
and U5999 (N_5999,N_1156,N_4046);
and U6000 (N_6000,N_845,N_2933);
nand U6001 (N_6001,N_2076,N_3317);
nor U6002 (N_6002,N_295,N_330);
and U6003 (N_6003,N_4532,N_4543);
nor U6004 (N_6004,N_89,N_1657);
or U6005 (N_6005,N_2826,N_1955);
or U6006 (N_6006,N_366,N_4937);
nor U6007 (N_6007,N_1923,N_346);
nor U6008 (N_6008,N_1849,N_1813);
nand U6009 (N_6009,N_1365,N_4103);
and U6010 (N_6010,N_3513,N_3860);
nand U6011 (N_6011,N_3437,N_2874);
or U6012 (N_6012,N_3526,N_4879);
and U6013 (N_6013,N_57,N_3688);
and U6014 (N_6014,N_4175,N_1681);
nor U6015 (N_6015,N_3198,N_3620);
nand U6016 (N_6016,N_3650,N_2089);
nand U6017 (N_6017,N_2771,N_2293);
nor U6018 (N_6018,N_2594,N_2743);
nand U6019 (N_6019,N_4501,N_492);
nor U6020 (N_6020,N_1191,N_692);
nor U6021 (N_6021,N_2591,N_4034);
and U6022 (N_6022,N_2388,N_2821);
and U6023 (N_6023,N_2021,N_477);
and U6024 (N_6024,N_1059,N_1825);
nor U6025 (N_6025,N_1739,N_196);
and U6026 (N_6026,N_2965,N_2491);
and U6027 (N_6027,N_2720,N_4355);
nor U6028 (N_6028,N_766,N_3741);
nor U6029 (N_6029,N_631,N_688);
or U6030 (N_6030,N_3873,N_2956);
and U6031 (N_6031,N_2420,N_749);
nand U6032 (N_6032,N_3280,N_1523);
or U6033 (N_6033,N_3367,N_431);
nand U6034 (N_6034,N_4372,N_3917);
and U6035 (N_6035,N_1733,N_1478);
nor U6036 (N_6036,N_2581,N_1412);
nor U6037 (N_6037,N_1793,N_4706);
nor U6038 (N_6038,N_2651,N_4351);
and U6039 (N_6039,N_3241,N_4871);
and U6040 (N_6040,N_4334,N_3421);
and U6041 (N_6041,N_2907,N_4490);
nand U6042 (N_6042,N_2829,N_534);
and U6043 (N_6043,N_3468,N_3362);
and U6044 (N_6044,N_4806,N_4645);
and U6045 (N_6045,N_4125,N_4120);
nand U6046 (N_6046,N_379,N_2477);
nand U6047 (N_6047,N_1810,N_3761);
and U6048 (N_6048,N_4862,N_2290);
nor U6049 (N_6049,N_1546,N_835);
and U6050 (N_6050,N_1055,N_1297);
nand U6051 (N_6051,N_3866,N_2784);
nand U6052 (N_6052,N_4914,N_3541);
nand U6053 (N_6053,N_252,N_4894);
nor U6054 (N_6054,N_1394,N_249);
or U6055 (N_6055,N_3550,N_3601);
nor U6056 (N_6056,N_939,N_4804);
nand U6057 (N_6057,N_2455,N_3602);
nand U6058 (N_6058,N_4995,N_3097);
or U6059 (N_6059,N_2527,N_3043);
nand U6060 (N_6060,N_91,N_3973);
or U6061 (N_6061,N_4481,N_410);
or U6062 (N_6062,N_4616,N_3777);
nand U6063 (N_6063,N_1071,N_3389);
xor U6064 (N_6064,N_4142,N_4867);
nor U6065 (N_6065,N_4448,N_3161);
and U6066 (N_6066,N_1160,N_2101);
nor U6067 (N_6067,N_1752,N_4343);
nor U6068 (N_6068,N_71,N_3686);
nand U6069 (N_6069,N_1689,N_2566);
nor U6070 (N_6070,N_3715,N_2248);
or U6071 (N_6071,N_2500,N_1110);
or U6072 (N_6072,N_3900,N_250);
and U6073 (N_6073,N_2630,N_1142);
and U6074 (N_6074,N_2810,N_2501);
nor U6075 (N_6075,N_2856,N_183);
nor U6076 (N_6076,N_4306,N_3764);
nand U6077 (N_6077,N_187,N_4119);
and U6078 (N_6078,N_342,N_3006);
and U6079 (N_6079,N_2173,N_2843);
nand U6080 (N_6080,N_3702,N_2695);
or U6081 (N_6081,N_1490,N_2105);
and U6082 (N_6082,N_4017,N_615);
nor U6083 (N_6083,N_851,N_4412);
and U6084 (N_6084,N_700,N_4725);
nor U6085 (N_6085,N_1829,N_703);
or U6086 (N_6086,N_4027,N_3040);
nor U6087 (N_6087,N_2067,N_3563);
nor U6088 (N_6088,N_1866,N_3335);
nor U6089 (N_6089,N_1135,N_4081);
and U6090 (N_6090,N_3087,N_3519);
and U6091 (N_6091,N_223,N_4160);
or U6092 (N_6092,N_2765,N_80);
and U6093 (N_6093,N_2413,N_3803);
or U6094 (N_6094,N_1576,N_1446);
xnor U6095 (N_6095,N_2217,N_2837);
and U6096 (N_6096,N_1564,N_713);
nand U6097 (N_6097,N_2745,N_3593);
and U6098 (N_6098,N_4903,N_1309);
nand U6099 (N_6099,N_1126,N_3422);
or U6100 (N_6100,N_1263,N_3116);
or U6101 (N_6101,N_4691,N_2209);
nand U6102 (N_6102,N_4104,N_2475);
and U6103 (N_6103,N_4624,N_4538);
nor U6104 (N_6104,N_967,N_2541);
nor U6105 (N_6105,N_2936,N_3621);
and U6106 (N_6106,N_694,N_3770);
nand U6107 (N_6107,N_1841,N_3815);
nor U6108 (N_6108,N_1502,N_3459);
or U6109 (N_6109,N_1354,N_702);
or U6110 (N_6110,N_4433,N_1883);
or U6111 (N_6111,N_2492,N_3655);
and U6112 (N_6112,N_293,N_1695);
and U6113 (N_6113,N_1425,N_3428);
or U6114 (N_6114,N_3282,N_1368);
or U6115 (N_6115,N_1645,N_868);
and U6116 (N_6116,N_1051,N_4528);
and U6117 (N_6117,N_2603,N_3018);
and U6118 (N_6118,N_2494,N_528);
nor U6119 (N_6119,N_64,N_2292);
and U6120 (N_6120,N_2662,N_2947);
nand U6121 (N_6121,N_412,N_4990);
or U6122 (N_6122,N_3313,N_4563);
and U6123 (N_6123,N_2314,N_1920);
nand U6124 (N_6124,N_4183,N_1245);
or U6125 (N_6125,N_1039,N_3906);
or U6126 (N_6126,N_1398,N_2834);
and U6127 (N_6127,N_1872,N_2411);
or U6128 (N_6128,N_4039,N_2268);
nand U6129 (N_6129,N_292,N_2115);
and U6130 (N_6130,N_4200,N_2621);
or U6131 (N_6131,N_269,N_4413);
nand U6132 (N_6132,N_1145,N_1756);
nor U6133 (N_6133,N_503,N_2924);
nor U6134 (N_6134,N_3375,N_4273);
and U6135 (N_6135,N_1304,N_3152);
or U6136 (N_6136,N_4422,N_1803);
or U6137 (N_6137,N_2943,N_4816);
nor U6138 (N_6138,N_747,N_3795);
and U6139 (N_6139,N_1981,N_959);
or U6140 (N_6140,N_1077,N_4618);
nand U6141 (N_6141,N_4936,N_160);
or U6142 (N_6142,N_1238,N_3706);
nor U6143 (N_6143,N_2362,N_586);
nor U6144 (N_6144,N_1693,N_1226);
or U6145 (N_6145,N_955,N_2839);
nand U6146 (N_6146,N_1288,N_3662);
nor U6147 (N_6147,N_3020,N_4688);
nand U6148 (N_6148,N_202,N_4499);
and U6149 (N_6149,N_2676,N_4658);
and U6150 (N_6150,N_1324,N_146);
nand U6151 (N_6151,N_864,N_3974);
nand U6152 (N_6152,N_217,N_3693);
and U6153 (N_6153,N_1921,N_3896);
and U6154 (N_6154,N_185,N_2599);
and U6155 (N_6155,N_4709,N_3867);
nand U6156 (N_6156,N_4962,N_2931);
nor U6157 (N_6157,N_3073,N_1790);
nor U6158 (N_6158,N_4231,N_2044);
or U6159 (N_6159,N_2656,N_1262);
or U6160 (N_6160,N_1994,N_3508);
and U6161 (N_6161,N_2706,N_3270);
or U6162 (N_6162,N_4799,N_1746);
and U6163 (N_6163,N_2050,N_460);
nand U6164 (N_6164,N_2155,N_1758);
or U6165 (N_6165,N_823,N_2780);
nand U6166 (N_6166,N_3157,N_2977);
nor U6167 (N_6167,N_642,N_1585);
or U6168 (N_6168,N_4076,N_3207);
nor U6169 (N_6169,N_910,N_4007);
nor U6170 (N_6170,N_1409,N_4493);
nor U6171 (N_6171,N_158,N_4762);
or U6172 (N_6172,N_3584,N_4716);
nor U6173 (N_6173,N_1663,N_743);
or U6174 (N_6174,N_779,N_152);
nand U6175 (N_6175,N_1653,N_2041);
or U6176 (N_6176,N_3210,N_4313);
nor U6177 (N_6177,N_3351,N_4827);
nand U6178 (N_6178,N_4310,N_3608);
nor U6179 (N_6179,N_2689,N_2270);
and U6180 (N_6180,N_4099,N_2551);
nand U6181 (N_6181,N_3933,N_729);
or U6182 (N_6182,N_4234,N_1580);
nor U6183 (N_6183,N_4166,N_1629);
and U6184 (N_6184,N_1598,N_3275);
and U6185 (N_6185,N_4619,N_3888);
nor U6186 (N_6186,N_3164,N_3450);
and U6187 (N_6187,N_232,N_2775);
nor U6188 (N_6188,N_1007,N_1305);
or U6189 (N_6189,N_1579,N_1839);
nor U6190 (N_6190,N_451,N_3964);
nand U6191 (N_6191,N_3133,N_611);
or U6192 (N_6192,N_994,N_1901);
nand U6193 (N_6193,N_4956,N_4247);
nor U6194 (N_6194,N_178,N_765);
nor U6195 (N_6195,N_4774,N_27);
nor U6196 (N_6196,N_3862,N_1140);
and U6197 (N_6197,N_2928,N_3403);
or U6198 (N_6198,N_4591,N_4275);
nor U6199 (N_6199,N_676,N_1817);
and U6200 (N_6200,N_589,N_4100);
or U6201 (N_6201,N_3670,N_2863);
and U6202 (N_6202,N_4610,N_1269);
nor U6203 (N_6203,N_1601,N_952);
or U6204 (N_6204,N_3891,N_1203);
nor U6205 (N_6205,N_2945,N_3869);
and U6206 (N_6206,N_559,N_2673);
and U6207 (N_6207,N_3982,N_605);
nand U6208 (N_6208,N_4882,N_1017);
or U6209 (N_6209,N_332,N_2557);
nor U6210 (N_6210,N_2595,N_4356);
and U6211 (N_6211,N_3791,N_2769);
nor U6212 (N_6212,N_3487,N_1824);
and U6213 (N_6213,N_1617,N_3357);
nand U6214 (N_6214,N_1562,N_504);
and U6215 (N_6215,N_4955,N_4404);
and U6216 (N_6216,N_1040,N_1186);
nand U6217 (N_6217,N_3482,N_24);
nand U6218 (N_6218,N_2614,N_4614);
nand U6219 (N_6219,N_21,N_3733);
nor U6220 (N_6220,N_4699,N_1078);
and U6221 (N_6221,N_860,N_3717);
or U6222 (N_6222,N_3660,N_3022);
nor U6223 (N_6223,N_4345,N_2483);
nand U6224 (N_6224,N_843,N_1228);
nand U6225 (N_6225,N_4846,N_2000);
or U6226 (N_6226,N_852,N_2312);
or U6227 (N_6227,N_1605,N_2007);
nor U6228 (N_6228,N_216,N_3158);
or U6229 (N_6229,N_906,N_2528);
and U6230 (N_6230,N_2845,N_3668);
or U6231 (N_6231,N_1837,N_409);
nor U6232 (N_6232,N_2060,N_2373);
nand U6233 (N_6233,N_2289,N_2473);
or U6234 (N_6234,N_1064,N_3811);
nand U6235 (N_6235,N_4311,N_4331);
nor U6236 (N_6236,N_486,N_4154);
or U6237 (N_6237,N_4753,N_927);
nor U6238 (N_6238,N_1864,N_355);
or U6239 (N_6239,N_281,N_3736);
nor U6240 (N_6240,N_2197,N_1656);
or U6241 (N_6241,N_658,N_896);
or U6242 (N_6242,N_4065,N_4047);
or U6243 (N_6243,N_4136,N_1748);
nor U6244 (N_6244,N_2188,N_4151);
or U6245 (N_6245,N_46,N_4797);
and U6246 (N_6246,N_885,N_1317);
nand U6247 (N_6247,N_144,N_4145);
nor U6248 (N_6248,N_4506,N_3377);
nand U6249 (N_6249,N_1181,N_4462);
nor U6250 (N_6250,N_3187,N_3792);
nand U6251 (N_6251,N_2572,N_4778);
or U6252 (N_6252,N_4187,N_2421);
and U6253 (N_6253,N_669,N_2518);
or U6254 (N_6254,N_426,N_2026);
and U6255 (N_6255,N_25,N_4741);
nor U6256 (N_6256,N_1643,N_1470);
or U6257 (N_6257,N_495,N_2303);
nand U6258 (N_6258,N_4479,N_1027);
nand U6259 (N_6259,N_1933,N_1282);
nand U6260 (N_6260,N_894,N_4875);
nor U6261 (N_6261,N_948,N_4766);
nand U6262 (N_6262,N_4035,N_461);
or U6263 (N_6263,N_357,N_2027);
nand U6264 (N_6264,N_1747,N_2187);
nand U6265 (N_6265,N_875,N_1970);
or U6266 (N_6266,N_3163,N_760);
and U6267 (N_6267,N_1088,N_1508);
xnor U6268 (N_6268,N_4393,N_2255);
or U6269 (N_6269,N_880,N_3096);
nor U6270 (N_6270,N_2576,N_1554);
nor U6271 (N_6271,N_2612,N_2309);
nand U6272 (N_6272,N_3689,N_1815);
nor U6273 (N_6273,N_2152,N_4915);
nand U6274 (N_6274,N_1086,N_1794);
nor U6275 (N_6275,N_734,N_2507);
nand U6276 (N_6276,N_846,N_2131);
and U6277 (N_6277,N_3354,N_2272);
nand U6278 (N_6278,N_2207,N_2917);
and U6279 (N_6279,N_3537,N_4423);
nand U6280 (N_6280,N_4400,N_65);
or U6281 (N_6281,N_2302,N_429);
and U6282 (N_6282,N_3879,N_3379);
or U6283 (N_6283,N_1252,N_2357);
nor U6284 (N_6284,N_4388,N_1163);
nand U6285 (N_6285,N_4170,N_84);
and U6286 (N_6286,N_963,N_3889);
and U6287 (N_6287,N_4964,N_3209);
nor U6288 (N_6288,N_4410,N_3120);
or U6289 (N_6289,N_2447,N_79);
nand U6290 (N_6290,N_1566,N_1439);
and U6291 (N_6291,N_809,N_1117);
nor U6292 (N_6292,N_1534,N_1500);
and U6293 (N_6293,N_413,N_1724);
nand U6294 (N_6294,N_2958,N_224);
nand U6295 (N_6295,N_337,N_2454);
nand U6296 (N_6296,N_1384,N_145);
xor U6297 (N_6297,N_1982,N_3870);
and U6298 (N_6298,N_1483,N_1330);
nand U6299 (N_6299,N_2708,N_4895);
and U6300 (N_6300,N_3848,N_791);
nor U6301 (N_6301,N_732,N_1886);
or U6302 (N_6302,N_1062,N_4403);
nor U6303 (N_6303,N_3290,N_587);
or U6304 (N_6304,N_636,N_4984);
or U6305 (N_6305,N_4,N_4734);
nand U6306 (N_6306,N_3001,N_2317);
nand U6307 (N_6307,N_4466,N_4615);
and U6308 (N_6308,N_552,N_1801);
nand U6309 (N_6309,N_2670,N_530);
and U6310 (N_6310,N_3199,N_2341);
nand U6311 (N_6311,N_3755,N_1178);
nor U6312 (N_6312,N_199,N_1042);
nand U6313 (N_6313,N_3344,N_3329);
and U6314 (N_6314,N_3002,N_4900);
and U6315 (N_6315,N_3385,N_3125);
and U6316 (N_6316,N_502,N_3980);
or U6317 (N_6317,N_1415,N_3047);
and U6318 (N_6318,N_1878,N_4259);
nor U6319 (N_6319,N_2162,N_433);
and U6320 (N_6320,N_2213,N_3258);
nor U6321 (N_6321,N_4298,N_2369);
or U6322 (N_6322,N_2428,N_2906);
nand U6323 (N_6323,N_1301,N_4026);
nor U6324 (N_6324,N_296,N_2825);
and U6325 (N_6325,N_4265,N_2807);
nor U6326 (N_6326,N_4432,N_4078);
or U6327 (N_6327,N_971,N_436);
nor U6328 (N_6328,N_626,N_3299);
or U6329 (N_6329,N_107,N_4603);
nand U6330 (N_6330,N_1894,N_2858);
nand U6331 (N_6331,N_4164,N_3759);
and U6332 (N_6332,N_1518,N_1227);
nand U6333 (N_6333,N_2683,N_60);
and U6334 (N_6334,N_3464,N_4139);
or U6335 (N_6335,N_4681,N_4507);
nor U6336 (N_6336,N_3934,N_4922);
or U6337 (N_6337,N_129,N_3153);
and U6338 (N_6338,N_3893,N_3885);
nor U6339 (N_6339,N_668,N_3136);
nand U6340 (N_6340,N_4219,N_656);
and U6341 (N_6341,N_1809,N_4760);
and U6342 (N_6342,N_2182,N_1165);
and U6343 (N_6343,N_4153,N_934);
nor U6344 (N_6344,N_726,N_3242);
xor U6345 (N_6345,N_4361,N_401);
and U6346 (N_6346,N_3516,N_2794);
and U6347 (N_6347,N_1290,N_2495);
nor U6348 (N_6348,N_2446,N_3998);
nand U6349 (N_6349,N_770,N_2786);
nand U6350 (N_6350,N_4661,N_2713);
or U6351 (N_6351,N_1003,N_900);
and U6352 (N_6352,N_3195,N_1116);
nor U6353 (N_6353,N_2376,N_3084);
and U6354 (N_6354,N_3677,N_3573);
nand U6355 (N_6355,N_4768,N_2499);
nand U6356 (N_6356,N_2584,N_4970);
or U6357 (N_6357,N_4385,N_2818);
nor U6358 (N_6358,N_1735,N_1764);
or U6359 (N_6359,N_18,N_3556);
nor U6360 (N_6360,N_3053,N_162);
nor U6361 (N_6361,N_629,N_2567);
and U6362 (N_6362,N_2479,N_3371);
and U6363 (N_6363,N_302,N_1914);
or U6364 (N_6364,N_2365,N_1607);
and U6365 (N_6365,N_2300,N_2978);
nor U6366 (N_6366,N_2795,N_2364);
and U6367 (N_6367,N_4285,N_2598);
and U6368 (N_6368,N_3606,N_2925);
and U6369 (N_6369,N_4594,N_4540);
nand U6370 (N_6370,N_2240,N_769);
and U6371 (N_6371,N_3877,N_4707);
nor U6372 (N_6372,N_977,N_4019);
nor U6373 (N_6373,N_2234,N_3875);
or U6374 (N_6374,N_2204,N_2161);
or U6375 (N_6375,N_494,N_772);
nand U6376 (N_6376,N_1240,N_390);
and U6377 (N_6377,N_976,N_4299);
and U6378 (N_6378,N_3747,N_2744);
nor U6379 (N_6379,N_4508,N_2685);
nor U6380 (N_6380,N_1127,N_4611);
and U6381 (N_6381,N_660,N_1056);
nand U6382 (N_6382,N_4271,N_3229);
xor U6383 (N_6383,N_3091,N_195);
or U6384 (N_6384,N_4752,N_4723);
nand U6385 (N_6385,N_1420,N_1833);
nor U6386 (N_6386,N_1335,N_1888);
and U6387 (N_6387,N_848,N_1138);
nand U6388 (N_6388,N_1922,N_2497);
nor U6389 (N_6389,N_2202,N_3854);
or U6390 (N_6390,N_2514,N_4593);
or U6391 (N_6391,N_1744,N_824);
nor U6392 (N_6392,N_1137,N_973);
or U6393 (N_6393,N_1143,N_363);
nor U6394 (N_6394,N_272,N_3590);
and U6395 (N_6395,N_3564,N_313);
or U6396 (N_6396,N_2449,N_4062);
and U6397 (N_6397,N_470,N_2560);
nor U6398 (N_6398,N_4592,N_1943);
nor U6399 (N_6399,N_4746,N_2866);
and U6400 (N_6400,N_2452,N_1666);
and U6401 (N_6401,N_3957,N_1599);
and U6402 (N_6402,N_1061,N_2770);
nor U6403 (N_6403,N_982,N_8);
nand U6404 (N_6404,N_226,N_1284);
nand U6405 (N_6405,N_2544,N_4148);
or U6406 (N_6406,N_1036,N_1010);
nor U6407 (N_6407,N_4206,N_3684);
nor U6408 (N_6408,N_958,N_3204);
nor U6409 (N_6409,N_116,N_944);
or U6410 (N_6410,N_11,N_691);
nand U6411 (N_6411,N_4150,N_2378);
and U6412 (N_6412,N_3636,N_2120);
and U6413 (N_6413,N_3000,N_2871);
or U6414 (N_6414,N_471,N_4988);
or U6415 (N_6415,N_1134,N_4788);
or U6416 (N_6416,N_189,N_3297);
and U6417 (N_6417,N_3481,N_4973);
nor U6418 (N_6418,N_1403,N_3374);
and U6419 (N_6419,N_1750,N_992);
nand U6420 (N_6420,N_1644,N_2265);
nand U6421 (N_6421,N_4536,N_16);
nand U6422 (N_6422,N_143,N_4985);
nor U6423 (N_6423,N_3404,N_2711);
nand U6424 (N_6424,N_193,N_807);
and U6425 (N_6425,N_4572,N_1340);
and U6426 (N_6426,N_2608,N_1545);
nand U6427 (N_6427,N_3346,N_2417);
nor U6428 (N_6428,N_4341,N_3080);
and U6429 (N_6429,N_4434,N_1692);
nand U6430 (N_6430,N_1400,N_4561);
and U6431 (N_6431,N_3390,N_3398);
nor U6432 (N_6432,N_3028,N_1231);
nor U6433 (N_6433,N_1869,N_1621);
nor U6434 (N_6434,N_4115,N_3498);
nor U6435 (N_6435,N_3220,N_4469);
nand U6436 (N_6436,N_4750,N_139);
nand U6437 (N_6437,N_3343,N_4771);
and U6438 (N_6438,N_1306,N_2275);
nor U6439 (N_6439,N_2489,N_2333);
nor U6440 (N_6440,N_541,N_1830);
nand U6441 (N_6441,N_802,N_4276);
nor U6442 (N_6442,N_458,N_3740);
xor U6443 (N_6443,N_505,N_724);
or U6444 (N_6444,N_2623,N_1535);
nand U6445 (N_6445,N_599,N_3710);
or U6446 (N_6446,N_3845,N_136);
nor U6447 (N_6447,N_1963,N_4781);
nand U6448 (N_6448,N_2055,N_3832);
or U6449 (N_6449,N_4841,N_3331);
or U6450 (N_6450,N_1388,N_1967);
nor U6451 (N_6451,N_2650,N_2935);
nand U6452 (N_6452,N_3947,N_456);
or U6453 (N_6453,N_4979,N_1454);
nor U6454 (N_6454,N_3609,N_933);
nor U6455 (N_6455,N_4016,N_4719);
and U6456 (N_6456,N_3180,N_3783);
nor U6457 (N_6457,N_1606,N_3068);
or U6458 (N_6458,N_2563,N_3466);
nand U6459 (N_6459,N_821,N_4870);
nand U6460 (N_6460,N_679,N_2748);
nor U6461 (N_6461,N_3872,N_3838);
and U6462 (N_6462,N_1172,N_297);
nor U6463 (N_6463,N_3173,N_2593);
and U6464 (N_6464,N_4292,N_4745);
nor U6465 (N_6465,N_4196,N_1312);
nand U6466 (N_6466,N_697,N_2269);
nand U6467 (N_6467,N_4702,N_2367);
nand U6468 (N_6468,N_1476,N_946);
and U6469 (N_6469,N_4191,N_1102);
nand U6470 (N_6470,N_1900,N_1323);
nor U6471 (N_6471,N_717,N_2709);
nand U6472 (N_6472,N_4949,N_2063);
and U6473 (N_6473,N_2018,N_2474);
or U6474 (N_6474,N_4892,N_2652);
xnor U6475 (N_6475,N_2408,N_1207);
and U6476 (N_6476,N_4470,N_1768);
or U6477 (N_6477,N_572,N_2718);
or U6478 (N_6478,N_1423,N_368);
nand U6479 (N_6479,N_2141,N_3975);
and U6480 (N_6480,N_4904,N_1393);
xnor U6481 (N_6481,N_2239,N_1241);
nand U6482 (N_6482,N_690,N_466);
nor U6483 (N_6483,N_1775,N_1604);
and U6484 (N_6484,N_4172,N_915);
nand U6485 (N_6485,N_1444,N_628);
and U6486 (N_6486,N_4555,N_4960);
and U6487 (N_6487,N_3085,N_4655);
and U6488 (N_6488,N_2140,N_449);
nor U6489 (N_6489,N_240,N_1270);
and U6490 (N_6490,N_655,N_3295);
and U6491 (N_6491,N_1385,N_2988);
or U6492 (N_6492,N_2508,N_2200);
or U6493 (N_6493,N_1597,N_3664);
nand U6494 (N_6494,N_473,N_4924);
nor U6495 (N_6495,N_4263,N_1919);
nor U6496 (N_6496,N_566,N_1079);
or U6497 (N_6497,N_2116,N_39);
xnor U6498 (N_6498,N_1107,N_3757);
nand U6499 (N_6499,N_3319,N_4184);
nor U6500 (N_6500,N_4067,N_2761);
and U6501 (N_6501,N_1477,N_3970);
nor U6502 (N_6502,N_3676,N_623);
nor U6503 (N_6503,N_2462,N_841);
nand U6504 (N_6504,N_276,N_957);
or U6505 (N_6505,N_3182,N_2296);
or U6506 (N_6506,N_459,N_1624);
or U6507 (N_6507,N_1774,N_905);
and U6508 (N_6508,N_2583,N_3016);
nor U6509 (N_6509,N_3212,N_1162);
or U6510 (N_6510,N_1486,N_2586);
or U6511 (N_6511,N_4548,N_829);
and U6512 (N_6512,N_3013,N_1391);
and U6513 (N_6513,N_3192,N_1846);
nor U6514 (N_6514,N_1024,N_3162);
nor U6515 (N_6515,N_1776,N_1119);
and U6516 (N_6516,N_4123,N_3445);
nor U6517 (N_6517,N_516,N_4896);
nor U6518 (N_6518,N_440,N_1014);
or U6519 (N_6519,N_4288,N_2220);
or U6520 (N_6520,N_3818,N_4089);
nor U6521 (N_6521,N_2537,N_2456);
and U6522 (N_6522,N_378,N_259);
and U6523 (N_6523,N_1935,N_4441);
nor U6524 (N_6524,N_2323,N_3108);
and U6525 (N_6525,N_2588,N_4934);
nand U6526 (N_6526,N_1753,N_633);
and U6527 (N_6527,N_4266,N_2872);
nand U6528 (N_6528,N_781,N_2110);
and U6529 (N_6529,N_3864,N_746);
or U6530 (N_6530,N_1382,N_359);
nand U6531 (N_6531,N_1936,N_1527);
and U6532 (N_6532,N_3285,N_4080);
or U6533 (N_6533,N_2661,N_1588);
or U6534 (N_6534,N_4395,N_1217);
and U6535 (N_6535,N_2017,N_3881);
or U6536 (N_6536,N_663,N_3092);
nor U6537 (N_6537,N_1043,N_2261);
nand U6538 (N_6538,N_3596,N_3079);
nand U6539 (N_6539,N_301,N_4919);
nand U6540 (N_6540,N_2322,N_1474);
nand U6541 (N_6541,N_4295,N_2097);
or U6542 (N_6542,N_2035,N_3387);
nand U6543 (N_6543,N_1402,N_4060);
or U6544 (N_6544,N_1276,N_755);
nand U6545 (N_6545,N_1503,N_3999);
nor U6546 (N_6546,N_4628,N_174);
nand U6547 (N_6547,N_2266,N_972);
and U6548 (N_6548,N_17,N_1983);
and U6549 (N_6549,N_3890,N_1033);
or U6550 (N_6550,N_680,N_2328);
nor U6551 (N_6551,N_3262,N_4143);
nor U6552 (N_6552,N_4981,N_2271);
nor U6553 (N_6553,N_1716,N_814);
and U6554 (N_6554,N_1495,N_3605);
nand U6555 (N_6555,N_4459,N_4792);
or U6556 (N_6556,N_2371,N_2543);
nor U6557 (N_6557,N_2051,N_3062);
nand U6558 (N_6558,N_1959,N_4106);
nand U6559 (N_6559,N_565,N_3347);
nand U6560 (N_6560,N_4813,N_3839);
and U6561 (N_6561,N_1762,N_1209);
and U6562 (N_6562,N_4367,N_3169);
nand U6563 (N_6563,N_4694,N_411);
nor U6564 (N_6564,N_4840,N_784);
and U6565 (N_6565,N_2419,N_3239);
nand U6566 (N_6566,N_2171,N_380);
or U6567 (N_6567,N_2389,N_2160);
nand U6568 (N_6568,N_4366,N_1611);
nand U6569 (N_6569,N_3141,N_2730);
nor U6570 (N_6570,N_34,N_4509);
or U6571 (N_6571,N_3372,N_2168);
or U6572 (N_6572,N_3427,N_2175);
or U6573 (N_6573,N_1139,N_4243);
nand U6574 (N_6574,N_1896,N_4677);
nor U6575 (N_6575,N_813,N_4359);
nand U6576 (N_6576,N_3175,N_3311);
nand U6577 (N_6577,N_539,N_704);
and U6578 (N_6578,N_4000,N_3981);
and U6579 (N_6579,N_529,N_1572);
nor U6580 (N_6580,N_1215,N_384);
nor U6581 (N_6581,N_3614,N_4976);
nor U6582 (N_6582,N_3775,N_3467);
or U6583 (N_6583,N_3887,N_100);
and U6584 (N_6584,N_4091,N_1731);
nand U6585 (N_6585,N_3434,N_2093);
and U6586 (N_6586,N_1034,N_2102);
or U6587 (N_6587,N_142,N_4821);
or U6588 (N_6588,N_4529,N_58);
or U6589 (N_6589,N_443,N_901);
nor U6590 (N_6590,N_2069,N_4004);
or U6591 (N_6591,N_2345,N_4819);
nand U6592 (N_6592,N_3265,N_4169);
nor U6593 (N_6593,N_4504,N_1353);
and U6594 (N_6594,N_2716,N_1094);
and U6595 (N_6595,N_1751,N_4031);
nor U6596 (N_6596,N_3599,N_2235);
and U6597 (N_6597,N_830,N_3176);
nand U6598 (N_6598,N_3396,N_364);
and U6599 (N_6599,N_2725,N_1928);
nand U6600 (N_6600,N_4075,N_2813);
nor U6601 (N_6601,N_1456,N_1068);
nand U6602 (N_6602,N_2975,N_1372);
nor U6603 (N_6603,N_4595,N_3916);
and U6604 (N_6604,N_1648,N_385);
nor U6605 (N_6605,N_2864,N_1868);
nor U6606 (N_6606,N_3748,N_2375);
and U6607 (N_6607,N_3552,N_2702);
or U6608 (N_6608,N_1969,N_563);
or U6609 (N_6609,N_588,N_2430);
nor U6610 (N_6610,N_4850,N_2405);
or U6611 (N_6611,N_3117,N_4648);
nand U6612 (N_6612,N_811,N_3820);
nand U6613 (N_6613,N_3350,N_3058);
and U6614 (N_6614,N_651,N_9);
and U6615 (N_6615,N_2867,N_1472);
and U6616 (N_6616,N_4742,N_2783);
or U6617 (N_6617,N_4803,N_4758);
and U6618 (N_6618,N_1244,N_448);
nand U6619 (N_6619,N_3753,N_2012);
or U6620 (N_6620,N_3325,N_161);
or U6621 (N_6621,N_1106,N_3103);
and U6622 (N_6622,N_3666,N_4282);
and U6623 (N_6623,N_370,N_4085);
nand U6624 (N_6624,N_1023,N_1249);
or U6625 (N_6625,N_2948,N_2088);
and U6626 (N_6626,N_1460,N_4986);
and U6627 (N_6627,N_1979,N_2208);
and U6628 (N_6628,N_4168,N_119);
nand U6629 (N_6629,N_3892,N_2972);
and U6630 (N_6630,N_3129,N_0);
nand U6631 (N_6631,N_4463,N_3420);
and U6632 (N_6632,N_321,N_4721);
nand U6633 (N_6633,N_1089,N_4880);
and U6634 (N_6634,N_491,N_3074);
nor U6635 (N_6635,N_1668,N_1898);
nor U6636 (N_6636,N_324,N_1053);
nor U6637 (N_6637,N_4925,N_1971);
and U6638 (N_6638,N_981,N_2802);
and U6639 (N_6639,N_643,N_4514);
or U6640 (N_6640,N_3612,N_1101);
nor U6641 (N_6641,N_156,N_3622);
nand U6642 (N_6642,N_1721,N_4232);
and U6643 (N_6643,N_1265,N_2237);
nand U6644 (N_6644,N_2090,N_97);
or U6645 (N_6645,N_3402,N_4108);
and U6646 (N_6646,N_4117,N_4510);
nand U6647 (N_6647,N_2046,N_3312);
nor U6648 (N_6648,N_899,N_2295);
and U6649 (N_6649,N_4631,N_722);
xor U6650 (N_6650,N_2659,N_4733);
nor U6651 (N_6651,N_3616,N_1264);
or U6652 (N_6652,N_2435,N_916);
nand U6653 (N_6653,N_4913,N_3951);
nor U6654 (N_6654,N_472,N_1326);
or U6655 (N_6655,N_4891,N_40);
nor U6656 (N_6656,N_674,N_1880);
or U6657 (N_6657,N_4301,N_1870);
nand U6658 (N_6658,N_2665,N_3086);
nand U6659 (N_6659,N_2047,N_2227);
and U6660 (N_6660,N_888,N_2383);
nor U6661 (N_6661,N_2667,N_3691);
and U6662 (N_6662,N_3972,N_3056);
xnor U6663 (N_6663,N_1759,N_2847);
nand U6664 (N_6664,N_1021,N_4800);
nor U6665 (N_6665,N_1311,N_4667);
or U6666 (N_6666,N_225,N_2574);
nand U6667 (N_6667,N_3919,N_4513);
or U6668 (N_6668,N_3069,N_3243);
nor U6669 (N_6669,N_1506,N_4185);
nor U6670 (N_6670,N_520,N_801);
nand U6671 (N_6671,N_2106,N_2777);
nor U6672 (N_6672,N_4765,N_2996);
and U6673 (N_6673,N_4676,N_670);
and U6674 (N_6674,N_2011,N_810);
or U6675 (N_6675,N_3812,N_3066);
and U6676 (N_6676,N_1885,N_1461);
nand U6677 (N_6677,N_3008,N_165);
nor U6678 (N_6678,N_859,N_2998);
nor U6679 (N_6679,N_1421,N_783);
nand U6680 (N_6680,N_3807,N_1469);
or U6681 (N_6681,N_2163,N_4671);
and U6682 (N_6682,N_4679,N_4669);
nand U6683 (N_6683,N_1344,N_4755);
nor U6684 (N_6684,N_4397,N_1646);
or U6685 (N_6685,N_2960,N_3661);
nand U6686 (N_6686,N_699,N_3692);
and U6687 (N_6687,N_3778,N_2014);
or U6688 (N_6688,N_3802,N_325);
and U6689 (N_6689,N_435,N_2895);
or U6690 (N_6690,N_2728,N_3629);
and U6691 (N_6691,N_2904,N_3721);
nand U6692 (N_6692,N_3738,N_673);
and U6693 (N_6693,N_3559,N_3588);
nor U6694 (N_6694,N_2320,N_3353);
nand U6695 (N_6695,N_1854,N_3928);
or U6696 (N_6696,N_3899,N_1623);
or U6697 (N_6697,N_1934,N_2400);
or U6698 (N_6698,N_4319,N_3395);
and U6699 (N_6699,N_4570,N_481);
and U6700 (N_6700,N_1408,N_3852);
or U6701 (N_6701,N_1876,N_2258);
and U6702 (N_6702,N_1492,N_523);
and U6703 (N_6703,N_3924,N_4450);
nand U6704 (N_6704,N_2203,N_4704);
nor U6705 (N_6705,N_3979,N_1287);
and U6706 (N_6706,N_3719,N_422);
xor U6707 (N_6707,N_3324,N_1530);
and U6708 (N_6708,N_2941,N_3446);
or U6709 (N_6709,N_4542,N_4300);
nand U6710 (N_6710,N_750,N_4494);
nor U6711 (N_6711,N_3865,N_4693);
nand U6712 (N_6712,N_2465,N_1093);
nand U6713 (N_6713,N_741,N_877);
nand U6714 (N_6714,N_2363,N_4417);
and U6715 (N_6715,N_1560,N_3911);
nor U6716 (N_6716,N_4070,N_3101);
or U6717 (N_6717,N_2001,N_3247);
nand U6718 (N_6718,N_1363,N_4712);
or U6719 (N_6719,N_2023,N_4967);
nor U6720 (N_6720,N_644,N_2888);
nand U6721 (N_6721,N_1154,N_3492);
nor U6722 (N_6722,N_4347,N_367);
or U6723 (N_6723,N_4638,N_2414);
or U6724 (N_6724,N_2156,N_132);
or U6725 (N_6725,N_568,N_2853);
nand U6726 (N_6726,N_2148,N_874);
and U6727 (N_6727,N_1012,N_2211);
or U6728 (N_6728,N_3985,N_4447);
nor U6729 (N_6729,N_753,N_2974);
or U6730 (N_6730,N_3682,N_3089);
xor U6731 (N_6731,N_3188,N_2355);
or U6732 (N_6732,N_251,N_1369);
nand U6733 (N_6733,N_3905,N_2733);
and U6734 (N_6734,N_3834,N_3017);
and U6735 (N_6735,N_4562,N_3007);
xor U6736 (N_6736,N_1291,N_4703);
and U6737 (N_6737,N_2167,N_1332);
nor U6738 (N_6738,N_3843,N_365);
and U6739 (N_6739,N_1908,N_735);
or U6740 (N_6740,N_38,N_1008);
nand U6741 (N_6741,N_1571,N_1112);
nand U6742 (N_6742,N_561,N_4437);
and U6743 (N_6743,N_3121,N_2185);
nor U6744 (N_6744,N_2391,N_3884);
nor U6745 (N_6745,N_4253,N_1536);
nor U6746 (N_6746,N_2441,N_1377);
and U6747 (N_6747,N_1987,N_1582);
nor U6748 (N_6748,N_548,N_2151);
nor U6749 (N_6749,N_1279,N_1882);
nor U6750 (N_6750,N_1903,N_3798);
and U6751 (N_6751,N_789,N_4051);
nand U6752 (N_6752,N_4118,N_1416);
or U6753 (N_6753,N_4182,N_1155);
and U6754 (N_6754,N_361,N_347);
and U6755 (N_6755,N_2688,N_3218);
and U6756 (N_6756,N_954,N_4511);
nor U6757 (N_6757,N_1141,N_2964);
or U6758 (N_6758,N_2037,N_3922);
or U6759 (N_6759,N_2332,N_2264);
nor U6760 (N_6760,N_1690,N_4844);
or U6761 (N_6761,N_464,N_2846);
nor U6762 (N_6762,N_2119,N_630);
or U6763 (N_6763,N_170,N_911);
nor U6764 (N_6764,N_1278,N_2982);
and U6765 (N_6765,N_1780,N_1816);
xor U6766 (N_6766,N_1075,N_943);
nand U6767 (N_6767,N_3814,N_1451);
and U6768 (N_6768,N_3515,N_2438);
nor U6769 (N_6769,N_733,N_3094);
nand U6770 (N_6770,N_334,N_1438);
or U6771 (N_6771,N_2198,N_2306);
or U6772 (N_6772,N_1455,N_2976);
nor U6773 (N_6773,N_1664,N_3456);
or U6774 (N_6774,N_3789,N_929);
and U6775 (N_6775,N_1070,N_1275);
nor U6776 (N_6776,N_4439,N_793);
nor U6777 (N_6777,N_218,N_1044);
and U6778 (N_6778,N_453,N_3111);
nor U6779 (N_6779,N_2043,N_3430);
nand U6780 (N_6780,N_1087,N_3773);
or U6781 (N_6781,N_3765,N_4852);
and U6782 (N_6782,N_4666,N_3326);
and U6783 (N_6783,N_1632,N_360);
and U6784 (N_6784,N_1205,N_1609);
or U6785 (N_6785,N_4722,N_2196);
nand U6786 (N_6786,N_3920,N_2176);
or U6787 (N_6787,N_2658,N_1931);
nor U6788 (N_6788,N_2993,N_3315);
and U6789 (N_6789,N_1011,N_546);
or U6790 (N_6790,N_2020,N_2195);
and U6791 (N_6791,N_222,N_2571);
nand U6792 (N_6792,N_920,N_968);
nand U6793 (N_6793,N_2913,N_3779);
nand U6794 (N_6794,N_1236,N_3529);
or U6795 (N_6795,N_2736,N_2607);
nor U6796 (N_6796,N_4582,N_3542);
nor U6797 (N_6797,N_3955,N_3965);
or U6798 (N_6798,N_2699,N_2146);
and U6799 (N_6799,N_3438,N_4848);
nand U6800 (N_6800,N_1773,N_4989);
and U6801 (N_6801,N_1001,N_780);
or U6802 (N_6802,N_209,N_1549);
or U6803 (N_6803,N_2918,N_172);
or U6804 (N_6804,N_4379,N_4633);
nor U6805 (N_6805,N_1341,N_2969);
or U6806 (N_6806,N_4773,N_3987);
and U6807 (N_6807,N_3435,N_935);
nor U6808 (N_6808,N_3339,N_234);
nor U6809 (N_6809,N_3024,N_4486);
nor U6810 (N_6810,N_1650,N_1652);
nand U6811 (N_6811,N_2406,N_394);
and U6812 (N_6812,N_4710,N_4997);
or U6813 (N_6813,N_354,N_4535);
or U6814 (N_6814,N_596,N_1434);
or U6815 (N_6815,N_737,N_87);
and U6816 (N_6816,N_2123,N_945);
and U6817 (N_6817,N_4203,N_1459);
nand U6818 (N_6818,N_2747,N_3252);
nand U6819 (N_6819,N_2981,N_212);
and U6820 (N_6820,N_3137,N_1463);
or U6821 (N_6821,N_371,N_1475);
and U6822 (N_6822,N_256,N_1229);
or U6823 (N_6823,N_4948,N_966);
or U6824 (N_6824,N_3268,N_3266);
nor U6825 (N_6825,N_2555,N_4932);
and U6826 (N_6826,N_1910,N_339);
and U6827 (N_6827,N_712,N_4554);
and U6828 (N_6828,N_4817,N_4653);
nand U6829 (N_6829,N_1875,N_4389);
or U6830 (N_6830,N_2177,N_2132);
or U6831 (N_6831,N_1729,N_2955);
or U6832 (N_6832,N_350,N_1083);
or U6833 (N_6833,N_4053,N_4084);
and U6834 (N_6834,N_1542,N_969);
and U6835 (N_6835,N_799,N_4673);
nor U6836 (N_6836,N_884,N_4269);
nand U6837 (N_6837,N_786,N_2191);
and U6838 (N_6838,N_1450,N_3310);
or U6839 (N_6839,N_1515,N_2480);
or U6840 (N_6840,N_1494,N_3727);
nor U6841 (N_6841,N_3749,N_2472);
nand U6842 (N_6842,N_3904,N_3716);
nor U6843 (N_6843,N_1941,N_1046);
or U6844 (N_6844,N_4996,N_1462);
and U6845 (N_6845,N_3944,N_4357);
or U6846 (N_6846,N_4478,N_4457);
nand U6847 (N_6847,N_4930,N_1250);
or U6848 (N_6848,N_2315,N_3907);
nand U6849 (N_6849,N_4453,N_2214);
nor U6850 (N_6850,N_3927,N_2999);
nand U6851 (N_6851,N_2842,N_562);
nor U6852 (N_6852,N_2129,N_4756);
and U6853 (N_6853,N_1221,N_457);
or U6854 (N_6854,N_891,N_940);
nor U6855 (N_6855,N_1581,N_1725);
and U6856 (N_6856,N_1471,N_918);
nor U6857 (N_6857,N_3640,N_3355);
nor U6858 (N_6858,N_1635,N_2524);
nor U6859 (N_6859,N_4312,N_1013);
xor U6860 (N_6860,N_4173,N_3384);
nor U6861 (N_6861,N_514,N_3216);
nor U6862 (N_6862,N_519,N_4107);
nor U6863 (N_6863,N_181,N_2953);
nor U6864 (N_6864,N_601,N_1673);
nor U6865 (N_6865,N_2696,N_1020);
or U6866 (N_6866,N_4305,N_3658);
and U6867 (N_6867,N_2233,N_2979);
nor U6868 (N_6868,N_1602,N_496);
nor U6869 (N_6869,N_815,N_4370);
and U6870 (N_6870,N_1328,N_3035);
or U6871 (N_6871,N_4877,N_667);
or U6872 (N_6872,N_3083,N_2727);
nor U6873 (N_6873,N_1891,N_3484);
and U6874 (N_6874,N_3675,N_3279);
or U6875 (N_6875,N_52,N_2815);
nor U6876 (N_6876,N_570,N_4886);
and U6877 (N_6877,N_4059,N_3555);
xnor U6878 (N_6878,N_879,N_3949);
or U6879 (N_6879,N_1998,N_1997);
nor U6880 (N_6880,N_341,N_2024);
and U6881 (N_6881,N_3014,N_4414);
and U6882 (N_6882,N_3090,N_415);
nor U6883 (N_6883,N_886,N_500);
nand U6884 (N_6884,N_4464,N_4360);
nand U6885 (N_6885,N_3690,N_1860);
and U6886 (N_6886,N_4283,N_797);
nor U6887 (N_6887,N_4421,N_4159);
nand U6888 (N_6888,N_1713,N_990);
and U6889 (N_6889,N_3333,N_3251);
or U6890 (N_6890,N_1578,N_1957);
or U6891 (N_6891,N_3051,N_3330);
and U6892 (N_6892,N_328,N_985);
or U6893 (N_6893,N_4325,N_778);
nand U6894 (N_6894,N_1895,N_604);
and U6895 (N_6895,N_3230,N_74);
nor U6896 (N_6896,N_2547,N_4045);
nand U6897 (N_6897,N_3100,N_103);
and U6898 (N_6898,N_2678,N_4726);
nand U6899 (N_6899,N_1066,N_253);
nor U6900 (N_6900,N_3825,N_3799);
or U6901 (N_6901,N_2513,N_188);
or U6902 (N_6902,N_1170,N_2754);
and U6903 (N_6903,N_4720,N_3156);
or U6904 (N_6904,N_574,N_1807);
nor U6905 (N_6905,N_1918,N_4517);
nor U6906 (N_6906,N_3150,N_2987);
nor U6907 (N_6907,N_4013,N_2801);
or U6908 (N_6908,N_4386,N_2221);
nor U6909 (N_6909,N_2215,N_1248);
nand U6910 (N_6910,N_3583,N_166);
or U6911 (N_6911,N_3857,N_721);
and U6912 (N_6912,N_3514,N_2995);
nor U6913 (N_6913,N_37,N_2534);
and U6914 (N_6914,N_1992,N_4971);
and U6915 (N_6915,N_3709,N_2062);
or U6916 (N_6916,N_3501,N_1568);
xor U6917 (N_6917,N_1873,N_4214);
nand U6918 (N_6918,N_382,N_1890);
nand U6919 (N_6919,N_134,N_2868);
and U6920 (N_6920,N_3626,N_4245);
nor U6921 (N_6921,N_1863,N_2739);
or U6922 (N_6922,N_2558,N_4537);
or U6923 (N_6923,N_2878,N_1065);
nor U6924 (N_6924,N_1299,N_2403);
and U6925 (N_6925,N_987,N_2337);
or U6926 (N_6926,N_4229,N_1831);
nor U6927 (N_6927,N_2199,N_754);
and U6928 (N_6928,N_4121,N_3244);
nor U6929 (N_6929,N_476,N_584);
nand U6930 (N_6930,N_785,N_3836);
nand U6931 (N_6931,N_77,N_1857);
and U6932 (N_6932,N_1823,N_1184);
nand U6933 (N_6933,N_3138,N_4680);
nor U6934 (N_6934,N_2881,N_2861);
and U6935 (N_6935,N_3722,N_4836);
nand U6936 (N_6936,N_4451,N_3208);
or U6937 (N_6937,N_4316,N_4387);
or U6938 (N_6938,N_2437,N_3673);
nor U6939 (N_6939,N_33,N_840);
and U6940 (N_6940,N_169,N_2412);
nor U6941 (N_6941,N_2792,N_2787);
nand U6942 (N_6942,N_2057,N_3547);
nand U6943 (N_6943,N_1374,N_3901);
nand U6944 (N_6944,N_1784,N_204);
and U6945 (N_6945,N_3469,N_41);
and U6946 (N_6946,N_1950,N_2549);
and U6947 (N_6947,N_4965,N_1442);
or U6948 (N_6948,N_1676,N_3880);
and U6949 (N_6949,N_4650,N_2655);
and U6950 (N_6950,N_1600,N_756);
nor U6951 (N_6951,N_1537,N_4747);
nor U6952 (N_6952,N_3273,N_4430);
and U6953 (N_6953,N_474,N_434);
and U6954 (N_6954,N_1466,N_1827);
or U6955 (N_6955,N_2384,N_3931);
or U6956 (N_6956,N_3106,N_731);
nand U6957 (N_6957,N_858,N_3010);
and U6958 (N_6958,N_2459,N_4632);
nor U6959 (N_6959,N_230,N_4575);
and U6960 (N_6960,N_1741,N_2638);
and U6961 (N_6961,N_4287,N_569);
nand U6962 (N_6962,N_2597,N_4791);
nand U6963 (N_6963,N_3167,N_598);
nor U6964 (N_6964,N_1387,N_2664);
nor U6965 (N_6965,N_4516,N_3809);
nand U6966 (N_6966,N_4678,N_3122);
nor U6967 (N_6967,N_806,N_114);
or U6968 (N_6968,N_682,N_2344);
nand U6969 (N_6969,N_3179,N_4888);
nand U6970 (N_6970,N_3539,N_1202);
and U6971 (N_6971,N_2143,N_4489);
and U6972 (N_6972,N_834,N_932);
and U6973 (N_6973,N_506,N_2121);
nor U6974 (N_6974,N_3611,N_792);
nand U6975 (N_6975,N_3821,N_4001);
or U6976 (N_6976,N_314,N_2254);
or U6977 (N_6977,N_3221,N_277);
and U6978 (N_6978,N_1834,N_1671);
or U6979 (N_6979,N_2440,N_2335);
nor U6980 (N_6980,N_2169,N_2700);
or U6981 (N_6981,N_701,N_2850);
nand U6982 (N_6982,N_3886,N_2095);
xor U6983 (N_6983,N_524,N_515);
or U6984 (N_6984,N_4866,N_2283);
nand U6985 (N_6985,N_4825,N_1204);
nand U6986 (N_6986,N_3032,N_4177);
and U6987 (N_6987,N_1912,N_3950);
nor U6988 (N_6988,N_3232,N_1858);
and U6989 (N_6989,N_4842,N_2084);
nor U6990 (N_6990,N_4697,N_1358);
nor U6991 (N_6991,N_425,N_2751);
and U6992 (N_6992,N_4130,N_2226);
nor U6993 (N_6993,N_997,N_469);
or U6994 (N_6994,N_609,N_271);
nor U6995 (N_6995,N_4344,N_3844);
or U6996 (N_6996,N_2086,N_1569);
nand U6997 (N_6997,N_2944,N_662);
nand U6998 (N_6998,N_4601,N_3088);
nor U6999 (N_6999,N_3240,N_4779);
nor U7000 (N_7000,N_1441,N_1268);
or U7001 (N_7001,N_2618,N_827);
and U7002 (N_7002,N_4381,N_1877);
or U7003 (N_7003,N_3148,N_2361);
nor U7004 (N_7004,N_554,N_2238);
nor U7005 (N_7005,N_4023,N_3392);
nand U7006 (N_7006,N_1499,N_2230);
and U7007 (N_7007,N_1360,N_1419);
or U7008 (N_7008,N_23,N_4515);
nor U7009 (N_7009,N_1874,N_4488);
or U7010 (N_7010,N_2694,N_4205);
and U7011 (N_7011,N_2301,N_3397);
nand U7012 (N_7012,N_2521,N_2545);
or U7013 (N_7013,N_4662,N_1277);
or U7014 (N_7014,N_4158,N_1909);
and U7015 (N_7015,N_2970,N_4286);
nand U7016 (N_7016,N_268,N_4659);
or U7017 (N_7017,N_3646,N_2640);
nor U7018 (N_7018,N_522,N_2714);
nand U7019 (N_7019,N_1120,N_255);
or U7020 (N_7020,N_1800,N_1984);
nand U7021 (N_7021,N_4910,N_369);
nand U7022 (N_7022,N_2030,N_3705);
nor U7023 (N_7023,N_3413,N_1792);
nor U7024 (N_7024,N_1573,N_1738);
nor U7025 (N_7025,N_4901,N_839);
nor U7026 (N_7026,N_962,N_1590);
nand U7027 (N_7027,N_1962,N_3874);
and U7028 (N_7028,N_468,N_2710);
and U7029 (N_7029,N_4029,N_284);
and U7030 (N_7030,N_1286,N_3318);
or U7031 (N_7031,N_2532,N_3011);
or U7032 (N_7032,N_2310,N_774);
nand U7033 (N_7033,N_4324,N_4220);
or U7034 (N_7034,N_416,N_32);
and U7035 (N_7035,N_2287,N_3763);
or U7036 (N_7036,N_2348,N_63);
and U7037 (N_7037,N_3323,N_4064);
or U7038 (N_7038,N_3142,N_3105);
or U7039 (N_7039,N_4378,N_4320);
nand U7040 (N_7040,N_3718,N_4577);
nor U7041 (N_7041,N_816,N_2231);
nor U7042 (N_7042,N_291,N_4605);
nand U7043 (N_7043,N_4446,N_1584);
nor U7044 (N_7044,N_3634,N_4772);
nor U7045 (N_7045,N_14,N_4188);
nand U7046 (N_7046,N_4587,N_3729);
and U7047 (N_7047,N_1544,N_4957);
or U7048 (N_7048,N_4947,N_2073);
nor U7049 (N_7049,N_1715,N_1285);
nor U7050 (N_7050,N_3057,N_687);
nand U7051 (N_7051,N_1255,N_3522);
nand U7052 (N_7052,N_4861,N_2256);
or U7053 (N_7053,N_1337,N_836);
or U7054 (N_7054,N_989,N_1113);
and U7055 (N_7055,N_1742,N_740);
and U7056 (N_7056,N_2321,N_3341);
nor U7057 (N_7057,N_4066,N_1283);
nand U7058 (N_7058,N_1654,N_309);
nand U7059 (N_7059,N_1422,N_2971);
or U7060 (N_7060,N_389,N_51);
or U7061 (N_7061,N_3647,N_4401);
nand U7062 (N_7062,N_970,N_3726);
nand U7063 (N_7063,N_4267,N_718);
and U7064 (N_7064,N_3288,N_4015);
or U7065 (N_7065,N_4622,N_1649);
nor U7066 (N_7066,N_83,N_1675);
or U7067 (N_7067,N_2466,N_2180);
nand U7068 (N_7068,N_2942,N_2915);
or U7069 (N_7069,N_4297,N_4093);
nand U7070 (N_7070,N_3077,N_776);
nor U7071 (N_7071,N_2691,N_650);
and U7072 (N_7072,N_1541,N_3963);
nor U7073 (N_7073,N_2511,N_335);
or U7074 (N_7074,N_2118,N_4566);
nand U7075 (N_7075,N_540,N_4037);
and U7076 (N_7076,N_101,N_3439);
nand U7077 (N_7077,N_3184,N_892);
and U7078 (N_7078,N_3642,N_4258);
xnor U7079 (N_7079,N_4775,N_4095);
and U7080 (N_7080,N_771,N_1951);
or U7081 (N_7081,N_3457,N_2016);
nand U7082 (N_7082,N_1539,N_3969);
or U7083 (N_7083,N_2923,N_1902);
and U7084 (N_7084,N_2707,N_1522);
and U7085 (N_7085,N_4972,N_2273);
and U7086 (N_7086,N_3352,N_3276);
nand U7087 (N_7087,N_2758,N_4522);
or U7088 (N_7088,N_4815,N_1897);
or U7089 (N_7089,N_1294,N_4250);
nor U7090 (N_7090,N_2219,N_1302);
nand U7091 (N_7091,N_4643,N_3511);
nor U7092 (N_7092,N_1405,N_2068);
nand U7093 (N_7093,N_2504,N_2880);
nand U7094 (N_7094,N_1174,N_265);
nand U7095 (N_7095,N_818,N_4942);
nor U7096 (N_7096,N_2490,N_2690);
and U7097 (N_7097,N_3630,N_3742);
nand U7098 (N_7098,N_1006,N_1740);
nand U7099 (N_7099,N_555,N_280);
or U7100 (N_7100,N_3443,N_4994);
and U7101 (N_7101,N_936,N_3441);
and U7102 (N_7102,N_3827,N_4260);
nand U7103 (N_7103,N_2172,N_3185);
nand U7104 (N_7104,N_4597,N_937);
nand U7105 (N_7105,N_2529,N_4737);
and U7106 (N_7106,N_2540,N_3174);
nand U7107 (N_7107,N_1171,N_396);
or U7108 (N_7108,N_1032,N_1627);
and U7109 (N_7109,N_826,N_3261);
nand U7110 (N_7110,N_1428,N_3236);
or U7111 (N_7111,N_4881,N_4178);
or U7112 (N_7112,N_1246,N_531);
nand U7113 (N_7113,N_758,N_4296);
nor U7114 (N_7114,N_131,N_2991);
or U7115 (N_7115,N_4890,N_3575);
nand U7116 (N_7116,N_4038,N_4606);
and U7117 (N_7117,N_4623,N_1836);
nand U7118 (N_7118,N_4759,N_3193);
or U7119 (N_7119,N_2107,N_1789);
nand U7120 (N_7120,N_164,N_4371);
nor U7121 (N_7121,N_4684,N_68);
nand U7122 (N_7122,N_1212,N_3135);
and U7123 (N_7123,N_4991,N_705);
nor U7124 (N_7124,N_3902,N_666);
nor U7125 (N_7125,N_393,N_4828);
or U7126 (N_7126,N_4249,N_4048);
nand U7127 (N_7127,N_2626,N_3264);
nor U7128 (N_7128,N_3744,N_808);
nand U7129 (N_7129,N_2189,N_286);
nor U7130 (N_7130,N_3694,N_1927);
nor U7131 (N_7131,N_804,N_4240);
nor U7132 (N_7132,N_3909,N_4435);
nand U7133 (N_7133,N_3189,N_853);
and U7134 (N_7134,N_4946,N_3052);
or U7135 (N_7135,N_4968,N_1976);
nand U7136 (N_7136,N_1973,N_1614);
or U7137 (N_7137,N_2415,N_600);
nor U7138 (N_7138,N_3419,N_728);
and U7139 (N_7139,N_4724,N_4365);
or U7140 (N_7140,N_3610,N_3414);
nor U7141 (N_7141,N_3061,N_2952);
and U7142 (N_7142,N_942,N_1211);
nand U7143 (N_7143,N_3678,N_3269);
and U7144 (N_7144,N_3667,N_4812);
and U7145 (N_7145,N_3465,N_3732);
or U7146 (N_7146,N_140,N_3340);
nand U7147 (N_7147,N_3418,N_2911);
and U7148 (N_7148,N_308,N_3711);
or U7149 (N_7149,N_3191,N_3458);
and U7150 (N_7150,N_3786,N_4621);
nand U7151 (N_7151,N_1783,N_4652);
or U7152 (N_7152,N_4318,N_61);
or U7153 (N_7153,N_356,N_2546);
or U7154 (N_7154,N_3059,N_1132);
or U7155 (N_7155,N_3038,N_1812);
or U7156 (N_7156,N_2356,N_2641);
nand U7157 (N_7157,N_133,N_1239);
nand U7158 (N_7158,N_4135,N_4465);
nand U7159 (N_7159,N_2639,N_1667);
nor U7160 (N_7160,N_2721,N_3768);
or U7161 (N_7161,N_130,N_1352);
and U7162 (N_7162,N_4217,N_4337);
and U7163 (N_7163,N_349,N_2228);
or U7164 (N_7164,N_1223,N_1179);
nand U7165 (N_7165,N_579,N_3300);
nand U7166 (N_7166,N_1243,N_4589);
nor U7167 (N_7167,N_4302,N_4651);
or U7168 (N_7168,N_1972,N_847);
and U7169 (N_7169,N_105,N_395);
nor U7170 (N_7170,N_2788,N_264);
or U7171 (N_7171,N_3391,N_4978);
nand U7172 (N_7172,N_931,N_4727);
or U7173 (N_7173,N_2622,N_849);
nor U7174 (N_7174,N_4407,N_4596);
or U7175 (N_7175,N_4649,N_1298);
nor U7176 (N_7176,N_3913,N_4620);
or U7177 (N_7177,N_1045,N_1930);
and U7178 (N_7178,N_924,N_2701);
nand U7179 (N_7179,N_266,N_3429);
nor U7180 (N_7180,N_3289,N_2005);
and U7181 (N_7181,N_4999,N_2875);
nand U7182 (N_7182,N_3752,N_1314);
nand U7183 (N_7183,N_4256,N_2862);
and U7184 (N_7184,N_1705,N_1778);
nand U7185 (N_7185,N_1808,N_3540);
nor U7186 (N_7186,N_4097,N_4380);
nand U7187 (N_7187,N_3447,N_3126);
or U7188 (N_7188,N_4731,N_177);
nand U7189 (N_7189,N_4859,N_1364);
and U7190 (N_7190,N_1637,N_1589);
nand U7191 (N_7191,N_2619,N_414);
and U7192 (N_7192,N_430,N_597);
or U7193 (N_7193,N_3203,N_4207);
and U7194 (N_7194,N_4496,N_2381);
nor U7195 (N_7195,N_283,N_1563);
and U7196 (N_7196,N_4165,N_2849);
nor U7197 (N_7197,N_4521,N_2824);
nand U7198 (N_7198,N_1433,N_1754);
nor U7199 (N_7199,N_1736,N_2873);
nor U7200 (N_7200,N_2879,N_2394);
nand U7201 (N_7201,N_2288,N_4333);
xnor U7202 (N_7202,N_3081,N_4897);
and U7203 (N_7203,N_4526,N_1361);
or U7204 (N_7204,N_2523,N_479);
nor U7205 (N_7205,N_1489,N_2281);
nor U7206 (N_7206,N_3277,N_2502);
or U7207 (N_7207,N_1709,N_3937);
or U7208 (N_7208,N_4445,N_913);
and U7209 (N_7209,N_4003,N_2326);
nand U7210 (N_7210,N_4739,N_1804);
and U7211 (N_7211,N_2857,N_2338);
and U7212 (N_7212,N_4943,N_3292);
nand U7213 (N_7213,N_3868,N_1795);
nand U7214 (N_7214,N_1685,N_3102);
and U7215 (N_7215,N_2625,N_3731);
and U7216 (N_7216,N_2085,N_2134);
nand U7217 (N_7217,N_2822,N_2039);
nand U7218 (N_7218,N_2178,N_261);
nor U7219 (N_7219,N_2819,N_1496);
and U7220 (N_7220,N_3031,N_4293);
or U7221 (N_7221,N_4807,N_4951);
nor U7222 (N_7222,N_1949,N_889);
nor U7223 (N_7223,N_305,N_1418);
or U7224 (N_7224,N_4354,N_1225);
nand U7225 (N_7225,N_1528,N_3226);
nor U7226 (N_7226,N_1401,N_406);
nand U7227 (N_7227,N_2396,N_3751);
or U7228 (N_7228,N_373,N_2729);
nand U7229 (N_7229,N_306,N_1114);
nand U7230 (N_7230,N_3490,N_203);
nor U7231 (N_7231,N_664,N_3112);
or U7232 (N_7232,N_1517,N_445);
and U7233 (N_7233,N_2553,N_1932);
nand U7234 (N_7234,N_3107,N_3746);
and U7235 (N_7235,N_1889,N_214);
and U7236 (N_7236,N_1613,N_1095);
nor U7237 (N_7237,N_4851,N_3597);
or U7238 (N_7238,N_1343,N_4927);
nor U7239 (N_7239,N_4585,N_4987);
or U7240 (N_7240,N_4114,N_3918);
or U7241 (N_7241,N_4340,N_549);
nor U7242 (N_7242,N_70,N_4952);
nor U7243 (N_7243,N_93,N_2424);
nor U7244 (N_7244,N_4028,N_1630);
and U7245 (N_7245,N_2519,N_999);
nand U7246 (N_7246,N_1467,N_2259);
nand U7247 (N_7247,N_2954,N_450);
and U7248 (N_7248,N_3935,N_544);
nand U7249 (N_7249,N_4626,N_3233);
or U7250 (N_7250,N_2891,N_4931);
and U7251 (N_7251,N_3517,N_3298);
or U7252 (N_7252,N_4399,N_2776);
nor U7253 (N_7253,N_2590,N_1881);
or U7254 (N_7254,N_661,N_1237);
and U7255 (N_7255,N_176,N_510);
or U7256 (N_7256,N_3222,N_4209);
and U7257 (N_7257,N_1956,N_4368);
or U7258 (N_7258,N_3945,N_4094);
nor U7259 (N_7259,N_92,N_405);
nand U7260 (N_7260,N_85,N_3534);
nor U7261 (N_7261,N_1300,N_4230);
and U7262 (N_7262,N_3452,N_1049);
nand U7263 (N_7263,N_4627,N_4547);
or U7264 (N_7264,N_2767,N_1041);
or U7265 (N_7265,N_1366,N_4682);
nand U7266 (N_7266,N_4426,N_2556);
or U7267 (N_7267,N_3012,N_4140);
nor U7268 (N_7268,N_4454,N_3304);
nand U7269 (N_7269,N_904,N_4284);
and U7270 (N_7270,N_3078,N_42);
nand U7271 (N_7271,N_1594,N_2263);
nor U7272 (N_7272,N_895,N_3245);
nor U7273 (N_7273,N_3932,N_69);
and U7274 (N_7274,N_543,N_4909);
and U7275 (N_7275,N_4144,N_3140);
and U7276 (N_7276,N_3557,N_19);
nor U7277 (N_7277,N_2352,N_3855);
nand U7278 (N_7278,N_2840,N_123);
and U7279 (N_7279,N_2379,N_4969);
nand U7280 (N_7280,N_4950,N_2568);
nor U7281 (N_7281,N_3303,N_1990);
or U7282 (N_7282,N_2520,N_4088);
or U7283 (N_7283,N_1197,N_2865);
nand U7284 (N_7284,N_1198,N_4705);
and U7285 (N_7285,N_4574,N_112);
or U7286 (N_7286,N_653,N_714);
and U7287 (N_7287,N_882,N_4129);
or U7288 (N_7288,N_3099,N_3730);
and U7289 (N_7289,N_4092,N_1867);
and U7290 (N_7290,N_2170,N_2034);
or U7291 (N_7291,N_3762,N_3697);
and U7292 (N_7292,N_922,N_3200);
nor U7293 (N_7293,N_4131,N_1073);
nand U7294 (N_7294,N_3470,N_1208);
nand U7295 (N_7295,N_2158,N_1947);
nor U7296 (N_7296,N_4189,N_706);
or U7297 (N_7297,N_3545,N_921);
or U7298 (N_7298,N_377,N_917);
nor U7299 (N_7299,N_2966,N_4090);
or U7300 (N_7300,N_3361,N_2579);
nor U7301 (N_7301,N_4754,N_3486);
and U7302 (N_7302,N_2277,N_696);
or U7303 (N_7303,N_4921,N_4137);
nor U7304 (N_7304,N_4715,N_2668);
and U7305 (N_7305,N_3197,N_878);
or U7306 (N_7306,N_3219,N_2968);
or U7307 (N_7307,N_2909,N_2799);
or U7308 (N_7308,N_775,N_1104);
or U7309 (N_7309,N_1620,N_4541);
nor U7310 (N_7310,N_2099,N_1550);
nand U7311 (N_7311,N_4223,N_2390);
nor U7312 (N_7312,N_3850,N_4042);
nand U7313 (N_7313,N_2100,N_3345);
nor U7314 (N_7314,N_4458,N_873);
or U7315 (N_7315,N_782,N_4257);
and U7316 (N_7316,N_3801,N_147);
nand U7317 (N_7317,N_4865,N_2899);
nor U7318 (N_7318,N_1861,N_2382);
or U7319 (N_7319,N_4583,N_2887);
or U7320 (N_7320,N_2859,N_1058);
and U7321 (N_7321,N_1271,N_2587);
nor U7322 (N_7322,N_3334,N_2329);
nand U7323 (N_7323,N_1396,N_4179);
or U7324 (N_7324,N_463,N_4823);
nand U7325 (N_7325,N_4375,N_1148);
or U7326 (N_7326,N_1274,N_683);
or U7327 (N_7327,N_1538,N_2133);
or U7328 (N_7328,N_1699,N_3524);
nor U7329 (N_7329,N_2916,N_3687);
nor U7330 (N_7330,N_4630,N_3381);
or U7331 (N_7331,N_719,N_1318);
nand U7332 (N_7332,N_3026,N_4941);
or U7333 (N_7333,N_2091,N_2245);
and U7334 (N_7334,N_3990,N_4141);
nand U7335 (N_7335,N_2457,N_3713);
or U7336 (N_7336,N_2327,N_4992);
and U7337 (N_7337,N_2604,N_4958);
or U7338 (N_7338,N_3796,N_578);
nand U7339 (N_7339,N_2386,N_953);
and U7340 (N_7340,N_3407,N_4246);
xnor U7341 (N_7341,N_29,N_2893);
nand U7342 (N_7342,N_1587,N_1149);
and U7343 (N_7343,N_3654,N_991);
and U7344 (N_7344,N_3202,N_4322);
nor U7345 (N_7345,N_2569,N_2157);
and U7346 (N_7346,N_3171,N_822);
nand U7347 (N_7347,N_2049,N_2542);
and U7348 (N_7348,N_1847,N_2232);
and U7349 (N_7349,N_2973,N_723);
nor U7350 (N_7350,N_1755,N_4884);
nand U7351 (N_7351,N_4558,N_2677);
xor U7352 (N_7352,N_689,N_1167);
nor U7353 (N_7353,N_1322,N_1293);
nor U7354 (N_7354,N_3521,N_614);
and U7355 (N_7355,N_210,N_236);
nor U7356 (N_7356,N_4152,N_2431);
nand U7357 (N_7357,N_3569,N_4420);
nor U7358 (N_7358,N_2305,N_2687);
and U7359 (N_7359,N_3953,N_1665);
and U7360 (N_7360,N_2444,N_3382);
nor U7361 (N_7361,N_4369,N_1123);
nor U7362 (N_7362,N_4218,N_1821);
nand U7363 (N_7363,N_3586,N_2884);
and U7364 (N_7364,N_122,N_3828);
and U7365 (N_7365,N_1190,N_4498);
nand U7366 (N_7366,N_343,N_2416);
nor U7367 (N_7367,N_2407,N_1638);
or U7368 (N_7368,N_4826,N_3504);
nor U7369 (N_7369,N_1166,N_4111);
nand U7370 (N_7370,N_30,N_2898);
and U7371 (N_7371,N_1559,N_1929);
nor U7372 (N_7372,N_2643,N_762);
or U7373 (N_7373,N_1926,N_4546);
nor U7374 (N_7374,N_4853,N_2735);
or U7375 (N_7375,N_2128,N_4161);
nor U7376 (N_7376,N_318,N_2216);
or U7377 (N_7377,N_3651,N_3914);
or U7378 (N_7378,N_1767,N_2992);
or U7379 (N_7379,N_2646,N_1641);
nand U7380 (N_7380,N_2186,N_2939);
nor U7381 (N_7381,N_2426,N_4923);
and U7382 (N_7382,N_3971,N_1960);
nor U7383 (N_7383,N_2343,N_2418);
or U7384 (N_7384,N_3337,N_627);
nand U7385 (N_7385,N_2516,N_148);
nor U7386 (N_7386,N_591,N_869);
or U7387 (N_7387,N_4174,N_3723);
and U7388 (N_7388,N_509,N_3720);
nor U7389 (N_7389,N_2536,N_3652);
and U7390 (N_7390,N_1350,N_4073);
nand U7391 (N_7391,N_2108,N_2719);
or U7392 (N_7392,N_3365,N_1626);
or U7393 (N_7393,N_381,N_2339);
and U7394 (N_7394,N_3145,N_710);
and U7395 (N_7395,N_3149,N_4077);
nand U7396 (N_7396,N_1786,N_151);
nor U7397 (N_7397,N_4564,N_262);
and U7398 (N_7398,N_3925,N_2145);
or U7399 (N_7399,N_154,N_787);
nor U7400 (N_7400,N_1781,N_902);
nor U7401 (N_7401,N_2353,N_2631);
or U7402 (N_7402,N_3817,N_1980);
or U7403 (N_7403,N_872,N_2548);
nand U7404 (N_7404,N_4714,N_1281);
and U7405 (N_7405,N_2989,N_507);
and U7406 (N_7406,N_4307,N_3128);
or U7407 (N_7407,N_1561,N_583);
and U7408 (N_7408,N_1761,N_1782);
nand U7409 (N_7409,N_2308,N_1917);
and U7410 (N_7410,N_2763,N_3871);
and U7411 (N_7411,N_736,N_923);
or U7412 (N_7412,N_2278,N_1526);
and U7413 (N_7413,N_3474,N_180);
nor U7414 (N_7414,N_576,N_909);
or U7415 (N_7415,N_1507,N_3205);
and U7416 (N_7416,N_315,N_1479);
nand U7417 (N_7417,N_2836,N_2835);
and U7418 (N_7418,N_3558,N_2104);
nor U7419 (N_7419,N_3363,N_2402);
or U7420 (N_7420,N_4696,N_3048);
nor U7421 (N_7421,N_323,N_1122);
nor U7422 (N_7422,N_1206,N_353);
or U7423 (N_7423,N_2410,N_1128);
nor U7424 (N_7424,N_59,N_4560);
nor U7425 (N_7425,N_788,N_4012);
nor U7426 (N_7426,N_4744,N_1152);
and U7427 (N_7427,N_624,N_2791);
nand U7428 (N_7428,N_237,N_513);
nand U7429 (N_7429,N_1968,N_2183);
nor U7430 (N_7430,N_2313,N_2717);
and U7431 (N_7431,N_4353,N_98);
and U7432 (N_7432,N_1251,N_1722);
nand U7433 (N_7433,N_3938,N_2052);
and U7434 (N_7434,N_2249,N_3613);
nand U7435 (N_7435,N_1082,N_317);
nor U7436 (N_7436,N_4308,N_4424);
or U7437 (N_7437,N_3776,N_4525);
or U7438 (N_7438,N_1510,N_838);
or U7439 (N_7439,N_1702,N_20);
or U7440 (N_7440,N_582,N_4262);
or U7441 (N_7441,N_2820,N_3327);
nor U7442 (N_7442,N_4617,N_267);
nor U7443 (N_7443,N_3895,N_1316);
nor U7444 (N_7444,N_1688,N_4580);
xnor U7445 (N_7445,N_2697,N_4335);
nand U7446 (N_7446,N_4251,N_1159);
and U7447 (N_7447,N_3213,N_96);
and U7448 (N_7448,N_2530,N_4040);
or U7449 (N_7449,N_2064,N_3358);
or U7450 (N_7450,N_2484,N_4050);
nor U7451 (N_7451,N_2071,N_1884);
and U7452 (N_7452,N_1397,N_3505);
nor U7453 (N_7453,N_300,N_2181);
or U7454 (N_7454,N_3986,N_2242);
nor U7455 (N_7455,N_90,N_3044);
and U7456 (N_7456,N_3224,N_3154);
nand U7457 (N_7457,N_3237,N_307);
and U7458 (N_7458,N_1907,N_4264);
xnor U7459 (N_7459,N_903,N_2048);
and U7460 (N_7460,N_2624,N_542);
nand U7461 (N_7461,N_3956,N_407);
and U7462 (N_7462,N_4963,N_4534);
nand U7463 (N_7463,N_1018,N_2724);
nand U7464 (N_7464,N_4809,N_2252);
and U7465 (N_7465,N_535,N_2961);
nor U7466 (N_7466,N_2028,N_1924);
and U7467 (N_7467,N_1404,N_417);
and U7468 (N_7468,N_1805,N_2434);
nand U7469 (N_7469,N_221,N_175);
nand U7470 (N_7470,N_4180,N_1840);
nand U7471 (N_7471,N_398,N_3548);
nand U7472 (N_7472,N_634,N_4640);
nand U7473 (N_7473,N_4289,N_1273);
or U7474 (N_7474,N_556,N_3568);
and U7475 (N_7475,N_618,N_438);
or U7476 (N_7476,N_3846,N_2889);
nor U7477 (N_7477,N_2855,N_3488);
and U7478 (N_7478,N_2336,N_1367);
nand U7479 (N_7479,N_3215,N_3633);
or U7480 (N_7480,N_1426,N_1548);
nor U7481 (N_7481,N_117,N_1772);
and U7482 (N_7482,N_2811,N_1253);
and U7483 (N_7483,N_4998,N_3448);
nor U7484 (N_7484,N_993,N_2307);
nand U7485 (N_7485,N_1214,N_2111);
nor U7486 (N_7486,N_1430,N_3543);
and U7487 (N_7487,N_2734,N_4056);
nor U7488 (N_7488,N_1925,N_2823);
or U7489 (N_7489,N_751,N_4396);
nand U7490 (N_7490,N_3388,N_1732);
and U7491 (N_7491,N_1966,N_2806);
and U7492 (N_7492,N_1080,N_3234);
nand U7493 (N_7493,N_1760,N_2201);
nor U7494 (N_7494,N_2669,N_1991);
nor U7495 (N_7495,N_1016,N_3805);
nor U7496 (N_7496,N_111,N_2509);
nand U7497 (N_7497,N_2755,N_4898);
and U7498 (N_7498,N_1406,N_1749);
and U7499 (N_7499,N_1448,N_2487);
nor U7500 (N_7500,N_3829,N_399);
and U7501 (N_7501,N_1471,N_3577);
nor U7502 (N_7502,N_4889,N_797);
nand U7503 (N_7503,N_2629,N_81);
or U7504 (N_7504,N_3731,N_3375);
nor U7505 (N_7505,N_663,N_1226);
nand U7506 (N_7506,N_727,N_4869);
nand U7507 (N_7507,N_1478,N_3037);
nand U7508 (N_7508,N_4402,N_762);
or U7509 (N_7509,N_4825,N_1683);
nand U7510 (N_7510,N_4878,N_3847);
or U7511 (N_7511,N_2602,N_4064);
and U7512 (N_7512,N_4282,N_3687);
or U7513 (N_7513,N_3132,N_1350);
nand U7514 (N_7514,N_1080,N_4300);
and U7515 (N_7515,N_342,N_1500);
nor U7516 (N_7516,N_1115,N_4564);
and U7517 (N_7517,N_1936,N_612);
or U7518 (N_7518,N_1134,N_2069);
and U7519 (N_7519,N_1892,N_510);
and U7520 (N_7520,N_3724,N_4193);
or U7521 (N_7521,N_1261,N_4486);
nand U7522 (N_7522,N_1751,N_831);
or U7523 (N_7523,N_1825,N_2845);
nand U7524 (N_7524,N_1595,N_3612);
nor U7525 (N_7525,N_724,N_3240);
or U7526 (N_7526,N_1945,N_3726);
or U7527 (N_7527,N_2166,N_527);
nor U7528 (N_7528,N_931,N_1746);
or U7529 (N_7529,N_2741,N_259);
or U7530 (N_7530,N_4273,N_2797);
and U7531 (N_7531,N_2105,N_2493);
or U7532 (N_7532,N_1288,N_683);
nor U7533 (N_7533,N_3730,N_2990);
and U7534 (N_7534,N_2478,N_517);
or U7535 (N_7535,N_200,N_1899);
nand U7536 (N_7536,N_1005,N_4375);
nor U7537 (N_7537,N_3642,N_2376);
and U7538 (N_7538,N_2049,N_3238);
nand U7539 (N_7539,N_1334,N_2525);
nor U7540 (N_7540,N_607,N_2040);
or U7541 (N_7541,N_1858,N_1965);
nor U7542 (N_7542,N_4811,N_4619);
nor U7543 (N_7543,N_73,N_2795);
and U7544 (N_7544,N_3135,N_4542);
or U7545 (N_7545,N_2460,N_348);
and U7546 (N_7546,N_4485,N_2078);
or U7547 (N_7547,N_2418,N_185);
nor U7548 (N_7548,N_3143,N_3000);
nand U7549 (N_7549,N_2587,N_4745);
and U7550 (N_7550,N_4052,N_2583);
and U7551 (N_7551,N_1401,N_2434);
nor U7552 (N_7552,N_1541,N_2057);
nand U7553 (N_7553,N_4060,N_2089);
nor U7554 (N_7554,N_1403,N_4366);
nand U7555 (N_7555,N_4585,N_159);
and U7556 (N_7556,N_2721,N_895);
nor U7557 (N_7557,N_1975,N_3755);
or U7558 (N_7558,N_2136,N_2876);
nand U7559 (N_7559,N_4900,N_4542);
nor U7560 (N_7560,N_1092,N_4679);
and U7561 (N_7561,N_2151,N_2673);
nand U7562 (N_7562,N_73,N_4972);
nand U7563 (N_7563,N_4276,N_3484);
nand U7564 (N_7564,N_2239,N_3770);
or U7565 (N_7565,N_887,N_3930);
nand U7566 (N_7566,N_4673,N_3249);
xnor U7567 (N_7567,N_189,N_3566);
nor U7568 (N_7568,N_3229,N_4229);
nand U7569 (N_7569,N_4052,N_1952);
nor U7570 (N_7570,N_2115,N_4593);
nor U7571 (N_7571,N_2764,N_4308);
and U7572 (N_7572,N_1399,N_1540);
and U7573 (N_7573,N_21,N_4351);
nor U7574 (N_7574,N_855,N_2679);
nor U7575 (N_7575,N_4057,N_4579);
xnor U7576 (N_7576,N_3342,N_489);
nor U7577 (N_7577,N_4784,N_3887);
nand U7578 (N_7578,N_4501,N_1047);
nand U7579 (N_7579,N_3404,N_699);
and U7580 (N_7580,N_128,N_3838);
nand U7581 (N_7581,N_4629,N_2343);
or U7582 (N_7582,N_3716,N_260);
nor U7583 (N_7583,N_1539,N_4068);
nor U7584 (N_7584,N_89,N_4402);
or U7585 (N_7585,N_4969,N_2933);
and U7586 (N_7586,N_4583,N_1732);
or U7587 (N_7587,N_294,N_3965);
and U7588 (N_7588,N_136,N_2771);
or U7589 (N_7589,N_4301,N_2805);
or U7590 (N_7590,N_155,N_1477);
and U7591 (N_7591,N_3272,N_1963);
nand U7592 (N_7592,N_603,N_690);
nand U7593 (N_7593,N_4068,N_758);
nor U7594 (N_7594,N_2523,N_4586);
and U7595 (N_7595,N_2184,N_4811);
or U7596 (N_7596,N_1128,N_2429);
or U7597 (N_7597,N_4974,N_2661);
and U7598 (N_7598,N_2244,N_1124);
or U7599 (N_7599,N_2600,N_515);
nand U7600 (N_7600,N_3125,N_120);
nor U7601 (N_7601,N_2728,N_2064);
or U7602 (N_7602,N_3127,N_4063);
nand U7603 (N_7603,N_4508,N_2226);
or U7604 (N_7604,N_2957,N_2582);
nor U7605 (N_7605,N_1622,N_2285);
and U7606 (N_7606,N_1370,N_1189);
and U7607 (N_7607,N_1438,N_4297);
or U7608 (N_7608,N_2624,N_1812);
and U7609 (N_7609,N_517,N_3777);
nor U7610 (N_7610,N_2797,N_2794);
or U7611 (N_7611,N_4853,N_902);
or U7612 (N_7612,N_3414,N_4980);
nand U7613 (N_7613,N_3477,N_3907);
nor U7614 (N_7614,N_1805,N_879);
and U7615 (N_7615,N_4307,N_4011);
and U7616 (N_7616,N_180,N_875);
and U7617 (N_7617,N_2188,N_3417);
nand U7618 (N_7618,N_3424,N_2461);
or U7619 (N_7619,N_633,N_3082);
or U7620 (N_7620,N_520,N_3127);
nand U7621 (N_7621,N_1584,N_4546);
nand U7622 (N_7622,N_2233,N_1051);
and U7623 (N_7623,N_4649,N_749);
nor U7624 (N_7624,N_4141,N_3731);
nand U7625 (N_7625,N_4492,N_1177);
nor U7626 (N_7626,N_214,N_68);
nor U7627 (N_7627,N_393,N_4729);
and U7628 (N_7628,N_404,N_4260);
and U7629 (N_7629,N_4036,N_1868);
or U7630 (N_7630,N_3460,N_1212);
nand U7631 (N_7631,N_901,N_1742);
or U7632 (N_7632,N_1500,N_401);
and U7633 (N_7633,N_3046,N_3974);
nand U7634 (N_7634,N_2310,N_3321);
nor U7635 (N_7635,N_1282,N_3563);
and U7636 (N_7636,N_2277,N_876);
and U7637 (N_7637,N_1372,N_2489);
nor U7638 (N_7638,N_2781,N_1239);
nand U7639 (N_7639,N_874,N_4019);
or U7640 (N_7640,N_144,N_2125);
or U7641 (N_7641,N_1187,N_2417);
nor U7642 (N_7642,N_4957,N_1303);
nand U7643 (N_7643,N_476,N_2804);
nor U7644 (N_7644,N_1888,N_1548);
xnor U7645 (N_7645,N_388,N_3286);
and U7646 (N_7646,N_4291,N_895);
or U7647 (N_7647,N_649,N_4559);
nand U7648 (N_7648,N_3148,N_2675);
xnor U7649 (N_7649,N_3272,N_1592);
or U7650 (N_7650,N_2807,N_4088);
or U7651 (N_7651,N_1794,N_1644);
and U7652 (N_7652,N_3272,N_2714);
nor U7653 (N_7653,N_4225,N_582);
or U7654 (N_7654,N_2639,N_4359);
nor U7655 (N_7655,N_223,N_4180);
nor U7656 (N_7656,N_3584,N_4858);
nand U7657 (N_7657,N_3141,N_4603);
and U7658 (N_7658,N_715,N_128);
nor U7659 (N_7659,N_2518,N_3697);
or U7660 (N_7660,N_2912,N_3926);
nand U7661 (N_7661,N_4931,N_2016);
and U7662 (N_7662,N_1090,N_4744);
or U7663 (N_7663,N_893,N_2792);
nor U7664 (N_7664,N_4823,N_1062);
and U7665 (N_7665,N_3631,N_350);
nand U7666 (N_7666,N_3433,N_3709);
or U7667 (N_7667,N_2023,N_4556);
and U7668 (N_7668,N_1711,N_2308);
nand U7669 (N_7669,N_3367,N_62);
nor U7670 (N_7670,N_4867,N_94);
or U7671 (N_7671,N_2761,N_4762);
and U7672 (N_7672,N_3924,N_1610);
and U7673 (N_7673,N_4116,N_4120);
nor U7674 (N_7674,N_3208,N_1985);
or U7675 (N_7675,N_2449,N_534);
nand U7676 (N_7676,N_3758,N_1787);
and U7677 (N_7677,N_4403,N_757);
or U7678 (N_7678,N_4223,N_3074);
nor U7679 (N_7679,N_3571,N_2699);
nor U7680 (N_7680,N_4128,N_136);
and U7681 (N_7681,N_1818,N_3826);
nand U7682 (N_7682,N_4861,N_3013);
and U7683 (N_7683,N_3265,N_381);
nor U7684 (N_7684,N_1063,N_2881);
nor U7685 (N_7685,N_2147,N_3945);
nand U7686 (N_7686,N_634,N_2379);
or U7687 (N_7687,N_3242,N_1026);
xor U7688 (N_7688,N_1765,N_1552);
nand U7689 (N_7689,N_3298,N_3310);
nand U7690 (N_7690,N_1264,N_2514);
nor U7691 (N_7691,N_2600,N_4880);
and U7692 (N_7692,N_2721,N_1359);
nand U7693 (N_7693,N_1555,N_1022);
nand U7694 (N_7694,N_3431,N_3600);
or U7695 (N_7695,N_2159,N_2766);
or U7696 (N_7696,N_734,N_4811);
nor U7697 (N_7697,N_402,N_2378);
and U7698 (N_7698,N_1545,N_1476);
and U7699 (N_7699,N_3765,N_4994);
nand U7700 (N_7700,N_550,N_3184);
xnor U7701 (N_7701,N_3725,N_729);
nand U7702 (N_7702,N_4297,N_4108);
nand U7703 (N_7703,N_928,N_2844);
and U7704 (N_7704,N_517,N_599);
nor U7705 (N_7705,N_2146,N_852);
nand U7706 (N_7706,N_4275,N_4221);
or U7707 (N_7707,N_706,N_2095);
nand U7708 (N_7708,N_1125,N_3924);
nand U7709 (N_7709,N_1848,N_3982);
or U7710 (N_7710,N_963,N_1112);
nor U7711 (N_7711,N_4294,N_556);
or U7712 (N_7712,N_536,N_4004);
and U7713 (N_7713,N_4100,N_22);
and U7714 (N_7714,N_626,N_4159);
nor U7715 (N_7715,N_4802,N_2979);
and U7716 (N_7716,N_2283,N_4421);
and U7717 (N_7717,N_3591,N_873);
nor U7718 (N_7718,N_2304,N_4135);
or U7719 (N_7719,N_3634,N_1934);
or U7720 (N_7720,N_4652,N_1403);
nand U7721 (N_7721,N_3899,N_4543);
xor U7722 (N_7722,N_4057,N_2584);
nor U7723 (N_7723,N_723,N_4916);
or U7724 (N_7724,N_4926,N_2240);
or U7725 (N_7725,N_3235,N_4556);
and U7726 (N_7726,N_161,N_2186);
nor U7727 (N_7727,N_2249,N_4339);
nand U7728 (N_7728,N_1079,N_4625);
nor U7729 (N_7729,N_2001,N_4802);
or U7730 (N_7730,N_2542,N_4240);
nand U7731 (N_7731,N_2529,N_1689);
nand U7732 (N_7732,N_353,N_2302);
nand U7733 (N_7733,N_301,N_344);
nand U7734 (N_7734,N_2289,N_1088);
and U7735 (N_7735,N_3289,N_1922);
nor U7736 (N_7736,N_294,N_4583);
or U7737 (N_7737,N_1021,N_3431);
or U7738 (N_7738,N_3408,N_2806);
nor U7739 (N_7739,N_4939,N_2129);
nor U7740 (N_7740,N_3233,N_4810);
and U7741 (N_7741,N_193,N_524);
or U7742 (N_7742,N_2732,N_1991);
or U7743 (N_7743,N_1940,N_2187);
nor U7744 (N_7744,N_733,N_3717);
or U7745 (N_7745,N_996,N_4947);
or U7746 (N_7746,N_175,N_530);
or U7747 (N_7747,N_2623,N_396);
nand U7748 (N_7748,N_2067,N_4663);
nand U7749 (N_7749,N_2297,N_225);
or U7750 (N_7750,N_4583,N_42);
nand U7751 (N_7751,N_3490,N_1959);
and U7752 (N_7752,N_3747,N_78);
or U7753 (N_7753,N_345,N_772);
or U7754 (N_7754,N_3590,N_3595);
or U7755 (N_7755,N_3961,N_3714);
or U7756 (N_7756,N_594,N_1070);
nand U7757 (N_7757,N_37,N_1191);
and U7758 (N_7758,N_3306,N_4042);
and U7759 (N_7759,N_631,N_156);
nand U7760 (N_7760,N_2576,N_899);
nand U7761 (N_7761,N_3230,N_522);
or U7762 (N_7762,N_4337,N_1048);
or U7763 (N_7763,N_67,N_4487);
nor U7764 (N_7764,N_2192,N_1646);
nor U7765 (N_7765,N_68,N_2436);
and U7766 (N_7766,N_834,N_3799);
nand U7767 (N_7767,N_1453,N_1162);
nand U7768 (N_7768,N_780,N_887);
nor U7769 (N_7769,N_2717,N_760);
nor U7770 (N_7770,N_2432,N_1768);
or U7771 (N_7771,N_221,N_551);
nor U7772 (N_7772,N_2814,N_2291);
and U7773 (N_7773,N_1402,N_898);
and U7774 (N_7774,N_1822,N_2142);
or U7775 (N_7775,N_1634,N_1300);
nor U7776 (N_7776,N_3843,N_1071);
or U7777 (N_7777,N_91,N_3304);
or U7778 (N_7778,N_3046,N_4139);
or U7779 (N_7779,N_2308,N_1691);
nor U7780 (N_7780,N_2722,N_356);
and U7781 (N_7781,N_3138,N_1582);
nor U7782 (N_7782,N_3271,N_612);
nor U7783 (N_7783,N_4920,N_2880);
nand U7784 (N_7784,N_3090,N_3290);
and U7785 (N_7785,N_1996,N_3340);
or U7786 (N_7786,N_3087,N_4339);
nand U7787 (N_7787,N_277,N_1398);
nor U7788 (N_7788,N_4782,N_1586);
nand U7789 (N_7789,N_1209,N_793);
or U7790 (N_7790,N_1317,N_3020);
nor U7791 (N_7791,N_1917,N_3625);
or U7792 (N_7792,N_1306,N_3301);
nand U7793 (N_7793,N_3145,N_1458);
nand U7794 (N_7794,N_4842,N_878);
nand U7795 (N_7795,N_1458,N_4599);
nor U7796 (N_7796,N_3987,N_888);
or U7797 (N_7797,N_3146,N_4834);
nor U7798 (N_7798,N_1889,N_3178);
or U7799 (N_7799,N_1351,N_1665);
nand U7800 (N_7800,N_3100,N_676);
nand U7801 (N_7801,N_3245,N_3949);
nand U7802 (N_7802,N_4046,N_1969);
nand U7803 (N_7803,N_4928,N_4694);
nor U7804 (N_7804,N_2931,N_2674);
nor U7805 (N_7805,N_320,N_4837);
or U7806 (N_7806,N_1878,N_946);
nor U7807 (N_7807,N_4106,N_4182);
nor U7808 (N_7808,N_865,N_4442);
and U7809 (N_7809,N_3068,N_485);
and U7810 (N_7810,N_1641,N_1391);
and U7811 (N_7811,N_4436,N_2298);
and U7812 (N_7812,N_585,N_4013);
nor U7813 (N_7813,N_220,N_923);
or U7814 (N_7814,N_1543,N_4455);
nand U7815 (N_7815,N_2754,N_3998);
nand U7816 (N_7816,N_2251,N_2511);
and U7817 (N_7817,N_2299,N_460);
nand U7818 (N_7818,N_1110,N_3332);
nor U7819 (N_7819,N_1426,N_501);
nand U7820 (N_7820,N_4720,N_2276);
nand U7821 (N_7821,N_2294,N_436);
nor U7822 (N_7822,N_326,N_1366);
nor U7823 (N_7823,N_1384,N_4777);
nor U7824 (N_7824,N_960,N_1198);
and U7825 (N_7825,N_169,N_3943);
and U7826 (N_7826,N_1130,N_476);
and U7827 (N_7827,N_3471,N_299);
nand U7828 (N_7828,N_4239,N_1961);
or U7829 (N_7829,N_2158,N_2264);
nand U7830 (N_7830,N_2590,N_673);
or U7831 (N_7831,N_1636,N_3024);
nor U7832 (N_7832,N_2678,N_3765);
or U7833 (N_7833,N_1356,N_2411);
nand U7834 (N_7834,N_4281,N_4205);
and U7835 (N_7835,N_3572,N_228);
nor U7836 (N_7836,N_3803,N_3074);
nor U7837 (N_7837,N_2368,N_2214);
nand U7838 (N_7838,N_4977,N_4250);
and U7839 (N_7839,N_2659,N_3880);
nand U7840 (N_7840,N_3827,N_3581);
nand U7841 (N_7841,N_1373,N_1668);
and U7842 (N_7842,N_3607,N_2583);
nand U7843 (N_7843,N_4310,N_947);
nand U7844 (N_7844,N_3304,N_2795);
nand U7845 (N_7845,N_4019,N_4399);
or U7846 (N_7846,N_484,N_3482);
or U7847 (N_7847,N_1784,N_4182);
nor U7848 (N_7848,N_1791,N_4064);
nor U7849 (N_7849,N_3045,N_3895);
and U7850 (N_7850,N_1343,N_2522);
and U7851 (N_7851,N_9,N_3318);
or U7852 (N_7852,N_60,N_331);
and U7853 (N_7853,N_955,N_2656);
and U7854 (N_7854,N_483,N_1164);
or U7855 (N_7855,N_669,N_2459);
and U7856 (N_7856,N_630,N_3757);
or U7857 (N_7857,N_3201,N_3786);
nor U7858 (N_7858,N_4076,N_3313);
nor U7859 (N_7859,N_2400,N_3487);
and U7860 (N_7860,N_397,N_4677);
and U7861 (N_7861,N_2742,N_2706);
and U7862 (N_7862,N_4073,N_997);
nor U7863 (N_7863,N_3400,N_892);
nor U7864 (N_7864,N_651,N_3241);
or U7865 (N_7865,N_3204,N_1836);
nand U7866 (N_7866,N_2113,N_856);
nor U7867 (N_7867,N_4099,N_1211);
nand U7868 (N_7868,N_3780,N_2430);
nand U7869 (N_7869,N_4952,N_2928);
and U7870 (N_7870,N_40,N_1457);
nand U7871 (N_7871,N_3220,N_122);
or U7872 (N_7872,N_2304,N_2021);
and U7873 (N_7873,N_84,N_1026);
nand U7874 (N_7874,N_612,N_2420);
nor U7875 (N_7875,N_1322,N_3129);
nor U7876 (N_7876,N_3057,N_2147);
nand U7877 (N_7877,N_1410,N_4889);
xnor U7878 (N_7878,N_2189,N_741);
nand U7879 (N_7879,N_261,N_609);
xor U7880 (N_7880,N_2167,N_1657);
nand U7881 (N_7881,N_4092,N_4165);
and U7882 (N_7882,N_3813,N_1488);
and U7883 (N_7883,N_199,N_3485);
nand U7884 (N_7884,N_2383,N_4601);
or U7885 (N_7885,N_1192,N_3690);
nand U7886 (N_7886,N_2943,N_1797);
nor U7887 (N_7887,N_4230,N_3677);
nand U7888 (N_7888,N_1802,N_1822);
nor U7889 (N_7889,N_3133,N_498);
nand U7890 (N_7890,N_322,N_942);
xnor U7891 (N_7891,N_387,N_202);
and U7892 (N_7892,N_3833,N_4334);
and U7893 (N_7893,N_3360,N_3825);
and U7894 (N_7894,N_2149,N_1429);
and U7895 (N_7895,N_3674,N_571);
or U7896 (N_7896,N_3902,N_2900);
nor U7897 (N_7897,N_205,N_1371);
nand U7898 (N_7898,N_4138,N_658);
nand U7899 (N_7899,N_854,N_1084);
nor U7900 (N_7900,N_4737,N_1585);
and U7901 (N_7901,N_1634,N_4848);
and U7902 (N_7902,N_3758,N_3244);
nand U7903 (N_7903,N_2997,N_1116);
nor U7904 (N_7904,N_715,N_2518);
nand U7905 (N_7905,N_2519,N_4790);
nor U7906 (N_7906,N_4173,N_783);
and U7907 (N_7907,N_3048,N_767);
nor U7908 (N_7908,N_2006,N_628);
and U7909 (N_7909,N_413,N_4244);
xor U7910 (N_7910,N_125,N_719);
nand U7911 (N_7911,N_3425,N_1534);
nand U7912 (N_7912,N_752,N_4251);
and U7913 (N_7913,N_4307,N_4903);
and U7914 (N_7914,N_3392,N_4408);
nand U7915 (N_7915,N_4659,N_4097);
or U7916 (N_7916,N_207,N_2603);
nand U7917 (N_7917,N_3622,N_1800);
and U7918 (N_7918,N_298,N_4589);
nand U7919 (N_7919,N_794,N_1034);
and U7920 (N_7920,N_4881,N_2233);
or U7921 (N_7921,N_298,N_4825);
nand U7922 (N_7922,N_2390,N_4373);
and U7923 (N_7923,N_2597,N_981);
and U7924 (N_7924,N_1764,N_341);
nor U7925 (N_7925,N_1349,N_226);
and U7926 (N_7926,N_4503,N_2056);
or U7927 (N_7927,N_4147,N_4564);
and U7928 (N_7928,N_581,N_211);
nor U7929 (N_7929,N_2240,N_2919);
nor U7930 (N_7930,N_4100,N_2484);
and U7931 (N_7931,N_4901,N_58);
nor U7932 (N_7932,N_22,N_2056);
or U7933 (N_7933,N_4913,N_1303);
nor U7934 (N_7934,N_464,N_4636);
nand U7935 (N_7935,N_3808,N_1207);
or U7936 (N_7936,N_2157,N_199);
nor U7937 (N_7937,N_809,N_1124);
xor U7938 (N_7938,N_2677,N_1875);
nor U7939 (N_7939,N_3765,N_2858);
or U7940 (N_7940,N_2254,N_4916);
nor U7941 (N_7941,N_337,N_1456);
nor U7942 (N_7942,N_1264,N_1716);
or U7943 (N_7943,N_792,N_2306);
nand U7944 (N_7944,N_4221,N_1449);
or U7945 (N_7945,N_4787,N_4845);
and U7946 (N_7946,N_4005,N_2166);
or U7947 (N_7947,N_632,N_1708);
and U7948 (N_7948,N_3406,N_4402);
and U7949 (N_7949,N_1974,N_2338);
or U7950 (N_7950,N_4500,N_1062);
nand U7951 (N_7951,N_4012,N_3130);
nand U7952 (N_7952,N_3777,N_3212);
and U7953 (N_7953,N_753,N_2221);
nand U7954 (N_7954,N_1931,N_1606);
or U7955 (N_7955,N_1323,N_2613);
or U7956 (N_7956,N_3826,N_3040);
nor U7957 (N_7957,N_2865,N_1412);
and U7958 (N_7958,N_157,N_2587);
and U7959 (N_7959,N_106,N_569);
nand U7960 (N_7960,N_711,N_330);
nor U7961 (N_7961,N_1934,N_902);
nand U7962 (N_7962,N_2565,N_1259);
or U7963 (N_7963,N_3662,N_2325);
or U7964 (N_7964,N_1437,N_3386);
nand U7965 (N_7965,N_4504,N_2543);
and U7966 (N_7966,N_331,N_4443);
and U7967 (N_7967,N_4823,N_2283);
or U7968 (N_7968,N_2959,N_2441);
nor U7969 (N_7969,N_3229,N_3044);
nor U7970 (N_7970,N_4771,N_4330);
nor U7971 (N_7971,N_2773,N_2449);
nor U7972 (N_7972,N_453,N_4501);
nand U7973 (N_7973,N_3831,N_2795);
nor U7974 (N_7974,N_3199,N_1508);
nand U7975 (N_7975,N_321,N_345);
nor U7976 (N_7976,N_659,N_626);
nand U7977 (N_7977,N_2573,N_1346);
nor U7978 (N_7978,N_3403,N_3173);
nand U7979 (N_7979,N_398,N_3249);
nand U7980 (N_7980,N_782,N_317);
and U7981 (N_7981,N_2262,N_4512);
or U7982 (N_7982,N_4827,N_4202);
nor U7983 (N_7983,N_2241,N_1157);
or U7984 (N_7984,N_334,N_2569);
and U7985 (N_7985,N_2721,N_964);
nor U7986 (N_7986,N_128,N_292);
nor U7987 (N_7987,N_3110,N_861);
or U7988 (N_7988,N_3063,N_3683);
and U7989 (N_7989,N_1958,N_4016);
or U7990 (N_7990,N_1813,N_581);
and U7991 (N_7991,N_2411,N_4384);
or U7992 (N_7992,N_2673,N_881);
nor U7993 (N_7993,N_530,N_1642);
and U7994 (N_7994,N_1836,N_4113);
and U7995 (N_7995,N_4296,N_4999);
nand U7996 (N_7996,N_1917,N_2742);
or U7997 (N_7997,N_2850,N_2961);
nor U7998 (N_7998,N_3106,N_2819);
nand U7999 (N_7999,N_2463,N_4377);
and U8000 (N_8000,N_4360,N_3582);
and U8001 (N_8001,N_3857,N_3352);
nor U8002 (N_8002,N_230,N_4411);
and U8003 (N_8003,N_4139,N_743);
nor U8004 (N_8004,N_193,N_3500);
or U8005 (N_8005,N_345,N_3236);
nand U8006 (N_8006,N_1961,N_2255);
nor U8007 (N_8007,N_4858,N_4519);
nand U8008 (N_8008,N_1247,N_2908);
and U8009 (N_8009,N_1081,N_2439);
nor U8010 (N_8010,N_546,N_2758);
nand U8011 (N_8011,N_2625,N_4768);
nand U8012 (N_8012,N_812,N_2312);
nand U8013 (N_8013,N_615,N_3575);
nor U8014 (N_8014,N_2389,N_3528);
or U8015 (N_8015,N_1767,N_3473);
or U8016 (N_8016,N_4114,N_3925);
nor U8017 (N_8017,N_211,N_1454);
and U8018 (N_8018,N_2918,N_366);
nand U8019 (N_8019,N_469,N_1189);
nand U8020 (N_8020,N_1252,N_4798);
nor U8021 (N_8021,N_1518,N_4618);
nand U8022 (N_8022,N_1203,N_2584);
nor U8023 (N_8023,N_4690,N_3720);
or U8024 (N_8024,N_4678,N_802);
nand U8025 (N_8025,N_3259,N_2328);
and U8026 (N_8026,N_881,N_3028);
nor U8027 (N_8027,N_3868,N_1448);
nor U8028 (N_8028,N_2377,N_4342);
and U8029 (N_8029,N_4636,N_4365);
and U8030 (N_8030,N_1173,N_1160);
or U8031 (N_8031,N_4228,N_2010);
nor U8032 (N_8032,N_1358,N_1907);
or U8033 (N_8033,N_495,N_4830);
nor U8034 (N_8034,N_3950,N_4252);
and U8035 (N_8035,N_2613,N_49);
nand U8036 (N_8036,N_3238,N_2331);
and U8037 (N_8037,N_2465,N_4798);
nand U8038 (N_8038,N_2849,N_2872);
or U8039 (N_8039,N_3475,N_1437);
nand U8040 (N_8040,N_3186,N_3756);
and U8041 (N_8041,N_1181,N_4176);
nand U8042 (N_8042,N_439,N_4767);
or U8043 (N_8043,N_1465,N_4930);
or U8044 (N_8044,N_4472,N_4412);
or U8045 (N_8045,N_1924,N_3496);
and U8046 (N_8046,N_669,N_3392);
nand U8047 (N_8047,N_650,N_2930);
or U8048 (N_8048,N_4922,N_4854);
nor U8049 (N_8049,N_4150,N_4474);
nand U8050 (N_8050,N_1682,N_2768);
and U8051 (N_8051,N_624,N_1480);
nand U8052 (N_8052,N_1158,N_4979);
or U8053 (N_8053,N_3398,N_3689);
or U8054 (N_8054,N_2585,N_1189);
or U8055 (N_8055,N_514,N_3870);
and U8056 (N_8056,N_1770,N_4271);
or U8057 (N_8057,N_459,N_566);
and U8058 (N_8058,N_3343,N_1761);
nor U8059 (N_8059,N_1115,N_3021);
nor U8060 (N_8060,N_30,N_4695);
nand U8061 (N_8061,N_1556,N_4857);
and U8062 (N_8062,N_4387,N_61);
or U8063 (N_8063,N_4401,N_601);
nor U8064 (N_8064,N_1936,N_2022);
or U8065 (N_8065,N_3869,N_4749);
nand U8066 (N_8066,N_1598,N_3836);
nor U8067 (N_8067,N_90,N_49);
nor U8068 (N_8068,N_1185,N_669);
nor U8069 (N_8069,N_3448,N_4493);
and U8070 (N_8070,N_901,N_1491);
nand U8071 (N_8071,N_3085,N_2626);
xnor U8072 (N_8072,N_2767,N_1973);
nand U8073 (N_8073,N_1519,N_2855);
nor U8074 (N_8074,N_1314,N_1949);
nor U8075 (N_8075,N_2626,N_3422);
nor U8076 (N_8076,N_2552,N_2536);
nand U8077 (N_8077,N_4709,N_1671);
and U8078 (N_8078,N_2466,N_3864);
nor U8079 (N_8079,N_3449,N_1699);
or U8080 (N_8080,N_2641,N_4430);
nor U8081 (N_8081,N_4549,N_4665);
nand U8082 (N_8082,N_4907,N_2781);
nor U8083 (N_8083,N_2344,N_2747);
nand U8084 (N_8084,N_1231,N_4717);
nand U8085 (N_8085,N_1212,N_3470);
nor U8086 (N_8086,N_3556,N_457);
nand U8087 (N_8087,N_664,N_1626);
nor U8088 (N_8088,N_1335,N_1359);
and U8089 (N_8089,N_4474,N_4117);
nor U8090 (N_8090,N_2971,N_2698);
and U8091 (N_8091,N_4480,N_4973);
nor U8092 (N_8092,N_308,N_346);
or U8093 (N_8093,N_1893,N_3222);
nor U8094 (N_8094,N_28,N_475);
nand U8095 (N_8095,N_1746,N_2087);
nor U8096 (N_8096,N_1804,N_3342);
nor U8097 (N_8097,N_3504,N_3721);
or U8098 (N_8098,N_344,N_1910);
or U8099 (N_8099,N_4822,N_2784);
nor U8100 (N_8100,N_752,N_2958);
and U8101 (N_8101,N_4294,N_694);
or U8102 (N_8102,N_2066,N_3955);
nor U8103 (N_8103,N_2838,N_1038);
nand U8104 (N_8104,N_2632,N_2504);
or U8105 (N_8105,N_2129,N_2982);
or U8106 (N_8106,N_2987,N_2616);
and U8107 (N_8107,N_9,N_1478);
and U8108 (N_8108,N_3309,N_3866);
nor U8109 (N_8109,N_166,N_3553);
nor U8110 (N_8110,N_521,N_3411);
or U8111 (N_8111,N_2453,N_3101);
nand U8112 (N_8112,N_3686,N_1268);
or U8113 (N_8113,N_3158,N_646);
and U8114 (N_8114,N_1613,N_3503);
and U8115 (N_8115,N_2322,N_4192);
nand U8116 (N_8116,N_3306,N_1616);
or U8117 (N_8117,N_4774,N_4996);
or U8118 (N_8118,N_4697,N_3500);
or U8119 (N_8119,N_3574,N_2621);
nor U8120 (N_8120,N_3359,N_1048);
or U8121 (N_8121,N_4730,N_3323);
nand U8122 (N_8122,N_4397,N_2509);
or U8123 (N_8123,N_1296,N_3399);
or U8124 (N_8124,N_1371,N_3915);
and U8125 (N_8125,N_1686,N_1568);
and U8126 (N_8126,N_3343,N_1728);
nand U8127 (N_8127,N_212,N_1440);
nor U8128 (N_8128,N_115,N_1605);
nor U8129 (N_8129,N_3534,N_2292);
and U8130 (N_8130,N_2404,N_4131);
or U8131 (N_8131,N_4000,N_2498);
or U8132 (N_8132,N_2742,N_1559);
nand U8133 (N_8133,N_424,N_3393);
nand U8134 (N_8134,N_3683,N_1694);
or U8135 (N_8135,N_368,N_4908);
or U8136 (N_8136,N_426,N_1629);
and U8137 (N_8137,N_4126,N_3961);
nor U8138 (N_8138,N_866,N_643);
nor U8139 (N_8139,N_949,N_4516);
nand U8140 (N_8140,N_3435,N_4512);
nand U8141 (N_8141,N_2342,N_2563);
nor U8142 (N_8142,N_2953,N_4573);
nand U8143 (N_8143,N_2952,N_4303);
and U8144 (N_8144,N_4735,N_433);
nand U8145 (N_8145,N_4287,N_2147);
xnor U8146 (N_8146,N_2530,N_3756);
nor U8147 (N_8147,N_4436,N_4258);
and U8148 (N_8148,N_3560,N_414);
nor U8149 (N_8149,N_1993,N_4493);
nand U8150 (N_8150,N_2227,N_4672);
or U8151 (N_8151,N_1436,N_4374);
nor U8152 (N_8152,N_522,N_1656);
nand U8153 (N_8153,N_1464,N_2555);
nor U8154 (N_8154,N_2837,N_965);
nor U8155 (N_8155,N_4244,N_343);
nor U8156 (N_8156,N_1064,N_4014);
or U8157 (N_8157,N_67,N_2646);
and U8158 (N_8158,N_533,N_3654);
nand U8159 (N_8159,N_41,N_3642);
nand U8160 (N_8160,N_3872,N_3092);
nor U8161 (N_8161,N_4707,N_201);
nor U8162 (N_8162,N_2857,N_219);
or U8163 (N_8163,N_3482,N_4460);
nand U8164 (N_8164,N_96,N_2378);
nand U8165 (N_8165,N_1984,N_3728);
nand U8166 (N_8166,N_4954,N_1793);
and U8167 (N_8167,N_4296,N_1493);
nand U8168 (N_8168,N_2390,N_545);
nand U8169 (N_8169,N_2040,N_3074);
or U8170 (N_8170,N_2269,N_3726);
nor U8171 (N_8171,N_2854,N_2409);
or U8172 (N_8172,N_3321,N_4997);
or U8173 (N_8173,N_979,N_2140);
and U8174 (N_8174,N_3798,N_3796);
and U8175 (N_8175,N_559,N_4163);
or U8176 (N_8176,N_4602,N_1781);
nor U8177 (N_8177,N_3810,N_4745);
nor U8178 (N_8178,N_307,N_2882);
nand U8179 (N_8179,N_1330,N_1433);
and U8180 (N_8180,N_924,N_2542);
xor U8181 (N_8181,N_3855,N_4266);
or U8182 (N_8182,N_860,N_3909);
or U8183 (N_8183,N_286,N_3465);
nand U8184 (N_8184,N_2129,N_2719);
and U8185 (N_8185,N_24,N_239);
or U8186 (N_8186,N_788,N_2648);
nor U8187 (N_8187,N_1380,N_4904);
and U8188 (N_8188,N_2461,N_1983);
and U8189 (N_8189,N_1719,N_3966);
xnor U8190 (N_8190,N_2341,N_1532);
nor U8191 (N_8191,N_699,N_856);
nor U8192 (N_8192,N_4344,N_3698);
or U8193 (N_8193,N_1063,N_2039);
or U8194 (N_8194,N_1393,N_2736);
and U8195 (N_8195,N_3922,N_1476);
or U8196 (N_8196,N_1752,N_1771);
and U8197 (N_8197,N_14,N_399);
xor U8198 (N_8198,N_3252,N_4013);
nand U8199 (N_8199,N_1707,N_2608);
nand U8200 (N_8200,N_4325,N_1741);
nand U8201 (N_8201,N_3894,N_3136);
or U8202 (N_8202,N_224,N_3495);
and U8203 (N_8203,N_4508,N_1327);
nor U8204 (N_8204,N_1664,N_4874);
or U8205 (N_8205,N_4276,N_3162);
nor U8206 (N_8206,N_3052,N_1718);
xor U8207 (N_8207,N_3076,N_3216);
nand U8208 (N_8208,N_937,N_3142);
nor U8209 (N_8209,N_40,N_2521);
and U8210 (N_8210,N_1382,N_4184);
or U8211 (N_8211,N_2970,N_2441);
nand U8212 (N_8212,N_4232,N_3962);
nor U8213 (N_8213,N_4627,N_2324);
or U8214 (N_8214,N_1280,N_2010);
or U8215 (N_8215,N_3645,N_1639);
or U8216 (N_8216,N_2468,N_2460);
or U8217 (N_8217,N_384,N_1232);
nor U8218 (N_8218,N_2482,N_3759);
or U8219 (N_8219,N_2075,N_761);
nor U8220 (N_8220,N_1496,N_2709);
or U8221 (N_8221,N_3602,N_1651);
or U8222 (N_8222,N_2886,N_4366);
nor U8223 (N_8223,N_1681,N_2285);
and U8224 (N_8224,N_140,N_265);
nand U8225 (N_8225,N_4544,N_946);
nand U8226 (N_8226,N_1656,N_3976);
or U8227 (N_8227,N_3655,N_1070);
and U8228 (N_8228,N_2572,N_2722);
or U8229 (N_8229,N_2128,N_2851);
or U8230 (N_8230,N_2328,N_3831);
nor U8231 (N_8231,N_1819,N_985);
and U8232 (N_8232,N_664,N_2800);
nor U8233 (N_8233,N_1709,N_213);
nor U8234 (N_8234,N_878,N_3442);
nor U8235 (N_8235,N_2187,N_110);
nand U8236 (N_8236,N_4838,N_272);
nor U8237 (N_8237,N_3269,N_3637);
nand U8238 (N_8238,N_1736,N_2845);
or U8239 (N_8239,N_72,N_3657);
or U8240 (N_8240,N_3088,N_1508);
nand U8241 (N_8241,N_2210,N_4096);
nor U8242 (N_8242,N_4887,N_1296);
nor U8243 (N_8243,N_3204,N_4371);
or U8244 (N_8244,N_55,N_417);
or U8245 (N_8245,N_3350,N_3883);
or U8246 (N_8246,N_2979,N_3170);
and U8247 (N_8247,N_4853,N_4576);
nand U8248 (N_8248,N_2615,N_4586);
nand U8249 (N_8249,N_3670,N_2259);
nor U8250 (N_8250,N_1133,N_469);
and U8251 (N_8251,N_4928,N_1849);
nand U8252 (N_8252,N_3102,N_391);
and U8253 (N_8253,N_278,N_4190);
nand U8254 (N_8254,N_2746,N_4553);
nor U8255 (N_8255,N_2456,N_2073);
and U8256 (N_8256,N_3615,N_1092);
nor U8257 (N_8257,N_4411,N_2259);
nand U8258 (N_8258,N_2845,N_1197);
nor U8259 (N_8259,N_4690,N_1868);
or U8260 (N_8260,N_1670,N_3279);
nor U8261 (N_8261,N_1441,N_1086);
nand U8262 (N_8262,N_4381,N_3585);
or U8263 (N_8263,N_4123,N_3005);
or U8264 (N_8264,N_1787,N_1347);
nand U8265 (N_8265,N_2636,N_2203);
nor U8266 (N_8266,N_4839,N_2522);
nand U8267 (N_8267,N_1130,N_4693);
and U8268 (N_8268,N_1142,N_4752);
and U8269 (N_8269,N_1940,N_2688);
nand U8270 (N_8270,N_3192,N_401);
nor U8271 (N_8271,N_1763,N_2336);
and U8272 (N_8272,N_2520,N_622);
nand U8273 (N_8273,N_1207,N_4778);
and U8274 (N_8274,N_361,N_1724);
or U8275 (N_8275,N_4375,N_995);
and U8276 (N_8276,N_3970,N_4595);
or U8277 (N_8277,N_2868,N_2735);
nand U8278 (N_8278,N_4360,N_182);
nor U8279 (N_8279,N_2881,N_384);
nand U8280 (N_8280,N_1741,N_1543);
or U8281 (N_8281,N_2484,N_1169);
xnor U8282 (N_8282,N_2178,N_3034);
nand U8283 (N_8283,N_3152,N_1163);
nor U8284 (N_8284,N_3969,N_1810);
nand U8285 (N_8285,N_4465,N_4023);
or U8286 (N_8286,N_482,N_186);
nor U8287 (N_8287,N_364,N_2470);
nand U8288 (N_8288,N_1751,N_2366);
and U8289 (N_8289,N_1276,N_2699);
and U8290 (N_8290,N_2819,N_1022);
or U8291 (N_8291,N_3767,N_1064);
and U8292 (N_8292,N_1446,N_1986);
nor U8293 (N_8293,N_1616,N_1560);
nand U8294 (N_8294,N_1431,N_2289);
or U8295 (N_8295,N_923,N_1043);
nor U8296 (N_8296,N_2356,N_768);
or U8297 (N_8297,N_4683,N_4245);
nor U8298 (N_8298,N_1513,N_531);
or U8299 (N_8299,N_2314,N_3795);
nand U8300 (N_8300,N_2622,N_4207);
and U8301 (N_8301,N_2422,N_3364);
nand U8302 (N_8302,N_2640,N_1685);
nor U8303 (N_8303,N_4759,N_2570);
nand U8304 (N_8304,N_2518,N_3839);
nand U8305 (N_8305,N_3727,N_3733);
and U8306 (N_8306,N_3407,N_317);
nand U8307 (N_8307,N_2704,N_929);
or U8308 (N_8308,N_2253,N_1084);
nand U8309 (N_8309,N_2556,N_1474);
and U8310 (N_8310,N_85,N_797);
nor U8311 (N_8311,N_3174,N_3600);
nor U8312 (N_8312,N_3873,N_1737);
nor U8313 (N_8313,N_2443,N_3019);
nor U8314 (N_8314,N_2561,N_3315);
and U8315 (N_8315,N_170,N_1362);
nand U8316 (N_8316,N_2701,N_4428);
and U8317 (N_8317,N_2813,N_3523);
nand U8318 (N_8318,N_4601,N_4469);
nor U8319 (N_8319,N_4128,N_376);
nand U8320 (N_8320,N_2619,N_288);
nor U8321 (N_8321,N_1003,N_1006);
and U8322 (N_8322,N_3545,N_1943);
and U8323 (N_8323,N_3262,N_4788);
nor U8324 (N_8324,N_4369,N_3700);
and U8325 (N_8325,N_1946,N_3738);
or U8326 (N_8326,N_4537,N_4038);
or U8327 (N_8327,N_3178,N_3792);
nor U8328 (N_8328,N_3788,N_2594);
nand U8329 (N_8329,N_3078,N_1402);
nand U8330 (N_8330,N_4288,N_51);
nor U8331 (N_8331,N_1020,N_4133);
nand U8332 (N_8332,N_957,N_362);
nand U8333 (N_8333,N_1825,N_3352);
nand U8334 (N_8334,N_1645,N_1921);
or U8335 (N_8335,N_2655,N_1560);
nor U8336 (N_8336,N_4372,N_3218);
and U8337 (N_8337,N_1756,N_3060);
nor U8338 (N_8338,N_1244,N_1382);
nand U8339 (N_8339,N_4021,N_15);
or U8340 (N_8340,N_4817,N_3021);
or U8341 (N_8341,N_474,N_4378);
or U8342 (N_8342,N_3809,N_4930);
nand U8343 (N_8343,N_565,N_3229);
and U8344 (N_8344,N_4742,N_3697);
and U8345 (N_8345,N_4621,N_4928);
and U8346 (N_8346,N_3901,N_2182);
nand U8347 (N_8347,N_1334,N_4250);
nand U8348 (N_8348,N_801,N_2163);
nand U8349 (N_8349,N_4469,N_3192);
nand U8350 (N_8350,N_1636,N_1491);
nor U8351 (N_8351,N_2249,N_3297);
nor U8352 (N_8352,N_2650,N_4373);
and U8353 (N_8353,N_107,N_4349);
or U8354 (N_8354,N_1581,N_4883);
or U8355 (N_8355,N_3730,N_277);
or U8356 (N_8356,N_213,N_890);
and U8357 (N_8357,N_4123,N_4207);
and U8358 (N_8358,N_12,N_3164);
nand U8359 (N_8359,N_815,N_3267);
and U8360 (N_8360,N_3877,N_4627);
nand U8361 (N_8361,N_1160,N_3233);
nor U8362 (N_8362,N_1684,N_2858);
and U8363 (N_8363,N_734,N_4453);
nand U8364 (N_8364,N_431,N_1216);
nand U8365 (N_8365,N_1001,N_4301);
nand U8366 (N_8366,N_2296,N_1800);
or U8367 (N_8367,N_1379,N_4084);
and U8368 (N_8368,N_3551,N_3126);
or U8369 (N_8369,N_2400,N_4063);
nand U8370 (N_8370,N_2016,N_1459);
nand U8371 (N_8371,N_3131,N_193);
nor U8372 (N_8372,N_3697,N_3196);
and U8373 (N_8373,N_1223,N_961);
or U8374 (N_8374,N_1568,N_2543);
nor U8375 (N_8375,N_4866,N_794);
or U8376 (N_8376,N_268,N_4503);
or U8377 (N_8377,N_2258,N_2095);
nand U8378 (N_8378,N_2439,N_3856);
and U8379 (N_8379,N_2174,N_1712);
or U8380 (N_8380,N_1240,N_3161);
nor U8381 (N_8381,N_116,N_302);
and U8382 (N_8382,N_678,N_2943);
and U8383 (N_8383,N_944,N_3815);
nor U8384 (N_8384,N_4412,N_3938);
or U8385 (N_8385,N_3421,N_4876);
or U8386 (N_8386,N_1029,N_2681);
nand U8387 (N_8387,N_1625,N_619);
or U8388 (N_8388,N_2747,N_28);
xor U8389 (N_8389,N_3761,N_4741);
and U8390 (N_8390,N_881,N_2208);
nor U8391 (N_8391,N_2574,N_1875);
nand U8392 (N_8392,N_2385,N_2592);
nor U8393 (N_8393,N_3514,N_4204);
nand U8394 (N_8394,N_2566,N_3102);
nand U8395 (N_8395,N_1666,N_116);
nand U8396 (N_8396,N_1779,N_3008);
and U8397 (N_8397,N_1420,N_2690);
nand U8398 (N_8398,N_15,N_4037);
nand U8399 (N_8399,N_1853,N_4428);
nand U8400 (N_8400,N_929,N_4453);
nor U8401 (N_8401,N_2056,N_2991);
nor U8402 (N_8402,N_2534,N_1795);
nor U8403 (N_8403,N_471,N_1724);
nand U8404 (N_8404,N_2846,N_3337);
and U8405 (N_8405,N_3288,N_3737);
nor U8406 (N_8406,N_704,N_3595);
nor U8407 (N_8407,N_4008,N_1282);
or U8408 (N_8408,N_4167,N_1994);
and U8409 (N_8409,N_361,N_3049);
nand U8410 (N_8410,N_4605,N_4671);
or U8411 (N_8411,N_975,N_209);
nand U8412 (N_8412,N_2074,N_2451);
and U8413 (N_8413,N_2842,N_2988);
and U8414 (N_8414,N_4322,N_1431);
and U8415 (N_8415,N_3949,N_856);
nand U8416 (N_8416,N_4129,N_3357);
and U8417 (N_8417,N_3435,N_887);
and U8418 (N_8418,N_77,N_290);
nand U8419 (N_8419,N_2699,N_524);
nor U8420 (N_8420,N_2570,N_2628);
and U8421 (N_8421,N_1014,N_4100);
nor U8422 (N_8422,N_1614,N_1322);
nand U8423 (N_8423,N_604,N_879);
nand U8424 (N_8424,N_2178,N_3294);
or U8425 (N_8425,N_2971,N_3583);
nor U8426 (N_8426,N_630,N_92);
and U8427 (N_8427,N_4815,N_2390);
nor U8428 (N_8428,N_3792,N_3522);
xnor U8429 (N_8429,N_294,N_2671);
nand U8430 (N_8430,N_2665,N_1164);
and U8431 (N_8431,N_2852,N_4845);
nand U8432 (N_8432,N_3787,N_4099);
nor U8433 (N_8433,N_3963,N_2871);
or U8434 (N_8434,N_1263,N_1494);
nand U8435 (N_8435,N_1737,N_3621);
nand U8436 (N_8436,N_525,N_3167);
or U8437 (N_8437,N_1925,N_4749);
nand U8438 (N_8438,N_3958,N_4772);
and U8439 (N_8439,N_3,N_4812);
nor U8440 (N_8440,N_1686,N_3360);
and U8441 (N_8441,N_1802,N_2688);
nor U8442 (N_8442,N_832,N_488);
and U8443 (N_8443,N_4346,N_4706);
nor U8444 (N_8444,N_2280,N_1005);
nand U8445 (N_8445,N_3366,N_927);
nor U8446 (N_8446,N_334,N_1132);
or U8447 (N_8447,N_2716,N_252);
or U8448 (N_8448,N_2633,N_3891);
nor U8449 (N_8449,N_4437,N_2478);
nand U8450 (N_8450,N_4081,N_2943);
nor U8451 (N_8451,N_3398,N_2857);
nand U8452 (N_8452,N_1621,N_3891);
nor U8453 (N_8453,N_973,N_770);
or U8454 (N_8454,N_669,N_1098);
or U8455 (N_8455,N_1306,N_4298);
and U8456 (N_8456,N_1277,N_23);
nor U8457 (N_8457,N_2590,N_3985);
nor U8458 (N_8458,N_1049,N_744);
or U8459 (N_8459,N_4714,N_916);
nor U8460 (N_8460,N_103,N_900);
or U8461 (N_8461,N_2591,N_2873);
nor U8462 (N_8462,N_4474,N_3206);
or U8463 (N_8463,N_983,N_388);
nand U8464 (N_8464,N_565,N_2569);
and U8465 (N_8465,N_898,N_96);
or U8466 (N_8466,N_1519,N_1183);
nor U8467 (N_8467,N_684,N_956);
or U8468 (N_8468,N_1552,N_2620);
nand U8469 (N_8469,N_2343,N_444);
and U8470 (N_8470,N_547,N_4647);
xnor U8471 (N_8471,N_1459,N_3265);
nand U8472 (N_8472,N_3004,N_4357);
nor U8473 (N_8473,N_1271,N_21);
nor U8474 (N_8474,N_2813,N_4032);
nand U8475 (N_8475,N_919,N_4855);
nor U8476 (N_8476,N_857,N_4244);
nand U8477 (N_8477,N_1085,N_843);
and U8478 (N_8478,N_3132,N_4980);
or U8479 (N_8479,N_4139,N_1839);
nor U8480 (N_8480,N_4165,N_2198);
and U8481 (N_8481,N_3834,N_810);
or U8482 (N_8482,N_4069,N_617);
nor U8483 (N_8483,N_4234,N_1071);
nand U8484 (N_8484,N_829,N_921);
or U8485 (N_8485,N_2554,N_362);
or U8486 (N_8486,N_591,N_569);
nor U8487 (N_8487,N_3110,N_1155);
nand U8488 (N_8488,N_1789,N_1161);
and U8489 (N_8489,N_1517,N_3798);
and U8490 (N_8490,N_3771,N_3787);
nand U8491 (N_8491,N_3205,N_2364);
nor U8492 (N_8492,N_1278,N_4697);
nand U8493 (N_8493,N_754,N_4455);
nor U8494 (N_8494,N_3715,N_3268);
nor U8495 (N_8495,N_2204,N_4215);
nand U8496 (N_8496,N_2492,N_4696);
and U8497 (N_8497,N_770,N_4291);
and U8498 (N_8498,N_941,N_1372);
nand U8499 (N_8499,N_3496,N_310);
and U8500 (N_8500,N_381,N_3041);
or U8501 (N_8501,N_210,N_2118);
nor U8502 (N_8502,N_1923,N_3674);
or U8503 (N_8503,N_831,N_4870);
nor U8504 (N_8504,N_4692,N_4501);
and U8505 (N_8505,N_2609,N_4921);
and U8506 (N_8506,N_3165,N_1669);
nor U8507 (N_8507,N_3180,N_4189);
or U8508 (N_8508,N_3261,N_3370);
or U8509 (N_8509,N_1261,N_3290);
or U8510 (N_8510,N_1923,N_556);
nand U8511 (N_8511,N_4499,N_1200);
or U8512 (N_8512,N_837,N_965);
and U8513 (N_8513,N_115,N_1288);
nor U8514 (N_8514,N_8,N_3355);
nor U8515 (N_8515,N_2321,N_4105);
nand U8516 (N_8516,N_1699,N_862);
and U8517 (N_8517,N_770,N_4843);
or U8518 (N_8518,N_1956,N_546);
and U8519 (N_8519,N_254,N_2820);
nand U8520 (N_8520,N_3940,N_1956);
nand U8521 (N_8521,N_3762,N_501);
or U8522 (N_8522,N_3242,N_3676);
nor U8523 (N_8523,N_1885,N_2304);
nand U8524 (N_8524,N_3860,N_1207);
and U8525 (N_8525,N_1908,N_1529);
nor U8526 (N_8526,N_494,N_1375);
or U8527 (N_8527,N_926,N_4204);
nor U8528 (N_8528,N_3045,N_3091);
and U8529 (N_8529,N_1530,N_1519);
or U8530 (N_8530,N_311,N_4544);
or U8531 (N_8531,N_2009,N_263);
nand U8532 (N_8532,N_2313,N_2629);
and U8533 (N_8533,N_584,N_4422);
or U8534 (N_8534,N_988,N_131);
nand U8535 (N_8535,N_4176,N_4420);
and U8536 (N_8536,N_297,N_2376);
nand U8537 (N_8537,N_2119,N_1882);
and U8538 (N_8538,N_996,N_4534);
and U8539 (N_8539,N_2874,N_4326);
nand U8540 (N_8540,N_2314,N_2280);
or U8541 (N_8541,N_3953,N_1396);
and U8542 (N_8542,N_2906,N_1074);
or U8543 (N_8543,N_1447,N_1830);
and U8544 (N_8544,N_4113,N_1317);
and U8545 (N_8545,N_208,N_507);
or U8546 (N_8546,N_3587,N_4441);
nor U8547 (N_8547,N_1562,N_2966);
or U8548 (N_8548,N_632,N_627);
or U8549 (N_8549,N_4514,N_3677);
or U8550 (N_8550,N_1488,N_902);
nand U8551 (N_8551,N_1258,N_1936);
and U8552 (N_8552,N_3488,N_161);
nand U8553 (N_8553,N_2765,N_4627);
xor U8554 (N_8554,N_1050,N_3275);
nor U8555 (N_8555,N_557,N_3936);
nand U8556 (N_8556,N_3816,N_4408);
or U8557 (N_8557,N_4415,N_4325);
xor U8558 (N_8558,N_1629,N_1541);
and U8559 (N_8559,N_82,N_4401);
and U8560 (N_8560,N_3348,N_1140);
and U8561 (N_8561,N_750,N_1370);
nor U8562 (N_8562,N_2319,N_2719);
and U8563 (N_8563,N_2797,N_256);
or U8564 (N_8564,N_603,N_4179);
and U8565 (N_8565,N_4590,N_1359);
or U8566 (N_8566,N_3694,N_425);
or U8567 (N_8567,N_2961,N_2873);
and U8568 (N_8568,N_3360,N_860);
and U8569 (N_8569,N_3219,N_2025);
nor U8570 (N_8570,N_2757,N_4137);
nor U8571 (N_8571,N_3001,N_762);
nor U8572 (N_8572,N_2693,N_1925);
nor U8573 (N_8573,N_1256,N_3925);
xor U8574 (N_8574,N_541,N_4239);
nand U8575 (N_8575,N_582,N_2943);
nand U8576 (N_8576,N_736,N_1188);
nor U8577 (N_8577,N_2350,N_2282);
nor U8578 (N_8578,N_2309,N_2717);
nor U8579 (N_8579,N_2928,N_1883);
nand U8580 (N_8580,N_4460,N_4352);
and U8581 (N_8581,N_781,N_4898);
nor U8582 (N_8582,N_1488,N_4789);
nor U8583 (N_8583,N_276,N_3504);
nor U8584 (N_8584,N_2868,N_2275);
or U8585 (N_8585,N_1159,N_1182);
nand U8586 (N_8586,N_2518,N_1679);
and U8587 (N_8587,N_2792,N_3561);
xnor U8588 (N_8588,N_444,N_962);
nand U8589 (N_8589,N_164,N_2006);
or U8590 (N_8590,N_534,N_1843);
or U8591 (N_8591,N_3220,N_658);
nand U8592 (N_8592,N_3206,N_4687);
nand U8593 (N_8593,N_4134,N_981);
nor U8594 (N_8594,N_3995,N_4734);
nand U8595 (N_8595,N_3282,N_2494);
nand U8596 (N_8596,N_1249,N_3154);
nand U8597 (N_8597,N_1389,N_4395);
nand U8598 (N_8598,N_4567,N_2042);
nor U8599 (N_8599,N_3349,N_4332);
nor U8600 (N_8600,N_4585,N_4346);
nand U8601 (N_8601,N_4955,N_2864);
nor U8602 (N_8602,N_3776,N_450);
nand U8603 (N_8603,N_531,N_3919);
or U8604 (N_8604,N_3302,N_2178);
nand U8605 (N_8605,N_2446,N_1532);
xor U8606 (N_8606,N_4637,N_3742);
and U8607 (N_8607,N_4163,N_4604);
nor U8608 (N_8608,N_2296,N_4863);
nand U8609 (N_8609,N_2390,N_2447);
and U8610 (N_8610,N_3151,N_1833);
and U8611 (N_8611,N_4428,N_3216);
or U8612 (N_8612,N_3418,N_1451);
or U8613 (N_8613,N_74,N_1834);
and U8614 (N_8614,N_4183,N_947);
or U8615 (N_8615,N_945,N_1611);
nand U8616 (N_8616,N_4212,N_1922);
nand U8617 (N_8617,N_2281,N_1341);
nand U8618 (N_8618,N_2780,N_881);
or U8619 (N_8619,N_2072,N_371);
nand U8620 (N_8620,N_4787,N_3724);
or U8621 (N_8621,N_2732,N_828);
and U8622 (N_8622,N_1431,N_3120);
or U8623 (N_8623,N_1297,N_649);
or U8624 (N_8624,N_2158,N_1325);
and U8625 (N_8625,N_4938,N_2661);
or U8626 (N_8626,N_4394,N_2640);
nor U8627 (N_8627,N_4721,N_1524);
nand U8628 (N_8628,N_127,N_3959);
or U8629 (N_8629,N_1833,N_1016);
and U8630 (N_8630,N_2897,N_3524);
nand U8631 (N_8631,N_4659,N_3396);
nand U8632 (N_8632,N_3313,N_4781);
nand U8633 (N_8633,N_4053,N_870);
or U8634 (N_8634,N_1342,N_187);
and U8635 (N_8635,N_2677,N_3123);
or U8636 (N_8636,N_4885,N_612);
and U8637 (N_8637,N_4175,N_2836);
and U8638 (N_8638,N_1286,N_3361);
nand U8639 (N_8639,N_1771,N_321);
nor U8640 (N_8640,N_2865,N_2975);
nor U8641 (N_8641,N_27,N_3118);
and U8642 (N_8642,N_3546,N_2231);
and U8643 (N_8643,N_1548,N_4145);
and U8644 (N_8644,N_2702,N_4470);
or U8645 (N_8645,N_3543,N_1524);
and U8646 (N_8646,N_747,N_539);
or U8647 (N_8647,N_1122,N_2312);
nand U8648 (N_8648,N_234,N_2839);
nor U8649 (N_8649,N_4370,N_1045);
nor U8650 (N_8650,N_170,N_4278);
nor U8651 (N_8651,N_202,N_1326);
and U8652 (N_8652,N_3647,N_4501);
and U8653 (N_8653,N_3722,N_3366);
nor U8654 (N_8654,N_3053,N_945);
nor U8655 (N_8655,N_394,N_250);
and U8656 (N_8656,N_4264,N_1254);
nand U8657 (N_8657,N_910,N_441);
nand U8658 (N_8658,N_1729,N_4194);
nor U8659 (N_8659,N_1434,N_1324);
or U8660 (N_8660,N_2281,N_1527);
nor U8661 (N_8661,N_4172,N_3713);
and U8662 (N_8662,N_954,N_2746);
nand U8663 (N_8663,N_2530,N_2844);
and U8664 (N_8664,N_4931,N_2337);
nor U8665 (N_8665,N_3968,N_590);
or U8666 (N_8666,N_2198,N_1046);
nand U8667 (N_8667,N_1633,N_4572);
nor U8668 (N_8668,N_3916,N_4280);
nor U8669 (N_8669,N_4744,N_4083);
and U8670 (N_8670,N_1897,N_2913);
nor U8671 (N_8671,N_4944,N_3418);
nor U8672 (N_8672,N_2956,N_65);
nor U8673 (N_8673,N_4396,N_3514);
and U8674 (N_8674,N_1946,N_751);
or U8675 (N_8675,N_1508,N_2623);
nand U8676 (N_8676,N_3638,N_657);
or U8677 (N_8677,N_636,N_2093);
or U8678 (N_8678,N_3513,N_3036);
or U8679 (N_8679,N_662,N_2329);
nand U8680 (N_8680,N_4859,N_1056);
and U8681 (N_8681,N_3675,N_1177);
nand U8682 (N_8682,N_1503,N_4223);
nand U8683 (N_8683,N_1943,N_1001);
nor U8684 (N_8684,N_3448,N_1397);
and U8685 (N_8685,N_1234,N_4667);
or U8686 (N_8686,N_1081,N_2938);
or U8687 (N_8687,N_2252,N_1328);
nor U8688 (N_8688,N_510,N_0);
nor U8689 (N_8689,N_3396,N_4123);
and U8690 (N_8690,N_1759,N_1069);
or U8691 (N_8691,N_2067,N_2782);
nand U8692 (N_8692,N_2322,N_2662);
nor U8693 (N_8693,N_3189,N_2153);
and U8694 (N_8694,N_3326,N_1143);
nand U8695 (N_8695,N_1173,N_570);
nor U8696 (N_8696,N_1752,N_873);
nor U8697 (N_8697,N_3865,N_1883);
and U8698 (N_8698,N_4860,N_4619);
nor U8699 (N_8699,N_3051,N_3788);
or U8700 (N_8700,N_2772,N_1866);
nand U8701 (N_8701,N_2539,N_4710);
or U8702 (N_8702,N_629,N_820);
nor U8703 (N_8703,N_3994,N_4275);
nor U8704 (N_8704,N_2690,N_750);
nor U8705 (N_8705,N_4009,N_487);
or U8706 (N_8706,N_982,N_614);
nor U8707 (N_8707,N_409,N_4549);
or U8708 (N_8708,N_3875,N_1366);
or U8709 (N_8709,N_3535,N_1183);
nor U8710 (N_8710,N_771,N_1313);
nand U8711 (N_8711,N_3773,N_2321);
and U8712 (N_8712,N_4345,N_4483);
or U8713 (N_8713,N_314,N_653);
or U8714 (N_8714,N_3836,N_4669);
nor U8715 (N_8715,N_3744,N_4554);
nor U8716 (N_8716,N_3844,N_1681);
nand U8717 (N_8717,N_943,N_1760);
and U8718 (N_8718,N_2544,N_1467);
nor U8719 (N_8719,N_3049,N_1009);
and U8720 (N_8720,N_285,N_1767);
nand U8721 (N_8721,N_1361,N_1453);
nand U8722 (N_8722,N_1667,N_4209);
nand U8723 (N_8723,N_2792,N_4519);
and U8724 (N_8724,N_580,N_4267);
or U8725 (N_8725,N_511,N_3793);
nand U8726 (N_8726,N_655,N_4940);
nand U8727 (N_8727,N_1808,N_4308);
and U8728 (N_8728,N_787,N_2390);
nand U8729 (N_8729,N_4828,N_4865);
and U8730 (N_8730,N_191,N_3002);
nand U8731 (N_8731,N_4503,N_735);
or U8732 (N_8732,N_4262,N_2317);
or U8733 (N_8733,N_3777,N_1849);
nor U8734 (N_8734,N_928,N_4541);
or U8735 (N_8735,N_996,N_3489);
or U8736 (N_8736,N_1544,N_4443);
nand U8737 (N_8737,N_2263,N_4348);
and U8738 (N_8738,N_3923,N_2522);
and U8739 (N_8739,N_4047,N_2927);
nand U8740 (N_8740,N_1794,N_225);
and U8741 (N_8741,N_2609,N_4638);
or U8742 (N_8742,N_1535,N_3078);
nor U8743 (N_8743,N_1359,N_4072);
xor U8744 (N_8744,N_2754,N_2247);
or U8745 (N_8745,N_4754,N_3206);
nand U8746 (N_8746,N_1037,N_2464);
or U8747 (N_8747,N_459,N_1775);
or U8748 (N_8748,N_1359,N_700);
nand U8749 (N_8749,N_351,N_3837);
nand U8750 (N_8750,N_224,N_3290);
nand U8751 (N_8751,N_3560,N_4444);
or U8752 (N_8752,N_687,N_2797);
nor U8753 (N_8753,N_1445,N_1919);
nand U8754 (N_8754,N_2898,N_802);
and U8755 (N_8755,N_4291,N_4296);
and U8756 (N_8756,N_4195,N_3894);
or U8757 (N_8757,N_2974,N_3666);
nand U8758 (N_8758,N_3783,N_3556);
and U8759 (N_8759,N_4851,N_1747);
nand U8760 (N_8760,N_2561,N_2764);
nand U8761 (N_8761,N_2676,N_1346);
nand U8762 (N_8762,N_4216,N_1064);
nand U8763 (N_8763,N_2823,N_3290);
and U8764 (N_8764,N_1370,N_867);
and U8765 (N_8765,N_535,N_4093);
nand U8766 (N_8766,N_1584,N_1146);
nor U8767 (N_8767,N_2960,N_3429);
nor U8768 (N_8768,N_4710,N_4336);
and U8769 (N_8769,N_4350,N_1793);
nand U8770 (N_8770,N_4778,N_1730);
or U8771 (N_8771,N_1988,N_874);
nand U8772 (N_8772,N_3480,N_3957);
nand U8773 (N_8773,N_2454,N_2499);
or U8774 (N_8774,N_419,N_3590);
nand U8775 (N_8775,N_1621,N_1278);
and U8776 (N_8776,N_1174,N_3484);
or U8777 (N_8777,N_624,N_1714);
or U8778 (N_8778,N_3522,N_1675);
nor U8779 (N_8779,N_4912,N_2799);
nand U8780 (N_8780,N_2660,N_3191);
and U8781 (N_8781,N_875,N_1564);
nor U8782 (N_8782,N_4160,N_3048);
and U8783 (N_8783,N_1537,N_836);
and U8784 (N_8784,N_3715,N_705);
and U8785 (N_8785,N_1036,N_1875);
and U8786 (N_8786,N_4885,N_3452);
nand U8787 (N_8787,N_1455,N_4927);
and U8788 (N_8788,N_2877,N_2537);
and U8789 (N_8789,N_924,N_959);
and U8790 (N_8790,N_4388,N_3258);
and U8791 (N_8791,N_4908,N_830);
or U8792 (N_8792,N_2318,N_1248);
nand U8793 (N_8793,N_406,N_605);
or U8794 (N_8794,N_4556,N_4048);
and U8795 (N_8795,N_1533,N_119);
or U8796 (N_8796,N_2286,N_4281);
nor U8797 (N_8797,N_85,N_3729);
nand U8798 (N_8798,N_2347,N_4510);
nand U8799 (N_8799,N_3713,N_2372);
nor U8800 (N_8800,N_1508,N_3788);
and U8801 (N_8801,N_101,N_3568);
nand U8802 (N_8802,N_2087,N_1169);
nand U8803 (N_8803,N_4365,N_4087);
or U8804 (N_8804,N_1845,N_4086);
nand U8805 (N_8805,N_3291,N_1952);
nor U8806 (N_8806,N_4136,N_4251);
nor U8807 (N_8807,N_4823,N_1017);
nor U8808 (N_8808,N_889,N_1133);
or U8809 (N_8809,N_1576,N_2410);
nor U8810 (N_8810,N_2104,N_1224);
nor U8811 (N_8811,N_378,N_4187);
nor U8812 (N_8812,N_890,N_3352);
nor U8813 (N_8813,N_674,N_4571);
nor U8814 (N_8814,N_3414,N_3608);
or U8815 (N_8815,N_2603,N_3297);
or U8816 (N_8816,N_3684,N_4510);
nor U8817 (N_8817,N_233,N_548);
and U8818 (N_8818,N_933,N_4994);
and U8819 (N_8819,N_670,N_2051);
and U8820 (N_8820,N_1220,N_3650);
nand U8821 (N_8821,N_2964,N_1560);
nand U8822 (N_8822,N_148,N_3315);
nor U8823 (N_8823,N_3762,N_214);
nor U8824 (N_8824,N_1768,N_28);
nor U8825 (N_8825,N_3891,N_1765);
and U8826 (N_8826,N_3522,N_2825);
and U8827 (N_8827,N_4592,N_3311);
nor U8828 (N_8828,N_549,N_3074);
and U8829 (N_8829,N_2825,N_4841);
and U8830 (N_8830,N_1295,N_4107);
and U8831 (N_8831,N_2183,N_3125);
nand U8832 (N_8832,N_1764,N_979);
or U8833 (N_8833,N_4358,N_2941);
and U8834 (N_8834,N_4422,N_3124);
nor U8835 (N_8835,N_2533,N_4792);
and U8836 (N_8836,N_4166,N_4538);
nor U8837 (N_8837,N_3879,N_1843);
or U8838 (N_8838,N_708,N_3384);
nor U8839 (N_8839,N_4363,N_3703);
or U8840 (N_8840,N_3548,N_2937);
and U8841 (N_8841,N_2116,N_1377);
nor U8842 (N_8842,N_191,N_2780);
nand U8843 (N_8843,N_4778,N_1999);
or U8844 (N_8844,N_2268,N_3275);
and U8845 (N_8845,N_3864,N_677);
nor U8846 (N_8846,N_4780,N_327);
or U8847 (N_8847,N_1589,N_1361);
nor U8848 (N_8848,N_1156,N_2122);
nor U8849 (N_8849,N_4941,N_4813);
nor U8850 (N_8850,N_1356,N_1226);
and U8851 (N_8851,N_3179,N_403);
and U8852 (N_8852,N_628,N_3865);
and U8853 (N_8853,N_3696,N_923);
xnor U8854 (N_8854,N_1238,N_775);
nor U8855 (N_8855,N_4419,N_2609);
nand U8856 (N_8856,N_4739,N_600);
nand U8857 (N_8857,N_1323,N_2467);
nor U8858 (N_8858,N_1447,N_3311);
nand U8859 (N_8859,N_3112,N_4297);
nand U8860 (N_8860,N_1919,N_2846);
nand U8861 (N_8861,N_2684,N_2107);
nand U8862 (N_8862,N_654,N_127);
nor U8863 (N_8863,N_78,N_4723);
or U8864 (N_8864,N_1949,N_2047);
or U8865 (N_8865,N_1036,N_605);
and U8866 (N_8866,N_3572,N_906);
nand U8867 (N_8867,N_1437,N_785);
nor U8868 (N_8868,N_1010,N_2601);
nor U8869 (N_8869,N_762,N_1611);
and U8870 (N_8870,N_376,N_129);
nand U8871 (N_8871,N_4069,N_605);
or U8872 (N_8872,N_4930,N_1227);
and U8873 (N_8873,N_1227,N_2609);
nand U8874 (N_8874,N_835,N_653);
and U8875 (N_8875,N_605,N_2472);
and U8876 (N_8876,N_665,N_1037);
or U8877 (N_8877,N_4065,N_164);
nor U8878 (N_8878,N_3141,N_1858);
nor U8879 (N_8879,N_385,N_4506);
or U8880 (N_8880,N_4430,N_279);
nand U8881 (N_8881,N_2521,N_3228);
nor U8882 (N_8882,N_295,N_176);
or U8883 (N_8883,N_2271,N_2016);
and U8884 (N_8884,N_4464,N_2908);
nor U8885 (N_8885,N_663,N_920);
or U8886 (N_8886,N_3859,N_293);
nor U8887 (N_8887,N_4059,N_4977);
nor U8888 (N_8888,N_4509,N_799);
and U8889 (N_8889,N_330,N_1717);
or U8890 (N_8890,N_2701,N_25);
nand U8891 (N_8891,N_2788,N_3125);
or U8892 (N_8892,N_4204,N_2347);
and U8893 (N_8893,N_4381,N_2618);
and U8894 (N_8894,N_4396,N_2016);
nor U8895 (N_8895,N_2192,N_2556);
nor U8896 (N_8896,N_3873,N_1169);
or U8897 (N_8897,N_845,N_2181);
or U8898 (N_8898,N_1131,N_65);
or U8899 (N_8899,N_887,N_1455);
or U8900 (N_8900,N_2541,N_2917);
nand U8901 (N_8901,N_2278,N_2407);
or U8902 (N_8902,N_454,N_4384);
or U8903 (N_8903,N_1901,N_3272);
or U8904 (N_8904,N_4114,N_1889);
or U8905 (N_8905,N_3833,N_1669);
nor U8906 (N_8906,N_2723,N_291);
and U8907 (N_8907,N_4993,N_3605);
or U8908 (N_8908,N_1178,N_2569);
nor U8909 (N_8909,N_3769,N_4826);
and U8910 (N_8910,N_3138,N_3076);
or U8911 (N_8911,N_2933,N_1588);
nand U8912 (N_8912,N_1510,N_1904);
or U8913 (N_8913,N_3811,N_315);
nand U8914 (N_8914,N_3599,N_1353);
nor U8915 (N_8915,N_3568,N_3537);
or U8916 (N_8916,N_2071,N_4850);
or U8917 (N_8917,N_304,N_2646);
and U8918 (N_8918,N_727,N_1913);
nor U8919 (N_8919,N_4313,N_1770);
or U8920 (N_8920,N_1149,N_3489);
nand U8921 (N_8921,N_1828,N_3508);
and U8922 (N_8922,N_379,N_4660);
or U8923 (N_8923,N_2069,N_3033);
nand U8924 (N_8924,N_99,N_94);
and U8925 (N_8925,N_1089,N_115);
and U8926 (N_8926,N_2770,N_1054);
nand U8927 (N_8927,N_2333,N_856);
and U8928 (N_8928,N_461,N_2230);
nand U8929 (N_8929,N_4560,N_3687);
nor U8930 (N_8930,N_2876,N_4454);
nand U8931 (N_8931,N_4468,N_2183);
and U8932 (N_8932,N_3512,N_44);
nor U8933 (N_8933,N_4148,N_1822);
and U8934 (N_8934,N_1453,N_897);
or U8935 (N_8935,N_4238,N_110);
and U8936 (N_8936,N_2218,N_2741);
or U8937 (N_8937,N_125,N_2359);
and U8938 (N_8938,N_2400,N_3762);
or U8939 (N_8939,N_2936,N_1061);
nor U8940 (N_8940,N_1433,N_2453);
or U8941 (N_8941,N_2463,N_186);
nand U8942 (N_8942,N_3085,N_194);
nor U8943 (N_8943,N_1751,N_3503);
and U8944 (N_8944,N_4597,N_77);
or U8945 (N_8945,N_424,N_1390);
nor U8946 (N_8946,N_1653,N_4656);
or U8947 (N_8947,N_4769,N_4054);
nor U8948 (N_8948,N_3860,N_4196);
or U8949 (N_8949,N_1571,N_1284);
or U8950 (N_8950,N_3506,N_2893);
nor U8951 (N_8951,N_2334,N_4299);
and U8952 (N_8952,N_3522,N_2776);
and U8953 (N_8953,N_1711,N_3620);
nand U8954 (N_8954,N_203,N_3720);
nand U8955 (N_8955,N_1530,N_3295);
nand U8956 (N_8956,N_3718,N_545);
nor U8957 (N_8957,N_592,N_755);
xor U8958 (N_8958,N_2255,N_2949);
nand U8959 (N_8959,N_4553,N_1648);
nor U8960 (N_8960,N_4313,N_1661);
and U8961 (N_8961,N_3797,N_1596);
and U8962 (N_8962,N_4607,N_1395);
nand U8963 (N_8963,N_1305,N_1806);
or U8964 (N_8964,N_4228,N_3213);
nand U8965 (N_8965,N_4218,N_1555);
and U8966 (N_8966,N_4686,N_1479);
nor U8967 (N_8967,N_2816,N_4775);
or U8968 (N_8968,N_593,N_3224);
and U8969 (N_8969,N_3352,N_682);
and U8970 (N_8970,N_4847,N_4361);
nand U8971 (N_8971,N_1429,N_474);
and U8972 (N_8972,N_3878,N_4427);
or U8973 (N_8973,N_915,N_4076);
nor U8974 (N_8974,N_4073,N_4163);
nor U8975 (N_8975,N_545,N_1839);
or U8976 (N_8976,N_3025,N_410);
or U8977 (N_8977,N_4334,N_274);
and U8978 (N_8978,N_4806,N_1049);
or U8979 (N_8979,N_3387,N_2409);
and U8980 (N_8980,N_1722,N_2516);
nor U8981 (N_8981,N_347,N_2234);
nor U8982 (N_8982,N_4513,N_4042);
nor U8983 (N_8983,N_4605,N_2433);
and U8984 (N_8984,N_2008,N_2019);
and U8985 (N_8985,N_1373,N_908);
and U8986 (N_8986,N_2018,N_4335);
and U8987 (N_8987,N_1308,N_2529);
nor U8988 (N_8988,N_899,N_4566);
or U8989 (N_8989,N_2451,N_4683);
or U8990 (N_8990,N_479,N_244);
nor U8991 (N_8991,N_4985,N_3841);
or U8992 (N_8992,N_721,N_3638);
nand U8993 (N_8993,N_3388,N_2311);
and U8994 (N_8994,N_3846,N_529);
and U8995 (N_8995,N_2619,N_2364);
nor U8996 (N_8996,N_770,N_3338);
or U8997 (N_8997,N_4226,N_3887);
nor U8998 (N_8998,N_3695,N_1577);
nor U8999 (N_8999,N_1396,N_4324);
and U9000 (N_9000,N_2369,N_3389);
or U9001 (N_9001,N_2898,N_1607);
nor U9002 (N_9002,N_765,N_2824);
and U9003 (N_9003,N_1937,N_1550);
nand U9004 (N_9004,N_4657,N_1860);
nand U9005 (N_9005,N_1925,N_3509);
and U9006 (N_9006,N_4030,N_2220);
and U9007 (N_9007,N_1461,N_4322);
and U9008 (N_9008,N_565,N_900);
or U9009 (N_9009,N_931,N_3870);
or U9010 (N_9010,N_3103,N_1197);
or U9011 (N_9011,N_3781,N_2774);
nor U9012 (N_9012,N_3435,N_1487);
nor U9013 (N_9013,N_4805,N_3814);
and U9014 (N_9014,N_1200,N_4092);
nand U9015 (N_9015,N_4993,N_3235);
nand U9016 (N_9016,N_3693,N_1085);
nor U9017 (N_9017,N_2407,N_1130);
and U9018 (N_9018,N_4379,N_1540);
nand U9019 (N_9019,N_4446,N_3192);
nand U9020 (N_9020,N_1953,N_2204);
nand U9021 (N_9021,N_3505,N_2572);
nand U9022 (N_9022,N_3166,N_2944);
nand U9023 (N_9023,N_3946,N_50);
or U9024 (N_9024,N_541,N_2629);
nor U9025 (N_9025,N_1961,N_815);
nor U9026 (N_9026,N_3660,N_2732);
or U9027 (N_9027,N_743,N_706);
nor U9028 (N_9028,N_2958,N_4385);
or U9029 (N_9029,N_3224,N_2194);
or U9030 (N_9030,N_2896,N_2091);
nand U9031 (N_9031,N_4512,N_1401);
and U9032 (N_9032,N_486,N_4464);
nand U9033 (N_9033,N_3832,N_2522);
nor U9034 (N_9034,N_3218,N_2652);
nand U9035 (N_9035,N_2713,N_2223);
nor U9036 (N_9036,N_3562,N_2252);
nand U9037 (N_9037,N_649,N_2595);
and U9038 (N_9038,N_3472,N_4220);
or U9039 (N_9039,N_3569,N_661);
nor U9040 (N_9040,N_3705,N_2447);
nor U9041 (N_9041,N_4602,N_3082);
and U9042 (N_9042,N_2709,N_4580);
nor U9043 (N_9043,N_1913,N_4378);
nor U9044 (N_9044,N_878,N_1931);
and U9045 (N_9045,N_3497,N_2320);
nor U9046 (N_9046,N_2115,N_3193);
nand U9047 (N_9047,N_3574,N_3793);
or U9048 (N_9048,N_94,N_508);
and U9049 (N_9049,N_4820,N_2865);
or U9050 (N_9050,N_3414,N_1575);
and U9051 (N_9051,N_2985,N_2772);
and U9052 (N_9052,N_556,N_2201);
nand U9053 (N_9053,N_3034,N_3447);
nor U9054 (N_9054,N_3554,N_3114);
nand U9055 (N_9055,N_4725,N_3681);
nor U9056 (N_9056,N_3535,N_3981);
and U9057 (N_9057,N_4605,N_904);
nor U9058 (N_9058,N_4616,N_11);
and U9059 (N_9059,N_1793,N_490);
nand U9060 (N_9060,N_3391,N_923);
and U9061 (N_9061,N_3887,N_2040);
nor U9062 (N_9062,N_457,N_4941);
and U9063 (N_9063,N_1483,N_1073);
nor U9064 (N_9064,N_4577,N_4853);
nand U9065 (N_9065,N_16,N_2819);
nand U9066 (N_9066,N_3152,N_844);
or U9067 (N_9067,N_3366,N_3268);
and U9068 (N_9068,N_931,N_105);
nand U9069 (N_9069,N_254,N_3382);
nor U9070 (N_9070,N_1941,N_4954);
nand U9071 (N_9071,N_3095,N_4423);
or U9072 (N_9072,N_3409,N_1774);
and U9073 (N_9073,N_3940,N_834);
or U9074 (N_9074,N_3369,N_4230);
nand U9075 (N_9075,N_4152,N_631);
nand U9076 (N_9076,N_563,N_3529);
nand U9077 (N_9077,N_2174,N_1720);
nor U9078 (N_9078,N_4714,N_2390);
or U9079 (N_9079,N_1769,N_1585);
nor U9080 (N_9080,N_3499,N_709);
nand U9081 (N_9081,N_4740,N_1343);
nor U9082 (N_9082,N_330,N_393);
and U9083 (N_9083,N_2752,N_3958);
nor U9084 (N_9084,N_3199,N_4993);
and U9085 (N_9085,N_1695,N_382);
nand U9086 (N_9086,N_2959,N_4192);
nand U9087 (N_9087,N_2458,N_3058);
or U9088 (N_9088,N_651,N_60);
or U9089 (N_9089,N_4803,N_1815);
nand U9090 (N_9090,N_1709,N_2787);
and U9091 (N_9091,N_2066,N_1368);
nor U9092 (N_9092,N_3317,N_529);
and U9093 (N_9093,N_4889,N_2289);
nand U9094 (N_9094,N_1600,N_3383);
or U9095 (N_9095,N_1474,N_3018);
nand U9096 (N_9096,N_1762,N_4817);
nor U9097 (N_9097,N_3158,N_4405);
nand U9098 (N_9098,N_1663,N_360);
nor U9099 (N_9099,N_2180,N_4832);
nand U9100 (N_9100,N_4695,N_2019);
or U9101 (N_9101,N_4523,N_2764);
xor U9102 (N_9102,N_1013,N_2224);
or U9103 (N_9103,N_1048,N_4845);
nor U9104 (N_9104,N_2841,N_2946);
or U9105 (N_9105,N_4760,N_4323);
nand U9106 (N_9106,N_708,N_3496);
nor U9107 (N_9107,N_911,N_1676);
and U9108 (N_9108,N_4185,N_2242);
or U9109 (N_9109,N_99,N_890);
or U9110 (N_9110,N_1621,N_677);
and U9111 (N_9111,N_634,N_3601);
or U9112 (N_9112,N_3874,N_939);
or U9113 (N_9113,N_4686,N_3925);
and U9114 (N_9114,N_2785,N_2367);
or U9115 (N_9115,N_996,N_833);
nand U9116 (N_9116,N_1945,N_102);
and U9117 (N_9117,N_3521,N_1859);
or U9118 (N_9118,N_447,N_3700);
and U9119 (N_9119,N_2779,N_3953);
nand U9120 (N_9120,N_1566,N_4323);
or U9121 (N_9121,N_3050,N_1573);
nand U9122 (N_9122,N_2838,N_4570);
nor U9123 (N_9123,N_2847,N_2769);
and U9124 (N_9124,N_972,N_1528);
or U9125 (N_9125,N_4633,N_4790);
or U9126 (N_9126,N_4519,N_1427);
nand U9127 (N_9127,N_4735,N_3345);
and U9128 (N_9128,N_2880,N_114);
and U9129 (N_9129,N_4902,N_1939);
nand U9130 (N_9130,N_4532,N_3153);
and U9131 (N_9131,N_2905,N_1062);
nor U9132 (N_9132,N_884,N_2394);
nor U9133 (N_9133,N_3475,N_4249);
nor U9134 (N_9134,N_3350,N_1993);
nor U9135 (N_9135,N_3187,N_1264);
and U9136 (N_9136,N_846,N_3806);
or U9137 (N_9137,N_1616,N_3624);
nor U9138 (N_9138,N_1549,N_2203);
and U9139 (N_9139,N_583,N_3263);
nand U9140 (N_9140,N_268,N_2088);
xor U9141 (N_9141,N_478,N_4789);
or U9142 (N_9142,N_2615,N_1142);
nor U9143 (N_9143,N_204,N_4052);
and U9144 (N_9144,N_159,N_3693);
and U9145 (N_9145,N_2365,N_708);
and U9146 (N_9146,N_3344,N_4642);
or U9147 (N_9147,N_2463,N_892);
or U9148 (N_9148,N_273,N_4750);
and U9149 (N_9149,N_2164,N_1256);
xnor U9150 (N_9150,N_1485,N_1795);
or U9151 (N_9151,N_739,N_2754);
nor U9152 (N_9152,N_4451,N_3168);
and U9153 (N_9153,N_4311,N_4051);
nand U9154 (N_9154,N_63,N_2869);
and U9155 (N_9155,N_3323,N_2521);
nand U9156 (N_9156,N_3044,N_3394);
nor U9157 (N_9157,N_495,N_2911);
nand U9158 (N_9158,N_1796,N_3776);
or U9159 (N_9159,N_4591,N_4387);
and U9160 (N_9160,N_4172,N_3396);
or U9161 (N_9161,N_4790,N_1540);
or U9162 (N_9162,N_3489,N_2926);
nand U9163 (N_9163,N_1588,N_4489);
or U9164 (N_9164,N_1805,N_506);
nor U9165 (N_9165,N_3971,N_2368);
and U9166 (N_9166,N_2937,N_4636);
or U9167 (N_9167,N_4293,N_3770);
or U9168 (N_9168,N_1842,N_13);
and U9169 (N_9169,N_4425,N_2143);
nand U9170 (N_9170,N_4836,N_3847);
nand U9171 (N_9171,N_541,N_3197);
and U9172 (N_9172,N_443,N_2668);
nand U9173 (N_9173,N_2366,N_3035);
nor U9174 (N_9174,N_2504,N_1759);
nand U9175 (N_9175,N_4232,N_401);
and U9176 (N_9176,N_3142,N_4050);
or U9177 (N_9177,N_4273,N_4796);
or U9178 (N_9178,N_2444,N_2669);
nor U9179 (N_9179,N_1938,N_3488);
nand U9180 (N_9180,N_1365,N_4583);
nor U9181 (N_9181,N_2781,N_3319);
nand U9182 (N_9182,N_20,N_4733);
nand U9183 (N_9183,N_244,N_1556);
nor U9184 (N_9184,N_420,N_2465);
nor U9185 (N_9185,N_4437,N_906);
or U9186 (N_9186,N_2916,N_462);
or U9187 (N_9187,N_3078,N_1510);
nand U9188 (N_9188,N_1115,N_695);
nand U9189 (N_9189,N_4467,N_2557);
and U9190 (N_9190,N_1007,N_1934);
and U9191 (N_9191,N_1753,N_1791);
and U9192 (N_9192,N_2790,N_98);
nand U9193 (N_9193,N_1802,N_4352);
nor U9194 (N_9194,N_999,N_3452);
nand U9195 (N_9195,N_2557,N_1062);
and U9196 (N_9196,N_662,N_800);
nand U9197 (N_9197,N_1991,N_1508);
or U9198 (N_9198,N_341,N_3431);
and U9199 (N_9199,N_3557,N_3497);
nor U9200 (N_9200,N_3751,N_840);
nor U9201 (N_9201,N_3917,N_1586);
and U9202 (N_9202,N_4947,N_4897);
nand U9203 (N_9203,N_4981,N_2391);
and U9204 (N_9204,N_1453,N_3930);
nor U9205 (N_9205,N_208,N_4344);
nand U9206 (N_9206,N_2795,N_2747);
and U9207 (N_9207,N_530,N_2196);
nand U9208 (N_9208,N_668,N_2852);
or U9209 (N_9209,N_4583,N_3371);
and U9210 (N_9210,N_2747,N_2350);
and U9211 (N_9211,N_1781,N_368);
and U9212 (N_9212,N_2206,N_3561);
nand U9213 (N_9213,N_1559,N_4517);
and U9214 (N_9214,N_2269,N_3957);
nand U9215 (N_9215,N_1047,N_253);
nor U9216 (N_9216,N_751,N_2913);
or U9217 (N_9217,N_4521,N_793);
and U9218 (N_9218,N_423,N_2129);
or U9219 (N_9219,N_1611,N_4551);
or U9220 (N_9220,N_804,N_1059);
or U9221 (N_9221,N_4999,N_2203);
nand U9222 (N_9222,N_2323,N_3061);
nor U9223 (N_9223,N_1451,N_4982);
nand U9224 (N_9224,N_242,N_3983);
and U9225 (N_9225,N_2987,N_1409);
and U9226 (N_9226,N_338,N_4120);
nand U9227 (N_9227,N_1238,N_784);
nand U9228 (N_9228,N_970,N_541);
and U9229 (N_9229,N_4827,N_2731);
nor U9230 (N_9230,N_4636,N_1791);
nor U9231 (N_9231,N_4997,N_3623);
nand U9232 (N_9232,N_4239,N_349);
nand U9233 (N_9233,N_820,N_3387);
nor U9234 (N_9234,N_2014,N_4592);
and U9235 (N_9235,N_647,N_4019);
or U9236 (N_9236,N_1564,N_4553);
nor U9237 (N_9237,N_4311,N_2510);
nand U9238 (N_9238,N_1629,N_4861);
nand U9239 (N_9239,N_1359,N_2452);
nand U9240 (N_9240,N_805,N_580);
nand U9241 (N_9241,N_1119,N_4316);
or U9242 (N_9242,N_4352,N_3365);
and U9243 (N_9243,N_1481,N_1765);
or U9244 (N_9244,N_4073,N_4667);
nor U9245 (N_9245,N_4387,N_419);
and U9246 (N_9246,N_3975,N_2158);
and U9247 (N_9247,N_3230,N_610);
or U9248 (N_9248,N_4582,N_518);
and U9249 (N_9249,N_3883,N_3393);
nand U9250 (N_9250,N_1456,N_3906);
nor U9251 (N_9251,N_2593,N_4000);
nor U9252 (N_9252,N_3811,N_3538);
or U9253 (N_9253,N_899,N_3738);
nand U9254 (N_9254,N_453,N_4155);
or U9255 (N_9255,N_3705,N_3423);
nor U9256 (N_9256,N_1257,N_2346);
nor U9257 (N_9257,N_2748,N_3421);
nor U9258 (N_9258,N_4745,N_4331);
or U9259 (N_9259,N_3570,N_1033);
or U9260 (N_9260,N_3730,N_2518);
nor U9261 (N_9261,N_178,N_1677);
and U9262 (N_9262,N_1032,N_3496);
and U9263 (N_9263,N_1501,N_996);
nand U9264 (N_9264,N_4864,N_4108);
nand U9265 (N_9265,N_1955,N_1992);
nor U9266 (N_9266,N_4402,N_1993);
nand U9267 (N_9267,N_682,N_3905);
nand U9268 (N_9268,N_1212,N_4668);
nand U9269 (N_9269,N_1607,N_2337);
and U9270 (N_9270,N_1054,N_4252);
and U9271 (N_9271,N_3039,N_782);
nand U9272 (N_9272,N_2636,N_2711);
nand U9273 (N_9273,N_2167,N_4053);
nand U9274 (N_9274,N_1157,N_2940);
and U9275 (N_9275,N_2233,N_4839);
or U9276 (N_9276,N_1830,N_4859);
and U9277 (N_9277,N_1433,N_3738);
xnor U9278 (N_9278,N_2715,N_37);
or U9279 (N_9279,N_3432,N_309);
or U9280 (N_9280,N_1089,N_2349);
nor U9281 (N_9281,N_1566,N_4670);
nand U9282 (N_9282,N_4200,N_2601);
nand U9283 (N_9283,N_3737,N_3335);
or U9284 (N_9284,N_861,N_1383);
or U9285 (N_9285,N_3117,N_4825);
nor U9286 (N_9286,N_2662,N_14);
or U9287 (N_9287,N_1555,N_608);
nand U9288 (N_9288,N_4294,N_334);
nor U9289 (N_9289,N_259,N_4200);
or U9290 (N_9290,N_243,N_1147);
xor U9291 (N_9291,N_1124,N_4088);
nand U9292 (N_9292,N_1863,N_4141);
and U9293 (N_9293,N_1152,N_3820);
nor U9294 (N_9294,N_953,N_267);
nand U9295 (N_9295,N_4415,N_3849);
or U9296 (N_9296,N_4596,N_1185);
and U9297 (N_9297,N_1468,N_4648);
nand U9298 (N_9298,N_1427,N_1863);
or U9299 (N_9299,N_3756,N_2460);
and U9300 (N_9300,N_2960,N_1932);
or U9301 (N_9301,N_739,N_1983);
nand U9302 (N_9302,N_4611,N_2944);
nand U9303 (N_9303,N_4256,N_2828);
nand U9304 (N_9304,N_1337,N_1052);
and U9305 (N_9305,N_3217,N_4297);
or U9306 (N_9306,N_4392,N_608);
or U9307 (N_9307,N_2538,N_4770);
and U9308 (N_9308,N_188,N_2858);
or U9309 (N_9309,N_2568,N_4699);
and U9310 (N_9310,N_2327,N_491);
nor U9311 (N_9311,N_1701,N_940);
or U9312 (N_9312,N_3123,N_2657);
nor U9313 (N_9313,N_4322,N_1166);
and U9314 (N_9314,N_1935,N_2723);
or U9315 (N_9315,N_2020,N_2928);
and U9316 (N_9316,N_2792,N_185);
nor U9317 (N_9317,N_956,N_4457);
nor U9318 (N_9318,N_1731,N_1086);
and U9319 (N_9319,N_121,N_4933);
nor U9320 (N_9320,N_1751,N_4051);
or U9321 (N_9321,N_2105,N_1293);
and U9322 (N_9322,N_4973,N_611);
and U9323 (N_9323,N_4769,N_3444);
and U9324 (N_9324,N_3015,N_2053);
or U9325 (N_9325,N_3079,N_4470);
nand U9326 (N_9326,N_1598,N_4745);
nor U9327 (N_9327,N_21,N_2280);
nand U9328 (N_9328,N_4525,N_4721);
nand U9329 (N_9329,N_2815,N_1621);
nor U9330 (N_9330,N_3421,N_3163);
or U9331 (N_9331,N_341,N_2384);
nor U9332 (N_9332,N_1159,N_1130);
nor U9333 (N_9333,N_424,N_1698);
and U9334 (N_9334,N_4189,N_2630);
or U9335 (N_9335,N_2613,N_598);
nor U9336 (N_9336,N_82,N_2126);
and U9337 (N_9337,N_4076,N_2804);
nand U9338 (N_9338,N_1405,N_3381);
and U9339 (N_9339,N_189,N_4658);
nor U9340 (N_9340,N_3724,N_2762);
and U9341 (N_9341,N_3657,N_1732);
and U9342 (N_9342,N_2422,N_3098);
nand U9343 (N_9343,N_3614,N_707);
or U9344 (N_9344,N_4459,N_2057);
and U9345 (N_9345,N_3613,N_3483);
nor U9346 (N_9346,N_3729,N_2933);
nand U9347 (N_9347,N_3294,N_4192);
nand U9348 (N_9348,N_61,N_4494);
nor U9349 (N_9349,N_1794,N_1518);
nand U9350 (N_9350,N_3364,N_3046);
or U9351 (N_9351,N_3660,N_4239);
nand U9352 (N_9352,N_4100,N_4104);
nand U9353 (N_9353,N_396,N_1342);
or U9354 (N_9354,N_3924,N_3248);
nor U9355 (N_9355,N_721,N_4779);
and U9356 (N_9356,N_1092,N_1896);
or U9357 (N_9357,N_2404,N_78);
or U9358 (N_9358,N_963,N_1918);
and U9359 (N_9359,N_1954,N_743);
or U9360 (N_9360,N_232,N_426);
nor U9361 (N_9361,N_4915,N_307);
or U9362 (N_9362,N_1967,N_4680);
and U9363 (N_9363,N_139,N_3704);
nand U9364 (N_9364,N_822,N_2174);
nand U9365 (N_9365,N_1121,N_875);
nor U9366 (N_9366,N_1060,N_3438);
and U9367 (N_9367,N_4712,N_2519);
and U9368 (N_9368,N_425,N_4699);
and U9369 (N_9369,N_3639,N_1615);
or U9370 (N_9370,N_793,N_152);
and U9371 (N_9371,N_3553,N_3755);
nor U9372 (N_9372,N_723,N_2103);
or U9373 (N_9373,N_3618,N_4937);
or U9374 (N_9374,N_922,N_2345);
nor U9375 (N_9375,N_3985,N_4431);
or U9376 (N_9376,N_4074,N_3404);
nor U9377 (N_9377,N_3746,N_3353);
or U9378 (N_9378,N_1229,N_3443);
nand U9379 (N_9379,N_438,N_4292);
or U9380 (N_9380,N_2400,N_1719);
nor U9381 (N_9381,N_1030,N_4942);
and U9382 (N_9382,N_3017,N_354);
nor U9383 (N_9383,N_2,N_563);
nand U9384 (N_9384,N_1771,N_1056);
nand U9385 (N_9385,N_1233,N_3426);
nand U9386 (N_9386,N_2847,N_4734);
nand U9387 (N_9387,N_2670,N_4004);
nor U9388 (N_9388,N_1445,N_49);
nand U9389 (N_9389,N_464,N_4720);
and U9390 (N_9390,N_1735,N_3105);
or U9391 (N_9391,N_3020,N_4795);
nand U9392 (N_9392,N_4890,N_3204);
nor U9393 (N_9393,N_4766,N_3252);
nor U9394 (N_9394,N_4861,N_4387);
nor U9395 (N_9395,N_786,N_2123);
and U9396 (N_9396,N_1038,N_1299);
or U9397 (N_9397,N_2769,N_450);
nor U9398 (N_9398,N_2781,N_2089);
nand U9399 (N_9399,N_1785,N_2023);
or U9400 (N_9400,N_3136,N_3870);
nor U9401 (N_9401,N_1495,N_4468);
nor U9402 (N_9402,N_4487,N_582);
nor U9403 (N_9403,N_4236,N_1499);
or U9404 (N_9404,N_3006,N_4396);
nand U9405 (N_9405,N_3499,N_4842);
nand U9406 (N_9406,N_4660,N_3838);
or U9407 (N_9407,N_604,N_1082);
nor U9408 (N_9408,N_4285,N_1924);
and U9409 (N_9409,N_4984,N_95);
and U9410 (N_9410,N_675,N_80);
nor U9411 (N_9411,N_4013,N_87);
nor U9412 (N_9412,N_4490,N_4722);
nand U9413 (N_9413,N_2249,N_108);
and U9414 (N_9414,N_1696,N_2719);
nor U9415 (N_9415,N_1169,N_3435);
nand U9416 (N_9416,N_1417,N_3050);
nand U9417 (N_9417,N_4361,N_3523);
nand U9418 (N_9418,N_3093,N_177);
and U9419 (N_9419,N_3184,N_1124);
xnor U9420 (N_9420,N_1442,N_2183);
or U9421 (N_9421,N_3972,N_3270);
nand U9422 (N_9422,N_1449,N_3493);
or U9423 (N_9423,N_2571,N_3597);
or U9424 (N_9424,N_4059,N_1764);
nor U9425 (N_9425,N_2309,N_1788);
nand U9426 (N_9426,N_4437,N_144);
nor U9427 (N_9427,N_2965,N_1687);
nor U9428 (N_9428,N_3068,N_2142);
nand U9429 (N_9429,N_1926,N_41);
or U9430 (N_9430,N_2511,N_4425);
nand U9431 (N_9431,N_4154,N_4648);
and U9432 (N_9432,N_4226,N_784);
nor U9433 (N_9433,N_4046,N_483);
nand U9434 (N_9434,N_1318,N_479);
or U9435 (N_9435,N_4721,N_3602);
and U9436 (N_9436,N_135,N_2957);
and U9437 (N_9437,N_3215,N_4462);
or U9438 (N_9438,N_4430,N_4636);
nor U9439 (N_9439,N_1264,N_4289);
nand U9440 (N_9440,N_145,N_359);
or U9441 (N_9441,N_3874,N_3109);
and U9442 (N_9442,N_2938,N_449);
or U9443 (N_9443,N_4322,N_3120);
and U9444 (N_9444,N_1053,N_2847);
nor U9445 (N_9445,N_3596,N_2826);
xor U9446 (N_9446,N_743,N_337);
nor U9447 (N_9447,N_2104,N_4572);
and U9448 (N_9448,N_885,N_4004);
nor U9449 (N_9449,N_1479,N_4106);
nor U9450 (N_9450,N_4255,N_837);
or U9451 (N_9451,N_2051,N_1369);
and U9452 (N_9452,N_842,N_403);
and U9453 (N_9453,N_4090,N_1174);
nand U9454 (N_9454,N_1022,N_3293);
nor U9455 (N_9455,N_444,N_4919);
nor U9456 (N_9456,N_2770,N_975);
nor U9457 (N_9457,N_2103,N_4401);
and U9458 (N_9458,N_857,N_4217);
or U9459 (N_9459,N_1409,N_967);
nand U9460 (N_9460,N_1990,N_4334);
nor U9461 (N_9461,N_4375,N_1609);
or U9462 (N_9462,N_4425,N_3811);
nor U9463 (N_9463,N_1333,N_1510);
nand U9464 (N_9464,N_3320,N_1406);
and U9465 (N_9465,N_506,N_4994);
and U9466 (N_9466,N_4111,N_859);
or U9467 (N_9467,N_981,N_4876);
nand U9468 (N_9468,N_3302,N_3703);
nand U9469 (N_9469,N_3652,N_1454);
or U9470 (N_9470,N_951,N_3202);
nand U9471 (N_9471,N_920,N_3793);
or U9472 (N_9472,N_209,N_114);
nand U9473 (N_9473,N_2710,N_1021);
and U9474 (N_9474,N_2100,N_2143);
or U9475 (N_9475,N_1483,N_4546);
or U9476 (N_9476,N_1206,N_2603);
or U9477 (N_9477,N_3457,N_805);
nand U9478 (N_9478,N_3492,N_3881);
nor U9479 (N_9479,N_671,N_3365);
nand U9480 (N_9480,N_3247,N_4893);
nor U9481 (N_9481,N_2980,N_2451);
or U9482 (N_9482,N_1688,N_3005);
nor U9483 (N_9483,N_1403,N_3484);
and U9484 (N_9484,N_2026,N_917);
nand U9485 (N_9485,N_3994,N_4308);
or U9486 (N_9486,N_265,N_889);
nand U9487 (N_9487,N_3909,N_1889);
nand U9488 (N_9488,N_3641,N_314);
nor U9489 (N_9489,N_2965,N_1638);
nand U9490 (N_9490,N_2085,N_11);
nand U9491 (N_9491,N_148,N_292);
or U9492 (N_9492,N_1207,N_4715);
or U9493 (N_9493,N_4468,N_2272);
nor U9494 (N_9494,N_4761,N_4458);
nor U9495 (N_9495,N_2419,N_2954);
or U9496 (N_9496,N_1755,N_46);
nor U9497 (N_9497,N_572,N_2246);
and U9498 (N_9498,N_1213,N_4420);
or U9499 (N_9499,N_4727,N_2188);
nor U9500 (N_9500,N_2587,N_2275);
nand U9501 (N_9501,N_4718,N_2210);
or U9502 (N_9502,N_3888,N_2374);
nand U9503 (N_9503,N_3924,N_4429);
and U9504 (N_9504,N_200,N_117);
and U9505 (N_9505,N_1685,N_4997);
nand U9506 (N_9506,N_3127,N_745);
nand U9507 (N_9507,N_3874,N_4526);
nor U9508 (N_9508,N_2026,N_800);
nor U9509 (N_9509,N_2563,N_4443);
and U9510 (N_9510,N_778,N_4039);
nor U9511 (N_9511,N_1741,N_4580);
nor U9512 (N_9512,N_2048,N_3995);
and U9513 (N_9513,N_1179,N_3703);
or U9514 (N_9514,N_3886,N_2188);
and U9515 (N_9515,N_1042,N_538);
or U9516 (N_9516,N_3671,N_3505);
and U9517 (N_9517,N_495,N_2537);
or U9518 (N_9518,N_2176,N_2915);
nand U9519 (N_9519,N_1086,N_2491);
and U9520 (N_9520,N_740,N_4548);
xnor U9521 (N_9521,N_1786,N_2360);
nor U9522 (N_9522,N_4833,N_3560);
nand U9523 (N_9523,N_4792,N_1159);
and U9524 (N_9524,N_2229,N_2755);
and U9525 (N_9525,N_3124,N_1312);
xor U9526 (N_9526,N_2465,N_99);
or U9527 (N_9527,N_737,N_4800);
and U9528 (N_9528,N_817,N_2473);
nand U9529 (N_9529,N_2944,N_606);
and U9530 (N_9530,N_736,N_236);
nand U9531 (N_9531,N_2218,N_1737);
and U9532 (N_9532,N_1923,N_3479);
and U9533 (N_9533,N_869,N_4016);
nor U9534 (N_9534,N_1375,N_249);
or U9535 (N_9535,N_2566,N_1900);
and U9536 (N_9536,N_1403,N_3411);
or U9537 (N_9537,N_1139,N_2347);
nand U9538 (N_9538,N_3307,N_4221);
and U9539 (N_9539,N_1367,N_2032);
or U9540 (N_9540,N_1919,N_2241);
and U9541 (N_9541,N_4446,N_67);
or U9542 (N_9542,N_996,N_2210);
nand U9543 (N_9543,N_4155,N_854);
or U9544 (N_9544,N_101,N_4148);
nand U9545 (N_9545,N_1857,N_2910);
nor U9546 (N_9546,N_59,N_1330);
or U9547 (N_9547,N_1296,N_1216);
or U9548 (N_9548,N_255,N_4113);
nor U9549 (N_9549,N_2113,N_4880);
nand U9550 (N_9550,N_2201,N_1498);
and U9551 (N_9551,N_3927,N_730);
nor U9552 (N_9552,N_829,N_2514);
nor U9553 (N_9553,N_4538,N_1760);
or U9554 (N_9554,N_2754,N_1202);
nand U9555 (N_9555,N_3872,N_2103);
or U9556 (N_9556,N_958,N_3447);
and U9557 (N_9557,N_1461,N_2012);
and U9558 (N_9558,N_3106,N_2472);
nor U9559 (N_9559,N_4251,N_74);
or U9560 (N_9560,N_1972,N_1581);
or U9561 (N_9561,N_4406,N_866);
or U9562 (N_9562,N_4112,N_1249);
or U9563 (N_9563,N_523,N_655);
and U9564 (N_9564,N_2389,N_411);
nand U9565 (N_9565,N_3705,N_3697);
and U9566 (N_9566,N_377,N_4167);
nand U9567 (N_9567,N_1373,N_2648);
nand U9568 (N_9568,N_1160,N_547);
nor U9569 (N_9569,N_2359,N_3691);
nor U9570 (N_9570,N_3284,N_2429);
or U9571 (N_9571,N_3864,N_662);
and U9572 (N_9572,N_352,N_159);
and U9573 (N_9573,N_1064,N_1822);
or U9574 (N_9574,N_1522,N_1154);
nand U9575 (N_9575,N_2776,N_2324);
or U9576 (N_9576,N_3021,N_901);
nand U9577 (N_9577,N_3030,N_662);
nand U9578 (N_9578,N_4786,N_2620);
nor U9579 (N_9579,N_2819,N_166);
or U9580 (N_9580,N_3704,N_2703);
xnor U9581 (N_9581,N_1265,N_3704);
and U9582 (N_9582,N_1485,N_145);
or U9583 (N_9583,N_633,N_4931);
nor U9584 (N_9584,N_2696,N_4603);
or U9585 (N_9585,N_537,N_1572);
nand U9586 (N_9586,N_4348,N_2195);
nor U9587 (N_9587,N_104,N_3593);
nand U9588 (N_9588,N_2103,N_2676);
nand U9589 (N_9589,N_3532,N_3742);
nand U9590 (N_9590,N_3251,N_2839);
or U9591 (N_9591,N_1916,N_4582);
nand U9592 (N_9592,N_3095,N_1088);
nor U9593 (N_9593,N_1868,N_2215);
and U9594 (N_9594,N_1445,N_4623);
nor U9595 (N_9595,N_3802,N_1286);
nor U9596 (N_9596,N_2549,N_2922);
nand U9597 (N_9597,N_2949,N_1665);
nand U9598 (N_9598,N_3595,N_4924);
and U9599 (N_9599,N_3235,N_4864);
nor U9600 (N_9600,N_4117,N_576);
nand U9601 (N_9601,N_3396,N_339);
nand U9602 (N_9602,N_2430,N_856);
or U9603 (N_9603,N_3591,N_355);
nand U9604 (N_9604,N_1603,N_3039);
nor U9605 (N_9605,N_1294,N_1106);
nor U9606 (N_9606,N_702,N_1584);
and U9607 (N_9607,N_1792,N_148);
nand U9608 (N_9608,N_348,N_2816);
nor U9609 (N_9609,N_1939,N_3527);
nor U9610 (N_9610,N_3878,N_4637);
nor U9611 (N_9611,N_1659,N_3497);
and U9612 (N_9612,N_2287,N_3463);
or U9613 (N_9613,N_1267,N_1076);
and U9614 (N_9614,N_3968,N_1568);
and U9615 (N_9615,N_4173,N_3454);
nor U9616 (N_9616,N_4754,N_3762);
nand U9617 (N_9617,N_3538,N_4239);
nor U9618 (N_9618,N_1616,N_337);
or U9619 (N_9619,N_3522,N_967);
nor U9620 (N_9620,N_1871,N_4723);
nand U9621 (N_9621,N_129,N_2850);
nand U9622 (N_9622,N_3274,N_4293);
and U9623 (N_9623,N_2936,N_783);
nand U9624 (N_9624,N_1425,N_1203);
and U9625 (N_9625,N_4538,N_2726);
nor U9626 (N_9626,N_4708,N_3631);
nor U9627 (N_9627,N_315,N_1090);
nand U9628 (N_9628,N_482,N_619);
nor U9629 (N_9629,N_2123,N_4153);
and U9630 (N_9630,N_2492,N_3968);
nor U9631 (N_9631,N_4743,N_3842);
nand U9632 (N_9632,N_1844,N_4673);
nor U9633 (N_9633,N_1175,N_2301);
nor U9634 (N_9634,N_1958,N_1838);
and U9635 (N_9635,N_2876,N_3239);
nand U9636 (N_9636,N_1586,N_3514);
nor U9637 (N_9637,N_1332,N_1493);
nor U9638 (N_9638,N_274,N_4444);
and U9639 (N_9639,N_3085,N_3697);
nand U9640 (N_9640,N_4117,N_366);
or U9641 (N_9641,N_1450,N_1735);
and U9642 (N_9642,N_4338,N_710);
nand U9643 (N_9643,N_2740,N_1038);
and U9644 (N_9644,N_3784,N_906);
or U9645 (N_9645,N_2474,N_4964);
or U9646 (N_9646,N_3272,N_2344);
or U9647 (N_9647,N_2921,N_3876);
and U9648 (N_9648,N_1525,N_260);
nor U9649 (N_9649,N_602,N_2228);
or U9650 (N_9650,N_1475,N_322);
nor U9651 (N_9651,N_1947,N_3606);
or U9652 (N_9652,N_3963,N_2427);
nor U9653 (N_9653,N_1477,N_1324);
or U9654 (N_9654,N_2762,N_4956);
or U9655 (N_9655,N_4191,N_387);
or U9656 (N_9656,N_42,N_636);
and U9657 (N_9657,N_1412,N_3687);
nand U9658 (N_9658,N_926,N_528);
and U9659 (N_9659,N_4328,N_3165);
nand U9660 (N_9660,N_1163,N_2342);
or U9661 (N_9661,N_2905,N_1192);
nand U9662 (N_9662,N_3473,N_4314);
or U9663 (N_9663,N_2643,N_1916);
nand U9664 (N_9664,N_4114,N_1456);
nand U9665 (N_9665,N_3107,N_807);
or U9666 (N_9666,N_3536,N_2684);
nor U9667 (N_9667,N_2453,N_2365);
nor U9668 (N_9668,N_4158,N_2900);
or U9669 (N_9669,N_4758,N_4807);
nand U9670 (N_9670,N_4956,N_3899);
nor U9671 (N_9671,N_4341,N_418);
nor U9672 (N_9672,N_2502,N_66);
nor U9673 (N_9673,N_1,N_4907);
nand U9674 (N_9674,N_4519,N_3776);
nor U9675 (N_9675,N_4553,N_216);
nor U9676 (N_9676,N_363,N_3626);
nor U9677 (N_9677,N_1135,N_3113);
or U9678 (N_9678,N_535,N_1538);
nand U9679 (N_9679,N_4729,N_320);
nor U9680 (N_9680,N_2499,N_4138);
xnor U9681 (N_9681,N_3418,N_4992);
xnor U9682 (N_9682,N_4132,N_96);
and U9683 (N_9683,N_2750,N_512);
nor U9684 (N_9684,N_633,N_2331);
nand U9685 (N_9685,N_166,N_4255);
and U9686 (N_9686,N_1140,N_3956);
nor U9687 (N_9687,N_3638,N_2110);
or U9688 (N_9688,N_4522,N_590);
and U9689 (N_9689,N_3948,N_4034);
or U9690 (N_9690,N_962,N_4324);
nand U9691 (N_9691,N_3757,N_1470);
or U9692 (N_9692,N_4475,N_273);
or U9693 (N_9693,N_4441,N_2945);
nand U9694 (N_9694,N_2534,N_1091);
nor U9695 (N_9695,N_4698,N_2391);
nor U9696 (N_9696,N_1813,N_3257);
nor U9697 (N_9697,N_2367,N_1465);
nand U9698 (N_9698,N_3430,N_964);
nor U9699 (N_9699,N_715,N_1929);
and U9700 (N_9700,N_2027,N_2279);
nor U9701 (N_9701,N_3944,N_2609);
and U9702 (N_9702,N_2732,N_4214);
nand U9703 (N_9703,N_61,N_1762);
and U9704 (N_9704,N_3331,N_1763);
nand U9705 (N_9705,N_2034,N_2634);
and U9706 (N_9706,N_4355,N_3361);
and U9707 (N_9707,N_4501,N_3820);
and U9708 (N_9708,N_1549,N_1473);
or U9709 (N_9709,N_3945,N_3787);
nand U9710 (N_9710,N_4261,N_4992);
or U9711 (N_9711,N_468,N_1797);
nor U9712 (N_9712,N_4579,N_2529);
or U9713 (N_9713,N_3211,N_756);
and U9714 (N_9714,N_3558,N_3906);
and U9715 (N_9715,N_4994,N_4577);
nand U9716 (N_9716,N_2712,N_1327);
and U9717 (N_9717,N_3785,N_4251);
nand U9718 (N_9718,N_4627,N_4608);
nor U9719 (N_9719,N_1200,N_3716);
nand U9720 (N_9720,N_4562,N_2910);
nor U9721 (N_9721,N_727,N_174);
nor U9722 (N_9722,N_2112,N_4);
nand U9723 (N_9723,N_75,N_576);
or U9724 (N_9724,N_35,N_3862);
nand U9725 (N_9725,N_4760,N_4101);
and U9726 (N_9726,N_2805,N_463);
nand U9727 (N_9727,N_675,N_1329);
or U9728 (N_9728,N_811,N_708);
nand U9729 (N_9729,N_4283,N_1524);
or U9730 (N_9730,N_991,N_104);
nand U9731 (N_9731,N_1352,N_1782);
and U9732 (N_9732,N_823,N_4661);
nand U9733 (N_9733,N_768,N_4684);
nand U9734 (N_9734,N_1148,N_2909);
nand U9735 (N_9735,N_2187,N_1761);
nor U9736 (N_9736,N_1168,N_4756);
and U9737 (N_9737,N_2936,N_2038);
and U9738 (N_9738,N_2968,N_2448);
nor U9739 (N_9739,N_858,N_481);
and U9740 (N_9740,N_2887,N_3974);
or U9741 (N_9741,N_4873,N_1709);
nor U9742 (N_9742,N_1303,N_4848);
nor U9743 (N_9743,N_2028,N_2632);
nand U9744 (N_9744,N_1391,N_2461);
or U9745 (N_9745,N_1278,N_4599);
or U9746 (N_9746,N_4031,N_2191);
nor U9747 (N_9747,N_1173,N_2734);
or U9748 (N_9748,N_1165,N_3166);
nand U9749 (N_9749,N_4522,N_2024);
nand U9750 (N_9750,N_2473,N_2395);
and U9751 (N_9751,N_413,N_751);
or U9752 (N_9752,N_2449,N_3730);
or U9753 (N_9753,N_4522,N_2341);
or U9754 (N_9754,N_4471,N_720);
or U9755 (N_9755,N_956,N_3207);
nand U9756 (N_9756,N_4480,N_790);
nand U9757 (N_9757,N_4146,N_538);
or U9758 (N_9758,N_2853,N_3263);
nand U9759 (N_9759,N_2738,N_2010);
and U9760 (N_9760,N_2248,N_1509);
or U9761 (N_9761,N_2502,N_2956);
and U9762 (N_9762,N_1930,N_1093);
nor U9763 (N_9763,N_3485,N_4986);
nor U9764 (N_9764,N_2800,N_4639);
nor U9765 (N_9765,N_2835,N_117);
nor U9766 (N_9766,N_2860,N_1272);
nor U9767 (N_9767,N_1185,N_2667);
or U9768 (N_9768,N_4574,N_1067);
or U9769 (N_9769,N_2307,N_2250);
nand U9770 (N_9770,N_2498,N_1783);
or U9771 (N_9771,N_3187,N_2661);
nor U9772 (N_9772,N_3497,N_966);
or U9773 (N_9773,N_2652,N_4115);
nand U9774 (N_9774,N_3075,N_3694);
and U9775 (N_9775,N_1022,N_3346);
nand U9776 (N_9776,N_4356,N_3948);
nor U9777 (N_9777,N_4225,N_3089);
nor U9778 (N_9778,N_1182,N_4670);
and U9779 (N_9779,N_729,N_1454);
and U9780 (N_9780,N_3040,N_4077);
and U9781 (N_9781,N_963,N_1351);
or U9782 (N_9782,N_4676,N_3352);
nor U9783 (N_9783,N_2297,N_4594);
nor U9784 (N_9784,N_1570,N_3874);
nand U9785 (N_9785,N_2973,N_3699);
xnor U9786 (N_9786,N_4527,N_2115);
and U9787 (N_9787,N_2421,N_3706);
nand U9788 (N_9788,N_1500,N_3326);
or U9789 (N_9789,N_95,N_487);
or U9790 (N_9790,N_2689,N_4870);
or U9791 (N_9791,N_2584,N_1255);
nand U9792 (N_9792,N_705,N_2852);
or U9793 (N_9793,N_2291,N_2908);
and U9794 (N_9794,N_1648,N_796);
or U9795 (N_9795,N_1342,N_2860);
or U9796 (N_9796,N_1852,N_4893);
nor U9797 (N_9797,N_519,N_296);
or U9798 (N_9798,N_2638,N_2621);
nor U9799 (N_9799,N_2881,N_4450);
nor U9800 (N_9800,N_3693,N_4244);
or U9801 (N_9801,N_354,N_137);
or U9802 (N_9802,N_1997,N_1574);
and U9803 (N_9803,N_4346,N_3960);
or U9804 (N_9804,N_3710,N_4689);
nand U9805 (N_9805,N_2583,N_1624);
and U9806 (N_9806,N_2489,N_3493);
nor U9807 (N_9807,N_4533,N_2521);
nand U9808 (N_9808,N_1340,N_3323);
and U9809 (N_9809,N_3551,N_798);
nor U9810 (N_9810,N_784,N_3956);
nand U9811 (N_9811,N_3288,N_3982);
or U9812 (N_9812,N_302,N_4415);
nand U9813 (N_9813,N_3633,N_2546);
and U9814 (N_9814,N_2812,N_4117);
and U9815 (N_9815,N_1958,N_1069);
nor U9816 (N_9816,N_3626,N_1954);
nand U9817 (N_9817,N_2461,N_500);
nand U9818 (N_9818,N_1423,N_4580);
nor U9819 (N_9819,N_2220,N_2690);
nor U9820 (N_9820,N_2824,N_3107);
and U9821 (N_9821,N_660,N_3941);
or U9822 (N_9822,N_1372,N_1280);
and U9823 (N_9823,N_2700,N_846);
or U9824 (N_9824,N_1563,N_1616);
nor U9825 (N_9825,N_1771,N_1313);
nor U9826 (N_9826,N_4384,N_4652);
nand U9827 (N_9827,N_1181,N_4538);
and U9828 (N_9828,N_1570,N_3966);
nand U9829 (N_9829,N_2569,N_1401);
nor U9830 (N_9830,N_1429,N_3773);
and U9831 (N_9831,N_4162,N_1022);
nand U9832 (N_9832,N_4586,N_1738);
or U9833 (N_9833,N_805,N_2657);
or U9834 (N_9834,N_2739,N_3448);
nand U9835 (N_9835,N_3182,N_527);
and U9836 (N_9836,N_4314,N_3618);
nor U9837 (N_9837,N_1732,N_3408);
and U9838 (N_9838,N_163,N_3862);
nand U9839 (N_9839,N_3723,N_4242);
nor U9840 (N_9840,N_4002,N_4128);
nor U9841 (N_9841,N_4408,N_3477);
or U9842 (N_9842,N_1599,N_1022);
nand U9843 (N_9843,N_1258,N_4847);
nor U9844 (N_9844,N_1479,N_2708);
nand U9845 (N_9845,N_649,N_4101);
or U9846 (N_9846,N_2708,N_3246);
or U9847 (N_9847,N_224,N_3727);
nand U9848 (N_9848,N_3947,N_1647);
nand U9849 (N_9849,N_3801,N_3001);
or U9850 (N_9850,N_4800,N_4620);
nand U9851 (N_9851,N_2544,N_3494);
or U9852 (N_9852,N_3512,N_3845);
nor U9853 (N_9853,N_2506,N_2084);
nor U9854 (N_9854,N_777,N_365);
nand U9855 (N_9855,N_1671,N_4236);
or U9856 (N_9856,N_1200,N_2277);
nand U9857 (N_9857,N_3410,N_456);
or U9858 (N_9858,N_3748,N_4166);
nand U9859 (N_9859,N_2783,N_2449);
or U9860 (N_9860,N_3921,N_2020);
nand U9861 (N_9861,N_4180,N_4040);
and U9862 (N_9862,N_3282,N_2613);
or U9863 (N_9863,N_1093,N_1503);
and U9864 (N_9864,N_576,N_4767);
or U9865 (N_9865,N_416,N_221);
nand U9866 (N_9866,N_4735,N_2911);
nor U9867 (N_9867,N_2464,N_4046);
and U9868 (N_9868,N_3398,N_4973);
and U9869 (N_9869,N_1554,N_1129);
or U9870 (N_9870,N_491,N_400);
nor U9871 (N_9871,N_4782,N_3437);
and U9872 (N_9872,N_2625,N_4856);
nor U9873 (N_9873,N_726,N_796);
nor U9874 (N_9874,N_4269,N_1384);
nand U9875 (N_9875,N_3463,N_4794);
and U9876 (N_9876,N_859,N_3627);
or U9877 (N_9877,N_4564,N_2192);
nand U9878 (N_9878,N_67,N_551);
and U9879 (N_9879,N_2332,N_3544);
and U9880 (N_9880,N_4964,N_3551);
or U9881 (N_9881,N_3126,N_1438);
nor U9882 (N_9882,N_4492,N_1926);
or U9883 (N_9883,N_168,N_101);
and U9884 (N_9884,N_1267,N_228);
nand U9885 (N_9885,N_474,N_4231);
or U9886 (N_9886,N_202,N_139);
and U9887 (N_9887,N_1495,N_125);
and U9888 (N_9888,N_3164,N_4117);
or U9889 (N_9889,N_1600,N_2733);
and U9890 (N_9890,N_963,N_2057);
nor U9891 (N_9891,N_602,N_2362);
nand U9892 (N_9892,N_3267,N_1214);
or U9893 (N_9893,N_634,N_3701);
nand U9894 (N_9894,N_2892,N_4396);
xor U9895 (N_9895,N_2657,N_1102);
nand U9896 (N_9896,N_3,N_3169);
nor U9897 (N_9897,N_4665,N_3878);
nand U9898 (N_9898,N_4572,N_2047);
and U9899 (N_9899,N_4829,N_3562);
and U9900 (N_9900,N_2169,N_195);
and U9901 (N_9901,N_1970,N_2736);
nand U9902 (N_9902,N_2081,N_602);
nand U9903 (N_9903,N_424,N_4146);
and U9904 (N_9904,N_4317,N_1429);
and U9905 (N_9905,N_3994,N_339);
nand U9906 (N_9906,N_1822,N_2993);
and U9907 (N_9907,N_2402,N_1691);
nand U9908 (N_9908,N_1438,N_2080);
or U9909 (N_9909,N_1889,N_4733);
and U9910 (N_9910,N_715,N_4300);
or U9911 (N_9911,N_4111,N_3709);
nor U9912 (N_9912,N_1821,N_4927);
nand U9913 (N_9913,N_4314,N_4430);
xnor U9914 (N_9914,N_3469,N_864);
or U9915 (N_9915,N_3927,N_2332);
or U9916 (N_9916,N_3594,N_4447);
nand U9917 (N_9917,N_4815,N_1141);
nand U9918 (N_9918,N_1105,N_2110);
nand U9919 (N_9919,N_4115,N_3901);
nor U9920 (N_9920,N_3207,N_3773);
nor U9921 (N_9921,N_3287,N_446);
and U9922 (N_9922,N_1338,N_3249);
nor U9923 (N_9923,N_1735,N_4594);
nand U9924 (N_9924,N_902,N_164);
nor U9925 (N_9925,N_2636,N_4094);
or U9926 (N_9926,N_846,N_4140);
or U9927 (N_9927,N_1657,N_4344);
nand U9928 (N_9928,N_4015,N_4184);
or U9929 (N_9929,N_3788,N_1948);
or U9930 (N_9930,N_2920,N_1149);
and U9931 (N_9931,N_4667,N_2886);
and U9932 (N_9932,N_4581,N_2687);
nand U9933 (N_9933,N_401,N_1977);
nand U9934 (N_9934,N_3101,N_4580);
and U9935 (N_9935,N_3552,N_1580);
and U9936 (N_9936,N_4792,N_3927);
and U9937 (N_9937,N_4460,N_1562);
and U9938 (N_9938,N_2242,N_521);
and U9939 (N_9939,N_52,N_2973);
nor U9940 (N_9940,N_1702,N_1484);
or U9941 (N_9941,N_4909,N_613);
or U9942 (N_9942,N_4752,N_4621);
and U9943 (N_9943,N_4705,N_1688);
nand U9944 (N_9944,N_4529,N_3802);
nand U9945 (N_9945,N_975,N_3067);
nor U9946 (N_9946,N_1008,N_1922);
or U9947 (N_9947,N_2486,N_2442);
and U9948 (N_9948,N_1500,N_4954);
and U9949 (N_9949,N_3525,N_3113);
xnor U9950 (N_9950,N_3780,N_1306);
and U9951 (N_9951,N_1439,N_2995);
nand U9952 (N_9952,N_4862,N_4519);
nor U9953 (N_9953,N_1104,N_1663);
nand U9954 (N_9954,N_3058,N_1945);
and U9955 (N_9955,N_3822,N_953);
or U9956 (N_9956,N_967,N_2728);
nand U9957 (N_9957,N_4056,N_2965);
nand U9958 (N_9958,N_55,N_2865);
nand U9959 (N_9959,N_4905,N_1451);
and U9960 (N_9960,N_653,N_3133);
nand U9961 (N_9961,N_1935,N_178);
or U9962 (N_9962,N_4033,N_4010);
or U9963 (N_9963,N_2585,N_2122);
and U9964 (N_9964,N_1685,N_4648);
or U9965 (N_9965,N_4439,N_4151);
nor U9966 (N_9966,N_3343,N_4853);
nand U9967 (N_9967,N_4862,N_1318);
and U9968 (N_9968,N_1331,N_4142);
or U9969 (N_9969,N_1468,N_4609);
nor U9970 (N_9970,N_2657,N_196);
or U9971 (N_9971,N_2189,N_4540);
and U9972 (N_9972,N_2499,N_705);
nand U9973 (N_9973,N_4929,N_1013);
and U9974 (N_9974,N_3822,N_4100);
nor U9975 (N_9975,N_4053,N_2154);
and U9976 (N_9976,N_4109,N_1900);
or U9977 (N_9977,N_4413,N_1018);
and U9978 (N_9978,N_2855,N_1777);
nand U9979 (N_9979,N_161,N_2963);
and U9980 (N_9980,N_2841,N_3811);
or U9981 (N_9981,N_4368,N_4620);
and U9982 (N_9982,N_1305,N_546);
and U9983 (N_9983,N_3488,N_4127);
and U9984 (N_9984,N_2753,N_2561);
and U9985 (N_9985,N_2185,N_86);
and U9986 (N_9986,N_2063,N_4658);
nor U9987 (N_9987,N_2114,N_514);
and U9988 (N_9988,N_3675,N_2482);
nor U9989 (N_9989,N_698,N_3602);
nor U9990 (N_9990,N_1539,N_3431);
and U9991 (N_9991,N_2147,N_987);
or U9992 (N_9992,N_2222,N_771);
and U9993 (N_9993,N_2312,N_4804);
and U9994 (N_9994,N_1664,N_577);
nor U9995 (N_9995,N_38,N_4365);
or U9996 (N_9996,N_45,N_3181);
and U9997 (N_9997,N_2138,N_21);
or U9998 (N_9998,N_3311,N_1250);
nand U9999 (N_9999,N_1089,N_414);
nor UO_0 (O_0,N_5799,N_6350);
and UO_1 (O_1,N_7551,N_9971);
nor UO_2 (O_2,N_6052,N_6875);
and UO_3 (O_3,N_9385,N_7675);
or UO_4 (O_4,N_7809,N_7371);
or UO_5 (O_5,N_6623,N_7729);
and UO_6 (O_6,N_9561,N_5700);
or UO_7 (O_7,N_6202,N_6323);
or UO_8 (O_8,N_9168,N_8515);
or UO_9 (O_9,N_5308,N_9607);
or UO_10 (O_10,N_9728,N_8941);
and UO_11 (O_11,N_7475,N_6830);
and UO_12 (O_12,N_6771,N_9225);
and UO_13 (O_13,N_9835,N_5552);
nand UO_14 (O_14,N_9635,N_8457);
nand UO_15 (O_15,N_7394,N_8434);
or UO_16 (O_16,N_7701,N_9141);
or UO_17 (O_17,N_5256,N_5759);
and UO_18 (O_18,N_8275,N_9642);
and UO_19 (O_19,N_9364,N_6157);
xor UO_20 (O_20,N_5020,N_6755);
nor UO_21 (O_21,N_6048,N_9548);
nor UO_22 (O_22,N_6769,N_7965);
nor UO_23 (O_23,N_7757,N_6540);
or UO_24 (O_24,N_8242,N_7251);
nor UO_25 (O_25,N_6774,N_5939);
and UO_26 (O_26,N_9263,N_9568);
nand UO_27 (O_27,N_5890,N_8176);
and UO_28 (O_28,N_7610,N_5584);
nor UO_29 (O_29,N_7092,N_9019);
and UO_30 (O_30,N_7973,N_9818);
nor UO_31 (O_31,N_6096,N_5068);
nor UO_32 (O_32,N_8088,N_7918);
xnor UO_33 (O_33,N_9485,N_7863);
and UO_34 (O_34,N_8148,N_7119);
or UO_35 (O_35,N_8637,N_7196);
nor UO_36 (O_36,N_8603,N_9554);
and UO_37 (O_37,N_9703,N_7690);
nor UO_38 (O_38,N_5972,N_7299);
nor UO_39 (O_39,N_6666,N_9391);
and UO_40 (O_40,N_8917,N_5781);
nand UO_41 (O_41,N_5875,N_6185);
nand UO_42 (O_42,N_8036,N_5475);
or UO_43 (O_43,N_6225,N_6715);
or UO_44 (O_44,N_8154,N_5187);
nand UO_45 (O_45,N_8921,N_9411);
nor UO_46 (O_46,N_8808,N_9220);
nor UO_47 (O_47,N_8943,N_6616);
nand UO_48 (O_48,N_8774,N_6186);
nand UO_49 (O_49,N_5124,N_5049);
or UO_50 (O_50,N_7012,N_9575);
and UO_51 (O_51,N_9000,N_7262);
nor UO_52 (O_52,N_9080,N_8200);
nand UO_53 (O_53,N_7031,N_5931);
or UO_54 (O_54,N_9005,N_9545);
nand UO_55 (O_55,N_9434,N_7400);
or UO_56 (O_56,N_7426,N_9377);
nor UO_57 (O_57,N_6878,N_9456);
or UO_58 (O_58,N_9161,N_7883);
nor UO_59 (O_59,N_9265,N_7068);
nand UO_60 (O_60,N_9597,N_8219);
nand UO_61 (O_61,N_9394,N_5166);
nor UO_62 (O_62,N_6823,N_7503);
and UO_63 (O_63,N_9400,N_8567);
nor UO_64 (O_64,N_5328,N_6836);
or UO_65 (O_65,N_6832,N_5871);
or UO_66 (O_66,N_7111,N_5226);
and UO_67 (O_67,N_5311,N_7354);
nand UO_68 (O_68,N_6377,N_9251);
or UO_69 (O_69,N_9665,N_7167);
and UO_70 (O_70,N_5095,N_5568);
nor UO_71 (O_71,N_8588,N_7615);
nor UO_72 (O_72,N_7294,N_8650);
and UO_73 (O_73,N_5180,N_8288);
and UO_74 (O_74,N_9913,N_5488);
nand UO_75 (O_75,N_5908,N_9882);
nand UO_76 (O_76,N_6608,N_6498);
or UO_77 (O_77,N_7810,N_5326);
nand UO_78 (O_78,N_8549,N_8656);
nor UO_79 (O_79,N_8764,N_6217);
nor UO_80 (O_80,N_8475,N_5697);
xnor UO_81 (O_81,N_6314,N_9224);
and UO_82 (O_82,N_7137,N_5899);
nor UO_83 (O_83,N_9738,N_8502);
and UO_84 (O_84,N_9431,N_5783);
or UO_85 (O_85,N_5719,N_5537);
or UO_86 (O_86,N_8957,N_8124);
and UO_87 (O_87,N_8987,N_7363);
and UO_88 (O_88,N_8198,N_8407);
and UO_89 (O_89,N_5796,N_8352);
nand UO_90 (O_90,N_6733,N_8900);
or UO_91 (O_91,N_7289,N_9062);
and UO_92 (O_92,N_5404,N_7380);
nand UO_93 (O_93,N_5075,N_7680);
or UO_94 (O_94,N_7901,N_8938);
and UO_95 (O_95,N_5852,N_8508);
nand UO_96 (O_96,N_5137,N_9743);
nor UO_97 (O_97,N_5248,N_7813);
nor UO_98 (O_98,N_9766,N_5986);
nor UO_99 (O_99,N_7310,N_9172);
and UO_100 (O_100,N_9550,N_8130);
or UO_101 (O_101,N_8117,N_8417);
nor UO_102 (O_102,N_7469,N_6238);
or UO_103 (O_103,N_6512,N_8296);
or UO_104 (O_104,N_5818,N_9118);
nor UO_105 (O_105,N_9292,N_5817);
nor UO_106 (O_106,N_8185,N_8826);
or UO_107 (O_107,N_5310,N_7976);
and UO_108 (O_108,N_6971,N_8641);
or UO_109 (O_109,N_9582,N_6164);
or UO_110 (O_110,N_7959,N_5678);
nor UO_111 (O_111,N_6353,N_5793);
or UO_112 (O_112,N_8918,N_9345);
nand UO_113 (O_113,N_8876,N_8583);
nor UO_114 (O_114,N_7742,N_5748);
nand UO_115 (O_115,N_7211,N_9159);
or UO_116 (O_116,N_8793,N_9775);
and UO_117 (O_117,N_9557,N_6452);
nand UO_118 (O_118,N_5619,N_5073);
or UO_119 (O_119,N_7879,N_9793);
nand UO_120 (O_120,N_6806,N_5634);
or UO_121 (O_121,N_7819,N_6169);
nand UO_122 (O_122,N_6459,N_6642);
or UO_123 (O_123,N_5699,N_5520);
or UO_124 (O_124,N_5878,N_7288);
nor UO_125 (O_125,N_7109,N_5048);
or UO_126 (O_126,N_6975,N_6473);
and UO_127 (O_127,N_9869,N_9537);
nor UO_128 (O_128,N_7279,N_6299);
or UO_129 (O_129,N_7921,N_9008);
or UO_130 (O_130,N_5622,N_9380);
nand UO_131 (O_131,N_7632,N_9821);
or UO_132 (O_132,N_7283,N_8230);
or UO_133 (O_133,N_5336,N_6132);
nor UO_134 (O_134,N_9959,N_8360);
nand UO_135 (O_135,N_5128,N_5444);
nor UO_136 (O_136,N_5009,N_8862);
nand UO_137 (O_137,N_6927,N_9951);
nor UO_138 (O_138,N_6248,N_9382);
and UO_139 (O_139,N_6092,N_7145);
nor UO_140 (O_140,N_7158,N_5333);
nand UO_141 (O_141,N_5195,N_7315);
and UO_142 (O_142,N_7892,N_7273);
and UO_143 (O_143,N_7596,N_7055);
nand UO_144 (O_144,N_7751,N_7466);
nor UO_145 (O_145,N_9235,N_8218);
nand UO_146 (O_146,N_8971,N_7062);
nor UO_147 (O_147,N_5578,N_7923);
or UO_148 (O_148,N_5366,N_9718);
and UO_149 (O_149,N_5795,N_7834);
and UO_150 (O_150,N_7799,N_9799);
or UO_151 (O_151,N_7606,N_7091);
nor UO_152 (O_152,N_7613,N_7874);
and UO_153 (O_153,N_5111,N_9095);
or UO_154 (O_154,N_5162,N_9916);
or UO_155 (O_155,N_9152,N_7491);
nor UO_156 (O_156,N_6308,N_5081);
nor UO_157 (O_157,N_8333,N_6680);
and UO_158 (O_158,N_9305,N_9993);
or UO_159 (O_159,N_5811,N_7847);
nand UO_160 (O_160,N_6589,N_5470);
nor UO_161 (O_161,N_8150,N_8528);
xor UO_162 (O_162,N_9867,N_9603);
or UO_163 (O_163,N_5865,N_7731);
nand UO_164 (O_164,N_9343,N_6790);
or UO_165 (O_165,N_6862,N_9990);
nand UO_166 (O_166,N_6604,N_9052);
and UO_167 (O_167,N_5508,N_8506);
and UO_168 (O_168,N_5561,N_9237);
nor UO_169 (O_169,N_9591,N_6824);
or UO_170 (O_170,N_5988,N_5624);
nand UO_171 (O_171,N_7479,N_7552);
nor UO_172 (O_172,N_9170,N_7090);
nor UO_173 (O_173,N_8949,N_7467);
and UO_174 (O_174,N_8817,N_8536);
and UO_175 (O_175,N_5181,N_9158);
or UO_176 (O_176,N_9074,N_7908);
nor UO_177 (O_177,N_6649,N_8960);
nand UO_178 (O_178,N_8510,N_6874);
nor UO_179 (O_179,N_5215,N_6326);
nand UO_180 (O_180,N_8615,N_8159);
or UO_181 (O_181,N_9525,N_9216);
nor UO_182 (O_182,N_8480,N_5178);
or UO_183 (O_183,N_7540,N_6112);
nand UO_184 (O_184,N_9218,N_6573);
and UO_185 (O_185,N_7318,N_8944);
nor UO_186 (O_186,N_6659,N_6732);
nor UO_187 (O_187,N_5758,N_7697);
or UO_188 (O_188,N_6490,N_6599);
or UO_189 (O_189,N_9488,N_7647);
nor UO_190 (O_190,N_6841,N_6791);
or UO_191 (O_191,N_9767,N_8035);
nor UO_192 (O_192,N_7766,N_9192);
or UO_193 (O_193,N_9994,N_5260);
nand UO_194 (O_194,N_7313,N_8334);
and UO_195 (O_195,N_6670,N_8748);
nand UO_196 (O_196,N_5625,N_7325);
nand UO_197 (O_197,N_8893,N_7465);
nand UO_198 (O_198,N_9397,N_7391);
nor UO_199 (O_199,N_8369,N_5567);
and UO_200 (O_200,N_6779,N_6190);
and UO_201 (O_201,N_6201,N_5421);
or UO_202 (O_202,N_9694,N_6356);
and UO_203 (O_203,N_5966,N_9533);
nand UO_204 (O_204,N_9330,N_8365);
nor UO_205 (O_205,N_7024,N_6433);
nor UO_206 (O_206,N_9198,N_6968);
and UO_207 (O_207,N_5347,N_9670);
and UO_208 (O_208,N_6244,N_6006);
nand UO_209 (O_209,N_9909,N_9287);
xnor UO_210 (O_210,N_8871,N_5098);
or UO_211 (O_211,N_9925,N_5126);
and UO_212 (O_212,N_5600,N_9090);
and UO_213 (O_213,N_7602,N_6800);
and UO_214 (O_214,N_5167,N_7468);
or UO_215 (O_215,N_9478,N_8073);
or UO_216 (O_216,N_6198,N_6026);
nand UO_217 (O_217,N_8595,N_7507);
nand UO_218 (O_218,N_9073,N_6767);
nor UO_219 (O_219,N_8857,N_7032);
and UO_220 (O_220,N_8736,N_5892);
or UO_221 (O_221,N_5635,N_9070);
nor UO_222 (O_222,N_6815,N_6517);
or UO_223 (O_223,N_5924,N_8520);
nand UO_224 (O_224,N_5206,N_6943);
or UO_225 (O_225,N_5334,N_6691);
and UO_226 (O_226,N_7240,N_5712);
and UO_227 (O_227,N_8580,N_5742);
nand UO_228 (O_228,N_8666,N_9915);
and UO_229 (O_229,N_9529,N_7800);
or UO_230 (O_230,N_6332,N_9418);
nand UO_231 (O_231,N_7352,N_8682);
and UO_232 (O_232,N_7036,N_5636);
or UO_233 (O_233,N_8497,N_5249);
and UO_234 (O_234,N_9658,N_9458);
or UO_235 (O_235,N_5094,N_9693);
nand UO_236 (O_236,N_6355,N_6120);
and UO_237 (O_237,N_6453,N_5405);
nand UO_238 (O_238,N_6743,N_6863);
nor UO_239 (O_239,N_5063,N_7726);
nor UO_240 (O_240,N_8694,N_9185);
or UO_241 (O_241,N_7624,N_8695);
or UO_242 (O_242,N_8988,N_5918);
or UO_243 (O_243,N_8420,N_9262);
or UO_244 (O_244,N_9029,N_5299);
and UO_245 (O_245,N_6482,N_7378);
nor UO_246 (O_246,N_7108,N_6828);
nand UO_247 (O_247,N_5343,N_7987);
nor UO_248 (O_248,N_7823,N_6899);
or UO_249 (O_249,N_8181,N_9716);
nand UO_250 (O_250,N_6457,N_6711);
or UO_251 (O_251,N_5529,N_5663);
nor UO_252 (O_252,N_8783,N_9715);
nor UO_253 (O_253,N_9276,N_8904);
and UO_254 (O_254,N_9247,N_7141);
nor UO_255 (O_255,N_6402,N_5264);
or UO_256 (O_256,N_9810,N_9891);
nor UO_257 (O_257,N_7360,N_6097);
or UO_258 (O_258,N_5403,N_7687);
nand UO_259 (O_259,N_6034,N_7260);
or UO_260 (O_260,N_6851,N_6362);
or UO_261 (O_261,N_8735,N_9641);
and UO_262 (O_262,N_5109,N_8912);
nand UO_263 (O_263,N_6083,N_6414);
or UO_264 (O_264,N_9519,N_9827);
or UO_265 (O_265,N_5282,N_8192);
and UO_266 (O_266,N_8493,N_8787);
and UO_267 (O_267,N_7753,N_5516);
nand UO_268 (O_268,N_6010,N_8687);
nand UO_269 (O_269,N_5024,N_9307);
and UO_270 (O_270,N_6989,N_8439);
nor UO_271 (O_271,N_8894,N_7885);
or UO_272 (O_272,N_6208,N_6763);
and UO_273 (O_273,N_5630,N_6384);
and UO_274 (O_274,N_5518,N_6565);
nor UO_275 (O_275,N_9874,N_9469);
and UO_276 (O_276,N_6619,N_7773);
and UO_277 (O_277,N_9174,N_8274);
or UO_278 (O_278,N_7180,N_7193);
and UO_279 (O_279,N_6893,N_8956);
nand UO_280 (O_280,N_5581,N_7236);
nand UO_281 (O_281,N_9864,N_8413);
or UO_282 (O_282,N_8010,N_7367);
nor UO_283 (O_283,N_8916,N_9296);
and UO_284 (O_284,N_9893,N_6984);
and UO_285 (O_285,N_5455,N_6243);
nor UO_286 (O_286,N_5410,N_9416);
and UO_287 (O_287,N_9309,N_5459);
nor UO_288 (O_288,N_6489,N_6954);
and UO_289 (O_289,N_5116,N_6627);
xnor UO_290 (O_290,N_7539,N_6741);
or UO_291 (O_291,N_9457,N_6122);
nor UO_292 (O_292,N_9843,N_6955);
or UO_293 (O_293,N_6161,N_6204);
nor UO_294 (O_294,N_8705,N_6579);
or UO_295 (O_295,N_6389,N_6896);
xnor UO_296 (O_296,N_8098,N_5042);
and UO_297 (O_297,N_8671,N_8196);
nand UO_298 (O_298,N_6015,N_5684);
nand UO_299 (O_299,N_9917,N_6031);
or UO_300 (O_300,N_7375,N_5609);
or UO_301 (O_301,N_6653,N_8831);
nor UO_302 (O_302,N_5373,N_7239);
and UO_303 (O_303,N_6068,N_7326);
nand UO_304 (O_304,N_6979,N_8527);
nand UO_305 (O_305,N_8039,N_5956);
and UO_306 (O_306,N_9183,N_6150);
and UO_307 (O_307,N_9369,N_8610);
and UO_308 (O_308,N_9816,N_6563);
or UO_309 (O_309,N_5493,N_8855);
or UO_310 (O_310,N_6193,N_6658);
nand UO_311 (O_311,N_8819,N_7870);
nand UO_312 (O_312,N_5669,N_7622);
nand UO_313 (O_313,N_7725,N_5171);
and UO_314 (O_314,N_6842,N_6032);
and UO_315 (O_315,N_6839,N_7616);
nand UO_316 (O_316,N_9765,N_9892);
or UO_317 (O_317,N_9717,N_6812);
nand UO_318 (O_318,N_6966,N_8560);
nand UO_319 (O_319,N_9374,N_9509);
or UO_320 (O_320,N_9272,N_7027);
nor UO_321 (O_321,N_7314,N_7774);
and UO_322 (O_322,N_5093,N_6641);
nor UO_323 (O_323,N_5453,N_9619);
nand UO_324 (O_324,N_5790,N_9534);
and UO_325 (O_325,N_5353,N_5190);
and UO_326 (O_326,N_9813,N_7078);
or UO_327 (O_327,N_7089,N_5262);
and UO_328 (O_328,N_7424,N_6182);
nor UO_329 (O_329,N_6757,N_6873);
nor UO_330 (O_330,N_5363,N_8491);
or UO_331 (O_331,N_5787,N_7714);
nand UO_332 (O_332,N_5329,N_5268);
or UO_333 (O_333,N_8645,N_7328);
nor UO_334 (O_334,N_9249,N_9792);
or UO_335 (O_335,N_8699,N_9884);
xnor UO_336 (O_336,N_9371,N_6534);
nor UO_337 (O_337,N_5968,N_9671);
or UO_338 (O_338,N_7286,N_9280);
nor UO_339 (O_339,N_6156,N_8727);
and UO_340 (O_340,N_8608,N_7496);
nand UO_341 (O_341,N_5200,N_6557);
nand UO_342 (O_342,N_6148,N_9521);
or UO_343 (O_343,N_7338,N_9201);
and UO_344 (O_344,N_9967,N_9678);
and UO_345 (O_345,N_9868,N_8553);
nand UO_346 (O_346,N_7607,N_8220);
nand UO_347 (O_347,N_8953,N_7020);
nor UO_348 (O_348,N_5885,N_6365);
nor UO_349 (O_349,N_6539,N_7112);
and UO_350 (O_350,N_9675,N_6087);
nand UO_351 (O_351,N_6992,N_6008);
and UO_352 (O_352,N_5204,N_9559);
or UO_353 (O_353,N_5577,N_5140);
and UO_354 (O_354,N_9099,N_7430);
nor UO_355 (O_355,N_8072,N_8366);
or UO_356 (O_356,N_6417,N_9384);
nor UO_357 (O_357,N_6478,N_8753);
nor UO_358 (O_358,N_5154,N_7826);
and UO_359 (O_359,N_7249,N_8972);
and UO_360 (O_360,N_6591,N_5036);
or UO_361 (O_361,N_9236,N_6716);
and UO_362 (O_362,N_8193,N_8326);
nand UO_363 (O_363,N_5134,N_9511);
nand UO_364 (O_364,N_8643,N_6380);
nor UO_365 (O_365,N_8305,N_8101);
or UO_366 (O_366,N_9025,N_6892);
nand UO_367 (O_367,N_8410,N_6569);
nand UO_368 (O_368,N_8054,N_6913);
nand UO_369 (O_369,N_8488,N_9754);
or UO_370 (O_370,N_7093,N_5431);
nor UO_371 (O_371,N_7254,N_6576);
nor UO_372 (O_372,N_9204,N_8759);
or UO_373 (O_373,N_9341,N_6342);
nand UO_374 (O_374,N_7347,N_6798);
and UO_375 (O_375,N_9549,N_7135);
nand UO_376 (O_376,N_8964,N_6094);
and UO_377 (O_377,N_9245,N_7985);
nand UO_378 (O_378,N_9282,N_7345);
xor UO_379 (O_379,N_9210,N_9209);
nor UO_380 (O_380,N_9072,N_6346);
nand UO_381 (O_381,N_6723,N_9636);
nand UO_382 (O_382,N_5536,N_5653);
nand UO_383 (O_383,N_6814,N_8486);
and UO_384 (O_384,N_6726,N_9285);
and UO_385 (O_385,N_9238,N_9705);
or UO_386 (O_386,N_6639,N_7612);
nor UO_387 (O_387,N_6996,N_6547);
or UO_388 (O_388,N_5779,N_6028);
nand UO_389 (O_389,N_7440,N_5246);
nor UO_390 (O_390,N_7472,N_6970);
or UO_391 (O_391,N_6136,N_9855);
and UO_392 (O_392,N_6797,N_5039);
nand UO_393 (O_393,N_8018,N_7657);
or UO_394 (O_394,N_5957,N_5293);
and UO_395 (O_395,N_8683,N_5125);
xor UO_396 (O_396,N_7603,N_7566);
or UO_397 (O_397,N_8109,N_8359);
nand UO_398 (O_398,N_7197,N_6536);
and UO_399 (O_399,N_5951,N_6153);
nor UO_400 (O_400,N_8848,N_6066);
and UO_401 (O_401,N_9100,N_8235);
and UO_402 (O_402,N_5047,N_8037);
nor UO_403 (O_403,N_7419,N_8057);
or UO_404 (O_404,N_7179,N_8380);
nand UO_405 (O_405,N_8702,N_5621);
or UO_406 (O_406,N_7428,N_7006);
nor UO_407 (O_407,N_8886,N_6110);
or UO_408 (O_408,N_8696,N_5244);
nor UO_409 (O_409,N_9190,N_8370);
nand UO_410 (O_410,N_7735,N_6251);
and UO_411 (O_411,N_5917,N_9217);
and UO_412 (O_412,N_7134,N_7629);
or UO_413 (O_413,N_8328,N_8089);
nand UO_414 (O_414,N_5524,N_9448);
or UO_415 (O_415,N_7098,N_9450);
or UO_416 (O_416,N_8128,N_8199);
and UO_417 (O_417,N_8224,N_8986);
nand UO_418 (O_418,N_7490,N_6415);
nor UO_419 (O_419,N_8276,N_7917);
and UO_420 (O_420,N_9667,N_5370);
nor UO_421 (O_421,N_6451,N_6631);
nor UO_422 (O_422,N_9232,N_6784);
and UO_423 (O_423,N_5550,N_9598);
and UO_424 (O_424,N_7295,N_8090);
nor UO_425 (O_425,N_9023,N_9535);
or UO_426 (O_426,N_7831,N_8070);
nor UO_427 (O_427,N_9009,N_9791);
nor UO_428 (O_428,N_9298,N_6191);
or UO_429 (O_429,N_9975,N_5401);
or UO_430 (O_430,N_5396,N_9358);
and UO_431 (O_431,N_6376,N_8190);
and UO_432 (O_432,N_6597,N_5915);
nor UO_433 (O_433,N_5191,N_6213);
or UO_434 (O_434,N_7999,N_8494);
and UO_435 (O_435,N_5977,N_5659);
or UO_436 (O_436,N_6124,N_7225);
or UO_437 (O_437,N_9252,N_8290);
nand UO_438 (O_438,N_6152,N_6129);
or UO_439 (O_439,N_7455,N_7206);
nor UO_440 (O_440,N_5618,N_5671);
and UO_441 (O_441,N_9423,N_9068);
nor UO_442 (O_442,N_7063,N_8909);
nor UO_443 (O_443,N_7480,N_8168);
nor UO_444 (O_444,N_5617,N_8183);
nor UO_445 (O_445,N_9101,N_6834);
and UO_446 (O_446,N_5598,N_5732);
nor UO_447 (O_447,N_5880,N_8788);
and UO_448 (O_448,N_9886,N_9699);
nand UO_449 (O_449,N_5668,N_5836);
nor UO_450 (O_450,N_5954,N_9605);
nor UO_451 (O_451,N_5743,N_6681);
nand UO_452 (O_452,N_5973,N_5005);
nor UO_453 (O_453,N_5948,N_7410);
nor UO_454 (O_454,N_6777,N_5008);
or UO_455 (O_455,N_7848,N_5198);
nand UO_456 (O_456,N_6025,N_7961);
or UO_457 (O_457,N_9383,N_6261);
nor UO_458 (O_458,N_9178,N_8464);
and UO_459 (O_459,N_7601,N_6170);
or UO_460 (O_460,N_9196,N_6808);
nand UO_461 (O_461,N_7221,N_8983);
nand UO_462 (O_462,N_8042,N_8362);
nand UO_463 (O_463,N_9091,N_8709);
or UO_464 (O_464,N_6949,N_8279);
or UO_465 (O_465,N_9077,N_5319);
and UO_466 (O_466,N_8927,N_5295);
xnor UO_467 (O_467,N_8299,N_6590);
nor UO_468 (O_468,N_7530,N_8593);
and UO_469 (O_469,N_9121,N_6381);
or UO_470 (O_470,N_7038,N_5057);
nand UO_471 (O_471,N_5704,N_8066);
nand UO_472 (O_472,N_8952,N_7693);
and UO_473 (O_473,N_7872,N_7948);
or UO_474 (O_474,N_8737,N_9965);
or UO_475 (O_475,N_5067,N_5970);
nor UO_476 (O_476,N_8127,N_6125);
nor UO_477 (O_477,N_9854,N_5656);
and UO_478 (O_478,N_9887,N_6656);
or UO_479 (O_479,N_9257,N_5883);
or UO_480 (O_480,N_5504,N_8845);
or UO_481 (O_481,N_6479,N_7264);
nand UO_482 (O_482,N_5006,N_6937);
nand UO_483 (O_483,N_6080,N_5562);
nand UO_484 (O_484,N_6009,N_8003);
nand UO_485 (O_485,N_7634,N_8357);
nand UO_486 (O_486,N_8264,N_7975);
and UO_487 (O_487,N_6543,N_6281);
and UO_488 (O_488,N_6177,N_8878);
nand UO_489 (O_489,N_8044,N_9471);
nor UO_490 (O_490,N_9093,N_6361);
and UO_491 (O_491,N_6054,N_8306);
nand UO_492 (O_492,N_7658,N_5576);
or UO_493 (O_493,N_5479,N_9815);
nor UO_494 (O_494,N_5448,N_8157);
and UO_495 (O_495,N_7291,N_7505);
nor UO_496 (O_496,N_9833,N_8985);
and UO_497 (O_497,N_6915,N_5253);
and UO_498 (O_498,N_5305,N_6042);
and UO_499 (O_499,N_7296,N_7045);
or UO_500 (O_500,N_9660,N_8445);
nand UO_501 (O_501,N_8040,N_8110);
nor UO_502 (O_502,N_7609,N_6022);
nand UO_503 (O_503,N_7567,N_8206);
and UO_504 (O_504,N_7856,N_9124);
and UO_505 (O_505,N_8269,N_9898);
or UO_506 (O_506,N_6803,N_9013);
or UO_507 (O_507,N_8634,N_6751);
or UO_508 (O_508,N_5202,N_9207);
nand UO_509 (O_509,N_7549,N_6036);
nor UO_510 (O_510,N_8227,N_7761);
and UO_511 (O_511,N_6312,N_5186);
and UO_512 (O_512,N_7889,N_5276);
and UO_513 (O_513,N_9803,N_7502);
and UO_514 (O_514,N_8355,N_8174);
or UO_515 (O_515,N_9714,N_9167);
and UO_516 (O_516,N_9612,N_9147);
nor UO_517 (O_517,N_7248,N_8984);
or UO_518 (O_518,N_5798,N_8460);
nand UO_519 (O_519,N_6718,N_8731);
and UO_520 (O_520,N_7526,N_8739);
or UO_521 (O_521,N_5102,N_8133);
nor UO_522 (O_522,N_9634,N_8842);
or UO_523 (O_523,N_8467,N_5117);
or UO_524 (O_524,N_7233,N_6820);
nor UO_525 (O_525,N_9331,N_9205);
nand UO_526 (O_526,N_6233,N_6371);
nor UO_527 (O_527,N_7172,N_8704);
or UO_528 (O_528,N_5078,N_8249);
and UO_529 (O_529,N_8301,N_8208);
nor UO_530 (O_530,N_9683,N_5105);
or UO_531 (O_531,N_8711,N_5457);
nand UO_532 (O_532,N_8936,N_6272);
or UO_533 (O_533,N_7285,N_7550);
nor UO_534 (O_534,N_8873,N_9691);
and UO_535 (O_535,N_5533,N_7929);
nor UO_536 (O_536,N_7498,N_5233);
nor UO_537 (O_537,N_6861,N_5472);
nand UO_538 (O_538,N_5808,N_6630);
or UO_539 (O_539,N_9365,N_8302);
nor UO_540 (O_540,N_9340,N_9761);
or UO_541 (O_541,N_5112,N_8119);
xnor UO_542 (O_542,N_9284,N_8945);
nand UO_543 (O_543,N_6160,N_5250);
and UO_544 (O_544,N_5823,N_9615);
or UO_545 (O_545,N_5484,N_6252);
nor UO_546 (O_546,N_8513,N_8202);
and UO_547 (O_547,N_7474,N_9175);
or UO_548 (O_548,N_7446,N_7899);
or UO_549 (O_549,N_7334,N_5088);
nand UO_550 (O_550,N_9063,N_9516);
or UO_551 (O_551,N_7591,N_5501);
and UO_552 (O_552,N_9392,N_8253);
nor UO_553 (O_553,N_9297,N_5633);
or UO_554 (O_554,N_6072,N_5344);
and UO_555 (O_555,N_6106,N_7843);
nor UO_556 (O_556,N_8710,N_5129);
and UO_557 (O_557,N_7011,N_9942);
nand UO_558 (O_558,N_7906,N_6840);
nand UO_559 (O_559,N_7708,N_9024);
nand UO_560 (O_560,N_8435,N_5538);
and UO_561 (O_561,N_5553,N_8246);
and UO_562 (O_562,N_7082,N_8005);
nor UO_563 (O_563,N_7348,N_6917);
or UO_564 (O_564,N_5054,N_5950);
nor UO_565 (O_565,N_5423,N_9674);
or UO_566 (O_566,N_9089,N_7662);
nor UO_567 (O_567,N_7035,N_7523);
nor UO_568 (O_568,N_5330,N_7927);
or UO_569 (O_569,N_9313,N_6327);
and UO_570 (O_570,N_6598,N_5407);
and UO_571 (O_571,N_7547,N_9075);
or UO_572 (O_572,N_5587,N_7081);
or UO_573 (O_573,N_7155,N_7064);
and UO_574 (O_574,N_5876,N_7127);
nor UO_575 (O_575,N_6848,N_8391);
nor UO_576 (O_576,N_5751,N_7317);
and UO_577 (O_577,N_7121,N_5820);
nor UO_578 (O_578,N_7633,N_8573);
and UO_579 (O_579,N_7007,N_5913);
or UO_580 (O_580,N_8384,N_5828);
nand UO_581 (O_581,N_8499,N_8555);
and UO_582 (O_582,N_8335,N_5464);
and UO_583 (O_583,N_6168,N_8062);
nand UO_584 (O_584,N_9921,N_6690);
nand UO_585 (O_585,N_8743,N_7942);
and UO_586 (O_586,N_9836,N_7306);
or UO_587 (O_587,N_6867,N_5136);
or UO_588 (O_588,N_5044,N_8382);
and UO_589 (O_589,N_5152,N_9439);
and UO_590 (O_590,N_8525,N_8343);
nor UO_591 (O_591,N_6322,N_8887);
nor UO_592 (O_592,N_6980,N_9896);
nor UO_593 (O_593,N_5051,N_9150);
or UO_594 (O_594,N_7638,N_6089);
and UO_595 (O_595,N_5335,N_7670);
nor UO_596 (O_596,N_6282,N_6293);
and UO_597 (O_597,N_8836,N_6044);
nand UO_598 (O_598,N_9532,N_8273);
xor UO_599 (O_599,N_9398,N_5143);
and UO_600 (O_600,N_9755,N_5211);
or UO_601 (O_601,N_5492,N_8009);
or UO_602 (O_602,N_9290,N_7369);
nand UO_603 (O_603,N_8978,N_5115);
nand UO_604 (O_604,N_9214,N_5971);
nand UO_605 (O_605,N_9333,N_6438);
or UO_606 (O_606,N_5245,N_5728);
and UO_607 (O_607,N_5946,N_9807);
and UO_608 (O_608,N_9149,N_8524);
or UO_609 (O_609,N_8993,N_8315);
and UO_610 (O_610,N_8547,N_6518);
nand UO_611 (O_611,N_5926,N_7003);
nor UO_612 (O_612,N_5733,N_6548);
nor UO_613 (O_613,N_6850,N_9842);
or UO_614 (O_614,N_6101,N_7494);
and UO_615 (O_615,N_9689,N_5938);
or UO_616 (O_616,N_8907,N_7780);
and UO_617 (O_617,N_5978,N_8387);
nor UO_618 (O_618,N_5774,N_5688);
nand UO_619 (O_619,N_9361,N_6249);
and UO_620 (O_620,N_7564,N_6964);
and UO_621 (O_621,N_8823,N_9651);
nand UO_622 (O_622,N_5123,N_9544);
and UO_623 (O_623,N_6626,N_5608);
xnor UO_624 (O_624,N_9289,N_5424);
nor UO_625 (O_625,N_5052,N_6963);
nor UO_626 (O_626,N_7432,N_5043);
and UO_627 (O_627,N_9490,N_8749);
and UO_628 (O_628,N_7794,N_9473);
and UO_629 (O_629,N_5845,N_5070);
and UO_630 (O_630,N_8373,N_7663);
and UO_631 (O_631,N_9031,N_6888);
and UO_632 (O_632,N_6852,N_7896);
nand UO_633 (O_633,N_6057,N_5523);
nor UO_634 (O_634,N_9259,N_6188);
nor UO_635 (O_635,N_5323,N_8222);
nand UO_636 (O_636,N_9740,N_9902);
nand UO_637 (O_637,N_6192,N_5531);
and UO_638 (O_638,N_6321,N_9904);
or UO_639 (O_639,N_9540,N_9536);
or UO_640 (O_640,N_5599,N_7671);
nor UO_641 (O_641,N_9638,N_5217);
and UO_642 (O_642,N_7877,N_6137);
or UO_643 (O_643,N_5682,N_6805);
or UO_644 (O_644,N_6687,N_5369);
and UO_645 (O_645,N_9270,N_8875);
or UO_646 (O_646,N_9437,N_5903);
nand UO_647 (O_647,N_6398,N_5786);
or UO_648 (O_648,N_6688,N_5432);
nand UO_649 (O_649,N_5437,N_8519);
nor UO_650 (O_650,N_5252,N_9066);
nor UO_651 (O_651,N_5119,N_9883);
or UO_652 (O_652,N_6683,N_9584);
nand UO_653 (O_653,N_9798,N_7924);
nand UO_654 (O_654,N_9943,N_7243);
and UO_655 (O_655,N_6462,N_8901);
or UO_656 (O_656,N_9539,N_6650);
nand UO_657 (O_657,N_7350,N_6033);
or UO_658 (O_658,N_7668,N_7459);
nand UO_659 (O_659,N_5565,N_5382);
nand UO_660 (O_660,N_7080,N_7113);
nor UO_661 (O_661,N_5650,N_8587);
nand UO_662 (O_662,N_7548,N_7593);
nand UO_663 (O_663,N_8940,N_5638);
and UO_664 (O_664,N_9961,N_5805);
nor UO_665 (O_665,N_9621,N_8883);
and UO_666 (O_666,N_5602,N_8265);
and UO_667 (O_667,N_9107,N_6684);
nor UO_668 (O_668,N_9659,N_7608);
or UO_669 (O_669,N_9856,N_9517);
or UO_670 (O_670,N_9112,N_7778);
or UO_671 (O_671,N_6702,N_9841);
nand UO_672 (O_672,N_5265,N_8026);
nor UO_673 (O_673,N_7083,N_9640);
and UO_674 (O_674,N_7431,N_8642);
and UO_675 (O_675,N_7255,N_6420);
nand UO_676 (O_676,N_5196,N_6219);
nand UO_677 (O_677,N_9599,N_7815);
or UO_678 (O_678,N_9199,N_6612);
or UO_679 (O_679,N_9753,N_6673);
or UO_680 (O_680,N_5461,N_8071);
or UO_681 (O_681,N_7851,N_8175);
or UO_682 (O_682,N_7739,N_7042);
or UO_683 (O_683,N_6341,N_9241);
xor UO_684 (O_684,N_8461,N_7037);
or UO_685 (O_685,N_9878,N_9769);
and UO_686 (O_686,N_7944,N_7510);
nand UO_687 (O_687,N_9905,N_7246);
or UO_688 (O_688,N_9770,N_8928);
nand UO_689 (O_689,N_8415,N_9645);
and UO_690 (O_690,N_9964,N_5259);
and UO_691 (O_691,N_6894,N_9105);
nor UO_692 (O_692,N_5945,N_8309);
nor UO_693 (O_693,N_9306,N_7344);
nor UO_694 (O_694,N_8981,N_7146);
nor UO_695 (O_695,N_6853,N_9507);
and UO_696 (O_696,N_8838,N_7228);
or UO_697 (O_697,N_7683,N_6047);
nand UO_698 (O_698,N_9056,N_9496);
nor UO_699 (O_699,N_6147,N_7120);
nand UO_700 (O_700,N_6750,N_6005);
or UO_701 (O_701,N_6035,N_5174);
and UO_702 (O_702,N_8780,N_7205);
nor UO_703 (O_703,N_9788,N_6298);
nand UO_704 (O_704,N_7666,N_7881);
or UO_705 (O_705,N_5844,N_5898);
and UO_706 (O_706,N_8910,N_7578);
and UO_707 (O_707,N_7095,N_7327);
nor UO_708 (O_708,N_7880,N_8217);
and UO_709 (O_709,N_6434,N_5646);
and UO_710 (O_710,N_7153,N_9482);
nor UO_711 (O_711,N_6973,N_7640);
or UO_712 (O_712,N_7335,N_8438);
nand UO_713 (O_713,N_7752,N_8933);
nand UO_714 (O_714,N_8679,N_9096);
nand UO_715 (O_715,N_9122,N_5216);
nand UO_716 (O_716,N_6064,N_7054);
and UO_717 (O_717,N_8619,N_7644);
and UO_718 (O_718,N_7835,N_7702);
nand UO_719 (O_719,N_5289,N_9823);
nor UO_720 (O_720,N_5548,N_6635);
or UO_721 (O_721,N_7241,N_7909);
nor UO_722 (O_722,N_8487,N_8742);
or UO_723 (O_723,N_7559,N_8019);
nor UO_724 (O_724,N_5381,N_5866);
nand UO_725 (O_725,N_5960,N_5490);
nand UO_726 (O_726,N_7546,N_5723);
or UO_727 (O_727,N_6477,N_7534);
or UO_728 (O_728,N_7316,N_6102);
or UO_729 (O_729,N_9129,N_5914);
and UO_730 (O_730,N_5270,N_7339);
nor UO_731 (O_731,N_8342,N_8926);
nand UO_732 (O_732,N_7676,N_5439);
and UO_733 (O_733,N_6821,N_8401);
nand UO_734 (O_734,N_8669,N_5554);
nand UO_735 (O_735,N_8451,N_7793);
nand UO_736 (O_736,N_5549,N_8958);
nor UO_737 (O_737,N_6301,N_8250);
and UO_738 (O_738,N_9461,N_9311);
nor UO_739 (O_739,N_5594,N_6532);
or UO_740 (O_740,N_6447,N_9275);
nand UO_741 (O_741,N_6972,N_7140);
and UO_742 (O_742,N_5833,N_9503);
nor UO_743 (O_743,N_6163,N_9433);
or UO_744 (O_744,N_6264,N_5583);
or UO_745 (O_745,N_7405,N_7076);
nand UO_746 (O_746,N_8496,N_6115);
and UO_747 (O_747,N_6255,N_5651);
or UO_748 (O_748,N_6288,N_5929);
or UO_749 (O_749,N_6449,N_8316);
nand UO_750 (O_750,N_8346,N_9593);
nor UO_751 (O_751,N_9502,N_9866);
nand UO_752 (O_752,N_8509,N_8134);
nor UO_753 (O_753,N_6319,N_6925);
nand UO_754 (O_754,N_5367,N_9255);
or UO_755 (O_755,N_9020,N_5050);
and UO_756 (O_756,N_8979,N_5815);
nor UO_757 (O_757,N_8108,N_6969);
nand UO_758 (O_758,N_7955,N_7132);
or UO_759 (O_759,N_5321,N_7801);
and UO_760 (O_760,N_6935,N_5254);
and UO_761 (O_761,N_9223,N_5118);
and UO_762 (O_762,N_8802,N_9162);
nand UO_763 (O_763,N_8621,N_8601);
nor UO_764 (O_764,N_5413,N_5251);
nor UO_765 (O_765,N_6638,N_6811);
and UO_766 (O_766,N_6421,N_6392);
or UO_767 (O_767,N_8162,N_9590);
and UO_768 (O_768,N_7284,N_6118);
nor UO_769 (O_769,N_7575,N_7058);
nand UO_770 (O_770,N_5307,N_5029);
nor UO_771 (O_771,N_8660,N_5711);
nor UO_772 (O_772,N_5976,N_5513);
and UO_773 (O_773,N_5034,N_7178);
nor UO_774 (O_774,N_5615,N_5184);
nor UO_775 (O_775,N_8430,N_8514);
and UO_776 (O_776,N_8446,N_7673);
and UO_777 (O_777,N_7244,N_7520);
nor UO_778 (O_778,N_9560,N_6885);
nor UO_779 (O_779,N_5272,N_6745);
nand UO_780 (O_780,N_5613,N_9650);
nand UO_781 (O_781,N_9945,N_6866);
or UO_782 (O_782,N_7340,N_5629);
or UO_783 (O_783,N_5673,N_7018);
nor UO_784 (O_784,N_8685,N_9937);
nor UO_785 (O_785,N_8568,N_8414);
and UO_786 (O_786,N_6002,N_9900);
nor UO_787 (O_787,N_8006,N_8312);
and UO_788 (O_788,N_7623,N_8495);
nand UO_789 (O_789,N_8550,N_6960);
xor UO_790 (O_790,N_7287,N_5144);
nor UO_791 (O_791,N_6744,N_6708);
or UO_792 (O_792,N_5555,N_5041);
nor UO_793 (O_793,N_5993,N_9176);
xor UO_794 (O_794,N_5468,N_7960);
and UO_795 (O_795,N_9723,N_9581);
and UO_796 (O_796,N_9087,N_9195);
nand UO_797 (O_797,N_7588,N_9267);
or UO_798 (O_798,N_5686,N_6831);
nor UO_799 (O_799,N_9393,N_7227);
nor UO_800 (O_800,N_5772,N_5491);
and UO_801 (O_801,N_5849,N_9677);
or UO_802 (O_802,N_8432,N_9200);
or UO_803 (O_803,N_9513,N_7538);
and UO_804 (O_804,N_6780,N_9801);
nand UO_805 (O_805,N_8511,N_7782);
nand UO_806 (O_806,N_7403,N_8692);
nor UO_807 (O_807,N_5467,N_7541);
nand UO_808 (O_808,N_9522,N_8512);
nand UO_809 (O_809,N_6625,N_7188);
or UO_810 (O_810,N_6320,N_8828);
and UO_811 (O_811,N_6354,N_9730);
and UO_812 (O_812,N_8698,N_8402);
and UO_813 (O_813,N_7128,N_5317);
nor UO_814 (O_814,N_9004,N_7099);
or UO_815 (O_815,N_5637,N_9144);
and UO_816 (O_816,N_9426,N_5741);
nor UO_817 (O_817,N_7628,N_7473);
nand UO_818 (O_818,N_7075,N_6061);
xnor UO_819 (O_819,N_5400,N_9876);
or UO_820 (O_820,N_9805,N_7416);
and UO_821 (O_821,N_9991,N_7056);
nand UO_822 (O_822,N_6879,N_7682);
nand UO_823 (O_823,N_6041,N_6029);
or UO_824 (O_824,N_7229,N_6333);
nor UO_825 (O_825,N_8500,N_5620);
nand UO_826 (O_826,N_5498,N_7312);
nor UO_827 (O_827,N_6485,N_8396);
nor UO_828 (O_828,N_9355,N_9222);
or UO_829 (O_829,N_5789,N_8903);
nor UO_830 (O_830,N_7689,N_7216);
xor UO_831 (O_831,N_6511,N_9334);
or UO_832 (O_832,N_7319,N_9362);
and UO_833 (O_833,N_9822,N_7964);
nor UO_834 (O_834,N_8304,N_5606);
and UO_835 (O_835,N_8171,N_5768);
or UO_836 (O_836,N_6692,N_5103);
and UO_837 (O_837,N_8537,N_6267);
nand UO_838 (O_838,N_5402,N_8233);
or UO_839 (O_839,N_9558,N_7788);
nor UO_840 (O_840,N_5436,N_8923);
nand UO_841 (O_841,N_9518,N_7277);
and UO_842 (O_842,N_7302,N_9098);
nand UO_843 (O_843,N_8074,N_5687);
nand UO_844 (O_844,N_7576,N_5928);
or UO_845 (O_845,N_8648,N_8061);
nand UO_846 (O_846,N_6444,N_8535);
nand UO_847 (O_847,N_7019,N_9221);
and UO_848 (O_848,N_5661,N_6753);
nor UO_849 (O_849,N_5130,N_9682);
and UO_850 (O_850,N_7458,N_9234);
and UO_851 (O_851,N_7298,N_5706);
nor UO_852 (O_852,N_9609,N_5419);
or UO_853 (O_853,N_5834,N_9781);
or UO_854 (O_854,N_8254,N_6325);
or UO_855 (O_855,N_5442,N_9113);
and UO_856 (O_856,N_9035,N_6086);
nor UO_857 (O_857,N_5406,N_7261);
nor UO_858 (O_858,N_7139,N_6962);
nor UO_859 (O_859,N_5019,N_6020);
nand UO_860 (O_860,N_7156,N_9646);
nor UO_861 (O_861,N_8100,N_8498);
and UO_862 (O_862,N_7297,N_7565);
or UO_863 (O_863,N_6429,N_9344);
nand UO_864 (O_864,N_8226,N_9278);
or UO_865 (O_865,N_8994,N_5004);
nor UO_866 (O_866,N_9908,N_6174);
nor UO_867 (O_867,N_7560,N_7792);
and UO_868 (O_868,N_7049,N_5384);
and UO_869 (O_869,N_5853,N_7438);
or UO_870 (O_870,N_5574,N_5551);
or UO_871 (O_871,N_7189,N_6487);
and UO_872 (O_872,N_9985,N_6145);
and UO_873 (O_873,N_8142,N_9865);
nor UO_874 (O_874,N_5585,N_6481);
and UO_875 (O_875,N_8968,N_9614);
and UO_876 (O_876,N_8757,N_9611);
and UO_877 (O_877,N_8184,N_7186);
and UO_878 (O_878,N_7652,N_6306);
nor UO_879 (O_879,N_8725,N_8096);
nand UO_880 (O_880,N_9153,N_5487);
and UO_881 (O_881,N_7366,N_8627);
or UO_882 (O_882,N_8598,N_6100);
nand UO_883 (O_883,N_7404,N_5953);
nor UO_884 (O_884,N_8188,N_6974);
or UO_885 (O_885,N_5023,N_8649);
and UO_886 (O_886,N_5021,N_5729);
and UO_887 (O_887,N_6721,N_7904);
and UO_888 (O_888,N_9594,N_9984);
nor UO_889 (O_889,N_6397,N_9727);
nor UO_890 (O_890,N_7535,N_5616);
xor UO_891 (O_891,N_9762,N_9226);
nand UO_892 (O_892,N_6941,N_9530);
and UO_893 (O_893,N_9662,N_8531);
and UO_894 (O_894,N_6921,N_7586);
or UO_895 (O_895,N_7065,N_9797);
and UO_896 (O_896,N_8892,N_9239);
and UO_897 (O_897,N_7353,N_7991);
nor UO_898 (O_898,N_8463,N_6253);
and UO_899 (O_899,N_5923,N_8644);
and UO_900 (O_900,N_7802,N_9684);
nand UO_901 (O_901,N_5446,N_5981);
and UO_902 (O_902,N_7421,N_9834);
and UO_903 (O_903,N_6646,N_8720);
or UO_904 (O_904,N_7516,N_7930);
nand UO_905 (O_905,N_8207,N_5519);
nand UO_906 (O_906,N_6317,N_6722);
or UO_907 (O_907,N_8622,N_9506);
nand UO_908 (O_908,N_5379,N_6567);
nand UO_909 (O_909,N_7723,N_6184);
or UO_910 (O_910,N_7425,N_9653);
and UO_911 (O_911,N_9729,N_7476);
or UO_912 (O_912,N_6286,N_9794);
nand UO_913 (O_913,N_7164,N_9814);
nand UO_914 (O_914,N_6297,N_7487);
and UO_915 (O_915,N_6581,N_8123);
or UO_916 (O_916,N_6224,N_7974);
nor UO_917 (O_917,N_9138,N_8424);
or UO_918 (O_918,N_5847,N_7484);
or UO_919 (O_919,N_8767,N_6357);
nand UO_920 (O_920,N_5175,N_6910);
nand UO_921 (O_921,N_6012,N_7518);
nand UO_922 (O_922,N_6358,N_6338);
and UO_923 (O_923,N_6367,N_9542);
nor UO_924 (O_924,N_5995,N_8541);
and UO_925 (O_925,N_7357,N_6644);
and UO_926 (O_926,N_5285,N_5512);
nor UO_927 (O_927,N_6551,N_5364);
nor UO_928 (O_928,N_7816,N_6731);
or UO_929 (O_929,N_8115,N_8925);
and UO_930 (O_930,N_5515,N_5930);
and UO_931 (O_931,N_9088,N_5893);
or UO_932 (O_932,N_5322,N_8085);
nor UO_933 (O_933,N_7720,N_8673);
nor UO_934 (O_934,N_8238,N_9681);
or UO_935 (O_935,N_9808,N_5026);
nor UO_936 (O_936,N_6023,N_8325);
nor UO_937 (O_937,N_6857,N_7213);
or UO_938 (O_938,N_7376,N_6407);
and UO_939 (O_939,N_8094,N_7182);
nor UO_940 (O_940,N_8745,N_7971);
and UO_941 (O_941,N_5110,N_8165);
or UO_942 (O_942,N_5694,N_7330);
nor UO_943 (O_943,N_8754,N_9145);
nand UO_944 (O_944,N_9403,N_7685);
nand UO_945 (O_945,N_8363,N_8616);
and UO_946 (O_946,N_5896,N_7875);
and UO_947 (O_947,N_6903,N_9500);
nor UO_948 (O_948,N_8442,N_6756);
nand UO_949 (O_949,N_5085,N_9120);
nand UO_950 (O_950,N_7086,N_9735);
or UO_951 (O_951,N_7125,N_5313);
and UO_952 (O_952,N_6998,N_7433);
nand UO_953 (O_953,N_8908,N_7053);
or UO_954 (O_954,N_6214,N_6363);
and UO_955 (O_955,N_9440,N_9036);
or UO_956 (O_956,N_5989,N_8045);
nor UO_957 (O_957,N_8516,N_6700);
nor UO_958 (O_958,N_7051,N_8955);
or UO_959 (O_959,N_8675,N_5752);
xnor UO_960 (O_960,N_5703,N_5922);
and UO_961 (O_961,N_7238,N_8723);
nor UO_962 (O_962,N_6944,N_6709);
or UO_963 (O_963,N_8017,N_8489);
nand UO_964 (O_964,N_7381,N_8470);
or UO_965 (O_965,N_8032,N_9127);
nor UO_966 (O_966,N_6436,N_5277);
nor UO_967 (O_967,N_5107,N_7759);
nor UO_968 (O_968,N_7967,N_8905);
xor UO_969 (O_969,N_9039,N_6845);
nand UO_970 (O_970,N_7159,N_8436);
nand UO_971 (O_971,N_8447,N_8283);
nor UO_972 (O_972,N_9969,N_5662);
and UO_973 (O_973,N_6396,N_6704);
nor UO_974 (O_974,N_9032,N_7148);
nand UO_975 (O_975,N_9050,N_6985);
nand UO_976 (O_976,N_5767,N_6637);
nand UO_977 (O_977,N_8962,N_7415);
nor UO_978 (O_978,N_7386,N_7215);
nor UO_979 (O_979,N_9360,N_5255);
and UO_980 (O_980,N_9912,N_6640);
nor UO_981 (O_981,N_6456,N_7060);
or UO_982 (O_982,N_6143,N_6056);
or UO_983 (O_983,N_8205,N_7272);
nand UO_984 (O_984,N_7300,N_9248);
or UO_985 (O_985,N_9627,N_5877);
nand UO_986 (O_986,N_9712,N_5089);
and UO_987 (O_987,N_9725,N_8213);
nor UO_988 (O_988,N_5570,N_8582);
nand UO_989 (O_989,N_9233,N_8025);
nor UO_990 (O_990,N_6724,N_8932);
and UO_991 (O_991,N_6099,N_9203);
or UO_992 (O_992,N_6940,N_9565);
and UO_993 (O_993,N_8824,N_8937);
nand UO_994 (O_994,N_5242,N_8490);
nor UO_995 (O_995,N_5274,N_8120);
or UO_996 (O_996,N_9373,N_7242);
and UO_997 (O_997,N_8995,N_6904);
nand UO_998 (O_998,N_7434,N_9460);
or UO_999 (O_999,N_6869,N_8681);
nand UO_1000 (O_1000,N_9698,N_5517);
and UO_1001 (O_1001,N_9497,N_5022);
and UO_1002 (O_1002,N_6562,N_5985);
nor UO_1003 (O_1003,N_9870,N_8503);
nor UO_1004 (O_1004,N_8517,N_8425);
and UO_1005 (O_1005,N_6409,N_5862);
or UO_1006 (O_1006,N_9163,N_5888);
or UO_1007 (O_1007,N_5604,N_6660);
nand UO_1008 (O_1008,N_9911,N_5059);
nand UO_1009 (O_1009,N_7071,N_5696);
nor UO_1010 (O_1010,N_7637,N_5283);
or UO_1011 (O_1011,N_8303,N_5422);
and UO_1012 (O_1012,N_6502,N_5176);
or UO_1013 (O_1013,N_9936,N_9230);
or UO_1014 (O_1014,N_8890,N_7916);
nand UO_1015 (O_1015,N_6419,N_9577);
nor UO_1016 (O_1016,N_7734,N_6296);
nand UO_1017 (O_1017,N_8350,N_8732);
nor UO_1018 (O_1018,N_7057,N_9354);
nor UO_1019 (O_1019,N_6114,N_9258);
and UO_1020 (O_1020,N_7010,N_7147);
and UO_1021 (O_1021,N_8914,N_8719);
nand UO_1022 (O_1022,N_5980,N_9131);
or UO_1023 (O_1023,N_5564,N_7649);
and UO_1024 (O_1024,N_9697,N_7293);
nor UO_1025 (O_1025,N_5388,N_9774);
nor UO_1026 (O_1026,N_5359,N_7849);
nor UO_1027 (O_1027,N_8204,N_6633);
nand UO_1028 (O_1028,N_7972,N_6496);
and UO_1029 (O_1029,N_9010,N_9739);
nand UO_1030 (O_1030,N_7590,N_9676);
and UO_1031 (O_1031,N_5352,N_6484);
xnor UO_1032 (O_1032,N_6383,N_5559);
nand UO_1033 (O_1033,N_8920,N_6559);
nor UO_1034 (O_1034,N_6792,N_6657);
nor UO_1035 (O_1035,N_6537,N_5440);
and UO_1036 (O_1036,N_6425,N_8866);
nand UO_1037 (O_1037,N_6263,N_5691);
or UO_1038 (O_1038,N_8965,N_8099);
or UO_1039 (O_1039,N_5001,N_8318);
and UO_1040 (O_1040,N_9773,N_6223);
nand UO_1041 (O_1041,N_5342,N_8126);
nor UO_1042 (O_1042,N_7253,N_5320);
and UO_1043 (O_1043,N_6729,N_8570);
nand UO_1044 (O_1044,N_9424,N_9044);
and UO_1045 (O_1045,N_6856,N_6183);
and UO_1046 (O_1046,N_6606,N_9587);
and UO_1047 (O_1047,N_9211,N_6694);
nor UO_1048 (O_1048,N_5061,N_9918);
nand UO_1049 (O_1049,N_9844,N_8095);
and UO_1050 (O_1050,N_6760,N_6603);
xnor UO_1051 (O_1051,N_7529,N_5709);
and UO_1052 (O_1052,N_7033,N_8911);
nand UO_1053 (O_1053,N_9633,N_6058);
nor UO_1054 (O_1054,N_7050,N_8331);
nand UO_1055 (O_1055,N_7660,N_5452);
nand UO_1056 (O_1056,N_9966,N_6081);
or UO_1057 (O_1057,N_8766,N_8336);
nor UO_1058 (O_1058,N_9139,N_6912);
or UO_1059 (O_1059,N_9757,N_6372);
or UO_1060 (O_1060,N_7678,N_7102);
nand UO_1061 (O_1061,N_8294,N_6762);
nor UO_1062 (O_1062,N_9021,N_8715);
or UO_1063 (O_1063,N_9531,N_7852);
nor UO_1064 (O_1064,N_6337,N_8889);
nor UO_1065 (O_1065,N_7919,N_5053);
nor UO_1066 (O_1066,N_8001,N_6503);
nor UO_1067 (O_1067,N_5675,N_9721);
nor UO_1068 (O_1068,N_7598,N_9076);
or UO_1069 (O_1069,N_7569,N_5183);
or UO_1070 (O_1070,N_6209,N_7324);
nor UO_1071 (O_1071,N_8700,N_5539);
or UO_1072 (O_1072,N_7895,N_5080);
nor UO_1073 (O_1073,N_6382,N_9231);
or UO_1074 (O_1074,N_8197,N_7373);
nand UO_1075 (O_1075,N_6999,N_5281);
nand UO_1076 (O_1076,N_5826,N_6159);
and UO_1077 (O_1077,N_8008,N_6084);
nand UO_1078 (O_1078,N_9480,N_9058);
nor UO_1079 (O_1079,N_5269,N_8386);
and UO_1080 (O_1080,N_8097,N_6515);
or UO_1081 (O_1081,N_9412,N_7384);
or UO_1082 (O_1082,N_7396,N_9086);
or UO_1083 (O_1083,N_7968,N_7014);
nor UO_1084 (O_1084,N_5769,N_8969);
nand UO_1085 (O_1085,N_7988,N_8562);
xor UO_1086 (O_1086,N_9795,N_9955);
or UO_1087 (O_1087,N_7700,N_7710);
and UO_1088 (O_1088,N_6829,N_9256);
nor UO_1089 (O_1089,N_9826,N_9279);
nor UO_1090 (O_1090,N_8846,N_9618);
and UO_1091 (O_1091,N_6220,N_6835);
and UO_1092 (O_1092,N_8469,N_8114);
nor UO_1093 (O_1093,N_5755,N_7508);
nor UO_1094 (O_1094,N_7085,N_5449);
and UO_1095 (O_1095,N_6596,N_7025);
nand UO_1096 (O_1096,N_7571,N_5365);
and UO_1097 (O_1097,N_8046,N_8722);
or UO_1098 (O_1098,N_7674,N_7463);
or UO_1099 (O_1099,N_6675,N_5965);
nor UO_1100 (O_1100,N_7194,N_7667);
and UO_1101 (O_1101,N_8324,N_6521);
nand UO_1102 (O_1102,N_5835,N_7536);
and UO_1103 (O_1103,N_7219,N_7544);
nor UO_1104 (O_1104,N_7000,N_5804);
and UO_1105 (O_1105,N_6549,N_6508);
or UO_1106 (O_1106,N_8913,N_5846);
nor UO_1107 (O_1107,N_6266,N_5420);
or UO_1108 (O_1108,N_7280,N_5851);
nand UO_1109 (O_1109,N_9041,N_9489);
nand UO_1110 (O_1110,N_9706,N_9779);
nor UO_1111 (O_1111,N_5220,N_9494);
nor UO_1112 (O_1112,N_6268,N_6529);
nand UO_1113 (O_1113,N_9978,N_8777);
and UO_1114 (O_1114,N_5497,N_8785);
or UO_1115 (O_1115,N_5652,N_5360);
or UO_1116 (O_1116,N_5750,N_5146);
nand UO_1117 (O_1117,N_5014,N_5816);
nor UO_1118 (O_1118,N_9995,N_9578);
nand UO_1119 (O_1119,N_5147,N_6158);
and UO_1120 (O_1120,N_7497,N_9219);
nand UO_1121 (O_1121,N_8180,N_7336);
or UO_1122 (O_1122,N_6331,N_8860);
or UO_1123 (O_1123,N_6366,N_8867);
nor UO_1124 (O_1124,N_7311,N_9094);
and UO_1125 (O_1125,N_8055,N_6175);
nand UO_1126 (O_1126,N_8297,N_9673);
nor UO_1127 (O_1127,N_9040,N_5037);
nand UO_1128 (O_1128,N_9786,N_9443);
and UO_1129 (O_1129,N_6908,N_8406);
nand UO_1130 (O_1130,N_7094,N_8449);
and UO_1131 (O_1131,N_5235,N_8740);
nor UO_1132 (O_1132,N_9475,N_7483);
and UO_1133 (O_1133,N_7361,N_5371);
or UO_1134 (O_1134,N_6501,N_5408);
or UO_1135 (O_1135,N_5734,N_7333);
and UO_1136 (O_1136,N_5627,N_5114);
nor UO_1137 (O_1137,N_5771,N_7639);
nor UO_1138 (O_1138,N_7409,N_7506);
and UO_1139 (O_1139,N_5891,N_9927);
nor UO_1140 (O_1140,N_7149,N_8015);
nand UO_1141 (O_1141,N_8999,N_5654);
and UO_1142 (O_1142,N_6965,N_9106);
or UO_1143 (O_1143,N_5563,N_8744);
or UO_1144 (O_1144,N_5996,N_8156);
nand UO_1145 (O_1145,N_7829,N_7855);
or UO_1146 (O_1146,N_7784,N_8416);
nand UO_1147 (O_1147,N_5417,N_7982);
and UO_1148 (O_1148,N_6672,N_7796);
nand UO_1149 (O_1149,N_5346,N_6600);
and UO_1150 (O_1150,N_6250,N_7871);
or UO_1151 (O_1151,N_9859,N_8915);
nor UO_1152 (O_1152,N_5465,N_5451);
and UO_1153 (O_1153,N_6847,N_6276);
nand UO_1154 (O_1154,N_7114,N_8686);
nand UO_1155 (O_1155,N_7531,N_8546);
or UO_1156 (O_1156,N_9312,N_5494);
xnor UO_1157 (O_1157,N_9543,N_9421);
or UO_1158 (O_1158,N_7160,N_5906);
and UO_1159 (O_1159,N_8630,N_8323);
and UO_1160 (O_1160,N_9151,N_7423);
or UO_1161 (O_1161,N_5603,N_8116);
or UO_1162 (O_1162,N_6883,N_5589);
and UO_1163 (O_1163,N_7915,N_9327);
or UO_1164 (O_1164,N_7737,N_5409);
nand UO_1165 (O_1165,N_7515,N_7437);
nor UO_1166 (O_1166,N_8472,N_7592);
nor UO_1167 (O_1167,N_9181,N_7825);
or UO_1168 (O_1168,N_7355,N_6404);
nor UO_1169 (O_1169,N_7620,N_9968);
nor UO_1170 (O_1170,N_7460,N_5925);
and UO_1171 (O_1171,N_7232,N_7980);
nor UO_1172 (O_1172,N_8829,N_8680);
nand UO_1173 (O_1173,N_5647,N_6505);
nand UO_1174 (O_1174,N_6117,N_8471);
or UO_1175 (O_1175,N_8431,N_5079);
nand UO_1176 (O_1176,N_5593,N_7767);
nand UO_1177 (O_1177,N_9254,N_9648);
or UO_1178 (O_1178,N_6624,N_7126);
or UO_1179 (O_1179,N_9310,N_6772);
nand UO_1180 (O_1180,N_6232,N_5735);
nor UO_1181 (O_1181,N_5990,N_9647);
or UO_1182 (O_1182,N_6900,N_9376);
and UO_1183 (O_1183,N_7138,N_7866);
nand UO_1184 (O_1184,N_6571,N_8081);
or UO_1185 (O_1185,N_8689,N_7897);
and UO_1186 (O_1186,N_9427,N_5998);
nor UO_1187 (O_1187,N_9060,N_5739);
nor UO_1188 (O_1188,N_6891,N_8284);
or UO_1189 (O_1189,N_7176,N_6686);
and UO_1190 (O_1190,N_9780,N_6021);
nand UO_1191 (O_1191,N_6854,N_7736);
nor UO_1192 (O_1192,N_8734,N_5131);
or UO_1193 (O_1193,N_8990,N_6959);
nand UO_1194 (O_1194,N_5380,N_6393);
and UO_1195 (O_1195,N_7274,N_8327);
and UO_1196 (O_1196,N_8141,N_6950);
nor UO_1197 (O_1197,N_9571,N_5749);
and UO_1198 (O_1198,N_5573,N_9498);
nand UO_1199 (O_1199,N_5076,N_7854);
and UO_1200 (O_1200,N_7712,N_7117);
nor UO_1201 (O_1201,N_7589,N_9319);
nand UO_1202 (O_1202,N_8093,N_7910);
nand UO_1203 (O_1203,N_9054,N_9110);
or UO_1204 (O_1204,N_7349,N_6460);
nor UO_1205 (O_1205,N_7021,N_9756);
nor UO_1206 (O_1206,N_8505,N_9523);
nand UO_1207 (O_1207,N_9399,N_9576);
nand UO_1208 (O_1208,N_9862,N_7898);
nor UO_1209 (O_1209,N_5447,N_8655);
or UO_1210 (O_1210,N_6318,N_9463);
xor UO_1211 (O_1211,N_5916,N_6728);
nor UO_1212 (O_1212,N_7512,N_6455);
nor UO_1213 (O_1213,N_7762,N_8807);
or UO_1214 (O_1214,N_8476,N_9451);
and UO_1215 (O_1215,N_8092,N_7724);
nor UO_1216 (O_1216,N_8868,N_8376);
nand UO_1217 (O_1217,N_8989,N_8048);
or UO_1218 (O_1218,N_7395,N_8899);
and UO_1219 (O_1219,N_6315,N_8724);
nor UO_1220 (O_1220,N_8078,N_8289);
nand UO_1221 (O_1221,N_5395,N_8606);
nor UO_1222 (O_1222,N_7343,N_6448);
and UO_1223 (O_1223,N_7061,N_5895);
and UO_1224 (O_1224,N_8349,N_7332);
nand UO_1225 (O_1225,N_9128,N_9977);
and UO_1226 (O_1226,N_8027,N_9631);
or UO_1227 (O_1227,N_7151,N_6442);
xnor UO_1228 (O_1228,N_8358,N_6330);
and UO_1229 (O_1229,N_9441,N_7716);
nor UO_1230 (O_1230,N_9547,N_7543);
and UO_1231 (O_1231,N_5429,N_7722);
nor UO_1232 (O_1232,N_6242,N_8521);
nor UO_1233 (O_1233,N_9796,N_5999);
and UO_1234 (O_1234,N_5967,N_6514);
or UO_1235 (O_1235,N_6558,N_6305);
nor UO_1236 (O_1236,N_6176,N_7769);
nand UO_1237 (O_1237,N_8419,N_9493);
nor UO_1238 (O_1238,N_9006,N_6535);
or UO_1239 (O_1239,N_6019,N_9299);
nor UO_1240 (O_1240,N_7978,N_6395);
nand UO_1241 (O_1241,N_8663,N_5848);
or UO_1242 (O_1242,N_7656,N_8172);
nor UO_1243 (O_1243,N_9784,N_7527);
and UO_1244 (O_1244,N_5974,N_7521);
nand UO_1245 (O_1245,N_8024,N_5975);
and UO_1246 (O_1246,N_6111,N_8189);
and UO_1247 (O_1247,N_9528,N_6570);
nand UO_1248 (O_1248,N_6568,N_9273);
nand UO_1249 (O_1249,N_9907,N_7887);
or UO_1250 (O_1250,N_8543,N_6967);
nor UO_1251 (O_1251,N_7902,N_7907);
and UO_1252 (O_1252,N_5454,N_9177);
and UO_1253 (O_1253,N_7307,N_5597);
nand UO_1254 (O_1254,N_6412,N_9580);
or UO_1255 (O_1255,N_9938,N_8007);
and UO_1256 (O_1256,N_6946,N_7356);
nor UO_1257 (O_1257,N_9137,N_7320);
and UO_1258 (O_1258,N_8166,N_7699);
nor UO_1259 (O_1259,N_6956,N_7116);
and UO_1260 (O_1260,N_9300,N_8229);
or UO_1261 (O_1261,N_8919,N_8388);
or UO_1262 (O_1262,N_8271,N_7684);
nor UO_1263 (O_1263,N_5840,N_8554);
or UO_1264 (O_1264,N_8670,N_8082);
or UO_1265 (O_1265,N_8636,N_9861);
and UO_1266 (O_1266,N_7746,N_6085);
and UO_1267 (O_1267,N_5230,N_9637);
xor UO_1268 (O_1268,N_9229,N_5316);
or UO_1269 (O_1269,N_5155,N_7711);
or UO_1270 (O_1270,N_8104,N_8539);
nand UO_1271 (O_1271,N_5239,N_6410);
nand UO_1272 (O_1272,N_8885,N_8930);
and UO_1273 (O_1273,N_5441,N_6575);
or UO_1274 (O_1274,N_7860,N_8839);
nor UO_1275 (O_1275,N_7997,N_6500);
nor UO_1276 (O_1276,N_8850,N_9595);
nand UO_1277 (O_1277,N_6030,N_7947);
or UO_1278 (O_1278,N_6717,N_5015);
and UO_1279 (O_1279,N_6230,N_8564);
and UO_1280 (O_1280,N_5397,N_8394);
or UO_1281 (O_1281,N_8640,N_7913);
xor UO_1282 (O_1282,N_8158,N_5222);
and UO_1283 (O_1283,N_8345,N_7554);
or UO_1284 (O_1284,N_8339,N_7806);
or UO_1285 (O_1285,N_7579,N_7202);
nand UO_1286 (O_1286,N_8236,N_7790);
or UO_1287 (O_1287,N_6123,N_7841);
nor UO_1288 (O_1288,N_8676,N_6045);
or UO_1289 (O_1289,N_5157,N_6428);
and UO_1290 (O_1290,N_8895,N_7732);
nand UO_1291 (O_1291,N_7185,N_9733);
nand UO_1292 (O_1292,N_8030,N_8161);
nor UO_1293 (O_1293,N_5267,N_5219);
nor UO_1294 (O_1294,N_7234,N_8551);
and UO_1295 (O_1295,N_8223,N_7226);
nor UO_1296 (O_1296,N_6822,N_6046);
nor UO_1297 (O_1297,N_5919,N_7144);
nand UO_1298 (O_1298,N_7008,N_6039);
or UO_1299 (O_1299,N_7618,N_5762);
and UO_1300 (O_1300,N_6127,N_5232);
or UO_1301 (O_1301,N_8771,N_5730);
and UO_1302 (O_1302,N_6335,N_6513);
nor UO_1303 (O_1303,N_8924,N_8245);
and UO_1304 (O_1304,N_5933,N_5203);
nand UO_1305 (O_1305,N_6400,N_5499);
or UO_1306 (O_1306,N_8322,N_5737);
or UO_1307 (O_1307,N_5902,N_8004);
nand UO_1308 (O_1308,N_8428,N_7641);
nor UO_1309 (O_1309,N_5530,N_9604);
nand UO_1310 (O_1310,N_9283,N_8620);
nand UO_1311 (O_1311,N_6654,N_9429);
xnor UO_1312 (O_1312,N_6520,N_6295);
or UO_1313 (O_1313,N_8340,N_8177);
and UO_1314 (O_1314,N_6663,N_9242);
and UO_1315 (O_1315,N_8800,N_9920);
nand UO_1316 (O_1316,N_6492,N_8481);
or UO_1317 (O_1317,N_5566,N_5987);
and UO_1318 (O_1318,N_8897,N_5544);
or UO_1319 (O_1319,N_8632,N_5309);
and UO_1320 (O_1320,N_9583,N_5161);
and UO_1321 (O_1321,N_8976,N_6423);
and UO_1322 (O_1322,N_5509,N_7392);
nor UO_1323 (O_1323,N_9123,N_6922);
nor UO_1324 (O_1324,N_5201,N_7203);
nor UO_1325 (O_1325,N_5821,N_5016);
nor UO_1326 (O_1326,N_6645,N_5314);
and UO_1327 (O_1327,N_9048,N_9988);
or UO_1328 (O_1328,N_5414,N_5765);
nand UO_1329 (O_1329,N_8825,N_5764);
nand UO_1330 (O_1330,N_8404,N_5361);
and UO_1331 (O_1331,N_5859,N_6289);
nor UO_1332 (O_1332,N_9407,N_6802);
or UO_1333 (O_1333,N_9574,N_9839);
and UO_1334 (O_1334,N_8533,N_8014);
nand UO_1335 (O_1335,N_8992,N_6454);
nand UO_1336 (O_1336,N_6119,N_7594);
nand UO_1337 (O_1337,N_9919,N_5889);
nand UO_1338 (O_1338,N_7453,N_8400);
or UO_1339 (O_1339,N_9749,N_9613);
nor UO_1340 (O_1340,N_7730,N_7136);
nor UO_1341 (O_1341,N_5169,N_8013);
nand UO_1342 (O_1342,N_5141,N_9164);
or UO_1343 (O_1343,N_8330,N_5375);
and UO_1344 (O_1344,N_5582,N_9987);
nor UO_1345 (O_1345,N_8792,N_9001);
nor UO_1346 (O_1346,N_7764,N_5944);
and UO_1347 (O_1347,N_5357,N_5349);
and UO_1348 (O_1348,N_7052,N_5474);
nor UO_1349 (O_1349,N_9804,N_9339);
or UO_1350 (O_1350,N_9903,N_8348);
and UO_1351 (O_1351,N_8248,N_5802);
and UO_1352 (O_1352,N_7200,N_6234);
or UO_1353 (O_1353,N_5476,N_6463);
nand UO_1354 (O_1354,N_5172,N_6788);
and UO_1355 (O_1355,N_5612,N_7177);
or UO_1356 (O_1356,N_6302,N_7704);
nor UO_1357 (O_1357,N_8086,N_5591);
nand UO_1358 (O_1358,N_8136,N_5792);
nand UO_1359 (O_1359,N_8065,N_8977);
nand UO_1360 (O_1360,N_9999,N_9324);
nor UO_1361 (O_1361,N_5189,N_9564);
nor UO_1362 (O_1362,N_7165,N_9308);
nand UO_1363 (O_1363,N_5084,N_8706);
nor UO_1364 (O_1364,N_6205,N_8738);
or UO_1365 (O_1365,N_7166,N_7462);
nor UO_1366 (O_1366,N_7499,N_7444);
nor UO_1367 (O_1367,N_6947,N_6953);
nor UO_1368 (O_1368,N_8647,N_9974);
nand UO_1369 (O_1369,N_5456,N_9169);
and UO_1370 (O_1370,N_9346,N_5667);
and UO_1371 (O_1371,N_9026,N_6671);
or UO_1372 (O_1372,N_8191,N_5886);
nand UO_1373 (O_1373,N_9625,N_7001);
or UO_1374 (O_1374,N_8851,N_9567);
and UO_1375 (O_1375,N_8980,N_8145);
or UO_1376 (O_1376,N_6173,N_5801);
xnor UO_1377 (O_1377,N_5692,N_6897);
nand UO_1378 (O_1378,N_7173,N_9819);
and UO_1379 (O_1379,N_8277,N_8996);
nor UO_1380 (O_1380,N_8076,N_5010);
or UO_1381 (O_1381,N_6775,N_8975);
and UO_1382 (O_1382,N_6151,N_7447);
or UO_1383 (O_1383,N_5376,N_9929);
nand UO_1384 (O_1384,N_8023,N_6695);
nand UO_1385 (O_1385,N_6825,N_5813);
nor UO_1386 (O_1386,N_6986,N_9447);
nand UO_1387 (O_1387,N_5108,N_9828);
or UO_1388 (O_1388,N_8665,N_7900);
and UO_1389 (O_1389,N_7183,N_9954);
nor UO_1390 (O_1390,N_9442,N_5433);
or UO_1391 (O_1391,N_8733,N_6300);
and UO_1392 (O_1392,N_9585,N_6431);
nor UO_1393 (O_1393,N_7891,N_5639);
nand UO_1394 (O_1394,N_8684,N_7758);
nand UO_1395 (O_1395,N_8967,N_5385);
nor UO_1396 (O_1396,N_9132,N_8902);
nand UO_1397 (O_1397,N_7199,N_8814);
xor UO_1398 (O_1398,N_6450,N_5332);
nor UO_1399 (O_1399,N_7937,N_6542);
nor UO_1400 (O_1400,N_7839,N_8653);
or UO_1401 (O_1401,N_5778,N_6817);
nor UO_1402 (O_1402,N_8000,N_8569);
and UO_1403 (O_1403,N_6613,N_7805);
nand UO_1404 (O_1404,N_8832,N_6530);
and UO_1405 (O_1405,N_8182,N_5677);
and UO_1406 (O_1406,N_6375,N_8841);
or UO_1407 (O_1407,N_9858,N_7747);
or UO_1408 (O_1408,N_6468,N_5099);
nor UO_1409 (O_1409,N_6877,N_6665);
and UO_1410 (O_1410,N_5506,N_7398);
nor UO_1411 (O_1411,N_5133,N_7648);
or UO_1412 (O_1412,N_5869,N_8029);
nand UO_1413 (O_1413,N_7524,N_8252);
or UO_1414 (O_1414,N_7368,N_7605);
and UO_1415 (O_1415,N_6471,N_7756);
nand UO_1416 (O_1416,N_8378,N_9832);
nand UO_1417 (O_1417,N_6507,N_9851);
nor UO_1418 (O_1418,N_6206,N_9348);
nor UO_1419 (O_1419,N_9850,N_8395);
and UO_1420 (O_1420,N_9713,N_5060);
or UO_1421 (O_1421,N_7781,N_8797);
or UO_1422 (O_1422,N_7946,N_5028);
nand UO_1423 (O_1423,N_9771,N_8043);
or UO_1424 (O_1424,N_8261,N_8592);
or UO_1425 (O_1425,N_9315,N_9135);
nand UO_1426 (O_1426,N_9387,N_5481);
or UO_1427 (O_1427,N_6065,N_7795);
nor UO_1428 (O_1428,N_6040,N_7864);
nand UO_1429 (O_1429,N_8884,N_6957);
and UO_1430 (O_1430,N_7493,N_7397);
or UO_1431 (O_1431,N_9314,N_7814);
nor UO_1432 (O_1432,N_6678,N_9422);
nor UO_1433 (O_1433,N_5722,N_6265);
or UO_1434 (O_1434,N_8799,N_9649);
nor UO_1435 (O_1435,N_5218,N_9165);
and UO_1436 (O_1436,N_8393,N_5532);
nand UO_1437 (O_1437,N_7448,N_5480);
nand UO_1438 (O_1438,N_9479,N_9379);
nand UO_1439 (O_1439,N_7838,N_5658);
nand UO_1440 (O_1440,N_8796,N_6095);
and UO_1441 (O_1441,N_9679,N_6311);
nand UO_1442 (O_1442,N_7600,N_7022);
and UO_1443 (O_1443,N_5701,N_5705);
and UO_1444 (O_1444,N_5992,N_8147);
nor UO_1445 (O_1445,N_9579,N_7106);
nand UO_1446 (O_1446,N_6126,N_6416);
nor UO_1447 (O_1447,N_7969,N_5858);
or UO_1448 (O_1448,N_7580,N_7545);
nor UO_1449 (O_1449,N_7115,N_6614);
nor UO_1450 (O_1450,N_9505,N_8639);
and UO_1451 (O_1451,N_7998,N_9515);
and UO_1452 (O_1452,N_5430,N_9935);
nand UO_1453 (O_1453,N_9409,N_7122);
or UO_1454 (O_1454,N_8050,N_8075);
and UO_1455 (O_1455,N_8295,N_8031);
nand UO_1456 (O_1456,N_8847,N_6475);
nand UO_1457 (O_1457,N_6062,N_7252);
nand UO_1458 (O_1458,N_7231,N_9389);
or UO_1459 (O_1459,N_8863,N_9115);
and UO_1460 (O_1460,N_8997,N_6785);
xnor UO_1461 (O_1461,N_7763,N_7265);
and UO_1462 (O_1462,N_7411,N_6776);
and UO_1463 (O_1463,N_7452,N_6783);
or UO_1464 (O_1464,N_8815,N_5715);
nor UO_1465 (O_1465,N_8590,N_8244);
nor UO_1466 (O_1466,N_5969,N_5165);
and UO_1467 (O_1467,N_6466,N_7894);
nand UO_1468 (O_1468,N_6430,N_6352);
nand UO_1469 (O_1469,N_5850,N_7886);
nand UO_1470 (O_1470,N_8341,N_8337);
and UO_1471 (O_1471,N_9863,N_5592);
nand UO_1472 (O_1472,N_9051,N_9092);
and UO_1473 (O_1473,N_8477,N_6813);
and UO_1474 (O_1474,N_8602,N_8118);
and UO_1475 (O_1475,N_6088,N_9274);
nor UO_1476 (O_1476,N_7028,N_7041);
or UO_1477 (O_1477,N_7949,N_8140);
and UO_1478 (O_1478,N_6411,N_8816);
nand UO_1479 (O_1479,N_8058,N_7562);
nor UO_1480 (O_1480,N_9405,N_6584);
nor UO_1481 (O_1481,N_9372,N_7853);
nor UO_1482 (O_1482,N_5055,N_5623);
or UO_1483 (O_1483,N_5934,N_5101);
and UO_1484 (O_1484,N_8452,N_5033);
nand UO_1485 (O_1485,N_9947,N_5294);
and UO_1486 (O_1486,N_8160,N_7771);
or UO_1487 (O_1487,N_9760,N_9228);
nand UO_1488 (O_1488,N_9622,N_8859);
nand UO_1489 (O_1489,N_8241,N_9924);
nand UO_1490 (O_1490,N_5300,N_8034);
nor UO_1491 (O_1491,N_5227,N_6531);
nor UO_1492 (O_1492,N_6316,N_8237);
or UO_1493 (O_1493,N_8822,N_7443);
nand UO_1494 (O_1494,N_5872,N_5192);
or UO_1495 (O_1495,N_9992,N_8820);
or UO_1496 (O_1496,N_6142,N_9710);
and UO_1497 (O_1497,N_6285,N_6222);
or UO_1498 (O_1498,N_6942,N_8747);
nand UO_1499 (O_1499,N_8611,N_6472);
endmodule