module basic_2500_25000_3000_40_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1931,In_477);
and U1 (N_1,In_1681,In_1440);
or U2 (N_2,In_336,In_319);
or U3 (N_3,In_1401,In_657);
nor U4 (N_4,In_485,In_1067);
nand U5 (N_5,In_719,In_1791);
or U6 (N_6,In_127,In_1157);
nor U7 (N_7,In_1825,In_1060);
or U8 (N_8,In_1322,In_1366);
and U9 (N_9,In_637,In_766);
or U10 (N_10,In_2125,In_242);
or U11 (N_11,In_1611,In_681);
and U12 (N_12,In_1076,In_850);
and U13 (N_13,In_1698,In_1985);
nand U14 (N_14,In_2299,In_824);
nand U15 (N_15,In_356,In_2457);
and U16 (N_16,In_22,In_411);
or U17 (N_17,In_2308,In_1237);
nand U18 (N_18,In_1392,In_1797);
or U19 (N_19,In_1396,In_1559);
and U20 (N_20,In_1566,In_1804);
nand U21 (N_21,In_2316,In_1318);
nand U22 (N_22,In_1297,In_148);
nand U23 (N_23,In_2398,In_2350);
nand U24 (N_24,In_1494,In_941);
xor U25 (N_25,In_865,In_1350);
nor U26 (N_26,In_1178,In_2216);
nand U27 (N_27,In_497,In_545);
or U28 (N_28,In_986,In_1997);
nand U29 (N_29,In_1296,In_1563);
xor U30 (N_30,In_770,In_555);
nor U31 (N_31,In_483,In_2315);
xnor U32 (N_32,In_1064,In_2245);
and U33 (N_33,In_2301,In_2082);
and U34 (N_34,In_1764,In_1195);
nor U35 (N_35,In_2377,In_2422);
or U36 (N_36,In_1523,In_2077);
nand U37 (N_37,In_1805,In_2184);
and U38 (N_38,In_1735,In_570);
nand U39 (N_39,In_392,In_2237);
nor U40 (N_40,In_458,In_358);
or U41 (N_41,In_1189,In_325);
and U42 (N_42,In_916,In_952);
and U43 (N_43,In_634,In_1836);
nand U44 (N_44,In_1204,In_1635);
nand U45 (N_45,In_2272,In_1705);
xnor U46 (N_46,In_1678,In_466);
or U47 (N_47,In_1348,In_1128);
xor U48 (N_48,In_665,In_1096);
nor U49 (N_49,In_843,In_1453);
nand U50 (N_50,In_1338,In_1818);
nor U51 (N_51,In_767,In_1225);
and U52 (N_52,In_80,In_408);
nand U53 (N_53,In_1715,In_167);
nand U54 (N_54,In_2265,In_2145);
nand U55 (N_55,In_895,In_396);
and U56 (N_56,In_1487,In_2415);
nor U57 (N_57,In_1892,In_321);
nand U58 (N_58,In_1493,In_1268);
xor U59 (N_59,In_1551,In_1267);
nand U60 (N_60,In_1404,In_974);
or U61 (N_61,In_1066,In_2179);
or U62 (N_62,In_513,In_1826);
nor U63 (N_63,In_1187,In_2343);
and U64 (N_64,In_2417,In_2222);
nand U65 (N_65,In_2273,In_654);
xnor U66 (N_66,In_2318,In_697);
or U67 (N_67,In_2193,In_970);
or U68 (N_68,In_1679,In_430);
xor U69 (N_69,In_1008,In_1053);
nor U70 (N_70,In_1755,In_2102);
xor U71 (N_71,In_2493,In_825);
or U72 (N_72,In_103,In_2100);
or U73 (N_73,In_1378,In_2479);
or U74 (N_74,In_2263,In_344);
and U75 (N_75,In_995,In_712);
nor U76 (N_76,In_1722,In_1479);
nand U77 (N_77,In_1449,In_2136);
nor U78 (N_78,In_1936,In_448);
and U79 (N_79,In_181,In_734);
or U80 (N_80,In_1704,In_1007);
nand U81 (N_81,In_2076,In_1358);
nor U82 (N_82,In_568,In_1497);
nor U83 (N_83,In_1245,In_1146);
nor U84 (N_84,In_1240,In_786);
and U85 (N_85,In_357,In_273);
nand U86 (N_86,In_214,In_937);
nand U87 (N_87,In_2135,In_1622);
nand U88 (N_88,In_1063,In_439);
or U89 (N_89,In_446,In_2049);
nand U90 (N_90,In_1749,In_1552);
or U91 (N_91,In_769,In_2058);
nand U92 (N_92,In_2367,In_1871);
nand U93 (N_93,In_2293,In_1044);
nand U94 (N_94,In_1671,In_2099);
nor U95 (N_95,In_2383,In_1959);
xnor U96 (N_96,In_2170,In_364);
and U97 (N_97,In_2023,In_1921);
nor U98 (N_98,In_2014,In_428);
nand U99 (N_99,In_2161,In_581);
nand U100 (N_100,In_1484,In_2194);
nand U101 (N_101,In_302,In_2494);
nor U102 (N_102,In_924,In_2052);
nand U103 (N_103,In_1317,In_1615);
or U104 (N_104,In_514,In_122);
nor U105 (N_105,In_136,In_94);
xor U106 (N_106,In_1475,In_1238);
nor U107 (N_107,In_280,In_30);
nand U108 (N_108,In_1284,In_915);
or U109 (N_109,In_1359,In_226);
or U110 (N_110,In_363,In_1107);
and U111 (N_111,In_297,In_388);
nor U112 (N_112,In_1194,In_1606);
or U113 (N_113,In_49,In_999);
and U114 (N_114,In_2064,In_487);
xnor U115 (N_115,In_417,In_849);
and U116 (N_116,In_2458,In_1380);
nor U117 (N_117,In_909,In_700);
or U118 (N_118,In_1160,In_1213);
and U119 (N_119,In_1341,In_1036);
nor U120 (N_120,In_1148,In_276);
xnor U121 (N_121,In_830,In_291);
nand U122 (N_122,In_899,In_2406);
nand U123 (N_123,In_609,In_1455);
xnor U124 (N_124,In_1032,In_1999);
or U125 (N_125,In_1618,In_1221);
or U126 (N_126,In_1509,In_1945);
and U127 (N_127,In_979,In_589);
or U128 (N_128,In_531,In_1336);
or U129 (N_129,In_1201,In_1402);
and U130 (N_130,In_2248,In_710);
nor U131 (N_131,In_1423,In_313);
or U132 (N_132,In_126,In_510);
or U133 (N_133,In_1695,In_1773);
nor U134 (N_134,In_1236,In_1332);
and U135 (N_135,In_1387,In_573);
nor U136 (N_136,In_535,In_1939);
nor U137 (N_137,In_761,In_81);
nand U138 (N_138,In_572,In_1644);
nor U139 (N_139,In_832,In_40);
nand U140 (N_140,In_402,In_2238);
nand U141 (N_141,In_1726,In_1090);
xnor U142 (N_142,In_1300,In_542);
and U143 (N_143,In_1272,In_1271);
nor U144 (N_144,In_1048,In_947);
nand U145 (N_145,In_473,In_1521);
nand U146 (N_146,In_1771,In_2017);
nand U147 (N_147,In_1820,In_1287);
nor U148 (N_148,In_566,In_1576);
or U149 (N_149,In_2478,In_853);
and U150 (N_150,In_966,In_1688);
nor U151 (N_151,In_2464,In_1274);
and U152 (N_152,In_2427,In_921);
nand U153 (N_153,In_86,In_595);
or U154 (N_154,In_1646,In_359);
or U155 (N_155,In_1210,In_2385);
nor U156 (N_156,In_746,In_2304);
nor U157 (N_157,In_375,In_162);
and U158 (N_158,In_1185,In_2234);
nor U159 (N_159,In_1376,In_471);
xnor U160 (N_160,In_2499,In_2280);
or U161 (N_161,In_164,In_2053);
nand U162 (N_162,In_1621,In_1425);
or U163 (N_163,In_1321,In_757);
nor U164 (N_164,In_268,In_349);
nor U165 (N_165,In_2462,In_1909);
nand U166 (N_166,In_1207,In_37);
nand U167 (N_167,In_1811,In_1544);
nand U168 (N_168,In_333,In_797);
nand U169 (N_169,In_2470,In_2105);
or U170 (N_170,In_119,In_2192);
and U171 (N_171,In_1460,In_1697);
nor U172 (N_172,In_78,In_106);
nor U173 (N_173,In_1738,In_2071);
or U174 (N_174,In_274,In_348);
or U175 (N_175,In_168,In_2101);
and U176 (N_176,In_2331,In_1492);
nor U177 (N_177,In_737,In_2405);
xor U178 (N_178,In_1441,In_685);
and U179 (N_179,In_586,In_2492);
nand U180 (N_180,In_1188,In_295);
or U181 (N_181,In_1609,In_166);
nor U182 (N_182,In_1205,In_722);
or U183 (N_183,In_2412,In_58);
and U184 (N_184,In_46,In_1311);
or U185 (N_185,In_42,In_331);
or U186 (N_186,In_1760,In_2460);
xnor U187 (N_187,In_2376,In_1852);
nor U188 (N_188,In_1897,In_97);
or U189 (N_189,In_0,In_1962);
nor U190 (N_190,In_1528,In_1718);
nor U191 (N_191,In_138,In_1355);
and U192 (N_192,In_1578,In_1694);
and U193 (N_193,In_1729,In_2190);
xor U194 (N_194,In_1292,In_1776);
nand U195 (N_195,In_2075,In_109);
nor U196 (N_196,In_306,In_640);
or U197 (N_197,In_2452,In_2418);
or U198 (N_198,In_2243,In_1168);
and U199 (N_199,In_118,In_311);
nor U200 (N_200,In_2326,In_957);
and U201 (N_201,In_83,In_845);
or U202 (N_202,In_869,In_582);
or U203 (N_203,In_1361,In_217);
nor U204 (N_204,In_253,In_669);
or U205 (N_205,In_1957,In_1742);
nand U206 (N_206,In_194,In_277);
or U207 (N_207,In_594,In_1603);
and U208 (N_208,In_1416,In_264);
nor U209 (N_209,In_1540,In_1106);
nor U210 (N_210,In_1250,In_1186);
nor U211 (N_211,In_725,In_1877);
and U212 (N_212,In_2208,In_744);
nor U213 (N_213,In_884,In_1581);
or U214 (N_214,In_1758,In_1261);
and U215 (N_215,In_1982,In_1410);
nand U216 (N_216,In_1613,In_171);
and U217 (N_217,In_1518,In_1277);
or U218 (N_218,In_1279,In_1354);
and U219 (N_219,In_32,In_678);
nor U220 (N_220,In_147,In_115);
or U221 (N_221,In_632,In_2340);
nor U222 (N_222,In_2404,In_1333);
xor U223 (N_223,In_2291,In_900);
and U224 (N_224,In_1232,In_316);
or U225 (N_225,In_2081,In_702);
nand U226 (N_226,In_2371,In_985);
and U227 (N_227,In_775,In_1550);
nor U228 (N_228,In_1055,In_879);
and U229 (N_229,In_837,In_1143);
and U230 (N_230,In_796,In_2109);
xor U231 (N_231,In_113,In_384);
nand U232 (N_232,In_2374,In_2360);
or U233 (N_233,In_1849,In_1794);
and U234 (N_234,In_1601,In_1971);
and U235 (N_235,In_990,In_557);
nor U236 (N_236,In_2410,In_1337);
or U237 (N_237,In_1612,In_793);
nand U238 (N_238,In_1069,In_1905);
or U239 (N_239,In_475,In_263);
or U240 (N_240,In_659,In_728);
or U241 (N_241,In_795,In_499);
nand U242 (N_242,In_826,In_1728);
and U243 (N_243,In_897,In_528);
nand U244 (N_244,In_1424,In_108);
nand U245 (N_245,In_1116,In_1891);
xor U246 (N_246,In_1763,In_29);
or U247 (N_247,In_861,In_765);
and U248 (N_248,In_493,In_523);
nor U249 (N_249,In_21,In_1964);
xor U250 (N_250,In_2096,In_773);
nor U251 (N_251,In_151,In_347);
nand U252 (N_252,In_1687,In_1103);
xor U253 (N_253,In_1832,In_2386);
nor U254 (N_254,In_1020,In_551);
or U255 (N_255,In_1500,In_1364);
and U256 (N_256,In_1113,In_288);
or U257 (N_257,In_836,In_1012);
nor U258 (N_258,In_256,In_2372);
nand U259 (N_259,In_862,In_1054);
nor U260 (N_260,In_2201,In_1122);
and U261 (N_261,In_1806,In_1822);
and U262 (N_262,In_68,In_628);
and U263 (N_263,In_1086,In_1680);
or U264 (N_264,In_548,In_1833);
nand U265 (N_265,In_1046,In_2214);
xor U266 (N_266,In_1912,In_1575);
and U267 (N_267,In_636,In_1556);
or U268 (N_268,In_2408,In_1884);
and U269 (N_269,In_1058,In_1074);
or U270 (N_270,In_2275,In_2338);
xnor U271 (N_271,In_1655,In_1);
nor U272 (N_272,In_991,In_1203);
xor U273 (N_273,In_420,In_1713);
xor U274 (N_274,In_1662,In_2393);
nand U275 (N_275,In_1693,In_1312);
and U276 (N_276,In_526,In_2488);
and U277 (N_277,In_1193,In_2495);
and U278 (N_278,In_426,In_142);
and U279 (N_279,In_1674,In_131);
or U280 (N_280,In_1748,In_498);
nor U281 (N_281,In_2233,In_982);
and U282 (N_282,In_804,In_1065);
and U283 (N_283,In_776,In_2011);
nor U284 (N_284,In_19,In_2031);
or U285 (N_285,In_1691,In_525);
nor U286 (N_286,In_791,In_2251);
and U287 (N_287,In_1451,In_383);
or U288 (N_288,In_445,In_207);
nor U289 (N_289,In_604,In_2468);
nand U290 (N_290,In_2416,In_726);
nor U291 (N_291,In_53,In_1562);
nand U292 (N_292,In_294,In_47);
and U293 (N_293,In_1141,In_2093);
nor U294 (N_294,In_495,In_1673);
or U295 (N_295,In_2313,In_1343);
or U296 (N_296,In_449,In_756);
nand U297 (N_297,In_2029,In_1770);
nand U298 (N_298,In_1281,In_158);
nand U299 (N_299,In_2079,In_1028);
or U300 (N_300,In_1352,In_155);
xnor U301 (N_301,In_529,In_1483);
nand U302 (N_302,In_662,In_976);
and U303 (N_303,In_1088,In_1288);
nand U304 (N_304,In_337,In_907);
or U305 (N_305,In_880,In_2439);
nor U306 (N_306,In_1430,In_543);
xor U307 (N_307,In_1432,In_1216);
xor U308 (N_308,In_1782,In_2483);
and U309 (N_309,In_1286,In_2120);
and U310 (N_310,In_809,In_645);
and U311 (N_311,In_806,In_1981);
or U312 (N_312,In_2039,In_972);
or U313 (N_313,In_2212,In_1541);
or U314 (N_314,In_1363,In_1270);
and U315 (N_315,In_1887,In_1447);
nand U316 (N_316,In_69,In_1672);
or U317 (N_317,In_312,In_1403);
nor U318 (N_318,In_639,In_416);
xnor U319 (N_319,In_431,In_2355);
and U320 (N_320,In_1061,In_889);
nand U321 (N_321,In_2111,In_1880);
or U322 (N_322,In_2176,In_267);
xor U323 (N_323,In_559,In_1158);
nor U324 (N_324,In_2287,In_1014);
nand U325 (N_325,In_2008,In_2080);
or U326 (N_326,In_1428,In_2061);
or U327 (N_327,In_2425,In_36);
or U328 (N_328,In_1934,In_2191);
or U329 (N_329,In_890,In_950);
or U330 (N_330,In_1126,In_215);
or U331 (N_331,In_534,In_2112);
nor U332 (N_332,In_590,In_650);
nand U333 (N_333,In_600,In_1918);
nand U334 (N_334,In_1522,In_2258);
nor U335 (N_335,In_1015,In_2186);
nand U336 (N_336,In_1446,In_1315);
xnor U337 (N_337,In_2220,In_964);
nor U338 (N_338,In_1434,In_282);
and U339 (N_339,In_2354,In_1724);
nor U340 (N_340,In_1040,In_2210);
nand U341 (N_341,In_183,In_554);
xnor U342 (N_342,In_1098,In_1789);
or U343 (N_343,In_803,In_1331);
nor U344 (N_344,In_783,In_868);
nand U345 (N_345,In_1623,In_701);
xnor U346 (N_346,In_1374,In_1263);
and U347 (N_347,In_456,In_1725);
nor U348 (N_348,In_309,In_2140);
nand U349 (N_349,In_1802,In_230);
and U350 (N_350,In_1645,In_1996);
and U351 (N_351,In_1056,In_2207);
or U352 (N_352,In_1235,In_633);
or U353 (N_353,In_1173,In_1083);
xor U354 (N_354,In_829,In_460);
and U355 (N_355,In_1377,In_827);
and U356 (N_356,In_2379,In_52);
xnor U357 (N_357,In_1745,In_77);
xor U358 (N_358,In_1721,In_1535);
or U359 (N_359,In_193,In_476);
or U360 (N_360,In_1133,In_1327);
nor U361 (N_361,In_1913,In_1369);
or U362 (N_362,In_720,In_896);
and U363 (N_363,In_31,In_926);
or U364 (N_364,In_2087,In_2228);
nand U365 (N_365,In_1382,In_1654);
and U366 (N_366,In_128,In_942);
and U367 (N_367,In_1488,In_258);
xor U368 (N_368,In_24,In_249);
nand U369 (N_369,In_35,In_187);
nand U370 (N_370,In_1843,In_1436);
nand U371 (N_371,In_851,In_782);
nor U372 (N_372,In_538,In_928);
nor U373 (N_373,In_904,In_1180);
and U374 (N_374,In_2158,In_1457);
and U375 (N_375,In_778,In_2188);
and U376 (N_376,In_1515,In_1587);
and U377 (N_377,In_847,In_661);
or U378 (N_378,In_1491,In_1386);
nand U379 (N_379,In_1524,In_57);
nand U380 (N_380,In_1254,In_211);
nor U381 (N_381,In_2142,In_434);
nand U382 (N_382,In_1591,In_2348);
nor U383 (N_383,In_2336,In_262);
or U384 (N_384,In_1313,In_2231);
and U385 (N_385,In_315,In_104);
or U386 (N_386,In_891,In_1192);
nor U387 (N_387,In_2303,In_62);
nand U388 (N_388,In_2341,In_386);
nor U389 (N_389,In_2068,In_1946);
and U390 (N_390,In_1823,In_703);
or U391 (N_391,In_160,In_2467);
and U392 (N_392,In_1091,In_620);
or U393 (N_393,In_1616,In_1812);
nor U394 (N_394,In_1231,In_1013);
and U395 (N_395,In_1799,In_839);
or U396 (N_396,In_1035,In_1022);
nand U397 (N_397,In_2226,In_1018);
or U398 (N_398,In_26,In_1970);
or U399 (N_399,In_2115,In_1876);
nand U400 (N_400,In_354,In_1372);
or U401 (N_401,In_680,In_2373);
and U402 (N_402,In_79,In_1075);
or U403 (N_403,In_1172,In_2388);
or U404 (N_404,In_1870,In_196);
nand U405 (N_405,In_1206,In_1628);
nand U406 (N_406,In_1114,In_1025);
nand U407 (N_407,In_980,In_292);
nand U408 (N_408,In_672,In_963);
xnor U409 (N_409,In_1998,In_742);
nand U410 (N_410,In_129,In_1775);
nor U411 (N_411,In_1458,In_614);
and U412 (N_412,In_2169,In_2289);
nor U413 (N_413,In_781,In_2054);
nor U414 (N_414,In_270,In_124);
nand U415 (N_415,In_1142,In_1659);
nor U416 (N_416,In_721,In_326);
nor U417 (N_417,In_480,In_197);
and U418 (N_418,In_2490,In_2218);
nor U419 (N_419,In_438,In_328);
nand U420 (N_420,In_93,In_500);
nor U421 (N_421,In_2413,In_814);
or U422 (N_422,In_2163,In_222);
or U423 (N_423,In_2453,In_561);
or U424 (N_424,In_823,In_143);
or U425 (N_425,In_1469,In_310);
nor U426 (N_426,In_1191,In_467);
or U427 (N_427,In_741,In_2361);
and U428 (N_428,In_2302,In_421);
and U429 (N_429,In_2127,In_546);
and U430 (N_430,In_875,In_705);
or U431 (N_431,In_1000,In_759);
xnor U432 (N_432,In_318,In_883);
or U433 (N_433,In_812,In_1042);
nor U434 (N_434,In_1077,In_687);
nand U435 (N_435,In_984,In_560);
and U436 (N_436,In_1684,In_810);
nor U437 (N_437,In_121,In_432);
nand U438 (N_438,In_1334,In_125);
or U439 (N_439,In_1765,In_1636);
and U440 (N_440,In_1813,In_652);
nand U441 (N_441,In_43,In_200);
or U442 (N_442,In_265,In_355);
and U443 (N_443,In_2399,In_1001);
nor U444 (N_444,In_1710,In_1490);
nor U445 (N_445,In_178,In_738);
nand U446 (N_446,In_1841,In_2429);
xor U447 (N_447,In_2235,In_1980);
or U448 (N_448,In_1633,In_724);
or U449 (N_449,In_317,In_1778);
nor U450 (N_450,In_1855,In_2268);
and U451 (N_451,In_818,In_1421);
or U452 (N_452,In_735,In_1399);
or U453 (N_453,In_1527,In_2202);
and U454 (N_454,In_474,In_1052);
and U455 (N_455,In_414,In_2187);
nor U456 (N_456,In_1306,In_1564);
and U457 (N_457,In_2156,In_715);
nand U458 (N_458,In_405,In_873);
nand U459 (N_459,In_1246,In_1023);
xor U460 (N_460,In_2365,In_56);
nand U461 (N_461,In_283,In_1149);
or U462 (N_462,In_1147,In_1808);
or U463 (N_463,In_1224,In_1498);
nand U464 (N_464,In_1070,In_989);
nand U465 (N_465,In_983,In_1648);
nor U466 (N_466,In_2271,In_1439);
nor U467 (N_467,In_578,In_339);
and U468 (N_468,In_208,In_539);
and U469 (N_469,In_1394,In_1124);
nand U470 (N_470,In_1426,In_1156);
or U471 (N_471,In_2421,In_1640);
and U472 (N_472,In_1928,In_1031);
nand U473 (N_473,In_1507,In_2284);
nand U474 (N_474,In_287,In_244);
xor U475 (N_475,In_1166,In_404);
and U476 (N_476,In_699,In_507);
nor U477 (N_477,In_395,In_565);
and U478 (N_478,In_1754,In_2329);
nor U479 (N_479,In_1155,In_2324);
nand U480 (N_480,In_1129,In_2349);
nand U481 (N_481,In_1907,In_682);
xnor U482 (N_482,In_754,In_1427);
and U483 (N_483,In_236,In_2062);
or U484 (N_484,In_758,In_1257);
nand U485 (N_485,In_468,In_919);
nand U486 (N_486,In_1125,In_1164);
or U487 (N_487,In_615,In_1516);
and U488 (N_488,In_452,In_1072);
nand U489 (N_489,In_472,In_2072);
or U490 (N_490,In_1783,In_1227);
or U491 (N_491,In_1711,In_1630);
nor U492 (N_492,In_727,In_2083);
and U493 (N_493,In_1381,In_260);
nor U494 (N_494,In_651,In_603);
or U495 (N_495,In_478,In_1838);
nand U496 (N_496,In_2476,In_149);
nand U497 (N_497,In_2141,In_973);
nand U498 (N_498,In_1223,In_303);
nor U499 (N_499,In_2409,In_1112);
nor U500 (N_500,In_2482,In_815);
nor U501 (N_501,In_1480,In_1229);
nand U502 (N_502,In_2276,In_360);
nand U503 (N_503,In_1159,In_406);
nor U504 (N_504,In_1894,In_1796);
xor U505 (N_505,In_2314,In_2042);
xor U506 (N_506,In_1809,In_73);
nand U507 (N_507,In_1130,In_1935);
xor U508 (N_508,In_1627,In_911);
nor U509 (N_509,In_110,In_1239);
xnor U510 (N_510,In_346,In_229);
nand U511 (N_511,In_944,In_2025);
nand U512 (N_512,In_2021,In_23);
and U513 (N_513,In_413,In_1733);
nor U514 (N_514,In_382,In_592);
nor U515 (N_515,In_367,In_1686);
or U516 (N_516,In_1743,In_1208);
nand U517 (N_517,In_1526,In_1356);
and U518 (N_518,In_1389,In_2198);
nor U519 (N_519,In_1269,In_771);
xnor U520 (N_520,In_1202,In_1226);
and U521 (N_521,In_1006,In_693);
and U522 (N_522,In_6,In_1730);
nand U523 (N_523,In_874,In_801);
and U524 (N_524,In_1873,In_141);
or U525 (N_525,In_1118,In_2209);
and U526 (N_526,In_1739,In_1251);
and U527 (N_527,In_1624,In_1976);
nor U528 (N_528,In_1991,In_925);
or U529 (N_529,In_1212,In_54);
xor U530 (N_530,In_718,In_2330);
and U531 (N_531,In_1198,In_2246);
nand U532 (N_532,In_1955,In_2262);
xnor U533 (N_533,In_453,In_2390);
or U534 (N_534,In_2426,In_2297);
or U535 (N_535,In_1868,In_170);
and U536 (N_536,In_191,In_707);
nand U537 (N_537,In_401,In_1740);
and U538 (N_538,In_394,In_863);
nand U539 (N_539,In_717,In_1407);
and U540 (N_540,In_623,In_1099);
or U541 (N_541,In_1585,In_673);
nor U542 (N_542,In_1276,In_25);
or U543 (N_543,In_1136,In_893);
or U544 (N_544,In_2183,In_596);
or U545 (N_545,In_2244,In_3);
nor U546 (N_546,In_1105,In_2300);
and U547 (N_547,In_114,In_247);
nand U548 (N_548,In_576,In_550);
or U549 (N_549,In_1506,In_2040);
nand U550 (N_550,In_1429,In_107);
nor U551 (N_551,In_532,In_1081);
and U552 (N_552,In_1625,In_329);
or U553 (N_553,In_1779,In_1266);
and U554 (N_554,In_2382,In_8);
nand U555 (N_555,In_642,In_1154);
nor U556 (N_556,In_1360,In_2463);
and U557 (N_557,In_789,In_1512);
xnor U558 (N_558,In_1406,In_1958);
xor U559 (N_559,In_747,In_502);
nand U560 (N_560,In_1917,In_271);
and U561 (N_561,In_975,In_1395);
nor U562 (N_562,In_1496,In_1417);
and U563 (N_563,In_1309,In_50);
and U564 (N_564,In_1589,In_1339);
and U565 (N_565,In_1438,In_366);
or U566 (N_566,In_479,In_2414);
xor U567 (N_567,In_99,In_2197);
and U568 (N_568,In_1335,In_1474);
or U569 (N_569,In_1788,In_690);
nor U570 (N_570,In_1769,In_1408);
nand U571 (N_571,In_1340,In_856);
and U572 (N_572,In_1570,In_2279);
nand U573 (N_573,In_255,In_1259);
nand U574 (N_574,In_1824,In_393);
or U575 (N_575,In_1599,In_2143);
and U576 (N_576,In_192,In_1415);
and U577 (N_577,In_788,In_956);
and U578 (N_578,In_463,In_923);
and U579 (N_579,In_190,In_2146);
xor U580 (N_580,In_962,In_1119);
or U581 (N_581,In_484,In_133);
and U582 (N_582,In_1600,In_2449);
and U583 (N_583,In_307,In_71);
or U584 (N_584,In_1911,In_353);
and U585 (N_585,In_1741,In_13);
nand U586 (N_586,In_7,In_2116);
or U587 (N_587,In_1508,In_1466);
or U588 (N_588,In_1353,In_2144);
nand U589 (N_589,In_1853,In_1561);
nand U590 (N_590,In_1533,In_1567);
nand U591 (N_591,In_993,In_648);
xnor U592 (N_592,In_2091,In_1298);
nor U593 (N_593,In_351,In_1829);
or U594 (N_594,In_848,In_1720);
nor U595 (N_595,In_2173,In_2257);
nand U596 (N_596,In_2441,In_2126);
xnor U597 (N_597,In_1167,In_1727);
nor U598 (N_598,In_522,In_2497);
or U599 (N_599,In_298,In_2496);
nor U600 (N_600,In_1850,In_14);
nor U601 (N_601,In_1950,In_503);
or U602 (N_602,In_1151,In_1247);
nand U603 (N_603,In_1846,In_1972);
nand U604 (N_604,In_286,In_949);
nor U605 (N_605,In_218,In_409);
nor U606 (N_606,In_1021,In_1594);
or U607 (N_607,In_506,In_1568);
nor U608 (N_608,In_465,In_1273);
nor U609 (N_609,In_1073,In_324);
nor U610 (N_610,In_641,In_1039);
nor U611 (N_611,In_655,In_1647);
nor U612 (N_612,In_1643,In_1790);
nand U613 (N_613,In_2151,In_140);
or U614 (N_614,In_1121,In_2148);
nor U615 (N_615,In_2319,In_48);
and U616 (N_616,In_605,In_2149);
and U617 (N_617,In_1943,In_1304);
or U618 (N_618,In_1951,In_120);
nor U619 (N_619,In_508,In_1653);
and U620 (N_620,In_914,In_188);
or U621 (N_621,In_55,In_340);
xor U622 (N_622,In_1127,In_216);
or U623 (N_623,In_2094,In_1089);
xor U624 (N_624,In_945,In_1637);
or U625 (N_625,In_1165,In_959);
and U626 (N_626,In_1784,In_1450);
nor U627 (N_627,In_2078,In_1736);
nor U628 (N_628,In_338,In_2380);
and U629 (N_629,In_1546,In_1351);
or U630 (N_630,In_1176,In_1530);
nor U631 (N_631,In_2147,In_1470);
nand U632 (N_632,In_1889,In_1803);
and U633 (N_633,In_1702,In_213);
and U634 (N_634,N_457,In_75);
nor U635 (N_635,In_1283,In_2339);
xnor U636 (N_636,In_2001,In_2255);
xor U637 (N_637,N_141,In_2305);
nor U638 (N_638,In_1329,N_151);
nor U639 (N_639,In_2403,In_987);
or U640 (N_640,In_2043,In_482);
nor U641 (N_641,In_1017,In_802);
and U642 (N_642,In_1639,In_549);
or U643 (N_643,In_2381,In_2098);
or U644 (N_644,In_2138,In_1983);
nand U645 (N_645,N_163,In_2213);
or U646 (N_646,In_1752,N_363);
or U647 (N_647,In_2278,N_11);
nor U648 (N_648,In_784,In_1255);
or U649 (N_649,In_1330,In_1893);
xnor U650 (N_650,In_794,In_38);
nor U651 (N_651,In_1316,In_597);
xor U652 (N_652,N_187,N_477);
or U653 (N_653,In_1463,In_2298);
nor U654 (N_654,N_145,N_27);
or U655 (N_655,In_464,N_362);
or U656 (N_656,In_2137,In_635);
and U657 (N_657,N_10,In_2165);
nor U658 (N_658,In_965,In_1839);
nand U659 (N_659,In_777,N_456);
nor U660 (N_660,N_416,N_267);
nand U661 (N_661,N_459,N_7);
nand U662 (N_662,In_1875,In_1517);
and U663 (N_663,In_939,N_123);
nand U664 (N_664,In_521,In_1869);
and U665 (N_665,In_199,N_138);
xor U666 (N_666,In_1898,In_1062);
or U667 (N_667,N_343,In_516);
nor U668 (N_668,N_67,In_1365);
and U669 (N_669,In_656,N_23);
nand U670 (N_670,In_1026,In_934);
or U671 (N_671,In_1454,In_219);
or U672 (N_672,In_1750,N_94);
nor U673 (N_673,In_616,In_204);
xnor U674 (N_674,In_2060,In_332);
nand U675 (N_675,In_85,In_692);
and U676 (N_676,In_1933,In_1471);
nor U677 (N_677,In_1104,In_1840);
nor U678 (N_678,In_2312,N_40);
nand U679 (N_679,N_566,N_367);
xor U680 (N_680,In_1501,N_212);
nand U681 (N_681,In_1994,In_1071);
nand U682 (N_682,In_2407,In_1218);
nand U683 (N_683,In_1320,N_481);
nor U684 (N_684,In_1431,In_2035);
nand U685 (N_685,In_2356,In_447);
and U686 (N_686,In_958,N_329);
and U687 (N_687,N_518,In_87);
and U688 (N_688,N_400,In_2437);
xor U689 (N_689,N_178,N_89);
xor U690 (N_690,N_394,N_31);
and U691 (N_691,In_1610,In_1258);
and U692 (N_692,N_374,In_1656);
nand U693 (N_693,In_932,N_517);
and U694 (N_694,N_135,In_227);
xor U695 (N_695,In_2095,In_259);
nand U696 (N_696,In_1572,In_1984);
or U697 (N_697,In_2000,N_238);
and U698 (N_698,In_1514,N_304);
nor U699 (N_699,In_330,N_217);
and U700 (N_700,In_252,In_2431);
nand U701 (N_701,In_1793,In_1759);
nand U702 (N_702,In_1029,In_407);
and U703 (N_703,In_1677,In_902);
or U704 (N_704,N_101,In_1941);
nor U705 (N_705,In_683,In_1511);
nor U706 (N_706,In_289,N_478);
nor U707 (N_707,N_25,In_704);
nand U708 (N_708,N_480,In_1828);
nand U709 (N_709,In_1414,In_492);
nand U710 (N_710,N_196,N_97);
or U711 (N_711,In_601,In_1989);
or U712 (N_712,N_544,N_202);
or U713 (N_713,In_1465,N_58);
nor U714 (N_714,In_1700,In_1649);
xor U715 (N_715,In_41,In_706);
and U716 (N_716,N_124,N_389);
or U717 (N_717,In_1153,In_2059);
or U718 (N_718,In_2387,N_167);
nor U719 (N_719,In_1992,In_870);
and U720 (N_720,In_1660,In_2155);
nor U721 (N_721,In_91,In_370);
and U722 (N_722,In_520,In_658);
and U723 (N_723,In_1370,In_558);
and U724 (N_724,N_179,In_1196);
and U725 (N_725,In_350,N_512);
and U726 (N_726,N_225,In_1177);
nand U727 (N_727,In_1596,N_149);
xnor U728 (N_728,In_165,N_539);
or U729 (N_729,N_264,In_111);
or U730 (N_730,In_198,In_679);
nand U731 (N_731,In_2424,N_222);
nor U732 (N_732,In_1024,In_574);
nand U733 (N_733,In_1590,N_75);
nand U734 (N_734,N_617,In_1145);
nor U735 (N_735,N_491,In_946);
nand U736 (N_736,In_981,N_282);
nand U737 (N_737,N_294,In_708);
xnor U738 (N_738,N_402,N_557);
or U739 (N_739,N_435,N_581);
and U740 (N_740,N_476,In_2241);
nand U741 (N_741,N_615,In_768);
or U742 (N_742,In_33,In_246);
and U743 (N_743,In_410,In_1398);
nand U744 (N_744,N_551,In_1282);
or U745 (N_745,In_2362,In_156);
or U746 (N_746,In_663,N_610);
nand U747 (N_747,In_1938,In_1707);
and U748 (N_748,N_513,In_1050);
or U749 (N_749,In_1816,In_5);
and U750 (N_750,N_467,N_601);
xor U751 (N_751,N_338,N_586);
nor U752 (N_752,In_1302,In_977);
nor U753 (N_753,In_257,N_39);
nor U754 (N_754,In_1731,In_2357);
nor U755 (N_755,In_66,N_79);
and U756 (N_756,N_391,In_1097);
nor U757 (N_757,In_748,In_1041);
nor U758 (N_758,N_208,In_1844);
nor U759 (N_759,In_1642,In_2123);
or U760 (N_760,In_1792,N_228);
nor U761 (N_761,N_414,In_1144);
xnor U762 (N_762,N_560,In_689);
and U763 (N_763,In_2166,In_76);
and U764 (N_764,In_2443,N_351);
and U765 (N_765,In_612,In_1882);
and U766 (N_766,In_2344,In_619);
and U767 (N_767,N_26,In_2139);
or U768 (N_768,In_179,In_835);
or U769 (N_769,N_144,In_1966);
nand U770 (N_770,In_2204,In_674);
and U771 (N_771,In_1027,In_2267);
nor U772 (N_772,In_1766,In_910);
or U773 (N_773,N_364,In_2065);
nor U774 (N_774,N_100,N_538);
nand U775 (N_775,In_2332,N_256);
nor U776 (N_776,In_611,N_440);
and U777 (N_777,N_419,In_1885);
or U778 (N_778,In_1293,In_2113);
nand U779 (N_779,In_1045,In_2428);
and U780 (N_780,In_992,In_2456);
nor U781 (N_781,N_587,In_284);
and U782 (N_782,N_112,N_170);
or U783 (N_783,N_583,N_327);
and U784 (N_784,In_2285,In_1448);
and U785 (N_785,N_474,N_137);
xor U786 (N_786,N_69,In_2046);
nand U787 (N_787,In_2402,In_1375);
and U788 (N_788,N_537,N_501);
nand U789 (N_789,N_511,In_820);
or U790 (N_790,In_800,N_608);
or U791 (N_791,In_39,In_562);
and U792 (N_792,In_838,In_1233);
or U793 (N_793,In_2436,In_308);
and U794 (N_794,N_563,In_2175);
nand U795 (N_795,In_281,In_515);
nand U796 (N_796,In_300,N_623);
xnor U797 (N_797,N_281,In_1362);
nor U798 (N_798,In_261,In_1602);
or U799 (N_799,In_1683,In_1010);
nand U800 (N_800,In_1478,N_115);
nor U801 (N_801,In_948,In_2092);
xnor U802 (N_802,N_54,In_567);
nor U803 (N_803,N_326,In_1435);
nor U804 (N_804,N_430,N_52);
and U805 (N_805,N_98,In_67);
nand U806 (N_806,In_1965,In_2445);
or U807 (N_807,In_785,N_312);
or U808 (N_808,In_2469,N_372);
xnor U809 (N_809,N_542,In_1379);
nor U810 (N_810,In_1472,In_1459);
nor U811 (N_811,In_1452,In_1510);
nor U812 (N_812,In_2178,In_1947);
nor U813 (N_813,N_356,In_1111);
xor U814 (N_814,In_1299,In_1214);
or U815 (N_815,In_369,In_221);
or U816 (N_816,In_527,In_1902);
nor U817 (N_817,In_4,In_998);
nand U818 (N_818,In_1685,In_2172);
or U819 (N_819,N_531,N_572);
and U820 (N_820,In_1139,In_713);
or U821 (N_821,In_442,In_1916);
or U822 (N_822,N_96,N_74);
and U823 (N_823,In_2107,In_1100);
xnor U824 (N_824,N_558,In_2004);
nand U825 (N_825,N_411,N_287);
or U826 (N_826,In_1264,In_2007);
or U827 (N_827,In_1604,In_2327);
and U828 (N_828,In_1413,In_385);
nand U829 (N_829,In_1692,In_1047);
or U830 (N_830,In_1301,In_1117);
xor U831 (N_831,N_359,N_505);
or U832 (N_832,In_2384,N_504);
nor U833 (N_833,N_269,In_1732);
and U834 (N_834,In_427,N_197);
nor U835 (N_835,In_1906,In_304);
xor U836 (N_836,In_1819,In_1927);
nand U837 (N_837,In_123,In_729);
or U838 (N_838,In_1979,N_200);
and U839 (N_839,In_1815,In_425);
xnor U840 (N_840,In_1078,In_1930);
or U841 (N_841,N_382,In_2181);
or U842 (N_842,N_139,In_955);
and U843 (N_843,In_2038,N_370);
xnor U844 (N_844,In_2337,In_352);
nand U845 (N_845,In_653,In_696);
or U846 (N_846,N_18,N_395);
xnor U847 (N_847,In_2032,N_22);
or U848 (N_848,In_1565,In_978);
or U849 (N_849,N_331,N_366);
and U850 (N_850,In_1094,N_334);
or U851 (N_851,N_33,In_714);
nor U852 (N_852,In_1038,N_381);
xor U853 (N_853,In_1525,In_1582);
and U854 (N_854,In_169,N_408);
nand U855 (N_855,N_588,In_2288);
nand U856 (N_856,In_1252,N_556);
and U857 (N_857,In_1973,In_234);
xor U858 (N_858,In_1135,In_2162);
and U859 (N_859,In_1346,N_494);
and U860 (N_860,In_100,N_234);
or U861 (N_861,In_322,N_580);
or U862 (N_862,In_1701,N_37);
or U863 (N_863,In_676,In_1504);
nor U864 (N_864,In_1059,In_130);
nand U865 (N_865,N_207,In_1886);
or U866 (N_866,In_2391,In_415);
or U867 (N_867,N_160,In_1954);
nand U868 (N_868,N_516,N_570);
nor U869 (N_869,N_316,N_506);
nand U870 (N_870,In_1170,In_2206);
and U871 (N_871,In_2307,N_297);
nand U872 (N_872,In_2066,N_384);
xor U873 (N_873,In_1342,N_148);
and U874 (N_874,N_360,N_263);
and U875 (N_875,In_811,In_443);
and U876 (N_876,In_967,In_279);
nand U877 (N_877,In_1409,In_1323);
xor U878 (N_878,In_1708,In_1305);
nor U879 (N_879,In_698,In_1520);
and U880 (N_880,In_488,N_130);
and U881 (N_881,In_2033,In_455);
nor U882 (N_882,In_504,N_519);
nand U883 (N_883,N_309,In_2351);
nand U884 (N_884,N_346,N_375);
nor U885 (N_885,In_418,In_1774);
xor U886 (N_886,In_157,N_589);
or U887 (N_887,N_399,In_1102);
and U888 (N_888,N_433,In_1665);
or U889 (N_889,N_348,In_621);
nand U890 (N_890,N_131,In_2203);
and U891 (N_891,N_158,N_447);
nor U892 (N_892,In_1942,In_541);
or U893 (N_893,In_2454,N_547);
nor U894 (N_894,N_607,In_2240);
and U895 (N_895,In_1080,In_2227);
nor U896 (N_896,N_274,In_2430);
or U897 (N_897,In_593,In_1217);
or U898 (N_898,In_245,In_1896);
xor U899 (N_899,In_381,N_515);
xor U900 (N_900,In_2450,In_469);
or U901 (N_901,In_1631,N_262);
nor U902 (N_902,In_174,In_1557);
xor U903 (N_903,In_1495,In_2295);
or U904 (N_904,In_1555,In_371);
and U905 (N_905,In_1549,In_2108);
or U906 (N_906,In_831,N_383);
nand U907 (N_907,N_32,N_192);
nor U908 (N_908,N_578,N_571);
and U909 (N_909,N_247,In_1975);
and U910 (N_910,In_1248,N_0);
nor U911 (N_911,In_1851,N_43);
nor U912 (N_912,In_2466,In_1547);
xor U913 (N_913,N_261,In_1539);
nor U914 (N_914,N_259,In_1230);
and U915 (N_915,In_1974,In_755);
nand U916 (N_916,In_866,In_563);
or U917 (N_917,In_2030,N_559);
and U918 (N_918,In_2420,In_1110);
nand U919 (N_919,In_1747,N_295);
and U920 (N_920,In_599,In_1658);
nor U921 (N_921,In_1291,N_498);
xnor U922 (N_922,N_248,In_647);
or U923 (N_923,In_233,N_114);
xnor U924 (N_924,In_2164,In_429);
nand U925 (N_925,In_1669,In_139);
nor U926 (N_926,N_584,In_2242);
or U927 (N_927,N_604,N_405);
or U928 (N_928,In_235,In_901);
nand U929 (N_929,In_1574,N_64);
nand U930 (N_930,In_2480,In_2160);
nand U931 (N_931,N_219,In_2200);
nand U932 (N_932,In_2006,In_763);
nand U933 (N_933,N_2,In_519);
and U934 (N_934,N_279,In_305);
or U935 (N_935,N_483,In_627);
nand U936 (N_936,In_1904,In_1663);
nor U937 (N_937,In_1101,In_664);
xor U938 (N_938,In_1583,N_596);
or U939 (N_939,In_792,In_1952);
nor U940 (N_940,In_16,N_470);
or U941 (N_941,N_49,N_218);
and U942 (N_942,In_2481,In_2252);
nand U943 (N_943,In_1915,In_1629);
nand U944 (N_944,N_324,In_223);
or U945 (N_945,In_2045,In_2346);
or U946 (N_946,In_20,In_1082);
or U947 (N_947,In_1859,N_308);
or U948 (N_948,In_1593,In_1920);
xor U949 (N_949,N_369,N_183);
nand U950 (N_950,In_1580,N_475);
nand U951 (N_951,In_943,N_466);
or U952 (N_952,N_62,N_428);
nor U953 (N_953,In_940,N_418);
nor U954 (N_954,In_840,N_479);
nand U955 (N_955,In_1542,In_28);
and U956 (N_956,In_285,In_44);
or U957 (N_957,In_1753,In_584);
and U958 (N_958,In_1827,In_1795);
or U959 (N_959,In_2199,In_1347);
nand U960 (N_960,In_580,In_1037);
nand U961 (N_961,In_930,In_2048);
nand U962 (N_962,In_459,In_750);
nand U963 (N_963,N_328,In_585);
and U964 (N_964,In_931,In_1993);
nand U965 (N_965,In_1786,In_971);
or U966 (N_966,In_2369,N_6);
nor U967 (N_967,N_215,N_458);
nor U968 (N_968,In_787,N_70);
nor U969 (N_969,N_520,In_2219);
xor U970 (N_970,In_745,N_301);
nor U971 (N_971,In_2152,N_464);
and U972 (N_972,N_386,In_2317);
or U973 (N_973,In_2097,N_181);
or U974 (N_974,N_83,In_799);
nor U975 (N_975,N_368,In_1641);
xnor U976 (N_976,In_2159,N_336);
and U977 (N_977,In_1184,N_619);
and U978 (N_978,In_2292,In_760);
or U979 (N_979,In_2286,N_550);
nand U980 (N_980,N_317,In_1132);
xnor U981 (N_981,N_299,N_582);
and U982 (N_982,In_1499,In_1482);
xnor U983 (N_983,In_2131,In_1807);
nand U984 (N_984,N_488,In_935);
and U985 (N_985,N_468,N_490);
nand U986 (N_986,N_189,In_583);
nor U987 (N_987,In_2270,N_251);
xor U988 (N_988,N_472,N_499);
nor U989 (N_989,In_2236,N_406);
nand U990 (N_990,N_404,In_1956);
nor U991 (N_991,In_454,In_1243);
or U992 (N_992,In_675,In_423);
nand U993 (N_993,In_2434,N_231);
or U994 (N_994,In_591,In_444);
nor U995 (N_995,In_272,N_165);
and U996 (N_996,In_17,In_2321);
nor U997 (N_997,In_1093,In_1878);
nand U998 (N_998,In_821,N_500);
nor U999 (N_999,In_335,N_485);
and U1000 (N_1000,N_390,N_162);
and U1001 (N_1001,In_1990,In_212);
nor U1002 (N_1002,In_1383,In_1175);
or U1003 (N_1003,In_936,N_453);
and U1004 (N_1004,In_666,N_258);
nor U1005 (N_1005,N_210,In_2073);
and U1006 (N_1006,In_2375,In_649);
nand U1007 (N_1007,N_579,In_1536);
and U1008 (N_1008,In_1411,In_2353);
or U1009 (N_1009,In_1171,N_275);
nand U1010 (N_1010,N_606,In_342);
nand U1011 (N_1011,In_1505,In_1534);
and U1012 (N_1012,In_378,In_2056);
nor U1013 (N_1013,N_357,In_2334);
nand U1014 (N_1014,N_126,In_1368);
or U1015 (N_1015,In_1537,N_339);
or U1016 (N_1016,In_1619,In_2018);
xor U1017 (N_1017,N_120,N_81);
nor U1018 (N_1018,In_2310,N_333);
nand U1019 (N_1019,N_620,In_1308);
xnor U1020 (N_1020,In_210,N_291);
nor U1021 (N_1021,In_101,In_1910);
nor U1022 (N_1022,In_887,N_80);
nor U1023 (N_1023,In_2063,N_482);
nand U1024 (N_1024,N_300,In_243);
nand U1025 (N_1025,In_1714,In_1190);
nor U1026 (N_1026,In_2026,In_808);
and U1027 (N_1027,N_552,In_569);
xnor U1028 (N_1028,In_2010,In_2129);
nor U1029 (N_1029,In_2474,In_2);
xnor U1030 (N_1030,N_310,N_450);
xor U1031 (N_1031,N_451,In_64);
or U1032 (N_1032,In_553,N_169);
nor U1033 (N_1033,In_1737,In_695);
nand U1034 (N_1034,N_3,In_2475);
nand U1035 (N_1035,N_56,In_881);
and U1036 (N_1036,N_448,In_844);
xor U1037 (N_1037,In_1650,N_320);
nand U1038 (N_1038,In_345,N_20);
and U1039 (N_1039,N_593,N_276);
nand U1040 (N_1040,N_93,In_2328);
and U1041 (N_1041,In_1588,N_1);
or U1042 (N_1042,In_2446,In_1543);
nor U1043 (N_1043,In_1473,N_42);
nor U1044 (N_1044,In_1638,In_954);
xnor U1045 (N_1045,In_2486,In_1123);
and U1046 (N_1046,In_2232,In_918);
and U1047 (N_1047,In_1883,In_2005);
and U1048 (N_1048,N_443,In_2223);
and U1049 (N_1049,N_307,In_1923);
nand U1050 (N_1050,N_214,N_455);
xnor U1051 (N_1051,In_1932,In_969);
nor U1052 (N_1052,In_2333,In_1513);
nor U1053 (N_1053,In_1706,In_1162);
or U1054 (N_1054,N_51,N_413);
or U1055 (N_1055,In_1467,N_224);
or U1056 (N_1056,In_575,In_1131);
nor U1057 (N_1057,In_852,In_2309);
and U1058 (N_1058,N_44,In_184);
nand U1059 (N_1059,In_1837,N_599);
nor U1060 (N_1060,In_225,In_2448);
nor U1061 (N_1061,N_103,In_278);
or U1062 (N_1062,In_172,In_1005);
and U1063 (N_1063,N_407,In_2320);
and U1064 (N_1064,In_1242,In_624);
xnor U1065 (N_1065,In_2358,In_2086);
nor U1066 (N_1066,In_805,N_146);
and U1067 (N_1067,N_420,In_2133);
nor U1068 (N_1068,In_739,In_18);
nand U1069 (N_1069,In_1831,N_355);
nor U1070 (N_1070,In_2342,N_352);
nand U1071 (N_1071,N_541,N_439);
and U1072 (N_1072,In_2306,In_2366);
nand U1073 (N_1073,N_201,In_857);
or U1074 (N_1074,In_892,N_527);
or U1075 (N_1075,In_953,In_643);
and U1076 (N_1076,N_220,In_2378);
nor U1077 (N_1077,In_2047,N_618);
xor U1078 (N_1078,In_398,N_590);
and U1079 (N_1079,In_1834,N_223);
and U1080 (N_1080,N_161,In_2411);
or U1081 (N_1081,N_84,In_1260);
nand U1082 (N_1082,N_595,In_231);
nor U1083 (N_1083,In_2168,In_323);
and U1084 (N_1084,N_342,In_2037);
and U1085 (N_1085,In_88,In_399);
xnor U1086 (N_1086,In_1872,In_1614);
xnor U1087 (N_1087,N_122,N_305);
nor U1088 (N_1088,N_344,N_271);
nor U1089 (N_1089,In_1757,In_512);
or U1090 (N_1090,In_1057,In_2019);
and U1091 (N_1091,In_368,In_314);
nor U1092 (N_1092,N_545,N_592);
xor U1093 (N_1093,In_59,In_1987);
and U1094 (N_1094,N_268,N_12);
xor U1095 (N_1095,In_716,In_1967);
nand U1096 (N_1096,N_171,In_1179);
nor U1097 (N_1097,N_315,In_299);
nor U1098 (N_1098,In_2260,N_330);
nor U1099 (N_1099,In_876,In_1503);
nor U1100 (N_1100,N_533,N_216);
and U1101 (N_1101,In_1456,N_432);
nor U1102 (N_1102,In_610,In_885);
or U1103 (N_1103,In_1961,In_501);
nor U1104 (N_1104,In_1888,In_1011);
nor U1105 (N_1105,N_495,N_422);
or U1106 (N_1106,N_36,In_2130);
and U1107 (N_1107,N_446,N_117);
xnor U1108 (N_1108,In_1785,In_908);
or U1109 (N_1109,In_1095,In_72);
nand U1110 (N_1110,In_2189,In_1349);
nand U1111 (N_1111,In_1800,In_733);
nor U1112 (N_1112,In_2195,In_730);
nor U1113 (N_1113,In_241,In_1777);
nand U1114 (N_1114,N_345,In_2364);
nand U1115 (N_1115,In_2121,In_2085);
and U1116 (N_1116,In_1461,In_1548);
and U1117 (N_1117,In_511,N_311);
or U1118 (N_1118,In_1634,In_2274);
nor U1119 (N_1119,N_106,In_1908);
or U1120 (N_1120,In_819,In_906);
nand U1121 (N_1121,N_487,In_2352);
and U1122 (N_1122,N_46,N_230);
and U1123 (N_1123,In_374,In_9);
nor U1124 (N_1124,N_150,In_1437);
nor U1125 (N_1125,In_1262,In_772);
nor U1126 (N_1126,In_1400,In_1901);
xnor U1127 (N_1127,In_1801,In_489);
and U1128 (N_1128,In_182,N_229);
and U1129 (N_1129,In_1385,N_16);
xnor U1130 (N_1130,In_1842,In_556);
nand U1131 (N_1131,In_390,N_561);
or U1132 (N_1132,In_571,In_2110);
nand U1133 (N_1133,N_349,In_1924);
and U1134 (N_1134,In_433,In_2250);
nor U1135 (N_1135,N_116,N_142);
nand U1136 (N_1136,In_301,In_1598);
nor U1137 (N_1137,In_751,In_1294);
nand U1138 (N_1138,In_1068,In_240);
nand U1139 (N_1139,In_376,In_691);
nand U1140 (N_1140,In_618,N_555);
and U1141 (N_1141,N_50,N_340);
nor U1142 (N_1142,In_1554,In_189);
nand U1143 (N_1143,N_48,In_731);
nand U1144 (N_1144,N_403,In_762);
and U1145 (N_1145,In_145,In_1858);
nand U1146 (N_1146,In_422,In_490);
nand U1147 (N_1147,In_743,N_436);
and U1148 (N_1148,In_1845,In_2484);
or U1149 (N_1149,In_95,In_1108);
and U1150 (N_1150,In_1303,In_2185);
or U1151 (N_1151,N_136,In_1289);
and U1152 (N_1152,N_277,N_543);
nor U1153 (N_1153,N_227,N_318);
nand U1154 (N_1154,N_29,In_2363);
nor U1155 (N_1155,N_8,In_1988);
or U1156 (N_1156,In_2359,In_2266);
and U1157 (N_1157,N_353,N_396);
nand U1158 (N_1158,N_575,N_105);
xor U1159 (N_1159,In_1326,In_486);
or U1160 (N_1160,In_1442,N_335);
nor U1161 (N_1161,In_2294,In_709);
xnor U1162 (N_1162,N_401,In_341);
nor U1163 (N_1163,N_452,In_1573);
and U1164 (N_1164,N_605,In_102);
nand U1165 (N_1165,N_57,In_1328);
and U1166 (N_1166,N_426,In_1835);
xnor U1167 (N_1167,In_764,N_204);
nor U1168 (N_1168,In_237,In_552);
nor U1169 (N_1169,In_2335,N_568);
or U1170 (N_1170,In_440,In_644);
nor U1171 (N_1171,In_2106,In_2117);
or U1172 (N_1172,In_2440,In_2498);
or U1173 (N_1173,In_2134,In_1900);
nand U1174 (N_1174,In_1532,N_361);
and U1175 (N_1175,In_1978,In_2461);
nor U1176 (N_1176,In_2455,In_180);
and U1177 (N_1177,N_166,N_241);
or U1178 (N_1178,N_242,In_1814);
nor U1179 (N_1179,N_393,In_1734);
and U1180 (N_1180,In_397,In_2119);
and U1181 (N_1181,In_1016,N_289);
and U1182 (N_1182,N_45,In_134);
or U1183 (N_1183,In_2034,In_205);
nand U1184 (N_1184,In_1689,In_1295);
and U1185 (N_1185,N_186,In_613);
nor U1186 (N_1186,In_1275,N_562);
xnor U1187 (N_1187,In_864,In_89);
nand U1188 (N_1188,In_296,In_2394);
nor U1189 (N_1189,N_536,In_2122);
nand U1190 (N_1190,In_1422,N_66);
or U1191 (N_1191,In_2132,In_1661);
xor U1192 (N_1192,In_2433,In_228);
nor U1193 (N_1193,In_1865,In_2104);
nor U1194 (N_1194,N_354,N_292);
or U1195 (N_1195,N_521,N_564);
or U1196 (N_1196,N_530,In_334);
and U1197 (N_1197,N_118,In_1558);
and U1198 (N_1198,In_1756,In_2296);
and U1199 (N_1199,In_1134,In_536);
nand U1200 (N_1200,In_361,In_1002);
nand U1201 (N_1201,N_341,In_27);
nor U1202 (N_1202,N_508,N_273);
and U1203 (N_1203,N_286,N_61);
or U1204 (N_1204,In_587,In_195);
and U1205 (N_1205,In_90,N_510);
and U1206 (N_1206,N_437,In_2057);
or U1207 (N_1207,In_1324,In_1418);
and U1208 (N_1208,In_1848,In_1995);
xnor U1209 (N_1209,N_534,N_460);
or U1210 (N_1210,In_1863,In_2036);
nand U1211 (N_1211,In_389,In_968);
or U1212 (N_1212,N_109,In_1899);
nand U1213 (N_1213,In_1109,In_269);
and U1214 (N_1214,In_248,N_303);
nor U1215 (N_1215,In_631,In_2465);
nand U1216 (N_1216,N_337,In_1699);
and U1217 (N_1217,N_332,In_2254);
or U1218 (N_1218,In_1597,In_927);
nand U1219 (N_1219,In_1682,In_1723);
or U1220 (N_1220,N_78,In_1084);
or U1221 (N_1221,N_194,In_2264);
and U1222 (N_1222,In_290,In_1717);
and U1223 (N_1223,In_1929,In_343);
or U1224 (N_1224,N_185,In_1620);
and U1225 (N_1225,N_616,In_667);
and U1226 (N_1226,In_1003,N_245);
nor U1227 (N_1227,In_988,In_577);
or U1228 (N_1228,N_272,N_350);
xor U1229 (N_1229,N_565,In_146);
nor U1230 (N_1230,N_108,In_1607);
and U1231 (N_1231,In_854,N_87);
nand U1232 (N_1232,In_517,In_435);
and U1233 (N_1233,In_1079,N_152);
nor U1234 (N_1234,In_1626,N_509);
nor U1235 (N_1235,N_524,In_437);
and U1236 (N_1236,In_688,In_1781);
or U1237 (N_1237,In_1004,N_240);
or U1238 (N_1238,In_2459,N_574);
nand U1239 (N_1239,In_185,In_951);
and U1240 (N_1240,In_96,In_377);
nor U1241 (N_1241,N_157,N_573);
and U1242 (N_1242,In_1211,In_63);
and U1243 (N_1243,N_47,In_533);
and U1244 (N_1244,In_380,In_1651);
or U1245 (N_1245,N_358,In_372);
nor U1246 (N_1246,N_529,In_1584);
nor U1247 (N_1247,N_206,N_60);
xnor U1248 (N_1248,N_90,N_298);
nand U1249 (N_1249,N_397,N_293);
nand U1250 (N_1250,In_2182,In_2084);
nand U1251 (N_1251,N_1176,N_497);
and U1252 (N_1252,N_644,In_2088);
xnor U1253 (N_1253,N_1118,N_1008);
and U1254 (N_1254,N_830,N_686);
xor U1255 (N_1255,N_652,N_86);
nand U1256 (N_1256,In_1666,N_1112);
nand U1257 (N_1257,N_1170,N_848);
or U1258 (N_1258,N_796,N_923);
nor U1259 (N_1259,N_429,In_749);
xor U1260 (N_1260,N_976,In_45);
nand U1261 (N_1261,In_1174,N_748);
or U1262 (N_1262,In_2423,N_891);
or U1263 (N_1263,N_525,N_864);
and U1264 (N_1264,N_1087,N_709);
nor U1265 (N_1265,In_105,In_1937);
xor U1266 (N_1266,N_1191,N_507);
or U1267 (N_1267,N_835,In_362);
nor U1268 (N_1268,In_1751,In_450);
nor U1269 (N_1269,In_1043,N_176);
nor U1270 (N_1270,N_648,N_1123);
or U1271 (N_1271,N_788,N_1110);
or U1272 (N_1272,N_177,N_977);
nor U1273 (N_1273,N_1230,N_1073);
nand U1274 (N_1274,In_2154,N_965);
nand U1275 (N_1275,N_968,N_205);
nand U1276 (N_1276,N_665,N_1014);
or U1277 (N_1277,In_2368,In_2070);
nand U1278 (N_1278,N_849,In_2322);
or U1279 (N_1279,In_112,N_789);
and U1280 (N_1280,In_547,N_1129);
nand U1281 (N_1281,In_807,N_1106);
nor U1282 (N_1282,N_925,N_1036);
xor U1283 (N_1283,N_1140,N_951);
nor U1284 (N_1284,In_2283,N_675);
and U1285 (N_1285,In_1137,N_1203);
nand U1286 (N_1286,N_441,N_790);
nand U1287 (N_1287,N_1150,N_916);
nand U1288 (N_1288,In_1433,N_1200);
or U1289 (N_1289,N_735,N_946);
or U1290 (N_1290,In_996,N_961);
nor U1291 (N_1291,N_907,N_1022);
nor U1292 (N_1292,In_912,N_594);
nand U1293 (N_1293,N_816,N_692);
nor U1294 (N_1294,N_948,N_71);
and U1295 (N_1295,N_750,N_1011);
nand U1296 (N_1296,In_834,In_1553);
nand U1297 (N_1297,In_373,N_679);
nor U1298 (N_1298,In_2016,In_203);
and U1299 (N_1299,N_260,N_621);
or U1300 (N_1300,In_232,In_1948);
and U1301 (N_1301,In_1879,In_579);
and U1302 (N_1302,N_658,In_1220);
or U1303 (N_1303,N_9,N_774);
nor U1304 (N_1304,In_1140,N_972);
xnor U1305 (N_1305,In_2028,In_1462);
nor U1306 (N_1306,N_1219,N_1031);
or U1307 (N_1307,N_1004,In_1579);
xnor U1308 (N_1308,In_2253,In_1412);
nand U1309 (N_1309,N_843,N_1032);
nand U1310 (N_1310,In_1034,N_1133);
xor U1311 (N_1311,N_782,N_540);
nand U1312 (N_1312,N_987,N_781);
and U1313 (N_1313,In_2224,N_1227);
and U1314 (N_1314,N_1098,N_489);
nor U1315 (N_1315,N_21,In_660);
nor U1316 (N_1316,In_736,In_1862);
and U1317 (N_1317,N_1030,N_88);
nand U1318 (N_1318,N_1119,N_184);
or U1319 (N_1319,N_65,N_983);
nor U1320 (N_1320,N_425,In_494);
nand U1321 (N_1321,N_756,In_1443);
nand U1322 (N_1322,N_982,N_807);
nand U1323 (N_1323,In_1919,N_1213);
or U1324 (N_1324,In_1249,N_1194);
nand U1325 (N_1325,In_2153,N_1162);
nor U1326 (N_1326,N_886,N_296);
or U1327 (N_1327,In_626,N_1006);
xor U1328 (N_1328,In_1444,N_969);
and U1329 (N_1329,In_251,N_1042);
nand U1330 (N_1330,N_978,N_745);
nor U1331 (N_1331,N_939,In_1033);
nand U1332 (N_1332,N_637,In_2221);
or U1333 (N_1333,In_152,In_606);
or U1334 (N_1334,In_2167,In_61);
and U1335 (N_1335,N_650,In_920);
and U1336 (N_1336,N_1063,N_1012);
nand U1337 (N_1337,N_897,N_1028);
and U1338 (N_1338,N_449,N_673);
and U1339 (N_1339,N_288,N_1010);
xor U1340 (N_1340,N_737,In_1914);
and U1341 (N_1341,In_2013,N_1013);
and U1342 (N_1342,N_903,N_918);
and U1343 (N_1343,N_19,In_1709);
or U1344 (N_1344,N_1206,N_91);
nor U1345 (N_1345,In_1676,In_15);
and U1346 (N_1346,In_2055,In_1890);
xnor U1347 (N_1347,N_822,N_598);
or U1348 (N_1348,N_874,In_153);
xnor U1349 (N_1349,N_804,N_1141);
nand U1350 (N_1350,In_1545,In_913);
nor U1351 (N_1351,In_2124,In_2491);
nand U1352 (N_1352,N_852,In_622);
nand U1353 (N_1353,N_1050,N_1156);
or U1354 (N_1354,N_173,N_964);
and U1355 (N_1355,N_765,In_1772);
and U1356 (N_1356,N_797,In_894);
nand U1357 (N_1357,In_2217,N_253);
xor U1358 (N_1358,In_1278,N_1000);
nor U1359 (N_1359,In_161,N_974);
and U1360 (N_1360,N_1053,N_674);
or U1361 (N_1361,N_779,N_423);
and U1362 (N_1362,N_254,N_1001);
nor U1363 (N_1363,In_1209,N_766);
nand U1364 (N_1364,N_643,N_1121);
or U1365 (N_1365,In_1577,N_626);
nand U1366 (N_1366,In_888,In_505);
xor U1367 (N_1367,N_1091,N_801);
xor U1368 (N_1368,N_1179,N_174);
nor U1369 (N_1369,N_1018,N_981);
nor U1370 (N_1370,In_2002,In_602);
nor U1371 (N_1371,N_1249,N_1215);
and U1372 (N_1372,N_738,N_1057);
nand U1373 (N_1373,N_1199,In_723);
and U1374 (N_1374,N_757,N_597);
and U1375 (N_1375,In_509,N_1064);
and U1376 (N_1376,N_1167,N_314);
or U1377 (N_1377,N_1033,N_924);
nand U1378 (N_1378,N_1082,N_1128);
nand U1379 (N_1379,N_821,In_387);
nand U1380 (N_1380,In_132,N_943);
nand U1381 (N_1381,N_182,In_898);
nand U1382 (N_1382,N_813,In_1969);
nand U1383 (N_1383,In_917,N_660);
or U1384 (N_1384,N_975,N_744);
or U1385 (N_1385,N_803,N_828);
and U1386 (N_1386,N_82,N_777);
or U1387 (N_1387,In_2473,In_817);
nand U1388 (N_1388,In_2432,N_1005);
nor U1389 (N_1389,In_1481,N_195);
or U1390 (N_1390,In_496,N_1122);
or U1391 (N_1391,N_629,In_2487);
xnor U1392 (N_1392,In_2311,In_2444);
nand U1393 (N_1393,N_1049,N_125);
nand U1394 (N_1394,N_986,In_774);
and U1395 (N_1395,N_603,In_1926);
or U1396 (N_1396,N_806,In_816);
nor U1397 (N_1397,N_1187,N_1038);
nor U1398 (N_1398,In_1200,N_1146);
nand U1399 (N_1399,N_970,N_1070);
nor U1400 (N_1400,N_929,In_1476);
nand U1401 (N_1401,N_129,In_1586);
nor U1402 (N_1402,In_1215,N_805);
and U1403 (N_1403,In_1949,N_63);
nor U1404 (N_1404,N_694,N_714);
or U1405 (N_1405,N_1069,N_880);
nand U1406 (N_1406,In_10,In_266);
or U1407 (N_1407,In_391,In_2067);
nand U1408 (N_1408,N_284,N_265);
or U1409 (N_1409,In_2128,In_1895);
xor U1410 (N_1410,In_1881,N_1061);
nand U1411 (N_1411,N_1231,N_1088);
and U1412 (N_1412,N_691,N_1158);
or U1413 (N_1413,N_940,N_1198);
nor U1414 (N_1414,In_1138,In_1228);
or U1415 (N_1415,N_237,In_159);
and U1416 (N_1416,In_1922,In_365);
nor U1417 (N_1417,N_1046,In_564);
or U1418 (N_1418,N_693,N_959);
or U1419 (N_1419,N_522,N_868);
and U1420 (N_1420,In_144,N_1034);
nor U1421 (N_1421,N_1025,N_1113);
nor U1422 (N_1422,N_387,N_1097);
nand U1423 (N_1423,N_257,In_1617);
nor U1424 (N_1424,N_659,N_1135);
or U1425 (N_1425,In_1388,In_1668);
or U1426 (N_1426,N_775,In_2015);
nand U1427 (N_1427,N_1177,N_795);
or U1428 (N_1428,N_759,N_250);
nor U1429 (N_1429,In_842,In_461);
and U1430 (N_1430,In_1489,In_1009);
and U1431 (N_1431,N_1145,In_2447);
nand U1432 (N_1432,In_630,In_275);
or U1433 (N_1433,N_492,N_764);
and U1434 (N_1434,N_1044,N_747);
nand U1435 (N_1435,N_754,In_1861);
nand U1436 (N_1436,In_84,N_863);
nand U1437 (N_1437,In_1464,N_1152);
nor U1438 (N_1438,N_535,In_1384);
and U1439 (N_1439,N_792,In_780);
nor U1440 (N_1440,N_388,N_950);
or U1441 (N_1441,N_703,In_34);
or U1442 (N_1442,In_2027,N_845);
nor U1443 (N_1443,In_2012,In_1285);
or U1444 (N_1444,N_1052,In_2395);
and U1445 (N_1445,In_436,In_1867);
and U1446 (N_1446,N_900,N_647);
nor U1447 (N_1447,N_1196,N_4);
and U1448 (N_1448,N_548,N_1148);
and U1449 (N_1449,N_784,N_651);
and U1450 (N_1450,N_252,N_945);
or U1451 (N_1451,N_155,In_1163);
and U1452 (N_1452,In_882,N_380);
nand U1453 (N_1453,N_898,N_1131);
nor U1454 (N_1454,In_1847,N_815);
nand U1455 (N_1455,N_875,In_220);
nor U1456 (N_1456,N_198,N_904);
or U1457 (N_1457,N_1139,In_1182);
and U1458 (N_1458,N_938,In_922);
nand U1459 (N_1459,In_2074,N_1101);
or U1460 (N_1460,N_726,In_419);
and U1461 (N_1461,N_1060,N_824);
nand U1462 (N_1462,In_878,N_484);
nand U1463 (N_1463,In_238,N_847);
nand U1464 (N_1464,N_895,N_153);
xor U1465 (N_1465,N_246,N_1095);
nor U1466 (N_1466,In_1419,N_378);
and U1467 (N_1467,N_662,In_1391);
nand U1468 (N_1468,N_1107,N_696);
xnor U1469 (N_1469,In_1538,N_1175);
and U1470 (N_1470,N_41,N_808);
nor U1471 (N_1471,N_915,In_2485);
nor U1472 (N_1472,N_721,In_2044);
nand U1473 (N_1473,N_1084,N_190);
nand U1474 (N_1474,In_2389,In_293);
and U1475 (N_1475,N_700,In_2229);
or U1476 (N_1476,In_116,N_628);
nand U1477 (N_1477,N_199,N_306);
or U1478 (N_1478,N_121,N_1149);
nor U1479 (N_1479,N_736,In_2438);
nor U1480 (N_1480,N_743,N_682);
and U1481 (N_1481,N_878,N_711);
or U1482 (N_1482,N_379,N_753);
and U1483 (N_1483,N_676,N_941);
nor U1484 (N_1484,N_133,N_462);
and U1485 (N_1485,N_1160,N_812);
or U1486 (N_1486,N_614,In_1768);
or U1487 (N_1487,In_1595,N_1037);
nand U1488 (N_1488,N_706,N_689);
nand U1489 (N_1489,N_671,N_34);
xnor U1490 (N_1490,In_2249,N_862);
and U1491 (N_1491,N_910,In_1657);
or U1492 (N_1492,N_1093,N_1075);
and U1493 (N_1493,N_68,N_1078);
xnor U1494 (N_1494,N_92,N_1043);
or U1495 (N_1495,N_612,In_98);
or U1496 (N_1496,In_732,N_739);
or U1497 (N_1497,In_2157,N_1157);
nor U1498 (N_1498,N_718,N_749);
nand U1499 (N_1499,N_1002,In_206);
nor U1500 (N_1500,N_809,N_110);
or U1501 (N_1501,In_424,N_613);
nor U1502 (N_1502,N_927,N_725);
nor U1503 (N_1503,In_1560,In_1810);
nand U1504 (N_1504,N_365,In_12);
nand U1505 (N_1505,In_1821,N_147);
and U1506 (N_1506,N_697,N_140);
and U1507 (N_1507,N_193,N_984);
nand U1508 (N_1508,In_1667,N_209);
nor U1509 (N_1509,N_839,N_892);
nand U1510 (N_1510,In_1569,N_95);
or U1511 (N_1511,In_540,N_85);
nand U1512 (N_1512,N_1124,N_872);
and U1513 (N_1513,In_886,N_820);
or U1514 (N_1514,N_1016,N_1237);
nor U1515 (N_1515,N_622,N_1243);
nand U1516 (N_1516,N_957,In_1963);
nor U1517 (N_1517,N_730,N_741);
and U1518 (N_1518,N_687,N_640);
or U1519 (N_1519,N_156,N_1247);
nand U1520 (N_1520,N_1181,N_1109);
nor U1521 (N_1521,N_1099,N_442);
and U1522 (N_1522,N_132,In_790);
nand U1523 (N_1523,N_630,N_77);
or U1524 (N_1524,In_2196,In_1120);
or U1525 (N_1525,N_826,N_873);
xnor U1526 (N_1526,In_177,N_503);
nor U1527 (N_1527,In_462,N_1027);
or U1528 (N_1528,N_1083,N_239);
and U1529 (N_1529,N_1071,N_1065);
xnor U1530 (N_1530,N_728,N_17);
and U1531 (N_1531,N_38,N_1143);
nand U1532 (N_1532,N_434,N_1234);
and U1533 (N_1533,N_908,In_779);
or U1534 (N_1534,N_1026,N_1081);
nand U1535 (N_1535,N_1190,In_173);
and U1536 (N_1536,N_729,In_2290);
and U1537 (N_1537,N_567,N_901);
or U1538 (N_1538,In_684,In_872);
or U1539 (N_1539,N_771,N_625);
nand U1540 (N_1540,N_960,N_1173);
or U1541 (N_1541,N_624,N_802);
nand U1542 (N_1542,N_856,In_1092);
nor U1543 (N_1543,N_786,N_654);
xnor U1544 (N_1544,N_1212,N_553);
or U1545 (N_1545,N_73,In_1716);
and U1546 (N_1546,N_695,N_791);
or U1547 (N_1547,N_278,N_935);
xor U1548 (N_1548,N_1021,In_2347);
and U1549 (N_1549,N_858,In_2323);
or U1550 (N_1550,N_732,N_634);
or U1551 (N_1551,N_866,N_893);
nor U1552 (N_1552,In_11,In_752);
and U1553 (N_1553,In_327,In_994);
and U1554 (N_1554,In_933,N_1127);
xor U1555 (N_1555,In_1675,In_530);
xnor U1556 (N_1556,N_486,In_2050);
or U1557 (N_1557,N_1189,In_753);
xnor U1558 (N_1558,In_1199,N_890);
xor U1559 (N_1559,N_837,N_932);
nand U1560 (N_1560,N_107,N_1184);
and U1561 (N_1561,N_1240,In_412);
and U1562 (N_1562,In_135,N_955);
and U1563 (N_1563,N_611,In_2150);
nand U1564 (N_1564,N_323,N_881);
or U1565 (N_1565,N_1180,N_104);
and U1566 (N_1566,N_1172,N_762);
nand U1567 (N_1567,N_1138,N_461);
nand U1568 (N_1568,In_1169,N_1074);
nor U1569 (N_1569,In_2451,N_119);
and U1570 (N_1570,In_1181,N_990);
nor U1571 (N_1571,N_888,N_670);
or U1572 (N_1572,In_2103,In_2090);
nor U1573 (N_1573,N_1244,N_532);
and U1574 (N_1574,N_15,In_2400);
xor U1575 (N_1575,N_471,In_2041);
nand U1576 (N_1576,N_1017,N_1066);
nand U1577 (N_1577,In_1830,N_834);
nor U1578 (N_1578,N_719,N_1114);
or U1579 (N_1579,In_1445,In_1087);
nor U1580 (N_1580,N_707,N_720);
nand U1581 (N_1581,In_60,In_2230);
xor U1582 (N_1582,N_926,N_347);
and U1583 (N_1583,In_1652,N_600);
nand U1584 (N_1584,In_470,N_1193);
nand U1585 (N_1585,In_2180,N_967);
nand U1586 (N_1586,N_1130,In_150);
or U1587 (N_1587,N_661,N_740);
and U1588 (N_1588,N_850,N_794);
and U1589 (N_1589,N_72,N_180);
xor U1590 (N_1590,In_1690,N_917);
xnor U1591 (N_1591,N_1168,In_2247);
nand U1592 (N_1592,In_92,N_684);
nor U1593 (N_1593,In_2020,N_798);
nor U1594 (N_1594,N_111,In_855);
xor U1595 (N_1595,N_1229,N_1155);
and U1596 (N_1596,N_642,N_713);
or U1597 (N_1597,In_1371,N_827);
and U1598 (N_1598,N_454,In_1817);
and U1599 (N_1599,In_625,N_496);
nand U1600 (N_1600,In_74,N_1216);
nor U1601 (N_1601,N_290,N_1154);
nand U1602 (N_1602,N_962,In_905);
nor U1603 (N_1603,N_127,N_270);
xnor U1604 (N_1604,N_1226,N_912);
xor U1605 (N_1605,In_2069,In_1420);
or U1606 (N_1606,In_671,N_742);
nor U1607 (N_1607,N_1192,In_1502);
nor U1608 (N_1608,N_663,In_163);
and U1609 (N_1609,N_933,In_2472);
nor U1610 (N_1610,N_723,N_1218);
and U1611 (N_1611,N_780,In_1325);
or U1612 (N_1612,N_1076,In_740);
nor U1613 (N_1613,N_1210,N_1105);
and U1614 (N_1614,In_1314,N_979);
xnor U1615 (N_1615,In_1290,In_2225);
nand U1616 (N_1616,N_701,In_638);
nor U1617 (N_1617,N_1178,In_646);
and U1618 (N_1618,In_1019,N_783);
and U1619 (N_1619,In_2442,N_752);
nand U1620 (N_1620,N_677,N_1116);
or U1621 (N_1621,N_840,N_1103);
nand U1622 (N_1622,N_905,N_463);
nor U1623 (N_1623,N_708,N_793);
xnor U1624 (N_1624,N_767,In_1477);
or U1625 (N_1625,In_1265,N_1164);
and U1626 (N_1626,N_1171,N_377);
nand U1627 (N_1627,N_678,N_226);
nand U1628 (N_1628,N_857,N_778);
nor U1629 (N_1629,N_1051,N_819);
and U1630 (N_1630,N_319,N_877);
nor U1631 (N_1631,N_322,N_853);
and U1632 (N_1632,N_772,In_154);
or U1633 (N_1633,N_667,N_632);
xor U1634 (N_1634,In_860,In_2281);
or U1635 (N_1635,In_2089,N_1239);
nand U1636 (N_1636,In_711,In_1030);
xor U1637 (N_1637,N_763,N_1019);
or U1638 (N_1638,N_851,N_865);
nand U1639 (N_1639,In_1115,N_704);
or U1640 (N_1640,N_1015,N_134);
or U1641 (N_1641,N_768,N_172);
or U1642 (N_1642,In_209,N_546);
or U1643 (N_1643,N_398,N_914);
or U1644 (N_1644,N_128,N_417);
nand U1645 (N_1645,In_798,N_733);
nand U1646 (N_1646,N_549,N_1086);
and U1647 (N_1647,N_1104,N_773);
nand U1648 (N_1648,N_526,In_1744);
or U1649 (N_1649,N_1223,N_998);
and U1650 (N_1650,In_544,N_645);
or U1651 (N_1651,In_1874,N_235);
nand U1652 (N_1652,N_1023,N_885);
nor U1653 (N_1653,In_2401,N_902);
nor U1654 (N_1654,N_702,N_1085);
and U1655 (N_1655,In_1256,In_1253);
and U1656 (N_1656,In_1222,N_666);
xor U1657 (N_1657,N_1147,N_995);
or U1658 (N_1658,N_867,In_2396);
xnor U1659 (N_1659,N_1111,N_712);
nand U1660 (N_1660,N_921,N_1054);
nor U1661 (N_1661,N_243,N_1222);
nand U1662 (N_1662,N_24,In_1944);
nor U1663 (N_1663,In_403,N_993);
nor U1664 (N_1664,N_444,N_609);
nor U1665 (N_1665,In_1608,N_949);
nand U1666 (N_1666,N_1142,N_14);
or U1667 (N_1667,N_1056,In_518);
or U1668 (N_1668,N_1079,N_930);
or U1669 (N_1669,N_937,N_879);
nor U1670 (N_1670,In_1051,N_683);
and U1671 (N_1671,N_1092,N_722);
nand U1672 (N_1672,N_232,N_944);
nand U1673 (N_1673,N_203,In_1780);
xor U1674 (N_1674,N_409,In_1856);
and U1675 (N_1675,In_1219,N_280);
xnor U1676 (N_1676,In_1468,N_1039);
or U1677 (N_1677,In_2397,N_823);
nor U1678 (N_1678,N_672,N_255);
and U1679 (N_1679,In_457,N_1188);
nor U1680 (N_1680,In_867,N_1166);
nand U1681 (N_1681,N_992,N_1115);
nand U1682 (N_1682,In_1405,N_922);
nand U1683 (N_1683,In_1085,In_1319);
and U1684 (N_1684,N_668,N_1100);
and U1685 (N_1685,N_635,N_1089);
nand U1686 (N_1686,In_2051,N_1144);
nand U1687 (N_1687,N_1125,In_137);
or U1688 (N_1688,In_1761,In_2471);
and U1689 (N_1689,N_1245,N_988);
or U1690 (N_1690,In_175,N_989);
nor U1691 (N_1691,In_1986,In_320);
or U1692 (N_1692,N_636,In_2282);
or U1693 (N_1693,N_1221,N_469);
and U1694 (N_1694,In_828,N_1047);
nand U1695 (N_1695,N_760,N_321);
or U1696 (N_1696,In_2003,N_731);
nand U1697 (N_1697,In_1241,N_1214);
nand U1698 (N_1698,N_958,N_554);
nand U1699 (N_1699,N_285,N_639);
or U1700 (N_1700,In_441,In_2325);
nand U1701 (N_1701,N_920,N_973);
and U1702 (N_1702,N_211,N_896);
nand U1703 (N_1703,N_159,In_2477);
nor U1704 (N_1704,N_664,N_889);
nor U1705 (N_1705,N_493,N_724);
xor U1706 (N_1706,N_35,In_929);
xnor U1707 (N_1707,N_1165,N_942);
or U1708 (N_1708,In_903,N_376);
xor U1709 (N_1709,N_373,In_1866);
or U1710 (N_1710,N_952,N_810);
and U1711 (N_1711,In_1183,In_481);
or U1712 (N_1712,N_53,N_1048);
and U1713 (N_1713,N_909,In_1854);
nor U1714 (N_1714,N_832,N_1183);
and U1715 (N_1715,In_1244,In_2205);
nor U1716 (N_1716,In_1531,In_1357);
and U1717 (N_1717,In_1486,N_5);
and U1718 (N_1718,N_1153,In_670);
and U1719 (N_1719,N_685,In_2269);
nand U1720 (N_1720,In_65,N_871);
nand U1721 (N_1721,N_412,N_1169);
or U1722 (N_1722,N_1062,N_716);
or U1723 (N_1723,In_961,N_919);
nand U1724 (N_1724,N_244,N_1207);
nor U1725 (N_1725,N_838,In_938);
nand U1726 (N_1726,N_681,N_825);
and U1727 (N_1727,N_221,N_894);
nand U1728 (N_1728,N_591,N_415);
and U1729 (N_1729,N_1136,N_313);
and U1730 (N_1730,N_906,In_2171);
or U1731 (N_1731,N_928,In_1664);
nor U1732 (N_1732,In_1860,N_842);
and U1733 (N_1733,In_1767,N_421);
nor U1734 (N_1734,N_1238,In_607);
nor U1735 (N_1735,In_588,N_831);
nand U1736 (N_1736,In_1605,N_577);
nor U1737 (N_1737,N_1009,In_2114);
and U1738 (N_1738,In_2419,N_997);
nand U1739 (N_1739,N_855,N_99);
and U1740 (N_1740,In_1903,N_213);
or U1741 (N_1741,N_1224,In_1161);
and U1742 (N_1742,N_569,In_2177);
or U1743 (N_1743,In_1798,In_997);
and U1744 (N_1744,N_59,N_836);
nand U1745 (N_1745,N_698,N_1217);
nor U1746 (N_1746,In_2215,N_249);
nand U1747 (N_1747,N_631,N_191);
nand U1748 (N_1748,N_746,N_1035);
and U1749 (N_1749,N_1055,In_629);
xnor U1750 (N_1750,N_655,N_1232);
and U1751 (N_1751,N_899,N_861);
or U1752 (N_1752,N_758,In_1307);
or U1753 (N_1753,N_1117,In_2239);
nand U1754 (N_1754,In_1787,In_2256);
or U1755 (N_1755,In_186,N_1067);
xnor U1756 (N_1756,N_1096,In_537);
or U1757 (N_1757,In_202,In_70);
and U1758 (N_1758,N_431,In_82);
and U1759 (N_1759,N_102,N_576);
or U1760 (N_1760,In_1150,N_1233);
and U1761 (N_1761,In_1632,N_947);
nor U1762 (N_1762,N_1132,In_813);
nand U1763 (N_1763,In_176,In_1719);
or U1764 (N_1764,N_883,N_410);
or U1765 (N_1765,N_999,In_1280);
nand U1766 (N_1766,N_1228,N_1108);
and U1767 (N_1767,In_2174,N_445);
or U1768 (N_1768,N_638,In_1049);
nor U1769 (N_1769,N_994,N_680);
or U1770 (N_1770,In_1344,N_175);
nor U1771 (N_1771,N_1241,N_1058);
or U1772 (N_1772,In_668,N_164);
nor U1773 (N_1773,In_1310,N_1197);
nand U1774 (N_1774,N_1201,In_608);
nand U1775 (N_1775,N_1040,N_641);
or U1776 (N_1776,N_438,N_936);
nand U1777 (N_1777,In_224,In_524);
and U1778 (N_1778,N_715,N_1045);
nor U1779 (N_1779,N_690,In_871);
or U1780 (N_1780,N_1220,N_841);
or U1781 (N_1781,In_1746,N_699);
and U1782 (N_1782,N_392,In_1397);
nand U1783 (N_1783,N_1102,N_800);
nor U1784 (N_1784,N_1090,N_887);
nor U1785 (N_1785,N_1080,In_1485);
and U1786 (N_1786,In_2024,In_250);
or U1787 (N_1787,N_818,N_956);
nand U1788 (N_1788,N_653,In_1670);
xor U1789 (N_1789,In_877,N_1003);
xnor U1790 (N_1790,N_869,In_1696);
nand U1791 (N_1791,N_13,N_734);
and U1792 (N_1792,N_236,N_751);
and U1793 (N_1793,N_1225,In_1529);
or U1794 (N_1794,In_1571,N_168);
nor U1795 (N_1795,N_1077,In_822);
xor U1796 (N_1796,In_694,N_1248);
nor U1797 (N_1797,In_1519,N_1029);
or U1798 (N_1798,N_1020,N_371);
and U1799 (N_1799,N_28,N_846);
and U1800 (N_1800,N_385,N_799);
nor U1801 (N_1801,N_1068,N_954);
and U1802 (N_1802,N_980,N_1134);
nor U1803 (N_1803,N_1137,In_2435);
nor U1804 (N_1804,N_776,N_911);
nor U1805 (N_1805,In_859,In_117);
or U1806 (N_1806,N_710,In_1373);
or U1807 (N_1807,N_113,In_491);
xnor U1808 (N_1808,N_934,N_233);
nand U1809 (N_1809,N_143,N_717);
or U1810 (N_1810,In_677,N_1208);
or U1811 (N_1811,In_2261,In_2489);
or U1812 (N_1812,N_76,N_1007);
nand U1813 (N_1813,N_1235,In_1390);
and U1814 (N_1814,N_1195,N_602);
and U1815 (N_1815,N_884,In_1367);
and U1816 (N_1816,N_302,N_913);
xnor U1817 (N_1817,In_2345,In_1234);
or U1818 (N_1818,In_2118,N_528);
xnor U1819 (N_1819,In_1977,N_727);
nand U1820 (N_1820,In_686,N_646);
nor U1821 (N_1821,N_649,In_833);
nor U1822 (N_1822,In_1968,N_963);
or U1823 (N_1823,N_188,In_1857);
and U1824 (N_1824,In_1152,N_1202);
nand U1825 (N_1825,N_1041,In_201);
nand U1826 (N_1826,N_1246,N_502);
or U1827 (N_1827,N_859,N_931);
nor U1828 (N_1828,N_814,N_787);
or U1829 (N_1829,N_876,In_841);
nor U1830 (N_1830,N_844,N_882);
and U1831 (N_1831,N_325,N_657);
or U1832 (N_1832,N_705,N_1163);
and U1833 (N_1833,In_858,In_1864);
nand U1834 (N_1834,In_1345,N_283);
or U1835 (N_1835,N_854,N_669);
or U1836 (N_1836,N_769,N_1186);
nand U1837 (N_1837,N_1094,N_1185);
and U1838 (N_1838,N_1126,N_1059);
nand U1839 (N_1839,In_400,N_656);
nand U1840 (N_1840,In_2211,N_870);
nand U1841 (N_1841,N_1236,N_860);
and U1842 (N_1842,N_1120,In_846);
nand U1843 (N_1843,N_627,In_1960);
nor U1844 (N_1844,In_1592,N_465);
nor U1845 (N_1845,N_817,In_2392);
or U1846 (N_1846,N_427,N_473);
nand U1847 (N_1847,In_254,N_966);
nor U1848 (N_1848,N_424,N_1242);
or U1849 (N_1849,In_1703,In_1940);
nand U1850 (N_1850,N_1151,In_2277);
and U1851 (N_1851,In_379,N_585);
nor U1852 (N_1852,N_266,In_239);
nor U1853 (N_1853,N_1182,N_770);
and U1854 (N_1854,N_833,N_1211);
xor U1855 (N_1855,In_2370,In_598);
and U1856 (N_1856,N_688,N_1159);
nor U1857 (N_1857,N_953,In_1393);
and U1858 (N_1858,N_1204,N_1209);
xor U1859 (N_1859,N_523,N_1174);
and U1860 (N_1860,N_829,N_1072);
and U1861 (N_1861,In_2022,N_971);
or U1862 (N_1862,N_514,In_1762);
and U1863 (N_1863,In_1953,In_2259);
nor U1864 (N_1864,N_1161,In_1925);
or U1865 (N_1865,N_985,In_2009);
nor U1866 (N_1866,N_55,In_1712);
nand U1867 (N_1867,In_960,N_785);
or U1868 (N_1868,N_1205,In_451);
nor U1869 (N_1869,N_996,In_1197);
nor U1870 (N_1870,N_30,N_991);
nand U1871 (N_1871,N_633,N_761);
nand U1872 (N_1872,In_51,N_755);
or U1873 (N_1873,N_811,N_154);
and U1874 (N_1874,In_617,N_1024);
or U1875 (N_1875,N_1329,N_1832);
nand U1876 (N_1876,N_1661,N_1567);
nand U1877 (N_1877,N_1628,N_1330);
and U1878 (N_1878,N_1496,N_1605);
nand U1879 (N_1879,N_1295,N_1586);
nor U1880 (N_1880,N_1429,N_1819);
and U1881 (N_1881,N_1717,N_1400);
and U1882 (N_1882,N_1509,N_1257);
and U1883 (N_1883,N_1572,N_1476);
nand U1884 (N_1884,N_1292,N_1564);
or U1885 (N_1885,N_1613,N_1415);
nand U1886 (N_1886,N_1540,N_1660);
nand U1887 (N_1887,N_1784,N_1419);
or U1888 (N_1888,N_1839,N_1270);
and U1889 (N_1889,N_1574,N_1376);
nand U1890 (N_1890,N_1386,N_1517);
or U1891 (N_1891,N_1640,N_1260);
nor U1892 (N_1892,N_1851,N_1473);
nand U1893 (N_1893,N_1579,N_1286);
and U1894 (N_1894,N_1543,N_1332);
and U1895 (N_1895,N_1825,N_1744);
or U1896 (N_1896,N_1826,N_1841);
nor U1897 (N_1897,N_1563,N_1384);
nand U1898 (N_1898,N_1364,N_1766);
nor U1899 (N_1899,N_1665,N_1449);
and U1900 (N_1900,N_1636,N_1498);
nor U1901 (N_1901,N_1763,N_1702);
nor U1902 (N_1902,N_1710,N_1278);
nor U1903 (N_1903,N_1647,N_1505);
nor U1904 (N_1904,N_1488,N_1420);
and U1905 (N_1905,N_1569,N_1444);
nor U1906 (N_1906,N_1456,N_1823);
nor U1907 (N_1907,N_1314,N_1606);
xnor U1908 (N_1908,N_1787,N_1409);
or U1909 (N_1909,N_1709,N_1447);
nand U1910 (N_1910,N_1525,N_1530);
or U1911 (N_1911,N_1304,N_1264);
and U1912 (N_1912,N_1822,N_1351);
nor U1913 (N_1913,N_1455,N_1287);
xnor U1914 (N_1914,N_1458,N_1688);
xnor U1915 (N_1915,N_1408,N_1664);
nor U1916 (N_1916,N_1635,N_1382);
nand U1917 (N_1917,N_1707,N_1849);
or U1918 (N_1918,N_1526,N_1536);
nor U1919 (N_1919,N_1815,N_1418);
or U1920 (N_1920,N_1343,N_1575);
nor U1921 (N_1921,N_1305,N_1381);
nand U1922 (N_1922,N_1266,N_1703);
nand U1923 (N_1923,N_1844,N_1322);
or U1924 (N_1924,N_1294,N_1803);
xor U1925 (N_1925,N_1261,N_1311);
nand U1926 (N_1926,N_1410,N_1735);
or U1927 (N_1927,N_1651,N_1805);
and U1928 (N_1928,N_1578,N_1860);
or U1929 (N_1929,N_1518,N_1609);
or U1930 (N_1930,N_1359,N_1788);
and U1931 (N_1931,N_1775,N_1315);
or U1932 (N_1932,N_1389,N_1439);
nand U1933 (N_1933,N_1462,N_1486);
or U1934 (N_1934,N_1399,N_1682);
xor U1935 (N_1935,N_1782,N_1556);
nand U1936 (N_1936,N_1341,N_1277);
nand U1937 (N_1937,N_1659,N_1417);
and U1938 (N_1938,N_1431,N_1691);
nand U1939 (N_1939,N_1291,N_1445);
or U1940 (N_1940,N_1837,N_1804);
nand U1941 (N_1941,N_1274,N_1650);
nand U1942 (N_1942,N_1437,N_1610);
nand U1943 (N_1943,N_1630,N_1396);
nand U1944 (N_1944,N_1489,N_1423);
nand U1945 (N_1945,N_1273,N_1771);
nor U1946 (N_1946,N_1412,N_1519);
and U1947 (N_1947,N_1406,N_1342);
nor U1948 (N_1948,N_1318,N_1807);
nor U1949 (N_1949,N_1678,N_1577);
or U1950 (N_1950,N_1495,N_1490);
or U1951 (N_1951,N_1279,N_1477);
nor U1952 (N_1952,N_1474,N_1840);
and U1953 (N_1953,N_1300,N_1809);
and U1954 (N_1954,N_1531,N_1510);
or U1955 (N_1955,N_1331,N_1634);
or U1956 (N_1956,N_1743,N_1559);
or U1957 (N_1957,N_1549,N_1850);
nor U1958 (N_1958,N_1629,N_1836);
nor U1959 (N_1959,N_1697,N_1546);
nor U1960 (N_1960,N_1785,N_1648);
or U1961 (N_1961,N_1720,N_1798);
nor U1962 (N_1962,N_1690,N_1778);
and U1963 (N_1963,N_1435,N_1786);
nand U1964 (N_1964,N_1633,N_1667);
or U1965 (N_1965,N_1334,N_1719);
nand U1966 (N_1966,N_1324,N_1463);
nor U1967 (N_1967,N_1770,N_1598);
and U1968 (N_1968,N_1482,N_1340);
and U1969 (N_1969,N_1362,N_1537);
or U1970 (N_1970,N_1643,N_1862);
or U1971 (N_1971,N_1453,N_1742);
xor U1972 (N_1972,N_1426,N_1459);
nand U1973 (N_1973,N_1584,N_1676);
xor U1974 (N_1974,N_1612,N_1621);
nor U1975 (N_1975,N_1773,N_1675);
nor U1976 (N_1976,N_1457,N_1639);
nand U1977 (N_1977,N_1325,N_1872);
nand U1978 (N_1978,N_1297,N_1668);
or U1979 (N_1979,N_1632,N_1452);
and U1980 (N_1980,N_1704,N_1712);
nand U1981 (N_1981,N_1827,N_1859);
or U1982 (N_1982,N_1600,N_1440);
xor U1983 (N_1983,N_1679,N_1741);
nand U1984 (N_1984,N_1383,N_1821);
or U1985 (N_1985,N_1796,N_1669);
and U1986 (N_1986,N_1581,N_1701);
xor U1987 (N_1987,N_1358,N_1696);
nor U1988 (N_1988,N_1620,N_1718);
nand U1989 (N_1989,N_1312,N_1566);
nor U1990 (N_1990,N_1595,N_1276);
nor U1991 (N_1991,N_1398,N_1316);
or U1992 (N_1992,N_1756,N_1721);
xor U1993 (N_1993,N_1655,N_1461);
and U1994 (N_1994,N_1855,N_1250);
nand U1995 (N_1995,N_1403,N_1732);
and U1996 (N_1996,N_1754,N_1861);
or U1997 (N_1997,N_1551,N_1834);
nor U1998 (N_1998,N_1319,N_1421);
xor U1999 (N_1999,N_1739,N_1251);
and U2000 (N_2000,N_1523,N_1533);
nor U2001 (N_2001,N_1871,N_1432);
and U2002 (N_2002,N_1768,N_1497);
and U2003 (N_2003,N_1538,N_1751);
nor U2004 (N_2004,N_1357,N_1857);
nand U2005 (N_2005,N_1781,N_1764);
nand U2006 (N_2006,N_1783,N_1683);
or U2007 (N_2007,N_1730,N_1414);
or U2008 (N_2008,N_1475,N_1622);
nor U2009 (N_2009,N_1740,N_1570);
nor U2010 (N_2010,N_1649,N_1654);
nor U2011 (N_2011,N_1366,N_1373);
xnor U2012 (N_2012,N_1797,N_1603);
and U2013 (N_2013,N_1824,N_1573);
nand U2014 (N_2014,N_1402,N_1761);
or U2015 (N_2015,N_1722,N_1363);
nor U2016 (N_2016,N_1694,N_1561);
and U2017 (N_2017,N_1293,N_1354);
nand U2018 (N_2018,N_1309,N_1731);
and U2019 (N_2019,N_1854,N_1657);
nand U2020 (N_2020,N_1438,N_1555);
nand U2021 (N_2021,N_1392,N_1835);
or U2022 (N_2022,N_1360,N_1856);
and U2023 (N_2023,N_1728,N_1820);
nor U2024 (N_2024,N_1700,N_1539);
nor U2025 (N_2025,N_1853,N_1256);
and U2026 (N_2026,N_1597,N_1638);
and U2027 (N_2027,N_1689,N_1789);
xor U2028 (N_2028,N_1795,N_1337);
or U2029 (N_2029,N_1548,N_1843);
nand U2030 (N_2030,N_1831,N_1338);
nor U2031 (N_2031,N_1607,N_1800);
and U2032 (N_2032,N_1507,N_1368);
nor U2033 (N_2033,N_1663,N_1395);
nand U2034 (N_2034,N_1298,N_1838);
nand U2035 (N_2035,N_1448,N_1441);
or U2036 (N_2036,N_1867,N_1816);
nor U2037 (N_2037,N_1799,N_1616);
or U2038 (N_2038,N_1749,N_1361);
nor U2039 (N_2039,N_1535,N_1503);
and U2040 (N_2040,N_1289,N_1253);
nand U2041 (N_2041,N_1356,N_1868);
or U2042 (N_2042,N_1374,N_1755);
and U2043 (N_2043,N_1752,N_1684);
or U2044 (N_2044,N_1594,N_1550);
nor U2045 (N_2045,N_1302,N_1480);
or U2046 (N_2046,N_1487,N_1738);
nand U2047 (N_2047,N_1865,N_1275);
nor U2048 (N_2048,N_1671,N_1848);
xnor U2049 (N_2049,N_1485,N_1387);
nand U2050 (N_2050,N_1470,N_1460);
nand U2051 (N_2051,N_1587,N_1748);
or U2052 (N_2052,N_1355,N_1336);
xnor U2053 (N_2053,N_1686,N_1802);
and U2054 (N_2054,N_1308,N_1451);
and U2055 (N_2055,N_1745,N_1858);
and U2056 (N_2056,N_1626,N_1642);
nor U2057 (N_2057,N_1511,N_1829);
and U2058 (N_2058,N_1442,N_1349);
nor U2059 (N_2059,N_1615,N_1759);
nand U2060 (N_2060,N_1469,N_1500);
nor U2061 (N_2061,N_1765,N_1596);
or U2062 (N_2062,N_1762,N_1812);
nor U2063 (N_2063,N_1619,N_1388);
and U2064 (N_2064,N_1321,N_1725);
nor U2065 (N_2065,N_1284,N_1472);
and U2066 (N_2066,N_1624,N_1604);
nand U2067 (N_2067,N_1541,N_1464);
or U2068 (N_2068,N_1767,N_1681);
nand U2069 (N_2069,N_1758,N_1637);
nor U2070 (N_2070,N_1576,N_1733);
xnor U2071 (N_2071,N_1588,N_1307);
nor U2072 (N_2072,N_1506,N_1347);
or U2073 (N_2073,N_1553,N_1601);
nand U2074 (N_2074,N_1269,N_1492);
nand U2075 (N_2075,N_1267,N_1792);
nand U2076 (N_2076,N_1545,N_1723);
and U2077 (N_2077,N_1692,N_1562);
nor U2078 (N_2078,N_1411,N_1680);
nand U2079 (N_2079,N_1580,N_1375);
nand U2080 (N_2080,N_1698,N_1673);
xor U2081 (N_2081,N_1774,N_1780);
and U2082 (N_2082,N_1801,N_1625);
nor U2083 (N_2083,N_1672,N_1339);
nand U2084 (N_2084,N_1810,N_1263);
or U2085 (N_2085,N_1811,N_1571);
nand U2086 (N_2086,N_1407,N_1641);
nor U2087 (N_2087,N_1662,N_1466);
xnor U2088 (N_2088,N_1422,N_1290);
nand U2089 (N_2089,N_1515,N_1369);
nand U2090 (N_2090,N_1873,N_1280);
and U2091 (N_2091,N_1446,N_1591);
nor U2092 (N_2092,N_1258,N_1527);
and U2093 (N_2093,N_1847,N_1736);
nand U2094 (N_2094,N_1599,N_1554);
or U2095 (N_2095,N_1413,N_1467);
xor U2096 (N_2096,N_1471,N_1808);
or U2097 (N_2097,N_1777,N_1714);
or U2098 (N_2098,N_1393,N_1352);
or U2099 (N_2099,N_1716,N_1254);
xor U2100 (N_2100,N_1544,N_1753);
and U2101 (N_2101,N_1769,N_1268);
nor U2102 (N_2102,N_1345,N_1560);
or U2103 (N_2103,N_1346,N_1602);
and U2104 (N_2104,N_1528,N_1468);
and U2105 (N_2105,N_1685,N_1552);
or U2106 (N_2106,N_1394,N_1425);
xnor U2107 (N_2107,N_1711,N_1813);
or U2108 (N_2108,N_1372,N_1379);
and U2109 (N_2109,N_1617,N_1757);
xor U2110 (N_2110,N_1869,N_1864);
nand U2111 (N_2111,N_1259,N_1385);
nand U2112 (N_2112,N_1760,N_1494);
nor U2113 (N_2113,N_1430,N_1695);
or U2114 (N_2114,N_1532,N_1501);
and U2115 (N_2115,N_1481,N_1303);
nor U2116 (N_2116,N_1283,N_1713);
xor U2117 (N_2117,N_1465,N_1817);
or U2118 (N_2118,N_1493,N_1288);
nand U2119 (N_2119,N_1252,N_1852);
and U2120 (N_2120,N_1729,N_1370);
or U2121 (N_2121,N_1265,N_1565);
nand U2122 (N_2122,N_1608,N_1520);
or U2123 (N_2123,N_1585,N_1734);
or U2124 (N_2124,N_1793,N_1365);
nand U2125 (N_2125,N_1776,N_1479);
xor U2126 (N_2126,N_1542,N_1644);
or U2127 (N_2127,N_1627,N_1317);
nor U2128 (N_2128,N_1313,N_1310);
or U2129 (N_2129,N_1296,N_1326);
nand U2130 (N_2130,N_1618,N_1658);
nor U2131 (N_2131,N_1397,N_1547);
nand U2132 (N_2132,N_1301,N_1750);
nor U2133 (N_2133,N_1434,N_1693);
nand U2134 (N_2134,N_1390,N_1327);
nand U2135 (N_2135,N_1478,N_1281);
and U2136 (N_2136,N_1484,N_1614);
or U2137 (N_2137,N_1522,N_1377);
or U2138 (N_2138,N_1806,N_1424);
nor U2139 (N_2139,N_1794,N_1404);
and U2140 (N_2140,N_1830,N_1866);
or U2141 (N_2141,N_1706,N_1323);
and U2142 (N_2142,N_1727,N_1715);
xnor U2143 (N_2143,N_1779,N_1699);
nand U2144 (N_2144,N_1724,N_1521);
nand U2145 (N_2145,N_1348,N_1299);
nor U2146 (N_2146,N_1405,N_1708);
and U2147 (N_2147,N_1380,N_1687);
and U2148 (N_2148,N_1557,N_1524);
nand U2149 (N_2149,N_1508,N_1772);
or U2150 (N_2150,N_1677,N_1726);
nand U2151 (N_2151,N_1353,N_1401);
and U2152 (N_2152,N_1367,N_1670);
nand U2153 (N_2153,N_1814,N_1592);
or U2154 (N_2154,N_1282,N_1454);
nand U2155 (N_2155,N_1791,N_1674);
and U2156 (N_2156,N_1870,N_1328);
nor U2157 (N_2157,N_1705,N_1450);
xnor U2158 (N_2158,N_1529,N_1262);
nor U2159 (N_2159,N_1583,N_1335);
nor U2160 (N_2160,N_1790,N_1653);
or U2161 (N_2161,N_1623,N_1666);
nor U2162 (N_2162,N_1513,N_1833);
nand U2163 (N_2163,N_1416,N_1306);
nand U2164 (N_2164,N_1371,N_1285);
nand U2165 (N_2165,N_1433,N_1646);
or U2166 (N_2166,N_1589,N_1514);
xnor U2167 (N_2167,N_1255,N_1333);
xnor U2168 (N_2168,N_1818,N_1512);
or U2169 (N_2169,N_1428,N_1272);
nand U2170 (N_2170,N_1874,N_1436);
and U2171 (N_2171,N_1631,N_1443);
and U2172 (N_2172,N_1846,N_1320);
nor U2173 (N_2173,N_1516,N_1502);
nor U2174 (N_2174,N_1483,N_1568);
or U2175 (N_2175,N_1842,N_1534);
nand U2176 (N_2176,N_1656,N_1582);
or U2177 (N_2177,N_1845,N_1427);
nor U2178 (N_2178,N_1504,N_1645);
nand U2179 (N_2179,N_1746,N_1590);
and U2180 (N_2180,N_1593,N_1271);
or U2181 (N_2181,N_1611,N_1391);
nor U2182 (N_2182,N_1378,N_1828);
xnor U2183 (N_2183,N_1747,N_1737);
and U2184 (N_2184,N_1558,N_1863);
nand U2185 (N_2185,N_1652,N_1491);
nor U2186 (N_2186,N_1350,N_1344);
or U2187 (N_2187,N_1499,N_1840);
nand U2188 (N_2188,N_1689,N_1637);
and U2189 (N_2189,N_1660,N_1298);
or U2190 (N_2190,N_1613,N_1410);
nor U2191 (N_2191,N_1265,N_1785);
and U2192 (N_2192,N_1781,N_1449);
and U2193 (N_2193,N_1404,N_1375);
nor U2194 (N_2194,N_1732,N_1680);
and U2195 (N_2195,N_1604,N_1290);
nand U2196 (N_2196,N_1810,N_1364);
nand U2197 (N_2197,N_1739,N_1863);
nor U2198 (N_2198,N_1521,N_1262);
and U2199 (N_2199,N_1758,N_1858);
or U2200 (N_2200,N_1556,N_1725);
nor U2201 (N_2201,N_1578,N_1745);
or U2202 (N_2202,N_1656,N_1753);
nand U2203 (N_2203,N_1408,N_1722);
xnor U2204 (N_2204,N_1314,N_1316);
and U2205 (N_2205,N_1322,N_1608);
and U2206 (N_2206,N_1433,N_1748);
and U2207 (N_2207,N_1414,N_1699);
nor U2208 (N_2208,N_1465,N_1717);
nor U2209 (N_2209,N_1655,N_1296);
nor U2210 (N_2210,N_1422,N_1702);
nor U2211 (N_2211,N_1384,N_1408);
and U2212 (N_2212,N_1452,N_1522);
nand U2213 (N_2213,N_1666,N_1475);
xnor U2214 (N_2214,N_1623,N_1322);
nand U2215 (N_2215,N_1279,N_1603);
and U2216 (N_2216,N_1429,N_1660);
nor U2217 (N_2217,N_1502,N_1609);
and U2218 (N_2218,N_1864,N_1530);
xor U2219 (N_2219,N_1801,N_1394);
nor U2220 (N_2220,N_1507,N_1533);
nand U2221 (N_2221,N_1818,N_1716);
nor U2222 (N_2222,N_1336,N_1682);
nand U2223 (N_2223,N_1759,N_1436);
and U2224 (N_2224,N_1763,N_1301);
and U2225 (N_2225,N_1636,N_1605);
nand U2226 (N_2226,N_1559,N_1294);
or U2227 (N_2227,N_1658,N_1698);
or U2228 (N_2228,N_1482,N_1641);
nor U2229 (N_2229,N_1264,N_1301);
nand U2230 (N_2230,N_1425,N_1351);
or U2231 (N_2231,N_1789,N_1462);
or U2232 (N_2232,N_1341,N_1492);
nand U2233 (N_2233,N_1874,N_1340);
and U2234 (N_2234,N_1781,N_1666);
and U2235 (N_2235,N_1351,N_1759);
nand U2236 (N_2236,N_1432,N_1434);
nand U2237 (N_2237,N_1456,N_1871);
and U2238 (N_2238,N_1392,N_1771);
xor U2239 (N_2239,N_1575,N_1508);
or U2240 (N_2240,N_1337,N_1775);
nor U2241 (N_2241,N_1615,N_1604);
and U2242 (N_2242,N_1333,N_1545);
or U2243 (N_2243,N_1716,N_1833);
and U2244 (N_2244,N_1515,N_1400);
or U2245 (N_2245,N_1517,N_1817);
or U2246 (N_2246,N_1638,N_1554);
nand U2247 (N_2247,N_1690,N_1704);
or U2248 (N_2248,N_1679,N_1322);
nand U2249 (N_2249,N_1444,N_1593);
nor U2250 (N_2250,N_1605,N_1264);
nor U2251 (N_2251,N_1671,N_1486);
nand U2252 (N_2252,N_1341,N_1448);
and U2253 (N_2253,N_1388,N_1697);
and U2254 (N_2254,N_1673,N_1298);
nor U2255 (N_2255,N_1865,N_1806);
and U2256 (N_2256,N_1451,N_1386);
and U2257 (N_2257,N_1338,N_1755);
and U2258 (N_2258,N_1530,N_1671);
and U2259 (N_2259,N_1529,N_1345);
nor U2260 (N_2260,N_1831,N_1373);
or U2261 (N_2261,N_1771,N_1507);
nor U2262 (N_2262,N_1600,N_1857);
or U2263 (N_2263,N_1453,N_1689);
xor U2264 (N_2264,N_1810,N_1475);
or U2265 (N_2265,N_1475,N_1301);
nand U2266 (N_2266,N_1872,N_1445);
nand U2267 (N_2267,N_1331,N_1303);
nand U2268 (N_2268,N_1272,N_1404);
nand U2269 (N_2269,N_1370,N_1347);
nor U2270 (N_2270,N_1599,N_1538);
nor U2271 (N_2271,N_1543,N_1423);
nand U2272 (N_2272,N_1593,N_1587);
nand U2273 (N_2273,N_1332,N_1851);
and U2274 (N_2274,N_1573,N_1691);
nor U2275 (N_2275,N_1603,N_1720);
or U2276 (N_2276,N_1330,N_1481);
and U2277 (N_2277,N_1583,N_1705);
nand U2278 (N_2278,N_1314,N_1736);
nor U2279 (N_2279,N_1604,N_1432);
and U2280 (N_2280,N_1408,N_1759);
and U2281 (N_2281,N_1806,N_1285);
nand U2282 (N_2282,N_1583,N_1702);
nor U2283 (N_2283,N_1675,N_1654);
nor U2284 (N_2284,N_1452,N_1306);
and U2285 (N_2285,N_1793,N_1593);
nand U2286 (N_2286,N_1659,N_1365);
nor U2287 (N_2287,N_1335,N_1872);
xnor U2288 (N_2288,N_1412,N_1478);
nor U2289 (N_2289,N_1820,N_1835);
nor U2290 (N_2290,N_1310,N_1444);
nand U2291 (N_2291,N_1303,N_1719);
nor U2292 (N_2292,N_1264,N_1486);
nand U2293 (N_2293,N_1376,N_1442);
nor U2294 (N_2294,N_1540,N_1409);
nand U2295 (N_2295,N_1872,N_1418);
nand U2296 (N_2296,N_1604,N_1573);
nor U2297 (N_2297,N_1291,N_1371);
nand U2298 (N_2298,N_1667,N_1476);
nor U2299 (N_2299,N_1570,N_1620);
xnor U2300 (N_2300,N_1668,N_1517);
or U2301 (N_2301,N_1614,N_1470);
nor U2302 (N_2302,N_1795,N_1392);
nor U2303 (N_2303,N_1466,N_1437);
nor U2304 (N_2304,N_1755,N_1713);
and U2305 (N_2305,N_1641,N_1457);
or U2306 (N_2306,N_1280,N_1798);
xor U2307 (N_2307,N_1264,N_1743);
and U2308 (N_2308,N_1492,N_1481);
or U2309 (N_2309,N_1762,N_1625);
nor U2310 (N_2310,N_1273,N_1428);
nor U2311 (N_2311,N_1320,N_1345);
and U2312 (N_2312,N_1647,N_1536);
nand U2313 (N_2313,N_1596,N_1314);
and U2314 (N_2314,N_1700,N_1713);
nor U2315 (N_2315,N_1791,N_1615);
nor U2316 (N_2316,N_1615,N_1775);
nor U2317 (N_2317,N_1333,N_1533);
nand U2318 (N_2318,N_1621,N_1753);
nand U2319 (N_2319,N_1521,N_1854);
nor U2320 (N_2320,N_1494,N_1342);
nor U2321 (N_2321,N_1666,N_1436);
and U2322 (N_2322,N_1269,N_1413);
and U2323 (N_2323,N_1558,N_1526);
nand U2324 (N_2324,N_1588,N_1853);
nand U2325 (N_2325,N_1450,N_1660);
nor U2326 (N_2326,N_1378,N_1518);
nand U2327 (N_2327,N_1459,N_1378);
nand U2328 (N_2328,N_1562,N_1431);
nor U2329 (N_2329,N_1638,N_1313);
nor U2330 (N_2330,N_1853,N_1559);
or U2331 (N_2331,N_1760,N_1527);
or U2332 (N_2332,N_1300,N_1837);
nand U2333 (N_2333,N_1486,N_1769);
nor U2334 (N_2334,N_1771,N_1344);
or U2335 (N_2335,N_1550,N_1449);
and U2336 (N_2336,N_1394,N_1720);
xor U2337 (N_2337,N_1635,N_1654);
and U2338 (N_2338,N_1447,N_1444);
or U2339 (N_2339,N_1546,N_1659);
or U2340 (N_2340,N_1304,N_1773);
and U2341 (N_2341,N_1427,N_1433);
and U2342 (N_2342,N_1541,N_1564);
nor U2343 (N_2343,N_1686,N_1307);
and U2344 (N_2344,N_1463,N_1280);
or U2345 (N_2345,N_1745,N_1869);
nand U2346 (N_2346,N_1478,N_1855);
xor U2347 (N_2347,N_1869,N_1435);
nor U2348 (N_2348,N_1502,N_1358);
nor U2349 (N_2349,N_1832,N_1579);
and U2350 (N_2350,N_1521,N_1361);
nor U2351 (N_2351,N_1442,N_1772);
or U2352 (N_2352,N_1806,N_1705);
xor U2353 (N_2353,N_1755,N_1853);
nor U2354 (N_2354,N_1287,N_1683);
nand U2355 (N_2355,N_1522,N_1862);
nand U2356 (N_2356,N_1700,N_1456);
or U2357 (N_2357,N_1536,N_1657);
and U2358 (N_2358,N_1274,N_1287);
and U2359 (N_2359,N_1600,N_1485);
and U2360 (N_2360,N_1374,N_1312);
xor U2361 (N_2361,N_1269,N_1381);
nand U2362 (N_2362,N_1365,N_1338);
and U2363 (N_2363,N_1274,N_1451);
nand U2364 (N_2364,N_1451,N_1276);
nor U2365 (N_2365,N_1336,N_1502);
or U2366 (N_2366,N_1549,N_1702);
nand U2367 (N_2367,N_1476,N_1412);
or U2368 (N_2368,N_1476,N_1823);
nand U2369 (N_2369,N_1326,N_1269);
and U2370 (N_2370,N_1381,N_1864);
and U2371 (N_2371,N_1259,N_1732);
nor U2372 (N_2372,N_1354,N_1297);
nand U2373 (N_2373,N_1499,N_1750);
or U2374 (N_2374,N_1365,N_1419);
nand U2375 (N_2375,N_1622,N_1867);
or U2376 (N_2376,N_1492,N_1692);
nor U2377 (N_2377,N_1450,N_1482);
xnor U2378 (N_2378,N_1320,N_1790);
xnor U2379 (N_2379,N_1662,N_1801);
nor U2380 (N_2380,N_1632,N_1345);
nand U2381 (N_2381,N_1277,N_1507);
nand U2382 (N_2382,N_1674,N_1796);
nand U2383 (N_2383,N_1521,N_1808);
and U2384 (N_2384,N_1270,N_1558);
nand U2385 (N_2385,N_1462,N_1540);
and U2386 (N_2386,N_1806,N_1507);
nand U2387 (N_2387,N_1828,N_1285);
and U2388 (N_2388,N_1270,N_1831);
nor U2389 (N_2389,N_1552,N_1268);
nand U2390 (N_2390,N_1620,N_1689);
or U2391 (N_2391,N_1526,N_1704);
nor U2392 (N_2392,N_1297,N_1310);
or U2393 (N_2393,N_1340,N_1664);
or U2394 (N_2394,N_1711,N_1678);
and U2395 (N_2395,N_1277,N_1399);
or U2396 (N_2396,N_1693,N_1477);
or U2397 (N_2397,N_1264,N_1386);
and U2398 (N_2398,N_1586,N_1746);
or U2399 (N_2399,N_1752,N_1440);
nand U2400 (N_2400,N_1695,N_1759);
nor U2401 (N_2401,N_1837,N_1871);
xor U2402 (N_2402,N_1385,N_1783);
or U2403 (N_2403,N_1844,N_1650);
or U2404 (N_2404,N_1278,N_1611);
or U2405 (N_2405,N_1573,N_1267);
xnor U2406 (N_2406,N_1710,N_1521);
and U2407 (N_2407,N_1360,N_1526);
nand U2408 (N_2408,N_1255,N_1414);
and U2409 (N_2409,N_1590,N_1641);
nor U2410 (N_2410,N_1469,N_1377);
or U2411 (N_2411,N_1295,N_1537);
nor U2412 (N_2412,N_1842,N_1428);
xnor U2413 (N_2413,N_1293,N_1378);
and U2414 (N_2414,N_1616,N_1767);
and U2415 (N_2415,N_1594,N_1714);
nand U2416 (N_2416,N_1763,N_1285);
nor U2417 (N_2417,N_1279,N_1557);
or U2418 (N_2418,N_1658,N_1864);
nor U2419 (N_2419,N_1442,N_1531);
nor U2420 (N_2420,N_1375,N_1865);
nor U2421 (N_2421,N_1483,N_1335);
or U2422 (N_2422,N_1694,N_1820);
nor U2423 (N_2423,N_1689,N_1591);
or U2424 (N_2424,N_1594,N_1519);
xnor U2425 (N_2425,N_1453,N_1468);
and U2426 (N_2426,N_1831,N_1849);
nand U2427 (N_2427,N_1827,N_1335);
nor U2428 (N_2428,N_1789,N_1561);
nor U2429 (N_2429,N_1569,N_1414);
nor U2430 (N_2430,N_1550,N_1375);
nor U2431 (N_2431,N_1301,N_1278);
xor U2432 (N_2432,N_1566,N_1529);
nor U2433 (N_2433,N_1590,N_1252);
or U2434 (N_2434,N_1733,N_1668);
or U2435 (N_2435,N_1271,N_1332);
nand U2436 (N_2436,N_1775,N_1406);
and U2437 (N_2437,N_1443,N_1669);
or U2438 (N_2438,N_1659,N_1296);
and U2439 (N_2439,N_1738,N_1362);
nor U2440 (N_2440,N_1392,N_1516);
and U2441 (N_2441,N_1417,N_1461);
or U2442 (N_2442,N_1270,N_1450);
or U2443 (N_2443,N_1464,N_1769);
or U2444 (N_2444,N_1826,N_1798);
nor U2445 (N_2445,N_1553,N_1491);
nand U2446 (N_2446,N_1758,N_1573);
nand U2447 (N_2447,N_1570,N_1665);
and U2448 (N_2448,N_1790,N_1642);
and U2449 (N_2449,N_1532,N_1704);
and U2450 (N_2450,N_1781,N_1572);
nor U2451 (N_2451,N_1486,N_1662);
or U2452 (N_2452,N_1521,N_1286);
nand U2453 (N_2453,N_1284,N_1843);
and U2454 (N_2454,N_1429,N_1765);
or U2455 (N_2455,N_1461,N_1840);
or U2456 (N_2456,N_1649,N_1676);
and U2457 (N_2457,N_1395,N_1785);
nor U2458 (N_2458,N_1285,N_1256);
nor U2459 (N_2459,N_1744,N_1550);
or U2460 (N_2460,N_1329,N_1695);
nand U2461 (N_2461,N_1626,N_1575);
nand U2462 (N_2462,N_1290,N_1582);
xor U2463 (N_2463,N_1391,N_1855);
nand U2464 (N_2464,N_1395,N_1456);
nor U2465 (N_2465,N_1344,N_1555);
or U2466 (N_2466,N_1470,N_1821);
and U2467 (N_2467,N_1782,N_1276);
and U2468 (N_2468,N_1814,N_1486);
nand U2469 (N_2469,N_1698,N_1766);
and U2470 (N_2470,N_1761,N_1451);
nor U2471 (N_2471,N_1481,N_1639);
xnor U2472 (N_2472,N_1780,N_1312);
or U2473 (N_2473,N_1750,N_1382);
and U2474 (N_2474,N_1361,N_1337);
and U2475 (N_2475,N_1764,N_1746);
xnor U2476 (N_2476,N_1676,N_1262);
nand U2477 (N_2477,N_1852,N_1748);
nor U2478 (N_2478,N_1525,N_1829);
or U2479 (N_2479,N_1686,N_1618);
nor U2480 (N_2480,N_1442,N_1642);
nand U2481 (N_2481,N_1522,N_1806);
and U2482 (N_2482,N_1611,N_1414);
nand U2483 (N_2483,N_1728,N_1419);
nor U2484 (N_2484,N_1839,N_1820);
and U2485 (N_2485,N_1770,N_1432);
nor U2486 (N_2486,N_1440,N_1525);
and U2487 (N_2487,N_1620,N_1258);
nor U2488 (N_2488,N_1481,N_1677);
nor U2489 (N_2489,N_1702,N_1765);
nor U2490 (N_2490,N_1520,N_1434);
and U2491 (N_2491,N_1318,N_1254);
and U2492 (N_2492,N_1587,N_1354);
nand U2493 (N_2493,N_1700,N_1709);
and U2494 (N_2494,N_1854,N_1329);
or U2495 (N_2495,N_1749,N_1734);
and U2496 (N_2496,N_1410,N_1497);
xnor U2497 (N_2497,N_1291,N_1772);
nand U2498 (N_2498,N_1794,N_1371);
xor U2499 (N_2499,N_1460,N_1698);
and U2500 (N_2500,N_2058,N_2467);
nor U2501 (N_2501,N_2415,N_2130);
xnor U2502 (N_2502,N_2476,N_2470);
or U2503 (N_2503,N_1880,N_2092);
or U2504 (N_2504,N_2481,N_2062);
nand U2505 (N_2505,N_2191,N_2414);
nor U2506 (N_2506,N_1932,N_2418);
nand U2507 (N_2507,N_2068,N_2320);
nor U2508 (N_2508,N_2104,N_2383);
nor U2509 (N_2509,N_1900,N_2143);
and U2510 (N_2510,N_2261,N_2405);
xor U2511 (N_2511,N_2382,N_2039);
nor U2512 (N_2512,N_2070,N_2216);
nor U2513 (N_2513,N_2228,N_2083);
nor U2514 (N_2514,N_2275,N_2100);
and U2515 (N_2515,N_2450,N_2489);
and U2516 (N_2516,N_2195,N_2443);
xor U2517 (N_2517,N_2357,N_2377);
or U2518 (N_2518,N_2018,N_2315);
or U2519 (N_2519,N_2378,N_2131);
nand U2520 (N_2520,N_2483,N_1917);
nor U2521 (N_2521,N_2333,N_2292);
nand U2522 (N_2522,N_2204,N_1918);
and U2523 (N_2523,N_2309,N_2186);
and U2524 (N_2524,N_1965,N_2269);
or U2525 (N_2525,N_2254,N_2102);
and U2526 (N_2526,N_2105,N_1936);
or U2527 (N_2527,N_2260,N_2486);
nor U2528 (N_2528,N_2087,N_2029);
or U2529 (N_2529,N_2167,N_2253);
nand U2530 (N_2530,N_2137,N_2229);
and U2531 (N_2531,N_2057,N_1958);
and U2532 (N_2532,N_2428,N_2093);
nor U2533 (N_2533,N_2053,N_2043);
nand U2534 (N_2534,N_2372,N_2111);
or U2535 (N_2535,N_2240,N_2350);
and U2536 (N_2536,N_2067,N_2471);
nand U2537 (N_2537,N_2288,N_1901);
or U2538 (N_2538,N_2017,N_2226);
nand U2539 (N_2539,N_2166,N_2252);
or U2540 (N_2540,N_2010,N_2199);
nand U2541 (N_2541,N_2213,N_2299);
or U2542 (N_2542,N_2146,N_2187);
nor U2543 (N_2543,N_2170,N_2215);
and U2544 (N_2544,N_2278,N_1927);
and U2545 (N_2545,N_2390,N_1897);
and U2546 (N_2546,N_1911,N_1984);
nor U2547 (N_2547,N_2453,N_2059);
nor U2548 (N_2548,N_2076,N_2014);
and U2549 (N_2549,N_2494,N_2395);
and U2550 (N_2550,N_2006,N_1997);
or U2551 (N_2551,N_2318,N_2074);
and U2552 (N_2552,N_2052,N_2360);
and U2553 (N_2553,N_2300,N_2343);
nor U2554 (N_2554,N_2132,N_2245);
or U2555 (N_2555,N_2060,N_1890);
nand U2556 (N_2556,N_2221,N_2123);
nor U2557 (N_2557,N_2160,N_2478);
nor U2558 (N_2558,N_2249,N_2126);
and U2559 (N_2559,N_2498,N_2273);
and U2560 (N_2560,N_2109,N_2247);
nand U2561 (N_2561,N_2487,N_2138);
nor U2562 (N_2562,N_2430,N_2466);
nand U2563 (N_2563,N_1981,N_1926);
xnor U2564 (N_2564,N_2118,N_2298);
nand U2565 (N_2565,N_2351,N_2003);
nand U2566 (N_2566,N_2075,N_2424);
or U2567 (N_2567,N_2293,N_2375);
and U2568 (N_2568,N_1899,N_2224);
nor U2569 (N_2569,N_2194,N_2331);
nand U2570 (N_2570,N_2180,N_2497);
nor U2571 (N_2571,N_2379,N_2141);
nand U2572 (N_2572,N_2369,N_2235);
nor U2573 (N_2573,N_2116,N_2363);
nand U2574 (N_2574,N_2172,N_1896);
nor U2575 (N_2575,N_2266,N_2000);
or U2576 (N_2576,N_2044,N_2230);
and U2577 (N_2577,N_1877,N_2295);
and U2578 (N_2578,N_2054,N_2150);
nand U2579 (N_2579,N_2165,N_2262);
or U2580 (N_2580,N_1923,N_2055);
xnor U2581 (N_2581,N_1971,N_1912);
or U2582 (N_2582,N_2308,N_2163);
nand U2583 (N_2583,N_2020,N_1980);
and U2584 (N_2584,N_2177,N_2162);
and U2585 (N_2585,N_1938,N_2297);
nand U2586 (N_2586,N_2251,N_2312);
nand U2587 (N_2587,N_2182,N_2242);
nand U2588 (N_2588,N_2041,N_2090);
and U2589 (N_2589,N_2038,N_2119);
nand U2590 (N_2590,N_2272,N_2339);
and U2591 (N_2591,N_1992,N_2304);
or U2592 (N_2592,N_2499,N_2460);
xor U2593 (N_2593,N_2197,N_2432);
nor U2594 (N_2594,N_2496,N_2371);
and U2595 (N_2595,N_2101,N_2337);
nand U2596 (N_2596,N_2473,N_2211);
nor U2597 (N_2597,N_2133,N_2362);
and U2598 (N_2598,N_2155,N_2189);
or U2599 (N_2599,N_2386,N_2484);
nand U2600 (N_2600,N_1875,N_1937);
and U2601 (N_2601,N_1895,N_2277);
and U2602 (N_2602,N_1940,N_2482);
nand U2603 (N_2603,N_2366,N_2113);
nor U2604 (N_2604,N_2169,N_2107);
nor U2605 (N_2605,N_2349,N_2411);
nand U2606 (N_2606,N_2238,N_1915);
or U2607 (N_2607,N_2144,N_2088);
nor U2608 (N_2608,N_1952,N_2358);
or U2609 (N_2609,N_2399,N_2417);
or U2610 (N_2610,N_2400,N_2079);
xor U2611 (N_2611,N_2294,N_1922);
and U2612 (N_2612,N_2050,N_2394);
nor U2613 (N_2613,N_1916,N_2056);
or U2614 (N_2614,N_2329,N_2196);
nor U2615 (N_2615,N_1907,N_2124);
and U2616 (N_2616,N_1930,N_2462);
or U2617 (N_2617,N_1882,N_1985);
and U2618 (N_2618,N_2396,N_1969);
xnor U2619 (N_2619,N_2422,N_2227);
xnor U2620 (N_2620,N_2434,N_2361);
nor U2621 (N_2621,N_2209,N_2457);
nor U2622 (N_2622,N_2158,N_2178);
xnor U2623 (N_2623,N_2220,N_2480);
nor U2624 (N_2624,N_2276,N_2225);
nand U2625 (N_2625,N_1974,N_1941);
nand U2626 (N_2626,N_1905,N_2112);
nand U2627 (N_2627,N_2491,N_2028);
nor U2628 (N_2628,N_2336,N_1995);
and U2629 (N_2629,N_2125,N_2461);
nand U2630 (N_2630,N_2449,N_2135);
or U2631 (N_2631,N_1904,N_2072);
xor U2632 (N_2632,N_2232,N_1892);
and U2633 (N_2633,N_1964,N_2202);
or U2634 (N_2634,N_2286,N_2246);
nor U2635 (N_2635,N_1948,N_2192);
nor U2636 (N_2636,N_2420,N_2136);
nor U2637 (N_2637,N_2139,N_2456);
or U2638 (N_2638,N_2179,N_2370);
xor U2639 (N_2639,N_1881,N_2392);
nor U2640 (N_2640,N_2183,N_2064);
nand U2641 (N_2641,N_2021,N_2485);
nor U2642 (N_2642,N_2475,N_2344);
or U2643 (N_2643,N_2368,N_2425);
xor U2644 (N_2644,N_1902,N_2103);
or U2645 (N_2645,N_2448,N_2340);
nor U2646 (N_2646,N_2347,N_2413);
nand U2647 (N_2647,N_1994,N_2019);
and U2648 (N_2648,N_2152,N_2419);
nand U2649 (N_2649,N_2151,N_2001);
xnor U2650 (N_2650,N_2009,N_2231);
and U2651 (N_2651,N_2374,N_1913);
and U2652 (N_2652,N_2463,N_2157);
nor U2653 (N_2653,N_2129,N_2200);
nor U2654 (N_2654,N_2237,N_1920);
nand U2655 (N_2655,N_2317,N_2048);
and U2656 (N_2656,N_2316,N_1998);
or U2657 (N_2657,N_2205,N_1963);
or U2658 (N_2658,N_2065,N_2081);
nor U2659 (N_2659,N_2441,N_2373);
nand U2660 (N_2660,N_2469,N_1943);
or U2661 (N_2661,N_2389,N_1956);
nor U2662 (N_2662,N_1959,N_2325);
nor U2663 (N_2663,N_2012,N_1960);
nor U2664 (N_2664,N_2433,N_2218);
or U2665 (N_2665,N_1977,N_2250);
nor U2666 (N_2666,N_2168,N_2359);
or U2667 (N_2667,N_2410,N_2032);
nor U2668 (N_2668,N_2330,N_2025);
nor U2669 (N_2669,N_2206,N_2270);
and U2670 (N_2670,N_1898,N_1942);
nor U2671 (N_2671,N_2036,N_2356);
or U2672 (N_2672,N_1925,N_2365);
nor U2673 (N_2673,N_2490,N_2134);
nand U2674 (N_2674,N_2352,N_2004);
nor U2675 (N_2675,N_2281,N_2442);
nand U2676 (N_2676,N_2397,N_2030);
and U2677 (N_2677,N_2338,N_2243);
and U2678 (N_2678,N_2007,N_2345);
nor U2679 (N_2679,N_2439,N_2033);
or U2680 (N_2680,N_2174,N_2259);
nand U2681 (N_2681,N_2284,N_2128);
or U2682 (N_2682,N_2042,N_1946);
nand U2683 (N_2683,N_2429,N_1909);
and U2684 (N_2684,N_2289,N_2106);
or U2685 (N_2685,N_2306,N_2114);
xor U2686 (N_2686,N_2069,N_2376);
nand U2687 (N_2687,N_2073,N_2279);
xor U2688 (N_2688,N_1894,N_2302);
and U2689 (N_2689,N_2207,N_2412);
or U2690 (N_2690,N_2334,N_1953);
nor U2691 (N_2691,N_2321,N_2203);
and U2692 (N_2692,N_2091,N_2263);
and U2693 (N_2693,N_2409,N_2437);
and U2694 (N_2694,N_1986,N_2353);
xor U2695 (N_2695,N_1954,N_2013);
nor U2696 (N_2696,N_1990,N_1944);
nand U2697 (N_2697,N_2035,N_2401);
and U2698 (N_2698,N_2346,N_2492);
and U2699 (N_2699,N_1983,N_2099);
nor U2700 (N_2700,N_1939,N_2154);
nand U2701 (N_2701,N_2431,N_2305);
or U2702 (N_2702,N_2078,N_1879);
nor U2703 (N_2703,N_2140,N_2061);
or U2704 (N_2704,N_2219,N_2464);
nor U2705 (N_2705,N_2193,N_1910);
nand U2706 (N_2706,N_1955,N_2444);
nor U2707 (N_2707,N_2217,N_2117);
xor U2708 (N_2708,N_2089,N_2016);
nand U2709 (N_2709,N_1949,N_2084);
and U2710 (N_2710,N_2427,N_2472);
or U2711 (N_2711,N_2233,N_2324);
nand U2712 (N_2712,N_2108,N_1968);
nand U2713 (N_2713,N_2326,N_2077);
nor U2714 (N_2714,N_2188,N_2436);
or U2715 (N_2715,N_2115,N_2313);
xnor U2716 (N_2716,N_2291,N_2267);
nand U2717 (N_2717,N_2208,N_2094);
xor U2718 (N_2718,N_2488,N_2301);
and U2719 (N_2719,N_1924,N_1886);
and U2720 (N_2720,N_1906,N_2381);
nor U2721 (N_2721,N_2348,N_2364);
nor U2722 (N_2722,N_1934,N_1950);
nor U2723 (N_2723,N_1891,N_2287);
and U2724 (N_2724,N_2011,N_2082);
nand U2725 (N_2725,N_2459,N_2223);
nand U2726 (N_2726,N_2264,N_2244);
xnor U2727 (N_2727,N_2047,N_1935);
and U2728 (N_2728,N_1903,N_1884);
nand U2729 (N_2729,N_2455,N_1921);
or U2730 (N_2730,N_2477,N_2282);
nand U2731 (N_2731,N_2495,N_2307);
and U2732 (N_2732,N_2127,N_1893);
or U2733 (N_2733,N_2098,N_2468);
nand U2734 (N_2734,N_2095,N_1979);
nand U2735 (N_2735,N_2319,N_2066);
and U2736 (N_2736,N_2008,N_1883);
and U2737 (N_2737,N_2274,N_2387);
nand U2738 (N_2738,N_2447,N_1982);
xor U2739 (N_2739,N_2406,N_2049);
or U2740 (N_2740,N_2239,N_2384);
nand U2741 (N_2741,N_1929,N_2451);
and U2742 (N_2742,N_2438,N_2142);
nor U2743 (N_2743,N_1888,N_1878);
or U2744 (N_2744,N_2148,N_2005);
nor U2745 (N_2745,N_2022,N_2423);
nand U2746 (N_2746,N_1978,N_2175);
nor U2747 (N_2747,N_1988,N_2421);
nand U2748 (N_2748,N_1975,N_1933);
nand U2749 (N_2749,N_2190,N_1973);
nand U2750 (N_2750,N_2290,N_2380);
nand U2751 (N_2751,N_2121,N_2474);
nand U2752 (N_2752,N_2173,N_2161);
and U2753 (N_2753,N_2285,N_2402);
nor U2754 (N_2754,N_2096,N_2322);
nand U2755 (N_2755,N_2002,N_2385);
and U2756 (N_2756,N_2446,N_2236);
nor U2757 (N_2757,N_2086,N_2388);
or U2758 (N_2758,N_2097,N_1889);
or U2759 (N_2759,N_1887,N_2452);
nor U2760 (N_2760,N_2164,N_2031);
or U2761 (N_2761,N_1951,N_2256);
xor U2762 (N_2762,N_2214,N_1972);
xnor U2763 (N_2763,N_2398,N_1885);
or U2764 (N_2764,N_2332,N_2335);
or U2765 (N_2765,N_2391,N_2147);
or U2766 (N_2766,N_1967,N_1876);
and U2767 (N_2767,N_2257,N_1962);
nand U2768 (N_2768,N_1966,N_2258);
or U2769 (N_2769,N_1996,N_2440);
xnor U2770 (N_2770,N_2110,N_2342);
and U2771 (N_2771,N_2328,N_2458);
nor U2772 (N_2772,N_2303,N_1991);
nor U2773 (N_2773,N_2210,N_2185);
nand U2774 (N_2774,N_2037,N_2063);
nand U2775 (N_2775,N_2255,N_2493);
nor U2776 (N_2776,N_2241,N_2046);
or U2777 (N_2777,N_2171,N_2407);
xnor U2778 (N_2778,N_2034,N_2341);
and U2779 (N_2779,N_2153,N_2181);
nor U2780 (N_2780,N_2045,N_2404);
and U2781 (N_2781,N_2367,N_1957);
nor U2782 (N_2782,N_2122,N_2015);
or U2783 (N_2783,N_2201,N_2234);
or U2784 (N_2784,N_1987,N_2040);
or U2785 (N_2785,N_2176,N_1947);
nor U2786 (N_2786,N_1914,N_2071);
or U2787 (N_2787,N_2479,N_2271);
nand U2788 (N_2788,N_2184,N_2355);
nor U2789 (N_2789,N_2159,N_2435);
and U2790 (N_2790,N_2354,N_2026);
nand U2791 (N_2791,N_2248,N_2323);
nor U2792 (N_2792,N_2156,N_1999);
or U2793 (N_2793,N_2296,N_1945);
and U2794 (N_2794,N_1993,N_1989);
and U2795 (N_2795,N_2393,N_2310);
nand U2796 (N_2796,N_2314,N_2023);
or U2797 (N_2797,N_1931,N_2426);
and U2798 (N_2798,N_2416,N_1961);
nand U2799 (N_2799,N_1919,N_2212);
nand U2800 (N_2800,N_1908,N_2085);
nor U2801 (N_2801,N_2149,N_2265);
nor U2802 (N_2802,N_2327,N_1928);
xnor U2803 (N_2803,N_2445,N_2027);
and U2804 (N_2804,N_2198,N_2454);
xnor U2805 (N_2805,N_2051,N_1976);
or U2806 (N_2806,N_2311,N_2280);
or U2807 (N_2807,N_2268,N_2408);
nand U2808 (N_2808,N_2283,N_2120);
and U2809 (N_2809,N_2080,N_2403);
or U2810 (N_2810,N_2145,N_2465);
nand U2811 (N_2811,N_2222,N_2024);
xnor U2812 (N_2812,N_1970,N_1951);
and U2813 (N_2813,N_2319,N_2206);
and U2814 (N_2814,N_1961,N_2012);
nor U2815 (N_2815,N_2208,N_2378);
or U2816 (N_2816,N_2139,N_2217);
and U2817 (N_2817,N_2182,N_1980);
nor U2818 (N_2818,N_2042,N_2415);
xnor U2819 (N_2819,N_2174,N_2104);
or U2820 (N_2820,N_1890,N_2256);
nand U2821 (N_2821,N_2329,N_2275);
or U2822 (N_2822,N_1992,N_1997);
and U2823 (N_2823,N_2118,N_1880);
nand U2824 (N_2824,N_1954,N_2362);
or U2825 (N_2825,N_2417,N_2361);
and U2826 (N_2826,N_1876,N_2298);
nor U2827 (N_2827,N_2393,N_2166);
xor U2828 (N_2828,N_2211,N_2486);
nand U2829 (N_2829,N_2104,N_2367);
nor U2830 (N_2830,N_2457,N_2249);
or U2831 (N_2831,N_2305,N_2287);
or U2832 (N_2832,N_2127,N_2215);
or U2833 (N_2833,N_2208,N_2464);
and U2834 (N_2834,N_2361,N_2227);
nor U2835 (N_2835,N_2321,N_1971);
and U2836 (N_2836,N_2242,N_2038);
nand U2837 (N_2837,N_2370,N_2386);
nor U2838 (N_2838,N_1947,N_1909);
nor U2839 (N_2839,N_2001,N_2319);
and U2840 (N_2840,N_2033,N_2238);
and U2841 (N_2841,N_2487,N_2086);
nor U2842 (N_2842,N_1883,N_2039);
nand U2843 (N_2843,N_1908,N_2403);
or U2844 (N_2844,N_2187,N_2345);
xor U2845 (N_2845,N_2049,N_1924);
or U2846 (N_2846,N_2126,N_2109);
and U2847 (N_2847,N_2053,N_2128);
xnor U2848 (N_2848,N_2414,N_2030);
nor U2849 (N_2849,N_2005,N_2196);
or U2850 (N_2850,N_2084,N_2070);
nor U2851 (N_2851,N_2008,N_2059);
nor U2852 (N_2852,N_2219,N_2439);
or U2853 (N_2853,N_1926,N_2381);
or U2854 (N_2854,N_1954,N_2024);
nor U2855 (N_2855,N_1962,N_2333);
nand U2856 (N_2856,N_2444,N_2129);
or U2857 (N_2857,N_2022,N_1908);
or U2858 (N_2858,N_2319,N_2371);
xnor U2859 (N_2859,N_2011,N_2307);
and U2860 (N_2860,N_2209,N_2056);
nor U2861 (N_2861,N_2326,N_2296);
and U2862 (N_2862,N_2431,N_2446);
nand U2863 (N_2863,N_2184,N_2494);
nor U2864 (N_2864,N_1900,N_2295);
nand U2865 (N_2865,N_1951,N_2345);
nand U2866 (N_2866,N_2284,N_2202);
nand U2867 (N_2867,N_2360,N_1916);
nor U2868 (N_2868,N_2022,N_2014);
nand U2869 (N_2869,N_2074,N_2097);
nand U2870 (N_2870,N_2339,N_1963);
nor U2871 (N_2871,N_2275,N_2219);
nand U2872 (N_2872,N_2445,N_2120);
and U2873 (N_2873,N_2200,N_1972);
xor U2874 (N_2874,N_2097,N_2445);
nand U2875 (N_2875,N_2457,N_2332);
xnor U2876 (N_2876,N_2236,N_2275);
and U2877 (N_2877,N_1931,N_2463);
or U2878 (N_2878,N_2292,N_2093);
or U2879 (N_2879,N_2443,N_1941);
and U2880 (N_2880,N_2440,N_2012);
or U2881 (N_2881,N_2242,N_2368);
nand U2882 (N_2882,N_2115,N_2220);
and U2883 (N_2883,N_1928,N_2287);
and U2884 (N_2884,N_2140,N_1918);
and U2885 (N_2885,N_2135,N_2413);
and U2886 (N_2886,N_2237,N_2030);
nor U2887 (N_2887,N_2144,N_2007);
or U2888 (N_2888,N_2349,N_2243);
nor U2889 (N_2889,N_1989,N_2436);
or U2890 (N_2890,N_2011,N_2047);
nand U2891 (N_2891,N_2307,N_2059);
nand U2892 (N_2892,N_2119,N_2275);
nor U2893 (N_2893,N_2119,N_2178);
and U2894 (N_2894,N_2474,N_2223);
nor U2895 (N_2895,N_2252,N_2186);
and U2896 (N_2896,N_2271,N_2409);
nand U2897 (N_2897,N_2431,N_1877);
nand U2898 (N_2898,N_1946,N_1926);
or U2899 (N_2899,N_2198,N_1909);
and U2900 (N_2900,N_2402,N_2471);
nand U2901 (N_2901,N_2366,N_2122);
xor U2902 (N_2902,N_1980,N_2152);
and U2903 (N_2903,N_2351,N_2214);
xor U2904 (N_2904,N_2417,N_2259);
and U2905 (N_2905,N_2000,N_2173);
nor U2906 (N_2906,N_2039,N_2129);
nor U2907 (N_2907,N_2355,N_2055);
and U2908 (N_2908,N_1895,N_2129);
and U2909 (N_2909,N_2485,N_2428);
nand U2910 (N_2910,N_1894,N_2214);
xor U2911 (N_2911,N_2054,N_1933);
nor U2912 (N_2912,N_2190,N_2428);
nor U2913 (N_2913,N_2182,N_1929);
and U2914 (N_2914,N_2496,N_2285);
nor U2915 (N_2915,N_2063,N_2492);
or U2916 (N_2916,N_2025,N_2077);
and U2917 (N_2917,N_2017,N_1946);
nand U2918 (N_2918,N_2465,N_2138);
or U2919 (N_2919,N_2241,N_1996);
nand U2920 (N_2920,N_2266,N_2214);
or U2921 (N_2921,N_1927,N_2366);
nor U2922 (N_2922,N_1905,N_2328);
nand U2923 (N_2923,N_2243,N_2329);
nor U2924 (N_2924,N_1913,N_2263);
nor U2925 (N_2925,N_1963,N_2120);
nor U2926 (N_2926,N_2087,N_2256);
and U2927 (N_2927,N_2129,N_2163);
or U2928 (N_2928,N_2184,N_2140);
or U2929 (N_2929,N_2029,N_2392);
or U2930 (N_2930,N_2267,N_2456);
or U2931 (N_2931,N_2347,N_2161);
or U2932 (N_2932,N_2366,N_2441);
or U2933 (N_2933,N_2372,N_2494);
nor U2934 (N_2934,N_1934,N_2259);
nand U2935 (N_2935,N_2259,N_2243);
and U2936 (N_2936,N_2278,N_2487);
and U2937 (N_2937,N_1984,N_2477);
or U2938 (N_2938,N_2036,N_2402);
nor U2939 (N_2939,N_2446,N_2464);
nand U2940 (N_2940,N_2213,N_2375);
nand U2941 (N_2941,N_2103,N_1966);
nor U2942 (N_2942,N_2409,N_2217);
nor U2943 (N_2943,N_2353,N_2149);
nand U2944 (N_2944,N_2417,N_2446);
or U2945 (N_2945,N_2032,N_2365);
or U2946 (N_2946,N_2355,N_2162);
and U2947 (N_2947,N_2234,N_2336);
or U2948 (N_2948,N_2275,N_2380);
nor U2949 (N_2949,N_2046,N_2354);
and U2950 (N_2950,N_1928,N_2435);
nand U2951 (N_2951,N_2020,N_2487);
nand U2952 (N_2952,N_2072,N_2050);
or U2953 (N_2953,N_1889,N_2200);
or U2954 (N_2954,N_2223,N_2426);
or U2955 (N_2955,N_2278,N_2306);
and U2956 (N_2956,N_2150,N_2099);
nor U2957 (N_2957,N_2088,N_1935);
nor U2958 (N_2958,N_2324,N_2115);
and U2959 (N_2959,N_2145,N_1906);
nand U2960 (N_2960,N_2363,N_2059);
or U2961 (N_2961,N_2459,N_2346);
nor U2962 (N_2962,N_2358,N_2416);
or U2963 (N_2963,N_2453,N_1943);
and U2964 (N_2964,N_2121,N_2429);
nor U2965 (N_2965,N_2490,N_2320);
and U2966 (N_2966,N_1885,N_2391);
xor U2967 (N_2967,N_2256,N_2167);
nand U2968 (N_2968,N_2262,N_2205);
and U2969 (N_2969,N_2453,N_1983);
xnor U2970 (N_2970,N_2499,N_2262);
nor U2971 (N_2971,N_2158,N_2029);
xnor U2972 (N_2972,N_2188,N_2016);
and U2973 (N_2973,N_2341,N_2195);
xnor U2974 (N_2974,N_2211,N_2333);
or U2975 (N_2975,N_2111,N_2004);
or U2976 (N_2976,N_2456,N_2360);
or U2977 (N_2977,N_2078,N_2470);
or U2978 (N_2978,N_1932,N_2476);
nand U2979 (N_2979,N_2392,N_2013);
or U2980 (N_2980,N_2187,N_2078);
nor U2981 (N_2981,N_1979,N_2129);
nor U2982 (N_2982,N_2298,N_2094);
nor U2983 (N_2983,N_1953,N_1951);
or U2984 (N_2984,N_2026,N_1927);
and U2985 (N_2985,N_2049,N_2060);
xnor U2986 (N_2986,N_2056,N_2240);
nand U2987 (N_2987,N_2311,N_2339);
xor U2988 (N_2988,N_2042,N_2412);
nand U2989 (N_2989,N_2302,N_2165);
xor U2990 (N_2990,N_2283,N_2295);
nand U2991 (N_2991,N_1879,N_2033);
or U2992 (N_2992,N_2041,N_2473);
nand U2993 (N_2993,N_2472,N_2166);
or U2994 (N_2994,N_1901,N_2385);
and U2995 (N_2995,N_2345,N_2057);
nand U2996 (N_2996,N_2213,N_2285);
nor U2997 (N_2997,N_2013,N_1917);
or U2998 (N_2998,N_2278,N_2202);
and U2999 (N_2999,N_2247,N_2226);
and U3000 (N_3000,N_1980,N_2381);
nand U3001 (N_3001,N_2482,N_2373);
and U3002 (N_3002,N_2008,N_2156);
nand U3003 (N_3003,N_2431,N_2117);
nand U3004 (N_3004,N_2321,N_1933);
nand U3005 (N_3005,N_2191,N_2261);
or U3006 (N_3006,N_2391,N_1966);
or U3007 (N_3007,N_2142,N_1944);
nor U3008 (N_3008,N_2447,N_2075);
nor U3009 (N_3009,N_1953,N_2250);
nand U3010 (N_3010,N_1927,N_2216);
nand U3011 (N_3011,N_2359,N_2068);
nand U3012 (N_3012,N_2275,N_2387);
xor U3013 (N_3013,N_2010,N_2312);
and U3014 (N_3014,N_2424,N_2257);
nand U3015 (N_3015,N_2239,N_2152);
nor U3016 (N_3016,N_2245,N_2135);
nor U3017 (N_3017,N_2452,N_2174);
and U3018 (N_3018,N_2378,N_2202);
and U3019 (N_3019,N_1946,N_2128);
nor U3020 (N_3020,N_2394,N_2224);
or U3021 (N_3021,N_2166,N_2000);
nand U3022 (N_3022,N_1958,N_1997);
nand U3023 (N_3023,N_2062,N_2188);
nand U3024 (N_3024,N_2094,N_2340);
nor U3025 (N_3025,N_2463,N_2313);
nor U3026 (N_3026,N_1887,N_2375);
nand U3027 (N_3027,N_1987,N_2059);
nand U3028 (N_3028,N_2403,N_2235);
nand U3029 (N_3029,N_1960,N_2179);
nor U3030 (N_3030,N_2208,N_1909);
or U3031 (N_3031,N_2476,N_2398);
nor U3032 (N_3032,N_1927,N_2159);
and U3033 (N_3033,N_2081,N_2132);
nor U3034 (N_3034,N_2248,N_2073);
or U3035 (N_3035,N_2131,N_2199);
and U3036 (N_3036,N_2187,N_2371);
or U3037 (N_3037,N_2304,N_2376);
or U3038 (N_3038,N_2139,N_1904);
nor U3039 (N_3039,N_2403,N_2200);
nor U3040 (N_3040,N_1969,N_1947);
nand U3041 (N_3041,N_2359,N_2207);
and U3042 (N_3042,N_2228,N_2428);
or U3043 (N_3043,N_1897,N_1914);
or U3044 (N_3044,N_1970,N_2327);
or U3045 (N_3045,N_2335,N_2005);
nand U3046 (N_3046,N_2073,N_2209);
xnor U3047 (N_3047,N_2329,N_2197);
xor U3048 (N_3048,N_2017,N_2280);
nand U3049 (N_3049,N_2289,N_1949);
and U3050 (N_3050,N_2485,N_2481);
nor U3051 (N_3051,N_2425,N_2400);
and U3052 (N_3052,N_1998,N_2492);
nand U3053 (N_3053,N_2258,N_2170);
or U3054 (N_3054,N_2304,N_1875);
or U3055 (N_3055,N_2312,N_1945);
nor U3056 (N_3056,N_2422,N_2150);
and U3057 (N_3057,N_2465,N_2203);
nor U3058 (N_3058,N_2377,N_2096);
and U3059 (N_3059,N_2485,N_1891);
nand U3060 (N_3060,N_2365,N_2266);
nor U3061 (N_3061,N_2437,N_2485);
and U3062 (N_3062,N_2300,N_1882);
xor U3063 (N_3063,N_1945,N_2301);
and U3064 (N_3064,N_1894,N_2002);
nand U3065 (N_3065,N_2161,N_2155);
nor U3066 (N_3066,N_2344,N_2346);
nand U3067 (N_3067,N_2236,N_2127);
nor U3068 (N_3068,N_2377,N_2064);
and U3069 (N_3069,N_2113,N_2440);
nor U3070 (N_3070,N_2275,N_2403);
or U3071 (N_3071,N_1992,N_2348);
and U3072 (N_3072,N_1882,N_2216);
xor U3073 (N_3073,N_2410,N_2466);
nand U3074 (N_3074,N_1946,N_2251);
nand U3075 (N_3075,N_2466,N_2258);
xnor U3076 (N_3076,N_2117,N_2127);
nand U3077 (N_3077,N_2157,N_2146);
nor U3078 (N_3078,N_2398,N_2416);
and U3079 (N_3079,N_1956,N_1904);
nand U3080 (N_3080,N_2117,N_2193);
nand U3081 (N_3081,N_2494,N_2140);
or U3082 (N_3082,N_2399,N_2401);
nand U3083 (N_3083,N_2422,N_1921);
or U3084 (N_3084,N_2034,N_2191);
nor U3085 (N_3085,N_2495,N_2174);
nand U3086 (N_3086,N_2481,N_2254);
nand U3087 (N_3087,N_2115,N_2416);
and U3088 (N_3088,N_1912,N_1891);
or U3089 (N_3089,N_2326,N_2091);
or U3090 (N_3090,N_2126,N_2216);
nor U3091 (N_3091,N_2163,N_2447);
and U3092 (N_3092,N_2256,N_2093);
and U3093 (N_3093,N_2471,N_2347);
nand U3094 (N_3094,N_2102,N_2289);
nor U3095 (N_3095,N_2213,N_1910);
nand U3096 (N_3096,N_1891,N_2275);
nand U3097 (N_3097,N_2485,N_2067);
and U3098 (N_3098,N_2453,N_1955);
nor U3099 (N_3099,N_2458,N_2071);
or U3100 (N_3100,N_2189,N_1988);
or U3101 (N_3101,N_2166,N_2081);
nand U3102 (N_3102,N_2445,N_2155);
or U3103 (N_3103,N_2057,N_2178);
nor U3104 (N_3104,N_2472,N_1969);
nor U3105 (N_3105,N_2219,N_2226);
or U3106 (N_3106,N_2142,N_1957);
or U3107 (N_3107,N_1918,N_1885);
nor U3108 (N_3108,N_2114,N_2352);
xor U3109 (N_3109,N_2283,N_1976);
nor U3110 (N_3110,N_2307,N_1984);
or U3111 (N_3111,N_2185,N_2220);
and U3112 (N_3112,N_2140,N_2466);
and U3113 (N_3113,N_2413,N_2328);
or U3114 (N_3114,N_2274,N_2402);
or U3115 (N_3115,N_2409,N_2418);
nand U3116 (N_3116,N_2052,N_2287);
or U3117 (N_3117,N_2382,N_1952);
nor U3118 (N_3118,N_2362,N_2348);
nor U3119 (N_3119,N_1948,N_2100);
and U3120 (N_3120,N_1887,N_2078);
or U3121 (N_3121,N_1878,N_2242);
nor U3122 (N_3122,N_2438,N_2236);
nand U3123 (N_3123,N_1883,N_2308);
and U3124 (N_3124,N_2017,N_2181);
nor U3125 (N_3125,N_2619,N_2939);
nor U3126 (N_3126,N_2931,N_3112);
or U3127 (N_3127,N_2683,N_2570);
xor U3128 (N_3128,N_2995,N_2775);
nor U3129 (N_3129,N_2998,N_3050);
or U3130 (N_3130,N_2624,N_2513);
nor U3131 (N_3131,N_2906,N_2527);
nand U3132 (N_3132,N_2980,N_2793);
or U3133 (N_3133,N_2714,N_2745);
nor U3134 (N_3134,N_2973,N_2728);
nor U3135 (N_3135,N_2936,N_2718);
or U3136 (N_3136,N_3015,N_2890);
and U3137 (N_3137,N_2934,N_2979);
nor U3138 (N_3138,N_3027,N_2815);
or U3139 (N_3139,N_2960,N_3076);
or U3140 (N_3140,N_2811,N_2644);
xnor U3141 (N_3141,N_3046,N_2523);
xor U3142 (N_3142,N_2877,N_2717);
nand U3143 (N_3143,N_2525,N_2804);
nor U3144 (N_3144,N_3007,N_2556);
or U3145 (N_3145,N_2514,N_2983);
nor U3146 (N_3146,N_2614,N_2836);
xnor U3147 (N_3147,N_2872,N_3065);
and U3148 (N_3148,N_2536,N_3040);
or U3149 (N_3149,N_2641,N_2774);
and U3150 (N_3150,N_2582,N_2542);
nor U3151 (N_3151,N_2835,N_2583);
and U3152 (N_3152,N_2638,N_2657);
and U3153 (N_3153,N_2511,N_2862);
and U3154 (N_3154,N_3092,N_2585);
nand U3155 (N_3155,N_2598,N_2561);
or U3156 (N_3156,N_2531,N_2984);
or U3157 (N_3157,N_3091,N_2504);
or U3158 (N_3158,N_2551,N_2682);
and U3159 (N_3159,N_2882,N_3104);
nand U3160 (N_3160,N_2897,N_2746);
and U3161 (N_3161,N_3022,N_2944);
xor U3162 (N_3162,N_2517,N_2950);
nand U3163 (N_3163,N_2956,N_3055);
nor U3164 (N_3164,N_2807,N_3036);
and U3165 (N_3165,N_2866,N_2978);
nor U3166 (N_3166,N_3048,N_2557);
nand U3167 (N_3167,N_2781,N_2613);
or U3168 (N_3168,N_2846,N_2732);
and U3169 (N_3169,N_2662,N_2798);
and U3170 (N_3170,N_2865,N_2850);
and U3171 (N_3171,N_2630,N_2658);
nor U3172 (N_3172,N_3062,N_3071);
and U3173 (N_3173,N_2819,N_2832);
nor U3174 (N_3174,N_3115,N_2792);
nor U3175 (N_3175,N_3008,N_2773);
nor U3176 (N_3176,N_2706,N_2867);
and U3177 (N_3177,N_2823,N_2675);
nand U3178 (N_3178,N_2629,N_2785);
or U3179 (N_3179,N_2711,N_2601);
nand U3180 (N_3180,N_2526,N_2818);
nand U3181 (N_3181,N_2584,N_2660);
nand U3182 (N_3182,N_2626,N_2989);
nor U3183 (N_3183,N_2666,N_2809);
and U3184 (N_3184,N_2903,N_2919);
nand U3185 (N_3185,N_2744,N_3069);
and U3186 (N_3186,N_3045,N_2516);
nand U3187 (N_3187,N_2668,N_3032);
and U3188 (N_3188,N_2825,N_2547);
nor U3189 (N_3189,N_2565,N_3090);
nand U3190 (N_3190,N_3074,N_3081);
and U3191 (N_3191,N_3026,N_2680);
nand U3192 (N_3192,N_2560,N_2749);
and U3193 (N_3193,N_3020,N_2889);
nor U3194 (N_3194,N_3005,N_3017);
nor U3195 (N_3195,N_2596,N_2620);
and U3196 (N_3196,N_3099,N_2945);
and U3197 (N_3197,N_2741,N_3052);
nor U3198 (N_3198,N_2697,N_2564);
and U3199 (N_3199,N_2966,N_2648);
nand U3200 (N_3200,N_2802,N_3039);
nor U3201 (N_3201,N_2821,N_2698);
and U3202 (N_3202,N_3021,N_2719);
and U3203 (N_3203,N_2722,N_2841);
nor U3204 (N_3204,N_2669,N_2827);
or U3205 (N_3205,N_3029,N_2948);
and U3206 (N_3206,N_2873,N_2767);
xnor U3207 (N_3207,N_2766,N_2856);
nor U3208 (N_3208,N_2876,N_2577);
or U3209 (N_3209,N_2656,N_2927);
or U3210 (N_3210,N_2911,N_2625);
xnor U3211 (N_3211,N_2687,N_2600);
nor U3212 (N_3212,N_2958,N_2685);
and U3213 (N_3213,N_2868,N_3035);
nor U3214 (N_3214,N_2587,N_2772);
nor U3215 (N_3215,N_2503,N_2521);
nor U3216 (N_3216,N_2691,N_2590);
nor U3217 (N_3217,N_2534,N_2591);
and U3218 (N_3218,N_2949,N_2705);
xor U3219 (N_3219,N_2935,N_2552);
xor U3220 (N_3220,N_2957,N_2729);
nand U3221 (N_3221,N_2593,N_2883);
and U3222 (N_3222,N_2992,N_2743);
nor U3223 (N_3223,N_2559,N_2954);
and U3224 (N_3224,N_2840,N_2864);
xnor U3225 (N_3225,N_3108,N_2830);
xor U3226 (N_3226,N_2797,N_2849);
and U3227 (N_3227,N_2971,N_2922);
nor U3228 (N_3228,N_3031,N_2893);
or U3229 (N_3229,N_2636,N_2932);
nand U3230 (N_3230,N_3094,N_2963);
and U3231 (N_3231,N_2887,N_2839);
nor U3232 (N_3232,N_2970,N_3058);
nand U3233 (N_3233,N_2814,N_2871);
or U3234 (N_3234,N_2885,N_2723);
nor U3235 (N_3235,N_3066,N_2908);
xor U3236 (N_3236,N_2533,N_2953);
or U3237 (N_3237,N_2817,N_2962);
xnor U3238 (N_3238,N_2579,N_2972);
nor U3239 (N_3239,N_2770,N_2920);
and U3240 (N_3240,N_3080,N_2747);
and U3241 (N_3241,N_2505,N_2771);
and U3242 (N_3242,N_2586,N_3087);
or U3243 (N_3243,N_3059,N_2681);
and U3244 (N_3244,N_2928,N_2667);
or U3245 (N_3245,N_2627,N_2813);
nand U3246 (N_3246,N_2721,N_2986);
nand U3247 (N_3247,N_2884,N_2639);
or U3248 (N_3248,N_3057,N_2941);
and U3249 (N_3249,N_2782,N_2575);
nor U3250 (N_3250,N_2951,N_2693);
and U3251 (N_3251,N_2750,N_2762);
and U3252 (N_3252,N_2837,N_2712);
nor U3253 (N_3253,N_3012,N_2589);
nand U3254 (N_3254,N_3096,N_3009);
nor U3255 (N_3255,N_2500,N_3061);
and U3256 (N_3256,N_2778,N_2554);
and U3257 (N_3257,N_2529,N_3053);
and U3258 (N_3258,N_3044,N_2631);
or U3259 (N_3259,N_2594,N_2822);
nand U3260 (N_3260,N_2917,N_2715);
nor U3261 (N_3261,N_2634,N_3033);
nand U3262 (N_3262,N_3102,N_2795);
and U3263 (N_3263,N_2780,N_2545);
or U3264 (N_3264,N_2899,N_2988);
and U3265 (N_3265,N_2786,N_2878);
and U3266 (N_3266,N_2716,N_3028);
and U3267 (N_3267,N_3078,N_2663);
nor U3268 (N_3268,N_2994,N_2679);
and U3269 (N_3269,N_2677,N_2555);
xnor U3270 (N_3270,N_2796,N_2976);
and U3271 (N_3271,N_2618,N_2896);
nor U3272 (N_3272,N_2946,N_3060);
and U3273 (N_3273,N_2898,N_2739);
nand U3274 (N_3274,N_2904,N_2673);
and U3275 (N_3275,N_2765,N_3072);
nor U3276 (N_3276,N_2758,N_2506);
and U3277 (N_3277,N_2510,N_2520);
nand U3278 (N_3278,N_2914,N_2858);
and U3279 (N_3279,N_2543,N_3086);
nand U3280 (N_3280,N_2562,N_2724);
or U3281 (N_3281,N_3042,N_3079);
or U3282 (N_3282,N_2703,N_2910);
nor U3283 (N_3283,N_2725,N_2707);
nand U3284 (N_3284,N_3105,N_3004);
and U3285 (N_3285,N_2530,N_2532);
or U3286 (N_3286,N_2623,N_2990);
nand U3287 (N_3287,N_2576,N_2993);
nor U3288 (N_3288,N_2735,N_2727);
nand U3289 (N_3289,N_2820,N_2794);
or U3290 (N_3290,N_2943,N_2757);
or U3291 (N_3291,N_2528,N_2678);
nor U3292 (N_3292,N_2548,N_2643);
xnor U3293 (N_3293,N_2621,N_3077);
nand U3294 (N_3294,N_2870,N_2645);
nand U3295 (N_3295,N_2838,N_3001);
nand U3296 (N_3296,N_2869,N_2874);
nand U3297 (N_3297,N_2790,N_2733);
or U3298 (N_3298,N_2895,N_3082);
nor U3299 (N_3299,N_2574,N_2930);
and U3300 (N_3300,N_2563,N_2764);
and U3301 (N_3301,N_2894,N_2915);
nand U3302 (N_3302,N_2863,N_2921);
and U3303 (N_3303,N_3123,N_2776);
nor U3304 (N_3304,N_2977,N_2605);
and U3305 (N_3305,N_2734,N_3024);
nor U3306 (N_3306,N_2912,N_2592);
nand U3307 (N_3307,N_2929,N_2507);
or U3308 (N_3308,N_3064,N_2695);
nor U3309 (N_3309,N_3002,N_2783);
and U3310 (N_3310,N_2861,N_2549);
and U3311 (N_3311,N_2606,N_2981);
xor U3312 (N_3312,N_2924,N_2646);
nor U3313 (N_3313,N_2686,N_2997);
and U3314 (N_3314,N_2654,N_2900);
or U3315 (N_3315,N_2933,N_2661);
xor U3316 (N_3316,N_2853,N_2664);
nand U3317 (N_3317,N_2801,N_3101);
and U3318 (N_3318,N_3038,N_3113);
and U3319 (N_3319,N_3110,N_2604);
xnor U3320 (N_3320,N_2905,N_3111);
or U3321 (N_3321,N_3041,N_2965);
and U3322 (N_3322,N_2855,N_2702);
or U3323 (N_3323,N_2599,N_3056);
nand U3324 (N_3324,N_2652,N_2969);
nor U3325 (N_3325,N_2726,N_2777);
and U3326 (N_3326,N_2642,N_2655);
nand U3327 (N_3327,N_2539,N_2751);
xnor U3328 (N_3328,N_2926,N_2955);
nor U3329 (N_3329,N_2799,N_2888);
nand U3330 (N_3330,N_2940,N_2967);
or U3331 (N_3331,N_3119,N_3073);
xor U3332 (N_3332,N_2824,N_2923);
and U3333 (N_3333,N_2709,N_3023);
nor U3334 (N_3334,N_2843,N_2701);
nor U3335 (N_3335,N_2632,N_2987);
and U3336 (N_3336,N_2688,N_3098);
or U3337 (N_3337,N_2760,N_2974);
nand U3338 (N_3338,N_2763,N_3067);
or U3339 (N_3339,N_2509,N_2834);
nor U3340 (N_3340,N_2522,N_2913);
nor U3341 (N_3341,N_2603,N_2515);
and U3342 (N_3342,N_2828,N_2806);
xor U3343 (N_3343,N_2736,N_2847);
nor U3344 (N_3344,N_2572,N_2852);
and U3345 (N_3345,N_3085,N_2881);
xor U3346 (N_3346,N_2694,N_2769);
nand U3347 (N_3347,N_2731,N_2860);
nand U3348 (N_3348,N_2637,N_2671);
and U3349 (N_3349,N_2519,N_3047);
nor U3350 (N_3350,N_3109,N_2985);
and U3351 (N_3351,N_2738,N_2740);
nor U3352 (N_3352,N_2937,N_2607);
nand U3353 (N_3353,N_2803,N_2787);
nor U3354 (N_3354,N_3088,N_2535);
xor U3355 (N_3355,N_2541,N_2544);
and U3356 (N_3356,N_2938,N_3122);
or U3357 (N_3357,N_2791,N_3051);
nor U3358 (N_3358,N_3118,N_2508);
nand U3359 (N_3359,N_2982,N_3063);
nor U3360 (N_3360,N_3043,N_2907);
nand U3361 (N_3361,N_2857,N_2672);
and U3362 (N_3362,N_2540,N_2676);
nand U3363 (N_3363,N_2615,N_2859);
nor U3364 (N_3364,N_2659,N_2754);
or U3365 (N_3365,N_3018,N_2961);
nand U3366 (N_3366,N_2810,N_3116);
or U3367 (N_3367,N_2826,N_3000);
or U3368 (N_3368,N_3068,N_2649);
and U3369 (N_3369,N_3084,N_2713);
and U3370 (N_3370,N_2952,N_2588);
nand U3371 (N_3371,N_3070,N_2568);
and U3372 (N_3372,N_2501,N_2569);
nor U3373 (N_3373,N_2848,N_2580);
nor U3374 (N_3374,N_3011,N_2805);
xnor U3375 (N_3375,N_2546,N_2690);
xor U3376 (N_3376,N_2784,N_2550);
and U3377 (N_3377,N_3107,N_2674);
nand U3378 (N_3378,N_2650,N_2975);
nand U3379 (N_3379,N_3097,N_2901);
xnor U3380 (N_3380,N_2578,N_3117);
or U3381 (N_3381,N_2902,N_2812);
nor U3382 (N_3382,N_2891,N_2670);
nor U3383 (N_3383,N_2611,N_2789);
nor U3384 (N_3384,N_2537,N_2779);
nand U3385 (N_3385,N_2602,N_2696);
nor U3386 (N_3386,N_2768,N_2609);
nand U3387 (N_3387,N_2538,N_2964);
nor U3388 (N_3388,N_2689,N_2567);
nand U3389 (N_3389,N_2831,N_2752);
nor U3390 (N_3390,N_3049,N_2816);
xnor U3391 (N_3391,N_2612,N_2916);
nand U3392 (N_3392,N_2761,N_2581);
nand U3393 (N_3393,N_2742,N_3124);
nand U3394 (N_3394,N_2879,N_3089);
or U3395 (N_3395,N_2710,N_2737);
xor U3396 (N_3396,N_2755,N_2512);
and U3397 (N_3397,N_3114,N_2759);
and U3398 (N_3398,N_3121,N_3054);
nand U3399 (N_3399,N_2628,N_2524);
nor U3400 (N_3400,N_2996,N_2968);
and U3401 (N_3401,N_3013,N_3075);
nand U3402 (N_3402,N_2610,N_2595);
or U3403 (N_3403,N_3010,N_2651);
nor U3404 (N_3404,N_2753,N_3120);
nand U3405 (N_3405,N_2959,N_3103);
nor U3406 (N_3406,N_2571,N_2947);
nand U3407 (N_3407,N_2518,N_2942);
or U3408 (N_3408,N_2616,N_2502);
xnor U3409 (N_3409,N_2608,N_2622);
nand U3410 (N_3410,N_3034,N_2720);
and U3411 (N_3411,N_2880,N_2704);
and U3412 (N_3412,N_2829,N_2842);
nor U3413 (N_3413,N_2918,N_2748);
nor U3414 (N_3414,N_2844,N_2566);
nand U3415 (N_3415,N_2617,N_2730);
nor U3416 (N_3416,N_2851,N_2925);
and U3417 (N_3417,N_3100,N_2708);
nand U3418 (N_3418,N_3030,N_2573);
and U3419 (N_3419,N_2892,N_2875);
or U3420 (N_3420,N_2647,N_2640);
and U3421 (N_3421,N_2788,N_2665);
and U3422 (N_3422,N_2558,N_3093);
nand U3423 (N_3423,N_2635,N_2909);
and U3424 (N_3424,N_2653,N_3016);
or U3425 (N_3425,N_2553,N_2991);
nand U3426 (N_3426,N_2700,N_3006);
xnor U3427 (N_3427,N_2854,N_2597);
or U3428 (N_3428,N_3106,N_2756);
or U3429 (N_3429,N_3037,N_3025);
nor U3430 (N_3430,N_2833,N_3003);
nand U3431 (N_3431,N_2699,N_3019);
nor U3432 (N_3432,N_2633,N_2808);
nor U3433 (N_3433,N_2692,N_3014);
and U3434 (N_3434,N_2886,N_3095);
and U3435 (N_3435,N_2800,N_2999);
and U3436 (N_3436,N_3083,N_2845);
or U3437 (N_3437,N_2684,N_2542);
and U3438 (N_3438,N_2958,N_2592);
and U3439 (N_3439,N_2999,N_2798);
nor U3440 (N_3440,N_3005,N_2687);
nor U3441 (N_3441,N_2635,N_2640);
nor U3442 (N_3442,N_2595,N_2856);
xor U3443 (N_3443,N_2728,N_2960);
nor U3444 (N_3444,N_2903,N_2680);
and U3445 (N_3445,N_2728,N_2786);
or U3446 (N_3446,N_2634,N_2978);
nand U3447 (N_3447,N_3000,N_2691);
or U3448 (N_3448,N_2783,N_2612);
and U3449 (N_3449,N_2882,N_2660);
nor U3450 (N_3450,N_3035,N_2632);
and U3451 (N_3451,N_2725,N_2687);
and U3452 (N_3452,N_2815,N_2655);
nand U3453 (N_3453,N_2680,N_3012);
nor U3454 (N_3454,N_2673,N_3045);
or U3455 (N_3455,N_2688,N_3048);
or U3456 (N_3456,N_2516,N_2618);
nor U3457 (N_3457,N_2541,N_2860);
nand U3458 (N_3458,N_2697,N_2933);
nor U3459 (N_3459,N_2994,N_2968);
or U3460 (N_3460,N_2632,N_3084);
and U3461 (N_3461,N_2695,N_2512);
nand U3462 (N_3462,N_3099,N_2947);
xnor U3463 (N_3463,N_2740,N_2984);
nor U3464 (N_3464,N_2758,N_2890);
xnor U3465 (N_3465,N_2648,N_2665);
nor U3466 (N_3466,N_2908,N_2898);
and U3467 (N_3467,N_2905,N_2672);
nor U3468 (N_3468,N_2783,N_2908);
or U3469 (N_3469,N_2934,N_2532);
xnor U3470 (N_3470,N_3084,N_2594);
nand U3471 (N_3471,N_2794,N_2577);
or U3472 (N_3472,N_3113,N_2621);
nand U3473 (N_3473,N_2650,N_2679);
nor U3474 (N_3474,N_2527,N_2917);
or U3475 (N_3475,N_2543,N_2729);
or U3476 (N_3476,N_3082,N_2939);
xnor U3477 (N_3477,N_2678,N_2592);
nand U3478 (N_3478,N_3105,N_2535);
nand U3479 (N_3479,N_3067,N_3102);
or U3480 (N_3480,N_2863,N_2673);
nor U3481 (N_3481,N_2715,N_2846);
xnor U3482 (N_3482,N_2678,N_2682);
nor U3483 (N_3483,N_2509,N_2684);
nand U3484 (N_3484,N_2726,N_3071);
and U3485 (N_3485,N_3002,N_2938);
nor U3486 (N_3486,N_2893,N_2661);
xor U3487 (N_3487,N_2534,N_2639);
or U3488 (N_3488,N_2932,N_2500);
and U3489 (N_3489,N_3098,N_2818);
nand U3490 (N_3490,N_2861,N_3057);
xnor U3491 (N_3491,N_2720,N_3037);
or U3492 (N_3492,N_2714,N_2700);
nand U3493 (N_3493,N_3021,N_2709);
or U3494 (N_3494,N_2878,N_3104);
xor U3495 (N_3495,N_2890,N_3101);
and U3496 (N_3496,N_2823,N_2672);
nor U3497 (N_3497,N_3078,N_2785);
and U3498 (N_3498,N_2508,N_2540);
xor U3499 (N_3499,N_2843,N_2593);
and U3500 (N_3500,N_3049,N_2986);
and U3501 (N_3501,N_2951,N_3052);
and U3502 (N_3502,N_2913,N_2759);
and U3503 (N_3503,N_2802,N_2708);
nor U3504 (N_3504,N_2631,N_2882);
nand U3505 (N_3505,N_2819,N_2959);
or U3506 (N_3506,N_3062,N_2718);
nand U3507 (N_3507,N_2758,N_2622);
nor U3508 (N_3508,N_2906,N_2736);
or U3509 (N_3509,N_2923,N_2723);
or U3510 (N_3510,N_3110,N_2724);
and U3511 (N_3511,N_3123,N_3117);
nor U3512 (N_3512,N_2643,N_3072);
nor U3513 (N_3513,N_2893,N_2599);
nor U3514 (N_3514,N_2879,N_2701);
nand U3515 (N_3515,N_3093,N_2523);
or U3516 (N_3516,N_2901,N_3017);
or U3517 (N_3517,N_2879,N_3124);
nor U3518 (N_3518,N_2667,N_2643);
or U3519 (N_3519,N_2689,N_2826);
nand U3520 (N_3520,N_2951,N_3039);
nor U3521 (N_3521,N_2865,N_3090);
or U3522 (N_3522,N_2963,N_2595);
or U3523 (N_3523,N_2555,N_2986);
nor U3524 (N_3524,N_2732,N_2889);
or U3525 (N_3525,N_2996,N_2995);
nand U3526 (N_3526,N_3124,N_2554);
and U3527 (N_3527,N_3059,N_3103);
or U3528 (N_3528,N_2796,N_2727);
nand U3529 (N_3529,N_2690,N_3006);
or U3530 (N_3530,N_3016,N_2914);
nor U3531 (N_3531,N_2610,N_2623);
nor U3532 (N_3532,N_2612,N_2961);
nand U3533 (N_3533,N_2957,N_2591);
and U3534 (N_3534,N_3060,N_2859);
xor U3535 (N_3535,N_2954,N_2845);
nor U3536 (N_3536,N_2631,N_2723);
nor U3537 (N_3537,N_2984,N_2860);
nand U3538 (N_3538,N_2503,N_3038);
nand U3539 (N_3539,N_2548,N_2513);
xor U3540 (N_3540,N_2942,N_2794);
xor U3541 (N_3541,N_2641,N_2977);
and U3542 (N_3542,N_2784,N_2534);
nand U3543 (N_3543,N_2840,N_2867);
and U3544 (N_3544,N_2755,N_2922);
and U3545 (N_3545,N_2687,N_2544);
xnor U3546 (N_3546,N_2677,N_2865);
or U3547 (N_3547,N_2729,N_3097);
nor U3548 (N_3548,N_2625,N_2609);
nand U3549 (N_3549,N_2863,N_2851);
and U3550 (N_3550,N_2992,N_3002);
nor U3551 (N_3551,N_2833,N_2649);
xnor U3552 (N_3552,N_3043,N_2596);
and U3553 (N_3553,N_2592,N_2846);
nor U3554 (N_3554,N_2793,N_2765);
nand U3555 (N_3555,N_2602,N_2844);
nand U3556 (N_3556,N_2938,N_2576);
nor U3557 (N_3557,N_2908,N_2568);
and U3558 (N_3558,N_2536,N_3092);
or U3559 (N_3559,N_2527,N_2945);
xor U3560 (N_3560,N_2796,N_2540);
and U3561 (N_3561,N_2539,N_2502);
or U3562 (N_3562,N_2504,N_2799);
nand U3563 (N_3563,N_2911,N_2688);
xor U3564 (N_3564,N_2693,N_2750);
or U3565 (N_3565,N_2618,N_2579);
xnor U3566 (N_3566,N_2830,N_2615);
nor U3567 (N_3567,N_2864,N_2972);
or U3568 (N_3568,N_3077,N_2797);
or U3569 (N_3569,N_3086,N_2938);
and U3570 (N_3570,N_2540,N_2615);
or U3571 (N_3571,N_2533,N_2645);
nor U3572 (N_3572,N_2535,N_2907);
nor U3573 (N_3573,N_3052,N_2955);
xor U3574 (N_3574,N_2836,N_3102);
nor U3575 (N_3575,N_2770,N_2768);
nor U3576 (N_3576,N_2823,N_2813);
nand U3577 (N_3577,N_2915,N_2935);
xnor U3578 (N_3578,N_2785,N_2710);
and U3579 (N_3579,N_2551,N_2604);
and U3580 (N_3580,N_2948,N_3064);
or U3581 (N_3581,N_2770,N_2866);
nand U3582 (N_3582,N_2698,N_3003);
or U3583 (N_3583,N_2748,N_2871);
nand U3584 (N_3584,N_2982,N_2658);
xnor U3585 (N_3585,N_2811,N_2716);
nand U3586 (N_3586,N_2881,N_2911);
and U3587 (N_3587,N_2601,N_2557);
and U3588 (N_3588,N_2985,N_3053);
or U3589 (N_3589,N_3006,N_2641);
or U3590 (N_3590,N_2891,N_2884);
nor U3591 (N_3591,N_2766,N_2714);
nor U3592 (N_3592,N_3016,N_2584);
nor U3593 (N_3593,N_2932,N_3109);
xor U3594 (N_3594,N_2805,N_2631);
or U3595 (N_3595,N_2508,N_2520);
and U3596 (N_3596,N_2504,N_2903);
nand U3597 (N_3597,N_2855,N_2835);
xor U3598 (N_3598,N_2530,N_2854);
or U3599 (N_3599,N_2799,N_2964);
or U3600 (N_3600,N_3111,N_2821);
nor U3601 (N_3601,N_2590,N_3007);
nand U3602 (N_3602,N_2770,N_2874);
nand U3603 (N_3603,N_2611,N_3040);
nor U3604 (N_3604,N_2541,N_2517);
nor U3605 (N_3605,N_2840,N_2745);
nor U3606 (N_3606,N_3014,N_2765);
or U3607 (N_3607,N_2784,N_2830);
or U3608 (N_3608,N_2981,N_2837);
xnor U3609 (N_3609,N_2715,N_2821);
or U3610 (N_3610,N_2570,N_2986);
nor U3611 (N_3611,N_2716,N_2819);
or U3612 (N_3612,N_2934,N_3066);
and U3613 (N_3613,N_2571,N_2522);
nand U3614 (N_3614,N_2873,N_3116);
nor U3615 (N_3615,N_2552,N_2933);
nand U3616 (N_3616,N_2603,N_3098);
xnor U3617 (N_3617,N_2824,N_2850);
xor U3618 (N_3618,N_3049,N_2765);
or U3619 (N_3619,N_2859,N_2845);
or U3620 (N_3620,N_3059,N_2502);
nor U3621 (N_3621,N_2509,N_2974);
nand U3622 (N_3622,N_2570,N_2883);
nand U3623 (N_3623,N_2875,N_2535);
nor U3624 (N_3624,N_2822,N_2649);
nand U3625 (N_3625,N_3117,N_2528);
nor U3626 (N_3626,N_2882,N_2934);
nor U3627 (N_3627,N_2768,N_3078);
nand U3628 (N_3628,N_2757,N_2603);
xor U3629 (N_3629,N_2690,N_2940);
xor U3630 (N_3630,N_2896,N_3072);
xnor U3631 (N_3631,N_2962,N_2915);
and U3632 (N_3632,N_3089,N_2868);
xor U3633 (N_3633,N_2827,N_2961);
nand U3634 (N_3634,N_2650,N_2754);
or U3635 (N_3635,N_2800,N_2749);
and U3636 (N_3636,N_2610,N_2570);
and U3637 (N_3637,N_2632,N_2594);
xnor U3638 (N_3638,N_2675,N_2925);
xor U3639 (N_3639,N_2925,N_2774);
xor U3640 (N_3640,N_2684,N_2585);
or U3641 (N_3641,N_2960,N_2981);
nor U3642 (N_3642,N_3073,N_3100);
and U3643 (N_3643,N_2956,N_2610);
or U3644 (N_3644,N_3015,N_2963);
and U3645 (N_3645,N_2670,N_3018);
or U3646 (N_3646,N_2714,N_2601);
and U3647 (N_3647,N_2911,N_2512);
nor U3648 (N_3648,N_2878,N_2830);
nor U3649 (N_3649,N_2770,N_2711);
or U3650 (N_3650,N_2910,N_2576);
or U3651 (N_3651,N_2798,N_2708);
nor U3652 (N_3652,N_3092,N_3034);
and U3653 (N_3653,N_2809,N_2907);
and U3654 (N_3654,N_2920,N_2734);
nor U3655 (N_3655,N_2869,N_2953);
and U3656 (N_3656,N_2949,N_2999);
nand U3657 (N_3657,N_2970,N_2538);
and U3658 (N_3658,N_2795,N_2985);
xnor U3659 (N_3659,N_2937,N_2864);
nor U3660 (N_3660,N_2784,N_2822);
nand U3661 (N_3661,N_2951,N_2737);
nor U3662 (N_3662,N_2617,N_2714);
nor U3663 (N_3663,N_2771,N_3071);
nand U3664 (N_3664,N_2818,N_2752);
or U3665 (N_3665,N_2946,N_3054);
nor U3666 (N_3666,N_2571,N_3067);
nand U3667 (N_3667,N_2786,N_3009);
or U3668 (N_3668,N_2964,N_2522);
nor U3669 (N_3669,N_3108,N_2986);
and U3670 (N_3670,N_2631,N_2643);
nor U3671 (N_3671,N_2703,N_2955);
and U3672 (N_3672,N_2607,N_2951);
nand U3673 (N_3673,N_2770,N_2719);
nor U3674 (N_3674,N_2576,N_2617);
and U3675 (N_3675,N_2503,N_2727);
nor U3676 (N_3676,N_2513,N_3059);
and U3677 (N_3677,N_2592,N_3065);
or U3678 (N_3678,N_2502,N_2601);
nand U3679 (N_3679,N_2675,N_2932);
nor U3680 (N_3680,N_2944,N_3069);
xor U3681 (N_3681,N_2615,N_2518);
nand U3682 (N_3682,N_3052,N_2944);
nor U3683 (N_3683,N_3068,N_2859);
and U3684 (N_3684,N_3124,N_2822);
nor U3685 (N_3685,N_2694,N_2711);
nand U3686 (N_3686,N_2959,N_2512);
xor U3687 (N_3687,N_2937,N_3087);
and U3688 (N_3688,N_2627,N_2532);
or U3689 (N_3689,N_2572,N_3087);
nor U3690 (N_3690,N_2949,N_2858);
xor U3691 (N_3691,N_2802,N_2527);
or U3692 (N_3692,N_2796,N_2827);
nor U3693 (N_3693,N_2964,N_2656);
and U3694 (N_3694,N_2851,N_2993);
or U3695 (N_3695,N_2663,N_3073);
nor U3696 (N_3696,N_3073,N_2995);
nor U3697 (N_3697,N_2845,N_3123);
and U3698 (N_3698,N_2723,N_2950);
or U3699 (N_3699,N_2851,N_2935);
and U3700 (N_3700,N_2694,N_3067);
nor U3701 (N_3701,N_2555,N_3006);
nand U3702 (N_3702,N_2605,N_2786);
nor U3703 (N_3703,N_2597,N_2939);
xor U3704 (N_3704,N_3018,N_2986);
xnor U3705 (N_3705,N_2723,N_2909);
and U3706 (N_3706,N_2817,N_2563);
nand U3707 (N_3707,N_2815,N_2879);
and U3708 (N_3708,N_3093,N_2996);
nand U3709 (N_3709,N_2860,N_2700);
and U3710 (N_3710,N_2814,N_2689);
nand U3711 (N_3711,N_2935,N_2622);
and U3712 (N_3712,N_3055,N_2961);
nand U3713 (N_3713,N_2971,N_2899);
and U3714 (N_3714,N_2676,N_2501);
or U3715 (N_3715,N_3015,N_2782);
or U3716 (N_3716,N_3091,N_2783);
and U3717 (N_3717,N_2602,N_2574);
or U3718 (N_3718,N_2739,N_2747);
or U3719 (N_3719,N_2663,N_2992);
nor U3720 (N_3720,N_2753,N_2814);
or U3721 (N_3721,N_2585,N_2866);
and U3722 (N_3722,N_2655,N_2631);
nand U3723 (N_3723,N_3054,N_2937);
nor U3724 (N_3724,N_2925,N_2523);
and U3725 (N_3725,N_2901,N_3089);
and U3726 (N_3726,N_2614,N_2994);
nand U3727 (N_3727,N_2997,N_2642);
nor U3728 (N_3728,N_2790,N_3017);
or U3729 (N_3729,N_2524,N_2533);
or U3730 (N_3730,N_3082,N_2637);
and U3731 (N_3731,N_3107,N_3108);
or U3732 (N_3732,N_3119,N_2975);
nor U3733 (N_3733,N_2950,N_2870);
nand U3734 (N_3734,N_2662,N_2889);
or U3735 (N_3735,N_2583,N_3094);
nor U3736 (N_3736,N_2528,N_2516);
nand U3737 (N_3737,N_2868,N_2965);
or U3738 (N_3738,N_2592,N_3048);
and U3739 (N_3739,N_2705,N_3077);
and U3740 (N_3740,N_3048,N_3071);
or U3741 (N_3741,N_3075,N_2633);
and U3742 (N_3742,N_3007,N_3051);
xor U3743 (N_3743,N_2852,N_2859);
nor U3744 (N_3744,N_2587,N_2833);
or U3745 (N_3745,N_2643,N_2677);
nor U3746 (N_3746,N_2999,N_2672);
nand U3747 (N_3747,N_2937,N_3016);
nor U3748 (N_3748,N_2780,N_2775);
nand U3749 (N_3749,N_2858,N_2787);
xor U3750 (N_3750,N_3283,N_3143);
or U3751 (N_3751,N_3170,N_3403);
and U3752 (N_3752,N_3568,N_3745);
xor U3753 (N_3753,N_3446,N_3247);
and U3754 (N_3754,N_3650,N_3214);
nand U3755 (N_3755,N_3460,N_3240);
nor U3756 (N_3756,N_3663,N_3677);
or U3757 (N_3757,N_3497,N_3200);
or U3758 (N_3758,N_3342,N_3252);
or U3759 (N_3759,N_3358,N_3661);
and U3760 (N_3760,N_3351,N_3380);
and U3761 (N_3761,N_3538,N_3296);
nand U3762 (N_3762,N_3306,N_3632);
or U3763 (N_3763,N_3537,N_3581);
xor U3764 (N_3764,N_3712,N_3494);
and U3765 (N_3765,N_3267,N_3203);
nor U3766 (N_3766,N_3589,N_3634);
xor U3767 (N_3767,N_3515,N_3559);
and U3768 (N_3768,N_3223,N_3280);
and U3769 (N_3769,N_3672,N_3207);
nand U3770 (N_3770,N_3630,N_3268);
nand U3771 (N_3771,N_3396,N_3449);
nand U3772 (N_3772,N_3593,N_3536);
nor U3773 (N_3773,N_3738,N_3313);
nor U3774 (N_3774,N_3250,N_3474);
and U3775 (N_3775,N_3441,N_3276);
nand U3776 (N_3776,N_3714,N_3558);
nand U3777 (N_3777,N_3179,N_3389);
nor U3778 (N_3778,N_3722,N_3418);
nor U3779 (N_3779,N_3264,N_3144);
or U3780 (N_3780,N_3597,N_3163);
nand U3781 (N_3781,N_3547,N_3324);
or U3782 (N_3782,N_3660,N_3680);
nand U3783 (N_3783,N_3265,N_3141);
nor U3784 (N_3784,N_3669,N_3426);
or U3785 (N_3785,N_3376,N_3488);
or U3786 (N_3786,N_3374,N_3657);
nand U3787 (N_3787,N_3739,N_3244);
or U3788 (N_3788,N_3472,N_3257);
nor U3789 (N_3789,N_3347,N_3431);
nor U3790 (N_3790,N_3225,N_3178);
or U3791 (N_3791,N_3604,N_3620);
nand U3792 (N_3792,N_3687,N_3564);
nor U3793 (N_3793,N_3540,N_3370);
nor U3794 (N_3794,N_3133,N_3691);
and U3795 (N_3795,N_3567,N_3174);
or U3796 (N_3796,N_3471,N_3666);
nand U3797 (N_3797,N_3219,N_3607);
and U3798 (N_3798,N_3198,N_3671);
nand U3799 (N_3799,N_3400,N_3408);
nand U3800 (N_3800,N_3550,N_3676);
nand U3801 (N_3801,N_3655,N_3224);
nor U3802 (N_3802,N_3470,N_3734);
nor U3803 (N_3803,N_3182,N_3624);
or U3804 (N_3804,N_3573,N_3667);
nand U3805 (N_3805,N_3373,N_3490);
or U3806 (N_3806,N_3165,N_3175);
or U3807 (N_3807,N_3628,N_3654);
xnor U3808 (N_3808,N_3381,N_3333);
nor U3809 (N_3809,N_3161,N_3384);
nor U3810 (N_3810,N_3433,N_3292);
or U3811 (N_3811,N_3332,N_3402);
nand U3812 (N_3812,N_3357,N_3631);
and U3813 (N_3813,N_3241,N_3259);
nand U3814 (N_3814,N_3355,N_3210);
nor U3815 (N_3815,N_3432,N_3295);
nor U3816 (N_3816,N_3235,N_3563);
or U3817 (N_3817,N_3234,N_3453);
and U3818 (N_3818,N_3438,N_3718);
and U3819 (N_3819,N_3246,N_3371);
and U3820 (N_3820,N_3270,N_3506);
nor U3821 (N_3821,N_3489,N_3614);
nor U3822 (N_3822,N_3397,N_3545);
or U3823 (N_3823,N_3321,N_3509);
nand U3824 (N_3824,N_3145,N_3549);
xor U3825 (N_3825,N_3623,N_3640);
nand U3826 (N_3826,N_3528,N_3361);
or U3827 (N_3827,N_3555,N_3566);
xnor U3828 (N_3828,N_3478,N_3125);
or U3829 (N_3829,N_3137,N_3637);
and U3830 (N_3830,N_3605,N_3378);
or U3831 (N_3831,N_3211,N_3166);
nor U3832 (N_3832,N_3706,N_3359);
xnor U3833 (N_3833,N_3372,N_3414);
or U3834 (N_3834,N_3421,N_3386);
or U3835 (N_3835,N_3723,N_3363);
or U3836 (N_3836,N_3304,N_3735);
or U3837 (N_3837,N_3301,N_3647);
and U3838 (N_3838,N_3642,N_3636);
and U3839 (N_3839,N_3254,N_3443);
nor U3840 (N_3840,N_3749,N_3275);
nand U3841 (N_3841,N_3613,N_3391);
xnor U3842 (N_3842,N_3557,N_3688);
and U3843 (N_3843,N_3656,N_3300);
nor U3844 (N_3844,N_3422,N_3277);
and U3845 (N_3845,N_3130,N_3533);
or U3846 (N_3846,N_3317,N_3187);
and U3847 (N_3847,N_3196,N_3274);
or U3848 (N_3848,N_3698,N_3456);
nand U3849 (N_3849,N_3588,N_3571);
xor U3850 (N_3850,N_3181,N_3385);
or U3851 (N_3851,N_3354,N_3286);
nand U3852 (N_3852,N_3584,N_3401);
and U3853 (N_3853,N_3675,N_3451);
and U3854 (N_3854,N_3448,N_3658);
or U3855 (N_3855,N_3684,N_3504);
nand U3856 (N_3856,N_3341,N_3694);
nor U3857 (N_3857,N_3279,N_3208);
nand U3858 (N_3858,N_3233,N_3319);
or U3859 (N_3859,N_3612,N_3475);
and U3860 (N_3860,N_3193,N_3410);
xor U3861 (N_3861,N_3330,N_3331);
nor U3862 (N_3862,N_3560,N_3340);
xnor U3863 (N_3863,N_3158,N_3516);
or U3864 (N_3864,N_3747,N_3173);
and U3865 (N_3865,N_3491,N_3189);
xor U3866 (N_3866,N_3399,N_3499);
and U3867 (N_3867,N_3700,N_3442);
and U3868 (N_3868,N_3154,N_3350);
nand U3869 (N_3869,N_3670,N_3258);
or U3870 (N_3870,N_3205,N_3465);
nand U3871 (N_3871,N_3217,N_3595);
and U3872 (N_3872,N_3546,N_3379);
and U3873 (N_3873,N_3334,N_3269);
or U3874 (N_3874,N_3689,N_3646);
nor U3875 (N_3875,N_3171,N_3483);
or U3876 (N_3876,N_3622,N_3216);
nor U3877 (N_3877,N_3713,N_3282);
nand U3878 (N_3878,N_3220,N_3464);
nand U3879 (N_3879,N_3338,N_3525);
nand U3880 (N_3880,N_3693,N_3575);
and U3881 (N_3881,N_3228,N_3232);
xnor U3882 (N_3882,N_3727,N_3479);
nand U3883 (N_3883,N_3619,N_3725);
nand U3884 (N_3884,N_3266,N_3195);
and U3885 (N_3885,N_3678,N_3184);
nand U3886 (N_3886,N_3352,N_3616);
nor U3887 (N_3887,N_3502,N_3554);
nor U3888 (N_3888,N_3172,N_3327);
or U3889 (N_3889,N_3387,N_3551);
nor U3890 (N_3890,N_3569,N_3503);
nor U3891 (N_3891,N_3263,N_3190);
nand U3892 (N_3892,N_3493,N_3531);
xor U3893 (N_3893,N_3262,N_3281);
xnor U3894 (N_3894,N_3512,N_3454);
xor U3895 (N_3895,N_3461,N_3218);
nand U3896 (N_3896,N_3285,N_3467);
and U3897 (N_3897,N_3416,N_3136);
or U3898 (N_3898,N_3458,N_3377);
or U3899 (N_3899,N_3312,N_3645);
or U3900 (N_3900,N_3445,N_3322);
nand U3901 (N_3901,N_3603,N_3339);
or U3902 (N_3902,N_3151,N_3229);
nor U3903 (N_3903,N_3699,N_3621);
nor U3904 (N_3904,N_3447,N_3673);
and U3905 (N_3905,N_3626,N_3519);
or U3906 (N_3906,N_3583,N_3495);
and U3907 (N_3907,N_3591,N_3393);
and U3908 (N_3908,N_3231,N_3682);
nand U3909 (N_3909,N_3197,N_3430);
nand U3910 (N_3910,N_3695,N_3487);
xnor U3911 (N_3911,N_3409,N_3518);
nor U3912 (N_3912,N_3226,N_3659);
and U3913 (N_3913,N_3526,N_3424);
xnor U3914 (N_3914,N_3419,N_3315);
and U3915 (N_3915,N_3169,N_3138);
nor U3916 (N_3916,N_3344,N_3153);
or U3917 (N_3917,N_3638,N_3237);
or U3918 (N_3918,N_3382,N_3587);
or U3919 (N_3919,N_3142,N_3548);
nand U3920 (N_3920,N_3362,N_3599);
xnor U3921 (N_3921,N_3434,N_3383);
nor U3922 (N_3922,N_3481,N_3552);
nor U3923 (N_3923,N_3251,N_3227);
or U3924 (N_3924,N_3177,N_3681);
nand U3925 (N_3925,N_3425,N_3696);
or U3926 (N_3926,N_3248,N_3649);
nand U3927 (N_3927,N_3744,N_3711);
and U3928 (N_3928,N_3462,N_3641);
xnor U3929 (N_3929,N_3505,N_3520);
or U3930 (N_3930,N_3420,N_3395);
and U3931 (N_3931,N_3202,N_3590);
or U3932 (N_3932,N_3349,N_3578);
and U3933 (N_3933,N_3375,N_3323);
nand U3934 (N_3934,N_3238,N_3466);
or U3935 (N_3935,N_3415,N_3436);
xnor U3936 (N_3936,N_3602,N_3743);
nand U3937 (N_3937,N_3293,N_3577);
xor U3938 (N_3938,N_3328,N_3716);
nor U3939 (N_3939,N_3608,N_3477);
nor U3940 (N_3940,N_3261,N_3260);
nor U3941 (N_3941,N_3299,N_3392);
xnor U3942 (N_3942,N_3343,N_3288);
nand U3943 (N_3943,N_3535,N_3435);
nand U3944 (N_3944,N_3160,N_3291);
nor U3945 (N_3945,N_3707,N_3708);
nand U3946 (N_3946,N_3302,N_3521);
or U3947 (N_3947,N_3580,N_3606);
or U3948 (N_3948,N_3287,N_3201);
nand U3949 (N_3949,N_3309,N_3176);
or U3950 (N_3950,N_3423,N_3586);
nand U3951 (N_3951,N_3709,N_3553);
or U3952 (N_3952,N_3484,N_3417);
or U3953 (N_3953,N_3147,N_3311);
and U3954 (N_3954,N_3480,N_3272);
or U3955 (N_3955,N_3501,N_3162);
nor U3956 (N_3956,N_3702,N_3188);
nor U3957 (N_3957,N_3368,N_3457);
and U3958 (N_3958,N_3513,N_3212);
and U3959 (N_3959,N_3611,N_3733);
and U3960 (N_3960,N_3307,N_3496);
and U3961 (N_3961,N_3326,N_3157);
nand U3962 (N_3962,N_3721,N_3284);
nor U3963 (N_3963,N_3668,N_3394);
nand U3964 (N_3964,N_3742,N_3440);
nand U3965 (N_3965,N_3697,N_3191);
or U3966 (N_3966,N_3705,N_3428);
or U3967 (N_3967,N_3625,N_3412);
nor U3968 (N_3968,N_3570,N_3128);
nor U3969 (N_3969,N_3701,N_3180);
nor U3970 (N_3970,N_3256,N_3305);
or U3971 (N_3971,N_3651,N_3134);
nand U3972 (N_3972,N_3192,N_3730);
nor U3973 (N_3973,N_3167,N_3482);
nand U3974 (N_3974,N_3664,N_3164);
or U3975 (N_3975,N_3325,N_3146);
xnor U3976 (N_3976,N_3574,N_3690);
or U3977 (N_3977,N_3345,N_3596);
nand U3978 (N_3978,N_3140,N_3455);
and U3979 (N_3979,N_3542,N_3585);
or U3980 (N_3980,N_3129,N_3253);
nand U3981 (N_3981,N_3522,N_3517);
and U3982 (N_3982,N_3437,N_3726);
nand U3983 (N_3983,N_3429,N_3439);
and U3984 (N_3984,N_3565,N_3230);
and U3985 (N_3985,N_3469,N_3610);
xor U3986 (N_3986,N_3168,N_3485);
nor U3987 (N_3987,N_3314,N_3127);
or U3988 (N_3988,N_3534,N_3703);
nor U3989 (N_3989,N_3511,N_3139);
and U3990 (N_3990,N_3633,N_3662);
or U3991 (N_3991,N_3746,N_3308);
or U3992 (N_3992,N_3627,N_3486);
and U3993 (N_3993,N_3303,N_3492);
or U3994 (N_3994,N_3346,N_3529);
and U3995 (N_3995,N_3508,N_3720);
xor U3996 (N_3996,N_3572,N_3500);
and U3997 (N_3997,N_3463,N_3148);
nand U3998 (N_3998,N_3562,N_3388);
or U3999 (N_3999,N_3717,N_3704);
or U4000 (N_4000,N_3579,N_3273);
or U4001 (N_4001,N_3348,N_3728);
xor U4002 (N_4002,N_3427,N_3204);
xor U4003 (N_4003,N_3271,N_3601);
and U4004 (N_4004,N_3635,N_3249);
or U4005 (N_4005,N_3715,N_3729);
nor U4006 (N_4006,N_3209,N_3674);
nor U4007 (N_4007,N_3155,N_3406);
nor U4008 (N_4008,N_3543,N_3206);
nand U4009 (N_4009,N_3369,N_3740);
and U4010 (N_4010,N_3530,N_3365);
or U4011 (N_4011,N_3199,N_3131);
nand U4012 (N_4012,N_3452,N_3748);
and U4013 (N_4013,N_3390,N_3222);
or U4014 (N_4014,N_3644,N_3367);
xnor U4015 (N_4015,N_3298,N_3665);
xor U4016 (N_4016,N_3527,N_3598);
or U4017 (N_4017,N_3639,N_3404);
nor U4018 (N_4018,N_3413,N_3194);
and U4019 (N_4019,N_3236,N_3468);
nor U4020 (N_4020,N_3683,N_3242);
or U4021 (N_4021,N_3510,N_3159);
nor U4022 (N_4022,N_3523,N_3473);
nand U4023 (N_4023,N_3150,N_3356);
nand U4024 (N_4024,N_3736,N_3732);
and U4025 (N_4025,N_3360,N_3126);
and U4026 (N_4026,N_3329,N_3149);
and U4027 (N_4027,N_3459,N_3679);
xnor U4028 (N_4028,N_3450,N_3353);
or U4029 (N_4029,N_3411,N_3336);
or U4030 (N_4030,N_3255,N_3245);
and U4031 (N_4031,N_3183,N_3648);
nor U4032 (N_4032,N_3294,N_3539);
nand U4033 (N_4033,N_3710,N_3444);
nor U4034 (N_4034,N_3215,N_3507);
and U4035 (N_4035,N_3643,N_3582);
nor U4036 (N_4036,N_3615,N_3692);
nor U4037 (N_4037,N_3561,N_3310);
xnor U4038 (N_4038,N_3617,N_3186);
nor U4039 (N_4039,N_3407,N_3290);
nor U4040 (N_4040,N_3335,N_3318);
nor U4041 (N_4041,N_3316,N_3278);
nor U4042 (N_4042,N_3600,N_3724);
xnor U4043 (N_4043,N_3239,N_3686);
nor U4044 (N_4044,N_3576,N_3532);
or U4045 (N_4045,N_3132,N_3156);
nor U4046 (N_4046,N_3594,N_3243);
nand U4047 (N_4047,N_3366,N_3514);
or U4048 (N_4048,N_3320,N_3405);
or U4049 (N_4049,N_3398,N_3737);
or U4050 (N_4050,N_3364,N_3152);
and U4051 (N_4051,N_3731,N_3629);
and U4052 (N_4052,N_3337,N_3221);
nor U4053 (N_4053,N_3524,N_3618);
and U4054 (N_4054,N_3297,N_3289);
nor U4055 (N_4055,N_3719,N_3609);
or U4056 (N_4056,N_3741,N_3544);
or U4057 (N_4057,N_3685,N_3213);
nor U4058 (N_4058,N_3592,N_3135);
or U4059 (N_4059,N_3652,N_3556);
nor U4060 (N_4060,N_3476,N_3185);
or U4061 (N_4061,N_3498,N_3541);
or U4062 (N_4062,N_3653,N_3553);
or U4063 (N_4063,N_3451,N_3566);
nand U4064 (N_4064,N_3422,N_3408);
xnor U4065 (N_4065,N_3267,N_3346);
and U4066 (N_4066,N_3147,N_3396);
nand U4067 (N_4067,N_3563,N_3429);
or U4068 (N_4068,N_3567,N_3569);
nand U4069 (N_4069,N_3166,N_3629);
nand U4070 (N_4070,N_3145,N_3266);
xor U4071 (N_4071,N_3631,N_3330);
and U4072 (N_4072,N_3182,N_3579);
nor U4073 (N_4073,N_3282,N_3645);
nor U4074 (N_4074,N_3329,N_3319);
and U4075 (N_4075,N_3679,N_3162);
xor U4076 (N_4076,N_3658,N_3269);
nand U4077 (N_4077,N_3487,N_3238);
and U4078 (N_4078,N_3465,N_3728);
or U4079 (N_4079,N_3740,N_3401);
xnor U4080 (N_4080,N_3572,N_3725);
nor U4081 (N_4081,N_3370,N_3432);
nand U4082 (N_4082,N_3567,N_3690);
or U4083 (N_4083,N_3276,N_3449);
nand U4084 (N_4084,N_3634,N_3213);
xnor U4085 (N_4085,N_3473,N_3558);
nor U4086 (N_4086,N_3395,N_3245);
nor U4087 (N_4087,N_3501,N_3288);
nand U4088 (N_4088,N_3538,N_3244);
nand U4089 (N_4089,N_3448,N_3134);
nand U4090 (N_4090,N_3418,N_3480);
nand U4091 (N_4091,N_3293,N_3320);
or U4092 (N_4092,N_3524,N_3172);
nand U4093 (N_4093,N_3599,N_3460);
and U4094 (N_4094,N_3513,N_3204);
and U4095 (N_4095,N_3284,N_3321);
nor U4096 (N_4096,N_3612,N_3600);
nor U4097 (N_4097,N_3341,N_3265);
or U4098 (N_4098,N_3495,N_3357);
nor U4099 (N_4099,N_3285,N_3336);
and U4100 (N_4100,N_3660,N_3415);
nor U4101 (N_4101,N_3205,N_3472);
or U4102 (N_4102,N_3336,N_3480);
and U4103 (N_4103,N_3555,N_3511);
and U4104 (N_4104,N_3299,N_3728);
nand U4105 (N_4105,N_3599,N_3225);
or U4106 (N_4106,N_3448,N_3532);
and U4107 (N_4107,N_3224,N_3317);
or U4108 (N_4108,N_3647,N_3402);
nor U4109 (N_4109,N_3668,N_3488);
and U4110 (N_4110,N_3181,N_3417);
or U4111 (N_4111,N_3707,N_3525);
xor U4112 (N_4112,N_3384,N_3387);
or U4113 (N_4113,N_3532,N_3614);
xor U4114 (N_4114,N_3315,N_3529);
and U4115 (N_4115,N_3318,N_3248);
and U4116 (N_4116,N_3537,N_3549);
and U4117 (N_4117,N_3325,N_3742);
and U4118 (N_4118,N_3492,N_3547);
or U4119 (N_4119,N_3744,N_3423);
or U4120 (N_4120,N_3531,N_3623);
nor U4121 (N_4121,N_3515,N_3534);
nor U4122 (N_4122,N_3156,N_3417);
nor U4123 (N_4123,N_3237,N_3588);
nor U4124 (N_4124,N_3660,N_3639);
nand U4125 (N_4125,N_3438,N_3141);
xnor U4126 (N_4126,N_3451,N_3327);
xor U4127 (N_4127,N_3514,N_3722);
or U4128 (N_4128,N_3134,N_3420);
nand U4129 (N_4129,N_3451,N_3212);
or U4130 (N_4130,N_3138,N_3558);
nand U4131 (N_4131,N_3552,N_3644);
and U4132 (N_4132,N_3497,N_3150);
nand U4133 (N_4133,N_3574,N_3227);
and U4134 (N_4134,N_3300,N_3306);
or U4135 (N_4135,N_3335,N_3709);
nor U4136 (N_4136,N_3738,N_3650);
or U4137 (N_4137,N_3570,N_3406);
nand U4138 (N_4138,N_3572,N_3609);
or U4139 (N_4139,N_3680,N_3391);
or U4140 (N_4140,N_3265,N_3351);
nor U4141 (N_4141,N_3410,N_3411);
and U4142 (N_4142,N_3212,N_3491);
nor U4143 (N_4143,N_3399,N_3335);
nor U4144 (N_4144,N_3658,N_3444);
and U4145 (N_4145,N_3663,N_3285);
nor U4146 (N_4146,N_3558,N_3467);
xor U4147 (N_4147,N_3476,N_3408);
or U4148 (N_4148,N_3555,N_3706);
and U4149 (N_4149,N_3716,N_3513);
nor U4150 (N_4150,N_3414,N_3411);
nor U4151 (N_4151,N_3660,N_3265);
nand U4152 (N_4152,N_3534,N_3212);
or U4153 (N_4153,N_3537,N_3482);
or U4154 (N_4154,N_3432,N_3618);
xor U4155 (N_4155,N_3555,N_3441);
xnor U4156 (N_4156,N_3614,N_3583);
and U4157 (N_4157,N_3679,N_3705);
nor U4158 (N_4158,N_3537,N_3282);
nand U4159 (N_4159,N_3709,N_3700);
or U4160 (N_4160,N_3222,N_3545);
and U4161 (N_4161,N_3411,N_3708);
or U4162 (N_4162,N_3544,N_3730);
or U4163 (N_4163,N_3184,N_3478);
or U4164 (N_4164,N_3706,N_3526);
and U4165 (N_4165,N_3639,N_3429);
and U4166 (N_4166,N_3438,N_3379);
and U4167 (N_4167,N_3327,N_3233);
nor U4168 (N_4168,N_3745,N_3137);
xor U4169 (N_4169,N_3193,N_3407);
nand U4170 (N_4170,N_3171,N_3402);
nor U4171 (N_4171,N_3688,N_3577);
nand U4172 (N_4172,N_3141,N_3147);
nand U4173 (N_4173,N_3243,N_3540);
nor U4174 (N_4174,N_3240,N_3590);
nor U4175 (N_4175,N_3739,N_3274);
nor U4176 (N_4176,N_3210,N_3462);
or U4177 (N_4177,N_3605,N_3672);
or U4178 (N_4178,N_3487,N_3523);
nor U4179 (N_4179,N_3490,N_3224);
or U4180 (N_4180,N_3630,N_3688);
or U4181 (N_4181,N_3468,N_3366);
and U4182 (N_4182,N_3674,N_3660);
nor U4183 (N_4183,N_3739,N_3699);
and U4184 (N_4184,N_3748,N_3373);
and U4185 (N_4185,N_3729,N_3157);
xnor U4186 (N_4186,N_3335,N_3428);
nor U4187 (N_4187,N_3676,N_3582);
and U4188 (N_4188,N_3200,N_3259);
nand U4189 (N_4189,N_3440,N_3593);
nor U4190 (N_4190,N_3466,N_3465);
nor U4191 (N_4191,N_3312,N_3572);
xor U4192 (N_4192,N_3631,N_3730);
and U4193 (N_4193,N_3631,N_3283);
xor U4194 (N_4194,N_3327,N_3494);
nor U4195 (N_4195,N_3496,N_3484);
and U4196 (N_4196,N_3618,N_3641);
nor U4197 (N_4197,N_3659,N_3311);
or U4198 (N_4198,N_3622,N_3731);
and U4199 (N_4199,N_3138,N_3517);
or U4200 (N_4200,N_3730,N_3436);
nand U4201 (N_4201,N_3584,N_3206);
nor U4202 (N_4202,N_3288,N_3211);
nand U4203 (N_4203,N_3366,N_3631);
and U4204 (N_4204,N_3561,N_3206);
and U4205 (N_4205,N_3149,N_3309);
and U4206 (N_4206,N_3137,N_3452);
nand U4207 (N_4207,N_3354,N_3658);
nand U4208 (N_4208,N_3245,N_3136);
and U4209 (N_4209,N_3324,N_3182);
or U4210 (N_4210,N_3195,N_3650);
nor U4211 (N_4211,N_3327,N_3374);
or U4212 (N_4212,N_3132,N_3483);
nand U4213 (N_4213,N_3673,N_3625);
and U4214 (N_4214,N_3714,N_3236);
or U4215 (N_4215,N_3684,N_3607);
nand U4216 (N_4216,N_3647,N_3241);
or U4217 (N_4217,N_3255,N_3292);
xor U4218 (N_4218,N_3360,N_3530);
or U4219 (N_4219,N_3508,N_3619);
or U4220 (N_4220,N_3480,N_3146);
or U4221 (N_4221,N_3429,N_3300);
nor U4222 (N_4222,N_3329,N_3472);
nand U4223 (N_4223,N_3498,N_3170);
and U4224 (N_4224,N_3384,N_3143);
nor U4225 (N_4225,N_3578,N_3155);
xnor U4226 (N_4226,N_3729,N_3337);
xor U4227 (N_4227,N_3416,N_3599);
or U4228 (N_4228,N_3204,N_3289);
nand U4229 (N_4229,N_3404,N_3378);
nand U4230 (N_4230,N_3351,N_3149);
nor U4231 (N_4231,N_3176,N_3470);
or U4232 (N_4232,N_3473,N_3129);
and U4233 (N_4233,N_3487,N_3388);
nor U4234 (N_4234,N_3726,N_3349);
and U4235 (N_4235,N_3666,N_3449);
or U4236 (N_4236,N_3459,N_3599);
and U4237 (N_4237,N_3441,N_3376);
nand U4238 (N_4238,N_3711,N_3158);
and U4239 (N_4239,N_3432,N_3561);
and U4240 (N_4240,N_3700,N_3193);
or U4241 (N_4241,N_3231,N_3378);
nor U4242 (N_4242,N_3305,N_3523);
or U4243 (N_4243,N_3406,N_3500);
nand U4244 (N_4244,N_3238,N_3652);
or U4245 (N_4245,N_3321,N_3709);
and U4246 (N_4246,N_3636,N_3422);
nor U4247 (N_4247,N_3571,N_3297);
nand U4248 (N_4248,N_3397,N_3284);
nand U4249 (N_4249,N_3478,N_3452);
nor U4250 (N_4250,N_3493,N_3296);
xor U4251 (N_4251,N_3196,N_3388);
nand U4252 (N_4252,N_3253,N_3746);
or U4253 (N_4253,N_3402,N_3301);
nand U4254 (N_4254,N_3675,N_3432);
and U4255 (N_4255,N_3481,N_3673);
or U4256 (N_4256,N_3334,N_3306);
nand U4257 (N_4257,N_3283,N_3647);
or U4258 (N_4258,N_3570,N_3530);
or U4259 (N_4259,N_3701,N_3172);
nand U4260 (N_4260,N_3705,N_3230);
nand U4261 (N_4261,N_3367,N_3612);
nor U4262 (N_4262,N_3334,N_3148);
xor U4263 (N_4263,N_3459,N_3554);
and U4264 (N_4264,N_3738,N_3353);
nand U4265 (N_4265,N_3518,N_3261);
and U4266 (N_4266,N_3603,N_3168);
xnor U4267 (N_4267,N_3221,N_3479);
and U4268 (N_4268,N_3182,N_3172);
nand U4269 (N_4269,N_3676,N_3390);
or U4270 (N_4270,N_3217,N_3400);
or U4271 (N_4271,N_3226,N_3637);
nor U4272 (N_4272,N_3438,N_3706);
and U4273 (N_4273,N_3156,N_3264);
nor U4274 (N_4274,N_3716,N_3346);
and U4275 (N_4275,N_3372,N_3373);
or U4276 (N_4276,N_3591,N_3516);
or U4277 (N_4277,N_3509,N_3711);
or U4278 (N_4278,N_3446,N_3636);
or U4279 (N_4279,N_3149,N_3193);
nor U4280 (N_4280,N_3650,N_3372);
and U4281 (N_4281,N_3379,N_3139);
xor U4282 (N_4282,N_3295,N_3171);
nor U4283 (N_4283,N_3158,N_3339);
nor U4284 (N_4284,N_3435,N_3259);
nor U4285 (N_4285,N_3671,N_3293);
and U4286 (N_4286,N_3572,N_3686);
and U4287 (N_4287,N_3293,N_3668);
nor U4288 (N_4288,N_3688,N_3652);
xnor U4289 (N_4289,N_3513,N_3369);
nor U4290 (N_4290,N_3433,N_3377);
or U4291 (N_4291,N_3346,N_3232);
or U4292 (N_4292,N_3303,N_3178);
nor U4293 (N_4293,N_3220,N_3340);
nand U4294 (N_4294,N_3174,N_3314);
xnor U4295 (N_4295,N_3282,N_3735);
nand U4296 (N_4296,N_3183,N_3690);
xor U4297 (N_4297,N_3626,N_3237);
nand U4298 (N_4298,N_3335,N_3457);
or U4299 (N_4299,N_3735,N_3513);
and U4300 (N_4300,N_3184,N_3360);
and U4301 (N_4301,N_3324,N_3411);
or U4302 (N_4302,N_3157,N_3209);
nand U4303 (N_4303,N_3622,N_3337);
nor U4304 (N_4304,N_3434,N_3376);
nand U4305 (N_4305,N_3196,N_3520);
nand U4306 (N_4306,N_3153,N_3164);
and U4307 (N_4307,N_3139,N_3631);
nand U4308 (N_4308,N_3555,N_3577);
nand U4309 (N_4309,N_3188,N_3504);
and U4310 (N_4310,N_3314,N_3521);
nand U4311 (N_4311,N_3606,N_3644);
nand U4312 (N_4312,N_3291,N_3128);
or U4313 (N_4313,N_3600,N_3588);
nor U4314 (N_4314,N_3300,N_3457);
xor U4315 (N_4315,N_3665,N_3495);
nand U4316 (N_4316,N_3126,N_3451);
xor U4317 (N_4317,N_3125,N_3322);
or U4318 (N_4318,N_3306,N_3455);
xnor U4319 (N_4319,N_3510,N_3305);
nor U4320 (N_4320,N_3466,N_3458);
nor U4321 (N_4321,N_3467,N_3148);
and U4322 (N_4322,N_3330,N_3303);
nand U4323 (N_4323,N_3312,N_3134);
nor U4324 (N_4324,N_3219,N_3332);
xor U4325 (N_4325,N_3472,N_3429);
and U4326 (N_4326,N_3696,N_3707);
nand U4327 (N_4327,N_3649,N_3564);
nand U4328 (N_4328,N_3612,N_3215);
nor U4329 (N_4329,N_3599,N_3386);
nor U4330 (N_4330,N_3226,N_3213);
and U4331 (N_4331,N_3358,N_3527);
or U4332 (N_4332,N_3243,N_3665);
xnor U4333 (N_4333,N_3240,N_3485);
nand U4334 (N_4334,N_3642,N_3432);
nor U4335 (N_4335,N_3692,N_3213);
and U4336 (N_4336,N_3353,N_3231);
or U4337 (N_4337,N_3390,N_3220);
xnor U4338 (N_4338,N_3713,N_3175);
and U4339 (N_4339,N_3314,N_3589);
or U4340 (N_4340,N_3287,N_3316);
nand U4341 (N_4341,N_3430,N_3699);
nand U4342 (N_4342,N_3663,N_3519);
and U4343 (N_4343,N_3601,N_3153);
xor U4344 (N_4344,N_3408,N_3672);
or U4345 (N_4345,N_3422,N_3157);
xnor U4346 (N_4346,N_3447,N_3599);
nand U4347 (N_4347,N_3494,N_3514);
nand U4348 (N_4348,N_3329,N_3675);
nor U4349 (N_4349,N_3584,N_3233);
or U4350 (N_4350,N_3673,N_3405);
or U4351 (N_4351,N_3702,N_3294);
or U4352 (N_4352,N_3332,N_3642);
or U4353 (N_4353,N_3513,N_3496);
nand U4354 (N_4354,N_3588,N_3341);
and U4355 (N_4355,N_3709,N_3380);
nor U4356 (N_4356,N_3249,N_3581);
and U4357 (N_4357,N_3624,N_3611);
or U4358 (N_4358,N_3130,N_3709);
xnor U4359 (N_4359,N_3211,N_3416);
nand U4360 (N_4360,N_3709,N_3747);
or U4361 (N_4361,N_3361,N_3536);
nor U4362 (N_4362,N_3148,N_3681);
nor U4363 (N_4363,N_3146,N_3733);
nand U4364 (N_4364,N_3562,N_3144);
or U4365 (N_4365,N_3294,N_3436);
xnor U4366 (N_4366,N_3567,N_3376);
xnor U4367 (N_4367,N_3703,N_3590);
and U4368 (N_4368,N_3425,N_3624);
xor U4369 (N_4369,N_3238,N_3725);
nand U4370 (N_4370,N_3192,N_3247);
nor U4371 (N_4371,N_3363,N_3612);
or U4372 (N_4372,N_3672,N_3405);
nor U4373 (N_4373,N_3594,N_3734);
nand U4374 (N_4374,N_3605,N_3329);
nor U4375 (N_4375,N_4168,N_4072);
xor U4376 (N_4376,N_3798,N_3916);
nor U4377 (N_4377,N_4036,N_3751);
nand U4378 (N_4378,N_4262,N_3838);
or U4379 (N_4379,N_4235,N_4027);
nand U4380 (N_4380,N_4311,N_3826);
nor U4381 (N_4381,N_4207,N_4154);
nand U4382 (N_4382,N_3781,N_3976);
and U4383 (N_4383,N_4218,N_4361);
or U4384 (N_4384,N_3753,N_3836);
or U4385 (N_4385,N_3914,N_3946);
nor U4386 (N_4386,N_4170,N_3839);
nor U4387 (N_4387,N_3789,N_3915);
and U4388 (N_4388,N_3938,N_4236);
and U4389 (N_4389,N_4232,N_4360);
and U4390 (N_4390,N_3876,N_4030);
and U4391 (N_4391,N_4108,N_4195);
nand U4392 (N_4392,N_4251,N_4272);
and U4393 (N_4393,N_4191,N_4045);
nor U4394 (N_4394,N_4369,N_3845);
or U4395 (N_4395,N_4127,N_4362);
and U4396 (N_4396,N_4265,N_4259);
nor U4397 (N_4397,N_4279,N_4355);
or U4398 (N_4398,N_3923,N_4142);
xor U4399 (N_4399,N_3887,N_4321);
nor U4400 (N_4400,N_3961,N_3981);
or U4401 (N_4401,N_4283,N_4303);
or U4402 (N_4402,N_4028,N_4084);
nor U4403 (N_4403,N_4131,N_3984);
and U4404 (N_4404,N_4284,N_4140);
nor U4405 (N_4405,N_4136,N_3899);
nand U4406 (N_4406,N_4271,N_4275);
nor U4407 (N_4407,N_4128,N_4346);
xnor U4408 (N_4408,N_3910,N_4367);
nor U4409 (N_4409,N_4242,N_3776);
nor U4410 (N_4410,N_4225,N_3891);
and U4411 (N_4411,N_3968,N_3985);
xor U4412 (N_4412,N_4181,N_3783);
nand U4413 (N_4413,N_4192,N_4281);
xor U4414 (N_4414,N_4081,N_3861);
nor U4415 (N_4415,N_3969,N_3955);
nor U4416 (N_4416,N_4290,N_3778);
nor U4417 (N_4417,N_3897,N_4282);
nand U4418 (N_4418,N_3900,N_3892);
or U4419 (N_4419,N_4101,N_4096);
and U4420 (N_4420,N_3756,N_3911);
nor U4421 (N_4421,N_3801,N_4021);
xnor U4422 (N_4422,N_4010,N_4014);
or U4423 (N_4423,N_3944,N_4009);
or U4424 (N_4424,N_3941,N_4292);
nor U4425 (N_4425,N_4374,N_3820);
xor U4426 (N_4426,N_3926,N_3952);
nand U4427 (N_4427,N_3912,N_3840);
and U4428 (N_4428,N_4188,N_4163);
nand U4429 (N_4429,N_4125,N_4050);
and U4430 (N_4430,N_3791,N_3805);
nor U4431 (N_4431,N_4370,N_3975);
nor U4432 (N_4432,N_3994,N_4352);
nor U4433 (N_4433,N_4075,N_4341);
nor U4434 (N_4434,N_4239,N_4147);
nor U4435 (N_4435,N_3764,N_4371);
or U4436 (N_4436,N_4260,N_3886);
nand U4437 (N_4437,N_4344,N_3823);
nand U4438 (N_4438,N_4059,N_4330);
and U4439 (N_4439,N_4230,N_4372);
nor U4440 (N_4440,N_4250,N_3990);
nand U4441 (N_4441,N_3959,N_4247);
and U4442 (N_4442,N_4106,N_3799);
and U4443 (N_4443,N_4245,N_4171);
or U4444 (N_4444,N_4306,N_4035);
xor U4445 (N_4445,N_3868,N_4209);
nor U4446 (N_4446,N_4308,N_4165);
and U4447 (N_4447,N_4336,N_4307);
nand U4448 (N_4448,N_4004,N_4095);
nor U4449 (N_4449,N_3812,N_4276);
or U4450 (N_4450,N_4020,N_4343);
nand U4451 (N_4451,N_4176,N_4196);
nand U4452 (N_4452,N_3935,N_4257);
nor U4453 (N_4453,N_4280,N_3875);
nor U4454 (N_4454,N_4324,N_4037);
nor U4455 (N_4455,N_4179,N_4120);
and U4456 (N_4456,N_4150,N_4193);
nand U4457 (N_4457,N_4286,N_3795);
nand U4458 (N_4458,N_4309,N_3962);
nand U4459 (N_4459,N_3752,N_4219);
nor U4460 (N_4460,N_3894,N_3794);
or U4461 (N_4461,N_3870,N_3869);
nor U4462 (N_4462,N_3804,N_3829);
and U4463 (N_4463,N_4363,N_3768);
and U4464 (N_4464,N_3879,N_4194);
or U4465 (N_4465,N_3754,N_4048);
nand U4466 (N_4466,N_3831,N_4186);
nor U4467 (N_4467,N_4214,N_4231);
xor U4468 (N_4468,N_4064,N_4001);
or U4469 (N_4469,N_3850,N_4203);
nand U4470 (N_4470,N_3878,N_4301);
nor U4471 (N_4471,N_4055,N_4200);
or U4472 (N_4472,N_3982,N_4118);
and U4473 (N_4473,N_3987,N_4228);
nor U4474 (N_4474,N_3785,N_3889);
and U4475 (N_4475,N_4085,N_3950);
nand U4476 (N_4476,N_4076,N_4318);
nand U4477 (N_4477,N_3880,N_3999);
nor U4478 (N_4478,N_4098,N_3821);
xor U4479 (N_4479,N_4305,N_4294);
xor U4480 (N_4480,N_3933,N_3943);
nor U4481 (N_4481,N_4172,N_3983);
and U4482 (N_4482,N_4152,N_4331);
and U4483 (N_4483,N_3874,N_4008);
and U4484 (N_4484,N_4099,N_3996);
or U4485 (N_4485,N_4089,N_4267);
or U4486 (N_4486,N_3810,N_3864);
nand U4487 (N_4487,N_3815,N_3967);
and U4488 (N_4488,N_4123,N_4146);
xnor U4489 (N_4489,N_3757,N_4220);
nor U4490 (N_4490,N_3860,N_4103);
and U4491 (N_4491,N_4326,N_4148);
or U4492 (N_4492,N_3951,N_3928);
nor U4493 (N_4493,N_4164,N_3947);
and U4494 (N_4494,N_3858,N_3929);
and U4495 (N_4495,N_4162,N_3792);
nor U4496 (N_4496,N_4046,N_3877);
nand U4497 (N_4497,N_4079,N_4051);
nor U4498 (N_4498,N_3822,N_3960);
and U4499 (N_4499,N_4077,N_4130);
nor U4500 (N_4500,N_3970,N_4047);
nand U4501 (N_4501,N_4080,N_4299);
and U4502 (N_4502,N_3787,N_4012);
and U4503 (N_4503,N_4356,N_4115);
and U4504 (N_4504,N_4145,N_3957);
nor U4505 (N_4505,N_3842,N_3883);
nor U4506 (N_4506,N_4011,N_4351);
nor U4507 (N_4507,N_4183,N_3991);
nand U4508 (N_4508,N_3818,N_4068);
nor U4509 (N_4509,N_4358,N_3817);
or U4510 (N_4510,N_3847,N_4062);
xnor U4511 (N_4511,N_4302,N_4082);
nor U4512 (N_4512,N_4222,N_3766);
and U4513 (N_4513,N_3846,N_4199);
nor U4514 (N_4514,N_4070,N_4138);
nand U4515 (N_4515,N_4015,N_3936);
and U4516 (N_4516,N_4052,N_4169);
nand U4517 (N_4517,N_3963,N_4003);
nand U4518 (N_4518,N_4058,N_4342);
or U4519 (N_4519,N_3909,N_4325);
nand U4520 (N_4520,N_4086,N_3898);
and U4521 (N_4521,N_3857,N_4041);
and U4522 (N_4522,N_4017,N_4285);
nand U4523 (N_4523,N_3828,N_3927);
or U4524 (N_4524,N_4365,N_3777);
nor U4525 (N_4525,N_4093,N_3977);
and U4526 (N_4526,N_3956,N_4110);
nor U4527 (N_4527,N_3906,N_3920);
nand U4528 (N_4528,N_4026,N_4274);
or U4529 (N_4529,N_4246,N_4069);
nor U4530 (N_4530,N_3881,N_4178);
nor U4531 (N_4531,N_4102,N_4024);
xnor U4532 (N_4532,N_3786,N_4073);
and U4533 (N_4533,N_3973,N_3964);
and U4534 (N_4534,N_3871,N_3827);
xor U4535 (N_4535,N_4354,N_3837);
nor U4536 (N_4536,N_3930,N_3953);
or U4537 (N_4537,N_4208,N_4189);
and U4538 (N_4538,N_4006,N_4206);
nand U4539 (N_4539,N_4252,N_3775);
or U4540 (N_4540,N_4078,N_4322);
and U4541 (N_4541,N_3770,N_4071);
and U4542 (N_4542,N_4323,N_3908);
nor U4543 (N_4543,N_4134,N_3948);
nand U4544 (N_4544,N_4234,N_4213);
or U4545 (N_4545,N_3852,N_4184);
and U4546 (N_4546,N_4107,N_4143);
nand U4547 (N_4547,N_3859,N_3767);
and U4548 (N_4548,N_3772,N_4105);
or U4549 (N_4549,N_3793,N_4278);
nand U4550 (N_4550,N_4122,N_3755);
nor U4551 (N_4551,N_4113,N_3882);
and U4552 (N_4552,N_4273,N_4157);
nand U4553 (N_4553,N_4111,N_4244);
or U4554 (N_4554,N_3763,N_4097);
and U4555 (N_4555,N_3790,N_4298);
nand U4556 (N_4556,N_3865,N_4335);
nor U4557 (N_4557,N_3867,N_3800);
and U4558 (N_4558,N_3934,N_4315);
and U4559 (N_4559,N_3972,N_4211);
nand U4560 (N_4560,N_3974,N_3945);
or U4561 (N_4561,N_4151,N_4087);
or U4562 (N_4562,N_4243,N_3843);
or U4563 (N_4563,N_4263,N_4060);
or U4564 (N_4564,N_3856,N_4061);
nor U4565 (N_4565,N_4197,N_4031);
nand U4566 (N_4566,N_3844,N_3803);
nor U4567 (N_4567,N_3966,N_4129);
nor U4568 (N_4568,N_4182,N_3758);
nor U4569 (N_4569,N_3807,N_4340);
xnor U4570 (N_4570,N_4187,N_3913);
or U4571 (N_4571,N_3940,N_3905);
and U4572 (N_4572,N_4039,N_4185);
and U4573 (N_4573,N_3816,N_4224);
xor U4574 (N_4574,N_3895,N_4177);
xor U4575 (N_4575,N_3902,N_4221);
or U4576 (N_4576,N_3841,N_4266);
and U4577 (N_4577,N_4054,N_4347);
and U4578 (N_4578,N_3808,N_4043);
or U4579 (N_4579,N_4166,N_3809);
and U4580 (N_4580,N_4233,N_4268);
xnor U4581 (N_4581,N_3997,N_4067);
nand U4582 (N_4582,N_4065,N_3971);
xor U4583 (N_4583,N_4114,N_4141);
nand U4584 (N_4584,N_3788,N_3896);
xnor U4585 (N_4585,N_3949,N_3922);
or U4586 (N_4586,N_4353,N_4173);
nor U4587 (N_4587,N_4319,N_4022);
nand U4588 (N_4588,N_3918,N_3782);
xor U4589 (N_4589,N_4332,N_3888);
nand U4590 (N_4590,N_4237,N_4180);
and U4591 (N_4591,N_3819,N_4212);
nand U4592 (N_4592,N_4345,N_4277);
or U4593 (N_4593,N_4159,N_4329);
nand U4594 (N_4594,N_4112,N_3863);
nand U4595 (N_4595,N_4057,N_4124);
and U4596 (N_4596,N_4204,N_4033);
and U4597 (N_4597,N_3761,N_4223);
nor U4598 (N_4598,N_4074,N_3773);
nor U4599 (N_4599,N_4100,N_4063);
nor U4600 (N_4600,N_4005,N_4155);
and U4601 (N_4601,N_4032,N_3884);
and U4602 (N_4602,N_3835,N_4132);
nand U4603 (N_4603,N_4025,N_3901);
nor U4604 (N_4604,N_4042,N_4190);
nand U4605 (N_4605,N_3903,N_3924);
nor U4606 (N_4606,N_4314,N_3995);
nand U4607 (N_4607,N_4119,N_4161);
and U4608 (N_4608,N_3796,N_3851);
and U4609 (N_4609,N_3769,N_4217);
nand U4610 (N_4610,N_4296,N_3872);
nand U4611 (N_4611,N_3832,N_4158);
nor U4612 (N_4612,N_3942,N_3954);
xor U4613 (N_4613,N_3925,N_3890);
nand U4614 (N_4614,N_4091,N_4040);
nor U4615 (N_4615,N_3771,N_3989);
nand U4616 (N_4616,N_4295,N_4349);
nor U4617 (N_4617,N_3921,N_4049);
nor U4618 (N_4618,N_4291,N_3907);
nor U4619 (N_4619,N_3762,N_4202);
nand U4620 (N_4620,N_4255,N_3774);
and U4621 (N_4621,N_3866,N_4104);
nand U4622 (N_4622,N_4216,N_3834);
and U4623 (N_4623,N_3806,N_4313);
and U4624 (N_4624,N_4248,N_3760);
nand U4625 (N_4625,N_3780,N_4320);
nor U4626 (N_4626,N_3917,N_3873);
and U4627 (N_4627,N_3814,N_4328);
and U4628 (N_4628,N_4368,N_4034);
and U4629 (N_4629,N_3978,N_4092);
or U4630 (N_4630,N_3824,N_4254);
or U4631 (N_4631,N_3988,N_4317);
or U4632 (N_4632,N_3853,N_4339);
and U4633 (N_4633,N_4334,N_4258);
xnor U4634 (N_4634,N_4269,N_4373);
nor U4635 (N_4635,N_3986,N_4000);
and U4636 (N_4636,N_4066,N_3779);
nor U4637 (N_4637,N_4153,N_4312);
and U4638 (N_4638,N_4016,N_4288);
nor U4639 (N_4639,N_4333,N_3797);
or U4640 (N_4640,N_3750,N_4149);
xor U4641 (N_4641,N_4241,N_3904);
and U4642 (N_4642,N_4287,N_4229);
or U4643 (N_4643,N_3765,N_4366);
and U4644 (N_4644,N_4327,N_3759);
nor U4645 (N_4645,N_3931,N_3811);
or U4646 (N_4646,N_3919,N_3939);
nand U4647 (N_4647,N_4044,N_3849);
nor U4648 (N_4648,N_4238,N_4175);
nand U4649 (N_4649,N_4310,N_4364);
or U4650 (N_4650,N_4264,N_4201);
and U4651 (N_4651,N_4240,N_4133);
nor U4652 (N_4652,N_4174,N_4297);
nand U4653 (N_4653,N_4023,N_4126);
nand U4654 (N_4654,N_4256,N_4359);
and U4655 (N_4655,N_4088,N_4135);
nor U4656 (N_4656,N_4304,N_4038);
and U4657 (N_4657,N_3958,N_3854);
and U4658 (N_4658,N_4293,N_3813);
or U4659 (N_4659,N_3802,N_3980);
and U4660 (N_4660,N_4109,N_4018);
or U4661 (N_4661,N_4337,N_4205);
and U4662 (N_4662,N_3965,N_3993);
nor U4663 (N_4663,N_4090,N_3893);
xnor U4664 (N_4664,N_3998,N_4094);
nand U4665 (N_4665,N_3992,N_3855);
xor U4666 (N_4666,N_4261,N_4160);
nand U4667 (N_4667,N_4270,N_4137);
nand U4668 (N_4668,N_4019,N_4007);
or U4669 (N_4669,N_4117,N_3833);
or U4670 (N_4670,N_4226,N_4198);
and U4671 (N_4671,N_4053,N_3862);
or U4672 (N_4672,N_3979,N_3825);
and U4673 (N_4673,N_4056,N_4338);
xor U4674 (N_4674,N_4116,N_4013);
nand U4675 (N_4675,N_4144,N_4253);
nor U4676 (N_4676,N_3830,N_4300);
nor U4677 (N_4677,N_4316,N_3784);
or U4678 (N_4678,N_4357,N_4215);
or U4679 (N_4679,N_4210,N_4029);
or U4680 (N_4680,N_4156,N_4167);
and U4681 (N_4681,N_4350,N_3932);
or U4682 (N_4682,N_3885,N_4249);
or U4683 (N_4683,N_4002,N_4227);
and U4684 (N_4684,N_4083,N_4121);
or U4685 (N_4685,N_3937,N_4289);
nor U4686 (N_4686,N_3848,N_4348);
and U4687 (N_4687,N_4139,N_3993);
xor U4688 (N_4688,N_4159,N_4212);
nor U4689 (N_4689,N_3854,N_4260);
nor U4690 (N_4690,N_4143,N_4159);
and U4691 (N_4691,N_4352,N_4046);
or U4692 (N_4692,N_4008,N_3939);
nand U4693 (N_4693,N_3777,N_4300);
nor U4694 (N_4694,N_3790,N_4318);
nand U4695 (N_4695,N_4155,N_4226);
and U4696 (N_4696,N_3756,N_4249);
nor U4697 (N_4697,N_4056,N_4171);
or U4698 (N_4698,N_4009,N_4223);
nor U4699 (N_4699,N_4265,N_4189);
nor U4700 (N_4700,N_3757,N_4147);
xor U4701 (N_4701,N_3917,N_4109);
nor U4702 (N_4702,N_3930,N_3809);
xor U4703 (N_4703,N_4262,N_4085);
nor U4704 (N_4704,N_3842,N_3972);
and U4705 (N_4705,N_4133,N_3785);
xnor U4706 (N_4706,N_3832,N_4062);
nor U4707 (N_4707,N_4129,N_3950);
xor U4708 (N_4708,N_3958,N_4058);
or U4709 (N_4709,N_4106,N_3833);
nand U4710 (N_4710,N_4367,N_4373);
and U4711 (N_4711,N_4218,N_4325);
or U4712 (N_4712,N_4113,N_4297);
and U4713 (N_4713,N_4086,N_4364);
and U4714 (N_4714,N_4040,N_4103);
nand U4715 (N_4715,N_3868,N_4232);
xnor U4716 (N_4716,N_3888,N_4345);
and U4717 (N_4717,N_3930,N_3873);
nor U4718 (N_4718,N_4022,N_4135);
nor U4719 (N_4719,N_3890,N_3878);
or U4720 (N_4720,N_4369,N_4283);
and U4721 (N_4721,N_4294,N_4028);
nor U4722 (N_4722,N_3929,N_3936);
and U4723 (N_4723,N_3790,N_4271);
nand U4724 (N_4724,N_4191,N_4041);
xor U4725 (N_4725,N_4247,N_3961);
and U4726 (N_4726,N_3881,N_4277);
nand U4727 (N_4727,N_3852,N_4065);
and U4728 (N_4728,N_4313,N_4200);
nand U4729 (N_4729,N_4280,N_4069);
xnor U4730 (N_4730,N_4224,N_3762);
or U4731 (N_4731,N_4341,N_4199);
or U4732 (N_4732,N_4190,N_4228);
nor U4733 (N_4733,N_3782,N_4291);
and U4734 (N_4734,N_4033,N_4218);
or U4735 (N_4735,N_4164,N_4124);
or U4736 (N_4736,N_3828,N_3783);
nor U4737 (N_4737,N_4260,N_4215);
nand U4738 (N_4738,N_4125,N_3876);
or U4739 (N_4739,N_3961,N_3863);
or U4740 (N_4740,N_3864,N_4299);
nand U4741 (N_4741,N_3847,N_4066);
or U4742 (N_4742,N_3984,N_4041);
and U4743 (N_4743,N_3963,N_4287);
or U4744 (N_4744,N_3963,N_3924);
nand U4745 (N_4745,N_3804,N_3971);
or U4746 (N_4746,N_4051,N_4261);
and U4747 (N_4747,N_4022,N_3819);
nand U4748 (N_4748,N_3765,N_3775);
or U4749 (N_4749,N_4127,N_4368);
and U4750 (N_4750,N_3824,N_4216);
xnor U4751 (N_4751,N_4360,N_4040);
or U4752 (N_4752,N_4225,N_3804);
and U4753 (N_4753,N_4040,N_4281);
nand U4754 (N_4754,N_3816,N_3768);
and U4755 (N_4755,N_4225,N_4292);
nand U4756 (N_4756,N_3816,N_3758);
nand U4757 (N_4757,N_4349,N_3877);
and U4758 (N_4758,N_4261,N_4155);
and U4759 (N_4759,N_4342,N_4345);
nand U4760 (N_4760,N_4081,N_3819);
nand U4761 (N_4761,N_4323,N_4086);
and U4762 (N_4762,N_3974,N_3789);
and U4763 (N_4763,N_4151,N_4230);
nor U4764 (N_4764,N_4306,N_3963);
xnor U4765 (N_4765,N_3805,N_4280);
nor U4766 (N_4766,N_4338,N_3816);
nor U4767 (N_4767,N_3861,N_3935);
or U4768 (N_4768,N_4066,N_4063);
nand U4769 (N_4769,N_3965,N_4194);
or U4770 (N_4770,N_4146,N_4002);
xor U4771 (N_4771,N_4212,N_4304);
xor U4772 (N_4772,N_4172,N_3776);
nor U4773 (N_4773,N_4079,N_4123);
or U4774 (N_4774,N_4343,N_4219);
nand U4775 (N_4775,N_3979,N_3899);
or U4776 (N_4776,N_4142,N_4166);
and U4777 (N_4777,N_3983,N_3963);
nand U4778 (N_4778,N_4253,N_4233);
nor U4779 (N_4779,N_4030,N_4099);
and U4780 (N_4780,N_4368,N_3968);
or U4781 (N_4781,N_3890,N_4341);
or U4782 (N_4782,N_4017,N_3993);
nor U4783 (N_4783,N_4213,N_3912);
nor U4784 (N_4784,N_4097,N_3888);
nand U4785 (N_4785,N_4183,N_4279);
nor U4786 (N_4786,N_3939,N_4327);
xnor U4787 (N_4787,N_3839,N_4269);
or U4788 (N_4788,N_4087,N_4081);
nor U4789 (N_4789,N_4353,N_3904);
nor U4790 (N_4790,N_3848,N_3779);
or U4791 (N_4791,N_3890,N_4081);
xor U4792 (N_4792,N_4039,N_3986);
and U4793 (N_4793,N_3986,N_3763);
and U4794 (N_4794,N_4034,N_3957);
or U4795 (N_4795,N_4136,N_3886);
and U4796 (N_4796,N_4017,N_4258);
and U4797 (N_4797,N_4107,N_4229);
nor U4798 (N_4798,N_3964,N_3885);
or U4799 (N_4799,N_4255,N_4260);
or U4800 (N_4800,N_4335,N_3900);
nor U4801 (N_4801,N_3992,N_3876);
nand U4802 (N_4802,N_3987,N_4033);
nor U4803 (N_4803,N_4307,N_3837);
and U4804 (N_4804,N_4144,N_4357);
nor U4805 (N_4805,N_4131,N_3929);
nor U4806 (N_4806,N_3991,N_3930);
and U4807 (N_4807,N_3965,N_4298);
or U4808 (N_4808,N_4075,N_4361);
nand U4809 (N_4809,N_3888,N_4153);
nor U4810 (N_4810,N_3992,N_4269);
nand U4811 (N_4811,N_3750,N_4039);
or U4812 (N_4812,N_4303,N_3778);
and U4813 (N_4813,N_3992,N_4139);
or U4814 (N_4814,N_3933,N_3774);
nor U4815 (N_4815,N_4340,N_3861);
nor U4816 (N_4816,N_4120,N_4012);
nor U4817 (N_4817,N_3931,N_4035);
nand U4818 (N_4818,N_4214,N_4066);
and U4819 (N_4819,N_4078,N_4269);
xor U4820 (N_4820,N_4077,N_3981);
and U4821 (N_4821,N_4168,N_3938);
xor U4822 (N_4822,N_4289,N_4342);
nand U4823 (N_4823,N_3962,N_4285);
xnor U4824 (N_4824,N_3892,N_4287);
and U4825 (N_4825,N_3817,N_4027);
and U4826 (N_4826,N_4341,N_4122);
nor U4827 (N_4827,N_3783,N_3877);
and U4828 (N_4828,N_3762,N_4305);
and U4829 (N_4829,N_3821,N_3850);
nand U4830 (N_4830,N_4148,N_4003);
nand U4831 (N_4831,N_4137,N_3939);
nor U4832 (N_4832,N_4328,N_3893);
or U4833 (N_4833,N_4151,N_3857);
and U4834 (N_4834,N_4359,N_4272);
or U4835 (N_4835,N_3789,N_4065);
and U4836 (N_4836,N_4374,N_3763);
or U4837 (N_4837,N_3854,N_4257);
and U4838 (N_4838,N_4251,N_4171);
nand U4839 (N_4839,N_4118,N_4366);
nand U4840 (N_4840,N_4262,N_4287);
or U4841 (N_4841,N_4325,N_4129);
nor U4842 (N_4842,N_3894,N_4296);
nor U4843 (N_4843,N_3934,N_3776);
xor U4844 (N_4844,N_4294,N_4324);
nor U4845 (N_4845,N_3786,N_4186);
or U4846 (N_4846,N_4316,N_4179);
nand U4847 (N_4847,N_4075,N_3912);
or U4848 (N_4848,N_4178,N_4116);
nor U4849 (N_4849,N_4006,N_4089);
or U4850 (N_4850,N_4082,N_4278);
nor U4851 (N_4851,N_4039,N_4045);
or U4852 (N_4852,N_3941,N_4136);
or U4853 (N_4853,N_4176,N_4146);
or U4854 (N_4854,N_3965,N_4358);
nand U4855 (N_4855,N_4246,N_3772);
nor U4856 (N_4856,N_3968,N_4004);
or U4857 (N_4857,N_4061,N_3901);
and U4858 (N_4858,N_3991,N_3977);
nand U4859 (N_4859,N_4117,N_3904);
or U4860 (N_4860,N_3900,N_4009);
nand U4861 (N_4861,N_4330,N_3800);
and U4862 (N_4862,N_3839,N_3751);
nor U4863 (N_4863,N_4335,N_3923);
and U4864 (N_4864,N_4357,N_4308);
and U4865 (N_4865,N_3843,N_4132);
nor U4866 (N_4866,N_4280,N_4219);
nor U4867 (N_4867,N_4081,N_4150);
or U4868 (N_4868,N_4038,N_3847);
or U4869 (N_4869,N_3813,N_4053);
nand U4870 (N_4870,N_4074,N_3904);
or U4871 (N_4871,N_4270,N_4240);
or U4872 (N_4872,N_3792,N_4039);
xnor U4873 (N_4873,N_4255,N_4162);
and U4874 (N_4874,N_3944,N_3829);
nand U4875 (N_4875,N_4040,N_4067);
nor U4876 (N_4876,N_4098,N_4113);
or U4877 (N_4877,N_4033,N_3816);
xor U4878 (N_4878,N_3891,N_3824);
or U4879 (N_4879,N_4041,N_4049);
or U4880 (N_4880,N_4312,N_3931);
or U4881 (N_4881,N_4314,N_4151);
nor U4882 (N_4882,N_3850,N_3849);
xnor U4883 (N_4883,N_4030,N_3963);
xor U4884 (N_4884,N_3961,N_4014);
or U4885 (N_4885,N_4126,N_4308);
and U4886 (N_4886,N_3803,N_4009);
nor U4887 (N_4887,N_4207,N_4284);
and U4888 (N_4888,N_4231,N_3803);
xnor U4889 (N_4889,N_3795,N_3970);
nand U4890 (N_4890,N_4210,N_4315);
nand U4891 (N_4891,N_4289,N_4339);
and U4892 (N_4892,N_4166,N_4028);
and U4893 (N_4893,N_3885,N_3855);
or U4894 (N_4894,N_4356,N_3931);
xnor U4895 (N_4895,N_3789,N_3896);
or U4896 (N_4896,N_3862,N_3925);
xor U4897 (N_4897,N_3956,N_4111);
and U4898 (N_4898,N_4329,N_4299);
nand U4899 (N_4899,N_4109,N_4318);
and U4900 (N_4900,N_4113,N_4172);
or U4901 (N_4901,N_4257,N_3967);
nand U4902 (N_4902,N_3914,N_3844);
and U4903 (N_4903,N_4304,N_3983);
or U4904 (N_4904,N_4305,N_4169);
or U4905 (N_4905,N_4173,N_3992);
xor U4906 (N_4906,N_4292,N_3820);
nand U4907 (N_4907,N_4169,N_3999);
nor U4908 (N_4908,N_3914,N_4263);
xor U4909 (N_4909,N_4048,N_4265);
nand U4910 (N_4910,N_4216,N_4160);
nand U4911 (N_4911,N_3842,N_4106);
nor U4912 (N_4912,N_4340,N_3885);
nor U4913 (N_4913,N_3775,N_4092);
and U4914 (N_4914,N_4106,N_4317);
or U4915 (N_4915,N_3773,N_4041);
or U4916 (N_4916,N_3800,N_4369);
and U4917 (N_4917,N_4157,N_4063);
nor U4918 (N_4918,N_3995,N_4292);
and U4919 (N_4919,N_3763,N_4050);
nand U4920 (N_4920,N_4046,N_4040);
or U4921 (N_4921,N_3981,N_4099);
nand U4922 (N_4922,N_3793,N_4347);
or U4923 (N_4923,N_4059,N_4057);
nor U4924 (N_4924,N_3860,N_4330);
xnor U4925 (N_4925,N_3839,N_3784);
and U4926 (N_4926,N_3751,N_4028);
nand U4927 (N_4927,N_4298,N_4324);
and U4928 (N_4928,N_4130,N_4098);
and U4929 (N_4929,N_4117,N_4265);
nand U4930 (N_4930,N_3867,N_4207);
or U4931 (N_4931,N_4071,N_4052);
nand U4932 (N_4932,N_4372,N_4171);
and U4933 (N_4933,N_4238,N_4016);
nor U4934 (N_4934,N_3956,N_4091);
nor U4935 (N_4935,N_3850,N_4126);
nor U4936 (N_4936,N_3977,N_4096);
or U4937 (N_4937,N_4237,N_3927);
nand U4938 (N_4938,N_3837,N_3934);
and U4939 (N_4939,N_4053,N_4295);
and U4940 (N_4940,N_4357,N_4102);
nand U4941 (N_4941,N_3835,N_4145);
and U4942 (N_4942,N_3955,N_3886);
nand U4943 (N_4943,N_3779,N_3866);
nor U4944 (N_4944,N_3846,N_3972);
nand U4945 (N_4945,N_4023,N_3853);
or U4946 (N_4946,N_4266,N_4158);
nor U4947 (N_4947,N_3938,N_4130);
nand U4948 (N_4948,N_3874,N_3812);
nand U4949 (N_4949,N_3991,N_3994);
nand U4950 (N_4950,N_3773,N_4135);
and U4951 (N_4951,N_4052,N_4217);
nand U4952 (N_4952,N_3794,N_3846);
nor U4953 (N_4953,N_3927,N_4082);
or U4954 (N_4954,N_4340,N_4039);
nor U4955 (N_4955,N_4064,N_3847);
and U4956 (N_4956,N_3800,N_4139);
or U4957 (N_4957,N_4334,N_4143);
nand U4958 (N_4958,N_3829,N_3949);
and U4959 (N_4959,N_4179,N_4185);
nand U4960 (N_4960,N_3996,N_3934);
nand U4961 (N_4961,N_4150,N_3935);
nand U4962 (N_4962,N_3860,N_4087);
and U4963 (N_4963,N_4235,N_4220);
nor U4964 (N_4964,N_3757,N_3827);
nor U4965 (N_4965,N_4098,N_4093);
or U4966 (N_4966,N_3952,N_4006);
or U4967 (N_4967,N_4297,N_3877);
or U4968 (N_4968,N_4297,N_4103);
xor U4969 (N_4969,N_3859,N_3751);
or U4970 (N_4970,N_4228,N_4373);
nand U4971 (N_4971,N_4336,N_4185);
and U4972 (N_4972,N_3958,N_3860);
nand U4973 (N_4973,N_4075,N_4068);
nand U4974 (N_4974,N_4323,N_4047);
nor U4975 (N_4975,N_3822,N_4139);
nand U4976 (N_4976,N_3883,N_4152);
nand U4977 (N_4977,N_3849,N_4007);
xnor U4978 (N_4978,N_4313,N_4017);
and U4979 (N_4979,N_3796,N_3941);
xor U4980 (N_4980,N_4145,N_3777);
and U4981 (N_4981,N_4246,N_4323);
nand U4982 (N_4982,N_4146,N_3916);
and U4983 (N_4983,N_4069,N_3987);
xor U4984 (N_4984,N_3926,N_4233);
nand U4985 (N_4985,N_3909,N_4056);
and U4986 (N_4986,N_4302,N_3998);
xor U4987 (N_4987,N_3962,N_4190);
or U4988 (N_4988,N_4209,N_4189);
nand U4989 (N_4989,N_4336,N_3754);
nor U4990 (N_4990,N_4222,N_3955);
or U4991 (N_4991,N_4037,N_4144);
or U4992 (N_4992,N_4354,N_4299);
and U4993 (N_4993,N_4365,N_4343);
xor U4994 (N_4994,N_3794,N_4373);
and U4995 (N_4995,N_4166,N_4032);
nand U4996 (N_4996,N_3936,N_3893);
and U4997 (N_4997,N_3964,N_4191);
and U4998 (N_4998,N_3921,N_4249);
nor U4999 (N_4999,N_4191,N_4072);
nor U5000 (N_5000,N_4933,N_4862);
nor U5001 (N_5001,N_4400,N_4528);
xor U5002 (N_5002,N_4410,N_4957);
or U5003 (N_5003,N_4585,N_4503);
xor U5004 (N_5004,N_4785,N_4834);
nor U5005 (N_5005,N_4449,N_4548);
and U5006 (N_5006,N_4611,N_4525);
nand U5007 (N_5007,N_4388,N_4599);
nor U5008 (N_5008,N_4586,N_4880);
or U5009 (N_5009,N_4536,N_4533);
and U5010 (N_5010,N_4502,N_4865);
xnor U5011 (N_5011,N_4382,N_4812);
nor U5012 (N_5012,N_4676,N_4402);
xnor U5013 (N_5013,N_4830,N_4538);
or U5014 (N_5014,N_4491,N_4658);
or U5015 (N_5015,N_4850,N_4390);
nor U5016 (N_5016,N_4967,N_4889);
nor U5017 (N_5017,N_4455,N_4392);
and U5018 (N_5018,N_4732,N_4387);
and U5019 (N_5019,N_4976,N_4484);
and U5020 (N_5020,N_4975,N_4762);
xor U5021 (N_5021,N_4621,N_4842);
and U5022 (N_5022,N_4747,N_4645);
xnor U5023 (N_5023,N_4495,N_4463);
xnor U5024 (N_5024,N_4913,N_4663);
or U5025 (N_5025,N_4813,N_4931);
nand U5026 (N_5026,N_4801,N_4760);
and U5027 (N_5027,N_4781,N_4987);
or U5028 (N_5028,N_4600,N_4576);
and U5029 (N_5029,N_4807,N_4997);
nor U5030 (N_5030,N_4632,N_4401);
nand U5031 (N_5031,N_4751,N_4968);
xor U5032 (N_5032,N_4529,N_4682);
or U5033 (N_5033,N_4809,N_4827);
nor U5034 (N_5034,N_4414,N_4718);
nor U5035 (N_5035,N_4746,N_4867);
or U5036 (N_5036,N_4664,N_4936);
nand U5037 (N_5037,N_4620,N_4730);
or U5038 (N_5038,N_4437,N_4767);
and U5039 (N_5039,N_4708,N_4646);
xnor U5040 (N_5040,N_4907,N_4754);
nor U5041 (N_5041,N_4772,N_4404);
and U5042 (N_5042,N_4421,N_4628);
or U5043 (N_5043,N_4728,N_4788);
and U5044 (N_5044,N_4970,N_4660);
or U5045 (N_5045,N_4474,N_4926);
nor U5046 (N_5046,N_4770,N_4740);
nor U5047 (N_5047,N_4555,N_4523);
or U5048 (N_5048,N_4651,N_4589);
nor U5049 (N_5049,N_4759,N_4377);
or U5050 (N_5050,N_4456,N_4899);
nand U5051 (N_5051,N_4532,N_4482);
and U5052 (N_5052,N_4983,N_4520);
and U5053 (N_5053,N_4443,N_4743);
or U5054 (N_5054,N_4550,N_4814);
nand U5055 (N_5055,N_4418,N_4783);
nand U5056 (N_5056,N_4854,N_4950);
nand U5057 (N_5057,N_4806,N_4613);
and U5058 (N_5058,N_4512,N_4614);
or U5059 (N_5059,N_4389,N_4541);
nand U5060 (N_5060,N_4775,N_4956);
and U5061 (N_5061,N_4624,N_4713);
and U5062 (N_5062,N_4489,N_4419);
nor U5063 (N_5063,N_4831,N_4859);
and U5064 (N_5064,N_4888,N_4724);
nand U5065 (N_5065,N_4438,N_4840);
nor U5066 (N_5066,N_4821,N_4451);
xor U5067 (N_5067,N_4923,N_4858);
or U5068 (N_5068,N_4659,N_4412);
and U5069 (N_5069,N_4988,N_4712);
nand U5070 (N_5070,N_4674,N_4804);
nor U5071 (N_5071,N_4929,N_4471);
and U5072 (N_5072,N_4979,N_4954);
or U5073 (N_5073,N_4617,N_4689);
nand U5074 (N_5074,N_4554,N_4459);
xnor U5075 (N_5075,N_4824,N_4846);
nand U5076 (N_5076,N_4974,N_4527);
or U5077 (N_5077,N_4839,N_4972);
and U5078 (N_5078,N_4667,N_4793);
and U5079 (N_5079,N_4588,N_4694);
nor U5080 (N_5080,N_4466,N_4477);
xor U5081 (N_5081,N_4887,N_4635);
or U5082 (N_5082,N_4995,N_4637);
and U5083 (N_5083,N_4593,N_4568);
or U5084 (N_5084,N_4745,N_4450);
nor U5085 (N_5085,N_4509,N_4756);
nor U5086 (N_5086,N_4861,N_4901);
and U5087 (N_5087,N_4462,N_4493);
or U5088 (N_5088,N_4436,N_4927);
and U5089 (N_5089,N_4710,N_4932);
or U5090 (N_5090,N_4940,N_4552);
nand U5091 (N_5091,N_4472,N_4490);
or U5092 (N_5092,N_4670,N_4590);
nor U5093 (N_5093,N_4794,N_4981);
or U5094 (N_5094,N_4883,N_4908);
nor U5095 (N_5095,N_4727,N_4431);
nor U5096 (N_5096,N_4508,N_4393);
xnor U5097 (N_5097,N_4557,N_4596);
nor U5098 (N_5098,N_4943,N_4764);
nand U5099 (N_5099,N_4582,N_4855);
nand U5100 (N_5100,N_4413,N_4871);
and U5101 (N_5101,N_4511,N_4882);
nor U5102 (N_5102,N_4469,N_4843);
xor U5103 (N_5103,N_4890,N_4734);
nand U5104 (N_5104,N_4623,N_4679);
and U5105 (N_5105,N_4542,N_4547);
xor U5106 (N_5106,N_4817,N_4597);
nand U5107 (N_5107,N_4748,N_4416);
or U5108 (N_5108,N_4953,N_4622);
and U5109 (N_5109,N_4969,N_4691);
nand U5110 (N_5110,N_4874,N_4941);
nand U5111 (N_5111,N_4828,N_4895);
nand U5112 (N_5112,N_4700,N_4429);
or U5113 (N_5113,N_4504,N_4709);
and U5114 (N_5114,N_4594,N_4584);
nand U5115 (N_5115,N_4722,N_4977);
xnor U5116 (N_5116,N_4787,N_4685);
nand U5117 (N_5117,N_4394,N_4612);
and U5118 (N_5118,N_4432,N_4440);
or U5119 (N_5119,N_4618,N_4385);
nand U5120 (N_5120,N_4522,N_4960);
and U5121 (N_5121,N_4869,N_4697);
xor U5122 (N_5122,N_4487,N_4765);
and U5123 (N_5123,N_4925,N_4980);
nand U5124 (N_5124,N_4841,N_4445);
nand U5125 (N_5125,N_4737,N_4938);
or U5126 (N_5126,N_4704,N_4497);
nor U5127 (N_5127,N_4833,N_4982);
nand U5128 (N_5128,N_4879,N_4711);
nor U5129 (N_5129,N_4836,N_4900);
and U5130 (N_5130,N_4399,N_4717);
or U5131 (N_5131,N_4777,N_4795);
nor U5132 (N_5132,N_4517,N_4905);
or U5133 (N_5133,N_4560,N_4857);
nor U5134 (N_5134,N_4897,N_4937);
nand U5135 (N_5135,N_4476,N_4848);
nand U5136 (N_5136,N_4894,N_4565);
nand U5137 (N_5137,N_4891,N_4629);
nand U5138 (N_5138,N_4725,N_4876);
and U5139 (N_5139,N_4766,N_4648);
xor U5140 (N_5140,N_4572,N_4716);
nor U5141 (N_5141,N_4942,N_4796);
nor U5142 (N_5142,N_4963,N_4898);
nor U5143 (N_5143,N_4702,N_4928);
nor U5144 (N_5144,N_4480,N_4672);
xor U5145 (N_5145,N_4731,N_4758);
and U5146 (N_5146,N_4407,N_4409);
nor U5147 (N_5147,N_4417,N_4516);
nor U5148 (N_5148,N_4993,N_4619);
nand U5149 (N_5149,N_4971,N_4381);
nand U5150 (N_5150,N_4973,N_4375);
and U5151 (N_5151,N_4992,N_4630);
nor U5152 (N_5152,N_4435,N_4473);
nand U5153 (N_5153,N_4615,N_4567);
or U5154 (N_5154,N_4696,N_4644);
nor U5155 (N_5155,N_4989,N_4998);
or U5156 (N_5156,N_4607,N_4608);
and U5157 (N_5157,N_4441,N_4881);
nand U5158 (N_5158,N_4442,N_4768);
or U5159 (N_5159,N_4699,N_4878);
and U5160 (N_5160,N_4778,N_4860);
and U5161 (N_5161,N_4934,N_4961);
nand U5162 (N_5162,N_4564,N_4653);
nand U5163 (N_5163,N_4738,N_4688);
and U5164 (N_5164,N_4591,N_4654);
and U5165 (N_5165,N_4657,N_4675);
or U5166 (N_5166,N_4822,N_4994);
and U5167 (N_5167,N_4687,N_4446);
nand U5168 (N_5168,N_4513,N_4403);
or U5169 (N_5169,N_4640,N_4884);
nand U5170 (N_5170,N_4524,N_4444);
nand U5171 (N_5171,N_4458,N_4551);
nand U5172 (N_5172,N_4483,N_4577);
and U5173 (N_5173,N_4433,N_4426);
or U5174 (N_5174,N_4396,N_4922);
or U5175 (N_5175,N_4605,N_4680);
xor U5176 (N_5176,N_4662,N_4815);
or U5177 (N_5177,N_4415,N_4539);
nand U5178 (N_5178,N_4604,N_4742);
xnor U5179 (N_5179,N_4499,N_4406);
or U5180 (N_5180,N_4427,N_4939);
nand U5181 (N_5181,N_4428,N_4966);
or U5182 (N_5182,N_4744,N_4677);
or U5183 (N_5183,N_4774,N_4505);
or U5184 (N_5184,N_4496,N_4634);
or U5185 (N_5185,N_4669,N_4475);
and U5186 (N_5186,N_4819,N_4515);
and U5187 (N_5187,N_4990,N_4453);
and U5188 (N_5188,N_4779,N_4769);
or U5189 (N_5189,N_4642,N_4510);
nand U5190 (N_5190,N_4703,N_4422);
or U5191 (N_5191,N_4818,N_4896);
nand U5192 (N_5192,N_4553,N_4918);
nand U5193 (N_5193,N_4780,N_4811);
xor U5194 (N_5194,N_4507,N_4917);
nand U5195 (N_5195,N_4959,N_4544);
nand U5196 (N_5196,N_4384,N_4603);
and U5197 (N_5197,N_4763,N_4837);
nand U5198 (N_5198,N_4569,N_4549);
nor U5199 (N_5199,N_4408,N_4581);
or U5200 (N_5200,N_4609,N_4639);
nand U5201 (N_5201,N_4506,N_4870);
or U5202 (N_5202,N_4964,N_4695);
nand U5203 (N_5203,N_4946,N_4559);
nor U5204 (N_5204,N_4531,N_4693);
or U5205 (N_5205,N_4601,N_4948);
and U5206 (N_5206,N_4518,N_4519);
nand U5207 (N_5207,N_4464,N_4457);
nor U5208 (N_5208,N_4985,N_4492);
nor U5209 (N_5209,N_4434,N_4430);
and U5210 (N_5210,N_4488,N_4666);
and U5211 (N_5211,N_4681,N_4800);
nor U5212 (N_5212,N_4398,N_4838);
nand U5213 (N_5213,N_4733,N_4991);
nand U5214 (N_5214,N_4752,N_4521);
nor U5215 (N_5215,N_4701,N_4784);
xor U5216 (N_5216,N_4829,N_4579);
nand U5217 (N_5217,N_4808,N_4892);
and U5218 (N_5218,N_4546,N_4465);
or U5219 (N_5219,N_4698,N_4835);
nand U5220 (N_5220,N_4706,N_4978);
or U5221 (N_5221,N_4984,N_4574);
or U5222 (N_5222,N_4545,N_4864);
nand U5223 (N_5223,N_4424,N_4949);
or U5224 (N_5224,N_4514,N_4755);
xnor U5225 (N_5225,N_4729,N_4944);
or U5226 (N_5226,N_4866,N_4911);
and U5227 (N_5227,N_4914,N_4735);
and U5228 (N_5228,N_4726,N_4606);
and U5229 (N_5229,N_4816,N_4665);
or U5230 (N_5230,N_4810,N_4877);
or U5231 (N_5231,N_4930,N_4636);
or U5232 (N_5232,N_4921,N_4916);
and U5233 (N_5233,N_4856,N_4425);
nor U5234 (N_5234,N_4376,N_4461);
xnor U5235 (N_5235,N_4955,N_4391);
xor U5236 (N_5236,N_4886,N_4478);
and U5237 (N_5237,N_4935,N_4655);
nand U5238 (N_5238,N_4500,N_4924);
xor U5239 (N_5239,N_4902,N_4562);
xor U5240 (N_5240,N_4535,N_4526);
nand U5241 (N_5241,N_4647,N_4986);
xor U5242 (N_5242,N_4671,N_4910);
xnor U5243 (N_5243,N_4958,N_4602);
and U5244 (N_5244,N_4598,N_4791);
and U5245 (N_5245,N_4739,N_4643);
and U5246 (N_5246,N_4873,N_4782);
and U5247 (N_5247,N_4631,N_4820);
and U5248 (N_5248,N_4397,N_4452);
and U5249 (N_5249,N_4789,N_4761);
and U5250 (N_5250,N_4537,N_4566);
and U5251 (N_5251,N_4379,N_4802);
or U5252 (N_5252,N_4797,N_4909);
and U5253 (N_5253,N_4919,N_4652);
nor U5254 (N_5254,N_4650,N_4868);
xor U5255 (N_5255,N_4952,N_4893);
nor U5256 (N_5256,N_4580,N_4904);
nor U5257 (N_5257,N_4656,N_4633);
nor U5258 (N_5258,N_4757,N_4498);
nand U5259 (N_5259,N_4420,N_4684);
and U5260 (N_5260,N_4673,N_4723);
nor U5261 (N_5261,N_4678,N_4962);
or U5262 (N_5262,N_4947,N_4915);
nor U5263 (N_5263,N_4690,N_4649);
or U5264 (N_5264,N_4851,N_4719);
nand U5265 (N_5265,N_4592,N_4720);
nor U5266 (N_5266,N_4996,N_4595);
or U5267 (N_5267,N_4558,N_4439);
nand U5268 (N_5268,N_4610,N_4885);
or U5269 (N_5269,N_4638,N_4741);
nor U5270 (N_5270,N_4543,N_4753);
nor U5271 (N_5271,N_4790,N_4454);
or U5272 (N_5272,N_4863,N_4786);
xor U5273 (N_5273,N_4383,N_4479);
xor U5274 (N_5274,N_4721,N_4561);
or U5275 (N_5275,N_4845,N_4852);
or U5276 (N_5276,N_4556,N_4749);
xor U5277 (N_5277,N_4792,N_4847);
xnor U5278 (N_5278,N_4715,N_4736);
or U5279 (N_5279,N_4773,N_4951);
or U5280 (N_5280,N_4903,N_4626);
xor U5281 (N_5281,N_4825,N_4750);
and U5282 (N_5282,N_4378,N_4460);
or U5283 (N_5283,N_4912,N_4494);
nand U5284 (N_5284,N_4799,N_4920);
and U5285 (N_5285,N_4641,N_4803);
or U5286 (N_5286,N_4405,N_4832);
and U5287 (N_5287,N_4448,N_4530);
nor U5288 (N_5288,N_4965,N_4798);
or U5289 (N_5289,N_4627,N_4776);
nor U5290 (N_5290,N_4826,N_4481);
and U5291 (N_5291,N_4470,N_4805);
nand U5292 (N_5292,N_4872,N_4616);
or U5293 (N_5293,N_4999,N_4468);
nor U5294 (N_5294,N_4395,N_4587);
nor U5295 (N_5295,N_4467,N_4540);
nor U5296 (N_5296,N_4485,N_4945);
and U5297 (N_5297,N_4661,N_4686);
or U5298 (N_5298,N_4563,N_4501);
nand U5299 (N_5299,N_4486,N_4853);
xor U5300 (N_5300,N_4683,N_4849);
nand U5301 (N_5301,N_4573,N_4386);
nor U5302 (N_5302,N_4411,N_4705);
xnor U5303 (N_5303,N_4447,N_4578);
nor U5304 (N_5304,N_4575,N_4906);
nand U5305 (N_5305,N_4692,N_4823);
nand U5306 (N_5306,N_4534,N_4583);
nor U5307 (N_5307,N_4571,N_4668);
and U5308 (N_5308,N_4714,N_4771);
nand U5309 (N_5309,N_4380,N_4423);
nand U5310 (N_5310,N_4570,N_4844);
and U5311 (N_5311,N_4707,N_4625);
xor U5312 (N_5312,N_4875,N_4896);
and U5313 (N_5313,N_4935,N_4688);
xor U5314 (N_5314,N_4446,N_4818);
nor U5315 (N_5315,N_4777,N_4418);
or U5316 (N_5316,N_4921,N_4509);
or U5317 (N_5317,N_4853,N_4651);
nand U5318 (N_5318,N_4885,N_4857);
or U5319 (N_5319,N_4453,N_4470);
nor U5320 (N_5320,N_4691,N_4769);
nand U5321 (N_5321,N_4416,N_4790);
or U5322 (N_5322,N_4936,N_4746);
and U5323 (N_5323,N_4448,N_4645);
and U5324 (N_5324,N_4939,N_4865);
xor U5325 (N_5325,N_4923,N_4870);
or U5326 (N_5326,N_4883,N_4380);
nand U5327 (N_5327,N_4707,N_4979);
nand U5328 (N_5328,N_4421,N_4862);
nand U5329 (N_5329,N_4959,N_4839);
and U5330 (N_5330,N_4968,N_4631);
or U5331 (N_5331,N_4388,N_4412);
xnor U5332 (N_5332,N_4403,N_4537);
nand U5333 (N_5333,N_4403,N_4961);
and U5334 (N_5334,N_4889,N_4548);
nand U5335 (N_5335,N_4662,N_4575);
nor U5336 (N_5336,N_4885,N_4805);
or U5337 (N_5337,N_4648,N_4710);
and U5338 (N_5338,N_4669,N_4741);
or U5339 (N_5339,N_4394,N_4922);
and U5340 (N_5340,N_4664,N_4634);
nor U5341 (N_5341,N_4419,N_4550);
nand U5342 (N_5342,N_4692,N_4979);
xor U5343 (N_5343,N_4582,N_4453);
and U5344 (N_5344,N_4802,N_4633);
and U5345 (N_5345,N_4405,N_4869);
or U5346 (N_5346,N_4795,N_4699);
and U5347 (N_5347,N_4772,N_4645);
and U5348 (N_5348,N_4898,N_4901);
nor U5349 (N_5349,N_4879,N_4530);
and U5350 (N_5350,N_4924,N_4979);
nand U5351 (N_5351,N_4479,N_4493);
nand U5352 (N_5352,N_4759,N_4990);
nand U5353 (N_5353,N_4406,N_4579);
or U5354 (N_5354,N_4984,N_4684);
and U5355 (N_5355,N_4773,N_4885);
and U5356 (N_5356,N_4995,N_4526);
nor U5357 (N_5357,N_4755,N_4722);
nor U5358 (N_5358,N_4729,N_4584);
and U5359 (N_5359,N_4451,N_4381);
and U5360 (N_5360,N_4617,N_4853);
nand U5361 (N_5361,N_4620,N_4933);
xnor U5362 (N_5362,N_4586,N_4709);
nor U5363 (N_5363,N_4439,N_4774);
nor U5364 (N_5364,N_4409,N_4514);
or U5365 (N_5365,N_4548,N_4383);
and U5366 (N_5366,N_4859,N_4567);
nand U5367 (N_5367,N_4523,N_4681);
or U5368 (N_5368,N_4589,N_4962);
xnor U5369 (N_5369,N_4855,N_4854);
nand U5370 (N_5370,N_4945,N_4386);
nand U5371 (N_5371,N_4578,N_4380);
or U5372 (N_5372,N_4506,N_4904);
or U5373 (N_5373,N_4694,N_4801);
xnor U5374 (N_5374,N_4964,N_4714);
nand U5375 (N_5375,N_4929,N_4615);
and U5376 (N_5376,N_4754,N_4903);
nand U5377 (N_5377,N_4414,N_4726);
or U5378 (N_5378,N_4376,N_4945);
nor U5379 (N_5379,N_4674,N_4685);
nor U5380 (N_5380,N_4421,N_4588);
nand U5381 (N_5381,N_4728,N_4438);
nand U5382 (N_5382,N_4636,N_4947);
nand U5383 (N_5383,N_4527,N_4886);
nand U5384 (N_5384,N_4960,N_4656);
nand U5385 (N_5385,N_4468,N_4449);
or U5386 (N_5386,N_4879,N_4976);
or U5387 (N_5387,N_4504,N_4382);
or U5388 (N_5388,N_4499,N_4457);
and U5389 (N_5389,N_4976,N_4592);
nor U5390 (N_5390,N_4375,N_4698);
and U5391 (N_5391,N_4438,N_4462);
and U5392 (N_5392,N_4404,N_4663);
nand U5393 (N_5393,N_4813,N_4799);
nor U5394 (N_5394,N_4416,N_4504);
nand U5395 (N_5395,N_4579,N_4776);
or U5396 (N_5396,N_4693,N_4505);
nor U5397 (N_5397,N_4842,N_4591);
nand U5398 (N_5398,N_4840,N_4873);
nand U5399 (N_5399,N_4824,N_4856);
and U5400 (N_5400,N_4504,N_4840);
and U5401 (N_5401,N_4997,N_4594);
nand U5402 (N_5402,N_4777,N_4804);
nand U5403 (N_5403,N_4811,N_4507);
and U5404 (N_5404,N_4393,N_4720);
nand U5405 (N_5405,N_4904,N_4993);
nand U5406 (N_5406,N_4607,N_4990);
nor U5407 (N_5407,N_4603,N_4590);
nand U5408 (N_5408,N_4810,N_4621);
xor U5409 (N_5409,N_4479,N_4719);
or U5410 (N_5410,N_4705,N_4828);
and U5411 (N_5411,N_4565,N_4469);
nand U5412 (N_5412,N_4983,N_4717);
xor U5413 (N_5413,N_4927,N_4977);
nor U5414 (N_5414,N_4943,N_4624);
and U5415 (N_5415,N_4721,N_4855);
nor U5416 (N_5416,N_4483,N_4840);
nor U5417 (N_5417,N_4805,N_4999);
and U5418 (N_5418,N_4493,N_4609);
and U5419 (N_5419,N_4538,N_4881);
nor U5420 (N_5420,N_4522,N_4375);
nor U5421 (N_5421,N_4603,N_4758);
xor U5422 (N_5422,N_4784,N_4943);
nand U5423 (N_5423,N_4717,N_4960);
and U5424 (N_5424,N_4819,N_4791);
and U5425 (N_5425,N_4977,N_4881);
or U5426 (N_5426,N_4865,N_4880);
nor U5427 (N_5427,N_4562,N_4901);
and U5428 (N_5428,N_4727,N_4782);
nand U5429 (N_5429,N_4978,N_4499);
and U5430 (N_5430,N_4412,N_4504);
or U5431 (N_5431,N_4792,N_4989);
and U5432 (N_5432,N_4404,N_4768);
nand U5433 (N_5433,N_4517,N_4688);
nand U5434 (N_5434,N_4907,N_4596);
nand U5435 (N_5435,N_4975,N_4611);
nor U5436 (N_5436,N_4884,N_4412);
nor U5437 (N_5437,N_4833,N_4682);
xnor U5438 (N_5438,N_4409,N_4948);
or U5439 (N_5439,N_4604,N_4769);
nand U5440 (N_5440,N_4403,N_4740);
or U5441 (N_5441,N_4791,N_4750);
or U5442 (N_5442,N_4924,N_4808);
or U5443 (N_5443,N_4845,N_4541);
nand U5444 (N_5444,N_4488,N_4910);
nand U5445 (N_5445,N_4602,N_4533);
or U5446 (N_5446,N_4593,N_4392);
nor U5447 (N_5447,N_4445,N_4464);
nor U5448 (N_5448,N_4382,N_4553);
nand U5449 (N_5449,N_4759,N_4869);
and U5450 (N_5450,N_4601,N_4469);
nand U5451 (N_5451,N_4486,N_4526);
nand U5452 (N_5452,N_4730,N_4537);
and U5453 (N_5453,N_4810,N_4494);
or U5454 (N_5454,N_4835,N_4379);
nor U5455 (N_5455,N_4702,N_4513);
nor U5456 (N_5456,N_4447,N_4600);
or U5457 (N_5457,N_4397,N_4976);
nand U5458 (N_5458,N_4746,N_4758);
nand U5459 (N_5459,N_4850,N_4547);
nor U5460 (N_5460,N_4505,N_4861);
nand U5461 (N_5461,N_4812,N_4935);
nand U5462 (N_5462,N_4708,N_4855);
nor U5463 (N_5463,N_4417,N_4472);
nand U5464 (N_5464,N_4618,N_4657);
or U5465 (N_5465,N_4861,N_4388);
xnor U5466 (N_5466,N_4946,N_4950);
and U5467 (N_5467,N_4526,N_4871);
nand U5468 (N_5468,N_4658,N_4666);
nand U5469 (N_5469,N_4586,N_4667);
or U5470 (N_5470,N_4972,N_4853);
or U5471 (N_5471,N_4800,N_4927);
or U5472 (N_5472,N_4629,N_4638);
and U5473 (N_5473,N_4890,N_4597);
nor U5474 (N_5474,N_4846,N_4655);
and U5475 (N_5475,N_4410,N_4689);
and U5476 (N_5476,N_4725,N_4952);
nand U5477 (N_5477,N_4754,N_4661);
and U5478 (N_5478,N_4382,N_4797);
nand U5479 (N_5479,N_4915,N_4684);
nor U5480 (N_5480,N_4658,N_4774);
or U5481 (N_5481,N_4612,N_4986);
and U5482 (N_5482,N_4590,N_4715);
or U5483 (N_5483,N_4774,N_4984);
and U5484 (N_5484,N_4537,N_4965);
nor U5485 (N_5485,N_4627,N_4826);
and U5486 (N_5486,N_4973,N_4634);
and U5487 (N_5487,N_4624,N_4494);
nand U5488 (N_5488,N_4579,N_4917);
xnor U5489 (N_5489,N_4588,N_4990);
nand U5490 (N_5490,N_4863,N_4423);
or U5491 (N_5491,N_4910,N_4853);
or U5492 (N_5492,N_4886,N_4392);
and U5493 (N_5493,N_4626,N_4761);
or U5494 (N_5494,N_4613,N_4785);
or U5495 (N_5495,N_4838,N_4780);
or U5496 (N_5496,N_4647,N_4866);
or U5497 (N_5497,N_4402,N_4978);
nor U5498 (N_5498,N_4552,N_4783);
and U5499 (N_5499,N_4936,N_4852);
nand U5500 (N_5500,N_4960,N_4750);
or U5501 (N_5501,N_4658,N_4791);
and U5502 (N_5502,N_4872,N_4765);
nand U5503 (N_5503,N_4627,N_4888);
nand U5504 (N_5504,N_4526,N_4831);
nor U5505 (N_5505,N_4948,N_4788);
nand U5506 (N_5506,N_4957,N_4616);
nand U5507 (N_5507,N_4581,N_4524);
nor U5508 (N_5508,N_4771,N_4890);
or U5509 (N_5509,N_4445,N_4480);
or U5510 (N_5510,N_4833,N_4495);
and U5511 (N_5511,N_4573,N_4667);
nand U5512 (N_5512,N_4430,N_4931);
nand U5513 (N_5513,N_4985,N_4445);
and U5514 (N_5514,N_4631,N_4889);
or U5515 (N_5515,N_4769,N_4856);
and U5516 (N_5516,N_4418,N_4528);
and U5517 (N_5517,N_4850,N_4859);
nor U5518 (N_5518,N_4562,N_4898);
or U5519 (N_5519,N_4861,N_4710);
nand U5520 (N_5520,N_4886,N_4717);
nand U5521 (N_5521,N_4788,N_4793);
nand U5522 (N_5522,N_4952,N_4896);
nor U5523 (N_5523,N_4684,N_4779);
and U5524 (N_5524,N_4429,N_4645);
or U5525 (N_5525,N_4453,N_4563);
nand U5526 (N_5526,N_4924,N_4845);
and U5527 (N_5527,N_4643,N_4621);
nand U5528 (N_5528,N_4681,N_4575);
xor U5529 (N_5529,N_4876,N_4459);
nor U5530 (N_5530,N_4515,N_4795);
nand U5531 (N_5531,N_4760,N_4472);
or U5532 (N_5532,N_4804,N_4975);
nand U5533 (N_5533,N_4775,N_4538);
xor U5534 (N_5534,N_4916,N_4521);
and U5535 (N_5535,N_4384,N_4667);
and U5536 (N_5536,N_4898,N_4988);
nand U5537 (N_5537,N_4408,N_4970);
or U5538 (N_5538,N_4879,N_4915);
nor U5539 (N_5539,N_4450,N_4602);
and U5540 (N_5540,N_4932,N_4892);
nor U5541 (N_5541,N_4846,N_4953);
and U5542 (N_5542,N_4929,N_4883);
xor U5543 (N_5543,N_4384,N_4784);
or U5544 (N_5544,N_4869,N_4955);
xnor U5545 (N_5545,N_4961,N_4512);
nor U5546 (N_5546,N_4726,N_4498);
nand U5547 (N_5547,N_4783,N_4497);
nor U5548 (N_5548,N_4444,N_4834);
and U5549 (N_5549,N_4739,N_4566);
nor U5550 (N_5550,N_4488,N_4832);
xnor U5551 (N_5551,N_4813,N_4671);
nor U5552 (N_5552,N_4378,N_4964);
or U5553 (N_5553,N_4868,N_4799);
or U5554 (N_5554,N_4525,N_4919);
or U5555 (N_5555,N_4752,N_4931);
nor U5556 (N_5556,N_4583,N_4978);
or U5557 (N_5557,N_4427,N_4665);
nand U5558 (N_5558,N_4743,N_4724);
or U5559 (N_5559,N_4814,N_4616);
or U5560 (N_5560,N_4429,N_4602);
nor U5561 (N_5561,N_4850,N_4770);
nor U5562 (N_5562,N_4401,N_4736);
nand U5563 (N_5563,N_4410,N_4904);
and U5564 (N_5564,N_4516,N_4495);
nor U5565 (N_5565,N_4837,N_4444);
and U5566 (N_5566,N_4633,N_4822);
or U5567 (N_5567,N_4455,N_4507);
nor U5568 (N_5568,N_4554,N_4907);
or U5569 (N_5569,N_4390,N_4709);
and U5570 (N_5570,N_4614,N_4469);
xnor U5571 (N_5571,N_4936,N_4445);
nand U5572 (N_5572,N_4799,N_4828);
nor U5573 (N_5573,N_4474,N_4588);
or U5574 (N_5574,N_4620,N_4482);
nor U5575 (N_5575,N_4708,N_4521);
xor U5576 (N_5576,N_4682,N_4379);
nand U5577 (N_5577,N_4964,N_4402);
and U5578 (N_5578,N_4574,N_4592);
and U5579 (N_5579,N_4945,N_4395);
nand U5580 (N_5580,N_4592,N_4605);
nor U5581 (N_5581,N_4527,N_4921);
nor U5582 (N_5582,N_4670,N_4721);
or U5583 (N_5583,N_4648,N_4772);
nand U5584 (N_5584,N_4424,N_4527);
nor U5585 (N_5585,N_4537,N_4377);
nand U5586 (N_5586,N_4759,N_4509);
or U5587 (N_5587,N_4482,N_4638);
and U5588 (N_5588,N_4615,N_4570);
and U5589 (N_5589,N_4448,N_4513);
nand U5590 (N_5590,N_4548,N_4402);
nand U5591 (N_5591,N_4844,N_4481);
or U5592 (N_5592,N_4986,N_4806);
nor U5593 (N_5593,N_4638,N_4646);
nand U5594 (N_5594,N_4986,N_4618);
and U5595 (N_5595,N_4953,N_4491);
nor U5596 (N_5596,N_4664,N_4748);
nor U5597 (N_5597,N_4506,N_4593);
nor U5598 (N_5598,N_4856,N_4758);
nand U5599 (N_5599,N_4591,N_4391);
nor U5600 (N_5600,N_4403,N_4785);
or U5601 (N_5601,N_4568,N_4429);
or U5602 (N_5602,N_4972,N_4832);
nand U5603 (N_5603,N_4475,N_4664);
or U5604 (N_5604,N_4695,N_4652);
nor U5605 (N_5605,N_4843,N_4479);
xor U5606 (N_5606,N_4739,N_4479);
and U5607 (N_5607,N_4834,N_4531);
nor U5608 (N_5608,N_4493,N_4522);
and U5609 (N_5609,N_4689,N_4604);
nand U5610 (N_5610,N_4813,N_4657);
nand U5611 (N_5611,N_4675,N_4711);
nor U5612 (N_5612,N_4975,N_4537);
or U5613 (N_5613,N_4942,N_4657);
nor U5614 (N_5614,N_4785,N_4713);
nor U5615 (N_5615,N_4656,N_4478);
or U5616 (N_5616,N_4658,N_4568);
xor U5617 (N_5617,N_4571,N_4756);
and U5618 (N_5618,N_4809,N_4402);
nand U5619 (N_5619,N_4736,N_4650);
or U5620 (N_5620,N_4861,N_4719);
nor U5621 (N_5621,N_4638,N_4949);
and U5622 (N_5622,N_4740,N_4725);
or U5623 (N_5623,N_4964,N_4464);
nand U5624 (N_5624,N_4571,N_4663);
or U5625 (N_5625,N_5107,N_5022);
nor U5626 (N_5626,N_5204,N_5350);
nor U5627 (N_5627,N_5331,N_5037);
and U5628 (N_5628,N_5384,N_5122);
or U5629 (N_5629,N_5285,N_5611);
or U5630 (N_5630,N_5024,N_5007);
or U5631 (N_5631,N_5262,N_5547);
nand U5632 (N_5632,N_5282,N_5571);
and U5633 (N_5633,N_5517,N_5556);
and U5634 (N_5634,N_5102,N_5187);
nor U5635 (N_5635,N_5238,N_5164);
and U5636 (N_5636,N_5562,N_5377);
and U5637 (N_5637,N_5396,N_5539);
or U5638 (N_5638,N_5463,N_5503);
nand U5639 (N_5639,N_5106,N_5074);
or U5640 (N_5640,N_5067,N_5128);
nor U5641 (N_5641,N_5297,N_5251);
and U5642 (N_5642,N_5118,N_5121);
nor U5643 (N_5643,N_5245,N_5335);
and U5644 (N_5644,N_5197,N_5445);
and U5645 (N_5645,N_5340,N_5530);
and U5646 (N_5646,N_5097,N_5048);
and U5647 (N_5647,N_5192,N_5129);
nor U5648 (N_5648,N_5535,N_5100);
nand U5649 (N_5649,N_5580,N_5230);
or U5650 (N_5650,N_5378,N_5143);
nand U5651 (N_5651,N_5462,N_5249);
nand U5652 (N_5652,N_5042,N_5587);
nand U5653 (N_5653,N_5555,N_5055);
and U5654 (N_5654,N_5582,N_5290);
and U5655 (N_5655,N_5438,N_5273);
and U5656 (N_5656,N_5542,N_5295);
or U5657 (N_5657,N_5259,N_5479);
nor U5658 (N_5658,N_5554,N_5172);
nor U5659 (N_5659,N_5306,N_5513);
and U5660 (N_5660,N_5344,N_5418);
xor U5661 (N_5661,N_5237,N_5575);
xnor U5662 (N_5662,N_5144,N_5054);
or U5663 (N_5663,N_5537,N_5491);
nand U5664 (N_5664,N_5454,N_5028);
xnor U5665 (N_5665,N_5349,N_5221);
xnor U5666 (N_5666,N_5576,N_5293);
or U5667 (N_5667,N_5526,N_5521);
or U5668 (N_5668,N_5601,N_5207);
nand U5669 (N_5669,N_5011,N_5534);
nand U5670 (N_5670,N_5206,N_5577);
nand U5671 (N_5671,N_5501,N_5313);
or U5672 (N_5672,N_5023,N_5317);
nor U5673 (N_5673,N_5281,N_5390);
nand U5674 (N_5674,N_5400,N_5280);
and U5675 (N_5675,N_5073,N_5568);
and U5676 (N_5676,N_5613,N_5357);
nand U5677 (N_5677,N_5508,N_5433);
xor U5678 (N_5678,N_5415,N_5602);
or U5679 (N_5679,N_5242,N_5525);
nor U5680 (N_5680,N_5296,N_5442);
and U5681 (N_5681,N_5600,N_5307);
nand U5682 (N_5682,N_5138,N_5116);
and U5683 (N_5683,N_5447,N_5234);
nor U5684 (N_5684,N_5361,N_5607);
nand U5685 (N_5685,N_5149,N_5132);
or U5686 (N_5686,N_5228,N_5165);
nor U5687 (N_5687,N_5174,N_5435);
nand U5688 (N_5688,N_5374,N_5599);
and U5689 (N_5689,N_5471,N_5021);
nand U5690 (N_5690,N_5189,N_5170);
or U5691 (N_5691,N_5423,N_5617);
or U5692 (N_5692,N_5597,N_5026);
and U5693 (N_5693,N_5289,N_5137);
and U5694 (N_5694,N_5009,N_5522);
or U5695 (N_5695,N_5232,N_5548);
or U5696 (N_5696,N_5181,N_5581);
and U5697 (N_5697,N_5298,N_5618);
nand U5698 (N_5698,N_5510,N_5010);
or U5699 (N_5699,N_5115,N_5446);
or U5700 (N_5700,N_5397,N_5443);
nor U5701 (N_5701,N_5236,N_5032);
and U5702 (N_5702,N_5001,N_5588);
xor U5703 (N_5703,N_5058,N_5202);
nand U5704 (N_5704,N_5018,N_5586);
nand U5705 (N_5705,N_5255,N_5185);
xor U5706 (N_5706,N_5531,N_5388);
nand U5707 (N_5707,N_5403,N_5252);
or U5708 (N_5708,N_5612,N_5362);
or U5709 (N_5709,N_5019,N_5482);
and U5710 (N_5710,N_5220,N_5099);
and U5711 (N_5711,N_5090,N_5416);
nor U5712 (N_5712,N_5399,N_5379);
nor U5713 (N_5713,N_5258,N_5040);
and U5714 (N_5714,N_5474,N_5114);
or U5715 (N_5715,N_5142,N_5124);
nor U5716 (N_5716,N_5079,N_5434);
and U5717 (N_5717,N_5034,N_5260);
xor U5718 (N_5718,N_5241,N_5188);
nor U5719 (N_5719,N_5466,N_5327);
and U5720 (N_5720,N_5359,N_5615);
nor U5721 (N_5721,N_5406,N_5609);
and U5722 (N_5722,N_5459,N_5421);
xnor U5723 (N_5723,N_5225,N_5093);
nor U5724 (N_5724,N_5256,N_5419);
or U5725 (N_5725,N_5385,N_5081);
or U5726 (N_5726,N_5348,N_5027);
and U5727 (N_5727,N_5215,N_5287);
nor U5728 (N_5728,N_5593,N_5005);
and U5729 (N_5729,N_5218,N_5614);
nor U5730 (N_5730,N_5578,N_5590);
and U5731 (N_5731,N_5227,N_5622);
nand U5732 (N_5732,N_5536,N_5383);
or U5733 (N_5733,N_5217,N_5325);
nand U5734 (N_5734,N_5239,N_5201);
or U5735 (N_5735,N_5305,N_5523);
nor U5736 (N_5736,N_5092,N_5150);
nand U5737 (N_5737,N_5050,N_5567);
and U5738 (N_5738,N_5069,N_5473);
or U5739 (N_5739,N_5498,N_5288);
nor U5740 (N_5740,N_5095,N_5179);
nand U5741 (N_5741,N_5424,N_5038);
nor U5742 (N_5742,N_5004,N_5075);
nand U5743 (N_5743,N_5047,N_5098);
and U5744 (N_5744,N_5518,N_5504);
xnor U5745 (N_5745,N_5162,N_5332);
nand U5746 (N_5746,N_5180,N_5169);
and U5747 (N_5747,N_5389,N_5088);
nor U5748 (N_5748,N_5353,N_5279);
nor U5749 (N_5749,N_5452,N_5065);
or U5750 (N_5750,N_5546,N_5564);
nand U5751 (N_5751,N_5541,N_5569);
or U5752 (N_5752,N_5440,N_5141);
or U5753 (N_5753,N_5254,N_5292);
and U5754 (N_5754,N_5222,N_5152);
nand U5755 (N_5755,N_5291,N_5064);
nor U5756 (N_5756,N_5008,N_5184);
xor U5757 (N_5757,N_5084,N_5270);
and U5758 (N_5758,N_5229,N_5351);
nor U5759 (N_5759,N_5060,N_5369);
nor U5760 (N_5760,N_5319,N_5465);
xnor U5761 (N_5761,N_5328,N_5366);
xor U5762 (N_5762,N_5493,N_5467);
nand U5763 (N_5763,N_5338,N_5085);
nand U5764 (N_5764,N_5014,N_5551);
nor U5765 (N_5765,N_5136,N_5127);
nand U5766 (N_5766,N_5515,N_5087);
or U5767 (N_5767,N_5528,N_5553);
and U5768 (N_5768,N_5373,N_5425);
nor U5769 (N_5769,N_5082,N_5314);
nor U5770 (N_5770,N_5043,N_5096);
and U5771 (N_5771,N_5158,N_5456);
or U5772 (N_5772,N_5382,N_5190);
nor U5773 (N_5773,N_5484,N_5550);
xnor U5774 (N_5774,N_5233,N_5231);
and U5775 (N_5775,N_5439,N_5160);
xor U5776 (N_5776,N_5140,N_5604);
nand U5777 (N_5777,N_5409,N_5046);
nand U5778 (N_5778,N_5219,N_5131);
and U5779 (N_5779,N_5594,N_5310);
or U5780 (N_5780,N_5346,N_5364);
nand U5781 (N_5781,N_5111,N_5312);
nor U5782 (N_5782,N_5352,N_5616);
nor U5783 (N_5783,N_5015,N_5422);
xnor U5784 (N_5784,N_5066,N_5372);
nand U5785 (N_5785,N_5560,N_5248);
or U5786 (N_5786,N_5476,N_5605);
or U5787 (N_5787,N_5608,N_5566);
or U5788 (N_5788,N_5450,N_5412);
nand U5789 (N_5789,N_5246,N_5516);
nand U5790 (N_5790,N_5025,N_5119);
nand U5791 (N_5791,N_5529,N_5205);
xor U5792 (N_5792,N_5276,N_5078);
or U5793 (N_5793,N_5483,N_5355);
or U5794 (N_5794,N_5458,N_5303);
and U5795 (N_5795,N_5570,N_5367);
xnor U5796 (N_5796,N_5300,N_5193);
or U5797 (N_5797,N_5156,N_5544);
nand U5798 (N_5798,N_5591,N_5035);
nand U5799 (N_5799,N_5153,N_5370);
xor U5800 (N_5800,N_5196,N_5126);
nand U5801 (N_5801,N_5134,N_5485);
nor U5802 (N_5802,N_5360,N_5089);
and U5803 (N_5803,N_5371,N_5395);
xor U5804 (N_5804,N_5182,N_5545);
nor U5805 (N_5805,N_5059,N_5203);
nand U5806 (N_5806,N_5146,N_5414);
nor U5807 (N_5807,N_5509,N_5572);
and U5808 (N_5808,N_5016,N_5387);
or U5809 (N_5809,N_5320,N_5457);
nand U5810 (N_5810,N_5573,N_5003);
or U5811 (N_5811,N_5363,N_5062);
xnor U5812 (N_5812,N_5514,N_5557);
nor U5813 (N_5813,N_5243,N_5226);
nor U5814 (N_5814,N_5077,N_5053);
nand U5815 (N_5815,N_5033,N_5481);
nor U5816 (N_5816,N_5444,N_5552);
nand U5817 (N_5817,N_5343,N_5497);
nor U5818 (N_5818,N_5441,N_5558);
or U5819 (N_5819,N_5209,N_5175);
or U5820 (N_5820,N_5268,N_5049);
nand U5821 (N_5821,N_5208,N_5155);
and U5822 (N_5822,N_5235,N_5502);
nor U5823 (N_5823,N_5480,N_5284);
and U5824 (N_5824,N_5091,N_5506);
or U5825 (N_5825,N_5341,N_5068);
or U5826 (N_5826,N_5329,N_5430);
nand U5827 (N_5827,N_5437,N_5365);
nor U5828 (N_5828,N_5533,N_5511);
xor U5829 (N_5829,N_5133,N_5606);
and U5830 (N_5830,N_5147,N_5030);
nand U5831 (N_5831,N_5486,N_5342);
nor U5832 (N_5832,N_5318,N_5505);
or U5833 (N_5833,N_5448,N_5210);
or U5834 (N_5834,N_5247,N_5411);
and U5835 (N_5835,N_5186,N_5080);
nor U5836 (N_5836,N_5212,N_5157);
nand U5837 (N_5837,N_5145,N_5094);
or U5838 (N_5838,N_5417,N_5358);
and U5839 (N_5839,N_5451,N_5161);
nor U5840 (N_5840,N_5103,N_5316);
nor U5841 (N_5841,N_5330,N_5354);
or U5842 (N_5842,N_5076,N_5431);
nand U5843 (N_5843,N_5519,N_5408);
nor U5844 (N_5844,N_5272,N_5393);
and U5845 (N_5845,N_5490,N_5002);
or U5846 (N_5846,N_5407,N_5083);
nand U5847 (N_5847,N_5006,N_5176);
and U5848 (N_5848,N_5278,N_5455);
or U5849 (N_5849,N_5478,N_5264);
nand U5850 (N_5850,N_5195,N_5598);
or U5851 (N_5851,N_5427,N_5151);
and U5852 (N_5852,N_5286,N_5429);
xor U5853 (N_5853,N_5211,N_5624);
nand U5854 (N_5854,N_5214,N_5584);
xnor U5855 (N_5855,N_5391,N_5428);
nor U5856 (N_5856,N_5610,N_5333);
and U5857 (N_5857,N_5347,N_5200);
nand U5858 (N_5858,N_5583,N_5585);
nand U5859 (N_5859,N_5420,N_5271);
and U5860 (N_5860,N_5269,N_5257);
nand U5861 (N_5861,N_5470,N_5168);
or U5862 (N_5862,N_5167,N_5380);
or U5863 (N_5863,N_5563,N_5324);
nand U5864 (N_5864,N_5125,N_5031);
xnor U5865 (N_5865,N_5299,N_5426);
or U5866 (N_5866,N_5520,N_5063);
xor U5867 (N_5867,N_5244,N_5477);
or U5868 (N_5868,N_5250,N_5579);
nand U5869 (N_5869,N_5339,N_5178);
nor U5870 (N_5870,N_5507,N_5592);
nand U5871 (N_5871,N_5392,N_5159);
nor U5872 (N_5872,N_5436,N_5620);
xor U5873 (N_5873,N_5540,N_5274);
nand U5874 (N_5874,N_5275,N_5044);
nand U5875 (N_5875,N_5216,N_5213);
nand U5876 (N_5876,N_5561,N_5224);
nand U5877 (N_5877,N_5029,N_5139);
nand U5878 (N_5878,N_5086,N_5623);
and U5879 (N_5879,N_5494,N_5301);
nand U5880 (N_5880,N_5148,N_5401);
and U5881 (N_5881,N_5398,N_5051);
or U5882 (N_5882,N_5461,N_5194);
nor U5883 (N_5883,N_5512,N_5302);
nand U5884 (N_5884,N_5596,N_5071);
and U5885 (N_5885,N_5120,N_5460);
or U5886 (N_5886,N_5135,N_5311);
and U5887 (N_5887,N_5163,N_5012);
or U5888 (N_5888,N_5041,N_5277);
nand U5889 (N_5889,N_5595,N_5070);
xnor U5890 (N_5890,N_5110,N_5402);
nand U5891 (N_5891,N_5253,N_5199);
and U5892 (N_5892,N_5045,N_5112);
and U5893 (N_5893,N_5294,N_5171);
and U5894 (N_5894,N_5173,N_5117);
or U5895 (N_5895,N_5105,N_5489);
nor U5896 (N_5896,N_5057,N_5017);
and U5897 (N_5897,N_5375,N_5404);
nand U5898 (N_5898,N_5527,N_5464);
or U5899 (N_5899,N_5321,N_5410);
nor U5900 (N_5900,N_5052,N_5472);
and U5901 (N_5901,N_5223,N_5265);
nand U5902 (N_5902,N_5496,N_5589);
nand U5903 (N_5903,N_5309,N_5240);
or U5904 (N_5904,N_5532,N_5113);
nand U5905 (N_5905,N_5376,N_5261);
and U5906 (N_5906,N_5322,N_5315);
nor U5907 (N_5907,N_5565,N_5323);
nand U5908 (N_5908,N_5267,N_5283);
nor U5909 (N_5909,N_5499,N_5559);
nor U5910 (N_5910,N_5381,N_5108);
and U5911 (N_5911,N_5345,N_5039);
xor U5912 (N_5912,N_5072,N_5475);
and U5913 (N_5913,N_5000,N_5154);
nor U5914 (N_5914,N_5020,N_5101);
or U5915 (N_5915,N_5334,N_5619);
nand U5916 (N_5916,N_5621,N_5574);
or U5917 (N_5917,N_5336,N_5356);
xnor U5918 (N_5918,N_5500,N_5266);
or U5919 (N_5919,N_5538,N_5432);
or U5920 (N_5920,N_5326,N_5337);
or U5921 (N_5921,N_5386,N_5549);
nor U5922 (N_5922,N_5198,N_5394);
nand U5923 (N_5923,N_5603,N_5191);
xor U5924 (N_5924,N_5413,N_5109);
and U5925 (N_5925,N_5013,N_5130);
nor U5926 (N_5926,N_5308,N_5449);
nor U5927 (N_5927,N_5487,N_5056);
xnor U5928 (N_5928,N_5123,N_5543);
or U5929 (N_5929,N_5061,N_5104);
or U5930 (N_5930,N_5495,N_5304);
or U5931 (N_5931,N_5468,N_5166);
nand U5932 (N_5932,N_5524,N_5263);
and U5933 (N_5933,N_5405,N_5036);
and U5934 (N_5934,N_5488,N_5469);
or U5935 (N_5935,N_5177,N_5368);
xnor U5936 (N_5936,N_5492,N_5183);
nor U5937 (N_5937,N_5453,N_5256);
nand U5938 (N_5938,N_5036,N_5327);
and U5939 (N_5939,N_5390,N_5413);
nor U5940 (N_5940,N_5153,N_5301);
or U5941 (N_5941,N_5437,N_5454);
or U5942 (N_5942,N_5298,N_5174);
and U5943 (N_5943,N_5324,N_5198);
or U5944 (N_5944,N_5556,N_5109);
xor U5945 (N_5945,N_5025,N_5456);
nand U5946 (N_5946,N_5414,N_5188);
nor U5947 (N_5947,N_5504,N_5533);
nand U5948 (N_5948,N_5613,N_5099);
and U5949 (N_5949,N_5302,N_5572);
or U5950 (N_5950,N_5137,N_5550);
or U5951 (N_5951,N_5302,N_5381);
nand U5952 (N_5952,N_5523,N_5088);
nand U5953 (N_5953,N_5506,N_5443);
nor U5954 (N_5954,N_5495,N_5001);
xnor U5955 (N_5955,N_5412,N_5241);
and U5956 (N_5956,N_5023,N_5464);
nand U5957 (N_5957,N_5064,N_5489);
nand U5958 (N_5958,N_5416,N_5513);
and U5959 (N_5959,N_5332,N_5156);
nand U5960 (N_5960,N_5086,N_5612);
nor U5961 (N_5961,N_5290,N_5466);
or U5962 (N_5962,N_5570,N_5258);
or U5963 (N_5963,N_5444,N_5203);
and U5964 (N_5964,N_5115,N_5118);
and U5965 (N_5965,N_5076,N_5492);
nand U5966 (N_5966,N_5594,N_5385);
or U5967 (N_5967,N_5205,N_5296);
or U5968 (N_5968,N_5195,N_5407);
and U5969 (N_5969,N_5473,N_5439);
nand U5970 (N_5970,N_5319,N_5208);
and U5971 (N_5971,N_5041,N_5535);
xor U5972 (N_5972,N_5608,N_5516);
nor U5973 (N_5973,N_5303,N_5375);
nand U5974 (N_5974,N_5536,N_5296);
and U5975 (N_5975,N_5428,N_5596);
or U5976 (N_5976,N_5583,N_5276);
xnor U5977 (N_5977,N_5085,N_5480);
and U5978 (N_5978,N_5395,N_5049);
and U5979 (N_5979,N_5136,N_5258);
nor U5980 (N_5980,N_5422,N_5173);
and U5981 (N_5981,N_5015,N_5049);
nor U5982 (N_5982,N_5477,N_5539);
or U5983 (N_5983,N_5218,N_5473);
nand U5984 (N_5984,N_5278,N_5381);
and U5985 (N_5985,N_5510,N_5576);
or U5986 (N_5986,N_5249,N_5421);
and U5987 (N_5987,N_5245,N_5424);
nand U5988 (N_5988,N_5214,N_5416);
nand U5989 (N_5989,N_5068,N_5448);
nor U5990 (N_5990,N_5554,N_5324);
or U5991 (N_5991,N_5282,N_5056);
nor U5992 (N_5992,N_5217,N_5187);
nor U5993 (N_5993,N_5387,N_5429);
and U5994 (N_5994,N_5508,N_5494);
and U5995 (N_5995,N_5122,N_5281);
nor U5996 (N_5996,N_5198,N_5056);
nand U5997 (N_5997,N_5205,N_5372);
nand U5998 (N_5998,N_5620,N_5606);
and U5999 (N_5999,N_5320,N_5397);
nor U6000 (N_6000,N_5398,N_5550);
xor U6001 (N_6001,N_5057,N_5040);
or U6002 (N_6002,N_5455,N_5045);
xor U6003 (N_6003,N_5071,N_5113);
nor U6004 (N_6004,N_5620,N_5094);
nand U6005 (N_6005,N_5478,N_5589);
nor U6006 (N_6006,N_5520,N_5325);
and U6007 (N_6007,N_5602,N_5615);
nand U6008 (N_6008,N_5006,N_5054);
nor U6009 (N_6009,N_5042,N_5521);
and U6010 (N_6010,N_5551,N_5458);
and U6011 (N_6011,N_5373,N_5214);
xnor U6012 (N_6012,N_5276,N_5060);
or U6013 (N_6013,N_5476,N_5155);
xor U6014 (N_6014,N_5111,N_5457);
or U6015 (N_6015,N_5566,N_5124);
or U6016 (N_6016,N_5094,N_5313);
xnor U6017 (N_6017,N_5439,N_5352);
nand U6018 (N_6018,N_5295,N_5339);
nand U6019 (N_6019,N_5469,N_5472);
nand U6020 (N_6020,N_5525,N_5495);
and U6021 (N_6021,N_5609,N_5322);
and U6022 (N_6022,N_5000,N_5106);
or U6023 (N_6023,N_5234,N_5108);
nor U6024 (N_6024,N_5156,N_5515);
and U6025 (N_6025,N_5277,N_5025);
or U6026 (N_6026,N_5209,N_5546);
or U6027 (N_6027,N_5410,N_5419);
nand U6028 (N_6028,N_5552,N_5434);
xor U6029 (N_6029,N_5133,N_5439);
nand U6030 (N_6030,N_5356,N_5067);
or U6031 (N_6031,N_5277,N_5404);
or U6032 (N_6032,N_5432,N_5330);
xnor U6033 (N_6033,N_5370,N_5272);
nand U6034 (N_6034,N_5526,N_5345);
and U6035 (N_6035,N_5040,N_5365);
nor U6036 (N_6036,N_5601,N_5497);
nor U6037 (N_6037,N_5032,N_5581);
nand U6038 (N_6038,N_5252,N_5374);
or U6039 (N_6039,N_5139,N_5000);
nand U6040 (N_6040,N_5191,N_5561);
nor U6041 (N_6041,N_5017,N_5493);
nand U6042 (N_6042,N_5030,N_5443);
xor U6043 (N_6043,N_5035,N_5601);
nor U6044 (N_6044,N_5135,N_5488);
or U6045 (N_6045,N_5258,N_5194);
or U6046 (N_6046,N_5337,N_5010);
nand U6047 (N_6047,N_5362,N_5150);
or U6048 (N_6048,N_5049,N_5123);
or U6049 (N_6049,N_5334,N_5067);
or U6050 (N_6050,N_5143,N_5131);
or U6051 (N_6051,N_5120,N_5116);
nand U6052 (N_6052,N_5500,N_5590);
and U6053 (N_6053,N_5130,N_5335);
xor U6054 (N_6054,N_5422,N_5124);
nand U6055 (N_6055,N_5418,N_5302);
xnor U6056 (N_6056,N_5006,N_5574);
or U6057 (N_6057,N_5233,N_5076);
and U6058 (N_6058,N_5184,N_5467);
or U6059 (N_6059,N_5053,N_5607);
nand U6060 (N_6060,N_5373,N_5259);
nand U6061 (N_6061,N_5108,N_5362);
nand U6062 (N_6062,N_5366,N_5521);
nand U6063 (N_6063,N_5247,N_5600);
and U6064 (N_6064,N_5382,N_5163);
nor U6065 (N_6065,N_5224,N_5347);
or U6066 (N_6066,N_5352,N_5236);
or U6067 (N_6067,N_5533,N_5536);
nand U6068 (N_6068,N_5274,N_5292);
and U6069 (N_6069,N_5518,N_5181);
nand U6070 (N_6070,N_5480,N_5610);
and U6071 (N_6071,N_5196,N_5149);
nand U6072 (N_6072,N_5164,N_5121);
or U6073 (N_6073,N_5468,N_5250);
and U6074 (N_6074,N_5461,N_5065);
nor U6075 (N_6075,N_5320,N_5383);
or U6076 (N_6076,N_5335,N_5235);
and U6077 (N_6077,N_5011,N_5351);
nand U6078 (N_6078,N_5416,N_5064);
nor U6079 (N_6079,N_5467,N_5078);
nor U6080 (N_6080,N_5409,N_5326);
and U6081 (N_6081,N_5227,N_5384);
or U6082 (N_6082,N_5260,N_5370);
or U6083 (N_6083,N_5412,N_5305);
or U6084 (N_6084,N_5114,N_5334);
nor U6085 (N_6085,N_5444,N_5150);
nor U6086 (N_6086,N_5062,N_5496);
and U6087 (N_6087,N_5014,N_5443);
nor U6088 (N_6088,N_5410,N_5536);
or U6089 (N_6089,N_5144,N_5418);
and U6090 (N_6090,N_5403,N_5364);
and U6091 (N_6091,N_5254,N_5476);
and U6092 (N_6092,N_5208,N_5176);
nor U6093 (N_6093,N_5552,N_5318);
nand U6094 (N_6094,N_5145,N_5039);
nor U6095 (N_6095,N_5510,N_5501);
nor U6096 (N_6096,N_5273,N_5069);
xnor U6097 (N_6097,N_5353,N_5123);
or U6098 (N_6098,N_5543,N_5312);
and U6099 (N_6099,N_5250,N_5261);
nand U6100 (N_6100,N_5309,N_5543);
nand U6101 (N_6101,N_5015,N_5362);
and U6102 (N_6102,N_5606,N_5103);
nor U6103 (N_6103,N_5614,N_5138);
and U6104 (N_6104,N_5098,N_5545);
nand U6105 (N_6105,N_5042,N_5130);
and U6106 (N_6106,N_5428,N_5059);
nor U6107 (N_6107,N_5429,N_5006);
and U6108 (N_6108,N_5199,N_5523);
or U6109 (N_6109,N_5100,N_5417);
nand U6110 (N_6110,N_5311,N_5557);
nand U6111 (N_6111,N_5310,N_5313);
and U6112 (N_6112,N_5477,N_5499);
nor U6113 (N_6113,N_5374,N_5291);
nor U6114 (N_6114,N_5259,N_5351);
or U6115 (N_6115,N_5619,N_5206);
and U6116 (N_6116,N_5151,N_5576);
or U6117 (N_6117,N_5038,N_5142);
nand U6118 (N_6118,N_5620,N_5061);
and U6119 (N_6119,N_5014,N_5472);
nor U6120 (N_6120,N_5442,N_5509);
nor U6121 (N_6121,N_5218,N_5423);
or U6122 (N_6122,N_5567,N_5341);
nand U6123 (N_6123,N_5480,N_5140);
nand U6124 (N_6124,N_5440,N_5246);
nand U6125 (N_6125,N_5421,N_5102);
nand U6126 (N_6126,N_5213,N_5324);
and U6127 (N_6127,N_5374,N_5595);
xnor U6128 (N_6128,N_5093,N_5061);
or U6129 (N_6129,N_5585,N_5212);
xor U6130 (N_6130,N_5082,N_5208);
or U6131 (N_6131,N_5444,N_5168);
nand U6132 (N_6132,N_5359,N_5256);
and U6133 (N_6133,N_5212,N_5269);
nor U6134 (N_6134,N_5454,N_5104);
nor U6135 (N_6135,N_5620,N_5011);
and U6136 (N_6136,N_5057,N_5380);
nand U6137 (N_6137,N_5117,N_5433);
or U6138 (N_6138,N_5120,N_5274);
nor U6139 (N_6139,N_5524,N_5366);
nor U6140 (N_6140,N_5518,N_5559);
nor U6141 (N_6141,N_5260,N_5242);
nand U6142 (N_6142,N_5616,N_5419);
nor U6143 (N_6143,N_5280,N_5567);
and U6144 (N_6144,N_5541,N_5377);
and U6145 (N_6145,N_5614,N_5455);
nand U6146 (N_6146,N_5348,N_5501);
nor U6147 (N_6147,N_5595,N_5001);
nand U6148 (N_6148,N_5487,N_5094);
nand U6149 (N_6149,N_5038,N_5012);
nor U6150 (N_6150,N_5314,N_5403);
nor U6151 (N_6151,N_5158,N_5201);
nor U6152 (N_6152,N_5275,N_5364);
nor U6153 (N_6153,N_5552,N_5148);
and U6154 (N_6154,N_5288,N_5121);
and U6155 (N_6155,N_5578,N_5183);
and U6156 (N_6156,N_5020,N_5276);
or U6157 (N_6157,N_5105,N_5400);
nand U6158 (N_6158,N_5257,N_5051);
nand U6159 (N_6159,N_5382,N_5503);
nand U6160 (N_6160,N_5153,N_5148);
and U6161 (N_6161,N_5509,N_5575);
or U6162 (N_6162,N_5517,N_5386);
and U6163 (N_6163,N_5413,N_5252);
nand U6164 (N_6164,N_5155,N_5296);
nor U6165 (N_6165,N_5454,N_5275);
nor U6166 (N_6166,N_5289,N_5028);
or U6167 (N_6167,N_5276,N_5403);
or U6168 (N_6168,N_5166,N_5473);
or U6169 (N_6169,N_5362,N_5158);
or U6170 (N_6170,N_5002,N_5468);
nand U6171 (N_6171,N_5427,N_5039);
nor U6172 (N_6172,N_5243,N_5170);
nor U6173 (N_6173,N_5350,N_5422);
nor U6174 (N_6174,N_5261,N_5421);
and U6175 (N_6175,N_5574,N_5604);
or U6176 (N_6176,N_5247,N_5395);
and U6177 (N_6177,N_5316,N_5517);
nand U6178 (N_6178,N_5455,N_5081);
and U6179 (N_6179,N_5608,N_5613);
xor U6180 (N_6180,N_5151,N_5368);
xor U6181 (N_6181,N_5210,N_5374);
or U6182 (N_6182,N_5336,N_5130);
nand U6183 (N_6183,N_5497,N_5174);
nand U6184 (N_6184,N_5204,N_5037);
nor U6185 (N_6185,N_5478,N_5508);
nand U6186 (N_6186,N_5230,N_5028);
or U6187 (N_6187,N_5376,N_5160);
nand U6188 (N_6188,N_5529,N_5335);
or U6189 (N_6189,N_5089,N_5134);
or U6190 (N_6190,N_5182,N_5018);
nor U6191 (N_6191,N_5289,N_5412);
nand U6192 (N_6192,N_5339,N_5399);
nor U6193 (N_6193,N_5385,N_5359);
or U6194 (N_6194,N_5220,N_5247);
and U6195 (N_6195,N_5304,N_5573);
or U6196 (N_6196,N_5596,N_5167);
nor U6197 (N_6197,N_5260,N_5562);
and U6198 (N_6198,N_5237,N_5304);
nor U6199 (N_6199,N_5049,N_5079);
nor U6200 (N_6200,N_5516,N_5046);
or U6201 (N_6201,N_5102,N_5189);
nand U6202 (N_6202,N_5232,N_5498);
nor U6203 (N_6203,N_5222,N_5312);
nand U6204 (N_6204,N_5301,N_5349);
nor U6205 (N_6205,N_5620,N_5520);
nand U6206 (N_6206,N_5309,N_5045);
and U6207 (N_6207,N_5055,N_5574);
nor U6208 (N_6208,N_5342,N_5491);
nor U6209 (N_6209,N_5222,N_5105);
nor U6210 (N_6210,N_5382,N_5486);
xor U6211 (N_6211,N_5342,N_5203);
or U6212 (N_6212,N_5518,N_5307);
or U6213 (N_6213,N_5375,N_5408);
or U6214 (N_6214,N_5383,N_5206);
nor U6215 (N_6215,N_5286,N_5244);
nand U6216 (N_6216,N_5515,N_5537);
nor U6217 (N_6217,N_5577,N_5015);
and U6218 (N_6218,N_5002,N_5365);
nand U6219 (N_6219,N_5152,N_5015);
nand U6220 (N_6220,N_5141,N_5256);
or U6221 (N_6221,N_5015,N_5463);
xor U6222 (N_6222,N_5295,N_5494);
or U6223 (N_6223,N_5607,N_5339);
nor U6224 (N_6224,N_5093,N_5294);
and U6225 (N_6225,N_5129,N_5264);
and U6226 (N_6226,N_5568,N_5107);
xnor U6227 (N_6227,N_5391,N_5516);
or U6228 (N_6228,N_5571,N_5544);
nor U6229 (N_6229,N_5275,N_5387);
nor U6230 (N_6230,N_5390,N_5575);
nor U6231 (N_6231,N_5455,N_5204);
nand U6232 (N_6232,N_5586,N_5616);
xor U6233 (N_6233,N_5102,N_5407);
xnor U6234 (N_6234,N_5263,N_5317);
or U6235 (N_6235,N_5022,N_5033);
nor U6236 (N_6236,N_5030,N_5564);
nand U6237 (N_6237,N_5003,N_5271);
xor U6238 (N_6238,N_5601,N_5527);
or U6239 (N_6239,N_5552,N_5501);
and U6240 (N_6240,N_5031,N_5139);
nand U6241 (N_6241,N_5610,N_5115);
or U6242 (N_6242,N_5596,N_5469);
or U6243 (N_6243,N_5406,N_5511);
nand U6244 (N_6244,N_5492,N_5182);
nor U6245 (N_6245,N_5485,N_5082);
or U6246 (N_6246,N_5331,N_5053);
nor U6247 (N_6247,N_5399,N_5518);
and U6248 (N_6248,N_5253,N_5535);
and U6249 (N_6249,N_5474,N_5127);
nor U6250 (N_6250,N_5845,N_5884);
xor U6251 (N_6251,N_5997,N_5824);
nor U6252 (N_6252,N_5757,N_5750);
xnor U6253 (N_6253,N_5742,N_6185);
or U6254 (N_6254,N_6191,N_5796);
xor U6255 (N_6255,N_6135,N_5926);
and U6256 (N_6256,N_5658,N_5665);
and U6257 (N_6257,N_5853,N_6146);
and U6258 (N_6258,N_5675,N_6022);
xor U6259 (N_6259,N_6005,N_5627);
or U6260 (N_6260,N_6036,N_5799);
nor U6261 (N_6261,N_6170,N_5850);
or U6262 (N_6262,N_6031,N_6240);
or U6263 (N_6263,N_5837,N_6079);
and U6264 (N_6264,N_5732,N_5925);
nor U6265 (N_6265,N_5829,N_5918);
nor U6266 (N_6266,N_5678,N_5780);
or U6267 (N_6267,N_6178,N_5857);
or U6268 (N_6268,N_6159,N_5789);
nor U6269 (N_6269,N_5977,N_5708);
or U6270 (N_6270,N_5896,N_5969);
nand U6271 (N_6271,N_5935,N_5721);
or U6272 (N_6272,N_5712,N_6216);
nand U6273 (N_6273,N_5930,N_6011);
xor U6274 (N_6274,N_5866,N_5746);
nand U6275 (N_6275,N_6035,N_5995);
nand U6276 (N_6276,N_5950,N_5921);
nand U6277 (N_6277,N_6129,N_6181);
nor U6278 (N_6278,N_5723,N_5931);
and U6279 (N_6279,N_5835,N_6149);
nand U6280 (N_6280,N_5970,N_6133);
and U6281 (N_6281,N_6233,N_5830);
or U6282 (N_6282,N_5741,N_6002);
nor U6283 (N_6283,N_6073,N_6143);
xor U6284 (N_6284,N_5916,N_6140);
and U6285 (N_6285,N_5764,N_5785);
or U6286 (N_6286,N_5719,N_6174);
xor U6287 (N_6287,N_6094,N_5646);
nand U6288 (N_6288,N_5941,N_5777);
or U6289 (N_6289,N_5791,N_6189);
nor U6290 (N_6290,N_5852,N_6012);
and U6291 (N_6291,N_6088,N_5864);
and U6292 (N_6292,N_5714,N_6072);
nand U6293 (N_6293,N_6059,N_6217);
xnor U6294 (N_6294,N_5945,N_5841);
and U6295 (N_6295,N_6119,N_6198);
nor U6296 (N_6296,N_5840,N_5983);
xor U6297 (N_6297,N_6049,N_5700);
and U6298 (N_6298,N_5980,N_5869);
nand U6299 (N_6299,N_6186,N_5752);
nor U6300 (N_6300,N_5988,N_6150);
nand U6301 (N_6301,N_5891,N_5671);
nor U6302 (N_6302,N_6228,N_6039);
and U6303 (N_6303,N_6065,N_5858);
or U6304 (N_6304,N_5677,N_5949);
nand U6305 (N_6305,N_5888,N_5848);
or U6306 (N_6306,N_5650,N_6025);
or U6307 (N_6307,N_5961,N_5703);
or U6308 (N_6308,N_5697,N_6082);
nand U6309 (N_6309,N_6184,N_6212);
nor U6310 (N_6310,N_5709,N_6144);
nand U6311 (N_6311,N_6008,N_6046);
xor U6312 (N_6312,N_6125,N_5689);
nor U6313 (N_6313,N_6175,N_5965);
nor U6314 (N_6314,N_5707,N_5812);
and U6315 (N_6315,N_5890,N_6029);
and U6316 (N_6316,N_6098,N_6014);
or U6317 (N_6317,N_5863,N_6118);
nor U6318 (N_6318,N_5762,N_6053);
nor U6319 (N_6319,N_6219,N_6225);
and U6320 (N_6320,N_6113,N_5701);
nand U6321 (N_6321,N_5745,N_6167);
nor U6322 (N_6322,N_5956,N_5635);
and U6323 (N_6323,N_6108,N_5993);
and U6324 (N_6324,N_5744,N_6067);
or U6325 (N_6325,N_5784,N_5914);
and U6326 (N_6326,N_5937,N_6075);
xnor U6327 (N_6327,N_6124,N_5797);
xnor U6328 (N_6328,N_6016,N_5656);
and U6329 (N_6329,N_6068,N_6069);
xnor U6330 (N_6330,N_6169,N_5927);
and U6331 (N_6331,N_5713,N_6131);
and U6332 (N_6332,N_6173,N_5978);
or U6333 (N_6333,N_5808,N_6218);
and U6334 (N_6334,N_6057,N_5690);
or U6335 (N_6335,N_6202,N_6033);
nor U6336 (N_6336,N_6078,N_6043);
nor U6337 (N_6337,N_5883,N_6117);
xnor U6338 (N_6338,N_5986,N_6206);
nor U6339 (N_6339,N_6214,N_5952);
nand U6340 (N_6340,N_6161,N_6199);
or U6341 (N_6341,N_6019,N_6086);
or U6342 (N_6342,N_5628,N_5661);
or U6343 (N_6343,N_6197,N_5892);
nand U6344 (N_6344,N_5818,N_5735);
and U6345 (N_6345,N_6234,N_5960);
or U6346 (N_6346,N_5976,N_6226);
xor U6347 (N_6347,N_5662,N_5885);
and U6348 (N_6348,N_6157,N_6164);
or U6349 (N_6349,N_5669,N_5836);
nand U6350 (N_6350,N_5639,N_5747);
and U6351 (N_6351,N_6000,N_6085);
nand U6352 (N_6352,N_5706,N_6021);
nand U6353 (N_6353,N_5946,N_6231);
or U6354 (N_6354,N_5679,N_5875);
nand U6355 (N_6355,N_5953,N_5938);
or U6356 (N_6356,N_5783,N_5668);
nand U6357 (N_6357,N_6142,N_6128);
and U6358 (N_6358,N_6077,N_6151);
and U6359 (N_6359,N_6051,N_5895);
or U6360 (N_6360,N_5838,N_5641);
nor U6361 (N_6361,N_5994,N_5958);
and U6362 (N_6362,N_5974,N_6101);
or U6363 (N_6363,N_5758,N_5693);
or U6364 (N_6364,N_5731,N_6213);
nand U6365 (N_6365,N_5975,N_6245);
nand U6366 (N_6366,N_5867,N_5851);
and U6367 (N_6367,N_6027,N_5922);
or U6368 (N_6368,N_5985,N_5692);
nand U6369 (N_6369,N_6210,N_6223);
nand U6370 (N_6370,N_5734,N_5910);
xor U6371 (N_6371,N_5694,N_5990);
or U6372 (N_6372,N_5902,N_5828);
and U6373 (N_6373,N_6238,N_5704);
xor U6374 (N_6374,N_5695,N_6044);
nand U6375 (N_6375,N_5827,N_5962);
nor U6376 (N_6376,N_5663,N_6114);
and U6377 (N_6377,N_6127,N_6132);
nand U6378 (N_6378,N_5873,N_6048);
and U6379 (N_6379,N_5972,N_6015);
nor U6380 (N_6380,N_6120,N_5640);
and U6381 (N_6381,N_5657,N_6080);
or U6382 (N_6382,N_5637,N_5907);
and U6383 (N_6383,N_5844,N_5859);
nand U6384 (N_6384,N_6121,N_5765);
nand U6385 (N_6385,N_5940,N_5681);
nand U6386 (N_6386,N_5673,N_6205);
or U6387 (N_6387,N_6055,N_5674);
or U6388 (N_6388,N_5802,N_6147);
nor U6389 (N_6389,N_5815,N_5899);
and U6390 (N_6390,N_5973,N_6116);
and U6391 (N_6391,N_6089,N_6062);
or U6392 (N_6392,N_6162,N_5810);
nor U6393 (N_6393,N_5979,N_6220);
nand U6394 (N_6394,N_5737,N_5908);
nand U6395 (N_6395,N_5736,N_5705);
and U6396 (N_6396,N_5776,N_6211);
or U6397 (N_6397,N_5932,N_6221);
or U6398 (N_6398,N_5963,N_5868);
nor U6399 (N_6399,N_5682,N_5655);
and U6400 (N_6400,N_5730,N_5727);
and U6401 (N_6401,N_5786,N_6097);
nor U6402 (N_6402,N_5722,N_5889);
and U6403 (N_6403,N_5687,N_5872);
nand U6404 (N_6404,N_5670,N_5842);
nor U6405 (N_6405,N_5846,N_5751);
or U6406 (N_6406,N_5644,N_5688);
or U6407 (N_6407,N_5774,N_6092);
or U6408 (N_6408,N_6138,N_6010);
or U6409 (N_6409,N_6242,N_5743);
or U6410 (N_6410,N_5654,N_6081);
or U6411 (N_6411,N_5800,N_5642);
nand U6412 (N_6412,N_5971,N_5766);
and U6413 (N_6413,N_6247,N_6060);
and U6414 (N_6414,N_5816,N_5683);
and U6415 (N_6415,N_5768,N_5893);
xnor U6416 (N_6416,N_6096,N_6163);
nor U6417 (N_6417,N_5767,N_6017);
and U6418 (N_6418,N_5987,N_6103);
nor U6419 (N_6419,N_5632,N_6070);
and U6420 (N_6420,N_5939,N_5809);
nor U6421 (N_6421,N_5648,N_5999);
nand U6422 (N_6422,N_5676,N_5934);
nand U6423 (N_6423,N_6248,N_5805);
or U6424 (N_6424,N_5924,N_5877);
nor U6425 (N_6425,N_5948,N_5726);
or U6426 (N_6426,N_5860,N_6195);
and U6427 (N_6427,N_5728,N_5702);
nor U6428 (N_6428,N_5847,N_5798);
nand U6429 (N_6429,N_6235,N_6026);
nor U6430 (N_6430,N_5964,N_5906);
and U6431 (N_6431,N_5634,N_5984);
xor U6432 (N_6432,N_5653,N_6155);
and U6433 (N_6433,N_5754,N_6004);
xor U6434 (N_6434,N_5710,N_5834);
nor U6435 (N_6435,N_5849,N_5666);
nor U6436 (N_6436,N_6194,N_6112);
or U6437 (N_6437,N_5718,N_5660);
nand U6438 (N_6438,N_6045,N_6152);
nand U6439 (N_6439,N_5643,N_5839);
and U6440 (N_6440,N_5820,N_6136);
nor U6441 (N_6441,N_5778,N_5626);
nor U6442 (N_6442,N_6100,N_5903);
nand U6443 (N_6443,N_5819,N_5915);
nor U6444 (N_6444,N_6204,N_5779);
nor U6445 (N_6445,N_6106,N_5720);
or U6446 (N_6446,N_6193,N_6009);
or U6447 (N_6447,N_5874,N_6034);
and U6448 (N_6448,N_6105,N_5898);
and U6449 (N_6449,N_5822,N_5923);
or U6450 (N_6450,N_5951,N_5792);
xor U6451 (N_6451,N_5667,N_5759);
or U6452 (N_6452,N_5711,N_6196);
nor U6453 (N_6453,N_6249,N_5724);
nor U6454 (N_6454,N_6076,N_6038);
nand U6455 (N_6455,N_6050,N_5912);
nand U6456 (N_6456,N_5801,N_5699);
and U6457 (N_6457,N_6001,N_6166);
xnor U6458 (N_6458,N_5862,N_6047);
and U6459 (N_6459,N_6182,N_5806);
nand U6460 (N_6460,N_5659,N_6153);
and U6461 (N_6461,N_5861,N_5775);
or U6462 (N_6462,N_6123,N_5817);
or U6463 (N_6463,N_5942,N_6111);
xor U6464 (N_6464,N_6040,N_5803);
nand U6465 (N_6465,N_5790,N_5716);
and U6466 (N_6466,N_6052,N_6222);
nand U6467 (N_6467,N_6165,N_6229);
nand U6468 (N_6468,N_5739,N_5981);
and U6469 (N_6469,N_6041,N_5833);
nor U6470 (N_6470,N_5717,N_5696);
and U6471 (N_6471,N_5771,N_5855);
nor U6472 (N_6472,N_6054,N_5904);
or U6473 (N_6473,N_6084,N_5871);
xnor U6474 (N_6474,N_5686,N_6071);
and U6475 (N_6475,N_5633,N_5821);
or U6476 (N_6476,N_5740,N_6102);
or U6477 (N_6477,N_5715,N_5879);
nand U6478 (N_6478,N_5947,N_5920);
xor U6479 (N_6479,N_5913,N_5664);
or U6480 (N_6480,N_5804,N_6095);
or U6481 (N_6481,N_5911,N_6074);
nor U6482 (N_6482,N_6203,N_5991);
and U6483 (N_6483,N_5966,N_6187);
or U6484 (N_6484,N_5773,N_6130);
and U6485 (N_6485,N_6176,N_6091);
and U6486 (N_6486,N_6104,N_5919);
and U6487 (N_6487,N_5807,N_5955);
nor U6488 (N_6488,N_6020,N_6188);
nand U6489 (N_6489,N_6007,N_5989);
nor U6490 (N_6490,N_5967,N_6244);
nor U6491 (N_6491,N_5831,N_5929);
nand U6492 (N_6492,N_6030,N_6018);
nand U6493 (N_6493,N_6093,N_5944);
nor U6494 (N_6494,N_6042,N_5886);
or U6495 (N_6495,N_5813,N_6243);
or U6496 (N_6496,N_5826,N_5685);
or U6497 (N_6497,N_6083,N_5900);
nor U6498 (N_6498,N_6006,N_5887);
and U6499 (N_6499,N_5636,N_5625);
or U6500 (N_6500,N_6110,N_5856);
nor U6501 (N_6501,N_5865,N_5825);
nor U6502 (N_6502,N_6232,N_6099);
nor U6503 (N_6503,N_6239,N_6148);
nor U6504 (N_6504,N_6087,N_6037);
or U6505 (N_6505,N_5917,N_5897);
nand U6506 (N_6506,N_5996,N_6179);
nor U6507 (N_6507,N_6115,N_6241);
and U6508 (N_6508,N_6246,N_5788);
and U6509 (N_6509,N_5770,N_5901);
nand U6510 (N_6510,N_6158,N_6180);
and U6511 (N_6511,N_6227,N_5652);
nor U6512 (N_6512,N_5733,N_6207);
nand U6513 (N_6513,N_5936,N_5992);
xnor U6514 (N_6514,N_5795,N_6208);
nor U6515 (N_6515,N_6160,N_5843);
or U6516 (N_6516,N_5781,N_6237);
nor U6517 (N_6517,N_5954,N_5691);
nand U6518 (N_6518,N_5631,N_6200);
nor U6519 (N_6519,N_6028,N_6177);
nor U6520 (N_6520,N_6230,N_5761);
or U6521 (N_6521,N_5645,N_6192);
nand U6522 (N_6522,N_6064,N_6201);
xor U6523 (N_6523,N_6063,N_6061);
and U6524 (N_6524,N_5968,N_5959);
nor U6525 (N_6525,N_6215,N_6209);
and U6526 (N_6526,N_5630,N_5748);
or U6527 (N_6527,N_6134,N_5772);
or U6528 (N_6528,N_6236,N_5725);
nor U6529 (N_6529,N_6090,N_6003);
nand U6530 (N_6530,N_6139,N_5753);
nand U6531 (N_6531,N_6172,N_5909);
nor U6532 (N_6532,N_6122,N_6024);
nand U6533 (N_6533,N_5629,N_5763);
nand U6534 (N_6534,N_5647,N_5782);
and U6535 (N_6535,N_5760,N_5998);
or U6536 (N_6536,N_6126,N_5882);
nor U6537 (N_6537,N_5769,N_6066);
nor U6538 (N_6538,N_6013,N_6190);
and U6539 (N_6539,N_5638,N_5928);
and U6540 (N_6540,N_5738,N_5811);
and U6541 (N_6541,N_6058,N_5729);
or U6542 (N_6542,N_6154,N_5823);
or U6543 (N_6543,N_5651,N_6141);
or U6544 (N_6544,N_5957,N_6183);
or U6545 (N_6545,N_5832,N_6023);
or U6546 (N_6546,N_6107,N_5943);
or U6547 (N_6547,N_5905,N_6156);
nand U6548 (N_6548,N_5894,N_5880);
or U6549 (N_6549,N_6168,N_6145);
and U6550 (N_6550,N_5876,N_5649);
and U6551 (N_6551,N_5672,N_5756);
and U6552 (N_6552,N_5680,N_5793);
or U6553 (N_6553,N_5749,N_5878);
nand U6554 (N_6554,N_5933,N_5870);
xor U6555 (N_6555,N_5684,N_5755);
and U6556 (N_6556,N_6032,N_6171);
nand U6557 (N_6557,N_6137,N_5794);
and U6558 (N_6558,N_6056,N_5814);
xnor U6559 (N_6559,N_5881,N_5854);
nor U6560 (N_6560,N_5787,N_6224);
nand U6561 (N_6561,N_5698,N_6109);
or U6562 (N_6562,N_5982,N_6107);
or U6563 (N_6563,N_6189,N_6134);
xor U6564 (N_6564,N_5945,N_5653);
nand U6565 (N_6565,N_5727,N_6006);
nand U6566 (N_6566,N_6234,N_5792);
and U6567 (N_6567,N_5648,N_6207);
nor U6568 (N_6568,N_5708,N_5874);
or U6569 (N_6569,N_6206,N_6135);
nand U6570 (N_6570,N_5641,N_5896);
or U6571 (N_6571,N_6050,N_5868);
and U6572 (N_6572,N_5866,N_6061);
nand U6573 (N_6573,N_5844,N_6221);
nand U6574 (N_6574,N_5847,N_6178);
xnor U6575 (N_6575,N_6111,N_5995);
nand U6576 (N_6576,N_5939,N_6238);
or U6577 (N_6577,N_5680,N_5884);
nor U6578 (N_6578,N_6150,N_5803);
or U6579 (N_6579,N_6159,N_6137);
nand U6580 (N_6580,N_5689,N_6234);
xor U6581 (N_6581,N_6179,N_5907);
nand U6582 (N_6582,N_5828,N_5994);
nand U6583 (N_6583,N_6159,N_5714);
or U6584 (N_6584,N_5633,N_5844);
or U6585 (N_6585,N_5657,N_6162);
nor U6586 (N_6586,N_6107,N_5665);
nor U6587 (N_6587,N_5758,N_5786);
or U6588 (N_6588,N_5952,N_5839);
and U6589 (N_6589,N_5950,N_5789);
nor U6590 (N_6590,N_5974,N_5780);
nor U6591 (N_6591,N_5756,N_5791);
nor U6592 (N_6592,N_6110,N_5899);
and U6593 (N_6593,N_5663,N_5755);
nand U6594 (N_6594,N_5951,N_6237);
nand U6595 (N_6595,N_5760,N_6228);
and U6596 (N_6596,N_5834,N_6110);
nand U6597 (N_6597,N_5865,N_6220);
or U6598 (N_6598,N_6151,N_5816);
nor U6599 (N_6599,N_5870,N_6079);
nor U6600 (N_6600,N_5866,N_6232);
or U6601 (N_6601,N_6013,N_6120);
and U6602 (N_6602,N_5726,N_5711);
xnor U6603 (N_6603,N_5720,N_6025);
and U6604 (N_6604,N_6109,N_5968);
xnor U6605 (N_6605,N_5744,N_5636);
nor U6606 (N_6606,N_5844,N_6124);
nor U6607 (N_6607,N_6046,N_5657);
xnor U6608 (N_6608,N_5706,N_5771);
nor U6609 (N_6609,N_6101,N_5887);
nor U6610 (N_6610,N_6127,N_5751);
nand U6611 (N_6611,N_6018,N_5990);
nand U6612 (N_6612,N_5687,N_5844);
and U6613 (N_6613,N_5826,N_6142);
nand U6614 (N_6614,N_6008,N_5739);
and U6615 (N_6615,N_5839,N_6117);
or U6616 (N_6616,N_5922,N_5827);
nor U6617 (N_6617,N_6111,N_5815);
nor U6618 (N_6618,N_6045,N_6151);
and U6619 (N_6619,N_6175,N_6128);
nor U6620 (N_6620,N_6099,N_5790);
nand U6621 (N_6621,N_5932,N_5837);
or U6622 (N_6622,N_5739,N_5867);
xnor U6623 (N_6623,N_6070,N_5643);
nor U6624 (N_6624,N_5706,N_6123);
nand U6625 (N_6625,N_5841,N_5974);
or U6626 (N_6626,N_6114,N_6093);
and U6627 (N_6627,N_5984,N_5724);
nand U6628 (N_6628,N_5735,N_6047);
nor U6629 (N_6629,N_5711,N_6043);
xor U6630 (N_6630,N_5960,N_5768);
xor U6631 (N_6631,N_5949,N_5780);
or U6632 (N_6632,N_5837,N_5924);
or U6633 (N_6633,N_5741,N_6020);
or U6634 (N_6634,N_6121,N_5867);
or U6635 (N_6635,N_5842,N_5920);
nor U6636 (N_6636,N_6153,N_5865);
nor U6637 (N_6637,N_6206,N_6195);
or U6638 (N_6638,N_6186,N_5668);
or U6639 (N_6639,N_5769,N_6208);
and U6640 (N_6640,N_5939,N_5681);
or U6641 (N_6641,N_5666,N_5979);
or U6642 (N_6642,N_5770,N_5952);
and U6643 (N_6643,N_6249,N_5801);
nand U6644 (N_6644,N_6070,N_5704);
or U6645 (N_6645,N_5961,N_5818);
nand U6646 (N_6646,N_6096,N_5961);
nand U6647 (N_6647,N_5713,N_5726);
nand U6648 (N_6648,N_5805,N_6096);
xor U6649 (N_6649,N_6178,N_5976);
and U6650 (N_6650,N_5887,N_6088);
and U6651 (N_6651,N_5636,N_5779);
nand U6652 (N_6652,N_5664,N_5976);
nor U6653 (N_6653,N_6098,N_5985);
or U6654 (N_6654,N_5754,N_5772);
nor U6655 (N_6655,N_6060,N_5929);
and U6656 (N_6656,N_6042,N_6201);
nor U6657 (N_6657,N_5777,N_5836);
nor U6658 (N_6658,N_5877,N_6060);
xor U6659 (N_6659,N_5956,N_5801);
xor U6660 (N_6660,N_5854,N_5707);
nor U6661 (N_6661,N_5719,N_6203);
or U6662 (N_6662,N_6030,N_6186);
nand U6663 (N_6663,N_5965,N_6108);
xnor U6664 (N_6664,N_6160,N_5769);
or U6665 (N_6665,N_5876,N_5678);
nand U6666 (N_6666,N_6223,N_5847);
nor U6667 (N_6667,N_5730,N_6076);
nand U6668 (N_6668,N_6175,N_5816);
or U6669 (N_6669,N_5706,N_6127);
nand U6670 (N_6670,N_5736,N_5772);
and U6671 (N_6671,N_5918,N_5898);
or U6672 (N_6672,N_6208,N_5944);
or U6673 (N_6673,N_5767,N_5981);
nand U6674 (N_6674,N_5950,N_6185);
and U6675 (N_6675,N_5625,N_5864);
nand U6676 (N_6676,N_6176,N_5759);
or U6677 (N_6677,N_6132,N_6112);
nand U6678 (N_6678,N_6199,N_5886);
or U6679 (N_6679,N_6040,N_5899);
nor U6680 (N_6680,N_5727,N_5869);
and U6681 (N_6681,N_5792,N_5886);
nor U6682 (N_6682,N_5884,N_5853);
or U6683 (N_6683,N_6152,N_6133);
xnor U6684 (N_6684,N_6028,N_6063);
or U6685 (N_6685,N_5910,N_5842);
nor U6686 (N_6686,N_5643,N_5802);
xor U6687 (N_6687,N_6029,N_6131);
or U6688 (N_6688,N_6220,N_5976);
and U6689 (N_6689,N_6224,N_6190);
nand U6690 (N_6690,N_5824,N_5789);
or U6691 (N_6691,N_5790,N_5714);
nor U6692 (N_6692,N_6050,N_6214);
xnor U6693 (N_6693,N_5814,N_5802);
and U6694 (N_6694,N_5954,N_6118);
or U6695 (N_6695,N_6208,N_6084);
or U6696 (N_6696,N_6094,N_5696);
xor U6697 (N_6697,N_6111,N_5909);
nand U6698 (N_6698,N_5669,N_5942);
and U6699 (N_6699,N_5904,N_5684);
nand U6700 (N_6700,N_6221,N_5861);
or U6701 (N_6701,N_5789,N_5715);
or U6702 (N_6702,N_6040,N_6203);
and U6703 (N_6703,N_6017,N_6115);
nor U6704 (N_6704,N_6229,N_5842);
and U6705 (N_6705,N_5813,N_6201);
nand U6706 (N_6706,N_6003,N_6249);
and U6707 (N_6707,N_5998,N_6022);
and U6708 (N_6708,N_5956,N_6236);
nor U6709 (N_6709,N_5897,N_5879);
or U6710 (N_6710,N_6226,N_5642);
or U6711 (N_6711,N_5890,N_6130);
xor U6712 (N_6712,N_5940,N_5696);
or U6713 (N_6713,N_6121,N_5910);
nand U6714 (N_6714,N_5661,N_5849);
nor U6715 (N_6715,N_5781,N_6244);
or U6716 (N_6716,N_6114,N_6136);
and U6717 (N_6717,N_5950,N_5669);
and U6718 (N_6718,N_5902,N_6045);
nor U6719 (N_6719,N_5957,N_5748);
nand U6720 (N_6720,N_6175,N_5944);
and U6721 (N_6721,N_5626,N_5720);
or U6722 (N_6722,N_5732,N_6056);
nor U6723 (N_6723,N_5725,N_5716);
nor U6724 (N_6724,N_6204,N_5751);
xnor U6725 (N_6725,N_5862,N_6202);
nor U6726 (N_6726,N_5767,N_5846);
nor U6727 (N_6727,N_5850,N_5877);
xor U6728 (N_6728,N_6145,N_5928);
nor U6729 (N_6729,N_5772,N_6234);
nor U6730 (N_6730,N_6242,N_6186);
and U6731 (N_6731,N_6235,N_5904);
nor U6732 (N_6732,N_5689,N_6128);
nand U6733 (N_6733,N_5889,N_5711);
nand U6734 (N_6734,N_5711,N_5649);
and U6735 (N_6735,N_6036,N_6155);
nor U6736 (N_6736,N_6174,N_6128);
nor U6737 (N_6737,N_6221,N_6153);
or U6738 (N_6738,N_5915,N_6063);
or U6739 (N_6739,N_5802,N_5669);
and U6740 (N_6740,N_5946,N_5980);
nor U6741 (N_6741,N_5836,N_6089);
and U6742 (N_6742,N_5753,N_5942);
and U6743 (N_6743,N_6002,N_6011);
and U6744 (N_6744,N_6086,N_5812);
nor U6745 (N_6745,N_6176,N_5772);
nor U6746 (N_6746,N_6192,N_5812);
or U6747 (N_6747,N_6216,N_6155);
nor U6748 (N_6748,N_6165,N_5911);
nand U6749 (N_6749,N_6114,N_5816);
or U6750 (N_6750,N_5652,N_5783);
or U6751 (N_6751,N_5689,N_5857);
nor U6752 (N_6752,N_5700,N_5990);
nor U6753 (N_6753,N_5859,N_6150);
and U6754 (N_6754,N_5924,N_6000);
or U6755 (N_6755,N_5942,N_6225);
nand U6756 (N_6756,N_5959,N_5745);
xnor U6757 (N_6757,N_6085,N_5759);
nor U6758 (N_6758,N_6092,N_5664);
nand U6759 (N_6759,N_5896,N_5648);
or U6760 (N_6760,N_6155,N_5686);
or U6761 (N_6761,N_6114,N_6222);
nor U6762 (N_6762,N_6060,N_5685);
nor U6763 (N_6763,N_5878,N_5646);
and U6764 (N_6764,N_5665,N_6096);
nor U6765 (N_6765,N_6063,N_5685);
nor U6766 (N_6766,N_5750,N_5802);
nor U6767 (N_6767,N_5779,N_6054);
and U6768 (N_6768,N_6122,N_6198);
nand U6769 (N_6769,N_5701,N_5697);
and U6770 (N_6770,N_6004,N_5940);
nor U6771 (N_6771,N_5779,N_5753);
xnor U6772 (N_6772,N_5829,N_5934);
nand U6773 (N_6773,N_5897,N_5780);
nand U6774 (N_6774,N_5994,N_5795);
nor U6775 (N_6775,N_6149,N_6184);
or U6776 (N_6776,N_6093,N_6028);
or U6777 (N_6777,N_5664,N_5906);
or U6778 (N_6778,N_5732,N_5881);
nand U6779 (N_6779,N_6057,N_6182);
or U6780 (N_6780,N_6134,N_5925);
xnor U6781 (N_6781,N_6127,N_5889);
or U6782 (N_6782,N_5847,N_6237);
and U6783 (N_6783,N_5894,N_6239);
nor U6784 (N_6784,N_5989,N_5866);
nor U6785 (N_6785,N_6009,N_6131);
and U6786 (N_6786,N_6131,N_5868);
xor U6787 (N_6787,N_5848,N_5630);
or U6788 (N_6788,N_5796,N_6123);
and U6789 (N_6789,N_5750,N_5844);
and U6790 (N_6790,N_5743,N_5806);
and U6791 (N_6791,N_5655,N_5959);
nor U6792 (N_6792,N_5670,N_5941);
nor U6793 (N_6793,N_6137,N_5717);
nor U6794 (N_6794,N_6136,N_6039);
nand U6795 (N_6795,N_6164,N_5659);
nand U6796 (N_6796,N_6040,N_6078);
nor U6797 (N_6797,N_6050,N_6239);
or U6798 (N_6798,N_6070,N_5980);
or U6799 (N_6799,N_6202,N_6232);
nor U6800 (N_6800,N_5832,N_5965);
or U6801 (N_6801,N_6200,N_5891);
or U6802 (N_6802,N_6125,N_6159);
or U6803 (N_6803,N_5990,N_5991);
nor U6804 (N_6804,N_5673,N_5843);
nor U6805 (N_6805,N_5739,N_5905);
nor U6806 (N_6806,N_5793,N_5914);
nand U6807 (N_6807,N_5852,N_5728);
nand U6808 (N_6808,N_5906,N_6066);
or U6809 (N_6809,N_5722,N_5772);
xor U6810 (N_6810,N_6126,N_5992);
nand U6811 (N_6811,N_5865,N_6065);
or U6812 (N_6812,N_6096,N_5774);
and U6813 (N_6813,N_5770,N_5851);
nand U6814 (N_6814,N_6090,N_6204);
nor U6815 (N_6815,N_5924,N_5797);
or U6816 (N_6816,N_6105,N_6206);
and U6817 (N_6817,N_5776,N_5887);
and U6818 (N_6818,N_5937,N_5865);
xor U6819 (N_6819,N_5800,N_6104);
and U6820 (N_6820,N_5977,N_5659);
nor U6821 (N_6821,N_6207,N_5776);
nor U6822 (N_6822,N_5853,N_6074);
nand U6823 (N_6823,N_5720,N_5850);
nor U6824 (N_6824,N_5931,N_5967);
and U6825 (N_6825,N_5633,N_6106);
and U6826 (N_6826,N_5817,N_6149);
or U6827 (N_6827,N_5830,N_5847);
nor U6828 (N_6828,N_5742,N_5736);
nor U6829 (N_6829,N_5775,N_6047);
or U6830 (N_6830,N_6102,N_6208);
or U6831 (N_6831,N_5810,N_6039);
or U6832 (N_6832,N_5909,N_5741);
nand U6833 (N_6833,N_5890,N_5884);
nor U6834 (N_6834,N_5867,N_5722);
nand U6835 (N_6835,N_6138,N_5899);
nand U6836 (N_6836,N_5828,N_5893);
or U6837 (N_6837,N_6074,N_5795);
nor U6838 (N_6838,N_6028,N_5731);
nor U6839 (N_6839,N_6047,N_6058);
and U6840 (N_6840,N_6087,N_6101);
or U6841 (N_6841,N_5880,N_5860);
or U6842 (N_6842,N_5968,N_5729);
xnor U6843 (N_6843,N_6031,N_5680);
nand U6844 (N_6844,N_5804,N_5673);
and U6845 (N_6845,N_6231,N_5767);
nand U6846 (N_6846,N_6188,N_5699);
nor U6847 (N_6847,N_6195,N_5647);
nor U6848 (N_6848,N_6195,N_5854);
xor U6849 (N_6849,N_5629,N_6216);
and U6850 (N_6850,N_5877,N_5799);
nor U6851 (N_6851,N_5786,N_5959);
nand U6852 (N_6852,N_5726,N_6195);
or U6853 (N_6853,N_5628,N_5691);
and U6854 (N_6854,N_6137,N_5887);
or U6855 (N_6855,N_6000,N_6196);
and U6856 (N_6856,N_6114,N_5749);
nor U6857 (N_6857,N_5883,N_6018);
nor U6858 (N_6858,N_6205,N_5887);
nand U6859 (N_6859,N_6198,N_6153);
and U6860 (N_6860,N_6085,N_6073);
or U6861 (N_6861,N_5940,N_5634);
nand U6862 (N_6862,N_5774,N_5746);
nand U6863 (N_6863,N_5699,N_5903);
xnor U6864 (N_6864,N_6117,N_5700);
xor U6865 (N_6865,N_5952,N_6052);
nand U6866 (N_6866,N_5819,N_6102);
nand U6867 (N_6867,N_5636,N_6097);
nor U6868 (N_6868,N_6143,N_6020);
and U6869 (N_6869,N_5853,N_6238);
or U6870 (N_6870,N_5653,N_6088);
nor U6871 (N_6871,N_5894,N_5744);
or U6872 (N_6872,N_5734,N_5791);
or U6873 (N_6873,N_6209,N_5786);
nor U6874 (N_6874,N_5981,N_5682);
or U6875 (N_6875,N_6734,N_6404);
or U6876 (N_6876,N_6272,N_6266);
nor U6877 (N_6877,N_6854,N_6618);
nand U6878 (N_6878,N_6324,N_6758);
or U6879 (N_6879,N_6619,N_6779);
nand U6880 (N_6880,N_6699,N_6262);
or U6881 (N_6881,N_6634,N_6674);
or U6882 (N_6882,N_6673,N_6525);
nand U6883 (N_6883,N_6306,N_6478);
nand U6884 (N_6884,N_6292,N_6279);
xnor U6885 (N_6885,N_6599,N_6724);
nand U6886 (N_6886,N_6851,N_6498);
nand U6887 (N_6887,N_6268,N_6356);
or U6888 (N_6888,N_6664,N_6718);
or U6889 (N_6889,N_6330,N_6757);
nor U6890 (N_6890,N_6644,N_6872);
nor U6891 (N_6891,N_6541,N_6586);
and U6892 (N_6892,N_6428,N_6472);
and U6893 (N_6893,N_6802,N_6832);
and U6894 (N_6894,N_6701,N_6742);
and U6895 (N_6895,N_6322,N_6829);
nand U6896 (N_6896,N_6861,N_6588);
nor U6897 (N_6897,N_6308,N_6693);
nand U6898 (N_6898,N_6390,N_6377);
nor U6899 (N_6899,N_6783,N_6833);
or U6900 (N_6900,N_6333,N_6679);
nand U6901 (N_6901,N_6696,N_6513);
and U6902 (N_6902,N_6766,N_6837);
nand U6903 (N_6903,N_6413,N_6780);
nor U6904 (N_6904,N_6274,N_6494);
nand U6905 (N_6905,N_6735,N_6489);
nand U6906 (N_6906,N_6560,N_6805);
nor U6907 (N_6907,N_6749,N_6566);
nor U6908 (N_6908,N_6380,N_6775);
nand U6909 (N_6909,N_6490,N_6553);
or U6910 (N_6910,N_6457,N_6339);
or U6911 (N_6911,N_6676,N_6311);
nand U6912 (N_6912,N_6425,N_6799);
nand U6913 (N_6913,N_6406,N_6350);
or U6914 (N_6914,N_6435,N_6710);
and U6915 (N_6915,N_6862,N_6420);
nor U6916 (N_6916,N_6508,N_6589);
and U6917 (N_6917,N_6819,N_6656);
nand U6918 (N_6918,N_6343,N_6442);
and U6919 (N_6919,N_6767,N_6329);
nor U6920 (N_6920,N_6482,N_6795);
nand U6921 (N_6921,N_6637,N_6546);
or U6922 (N_6922,N_6352,N_6858);
nor U6923 (N_6923,N_6410,N_6869);
nor U6924 (N_6924,N_6743,N_6764);
nand U6925 (N_6925,N_6373,N_6446);
or U6926 (N_6926,N_6526,N_6838);
xor U6927 (N_6927,N_6815,N_6276);
nand U6928 (N_6928,N_6521,N_6709);
nand U6929 (N_6929,N_6405,N_6667);
nand U6930 (N_6930,N_6627,N_6579);
xor U6931 (N_6931,N_6790,N_6340);
or U6932 (N_6932,N_6839,N_6641);
nand U6933 (N_6933,N_6323,N_6778);
or U6934 (N_6934,N_6290,N_6635);
nand U6935 (N_6935,N_6830,N_6721);
xnor U6936 (N_6936,N_6313,N_6584);
and U6937 (N_6937,N_6573,N_6580);
and U6938 (N_6938,N_6448,N_6865);
and U6939 (N_6939,N_6273,N_6629);
nor U6940 (N_6940,N_6355,N_6471);
nand U6941 (N_6941,N_6737,N_6504);
or U6942 (N_6942,N_6361,N_6314);
or U6943 (N_6943,N_6828,N_6259);
nor U6944 (N_6944,N_6711,N_6852);
nand U6945 (N_6945,N_6611,N_6787);
and U6946 (N_6946,N_6319,N_6336);
or U6947 (N_6947,N_6260,N_6871);
nor U6948 (N_6948,N_6285,N_6646);
nor U6949 (N_6949,N_6762,N_6844);
and U6950 (N_6950,N_6581,N_6782);
nand U6951 (N_6951,N_6368,N_6370);
or U6952 (N_6952,N_6297,N_6789);
or U6953 (N_6953,N_6557,N_6280);
nor U6954 (N_6954,N_6597,N_6376);
or U6955 (N_6955,N_6744,N_6493);
nand U6956 (N_6956,N_6296,N_6874);
nand U6957 (N_6957,N_6661,N_6564);
and U6958 (N_6958,N_6432,N_6495);
nor U6959 (N_6959,N_6607,N_6717);
nor U6960 (N_6960,N_6807,N_6347);
and U6961 (N_6961,N_6626,N_6283);
nand U6962 (N_6962,N_6451,N_6590);
xor U6963 (N_6963,N_6592,N_6258);
and U6964 (N_6964,N_6388,N_6543);
or U6965 (N_6965,N_6542,N_6403);
and U6966 (N_6966,N_6687,N_6264);
or U6967 (N_6967,N_6344,N_6555);
and U6968 (N_6968,N_6514,N_6371);
and U6969 (N_6969,N_6554,N_6394);
and U6970 (N_6970,N_6824,N_6253);
nand U6971 (N_6971,N_6715,N_6840);
and U6972 (N_6972,N_6797,N_6353);
nor U6973 (N_6973,N_6278,N_6583);
nand U6974 (N_6974,N_6796,N_6469);
or U6975 (N_6975,N_6746,N_6295);
nor U6976 (N_6976,N_6366,N_6843);
xnor U6977 (N_6977,N_6315,N_6801);
nand U6978 (N_6978,N_6518,N_6770);
nand U6979 (N_6979,N_6302,N_6614);
nor U6980 (N_6980,N_6341,N_6299);
or U6981 (N_6981,N_6659,N_6603);
nor U6982 (N_6982,N_6456,N_6683);
or U6983 (N_6983,N_6825,N_6503);
and U6984 (N_6984,N_6288,N_6692);
and U6985 (N_6985,N_6548,N_6332);
and U6986 (N_6986,N_6400,N_6427);
nand U6987 (N_6987,N_6385,N_6447);
and U6988 (N_6988,N_6678,N_6537);
nor U6989 (N_6989,N_6433,N_6873);
and U6990 (N_6990,N_6487,N_6765);
nand U6991 (N_6991,N_6424,N_6691);
nor U6992 (N_6992,N_6863,N_6856);
nor U6993 (N_6993,N_6816,N_6587);
or U6994 (N_6994,N_6294,N_6270);
and U6995 (N_6995,N_6458,N_6731);
nor U6996 (N_6996,N_6608,N_6642);
nor U6997 (N_6997,N_6545,N_6534);
and U6998 (N_6998,N_6741,N_6640);
xnor U6999 (N_6999,N_6577,N_6499);
nor U7000 (N_7000,N_6853,N_6567);
nor U7001 (N_7001,N_6519,N_6609);
nand U7002 (N_7002,N_6475,N_6658);
nor U7003 (N_7003,N_6360,N_6254);
nand U7004 (N_7004,N_6625,N_6289);
or U7005 (N_7005,N_6857,N_6615);
and U7006 (N_7006,N_6655,N_6491);
and U7007 (N_7007,N_6275,N_6335);
and U7008 (N_7008,N_6723,N_6812);
nor U7009 (N_7009,N_6751,N_6349);
nand U7010 (N_7010,N_6798,N_6663);
and U7011 (N_7011,N_6831,N_6455);
xnor U7012 (N_7012,N_6649,N_6814);
xor U7013 (N_7013,N_6675,N_6565);
and U7014 (N_7014,N_6530,N_6774);
nand U7015 (N_7015,N_6510,N_6505);
nor U7016 (N_7016,N_6415,N_6466);
or U7017 (N_7017,N_6484,N_6287);
or U7018 (N_7018,N_6794,N_6739);
nor U7019 (N_7019,N_6422,N_6511);
and U7020 (N_7020,N_6585,N_6321);
or U7021 (N_7021,N_6301,N_6777);
or U7022 (N_7022,N_6345,N_6492);
nand U7023 (N_7023,N_6485,N_6791);
xnor U7024 (N_7024,N_6680,N_6453);
and U7025 (N_7025,N_6378,N_6317);
nand U7026 (N_7026,N_6617,N_6716);
or U7027 (N_7027,N_6776,N_6357);
or U7028 (N_7028,N_6506,N_6808);
nor U7029 (N_7029,N_6535,N_6702);
nor U7030 (N_7030,N_6686,N_6396);
nor U7031 (N_7031,N_6439,N_6849);
xor U7032 (N_7032,N_6576,N_6327);
and U7033 (N_7033,N_6533,N_6509);
or U7034 (N_7034,N_6601,N_6395);
nor U7035 (N_7035,N_6517,N_6501);
nor U7036 (N_7036,N_6414,N_6417);
xnor U7037 (N_7037,N_6527,N_6441);
nand U7038 (N_7038,N_6729,N_6271);
nor U7039 (N_7039,N_6745,N_6684);
and U7040 (N_7040,N_6841,N_6563);
and U7041 (N_7041,N_6346,N_6267);
and U7042 (N_7042,N_6689,N_6773);
xnor U7043 (N_7043,N_6714,N_6497);
nor U7044 (N_7044,N_6756,N_6393);
nand U7045 (N_7045,N_6444,N_6769);
or U7046 (N_7046,N_6593,N_6720);
nor U7047 (N_7047,N_6544,N_6364);
nand U7048 (N_7048,N_6250,N_6648);
or U7049 (N_7049,N_6834,N_6612);
and U7050 (N_7050,N_6747,N_6540);
nand U7051 (N_7051,N_6402,N_6470);
nor U7052 (N_7052,N_6284,N_6558);
or U7053 (N_7053,N_6468,N_6507);
or U7054 (N_7054,N_6461,N_6662);
or U7055 (N_7055,N_6325,N_6685);
or U7056 (N_7056,N_6652,N_6620);
xor U7057 (N_7057,N_6320,N_6529);
or U7058 (N_7058,N_6318,N_6551);
nand U7059 (N_7059,N_6342,N_6465);
xor U7060 (N_7060,N_6632,N_6528);
or U7061 (N_7061,N_6855,N_6477);
nand U7062 (N_7062,N_6450,N_6610);
nor U7063 (N_7063,N_6677,N_6556);
nand U7064 (N_7064,N_6639,N_6363);
nor U7065 (N_7065,N_6867,N_6719);
or U7066 (N_7066,N_6647,N_6571);
nor U7067 (N_7067,N_6730,N_6500);
or U7068 (N_7068,N_6359,N_6752);
or U7069 (N_7069,N_6516,N_6572);
and U7070 (N_7070,N_6600,N_6362);
nand U7071 (N_7071,N_6547,N_6522);
nor U7072 (N_7072,N_6460,N_6672);
and U7073 (N_7073,N_6622,N_6616);
nor U7074 (N_7074,N_6643,N_6552);
nand U7075 (N_7075,N_6864,N_6256);
xnor U7076 (N_7076,N_6300,N_6426);
or U7077 (N_7077,N_6826,N_6419);
and U7078 (N_7078,N_6559,N_6381);
nor U7079 (N_7079,N_6624,N_6454);
nand U7080 (N_7080,N_6578,N_6358);
nand U7081 (N_7081,N_6502,N_6860);
or U7082 (N_7082,N_6866,N_6606);
nor U7083 (N_7083,N_6348,N_6265);
nand U7084 (N_7084,N_6631,N_6850);
nand U7085 (N_7085,N_6462,N_6712);
nor U7086 (N_7086,N_6705,N_6416);
or U7087 (N_7087,N_6707,N_6836);
nor U7088 (N_7088,N_6792,N_6401);
and U7089 (N_7089,N_6269,N_6549);
and U7090 (N_7090,N_6411,N_6387);
or U7091 (N_7091,N_6440,N_6310);
and U7092 (N_7092,N_6682,N_6391);
or U7093 (N_7093,N_6623,N_6842);
nand U7094 (N_7094,N_6392,N_6602);
or U7095 (N_7095,N_6331,N_6397);
nand U7096 (N_7096,N_6326,N_6868);
nor U7097 (N_7097,N_6480,N_6645);
xor U7098 (N_7098,N_6354,N_6698);
or U7099 (N_7099,N_6800,N_6409);
or U7100 (N_7100,N_6464,N_6657);
or U7101 (N_7101,N_6727,N_6605);
xor U7102 (N_7102,N_6628,N_6694);
xnor U7103 (N_7103,N_6732,N_6845);
nand U7104 (N_7104,N_6538,N_6793);
nand U7105 (N_7105,N_6316,N_6474);
or U7106 (N_7106,N_6430,N_6688);
nor U7107 (N_7107,N_6379,N_6809);
nand U7108 (N_7108,N_6367,N_6820);
or U7109 (N_7109,N_6591,N_6436);
and U7110 (N_7110,N_6725,N_6713);
xnor U7111 (N_7111,N_6613,N_6810);
nor U7112 (N_7112,N_6681,N_6277);
or U7113 (N_7113,N_6784,N_6452);
xnor U7114 (N_7114,N_6736,N_6337);
or U7115 (N_7115,N_6304,N_6594);
or U7116 (N_7116,N_6759,N_6660);
and U7117 (N_7117,N_6496,N_6650);
nand U7118 (N_7118,N_6722,N_6728);
nor U7119 (N_7119,N_6286,N_6598);
nor U7120 (N_7120,N_6374,N_6700);
nor U7121 (N_7121,N_6291,N_6515);
nand U7122 (N_7122,N_6703,N_6847);
and U7123 (N_7123,N_6365,N_6298);
and U7124 (N_7124,N_6811,N_6595);
nor U7125 (N_7125,N_6668,N_6255);
nor U7126 (N_7126,N_6386,N_6785);
or U7127 (N_7127,N_6582,N_6786);
nand U7128 (N_7128,N_6369,N_6383);
or U7129 (N_7129,N_6670,N_6338);
and U7130 (N_7130,N_6818,N_6813);
nand U7131 (N_7131,N_6669,N_6621);
nor U7132 (N_7132,N_6536,N_6575);
and U7133 (N_7133,N_6483,N_6754);
nor U7134 (N_7134,N_6569,N_6768);
nand U7135 (N_7135,N_6418,N_6445);
or U7136 (N_7136,N_6539,N_6550);
nand U7137 (N_7137,N_6412,N_6282);
nor U7138 (N_7138,N_6562,N_6708);
nand U7139 (N_7139,N_6772,N_6473);
nor U7140 (N_7140,N_6398,N_6568);
or U7141 (N_7141,N_6704,N_6384);
nand U7142 (N_7142,N_6654,N_6561);
nor U7143 (N_7143,N_6443,N_6375);
or U7144 (N_7144,N_6706,N_6763);
and U7145 (N_7145,N_6312,N_6479);
nand U7146 (N_7146,N_6846,N_6753);
nand U7147 (N_7147,N_6788,N_6434);
or U7148 (N_7148,N_6512,N_6334);
and U7149 (N_7149,N_6761,N_6806);
nor U7150 (N_7150,N_6604,N_6740);
nor U7151 (N_7151,N_6520,N_6823);
or U7152 (N_7152,N_6859,N_6372);
or U7153 (N_7153,N_6431,N_6305);
or U7154 (N_7154,N_6822,N_6636);
or U7155 (N_7155,N_6817,N_6665);
nor U7156 (N_7156,N_6399,N_6532);
nand U7157 (N_7157,N_6252,N_6407);
and U7158 (N_7158,N_6570,N_6421);
and U7159 (N_7159,N_6389,N_6486);
and U7160 (N_7160,N_6666,N_6524);
and U7161 (N_7161,N_6671,N_6835);
and U7162 (N_7162,N_6281,N_6750);
xnor U7163 (N_7163,N_6307,N_6821);
nand U7164 (N_7164,N_6804,N_6827);
xor U7165 (N_7165,N_6574,N_6690);
nor U7166 (N_7166,N_6382,N_6726);
nand U7167 (N_7167,N_6476,N_6263);
xor U7168 (N_7168,N_6651,N_6748);
xnor U7169 (N_7169,N_6423,N_6309);
or U7170 (N_7170,N_6760,N_6870);
or U7171 (N_7171,N_6755,N_6429);
nor U7172 (N_7172,N_6261,N_6438);
or U7173 (N_7173,N_6408,N_6633);
nand U7174 (N_7174,N_6738,N_6467);
and U7175 (N_7175,N_6630,N_6803);
nor U7176 (N_7176,N_6697,N_6463);
nor U7177 (N_7177,N_6351,N_6733);
xnor U7178 (N_7178,N_6257,N_6437);
nor U7179 (N_7179,N_6531,N_6848);
and U7180 (N_7180,N_6596,N_6459);
and U7181 (N_7181,N_6771,N_6293);
or U7182 (N_7182,N_6695,N_6449);
and U7183 (N_7183,N_6303,N_6488);
and U7184 (N_7184,N_6781,N_6251);
nor U7185 (N_7185,N_6638,N_6328);
nand U7186 (N_7186,N_6481,N_6523);
nor U7187 (N_7187,N_6653,N_6594);
or U7188 (N_7188,N_6373,N_6735);
and U7189 (N_7189,N_6562,N_6442);
nand U7190 (N_7190,N_6727,N_6266);
nor U7191 (N_7191,N_6862,N_6334);
nand U7192 (N_7192,N_6754,N_6657);
or U7193 (N_7193,N_6653,N_6456);
nand U7194 (N_7194,N_6483,N_6321);
and U7195 (N_7195,N_6310,N_6319);
and U7196 (N_7196,N_6444,N_6250);
and U7197 (N_7197,N_6727,N_6362);
nand U7198 (N_7198,N_6543,N_6434);
and U7199 (N_7199,N_6563,N_6556);
nand U7200 (N_7200,N_6322,N_6841);
or U7201 (N_7201,N_6282,N_6349);
nor U7202 (N_7202,N_6471,N_6554);
nand U7203 (N_7203,N_6561,N_6795);
xor U7204 (N_7204,N_6353,N_6735);
or U7205 (N_7205,N_6544,N_6767);
nand U7206 (N_7206,N_6663,N_6484);
nand U7207 (N_7207,N_6656,N_6417);
nor U7208 (N_7208,N_6408,N_6554);
or U7209 (N_7209,N_6284,N_6468);
xnor U7210 (N_7210,N_6579,N_6641);
or U7211 (N_7211,N_6359,N_6331);
or U7212 (N_7212,N_6286,N_6847);
xnor U7213 (N_7213,N_6663,N_6785);
and U7214 (N_7214,N_6854,N_6774);
and U7215 (N_7215,N_6649,N_6397);
nor U7216 (N_7216,N_6452,N_6835);
or U7217 (N_7217,N_6677,N_6434);
and U7218 (N_7218,N_6796,N_6530);
nor U7219 (N_7219,N_6607,N_6469);
or U7220 (N_7220,N_6817,N_6347);
nor U7221 (N_7221,N_6308,N_6327);
or U7222 (N_7222,N_6331,N_6353);
or U7223 (N_7223,N_6656,N_6296);
nand U7224 (N_7224,N_6334,N_6400);
or U7225 (N_7225,N_6311,N_6429);
or U7226 (N_7226,N_6461,N_6826);
nor U7227 (N_7227,N_6601,N_6530);
or U7228 (N_7228,N_6835,N_6291);
or U7229 (N_7229,N_6751,N_6676);
and U7230 (N_7230,N_6298,N_6750);
nand U7231 (N_7231,N_6762,N_6269);
xnor U7232 (N_7232,N_6771,N_6642);
nor U7233 (N_7233,N_6494,N_6412);
nor U7234 (N_7234,N_6268,N_6271);
or U7235 (N_7235,N_6681,N_6413);
nand U7236 (N_7236,N_6545,N_6364);
or U7237 (N_7237,N_6792,N_6416);
nand U7238 (N_7238,N_6530,N_6315);
and U7239 (N_7239,N_6447,N_6370);
nor U7240 (N_7240,N_6664,N_6480);
nand U7241 (N_7241,N_6341,N_6252);
or U7242 (N_7242,N_6365,N_6255);
nor U7243 (N_7243,N_6342,N_6427);
nor U7244 (N_7244,N_6745,N_6765);
nand U7245 (N_7245,N_6300,N_6364);
or U7246 (N_7246,N_6549,N_6751);
nor U7247 (N_7247,N_6690,N_6389);
xor U7248 (N_7248,N_6485,N_6350);
or U7249 (N_7249,N_6823,N_6463);
and U7250 (N_7250,N_6287,N_6787);
nand U7251 (N_7251,N_6259,N_6437);
or U7252 (N_7252,N_6362,N_6321);
nor U7253 (N_7253,N_6824,N_6524);
or U7254 (N_7254,N_6356,N_6852);
xor U7255 (N_7255,N_6575,N_6327);
nand U7256 (N_7256,N_6361,N_6350);
nor U7257 (N_7257,N_6788,N_6589);
and U7258 (N_7258,N_6685,N_6824);
and U7259 (N_7259,N_6275,N_6496);
and U7260 (N_7260,N_6845,N_6497);
nand U7261 (N_7261,N_6780,N_6643);
or U7262 (N_7262,N_6607,N_6405);
and U7263 (N_7263,N_6668,N_6523);
or U7264 (N_7264,N_6467,N_6397);
nor U7265 (N_7265,N_6808,N_6565);
and U7266 (N_7266,N_6454,N_6825);
nand U7267 (N_7267,N_6475,N_6488);
nor U7268 (N_7268,N_6481,N_6857);
nor U7269 (N_7269,N_6430,N_6329);
nand U7270 (N_7270,N_6640,N_6367);
and U7271 (N_7271,N_6853,N_6438);
nand U7272 (N_7272,N_6385,N_6596);
or U7273 (N_7273,N_6311,N_6313);
xnor U7274 (N_7274,N_6455,N_6511);
nor U7275 (N_7275,N_6572,N_6555);
nor U7276 (N_7276,N_6631,N_6784);
or U7277 (N_7277,N_6549,N_6852);
or U7278 (N_7278,N_6655,N_6647);
and U7279 (N_7279,N_6353,N_6467);
and U7280 (N_7280,N_6580,N_6313);
nand U7281 (N_7281,N_6838,N_6381);
or U7282 (N_7282,N_6391,N_6346);
or U7283 (N_7283,N_6802,N_6516);
and U7284 (N_7284,N_6333,N_6554);
and U7285 (N_7285,N_6621,N_6657);
nand U7286 (N_7286,N_6434,N_6774);
nand U7287 (N_7287,N_6587,N_6814);
or U7288 (N_7288,N_6835,N_6492);
and U7289 (N_7289,N_6699,N_6406);
nand U7290 (N_7290,N_6621,N_6437);
nand U7291 (N_7291,N_6469,N_6257);
xnor U7292 (N_7292,N_6672,N_6785);
and U7293 (N_7293,N_6283,N_6849);
and U7294 (N_7294,N_6308,N_6468);
and U7295 (N_7295,N_6652,N_6514);
or U7296 (N_7296,N_6467,N_6443);
nand U7297 (N_7297,N_6576,N_6500);
and U7298 (N_7298,N_6775,N_6813);
and U7299 (N_7299,N_6464,N_6782);
or U7300 (N_7300,N_6836,N_6454);
xor U7301 (N_7301,N_6377,N_6292);
xnor U7302 (N_7302,N_6826,N_6311);
nor U7303 (N_7303,N_6282,N_6586);
and U7304 (N_7304,N_6468,N_6587);
nor U7305 (N_7305,N_6758,N_6787);
or U7306 (N_7306,N_6606,N_6502);
nor U7307 (N_7307,N_6681,N_6628);
xor U7308 (N_7308,N_6695,N_6333);
nand U7309 (N_7309,N_6530,N_6382);
xor U7310 (N_7310,N_6708,N_6604);
nand U7311 (N_7311,N_6660,N_6633);
nand U7312 (N_7312,N_6680,N_6796);
xor U7313 (N_7313,N_6817,N_6747);
and U7314 (N_7314,N_6364,N_6600);
or U7315 (N_7315,N_6373,N_6362);
or U7316 (N_7316,N_6446,N_6298);
and U7317 (N_7317,N_6503,N_6704);
and U7318 (N_7318,N_6616,N_6765);
and U7319 (N_7319,N_6598,N_6455);
or U7320 (N_7320,N_6713,N_6873);
xnor U7321 (N_7321,N_6442,N_6793);
or U7322 (N_7322,N_6672,N_6323);
and U7323 (N_7323,N_6623,N_6820);
xnor U7324 (N_7324,N_6464,N_6385);
nand U7325 (N_7325,N_6355,N_6785);
nor U7326 (N_7326,N_6345,N_6827);
nand U7327 (N_7327,N_6650,N_6826);
nand U7328 (N_7328,N_6371,N_6562);
xnor U7329 (N_7329,N_6498,N_6736);
nand U7330 (N_7330,N_6393,N_6253);
nor U7331 (N_7331,N_6265,N_6751);
and U7332 (N_7332,N_6578,N_6374);
nor U7333 (N_7333,N_6395,N_6489);
nand U7334 (N_7334,N_6548,N_6673);
or U7335 (N_7335,N_6407,N_6665);
and U7336 (N_7336,N_6824,N_6596);
and U7337 (N_7337,N_6337,N_6571);
or U7338 (N_7338,N_6295,N_6572);
nor U7339 (N_7339,N_6765,N_6612);
nand U7340 (N_7340,N_6610,N_6836);
or U7341 (N_7341,N_6270,N_6363);
nor U7342 (N_7342,N_6822,N_6803);
nand U7343 (N_7343,N_6678,N_6450);
xor U7344 (N_7344,N_6806,N_6788);
or U7345 (N_7345,N_6568,N_6272);
or U7346 (N_7346,N_6713,N_6869);
xnor U7347 (N_7347,N_6729,N_6634);
and U7348 (N_7348,N_6471,N_6311);
or U7349 (N_7349,N_6478,N_6871);
and U7350 (N_7350,N_6468,N_6519);
nor U7351 (N_7351,N_6428,N_6556);
nand U7352 (N_7352,N_6870,N_6552);
nand U7353 (N_7353,N_6556,N_6295);
nor U7354 (N_7354,N_6357,N_6824);
nand U7355 (N_7355,N_6727,N_6281);
xor U7356 (N_7356,N_6366,N_6825);
nor U7357 (N_7357,N_6476,N_6685);
or U7358 (N_7358,N_6519,N_6574);
or U7359 (N_7359,N_6864,N_6761);
and U7360 (N_7360,N_6584,N_6620);
or U7361 (N_7361,N_6790,N_6820);
nor U7362 (N_7362,N_6653,N_6473);
or U7363 (N_7363,N_6837,N_6367);
and U7364 (N_7364,N_6350,N_6347);
or U7365 (N_7365,N_6267,N_6574);
nand U7366 (N_7366,N_6633,N_6857);
nand U7367 (N_7367,N_6677,N_6264);
xnor U7368 (N_7368,N_6558,N_6541);
nor U7369 (N_7369,N_6759,N_6741);
or U7370 (N_7370,N_6759,N_6510);
xnor U7371 (N_7371,N_6554,N_6421);
xnor U7372 (N_7372,N_6580,N_6528);
nor U7373 (N_7373,N_6282,N_6524);
and U7374 (N_7374,N_6505,N_6384);
or U7375 (N_7375,N_6567,N_6375);
and U7376 (N_7376,N_6326,N_6815);
nand U7377 (N_7377,N_6354,N_6733);
nor U7378 (N_7378,N_6454,N_6542);
and U7379 (N_7379,N_6341,N_6865);
or U7380 (N_7380,N_6647,N_6357);
or U7381 (N_7381,N_6613,N_6783);
or U7382 (N_7382,N_6745,N_6426);
or U7383 (N_7383,N_6287,N_6872);
nor U7384 (N_7384,N_6717,N_6347);
and U7385 (N_7385,N_6326,N_6738);
nand U7386 (N_7386,N_6807,N_6506);
or U7387 (N_7387,N_6737,N_6505);
and U7388 (N_7388,N_6506,N_6284);
nand U7389 (N_7389,N_6517,N_6602);
xnor U7390 (N_7390,N_6783,N_6569);
xnor U7391 (N_7391,N_6685,N_6769);
nand U7392 (N_7392,N_6605,N_6387);
or U7393 (N_7393,N_6503,N_6754);
nor U7394 (N_7394,N_6645,N_6261);
and U7395 (N_7395,N_6633,N_6809);
nor U7396 (N_7396,N_6523,N_6795);
xor U7397 (N_7397,N_6313,N_6593);
nor U7398 (N_7398,N_6641,N_6449);
nor U7399 (N_7399,N_6280,N_6745);
and U7400 (N_7400,N_6278,N_6446);
nand U7401 (N_7401,N_6296,N_6371);
nor U7402 (N_7402,N_6508,N_6265);
nor U7403 (N_7403,N_6818,N_6672);
or U7404 (N_7404,N_6679,N_6753);
or U7405 (N_7405,N_6658,N_6560);
xor U7406 (N_7406,N_6751,N_6477);
or U7407 (N_7407,N_6496,N_6274);
nand U7408 (N_7408,N_6430,N_6464);
or U7409 (N_7409,N_6375,N_6722);
nand U7410 (N_7410,N_6574,N_6791);
nand U7411 (N_7411,N_6819,N_6739);
or U7412 (N_7412,N_6301,N_6273);
or U7413 (N_7413,N_6612,N_6838);
or U7414 (N_7414,N_6368,N_6620);
and U7415 (N_7415,N_6672,N_6533);
or U7416 (N_7416,N_6371,N_6262);
nor U7417 (N_7417,N_6668,N_6452);
and U7418 (N_7418,N_6330,N_6814);
nand U7419 (N_7419,N_6758,N_6437);
nor U7420 (N_7420,N_6711,N_6561);
nor U7421 (N_7421,N_6461,N_6487);
nand U7422 (N_7422,N_6821,N_6416);
and U7423 (N_7423,N_6775,N_6777);
and U7424 (N_7424,N_6455,N_6313);
or U7425 (N_7425,N_6287,N_6565);
nor U7426 (N_7426,N_6393,N_6261);
or U7427 (N_7427,N_6557,N_6612);
and U7428 (N_7428,N_6282,N_6525);
nor U7429 (N_7429,N_6518,N_6389);
xnor U7430 (N_7430,N_6514,N_6726);
or U7431 (N_7431,N_6269,N_6529);
nor U7432 (N_7432,N_6872,N_6506);
and U7433 (N_7433,N_6456,N_6821);
nor U7434 (N_7434,N_6337,N_6666);
and U7435 (N_7435,N_6342,N_6524);
or U7436 (N_7436,N_6484,N_6497);
nor U7437 (N_7437,N_6503,N_6845);
or U7438 (N_7438,N_6419,N_6351);
nor U7439 (N_7439,N_6752,N_6478);
and U7440 (N_7440,N_6402,N_6804);
nand U7441 (N_7441,N_6572,N_6372);
nor U7442 (N_7442,N_6594,N_6360);
nor U7443 (N_7443,N_6438,N_6805);
and U7444 (N_7444,N_6653,N_6449);
or U7445 (N_7445,N_6627,N_6541);
or U7446 (N_7446,N_6550,N_6407);
and U7447 (N_7447,N_6415,N_6612);
xor U7448 (N_7448,N_6605,N_6328);
or U7449 (N_7449,N_6734,N_6557);
nand U7450 (N_7450,N_6391,N_6297);
nor U7451 (N_7451,N_6677,N_6705);
nor U7452 (N_7452,N_6744,N_6667);
xnor U7453 (N_7453,N_6767,N_6660);
or U7454 (N_7454,N_6261,N_6712);
nand U7455 (N_7455,N_6640,N_6376);
nor U7456 (N_7456,N_6866,N_6411);
and U7457 (N_7457,N_6683,N_6331);
nand U7458 (N_7458,N_6835,N_6321);
or U7459 (N_7459,N_6601,N_6286);
nor U7460 (N_7460,N_6681,N_6298);
nor U7461 (N_7461,N_6862,N_6606);
nand U7462 (N_7462,N_6474,N_6655);
nand U7463 (N_7463,N_6808,N_6355);
and U7464 (N_7464,N_6645,N_6281);
or U7465 (N_7465,N_6501,N_6516);
nor U7466 (N_7466,N_6542,N_6376);
and U7467 (N_7467,N_6405,N_6827);
xor U7468 (N_7468,N_6463,N_6456);
and U7469 (N_7469,N_6280,N_6787);
or U7470 (N_7470,N_6339,N_6722);
nand U7471 (N_7471,N_6645,N_6567);
xor U7472 (N_7472,N_6268,N_6285);
nand U7473 (N_7473,N_6413,N_6415);
nand U7474 (N_7474,N_6796,N_6466);
nand U7475 (N_7475,N_6413,N_6548);
nor U7476 (N_7476,N_6576,N_6850);
xnor U7477 (N_7477,N_6604,N_6611);
nor U7478 (N_7478,N_6613,N_6355);
nand U7479 (N_7479,N_6312,N_6594);
xor U7480 (N_7480,N_6405,N_6822);
xnor U7481 (N_7481,N_6509,N_6467);
nor U7482 (N_7482,N_6488,N_6729);
nand U7483 (N_7483,N_6790,N_6569);
nor U7484 (N_7484,N_6725,N_6754);
xnor U7485 (N_7485,N_6254,N_6345);
nand U7486 (N_7486,N_6583,N_6699);
xnor U7487 (N_7487,N_6257,N_6373);
xnor U7488 (N_7488,N_6271,N_6346);
or U7489 (N_7489,N_6652,N_6575);
nand U7490 (N_7490,N_6296,N_6760);
xor U7491 (N_7491,N_6745,N_6265);
nand U7492 (N_7492,N_6804,N_6770);
and U7493 (N_7493,N_6852,N_6580);
nor U7494 (N_7494,N_6865,N_6324);
and U7495 (N_7495,N_6815,N_6263);
or U7496 (N_7496,N_6568,N_6812);
or U7497 (N_7497,N_6374,N_6658);
or U7498 (N_7498,N_6843,N_6332);
or U7499 (N_7499,N_6422,N_6332);
or U7500 (N_7500,N_7053,N_6906);
xor U7501 (N_7501,N_7137,N_7162);
or U7502 (N_7502,N_6981,N_6929);
nand U7503 (N_7503,N_6967,N_7394);
nor U7504 (N_7504,N_7485,N_7408);
and U7505 (N_7505,N_6994,N_7396);
nor U7506 (N_7506,N_7212,N_7089);
and U7507 (N_7507,N_6936,N_7406);
nand U7508 (N_7508,N_6979,N_7459);
nand U7509 (N_7509,N_7361,N_7470);
nand U7510 (N_7510,N_6974,N_7472);
and U7511 (N_7511,N_7224,N_6992);
nor U7512 (N_7512,N_7060,N_7287);
nand U7513 (N_7513,N_7034,N_7016);
or U7514 (N_7514,N_7302,N_7483);
nor U7515 (N_7515,N_6965,N_7079);
nor U7516 (N_7516,N_7109,N_7223);
nor U7517 (N_7517,N_7451,N_7431);
or U7518 (N_7518,N_6940,N_7471);
or U7519 (N_7519,N_7325,N_7036);
xnor U7520 (N_7520,N_7203,N_6950);
and U7521 (N_7521,N_7012,N_6968);
nor U7522 (N_7522,N_7161,N_7401);
nand U7523 (N_7523,N_6986,N_7388);
nor U7524 (N_7524,N_7186,N_7381);
or U7525 (N_7525,N_6895,N_7099);
and U7526 (N_7526,N_7258,N_7094);
or U7527 (N_7527,N_6921,N_7221);
and U7528 (N_7528,N_7321,N_7183);
nor U7529 (N_7529,N_6980,N_7192);
or U7530 (N_7530,N_6898,N_7081);
or U7531 (N_7531,N_7430,N_7250);
nand U7532 (N_7532,N_6947,N_6955);
and U7533 (N_7533,N_7432,N_7115);
nand U7534 (N_7534,N_7481,N_7433);
or U7535 (N_7535,N_7176,N_7142);
and U7536 (N_7536,N_7141,N_7469);
nand U7537 (N_7537,N_7309,N_7172);
and U7538 (N_7538,N_7131,N_7277);
xnor U7539 (N_7539,N_7157,N_7202);
nand U7540 (N_7540,N_7173,N_7316);
xor U7541 (N_7541,N_7256,N_7386);
xnor U7542 (N_7542,N_7140,N_7284);
xnor U7543 (N_7543,N_7123,N_7324);
and U7544 (N_7544,N_7415,N_6886);
nand U7545 (N_7545,N_7073,N_7083);
and U7546 (N_7546,N_6885,N_6908);
and U7547 (N_7547,N_7178,N_7063);
xnor U7548 (N_7548,N_7128,N_7006);
and U7549 (N_7549,N_7004,N_7498);
nor U7550 (N_7550,N_7370,N_7225);
or U7551 (N_7551,N_6878,N_7023);
or U7552 (N_7552,N_6995,N_7251);
and U7553 (N_7553,N_6917,N_7437);
xor U7554 (N_7554,N_6951,N_6931);
nor U7555 (N_7555,N_7477,N_7414);
and U7556 (N_7556,N_7475,N_7000);
or U7557 (N_7557,N_7416,N_7113);
nand U7558 (N_7558,N_6958,N_7064);
nor U7559 (N_7559,N_7241,N_7344);
and U7560 (N_7560,N_7228,N_7027);
nor U7561 (N_7561,N_7383,N_7208);
or U7562 (N_7562,N_7096,N_7299);
nand U7563 (N_7563,N_7440,N_7249);
nor U7564 (N_7564,N_7144,N_6920);
or U7565 (N_7565,N_7465,N_7378);
nand U7566 (N_7566,N_7181,N_7046);
nand U7567 (N_7567,N_6942,N_7118);
nor U7568 (N_7568,N_7008,N_6875);
nand U7569 (N_7569,N_6912,N_6930);
or U7570 (N_7570,N_7360,N_7418);
nor U7571 (N_7571,N_6991,N_6897);
xor U7572 (N_7572,N_7468,N_7400);
or U7573 (N_7573,N_7138,N_6879);
xnor U7574 (N_7574,N_7165,N_7281);
nand U7575 (N_7575,N_7493,N_7317);
nor U7576 (N_7576,N_7122,N_7411);
nor U7577 (N_7577,N_7276,N_7114);
xor U7578 (N_7578,N_7391,N_7037);
or U7579 (N_7579,N_7197,N_7043);
and U7580 (N_7580,N_7233,N_7005);
xnor U7581 (N_7581,N_7112,N_7319);
and U7582 (N_7582,N_6890,N_7308);
nor U7583 (N_7583,N_7413,N_7159);
nor U7584 (N_7584,N_6973,N_7442);
or U7585 (N_7585,N_6997,N_7438);
nand U7586 (N_7586,N_7078,N_7047);
and U7587 (N_7587,N_7369,N_7133);
and U7588 (N_7588,N_7041,N_6887);
and U7589 (N_7589,N_7048,N_7179);
nand U7590 (N_7590,N_7206,N_7279);
nor U7591 (N_7591,N_7232,N_6932);
nor U7592 (N_7592,N_7194,N_6959);
nor U7593 (N_7593,N_7017,N_7397);
nor U7594 (N_7594,N_7260,N_6978);
nor U7595 (N_7595,N_7007,N_7158);
and U7596 (N_7596,N_6952,N_7211);
and U7597 (N_7597,N_7262,N_7195);
nand U7598 (N_7598,N_7214,N_7387);
or U7599 (N_7599,N_7288,N_7134);
xor U7600 (N_7600,N_7356,N_7105);
nand U7601 (N_7601,N_7039,N_7090);
nor U7602 (N_7602,N_6934,N_7289);
nand U7603 (N_7603,N_7269,N_7296);
xor U7604 (N_7604,N_7188,N_7095);
nor U7605 (N_7605,N_7343,N_7051);
nor U7606 (N_7606,N_7312,N_7151);
or U7607 (N_7607,N_6933,N_7322);
or U7608 (N_7608,N_7375,N_7120);
nor U7609 (N_7609,N_7059,N_7033);
nand U7610 (N_7610,N_6998,N_6928);
or U7611 (N_7611,N_7399,N_7132);
or U7612 (N_7612,N_6901,N_6939);
and U7613 (N_7613,N_7110,N_7061);
nor U7614 (N_7614,N_6914,N_7290);
or U7615 (N_7615,N_7014,N_7499);
nand U7616 (N_7616,N_7353,N_7446);
and U7617 (N_7617,N_7291,N_7488);
nor U7618 (N_7618,N_7097,N_7001);
nand U7619 (N_7619,N_7200,N_7019);
or U7620 (N_7620,N_6888,N_7467);
and U7621 (N_7621,N_6883,N_7448);
xnor U7622 (N_7622,N_7462,N_7347);
nand U7623 (N_7623,N_6970,N_7272);
and U7624 (N_7624,N_7393,N_7247);
and U7625 (N_7625,N_7346,N_7489);
nor U7626 (N_7626,N_7243,N_7458);
nor U7627 (N_7627,N_6884,N_7231);
nand U7628 (N_7628,N_7242,N_6963);
and U7629 (N_7629,N_7328,N_7274);
xnor U7630 (N_7630,N_7234,N_6984);
xnor U7631 (N_7631,N_6922,N_7404);
xnor U7632 (N_7632,N_7170,N_6954);
nand U7633 (N_7633,N_6975,N_7320);
xnor U7634 (N_7634,N_7389,N_6961);
and U7635 (N_7635,N_7280,N_7169);
nor U7636 (N_7636,N_7246,N_7153);
nand U7637 (N_7637,N_7336,N_7257);
xnor U7638 (N_7638,N_7327,N_7003);
nor U7639 (N_7639,N_7310,N_7351);
nand U7640 (N_7640,N_6957,N_6880);
and U7641 (N_7641,N_6977,N_7130);
nand U7642 (N_7642,N_6988,N_7464);
xor U7643 (N_7643,N_7057,N_6949);
nand U7644 (N_7644,N_7456,N_7135);
nand U7645 (N_7645,N_7182,N_7248);
nor U7646 (N_7646,N_7439,N_7227);
and U7647 (N_7647,N_7392,N_7164);
nand U7648 (N_7648,N_7050,N_7149);
nor U7649 (N_7649,N_7226,N_7150);
or U7650 (N_7650,N_7075,N_6982);
nand U7651 (N_7651,N_7009,N_7354);
and U7652 (N_7652,N_7267,N_7038);
or U7653 (N_7653,N_7371,N_6935);
nor U7654 (N_7654,N_7230,N_7407);
or U7655 (N_7655,N_7055,N_6946);
or U7656 (N_7656,N_7330,N_7455);
nand U7657 (N_7657,N_7245,N_7444);
or U7658 (N_7658,N_7139,N_7434);
or U7659 (N_7659,N_7304,N_7395);
xnor U7660 (N_7660,N_7156,N_7306);
nand U7661 (N_7661,N_6923,N_7025);
nand U7662 (N_7662,N_7101,N_7349);
nand U7663 (N_7663,N_7201,N_7026);
nand U7664 (N_7664,N_7490,N_7103);
nor U7665 (N_7665,N_7368,N_7253);
and U7666 (N_7666,N_7457,N_7390);
and U7667 (N_7667,N_7146,N_7450);
nand U7668 (N_7668,N_7238,N_7335);
nor U7669 (N_7669,N_7239,N_7255);
nand U7670 (N_7670,N_7382,N_7205);
and U7671 (N_7671,N_7002,N_7196);
nand U7672 (N_7672,N_7365,N_7098);
nand U7673 (N_7673,N_6910,N_7152);
nand U7674 (N_7674,N_7031,N_7340);
xor U7675 (N_7675,N_7435,N_7424);
nand U7676 (N_7676,N_7069,N_7010);
or U7677 (N_7677,N_7492,N_6987);
nand U7678 (N_7678,N_7207,N_7417);
nand U7679 (N_7679,N_7121,N_7129);
nand U7680 (N_7680,N_6926,N_7405);
xor U7681 (N_7681,N_7385,N_7292);
nand U7682 (N_7682,N_7028,N_7236);
nor U7683 (N_7683,N_6941,N_6989);
nand U7684 (N_7684,N_7426,N_6971);
and U7685 (N_7685,N_7333,N_7486);
nor U7686 (N_7686,N_7314,N_7092);
xnor U7687 (N_7687,N_7445,N_7199);
xor U7688 (N_7688,N_6976,N_7358);
nand U7689 (N_7689,N_7478,N_7266);
or U7690 (N_7690,N_6944,N_6945);
xnor U7691 (N_7691,N_7022,N_7357);
xor U7692 (N_7692,N_6907,N_7240);
or U7693 (N_7693,N_7072,N_7348);
nor U7694 (N_7694,N_7254,N_7185);
nand U7695 (N_7695,N_7111,N_7222);
or U7696 (N_7696,N_7497,N_7070);
xor U7697 (N_7697,N_7373,N_7029);
xor U7698 (N_7698,N_7337,N_7119);
nor U7699 (N_7699,N_7436,N_7275);
and U7700 (N_7700,N_7155,N_7487);
or U7701 (N_7701,N_7303,N_7187);
and U7702 (N_7702,N_7077,N_7174);
and U7703 (N_7703,N_7482,N_7116);
or U7704 (N_7704,N_7315,N_7474);
or U7705 (N_7705,N_6889,N_7024);
or U7706 (N_7706,N_7035,N_7419);
and U7707 (N_7707,N_7447,N_7441);
and U7708 (N_7708,N_7218,N_7127);
nand U7709 (N_7709,N_6902,N_7409);
xor U7710 (N_7710,N_7147,N_7429);
or U7711 (N_7711,N_7449,N_7091);
and U7712 (N_7712,N_7124,N_7421);
and U7713 (N_7713,N_7367,N_7331);
or U7714 (N_7714,N_7329,N_7190);
or U7715 (N_7715,N_7496,N_7076);
nor U7716 (N_7716,N_7494,N_6913);
nor U7717 (N_7717,N_7282,N_7184);
nand U7718 (N_7718,N_7332,N_7220);
nand U7719 (N_7719,N_7452,N_7189);
xor U7720 (N_7720,N_6962,N_7460);
nand U7721 (N_7721,N_7160,N_7476);
nor U7722 (N_7722,N_7093,N_6916);
nand U7723 (N_7723,N_7366,N_7300);
and U7724 (N_7724,N_7219,N_6905);
nand U7725 (N_7725,N_7177,N_6948);
xnor U7726 (N_7726,N_7273,N_7066);
nand U7727 (N_7727,N_7334,N_6911);
nand U7728 (N_7728,N_7350,N_7052);
and U7729 (N_7729,N_7237,N_6915);
nand U7730 (N_7730,N_6938,N_6985);
nor U7731 (N_7731,N_7355,N_6927);
and U7732 (N_7732,N_7425,N_7215);
nand U7733 (N_7733,N_7056,N_7217);
nand U7734 (N_7734,N_7163,N_7252);
nor U7735 (N_7735,N_7085,N_7326);
nor U7736 (N_7736,N_7168,N_7484);
nand U7737 (N_7737,N_7032,N_7084);
and U7738 (N_7738,N_7108,N_6881);
xnor U7739 (N_7739,N_7209,N_7305);
and U7740 (N_7740,N_7293,N_6972);
nor U7741 (N_7741,N_7175,N_7244);
nand U7742 (N_7742,N_7145,N_7363);
nand U7743 (N_7743,N_6925,N_7270);
or U7744 (N_7744,N_7171,N_7067);
nor U7745 (N_7745,N_7479,N_7271);
or U7746 (N_7746,N_7454,N_7427);
nor U7747 (N_7747,N_7412,N_7384);
nand U7748 (N_7748,N_7107,N_7210);
nor U7749 (N_7749,N_6877,N_7313);
and U7750 (N_7750,N_7088,N_7443);
nor U7751 (N_7751,N_7082,N_7285);
and U7752 (N_7752,N_7264,N_6909);
nor U7753 (N_7753,N_6999,N_7420);
xor U7754 (N_7754,N_7154,N_7461);
and U7755 (N_7755,N_7278,N_7087);
nor U7756 (N_7756,N_7374,N_7044);
xnor U7757 (N_7757,N_6918,N_7229);
or U7758 (N_7758,N_6893,N_7402);
or U7759 (N_7759,N_6996,N_6993);
xnor U7760 (N_7760,N_7311,N_7125);
and U7761 (N_7761,N_7359,N_7198);
and U7762 (N_7762,N_7259,N_7398);
and U7763 (N_7763,N_7377,N_7216);
or U7764 (N_7764,N_7167,N_7191);
nand U7765 (N_7765,N_7065,N_6990);
or U7766 (N_7766,N_6899,N_7166);
and U7767 (N_7767,N_6876,N_7018);
nor U7768 (N_7768,N_7015,N_7042);
or U7769 (N_7769,N_7491,N_6900);
nand U7770 (N_7770,N_7283,N_7045);
or U7771 (N_7771,N_7054,N_7058);
and U7772 (N_7772,N_7193,N_6903);
or U7773 (N_7773,N_7339,N_7148);
or U7774 (N_7774,N_7213,N_7013);
nand U7775 (N_7775,N_7380,N_7074);
and U7776 (N_7776,N_7341,N_7071);
or U7777 (N_7777,N_6953,N_7463);
and U7778 (N_7778,N_7080,N_6892);
or U7779 (N_7779,N_7345,N_6956);
nor U7780 (N_7780,N_6894,N_7466);
or U7781 (N_7781,N_7453,N_7235);
or U7782 (N_7782,N_7263,N_7480);
nand U7783 (N_7783,N_7030,N_7410);
nand U7784 (N_7784,N_7352,N_7143);
nand U7785 (N_7785,N_6964,N_7265);
nor U7786 (N_7786,N_7102,N_7104);
nand U7787 (N_7787,N_7126,N_7180);
or U7788 (N_7788,N_7376,N_6924);
or U7789 (N_7789,N_6891,N_6969);
nor U7790 (N_7790,N_7423,N_7100);
or U7791 (N_7791,N_7379,N_7307);
nand U7792 (N_7792,N_7261,N_7318);
and U7793 (N_7793,N_7049,N_7428);
nor U7794 (N_7794,N_7020,N_6960);
xnor U7795 (N_7795,N_7323,N_6882);
or U7796 (N_7796,N_7338,N_7473);
and U7797 (N_7797,N_7286,N_6937);
nand U7798 (N_7798,N_7294,N_7040);
nor U7799 (N_7799,N_6983,N_7117);
or U7800 (N_7800,N_7298,N_7495);
and U7801 (N_7801,N_7372,N_7086);
nor U7802 (N_7802,N_7422,N_7268);
xnor U7803 (N_7803,N_7403,N_7021);
nand U7804 (N_7804,N_7297,N_7204);
nand U7805 (N_7805,N_7295,N_7068);
or U7806 (N_7806,N_6919,N_6943);
or U7807 (N_7807,N_6904,N_7301);
nor U7808 (N_7808,N_7362,N_7011);
or U7809 (N_7809,N_7364,N_6966);
nor U7810 (N_7810,N_7342,N_7062);
nor U7811 (N_7811,N_7106,N_7136);
nand U7812 (N_7812,N_6896,N_7220);
and U7813 (N_7813,N_7115,N_7485);
xnor U7814 (N_7814,N_7428,N_6928);
or U7815 (N_7815,N_7044,N_7258);
or U7816 (N_7816,N_7124,N_6914);
or U7817 (N_7817,N_6929,N_6966);
xnor U7818 (N_7818,N_7071,N_7249);
or U7819 (N_7819,N_7395,N_7355);
and U7820 (N_7820,N_7172,N_6926);
nand U7821 (N_7821,N_7185,N_7238);
or U7822 (N_7822,N_7290,N_7269);
nor U7823 (N_7823,N_7396,N_7188);
nand U7824 (N_7824,N_7111,N_7419);
nor U7825 (N_7825,N_7346,N_7340);
nand U7826 (N_7826,N_6950,N_7238);
and U7827 (N_7827,N_7474,N_6917);
and U7828 (N_7828,N_7092,N_7231);
and U7829 (N_7829,N_7434,N_7171);
nor U7830 (N_7830,N_6911,N_6908);
and U7831 (N_7831,N_7288,N_7249);
nand U7832 (N_7832,N_6914,N_7229);
and U7833 (N_7833,N_7116,N_7104);
xor U7834 (N_7834,N_7249,N_7018);
or U7835 (N_7835,N_7090,N_7450);
or U7836 (N_7836,N_7415,N_7456);
or U7837 (N_7837,N_7459,N_7013);
nor U7838 (N_7838,N_7034,N_7358);
nand U7839 (N_7839,N_7032,N_7240);
and U7840 (N_7840,N_7191,N_6997);
or U7841 (N_7841,N_6924,N_7091);
and U7842 (N_7842,N_6982,N_6975);
or U7843 (N_7843,N_7441,N_7462);
xor U7844 (N_7844,N_7183,N_7004);
nor U7845 (N_7845,N_7134,N_7377);
nor U7846 (N_7846,N_7218,N_6886);
nand U7847 (N_7847,N_7056,N_6979);
xor U7848 (N_7848,N_6926,N_7468);
or U7849 (N_7849,N_7468,N_7451);
or U7850 (N_7850,N_7090,N_7127);
nand U7851 (N_7851,N_6951,N_7155);
or U7852 (N_7852,N_7337,N_6999);
nand U7853 (N_7853,N_7410,N_7362);
nand U7854 (N_7854,N_7093,N_7436);
nor U7855 (N_7855,N_7479,N_7160);
nand U7856 (N_7856,N_7243,N_6995);
and U7857 (N_7857,N_7271,N_7452);
and U7858 (N_7858,N_7296,N_7422);
and U7859 (N_7859,N_7223,N_7145);
nand U7860 (N_7860,N_6976,N_7285);
nor U7861 (N_7861,N_7320,N_6987);
nand U7862 (N_7862,N_7021,N_6987);
nand U7863 (N_7863,N_7427,N_7166);
and U7864 (N_7864,N_7178,N_7040);
nand U7865 (N_7865,N_6999,N_7147);
and U7866 (N_7866,N_7134,N_7037);
and U7867 (N_7867,N_7322,N_7467);
or U7868 (N_7868,N_6977,N_6953);
and U7869 (N_7869,N_7397,N_7363);
and U7870 (N_7870,N_6951,N_7378);
nand U7871 (N_7871,N_7014,N_7476);
or U7872 (N_7872,N_7445,N_7359);
xnor U7873 (N_7873,N_7150,N_7201);
and U7874 (N_7874,N_7301,N_7019);
or U7875 (N_7875,N_7257,N_7260);
and U7876 (N_7876,N_7116,N_7410);
nand U7877 (N_7877,N_7199,N_7017);
or U7878 (N_7878,N_6943,N_7408);
and U7879 (N_7879,N_7374,N_7446);
nand U7880 (N_7880,N_7260,N_7008);
nor U7881 (N_7881,N_7247,N_7468);
or U7882 (N_7882,N_7498,N_6888);
nor U7883 (N_7883,N_6881,N_7163);
nor U7884 (N_7884,N_7189,N_7352);
nand U7885 (N_7885,N_6935,N_7131);
nor U7886 (N_7886,N_7251,N_7312);
xor U7887 (N_7887,N_7259,N_6939);
xnor U7888 (N_7888,N_7281,N_6984);
nor U7889 (N_7889,N_7398,N_7104);
and U7890 (N_7890,N_7192,N_7350);
xor U7891 (N_7891,N_7003,N_7132);
nand U7892 (N_7892,N_7243,N_6948);
and U7893 (N_7893,N_6986,N_6941);
and U7894 (N_7894,N_6895,N_7185);
and U7895 (N_7895,N_7096,N_7119);
xnor U7896 (N_7896,N_6962,N_7162);
or U7897 (N_7897,N_7393,N_7076);
nor U7898 (N_7898,N_7278,N_7318);
and U7899 (N_7899,N_6876,N_7152);
or U7900 (N_7900,N_7102,N_7368);
nor U7901 (N_7901,N_7099,N_7070);
and U7902 (N_7902,N_7316,N_7229);
or U7903 (N_7903,N_6933,N_7032);
or U7904 (N_7904,N_7246,N_6998);
and U7905 (N_7905,N_7184,N_7120);
nor U7906 (N_7906,N_6962,N_7417);
xnor U7907 (N_7907,N_7379,N_6920);
and U7908 (N_7908,N_6976,N_7348);
nand U7909 (N_7909,N_7283,N_6938);
xor U7910 (N_7910,N_7219,N_6962);
or U7911 (N_7911,N_7434,N_6999);
or U7912 (N_7912,N_7084,N_7230);
or U7913 (N_7913,N_7378,N_6942);
nor U7914 (N_7914,N_7160,N_7214);
nor U7915 (N_7915,N_6910,N_7170);
nor U7916 (N_7916,N_7045,N_7083);
or U7917 (N_7917,N_6917,N_7296);
nor U7918 (N_7918,N_7160,N_7262);
nor U7919 (N_7919,N_7369,N_7045);
nor U7920 (N_7920,N_7361,N_6952);
nand U7921 (N_7921,N_7030,N_7472);
nor U7922 (N_7922,N_7298,N_7267);
or U7923 (N_7923,N_7221,N_7203);
nor U7924 (N_7924,N_7135,N_6978);
or U7925 (N_7925,N_7133,N_7466);
and U7926 (N_7926,N_7346,N_7218);
nand U7927 (N_7927,N_7347,N_6985);
and U7928 (N_7928,N_7254,N_6997);
and U7929 (N_7929,N_7399,N_7081);
nand U7930 (N_7930,N_7363,N_6953);
and U7931 (N_7931,N_7314,N_7263);
nand U7932 (N_7932,N_7218,N_6972);
nor U7933 (N_7933,N_7475,N_6966);
or U7934 (N_7934,N_7318,N_7204);
or U7935 (N_7935,N_7076,N_7236);
nand U7936 (N_7936,N_7193,N_7060);
nand U7937 (N_7937,N_7319,N_7080);
xor U7938 (N_7938,N_7362,N_7190);
and U7939 (N_7939,N_7290,N_7141);
nand U7940 (N_7940,N_7306,N_7076);
or U7941 (N_7941,N_7173,N_7384);
nor U7942 (N_7942,N_6910,N_6892);
and U7943 (N_7943,N_7216,N_7073);
and U7944 (N_7944,N_7342,N_7272);
and U7945 (N_7945,N_7074,N_7240);
xor U7946 (N_7946,N_7129,N_7120);
nand U7947 (N_7947,N_6995,N_7026);
nand U7948 (N_7948,N_7439,N_7287);
nor U7949 (N_7949,N_7427,N_7297);
and U7950 (N_7950,N_6971,N_7413);
or U7951 (N_7951,N_7151,N_7063);
nor U7952 (N_7952,N_7311,N_7263);
nand U7953 (N_7953,N_7202,N_7178);
and U7954 (N_7954,N_7226,N_7345);
nand U7955 (N_7955,N_7050,N_7266);
or U7956 (N_7956,N_7318,N_7274);
and U7957 (N_7957,N_6973,N_7436);
and U7958 (N_7958,N_6941,N_6953);
nor U7959 (N_7959,N_6880,N_6893);
nand U7960 (N_7960,N_7304,N_7338);
or U7961 (N_7961,N_7237,N_7400);
and U7962 (N_7962,N_7049,N_7469);
nand U7963 (N_7963,N_7471,N_7027);
and U7964 (N_7964,N_7418,N_7122);
or U7965 (N_7965,N_7154,N_7447);
nor U7966 (N_7966,N_7079,N_7344);
and U7967 (N_7967,N_6926,N_6884);
nand U7968 (N_7968,N_7264,N_7034);
and U7969 (N_7969,N_7009,N_7179);
and U7970 (N_7970,N_7149,N_6931);
nand U7971 (N_7971,N_7363,N_6978);
or U7972 (N_7972,N_6893,N_6968);
nand U7973 (N_7973,N_7352,N_7058);
xnor U7974 (N_7974,N_7412,N_6957);
and U7975 (N_7975,N_7372,N_7300);
or U7976 (N_7976,N_6996,N_7148);
nand U7977 (N_7977,N_6966,N_7341);
nand U7978 (N_7978,N_7247,N_7074);
or U7979 (N_7979,N_7162,N_7443);
and U7980 (N_7980,N_7362,N_7080);
nand U7981 (N_7981,N_6922,N_7102);
and U7982 (N_7982,N_7431,N_6979);
or U7983 (N_7983,N_7191,N_7057);
xnor U7984 (N_7984,N_7129,N_7300);
nand U7985 (N_7985,N_7276,N_7020);
nand U7986 (N_7986,N_6953,N_7216);
and U7987 (N_7987,N_7227,N_7447);
xnor U7988 (N_7988,N_7085,N_7494);
and U7989 (N_7989,N_7127,N_6993);
and U7990 (N_7990,N_7457,N_7466);
or U7991 (N_7991,N_7171,N_7376);
or U7992 (N_7992,N_7293,N_7429);
nand U7993 (N_7993,N_7358,N_7055);
or U7994 (N_7994,N_7429,N_7077);
or U7995 (N_7995,N_7259,N_7387);
or U7996 (N_7996,N_7236,N_7195);
nor U7997 (N_7997,N_7046,N_7146);
nand U7998 (N_7998,N_7423,N_7168);
nand U7999 (N_7999,N_6964,N_7253);
or U8000 (N_8000,N_7434,N_7405);
or U8001 (N_8001,N_6975,N_7175);
or U8002 (N_8002,N_6950,N_7127);
nand U8003 (N_8003,N_7482,N_7114);
nand U8004 (N_8004,N_7100,N_7430);
and U8005 (N_8005,N_7103,N_6976);
nor U8006 (N_8006,N_7074,N_7037);
xnor U8007 (N_8007,N_6891,N_7345);
or U8008 (N_8008,N_7426,N_7129);
and U8009 (N_8009,N_6999,N_7063);
or U8010 (N_8010,N_6954,N_7016);
and U8011 (N_8011,N_7347,N_7090);
and U8012 (N_8012,N_7341,N_7255);
and U8013 (N_8013,N_7225,N_7306);
and U8014 (N_8014,N_7033,N_7090);
and U8015 (N_8015,N_7309,N_7239);
xor U8016 (N_8016,N_7294,N_7362);
nand U8017 (N_8017,N_7008,N_7215);
or U8018 (N_8018,N_6892,N_7386);
nor U8019 (N_8019,N_7036,N_7432);
and U8020 (N_8020,N_7167,N_7333);
or U8021 (N_8021,N_6941,N_6896);
nand U8022 (N_8022,N_6972,N_7144);
and U8023 (N_8023,N_7481,N_7198);
nor U8024 (N_8024,N_7447,N_7140);
nor U8025 (N_8025,N_7021,N_7236);
or U8026 (N_8026,N_7038,N_7032);
or U8027 (N_8027,N_7176,N_7001);
or U8028 (N_8028,N_7400,N_7241);
nand U8029 (N_8029,N_7017,N_6970);
nand U8030 (N_8030,N_7118,N_7082);
nor U8031 (N_8031,N_6960,N_7101);
nand U8032 (N_8032,N_7450,N_7028);
or U8033 (N_8033,N_7202,N_6920);
or U8034 (N_8034,N_6961,N_7335);
or U8035 (N_8035,N_7373,N_6896);
or U8036 (N_8036,N_7289,N_7181);
nand U8037 (N_8037,N_7196,N_6963);
and U8038 (N_8038,N_7137,N_7161);
nand U8039 (N_8039,N_6979,N_6926);
nand U8040 (N_8040,N_7268,N_7035);
and U8041 (N_8041,N_7187,N_7318);
nand U8042 (N_8042,N_7436,N_7434);
and U8043 (N_8043,N_7457,N_6966);
nand U8044 (N_8044,N_6988,N_7247);
nand U8045 (N_8045,N_7040,N_7108);
nor U8046 (N_8046,N_6930,N_6993);
nand U8047 (N_8047,N_7333,N_7373);
nor U8048 (N_8048,N_7270,N_7053);
or U8049 (N_8049,N_6899,N_7428);
nor U8050 (N_8050,N_6939,N_7253);
nor U8051 (N_8051,N_7063,N_7225);
xor U8052 (N_8052,N_7306,N_7087);
nor U8053 (N_8053,N_7286,N_7466);
and U8054 (N_8054,N_7196,N_6945);
and U8055 (N_8055,N_7366,N_7288);
and U8056 (N_8056,N_7438,N_6893);
and U8057 (N_8057,N_7125,N_6878);
nand U8058 (N_8058,N_7493,N_7314);
or U8059 (N_8059,N_7261,N_7243);
xnor U8060 (N_8060,N_7476,N_6970);
nor U8061 (N_8061,N_7140,N_6943);
nand U8062 (N_8062,N_7382,N_7418);
and U8063 (N_8063,N_7327,N_7474);
nor U8064 (N_8064,N_6922,N_6903);
or U8065 (N_8065,N_7197,N_7099);
or U8066 (N_8066,N_7044,N_7113);
or U8067 (N_8067,N_7127,N_7213);
and U8068 (N_8068,N_6886,N_7405);
xnor U8069 (N_8069,N_7163,N_7261);
and U8070 (N_8070,N_7165,N_7123);
nor U8071 (N_8071,N_7487,N_7330);
and U8072 (N_8072,N_7349,N_7014);
nor U8073 (N_8073,N_7246,N_7410);
or U8074 (N_8074,N_7050,N_7234);
or U8075 (N_8075,N_7129,N_7078);
or U8076 (N_8076,N_7438,N_6952);
nor U8077 (N_8077,N_7141,N_7188);
xor U8078 (N_8078,N_7205,N_6998);
nor U8079 (N_8079,N_7244,N_7355);
nand U8080 (N_8080,N_7224,N_7432);
nor U8081 (N_8081,N_7055,N_7197);
or U8082 (N_8082,N_6958,N_7243);
nand U8083 (N_8083,N_7270,N_7463);
or U8084 (N_8084,N_6958,N_7466);
and U8085 (N_8085,N_7397,N_7499);
xnor U8086 (N_8086,N_7186,N_7203);
nand U8087 (N_8087,N_7004,N_7275);
nor U8088 (N_8088,N_7046,N_7285);
or U8089 (N_8089,N_6877,N_7489);
nand U8090 (N_8090,N_7244,N_7077);
or U8091 (N_8091,N_7416,N_7193);
xor U8092 (N_8092,N_7463,N_7101);
nand U8093 (N_8093,N_7053,N_7259);
or U8094 (N_8094,N_7138,N_7122);
or U8095 (N_8095,N_7403,N_7250);
and U8096 (N_8096,N_7454,N_7179);
or U8097 (N_8097,N_7396,N_7280);
or U8098 (N_8098,N_7444,N_6927);
or U8099 (N_8099,N_7156,N_7186);
nor U8100 (N_8100,N_7478,N_6914);
nor U8101 (N_8101,N_7075,N_7337);
nor U8102 (N_8102,N_7404,N_6879);
and U8103 (N_8103,N_6932,N_7402);
nor U8104 (N_8104,N_7023,N_7180);
and U8105 (N_8105,N_7058,N_7411);
nor U8106 (N_8106,N_7257,N_7310);
nor U8107 (N_8107,N_7219,N_7436);
xor U8108 (N_8108,N_6929,N_7373);
nor U8109 (N_8109,N_7296,N_7136);
nor U8110 (N_8110,N_7410,N_7216);
or U8111 (N_8111,N_7399,N_7216);
nand U8112 (N_8112,N_6958,N_7086);
nand U8113 (N_8113,N_7311,N_6883);
and U8114 (N_8114,N_7109,N_6894);
nor U8115 (N_8115,N_7094,N_6952);
and U8116 (N_8116,N_7192,N_7273);
nand U8117 (N_8117,N_7381,N_7485);
nor U8118 (N_8118,N_7377,N_7180);
and U8119 (N_8119,N_7313,N_7010);
or U8120 (N_8120,N_7372,N_7016);
or U8121 (N_8121,N_7376,N_7313);
xnor U8122 (N_8122,N_7433,N_7215);
or U8123 (N_8123,N_7379,N_7346);
nor U8124 (N_8124,N_7159,N_7161);
and U8125 (N_8125,N_8054,N_8052);
xnor U8126 (N_8126,N_7814,N_7743);
xor U8127 (N_8127,N_7580,N_7761);
nor U8128 (N_8128,N_7944,N_7513);
and U8129 (N_8129,N_7689,N_7598);
nor U8130 (N_8130,N_7991,N_7934);
and U8131 (N_8131,N_7565,N_7587);
nand U8132 (N_8132,N_7854,N_8078);
nand U8133 (N_8133,N_7764,N_7521);
or U8134 (N_8134,N_7878,N_7635);
nand U8135 (N_8135,N_7977,N_7947);
or U8136 (N_8136,N_7683,N_7926);
nor U8137 (N_8137,N_8014,N_7954);
nor U8138 (N_8138,N_7584,N_7540);
or U8139 (N_8139,N_7653,N_7523);
xnor U8140 (N_8140,N_7789,N_7674);
and U8141 (N_8141,N_7711,N_7591);
xor U8142 (N_8142,N_7697,N_8081);
or U8143 (N_8143,N_7757,N_7881);
nand U8144 (N_8144,N_7514,N_7614);
and U8145 (N_8145,N_7869,N_7571);
nand U8146 (N_8146,N_7824,N_7604);
or U8147 (N_8147,N_7634,N_8109);
nand U8148 (N_8148,N_7682,N_7811);
nor U8149 (N_8149,N_7507,N_7626);
and U8150 (N_8150,N_7930,N_7651);
and U8151 (N_8151,N_7864,N_7596);
xnor U8152 (N_8152,N_8001,N_7517);
xor U8153 (N_8153,N_8107,N_7581);
or U8154 (N_8154,N_8119,N_7766);
or U8155 (N_8155,N_7974,N_7975);
nor U8156 (N_8156,N_7841,N_8008);
nor U8157 (N_8157,N_8029,N_7821);
or U8158 (N_8158,N_7780,N_7957);
nand U8159 (N_8159,N_8010,N_7891);
and U8160 (N_8160,N_7852,N_7893);
or U8161 (N_8161,N_7510,N_7818);
and U8162 (N_8162,N_7883,N_8103);
or U8163 (N_8163,N_7972,N_7532);
nand U8164 (N_8164,N_7589,N_7758);
xnor U8165 (N_8165,N_7552,N_7553);
nand U8166 (N_8166,N_7545,N_7943);
and U8167 (N_8167,N_7834,N_7680);
nand U8168 (N_8168,N_7809,N_8059);
nor U8169 (N_8169,N_7570,N_7833);
and U8170 (N_8170,N_7887,N_7739);
nor U8171 (N_8171,N_7942,N_8100);
nand U8172 (N_8172,N_8012,N_7950);
or U8173 (N_8173,N_7769,N_7686);
nor U8174 (N_8174,N_7923,N_7948);
nor U8175 (N_8175,N_7594,N_7906);
nor U8176 (N_8176,N_7855,N_8116);
and U8177 (N_8177,N_7667,N_8062);
nor U8178 (N_8178,N_7629,N_7772);
nand U8179 (N_8179,N_7694,N_7924);
or U8180 (N_8180,N_7753,N_7968);
xnor U8181 (N_8181,N_8011,N_8030);
nor U8182 (N_8182,N_8105,N_8117);
and U8183 (N_8183,N_8049,N_7831);
or U8184 (N_8184,N_7648,N_7819);
or U8185 (N_8185,N_7803,N_7666);
or U8186 (N_8186,N_7922,N_8053);
xor U8187 (N_8187,N_7982,N_7762);
or U8188 (N_8188,N_8077,N_7901);
and U8189 (N_8189,N_8047,N_7538);
and U8190 (N_8190,N_7732,N_7675);
or U8191 (N_8191,N_7765,N_7965);
nand U8192 (N_8192,N_7652,N_7701);
nor U8193 (N_8193,N_7700,N_7911);
or U8194 (N_8194,N_7870,N_7522);
or U8195 (N_8195,N_7506,N_7593);
or U8196 (N_8196,N_7736,N_7549);
nand U8197 (N_8197,N_7727,N_8006);
nor U8198 (N_8198,N_7610,N_8090);
nand U8199 (N_8199,N_8040,N_8036);
xnor U8200 (N_8200,N_7737,N_7751);
or U8201 (N_8201,N_7639,N_7823);
nor U8202 (N_8202,N_8041,N_7939);
nand U8203 (N_8203,N_7691,N_8114);
or U8204 (N_8204,N_7741,N_7961);
nor U8205 (N_8205,N_8028,N_7993);
nand U8206 (N_8206,N_8123,N_8021);
or U8207 (N_8207,N_8087,N_7734);
nor U8208 (N_8208,N_7778,N_7566);
nand U8209 (N_8209,N_7847,N_7768);
and U8210 (N_8210,N_7816,N_7738);
nor U8211 (N_8211,N_7949,N_8024);
nor U8212 (N_8212,N_7558,N_7546);
nor U8213 (N_8213,N_7815,N_7866);
or U8214 (N_8214,N_7863,N_8072);
or U8215 (N_8215,N_7735,N_7564);
xor U8216 (N_8216,N_7921,N_8018);
nor U8217 (N_8217,N_7868,N_7917);
or U8218 (N_8218,N_8073,N_7693);
and U8219 (N_8219,N_7657,N_7539);
nor U8220 (N_8220,N_7668,N_7642);
or U8221 (N_8221,N_8110,N_7937);
or U8222 (N_8222,N_7895,N_7919);
nor U8223 (N_8223,N_7918,N_8101);
nor U8224 (N_8224,N_7835,N_7588);
nand U8225 (N_8225,N_8102,N_8022);
and U8226 (N_8226,N_7952,N_7722);
nor U8227 (N_8227,N_7846,N_7608);
xnor U8228 (N_8228,N_8061,N_7621);
xor U8229 (N_8229,N_7720,N_7782);
or U8230 (N_8230,N_8113,N_7748);
nand U8231 (N_8231,N_7503,N_7873);
or U8232 (N_8232,N_7568,N_8060);
nand U8233 (N_8233,N_7533,N_8079);
nor U8234 (N_8234,N_7677,N_7801);
and U8235 (N_8235,N_7687,N_7670);
nand U8236 (N_8236,N_8120,N_7898);
or U8237 (N_8237,N_7663,N_7787);
or U8238 (N_8238,N_7638,N_7980);
nor U8239 (N_8239,N_8069,N_7890);
nor U8240 (N_8240,N_7829,N_8092);
xor U8241 (N_8241,N_8097,N_8046);
nor U8242 (N_8242,N_7632,N_7777);
and U8243 (N_8243,N_7573,N_7535);
nor U8244 (N_8244,N_7981,N_8082);
and U8245 (N_8245,N_8076,N_7690);
or U8246 (N_8246,N_7867,N_7526);
nor U8247 (N_8247,N_8118,N_8094);
nor U8248 (N_8248,N_7885,N_7515);
nand U8249 (N_8249,N_7994,N_7527);
xnor U8250 (N_8250,N_8074,N_7963);
nor U8251 (N_8251,N_7790,N_7628);
or U8252 (N_8252,N_7551,N_8065);
nor U8253 (N_8253,N_7894,N_7520);
nand U8254 (N_8254,N_7941,N_7665);
nand U8255 (N_8255,N_7599,N_7827);
nor U8256 (N_8256,N_7585,N_7574);
or U8257 (N_8257,N_7650,N_7932);
nand U8258 (N_8258,N_7595,N_7853);
or U8259 (N_8259,N_7724,N_7861);
or U8260 (N_8260,N_7547,N_7946);
or U8261 (N_8261,N_7541,N_7862);
nor U8262 (N_8262,N_7713,N_7910);
nand U8263 (N_8263,N_7630,N_7554);
nor U8264 (N_8264,N_7719,N_7605);
nor U8265 (N_8265,N_8095,N_7978);
nand U8266 (N_8266,N_7907,N_7904);
or U8267 (N_8267,N_7928,N_7839);
nand U8268 (N_8268,N_7899,N_8111);
nor U8269 (N_8269,N_8057,N_7583);
or U8270 (N_8270,N_7920,N_7804);
or U8271 (N_8271,N_7692,N_8017);
xor U8272 (N_8272,N_7637,N_8031);
nor U8273 (N_8273,N_7612,N_7592);
nor U8274 (N_8274,N_7783,N_7622);
nor U8275 (N_8275,N_7775,N_7579);
nor U8276 (N_8276,N_7643,N_8066);
and U8277 (N_8277,N_8013,N_7733);
or U8278 (N_8278,N_7703,N_8027);
and U8279 (N_8279,N_7791,N_7746);
nor U8280 (N_8280,N_7959,N_7865);
nor U8281 (N_8281,N_7685,N_7905);
nor U8282 (N_8282,N_7969,N_7884);
or U8283 (N_8283,N_8096,N_7618);
nand U8284 (N_8284,N_7500,N_7715);
nor U8285 (N_8285,N_7613,N_7970);
and U8286 (N_8286,N_7807,N_7508);
or U8287 (N_8287,N_8003,N_7509);
nand U8288 (N_8288,N_7914,N_7752);
nor U8289 (N_8289,N_8048,N_7984);
nor U8290 (N_8290,N_7813,N_7915);
nor U8291 (N_8291,N_7676,N_7976);
nor U8292 (N_8292,N_8115,N_7704);
nor U8293 (N_8293,N_7967,N_7874);
nand U8294 (N_8294,N_7543,N_7501);
or U8295 (N_8295,N_7792,N_7729);
nor U8296 (N_8296,N_7794,N_7616);
nor U8297 (N_8297,N_7871,N_7710);
or U8298 (N_8298,N_7983,N_7646);
nor U8299 (N_8299,N_7684,N_7875);
xnor U8300 (N_8300,N_7966,N_7913);
and U8301 (N_8301,N_7810,N_7808);
xor U8302 (N_8302,N_7945,N_7721);
or U8303 (N_8303,N_7857,N_7615);
and U8304 (N_8304,N_7902,N_8075);
or U8305 (N_8305,N_8083,N_7820);
nor U8306 (N_8306,N_8067,N_7623);
nor U8307 (N_8307,N_7633,N_7645);
nor U8308 (N_8308,N_7838,N_7900);
nor U8309 (N_8309,N_7601,N_8042);
or U8310 (N_8310,N_7531,N_7909);
or U8311 (N_8311,N_7837,N_7802);
xor U8312 (N_8312,N_7955,N_7673);
nand U8313 (N_8313,N_7577,N_7617);
and U8314 (N_8314,N_7903,N_7611);
and U8315 (N_8315,N_7848,N_7940);
nand U8316 (N_8316,N_7797,N_7962);
xnor U8317 (N_8317,N_8089,N_7896);
or U8318 (N_8318,N_7796,N_7826);
nor U8319 (N_8319,N_7858,N_7876);
nor U8320 (N_8320,N_7709,N_7785);
or U8321 (N_8321,N_7779,N_7985);
xnor U8322 (N_8322,N_7708,N_7516);
nor U8323 (N_8323,N_7597,N_7716);
nand U8324 (N_8324,N_7688,N_7951);
and U8325 (N_8325,N_7886,N_8038);
or U8326 (N_8326,N_7840,N_7747);
and U8327 (N_8327,N_7845,N_7851);
or U8328 (N_8328,N_7859,N_7992);
and U8329 (N_8329,N_7931,N_7882);
nor U8330 (N_8330,N_8000,N_7756);
nand U8331 (N_8331,N_7798,N_7936);
and U8332 (N_8332,N_8032,N_7781);
nand U8333 (N_8333,N_7759,N_8016);
nor U8334 (N_8334,N_7627,N_8063);
or U8335 (N_8335,N_7836,N_8108);
nor U8336 (N_8336,N_7609,N_7528);
and U8337 (N_8337,N_7695,N_7679);
nor U8338 (N_8338,N_8068,N_7519);
nor U8339 (N_8339,N_7832,N_7795);
nand U8340 (N_8340,N_7825,N_7561);
and U8341 (N_8341,N_7644,N_7767);
nor U8342 (N_8342,N_8035,N_7938);
nor U8343 (N_8343,N_7872,N_7760);
nor U8344 (N_8344,N_7830,N_7953);
or U8345 (N_8345,N_7534,N_7771);
nor U8346 (N_8346,N_7625,N_7712);
nor U8347 (N_8347,N_7860,N_7671);
nor U8348 (N_8348,N_8086,N_7569);
or U8349 (N_8349,N_7536,N_7925);
nand U8350 (N_8350,N_8055,N_8112);
nor U8351 (N_8351,N_7660,N_7927);
nor U8352 (N_8352,N_7559,N_7731);
nand U8353 (N_8353,N_7603,N_7850);
xnor U8354 (N_8354,N_7742,N_7664);
nand U8355 (N_8355,N_8088,N_7989);
and U8356 (N_8356,N_7842,N_7698);
and U8357 (N_8357,N_7640,N_7935);
nor U8358 (N_8358,N_8106,N_7662);
or U8359 (N_8359,N_7672,N_7696);
or U8360 (N_8360,N_7705,N_7754);
nand U8361 (N_8361,N_7631,N_8056);
nor U8362 (N_8362,N_7586,N_7897);
nor U8363 (N_8363,N_7706,N_8026);
and U8364 (N_8364,N_7805,N_7929);
and U8365 (N_8365,N_8071,N_7560);
or U8366 (N_8366,N_7770,N_7658);
xnor U8367 (N_8367,N_7544,N_8124);
and U8368 (N_8368,N_7518,N_8099);
xnor U8369 (N_8369,N_8005,N_7788);
or U8370 (N_8370,N_8015,N_8033);
and U8371 (N_8371,N_8007,N_7996);
and U8372 (N_8372,N_7933,N_7505);
or U8373 (N_8373,N_7793,N_7600);
xnor U8374 (N_8374,N_8045,N_7822);
nand U8375 (N_8375,N_7964,N_7988);
xor U8376 (N_8376,N_7843,N_7624);
or U8377 (N_8377,N_7723,N_7576);
nand U8378 (N_8378,N_8019,N_7542);
nand U8379 (N_8379,N_7678,N_7844);
and U8380 (N_8380,N_7773,N_7744);
and U8381 (N_8381,N_7956,N_7892);
nand U8382 (N_8382,N_7530,N_7828);
nand U8383 (N_8383,N_7971,N_7529);
or U8384 (N_8384,N_7774,N_8098);
nand U8385 (N_8385,N_7997,N_7567);
nand U8386 (N_8386,N_7979,N_7607);
and U8387 (N_8387,N_7656,N_8039);
xor U8388 (N_8388,N_7649,N_8051);
or U8389 (N_8389,N_7889,N_8085);
xor U8390 (N_8390,N_7990,N_7740);
and U8391 (N_8391,N_7669,N_8080);
xor U8392 (N_8392,N_7987,N_8093);
or U8393 (N_8393,N_7730,N_7888);
nand U8394 (N_8394,N_8044,N_7502);
or U8395 (N_8395,N_7750,N_7636);
xor U8396 (N_8396,N_7755,N_7582);
nand U8397 (N_8397,N_7986,N_7556);
or U8398 (N_8398,N_7877,N_7524);
nor U8399 (N_8399,N_7806,N_7749);
or U8400 (N_8400,N_7572,N_7812);
and U8401 (N_8401,N_8004,N_7563);
nand U8402 (N_8402,N_7856,N_7602);
nor U8403 (N_8403,N_7699,N_7973);
and U8404 (N_8404,N_7511,N_7800);
nor U8405 (N_8405,N_7578,N_7681);
nand U8406 (N_8406,N_8025,N_7799);
and U8407 (N_8407,N_7661,N_7784);
and U8408 (N_8408,N_8034,N_7958);
xor U8409 (N_8409,N_7575,N_8043);
or U8410 (N_8410,N_7590,N_7998);
and U8411 (N_8411,N_7562,N_7717);
xnor U8412 (N_8412,N_7504,N_7786);
nand U8413 (N_8413,N_7879,N_7718);
or U8414 (N_8414,N_8122,N_8058);
and U8415 (N_8415,N_7995,N_7550);
and U8416 (N_8416,N_7647,N_8020);
or U8417 (N_8417,N_7619,N_8121);
and U8418 (N_8418,N_8009,N_7912);
or U8419 (N_8419,N_7659,N_7548);
and U8420 (N_8420,N_8070,N_7525);
nor U8421 (N_8421,N_7555,N_7606);
or U8422 (N_8422,N_7916,N_7654);
or U8423 (N_8423,N_8050,N_7960);
and U8424 (N_8424,N_7641,N_8002);
or U8425 (N_8425,N_7745,N_7728);
or U8426 (N_8426,N_7702,N_7880);
and U8427 (N_8427,N_7726,N_7714);
or U8428 (N_8428,N_7763,N_8104);
xnor U8429 (N_8429,N_7817,N_7537);
or U8430 (N_8430,N_7707,N_7776);
and U8431 (N_8431,N_7655,N_7908);
and U8432 (N_8432,N_7620,N_7512);
and U8433 (N_8433,N_7999,N_7557);
nor U8434 (N_8434,N_7725,N_8023);
or U8435 (N_8435,N_8084,N_8064);
nand U8436 (N_8436,N_7849,N_8091);
and U8437 (N_8437,N_8037,N_7673);
and U8438 (N_8438,N_7800,N_7805);
xnor U8439 (N_8439,N_7575,N_7811);
nand U8440 (N_8440,N_7973,N_7728);
or U8441 (N_8441,N_7521,N_7810);
nand U8442 (N_8442,N_8054,N_7835);
nor U8443 (N_8443,N_7698,N_7516);
nand U8444 (N_8444,N_7831,N_8027);
or U8445 (N_8445,N_8015,N_7960);
nor U8446 (N_8446,N_7576,N_7656);
or U8447 (N_8447,N_7734,N_7586);
nand U8448 (N_8448,N_7783,N_7523);
nand U8449 (N_8449,N_7862,N_8124);
or U8450 (N_8450,N_7678,N_7985);
or U8451 (N_8451,N_8093,N_7591);
nand U8452 (N_8452,N_7517,N_7634);
and U8453 (N_8453,N_7619,N_7560);
nand U8454 (N_8454,N_7986,N_8050);
and U8455 (N_8455,N_7976,N_7807);
or U8456 (N_8456,N_7803,N_7556);
or U8457 (N_8457,N_8080,N_7956);
nor U8458 (N_8458,N_7991,N_7540);
nand U8459 (N_8459,N_8012,N_7514);
nand U8460 (N_8460,N_7771,N_7552);
nor U8461 (N_8461,N_7861,N_7905);
nor U8462 (N_8462,N_8102,N_7598);
xor U8463 (N_8463,N_7799,N_8124);
nand U8464 (N_8464,N_8035,N_7890);
and U8465 (N_8465,N_8067,N_7940);
and U8466 (N_8466,N_7551,N_7869);
nor U8467 (N_8467,N_7745,N_7977);
nor U8468 (N_8468,N_7950,N_7523);
nand U8469 (N_8469,N_7565,N_7814);
nor U8470 (N_8470,N_7742,N_8071);
nor U8471 (N_8471,N_7964,N_8093);
and U8472 (N_8472,N_8116,N_7967);
xor U8473 (N_8473,N_7547,N_7587);
and U8474 (N_8474,N_7601,N_7884);
nor U8475 (N_8475,N_7735,N_7782);
nor U8476 (N_8476,N_7980,N_7526);
or U8477 (N_8477,N_7683,N_7603);
and U8478 (N_8478,N_7701,N_7863);
and U8479 (N_8479,N_8049,N_7985);
nor U8480 (N_8480,N_7857,N_7689);
and U8481 (N_8481,N_7792,N_7878);
nor U8482 (N_8482,N_8074,N_7827);
xor U8483 (N_8483,N_7643,N_8091);
xnor U8484 (N_8484,N_7819,N_7902);
nor U8485 (N_8485,N_8047,N_7800);
or U8486 (N_8486,N_7985,N_8102);
xnor U8487 (N_8487,N_7927,N_7558);
and U8488 (N_8488,N_7711,N_7607);
nor U8489 (N_8489,N_7529,N_7819);
or U8490 (N_8490,N_7798,N_8023);
nand U8491 (N_8491,N_7689,N_7794);
or U8492 (N_8492,N_7797,N_7718);
nor U8493 (N_8493,N_7595,N_8046);
or U8494 (N_8494,N_7540,N_7712);
nor U8495 (N_8495,N_7840,N_7785);
and U8496 (N_8496,N_8008,N_7519);
nand U8497 (N_8497,N_7722,N_8063);
or U8498 (N_8498,N_7519,N_7663);
or U8499 (N_8499,N_7951,N_7812);
and U8500 (N_8500,N_7952,N_8067);
nor U8501 (N_8501,N_7765,N_8016);
nor U8502 (N_8502,N_7934,N_7962);
and U8503 (N_8503,N_8105,N_7740);
and U8504 (N_8504,N_7914,N_8117);
and U8505 (N_8505,N_7872,N_7550);
or U8506 (N_8506,N_7771,N_8040);
nor U8507 (N_8507,N_7583,N_7661);
nor U8508 (N_8508,N_7802,N_8087);
nor U8509 (N_8509,N_8048,N_7995);
nand U8510 (N_8510,N_8028,N_7715);
or U8511 (N_8511,N_7624,N_7618);
nor U8512 (N_8512,N_7951,N_7723);
nor U8513 (N_8513,N_7508,N_8089);
nand U8514 (N_8514,N_7559,N_7820);
and U8515 (N_8515,N_7901,N_7991);
xnor U8516 (N_8516,N_8060,N_7676);
nor U8517 (N_8517,N_8047,N_7987);
or U8518 (N_8518,N_8050,N_7669);
xor U8519 (N_8519,N_8023,N_8061);
or U8520 (N_8520,N_7905,N_8122);
nand U8521 (N_8521,N_7616,N_7980);
xor U8522 (N_8522,N_7974,N_7917);
nor U8523 (N_8523,N_7587,N_7556);
nand U8524 (N_8524,N_8008,N_7609);
xnor U8525 (N_8525,N_7745,N_7549);
or U8526 (N_8526,N_8107,N_7527);
nor U8527 (N_8527,N_8044,N_8009);
xnor U8528 (N_8528,N_7953,N_7904);
nand U8529 (N_8529,N_8013,N_7615);
and U8530 (N_8530,N_7919,N_7944);
nor U8531 (N_8531,N_7717,N_7894);
nor U8532 (N_8532,N_7592,N_8118);
nor U8533 (N_8533,N_7876,N_7726);
nand U8534 (N_8534,N_7675,N_7848);
and U8535 (N_8535,N_7802,N_7726);
nand U8536 (N_8536,N_7987,N_7997);
or U8537 (N_8537,N_7524,N_7799);
nor U8538 (N_8538,N_7918,N_7904);
nor U8539 (N_8539,N_8026,N_8080);
nor U8540 (N_8540,N_7556,N_7877);
or U8541 (N_8541,N_7794,N_7795);
or U8542 (N_8542,N_7920,N_7860);
and U8543 (N_8543,N_7828,N_7808);
nand U8544 (N_8544,N_7735,N_8019);
nor U8545 (N_8545,N_7578,N_8120);
nand U8546 (N_8546,N_7823,N_8064);
nand U8547 (N_8547,N_7800,N_7975);
or U8548 (N_8548,N_7623,N_7550);
nand U8549 (N_8549,N_7823,N_7659);
nor U8550 (N_8550,N_7887,N_8053);
nand U8551 (N_8551,N_7886,N_8076);
and U8552 (N_8552,N_7660,N_7754);
nor U8553 (N_8553,N_7720,N_7673);
and U8554 (N_8554,N_7717,N_8117);
or U8555 (N_8555,N_7915,N_7508);
or U8556 (N_8556,N_7693,N_7685);
xnor U8557 (N_8557,N_7711,N_7971);
and U8558 (N_8558,N_7584,N_8003);
nor U8559 (N_8559,N_7554,N_8080);
or U8560 (N_8560,N_7913,N_7901);
or U8561 (N_8561,N_8065,N_8068);
nand U8562 (N_8562,N_7938,N_7911);
and U8563 (N_8563,N_7596,N_7577);
nor U8564 (N_8564,N_7527,N_7813);
nand U8565 (N_8565,N_7560,N_7537);
or U8566 (N_8566,N_7841,N_7767);
or U8567 (N_8567,N_7821,N_7559);
nor U8568 (N_8568,N_7620,N_8039);
nand U8569 (N_8569,N_7795,N_8079);
nand U8570 (N_8570,N_7564,N_7820);
nor U8571 (N_8571,N_8089,N_7735);
and U8572 (N_8572,N_8069,N_7745);
or U8573 (N_8573,N_7987,N_7519);
or U8574 (N_8574,N_7587,N_7768);
xnor U8575 (N_8575,N_8062,N_7822);
nor U8576 (N_8576,N_7984,N_7822);
nor U8577 (N_8577,N_7603,N_8053);
and U8578 (N_8578,N_7853,N_7574);
and U8579 (N_8579,N_7974,N_7964);
or U8580 (N_8580,N_8054,N_7710);
and U8581 (N_8581,N_8048,N_7502);
and U8582 (N_8582,N_7577,N_7552);
nand U8583 (N_8583,N_7556,N_7931);
and U8584 (N_8584,N_7583,N_7516);
xnor U8585 (N_8585,N_7629,N_7680);
nand U8586 (N_8586,N_7979,N_8021);
nor U8587 (N_8587,N_7801,N_8049);
and U8588 (N_8588,N_7646,N_7795);
xor U8589 (N_8589,N_7667,N_8048);
nand U8590 (N_8590,N_7954,N_7825);
nand U8591 (N_8591,N_8073,N_7601);
and U8592 (N_8592,N_7899,N_7677);
or U8593 (N_8593,N_7761,N_7560);
nand U8594 (N_8594,N_7693,N_7675);
nor U8595 (N_8595,N_7623,N_7520);
nand U8596 (N_8596,N_8046,N_7587);
or U8597 (N_8597,N_7981,N_7558);
or U8598 (N_8598,N_7970,N_8068);
nor U8599 (N_8599,N_7753,N_7706);
or U8600 (N_8600,N_7829,N_8035);
or U8601 (N_8601,N_7947,N_7573);
or U8602 (N_8602,N_7933,N_7694);
or U8603 (N_8603,N_7933,N_7908);
and U8604 (N_8604,N_7591,N_7635);
nor U8605 (N_8605,N_7983,N_7879);
and U8606 (N_8606,N_7881,N_7618);
and U8607 (N_8607,N_7953,N_7609);
and U8608 (N_8608,N_7947,N_7830);
nand U8609 (N_8609,N_8050,N_7538);
nor U8610 (N_8610,N_7854,N_7994);
nor U8611 (N_8611,N_7514,N_7596);
and U8612 (N_8612,N_7725,N_7613);
or U8613 (N_8613,N_7563,N_7719);
or U8614 (N_8614,N_7862,N_7566);
nand U8615 (N_8615,N_7595,N_7839);
nand U8616 (N_8616,N_7827,N_8035);
nand U8617 (N_8617,N_7816,N_7996);
and U8618 (N_8618,N_7748,N_8072);
or U8619 (N_8619,N_8111,N_7699);
nand U8620 (N_8620,N_8062,N_7716);
nand U8621 (N_8621,N_7734,N_8056);
xor U8622 (N_8622,N_7587,N_7988);
or U8623 (N_8623,N_7688,N_7929);
nand U8624 (N_8624,N_7554,N_7915);
nor U8625 (N_8625,N_7716,N_7719);
xor U8626 (N_8626,N_8065,N_7787);
or U8627 (N_8627,N_7506,N_7616);
xnor U8628 (N_8628,N_7696,N_7823);
nor U8629 (N_8629,N_7717,N_7502);
nor U8630 (N_8630,N_7801,N_8009);
nor U8631 (N_8631,N_7885,N_7598);
nand U8632 (N_8632,N_8098,N_7864);
nand U8633 (N_8633,N_7801,N_7752);
and U8634 (N_8634,N_7990,N_7889);
and U8635 (N_8635,N_7934,N_7930);
nand U8636 (N_8636,N_7877,N_7640);
or U8637 (N_8637,N_7695,N_7584);
nand U8638 (N_8638,N_7800,N_7763);
or U8639 (N_8639,N_7866,N_7895);
and U8640 (N_8640,N_7529,N_7951);
and U8641 (N_8641,N_7587,N_8026);
or U8642 (N_8642,N_8087,N_8119);
nor U8643 (N_8643,N_7986,N_7687);
and U8644 (N_8644,N_7729,N_7714);
nand U8645 (N_8645,N_7559,N_8098);
or U8646 (N_8646,N_7758,N_8105);
nand U8647 (N_8647,N_7892,N_7584);
nand U8648 (N_8648,N_8099,N_7867);
nand U8649 (N_8649,N_8043,N_7590);
nor U8650 (N_8650,N_7503,N_7575);
nor U8651 (N_8651,N_7664,N_7619);
or U8652 (N_8652,N_8100,N_7937);
xor U8653 (N_8653,N_7766,N_7870);
nor U8654 (N_8654,N_7704,N_8046);
nand U8655 (N_8655,N_8005,N_7934);
nand U8656 (N_8656,N_8081,N_7586);
nand U8657 (N_8657,N_7771,N_7512);
nand U8658 (N_8658,N_7688,N_8097);
nor U8659 (N_8659,N_7636,N_7729);
or U8660 (N_8660,N_7988,N_7978);
or U8661 (N_8661,N_7745,N_7691);
xnor U8662 (N_8662,N_8041,N_7751);
xor U8663 (N_8663,N_7932,N_7653);
nand U8664 (N_8664,N_7718,N_7769);
nor U8665 (N_8665,N_7554,N_7566);
nor U8666 (N_8666,N_7857,N_7745);
nor U8667 (N_8667,N_7793,N_7722);
nor U8668 (N_8668,N_7802,N_8073);
xor U8669 (N_8669,N_7903,N_7945);
or U8670 (N_8670,N_7757,N_7641);
or U8671 (N_8671,N_7896,N_8110);
or U8672 (N_8672,N_7530,N_7896);
nor U8673 (N_8673,N_8056,N_7942);
xnor U8674 (N_8674,N_7807,N_8020);
nor U8675 (N_8675,N_7653,N_7604);
nor U8676 (N_8676,N_7910,N_7840);
nor U8677 (N_8677,N_7953,N_8097);
and U8678 (N_8678,N_7839,N_7830);
or U8679 (N_8679,N_7640,N_7772);
or U8680 (N_8680,N_7555,N_8111);
nor U8681 (N_8681,N_7955,N_8022);
nand U8682 (N_8682,N_7914,N_7636);
nand U8683 (N_8683,N_7953,N_7922);
nand U8684 (N_8684,N_7611,N_7935);
and U8685 (N_8685,N_7502,N_7740);
and U8686 (N_8686,N_7768,N_7930);
nand U8687 (N_8687,N_7959,N_7658);
or U8688 (N_8688,N_7664,N_7504);
nor U8689 (N_8689,N_7727,N_7550);
and U8690 (N_8690,N_7621,N_7777);
nand U8691 (N_8691,N_7790,N_7718);
nand U8692 (N_8692,N_7593,N_7917);
nand U8693 (N_8693,N_7634,N_7584);
nand U8694 (N_8694,N_7519,N_7532);
or U8695 (N_8695,N_7710,N_7895);
or U8696 (N_8696,N_7592,N_7950);
nand U8697 (N_8697,N_8111,N_7553);
nor U8698 (N_8698,N_7810,N_7790);
or U8699 (N_8699,N_7837,N_7968);
nand U8700 (N_8700,N_7654,N_7848);
and U8701 (N_8701,N_7674,N_7675);
nand U8702 (N_8702,N_7546,N_7722);
or U8703 (N_8703,N_7959,N_7750);
and U8704 (N_8704,N_7807,N_7796);
and U8705 (N_8705,N_7570,N_7541);
and U8706 (N_8706,N_8000,N_7964);
and U8707 (N_8707,N_7977,N_7786);
and U8708 (N_8708,N_7687,N_7648);
nor U8709 (N_8709,N_7829,N_7799);
or U8710 (N_8710,N_7849,N_7864);
nand U8711 (N_8711,N_7807,N_7648);
or U8712 (N_8712,N_8103,N_7717);
nand U8713 (N_8713,N_7759,N_8088);
xnor U8714 (N_8714,N_8011,N_7508);
and U8715 (N_8715,N_8080,N_8120);
and U8716 (N_8716,N_7995,N_8033);
or U8717 (N_8717,N_7508,N_7854);
nor U8718 (N_8718,N_7775,N_7689);
nand U8719 (N_8719,N_7542,N_7850);
nor U8720 (N_8720,N_7853,N_7514);
nand U8721 (N_8721,N_7775,N_8110);
and U8722 (N_8722,N_7918,N_7857);
xnor U8723 (N_8723,N_7900,N_7880);
nor U8724 (N_8724,N_7527,N_7958);
nor U8725 (N_8725,N_7578,N_7594);
xor U8726 (N_8726,N_7817,N_7856);
or U8727 (N_8727,N_8084,N_7986);
and U8728 (N_8728,N_8113,N_7920);
nor U8729 (N_8729,N_7664,N_8053);
nand U8730 (N_8730,N_8031,N_7619);
or U8731 (N_8731,N_7563,N_7641);
nand U8732 (N_8732,N_7626,N_7707);
xnor U8733 (N_8733,N_7789,N_7627);
and U8734 (N_8734,N_8016,N_7745);
nor U8735 (N_8735,N_7597,N_7680);
or U8736 (N_8736,N_7612,N_7718);
and U8737 (N_8737,N_7642,N_7957);
xor U8738 (N_8738,N_7627,N_7994);
or U8739 (N_8739,N_8103,N_7762);
nand U8740 (N_8740,N_7620,N_8083);
nand U8741 (N_8741,N_7802,N_7799);
nand U8742 (N_8742,N_8044,N_7924);
nand U8743 (N_8743,N_7819,N_7513);
nand U8744 (N_8744,N_7887,N_7759);
nor U8745 (N_8745,N_7727,N_7547);
nor U8746 (N_8746,N_8052,N_7591);
nor U8747 (N_8747,N_7588,N_7628);
and U8748 (N_8748,N_7654,N_7751);
or U8749 (N_8749,N_7636,N_7569);
nor U8750 (N_8750,N_8463,N_8514);
xnor U8751 (N_8751,N_8359,N_8737);
and U8752 (N_8752,N_8268,N_8392);
or U8753 (N_8753,N_8493,N_8420);
nor U8754 (N_8754,N_8425,N_8656);
nor U8755 (N_8755,N_8485,N_8572);
xor U8756 (N_8756,N_8381,N_8500);
nand U8757 (N_8757,N_8202,N_8263);
nor U8758 (N_8758,N_8167,N_8154);
nor U8759 (N_8759,N_8378,N_8642);
nand U8760 (N_8760,N_8497,N_8242);
or U8761 (N_8761,N_8413,N_8264);
nand U8762 (N_8762,N_8362,N_8182);
nor U8763 (N_8763,N_8716,N_8593);
nor U8764 (N_8764,N_8467,N_8351);
nor U8765 (N_8765,N_8501,N_8513);
nand U8766 (N_8766,N_8221,N_8416);
nand U8767 (N_8767,N_8130,N_8733);
xor U8768 (N_8768,N_8406,N_8335);
nand U8769 (N_8769,N_8295,N_8371);
and U8770 (N_8770,N_8526,N_8709);
nand U8771 (N_8771,N_8645,N_8449);
nor U8772 (N_8772,N_8403,N_8507);
or U8773 (N_8773,N_8715,N_8739);
nand U8774 (N_8774,N_8290,N_8292);
nand U8775 (N_8775,N_8330,N_8627);
or U8776 (N_8776,N_8260,N_8749);
and U8777 (N_8777,N_8603,N_8294);
xor U8778 (N_8778,N_8168,N_8414);
or U8779 (N_8779,N_8320,N_8280);
nor U8780 (N_8780,N_8655,N_8470);
nor U8781 (N_8781,N_8651,N_8411);
xor U8782 (N_8782,N_8325,N_8271);
or U8783 (N_8783,N_8602,N_8194);
or U8784 (N_8784,N_8172,N_8691);
or U8785 (N_8785,N_8701,N_8375);
or U8786 (N_8786,N_8592,N_8402);
nor U8787 (N_8787,N_8744,N_8620);
or U8788 (N_8788,N_8678,N_8451);
xnor U8789 (N_8789,N_8486,N_8708);
and U8790 (N_8790,N_8207,N_8309);
or U8791 (N_8791,N_8609,N_8660);
nand U8792 (N_8792,N_8265,N_8272);
nand U8793 (N_8793,N_8253,N_8353);
and U8794 (N_8794,N_8519,N_8647);
or U8795 (N_8795,N_8509,N_8588);
nor U8796 (N_8796,N_8719,N_8595);
nand U8797 (N_8797,N_8574,N_8350);
or U8798 (N_8798,N_8631,N_8312);
or U8799 (N_8799,N_8633,N_8545);
nor U8800 (N_8800,N_8596,N_8316);
or U8801 (N_8801,N_8398,N_8148);
or U8802 (N_8802,N_8462,N_8517);
or U8803 (N_8803,N_8480,N_8275);
nand U8804 (N_8804,N_8146,N_8421);
xnor U8805 (N_8805,N_8210,N_8319);
nor U8806 (N_8806,N_8198,N_8313);
or U8807 (N_8807,N_8630,N_8686);
nand U8808 (N_8808,N_8576,N_8504);
nor U8809 (N_8809,N_8632,N_8689);
nor U8810 (N_8810,N_8615,N_8674);
nand U8811 (N_8811,N_8446,N_8156);
nand U8812 (N_8812,N_8555,N_8441);
nand U8813 (N_8813,N_8274,N_8508);
nor U8814 (N_8814,N_8569,N_8372);
and U8815 (N_8815,N_8166,N_8525);
nand U8816 (N_8816,N_8583,N_8579);
or U8817 (N_8817,N_8426,N_8190);
and U8818 (N_8818,N_8277,N_8464);
nor U8819 (N_8819,N_8561,N_8183);
nand U8820 (N_8820,N_8684,N_8358);
or U8821 (N_8821,N_8237,N_8394);
and U8822 (N_8822,N_8582,N_8531);
or U8823 (N_8823,N_8400,N_8624);
xor U8824 (N_8824,N_8374,N_8456);
nor U8825 (N_8825,N_8738,N_8562);
and U8826 (N_8826,N_8422,N_8713);
xor U8827 (N_8827,N_8306,N_8393);
nand U8828 (N_8828,N_8566,N_8554);
and U8829 (N_8829,N_8439,N_8613);
xnor U8830 (N_8830,N_8494,N_8506);
nand U8831 (N_8831,N_8254,N_8160);
nor U8832 (N_8832,N_8587,N_8687);
or U8833 (N_8833,N_8502,N_8363);
nor U8834 (N_8834,N_8721,N_8412);
and U8835 (N_8835,N_8440,N_8409);
nor U8836 (N_8836,N_8401,N_8543);
and U8837 (N_8837,N_8257,N_8235);
nand U8838 (N_8838,N_8189,N_8226);
nand U8839 (N_8839,N_8356,N_8735);
or U8840 (N_8840,N_8720,N_8157);
nor U8841 (N_8841,N_8225,N_8734);
nand U8842 (N_8842,N_8155,N_8153);
nand U8843 (N_8843,N_8339,N_8246);
or U8844 (N_8844,N_8340,N_8193);
or U8845 (N_8845,N_8455,N_8380);
and U8846 (N_8846,N_8307,N_8383);
nor U8847 (N_8847,N_8216,N_8315);
or U8848 (N_8848,N_8410,N_8331);
or U8849 (N_8849,N_8186,N_8327);
nand U8850 (N_8850,N_8149,N_8418);
nand U8851 (N_8851,N_8657,N_8717);
nand U8852 (N_8852,N_8430,N_8597);
or U8853 (N_8853,N_8673,N_8283);
nand U8854 (N_8854,N_8250,N_8606);
xnor U8855 (N_8855,N_8432,N_8136);
nor U8856 (N_8856,N_8305,N_8177);
and U8857 (N_8857,N_8334,N_8668);
xor U8858 (N_8858,N_8669,N_8191);
nand U8859 (N_8859,N_8725,N_8236);
xnor U8860 (N_8860,N_8288,N_8165);
and U8861 (N_8861,N_8707,N_8693);
nor U8862 (N_8862,N_8259,N_8389);
nand U8863 (N_8863,N_8591,N_8747);
nand U8864 (N_8864,N_8466,N_8397);
and U8865 (N_8865,N_8293,N_8296);
and U8866 (N_8866,N_8220,N_8147);
nor U8867 (N_8867,N_8352,N_8141);
or U8868 (N_8868,N_8289,N_8698);
nor U8869 (N_8869,N_8303,N_8458);
and U8870 (N_8870,N_8249,N_8213);
nand U8871 (N_8871,N_8454,N_8310);
and U8872 (N_8872,N_8512,N_8524);
and U8873 (N_8873,N_8518,N_8269);
nand U8874 (N_8874,N_8457,N_8623);
or U8875 (N_8875,N_8344,N_8304);
or U8876 (N_8876,N_8557,N_8131);
nand U8877 (N_8877,N_8170,N_8675);
nor U8878 (N_8878,N_8585,N_8437);
nand U8879 (N_8879,N_8227,N_8533);
nand U8880 (N_8880,N_8270,N_8499);
or U8881 (N_8881,N_8492,N_8178);
nand U8882 (N_8882,N_8360,N_8276);
nor U8883 (N_8883,N_8142,N_8710);
or U8884 (N_8884,N_8560,N_8450);
nor U8885 (N_8885,N_8740,N_8549);
nand U8886 (N_8886,N_8284,N_8646);
or U8887 (N_8887,N_8228,N_8590);
nor U8888 (N_8888,N_8217,N_8677);
nand U8889 (N_8889,N_8143,N_8407);
nand U8890 (N_8890,N_8644,N_8471);
and U8891 (N_8891,N_8681,N_8598);
and U8892 (N_8892,N_8638,N_8152);
or U8893 (N_8893,N_8702,N_8298);
nor U8894 (N_8894,N_8245,N_8722);
nand U8895 (N_8895,N_8438,N_8247);
and U8896 (N_8896,N_8629,N_8662);
nor U8897 (N_8897,N_8619,N_8212);
nand U8898 (N_8898,N_8215,N_8175);
and U8899 (N_8899,N_8337,N_8195);
nor U8900 (N_8900,N_8688,N_8343);
nor U8901 (N_8901,N_8666,N_8251);
or U8902 (N_8902,N_8333,N_8329);
and U8903 (N_8903,N_8164,N_8643);
nor U8904 (N_8904,N_8435,N_8390);
or U8905 (N_8905,N_8649,N_8553);
nand U8906 (N_8906,N_8511,N_8634);
nor U8907 (N_8907,N_8529,N_8382);
nand U8908 (N_8908,N_8726,N_8234);
nor U8909 (N_8909,N_8162,N_8445);
nor U8910 (N_8910,N_8498,N_8433);
and U8911 (N_8911,N_8637,N_8302);
nor U8912 (N_8912,N_8266,N_8127);
and U8913 (N_8913,N_8711,N_8523);
or U8914 (N_8914,N_8336,N_8324);
or U8915 (N_8915,N_8653,N_8604);
or U8916 (N_8916,N_8682,N_8408);
and U8917 (N_8917,N_8540,N_8125);
xor U8918 (N_8918,N_8161,N_8460);
nand U8919 (N_8919,N_8484,N_8599);
or U8920 (N_8920,N_8448,N_8184);
nand U8921 (N_8921,N_8159,N_8652);
and U8922 (N_8922,N_8536,N_8308);
nor U8923 (N_8923,N_8469,N_8395);
nand U8924 (N_8924,N_8522,N_8559);
nand U8925 (N_8925,N_8636,N_8238);
nand U8926 (N_8926,N_8661,N_8200);
nor U8927 (N_8927,N_8654,N_8368);
xnor U8928 (N_8928,N_8206,N_8384);
nor U8929 (N_8929,N_8145,N_8328);
nand U8930 (N_8930,N_8743,N_8472);
nor U8931 (N_8931,N_8584,N_8405);
nor U8932 (N_8932,N_8612,N_8132);
and U8933 (N_8933,N_8601,N_8683);
nand U8934 (N_8934,N_8424,N_8199);
and U8935 (N_8935,N_8690,N_8544);
nor U8936 (N_8936,N_8580,N_8704);
nor U8937 (N_8937,N_8126,N_8427);
xnor U8938 (N_8938,N_8481,N_8391);
nand U8939 (N_8939,N_8151,N_8388);
and U8940 (N_8940,N_8137,N_8219);
nand U8941 (N_8941,N_8347,N_8285);
nor U8942 (N_8942,N_8729,N_8510);
and U8943 (N_8943,N_8176,N_8317);
nor U8944 (N_8944,N_8273,N_8703);
nand U8945 (N_8945,N_8685,N_8474);
nand U8946 (N_8946,N_8699,N_8291);
nand U8947 (N_8947,N_8479,N_8173);
or U8948 (N_8948,N_8639,N_8279);
nand U8949 (N_8949,N_8745,N_8692);
nand U8950 (N_8950,N_8341,N_8150);
nor U8951 (N_8951,N_8248,N_8434);
and U8952 (N_8952,N_8214,N_8581);
xor U8953 (N_8953,N_8244,N_8267);
xor U8954 (N_8954,N_8443,N_8261);
and U8955 (N_8955,N_8730,N_8346);
nand U8956 (N_8956,N_8558,N_8197);
xor U8957 (N_8957,N_8223,N_8622);
nand U8958 (N_8958,N_8565,N_8700);
nand U8959 (N_8959,N_8551,N_8299);
and U8960 (N_8960,N_8366,N_8748);
and U8961 (N_8961,N_8680,N_8354);
nand U8962 (N_8962,N_8192,N_8431);
and U8963 (N_8963,N_8618,N_8663);
xnor U8964 (N_8964,N_8240,N_8256);
nor U8965 (N_8965,N_8659,N_8286);
xor U8966 (N_8966,N_8625,N_8530);
and U8967 (N_8967,N_8736,N_8187);
nor U8968 (N_8968,N_8428,N_8376);
or U8969 (N_8969,N_8300,N_8664);
and U8970 (N_8970,N_8365,N_8600);
nand U8971 (N_8971,N_8527,N_8342);
and U8972 (N_8972,N_8594,N_8746);
and U8973 (N_8973,N_8573,N_8496);
or U8974 (N_8974,N_8488,N_8239);
and U8975 (N_8975,N_8586,N_8321);
nand U8976 (N_8976,N_8505,N_8231);
nand U8977 (N_8977,N_8490,N_8658);
nand U8978 (N_8978,N_8714,N_8548);
nor U8979 (N_8979,N_8728,N_8255);
nor U8980 (N_8980,N_8552,N_8465);
nor U8981 (N_8981,N_8287,N_8282);
xnor U8982 (N_8982,N_8205,N_8396);
nor U8983 (N_8983,N_8589,N_8318);
or U8984 (N_8984,N_8196,N_8671);
nand U8985 (N_8985,N_8230,N_8539);
nand U8986 (N_8986,N_8163,N_8571);
and U8987 (N_8987,N_8211,N_8741);
nand U8988 (N_8988,N_8224,N_8635);
nor U8989 (N_8989,N_8209,N_8535);
xor U8990 (N_8990,N_8578,N_8222);
xor U8991 (N_8991,N_8694,N_8563);
nor U8992 (N_8992,N_8323,N_8444);
xnor U8993 (N_8993,N_8621,N_8537);
nor U8994 (N_8994,N_8181,N_8487);
or U8995 (N_8995,N_8705,N_8326);
and U8996 (N_8996,N_8369,N_8532);
or U8997 (N_8997,N_8477,N_8489);
nand U8998 (N_8998,N_8361,N_8516);
and U8999 (N_8999,N_8607,N_8570);
nand U9000 (N_9000,N_8575,N_8528);
and U9001 (N_9001,N_8218,N_8476);
or U9002 (N_9002,N_8387,N_8568);
nor U9003 (N_9003,N_8731,N_8712);
xor U9004 (N_9004,N_8468,N_8605);
or U9005 (N_9005,N_8732,N_8201);
and U9006 (N_9006,N_8676,N_8232);
nand U9007 (N_9007,N_8696,N_8417);
nand U9008 (N_9008,N_8648,N_8447);
xnor U9009 (N_9009,N_8567,N_8442);
xor U9010 (N_9010,N_8577,N_8550);
nor U9011 (N_9011,N_8534,N_8399);
or U9012 (N_9012,N_8616,N_8461);
xnor U9013 (N_9013,N_8278,N_8129);
or U9014 (N_9014,N_8204,N_8641);
xnor U9015 (N_9015,N_8241,N_8348);
nor U9016 (N_9016,N_8338,N_8144);
and U9017 (N_9017,N_8723,N_8262);
and U9018 (N_9018,N_8281,N_8203);
and U9019 (N_9019,N_8520,N_8650);
nand U9020 (N_9020,N_8495,N_8301);
nor U9021 (N_9021,N_8640,N_8139);
and U9022 (N_9022,N_8742,N_8706);
xor U9023 (N_9023,N_8419,N_8174);
nor U9024 (N_9024,N_8429,N_8373);
nand U9025 (N_9025,N_8718,N_8617);
or U9026 (N_9026,N_8138,N_8459);
and U9027 (N_9027,N_8697,N_8473);
xor U9028 (N_9028,N_8357,N_8311);
nor U9029 (N_9029,N_8252,N_8672);
or U9030 (N_9030,N_8370,N_8503);
and U9031 (N_9031,N_8332,N_8491);
nor U9032 (N_9032,N_8628,N_8322);
or U9033 (N_9033,N_8243,N_8564);
nor U9034 (N_9034,N_8345,N_8297);
nand U9035 (N_9035,N_8436,N_8665);
nand U9036 (N_9036,N_8478,N_8188);
nand U9037 (N_9037,N_8233,N_8611);
nand U9038 (N_9038,N_8546,N_8314);
nor U9039 (N_9039,N_8169,N_8541);
nand U9040 (N_9040,N_8208,N_8133);
nand U9041 (N_9041,N_8158,N_8483);
nor U9042 (N_9042,N_8364,N_8667);
and U9043 (N_9043,N_8610,N_8135);
nand U9044 (N_9044,N_8185,N_8179);
nor U9045 (N_9045,N_8349,N_8515);
and U9046 (N_9046,N_8377,N_8452);
and U9047 (N_9047,N_8180,N_8171);
and U9048 (N_9048,N_8626,N_8453);
nor U9049 (N_9049,N_8614,N_8415);
or U9050 (N_9050,N_8556,N_8386);
nor U9051 (N_9051,N_8423,N_8538);
and U9052 (N_9052,N_8258,N_8128);
or U9053 (N_9053,N_8379,N_8355);
and U9054 (N_9054,N_8140,N_8727);
nor U9055 (N_9055,N_8679,N_8695);
nor U9056 (N_9056,N_8404,N_8385);
or U9057 (N_9057,N_8482,N_8475);
nor U9058 (N_9058,N_8724,N_8521);
or U9059 (N_9059,N_8542,N_8367);
and U9060 (N_9060,N_8670,N_8134);
xnor U9061 (N_9061,N_8608,N_8547);
or U9062 (N_9062,N_8229,N_8675);
nand U9063 (N_9063,N_8371,N_8550);
and U9064 (N_9064,N_8340,N_8406);
nor U9065 (N_9065,N_8658,N_8586);
and U9066 (N_9066,N_8399,N_8598);
or U9067 (N_9067,N_8359,N_8720);
nand U9068 (N_9068,N_8364,N_8648);
and U9069 (N_9069,N_8354,N_8723);
nor U9070 (N_9070,N_8639,N_8206);
or U9071 (N_9071,N_8675,N_8705);
and U9072 (N_9072,N_8279,N_8126);
and U9073 (N_9073,N_8490,N_8534);
nand U9074 (N_9074,N_8296,N_8339);
xor U9075 (N_9075,N_8567,N_8356);
and U9076 (N_9076,N_8487,N_8217);
nor U9077 (N_9077,N_8431,N_8416);
nor U9078 (N_9078,N_8454,N_8597);
or U9079 (N_9079,N_8155,N_8633);
nor U9080 (N_9080,N_8520,N_8189);
or U9081 (N_9081,N_8502,N_8480);
nor U9082 (N_9082,N_8241,N_8687);
xor U9083 (N_9083,N_8717,N_8297);
and U9084 (N_9084,N_8544,N_8163);
nor U9085 (N_9085,N_8132,N_8554);
and U9086 (N_9086,N_8298,N_8276);
or U9087 (N_9087,N_8667,N_8620);
nand U9088 (N_9088,N_8466,N_8604);
xor U9089 (N_9089,N_8206,N_8386);
xnor U9090 (N_9090,N_8398,N_8596);
or U9091 (N_9091,N_8300,N_8736);
nand U9092 (N_9092,N_8276,N_8323);
or U9093 (N_9093,N_8265,N_8615);
and U9094 (N_9094,N_8453,N_8458);
nor U9095 (N_9095,N_8467,N_8164);
or U9096 (N_9096,N_8233,N_8247);
or U9097 (N_9097,N_8733,N_8162);
or U9098 (N_9098,N_8246,N_8586);
xnor U9099 (N_9099,N_8200,N_8352);
or U9100 (N_9100,N_8682,N_8380);
nand U9101 (N_9101,N_8395,N_8663);
nor U9102 (N_9102,N_8270,N_8374);
nor U9103 (N_9103,N_8241,N_8165);
nor U9104 (N_9104,N_8474,N_8281);
nor U9105 (N_9105,N_8591,N_8184);
nor U9106 (N_9106,N_8296,N_8522);
and U9107 (N_9107,N_8489,N_8541);
or U9108 (N_9108,N_8337,N_8712);
and U9109 (N_9109,N_8507,N_8434);
and U9110 (N_9110,N_8580,N_8699);
nor U9111 (N_9111,N_8153,N_8180);
nand U9112 (N_9112,N_8667,N_8313);
nand U9113 (N_9113,N_8181,N_8715);
nand U9114 (N_9114,N_8653,N_8739);
xor U9115 (N_9115,N_8710,N_8464);
nand U9116 (N_9116,N_8189,N_8303);
nor U9117 (N_9117,N_8602,N_8337);
or U9118 (N_9118,N_8130,N_8336);
nor U9119 (N_9119,N_8565,N_8488);
nand U9120 (N_9120,N_8621,N_8339);
nor U9121 (N_9121,N_8477,N_8466);
and U9122 (N_9122,N_8312,N_8353);
or U9123 (N_9123,N_8495,N_8749);
and U9124 (N_9124,N_8709,N_8282);
and U9125 (N_9125,N_8262,N_8565);
or U9126 (N_9126,N_8347,N_8129);
or U9127 (N_9127,N_8466,N_8388);
nor U9128 (N_9128,N_8412,N_8275);
and U9129 (N_9129,N_8140,N_8596);
xor U9130 (N_9130,N_8363,N_8241);
or U9131 (N_9131,N_8499,N_8369);
nor U9132 (N_9132,N_8678,N_8607);
and U9133 (N_9133,N_8426,N_8685);
and U9134 (N_9134,N_8131,N_8672);
nor U9135 (N_9135,N_8456,N_8270);
and U9136 (N_9136,N_8423,N_8589);
nor U9137 (N_9137,N_8224,N_8599);
xor U9138 (N_9138,N_8631,N_8726);
nor U9139 (N_9139,N_8552,N_8656);
nor U9140 (N_9140,N_8483,N_8650);
and U9141 (N_9141,N_8407,N_8267);
and U9142 (N_9142,N_8220,N_8505);
nor U9143 (N_9143,N_8164,N_8474);
nor U9144 (N_9144,N_8489,N_8665);
or U9145 (N_9145,N_8229,N_8174);
and U9146 (N_9146,N_8624,N_8534);
nand U9147 (N_9147,N_8278,N_8713);
and U9148 (N_9148,N_8280,N_8304);
and U9149 (N_9149,N_8248,N_8713);
nand U9150 (N_9150,N_8451,N_8541);
and U9151 (N_9151,N_8426,N_8653);
and U9152 (N_9152,N_8698,N_8527);
nand U9153 (N_9153,N_8138,N_8481);
nand U9154 (N_9154,N_8606,N_8580);
and U9155 (N_9155,N_8725,N_8516);
xnor U9156 (N_9156,N_8295,N_8293);
xor U9157 (N_9157,N_8244,N_8381);
or U9158 (N_9158,N_8562,N_8282);
or U9159 (N_9159,N_8401,N_8729);
nand U9160 (N_9160,N_8728,N_8486);
or U9161 (N_9161,N_8332,N_8475);
or U9162 (N_9162,N_8716,N_8228);
nor U9163 (N_9163,N_8406,N_8175);
and U9164 (N_9164,N_8144,N_8614);
or U9165 (N_9165,N_8628,N_8202);
nand U9166 (N_9166,N_8565,N_8655);
and U9167 (N_9167,N_8579,N_8227);
or U9168 (N_9168,N_8463,N_8525);
xnor U9169 (N_9169,N_8654,N_8132);
xor U9170 (N_9170,N_8747,N_8481);
xnor U9171 (N_9171,N_8280,N_8417);
or U9172 (N_9172,N_8331,N_8188);
xnor U9173 (N_9173,N_8502,N_8169);
or U9174 (N_9174,N_8439,N_8318);
xnor U9175 (N_9175,N_8459,N_8672);
xnor U9176 (N_9176,N_8605,N_8514);
nand U9177 (N_9177,N_8300,N_8233);
nand U9178 (N_9178,N_8523,N_8406);
and U9179 (N_9179,N_8557,N_8558);
and U9180 (N_9180,N_8624,N_8193);
and U9181 (N_9181,N_8734,N_8685);
or U9182 (N_9182,N_8137,N_8675);
or U9183 (N_9183,N_8694,N_8337);
or U9184 (N_9184,N_8686,N_8426);
and U9185 (N_9185,N_8259,N_8304);
or U9186 (N_9186,N_8274,N_8557);
xor U9187 (N_9187,N_8664,N_8507);
nor U9188 (N_9188,N_8456,N_8434);
nor U9189 (N_9189,N_8515,N_8737);
xnor U9190 (N_9190,N_8321,N_8587);
and U9191 (N_9191,N_8230,N_8534);
and U9192 (N_9192,N_8711,N_8395);
xor U9193 (N_9193,N_8275,N_8541);
nor U9194 (N_9194,N_8220,N_8190);
or U9195 (N_9195,N_8638,N_8492);
and U9196 (N_9196,N_8291,N_8401);
xnor U9197 (N_9197,N_8550,N_8603);
or U9198 (N_9198,N_8388,N_8386);
nor U9199 (N_9199,N_8672,N_8300);
or U9200 (N_9200,N_8229,N_8270);
xor U9201 (N_9201,N_8243,N_8237);
or U9202 (N_9202,N_8733,N_8158);
or U9203 (N_9203,N_8167,N_8330);
nor U9204 (N_9204,N_8745,N_8653);
and U9205 (N_9205,N_8127,N_8454);
nand U9206 (N_9206,N_8210,N_8321);
nand U9207 (N_9207,N_8190,N_8729);
nor U9208 (N_9208,N_8376,N_8627);
nor U9209 (N_9209,N_8182,N_8467);
or U9210 (N_9210,N_8391,N_8246);
xnor U9211 (N_9211,N_8423,N_8696);
xnor U9212 (N_9212,N_8333,N_8555);
xor U9213 (N_9213,N_8669,N_8338);
nand U9214 (N_9214,N_8330,N_8676);
or U9215 (N_9215,N_8237,N_8512);
and U9216 (N_9216,N_8646,N_8333);
nor U9217 (N_9217,N_8651,N_8367);
nor U9218 (N_9218,N_8241,N_8737);
and U9219 (N_9219,N_8377,N_8533);
or U9220 (N_9220,N_8745,N_8192);
nand U9221 (N_9221,N_8737,N_8199);
nand U9222 (N_9222,N_8159,N_8518);
nor U9223 (N_9223,N_8375,N_8390);
and U9224 (N_9224,N_8552,N_8596);
or U9225 (N_9225,N_8671,N_8458);
or U9226 (N_9226,N_8146,N_8311);
and U9227 (N_9227,N_8565,N_8710);
nor U9228 (N_9228,N_8593,N_8675);
xnor U9229 (N_9229,N_8309,N_8375);
nor U9230 (N_9230,N_8259,N_8305);
nand U9231 (N_9231,N_8515,N_8313);
and U9232 (N_9232,N_8228,N_8199);
nor U9233 (N_9233,N_8381,N_8167);
xor U9234 (N_9234,N_8247,N_8631);
or U9235 (N_9235,N_8189,N_8297);
nand U9236 (N_9236,N_8565,N_8625);
nand U9237 (N_9237,N_8326,N_8332);
or U9238 (N_9238,N_8529,N_8648);
nor U9239 (N_9239,N_8714,N_8428);
or U9240 (N_9240,N_8206,N_8715);
or U9241 (N_9241,N_8647,N_8344);
or U9242 (N_9242,N_8348,N_8496);
nor U9243 (N_9243,N_8308,N_8386);
or U9244 (N_9244,N_8140,N_8670);
nand U9245 (N_9245,N_8659,N_8570);
nand U9246 (N_9246,N_8449,N_8415);
xor U9247 (N_9247,N_8310,N_8358);
nor U9248 (N_9248,N_8743,N_8535);
nand U9249 (N_9249,N_8136,N_8234);
nor U9250 (N_9250,N_8191,N_8223);
nand U9251 (N_9251,N_8474,N_8259);
nand U9252 (N_9252,N_8140,N_8690);
nor U9253 (N_9253,N_8707,N_8380);
or U9254 (N_9254,N_8359,N_8242);
nor U9255 (N_9255,N_8577,N_8490);
nor U9256 (N_9256,N_8294,N_8330);
nand U9257 (N_9257,N_8172,N_8176);
nand U9258 (N_9258,N_8564,N_8246);
nor U9259 (N_9259,N_8476,N_8539);
or U9260 (N_9260,N_8172,N_8639);
nor U9261 (N_9261,N_8510,N_8219);
and U9262 (N_9262,N_8620,N_8593);
nand U9263 (N_9263,N_8152,N_8316);
nor U9264 (N_9264,N_8499,N_8602);
and U9265 (N_9265,N_8535,N_8226);
and U9266 (N_9266,N_8384,N_8652);
nor U9267 (N_9267,N_8457,N_8308);
and U9268 (N_9268,N_8740,N_8171);
nand U9269 (N_9269,N_8384,N_8477);
or U9270 (N_9270,N_8589,N_8217);
nor U9271 (N_9271,N_8622,N_8295);
nor U9272 (N_9272,N_8595,N_8451);
or U9273 (N_9273,N_8472,N_8393);
nor U9274 (N_9274,N_8683,N_8315);
nor U9275 (N_9275,N_8344,N_8372);
and U9276 (N_9276,N_8726,N_8163);
nor U9277 (N_9277,N_8574,N_8341);
and U9278 (N_9278,N_8631,N_8637);
or U9279 (N_9279,N_8145,N_8497);
nor U9280 (N_9280,N_8666,N_8724);
nand U9281 (N_9281,N_8733,N_8166);
or U9282 (N_9282,N_8165,N_8470);
and U9283 (N_9283,N_8507,N_8215);
and U9284 (N_9284,N_8156,N_8159);
xor U9285 (N_9285,N_8527,N_8559);
or U9286 (N_9286,N_8143,N_8596);
nor U9287 (N_9287,N_8175,N_8723);
nor U9288 (N_9288,N_8352,N_8451);
or U9289 (N_9289,N_8171,N_8603);
or U9290 (N_9290,N_8180,N_8338);
or U9291 (N_9291,N_8700,N_8661);
or U9292 (N_9292,N_8478,N_8511);
and U9293 (N_9293,N_8171,N_8377);
xnor U9294 (N_9294,N_8353,N_8668);
or U9295 (N_9295,N_8475,N_8511);
and U9296 (N_9296,N_8255,N_8611);
and U9297 (N_9297,N_8578,N_8379);
nor U9298 (N_9298,N_8383,N_8414);
nor U9299 (N_9299,N_8588,N_8473);
or U9300 (N_9300,N_8705,N_8572);
or U9301 (N_9301,N_8555,N_8537);
or U9302 (N_9302,N_8188,N_8397);
and U9303 (N_9303,N_8339,N_8367);
nand U9304 (N_9304,N_8449,N_8607);
nand U9305 (N_9305,N_8368,N_8515);
and U9306 (N_9306,N_8232,N_8289);
or U9307 (N_9307,N_8401,N_8608);
nor U9308 (N_9308,N_8546,N_8703);
nor U9309 (N_9309,N_8566,N_8739);
xor U9310 (N_9310,N_8718,N_8347);
nor U9311 (N_9311,N_8731,N_8405);
xnor U9312 (N_9312,N_8703,N_8182);
nand U9313 (N_9313,N_8213,N_8442);
and U9314 (N_9314,N_8497,N_8629);
nor U9315 (N_9315,N_8315,N_8678);
nor U9316 (N_9316,N_8491,N_8199);
nand U9317 (N_9317,N_8599,N_8636);
xor U9318 (N_9318,N_8617,N_8132);
or U9319 (N_9319,N_8367,N_8232);
and U9320 (N_9320,N_8725,N_8298);
nor U9321 (N_9321,N_8350,N_8748);
xnor U9322 (N_9322,N_8536,N_8503);
and U9323 (N_9323,N_8493,N_8254);
nor U9324 (N_9324,N_8706,N_8194);
xor U9325 (N_9325,N_8520,N_8271);
or U9326 (N_9326,N_8396,N_8273);
and U9327 (N_9327,N_8128,N_8343);
or U9328 (N_9328,N_8633,N_8604);
xnor U9329 (N_9329,N_8625,N_8164);
nor U9330 (N_9330,N_8686,N_8627);
or U9331 (N_9331,N_8125,N_8185);
nand U9332 (N_9332,N_8397,N_8358);
and U9333 (N_9333,N_8694,N_8686);
nor U9334 (N_9334,N_8503,N_8446);
nor U9335 (N_9335,N_8375,N_8176);
xor U9336 (N_9336,N_8370,N_8679);
nand U9337 (N_9337,N_8509,N_8153);
or U9338 (N_9338,N_8723,N_8610);
nand U9339 (N_9339,N_8731,N_8226);
nor U9340 (N_9340,N_8703,N_8448);
nand U9341 (N_9341,N_8128,N_8213);
or U9342 (N_9342,N_8466,N_8371);
nand U9343 (N_9343,N_8439,N_8181);
nor U9344 (N_9344,N_8389,N_8736);
nor U9345 (N_9345,N_8378,N_8674);
nor U9346 (N_9346,N_8317,N_8621);
nor U9347 (N_9347,N_8366,N_8377);
and U9348 (N_9348,N_8285,N_8396);
nand U9349 (N_9349,N_8230,N_8151);
and U9350 (N_9350,N_8202,N_8322);
or U9351 (N_9351,N_8475,N_8254);
nand U9352 (N_9352,N_8746,N_8187);
and U9353 (N_9353,N_8529,N_8371);
and U9354 (N_9354,N_8241,N_8659);
or U9355 (N_9355,N_8640,N_8679);
nand U9356 (N_9356,N_8712,N_8611);
nor U9357 (N_9357,N_8514,N_8171);
and U9358 (N_9358,N_8714,N_8156);
nor U9359 (N_9359,N_8445,N_8209);
and U9360 (N_9360,N_8706,N_8554);
or U9361 (N_9361,N_8274,N_8296);
and U9362 (N_9362,N_8202,N_8443);
nor U9363 (N_9363,N_8542,N_8560);
nand U9364 (N_9364,N_8659,N_8663);
and U9365 (N_9365,N_8309,N_8747);
nand U9366 (N_9366,N_8412,N_8235);
nor U9367 (N_9367,N_8290,N_8223);
nand U9368 (N_9368,N_8395,N_8606);
and U9369 (N_9369,N_8390,N_8262);
nor U9370 (N_9370,N_8375,N_8473);
and U9371 (N_9371,N_8279,N_8511);
nand U9372 (N_9372,N_8240,N_8336);
nand U9373 (N_9373,N_8169,N_8131);
and U9374 (N_9374,N_8407,N_8472);
nand U9375 (N_9375,N_8811,N_9373);
or U9376 (N_9376,N_9163,N_9333);
and U9377 (N_9377,N_9087,N_9152);
nand U9378 (N_9378,N_9208,N_8902);
or U9379 (N_9379,N_9191,N_8840);
nand U9380 (N_9380,N_9094,N_9291);
or U9381 (N_9381,N_8918,N_9196);
nand U9382 (N_9382,N_8927,N_8890);
and U9383 (N_9383,N_9008,N_9283);
or U9384 (N_9384,N_8973,N_9274);
and U9385 (N_9385,N_8858,N_8767);
nor U9386 (N_9386,N_9200,N_9019);
and U9387 (N_9387,N_9162,N_9301);
nor U9388 (N_9388,N_8916,N_8929);
nand U9389 (N_9389,N_9088,N_9022);
or U9390 (N_9390,N_9270,N_9300);
nor U9391 (N_9391,N_9329,N_9172);
nor U9392 (N_9392,N_9254,N_9101);
or U9393 (N_9393,N_9272,N_9319);
nor U9394 (N_9394,N_9238,N_9122);
nor U9395 (N_9395,N_9137,N_8843);
and U9396 (N_9396,N_9289,N_9044);
nor U9397 (N_9397,N_8752,N_9117);
nand U9398 (N_9398,N_8839,N_9089);
nor U9399 (N_9399,N_9280,N_8938);
nand U9400 (N_9400,N_9212,N_9339);
nand U9401 (N_9401,N_8987,N_9343);
or U9402 (N_9402,N_9344,N_9083);
or U9403 (N_9403,N_8755,N_9129);
and U9404 (N_9404,N_9056,N_9158);
nor U9405 (N_9405,N_9345,N_9322);
nor U9406 (N_9406,N_9355,N_8917);
nor U9407 (N_9407,N_9231,N_9215);
nor U9408 (N_9408,N_9228,N_8930);
or U9409 (N_9409,N_9264,N_8985);
nand U9410 (N_9410,N_8812,N_8928);
nand U9411 (N_9411,N_9335,N_9229);
or U9412 (N_9412,N_8763,N_9029);
or U9413 (N_9413,N_8813,N_9055);
nand U9414 (N_9414,N_9247,N_9020);
and U9415 (N_9415,N_8941,N_9279);
nor U9416 (N_9416,N_9311,N_9031);
nor U9417 (N_9417,N_9276,N_9351);
and U9418 (N_9418,N_8801,N_9237);
or U9419 (N_9419,N_9116,N_8889);
and U9420 (N_9420,N_8807,N_9104);
and U9421 (N_9421,N_9001,N_9060);
xnor U9422 (N_9422,N_8977,N_9077);
nand U9423 (N_9423,N_9364,N_9176);
or U9424 (N_9424,N_9041,N_8814);
and U9425 (N_9425,N_9277,N_8903);
or U9426 (N_9426,N_8923,N_8764);
and U9427 (N_9427,N_8900,N_9282);
or U9428 (N_9428,N_8794,N_8921);
nand U9429 (N_9429,N_8831,N_8966);
nand U9430 (N_9430,N_9002,N_8782);
nand U9431 (N_9431,N_8957,N_9256);
and U9432 (N_9432,N_9181,N_8924);
nand U9433 (N_9433,N_9051,N_9246);
nor U9434 (N_9434,N_8787,N_9033);
nor U9435 (N_9435,N_8778,N_8759);
and U9436 (N_9436,N_9188,N_9170);
nand U9437 (N_9437,N_9120,N_9128);
nor U9438 (N_9438,N_9146,N_9302);
nand U9439 (N_9439,N_9253,N_8896);
xor U9440 (N_9440,N_9349,N_8974);
and U9441 (N_9441,N_8848,N_8783);
xnor U9442 (N_9442,N_8994,N_9049);
or U9443 (N_9443,N_9211,N_9261);
nand U9444 (N_9444,N_9216,N_9086);
nand U9445 (N_9445,N_9227,N_9014);
nor U9446 (N_9446,N_8835,N_9263);
xor U9447 (N_9447,N_8969,N_9091);
nand U9448 (N_9448,N_9371,N_8789);
or U9449 (N_9449,N_8982,N_8798);
nor U9450 (N_9450,N_8857,N_9037);
or U9451 (N_9451,N_8867,N_8976);
or U9452 (N_9452,N_9245,N_8965);
and U9453 (N_9453,N_8954,N_8815);
and U9454 (N_9454,N_8873,N_8905);
nand U9455 (N_9455,N_9140,N_8754);
nand U9456 (N_9456,N_8955,N_8868);
nand U9457 (N_9457,N_8980,N_9007);
nand U9458 (N_9458,N_9171,N_8834);
and U9459 (N_9459,N_8855,N_9076);
or U9460 (N_9460,N_8978,N_9219);
nor U9461 (N_9461,N_8971,N_9090);
nor U9462 (N_9462,N_9178,N_9205);
or U9463 (N_9463,N_9063,N_9017);
or U9464 (N_9464,N_9099,N_9258);
and U9465 (N_9465,N_8911,N_8849);
or U9466 (N_9466,N_9092,N_9348);
nor U9467 (N_9467,N_9106,N_9326);
or U9468 (N_9468,N_9127,N_8963);
and U9469 (N_9469,N_8786,N_8962);
and U9470 (N_9470,N_9287,N_8845);
and U9471 (N_9471,N_9134,N_9187);
and U9472 (N_9472,N_8934,N_8997);
and U9473 (N_9473,N_8960,N_9290);
and U9474 (N_9474,N_9168,N_8940);
or U9475 (N_9475,N_9241,N_8820);
or U9476 (N_9476,N_8784,N_9011);
and U9477 (N_9477,N_9043,N_9341);
nor U9478 (N_9478,N_8829,N_8853);
or U9479 (N_9479,N_9251,N_9233);
nand U9480 (N_9480,N_8931,N_9038);
nor U9481 (N_9481,N_9209,N_9213);
or U9482 (N_9482,N_9367,N_9295);
xor U9483 (N_9483,N_9347,N_9123);
or U9484 (N_9484,N_8768,N_9308);
nor U9485 (N_9485,N_9198,N_9113);
xnor U9486 (N_9486,N_9214,N_8959);
and U9487 (N_9487,N_8950,N_9052);
and U9488 (N_9488,N_9275,N_9000);
or U9489 (N_9489,N_8935,N_9066);
and U9490 (N_9490,N_9336,N_8964);
nor U9491 (N_9491,N_9353,N_9081);
and U9492 (N_9492,N_8888,N_9201);
and U9493 (N_9493,N_8975,N_9357);
nor U9494 (N_9494,N_8785,N_9374);
or U9495 (N_9495,N_8810,N_9299);
nor U9496 (N_9496,N_8972,N_9346);
and U9497 (N_9497,N_9139,N_9225);
xor U9498 (N_9498,N_9165,N_8949);
nor U9499 (N_9499,N_8753,N_9065);
and U9500 (N_9500,N_8750,N_8979);
xnor U9501 (N_9501,N_8799,N_9332);
nor U9502 (N_9502,N_8875,N_8821);
nand U9503 (N_9503,N_8886,N_8922);
and U9504 (N_9504,N_8866,N_8894);
and U9505 (N_9505,N_9175,N_8989);
nor U9506 (N_9506,N_9135,N_9136);
nand U9507 (N_9507,N_9222,N_9255);
nor U9508 (N_9508,N_9138,N_9284);
or U9509 (N_9509,N_9054,N_9061);
nand U9510 (N_9510,N_9110,N_9350);
nand U9511 (N_9511,N_9325,N_9318);
xnor U9512 (N_9512,N_8915,N_9169);
xor U9513 (N_9513,N_9012,N_9015);
and U9514 (N_9514,N_9234,N_9124);
or U9515 (N_9515,N_9070,N_9132);
or U9516 (N_9516,N_8774,N_8912);
and U9517 (N_9517,N_8939,N_9189);
nand U9518 (N_9518,N_8968,N_9100);
and U9519 (N_9519,N_9072,N_8914);
nor U9520 (N_9520,N_8961,N_8762);
nor U9521 (N_9521,N_9257,N_9036);
nor U9522 (N_9522,N_9159,N_8932);
or U9523 (N_9523,N_9224,N_8808);
or U9524 (N_9524,N_8956,N_9317);
and U9525 (N_9525,N_9309,N_9085);
nand U9526 (N_9526,N_9082,N_9179);
nor U9527 (N_9527,N_8942,N_9084);
nand U9528 (N_9528,N_8862,N_9292);
and U9529 (N_9529,N_9243,N_9330);
nor U9530 (N_9530,N_8993,N_9018);
or U9531 (N_9531,N_9267,N_9078);
and U9532 (N_9532,N_8816,N_9260);
and U9533 (N_9533,N_9195,N_9107);
nor U9534 (N_9534,N_9236,N_9126);
nand U9535 (N_9535,N_9230,N_9361);
nand U9536 (N_9536,N_8995,N_9217);
xor U9537 (N_9537,N_9109,N_9321);
nor U9538 (N_9538,N_9358,N_8756);
and U9539 (N_9539,N_9304,N_9111);
or U9540 (N_9540,N_8766,N_9006);
nor U9541 (N_9541,N_9337,N_9142);
xnor U9542 (N_9542,N_9320,N_8830);
nand U9543 (N_9543,N_8871,N_9183);
or U9544 (N_9544,N_8908,N_8906);
nor U9545 (N_9545,N_9003,N_8832);
nor U9546 (N_9546,N_9206,N_8802);
nand U9547 (N_9547,N_9324,N_9210);
nand U9548 (N_9548,N_9125,N_8856);
nand U9549 (N_9549,N_8952,N_8945);
and U9550 (N_9550,N_9197,N_9312);
nor U9551 (N_9551,N_9259,N_9194);
and U9552 (N_9552,N_9298,N_9069);
and U9553 (N_9553,N_8991,N_9306);
nand U9554 (N_9554,N_9164,N_9133);
xor U9555 (N_9555,N_8898,N_9368);
xor U9556 (N_9556,N_9080,N_9369);
and U9557 (N_9557,N_8877,N_9173);
xor U9558 (N_9558,N_9067,N_8988);
nor U9559 (N_9559,N_9232,N_9244);
and U9560 (N_9560,N_9262,N_9064);
and U9561 (N_9561,N_8919,N_8836);
and U9562 (N_9562,N_9004,N_9204);
and U9563 (N_9563,N_9016,N_9248);
nor U9564 (N_9564,N_8761,N_9294);
and U9565 (N_9565,N_9121,N_9340);
nor U9566 (N_9566,N_8775,N_8792);
nor U9567 (N_9567,N_8805,N_9093);
nor U9568 (N_9568,N_9160,N_8951);
nor U9569 (N_9569,N_8854,N_9156);
nor U9570 (N_9570,N_9153,N_9058);
and U9571 (N_9571,N_9118,N_8946);
and U9572 (N_9572,N_8891,N_8795);
nor U9573 (N_9573,N_8850,N_9108);
nand U9574 (N_9574,N_9186,N_9334);
nand U9575 (N_9575,N_9226,N_9150);
nand U9576 (N_9576,N_8851,N_9147);
nand U9577 (N_9577,N_9269,N_9218);
xnor U9578 (N_9578,N_9073,N_8899);
and U9579 (N_9579,N_8874,N_9313);
nor U9580 (N_9580,N_8758,N_9202);
and U9581 (N_9581,N_9105,N_8992);
nand U9582 (N_9582,N_9266,N_9161);
nand U9583 (N_9583,N_9119,N_9207);
nor U9584 (N_9584,N_9250,N_8937);
or U9585 (N_9585,N_8804,N_8844);
nand U9586 (N_9586,N_8953,N_8859);
and U9587 (N_9587,N_9285,N_8885);
xnor U9588 (N_9588,N_8852,N_9115);
nand U9589 (N_9589,N_9028,N_9039);
nand U9590 (N_9590,N_9013,N_9167);
nor U9591 (N_9591,N_9102,N_9112);
xnor U9592 (N_9592,N_9045,N_9323);
nor U9593 (N_9593,N_8860,N_9235);
and U9594 (N_9594,N_9268,N_8773);
nand U9595 (N_9595,N_8878,N_9166);
or U9596 (N_9596,N_8925,N_9095);
nand U9597 (N_9597,N_9221,N_9370);
or U9598 (N_9598,N_9252,N_8800);
and U9599 (N_9599,N_9303,N_8863);
or U9600 (N_9600,N_9075,N_9356);
nand U9601 (N_9601,N_8892,N_9372);
or U9602 (N_9602,N_9316,N_9293);
nor U9603 (N_9603,N_8781,N_9149);
and U9604 (N_9604,N_8779,N_8788);
and U9605 (N_9605,N_8999,N_9145);
and U9606 (N_9606,N_8948,N_9046);
nand U9607 (N_9607,N_8796,N_8895);
and U9608 (N_9608,N_8826,N_9114);
or U9609 (N_9609,N_9366,N_9062);
nor U9610 (N_9610,N_8825,N_8827);
nand U9611 (N_9611,N_8757,N_9151);
and U9612 (N_9612,N_8819,N_8824);
nand U9613 (N_9613,N_8970,N_9297);
nor U9614 (N_9614,N_9286,N_9193);
and U9615 (N_9615,N_9071,N_8984);
nor U9616 (N_9616,N_8791,N_8909);
nand U9617 (N_9617,N_8864,N_8881);
or U9618 (N_9618,N_8828,N_8842);
nor U9619 (N_9619,N_9050,N_9131);
nand U9620 (N_9620,N_9199,N_9310);
xnor U9621 (N_9621,N_9034,N_8780);
nand U9622 (N_9622,N_9010,N_8771);
nor U9623 (N_9623,N_8803,N_8838);
nand U9624 (N_9624,N_9360,N_8887);
or U9625 (N_9625,N_9103,N_8947);
and U9626 (N_9626,N_9155,N_8933);
and U9627 (N_9627,N_9338,N_9240);
or U9628 (N_9628,N_9154,N_9185);
nor U9629 (N_9629,N_8846,N_9362);
nor U9630 (N_9630,N_8861,N_9024);
nand U9631 (N_9631,N_9030,N_8772);
or U9632 (N_9632,N_8876,N_9192);
or U9633 (N_9633,N_9203,N_9327);
nor U9634 (N_9634,N_8770,N_8882);
and U9635 (N_9635,N_9288,N_9365);
nor U9636 (N_9636,N_9068,N_9220);
nand U9637 (N_9637,N_9021,N_8967);
xnor U9638 (N_9638,N_9074,N_8913);
nand U9639 (N_9639,N_8823,N_9059);
nor U9640 (N_9640,N_8926,N_8793);
nor U9641 (N_9641,N_8777,N_8883);
and U9642 (N_9642,N_9130,N_9177);
or U9643 (N_9643,N_9184,N_8879);
nand U9644 (N_9644,N_9035,N_9025);
nor U9645 (N_9645,N_9032,N_9180);
nor U9646 (N_9646,N_9042,N_9182);
xnor U9647 (N_9647,N_8833,N_8776);
xor U9648 (N_9648,N_8817,N_9190);
xnor U9649 (N_9649,N_9359,N_9296);
nand U9650 (N_9650,N_9331,N_8769);
and U9651 (N_9651,N_8809,N_9098);
or U9652 (N_9652,N_9239,N_8958);
nor U9653 (N_9653,N_9097,N_9148);
nand U9654 (N_9654,N_8872,N_9223);
xor U9655 (N_9655,N_9281,N_9305);
or U9656 (N_9656,N_8818,N_8751);
nor U9657 (N_9657,N_9157,N_9315);
and U9658 (N_9658,N_8822,N_8990);
nand U9659 (N_9659,N_8904,N_9023);
and U9660 (N_9660,N_9307,N_9040);
or U9661 (N_9661,N_8841,N_9048);
or U9662 (N_9662,N_8943,N_8806);
or U9663 (N_9663,N_8996,N_8986);
and U9664 (N_9664,N_9026,N_8981);
nand U9665 (N_9665,N_9053,N_8847);
nor U9666 (N_9666,N_8983,N_8865);
xor U9667 (N_9667,N_9143,N_8880);
nand U9668 (N_9668,N_9079,N_8797);
or U9669 (N_9669,N_9363,N_8998);
or U9670 (N_9670,N_8760,N_8893);
or U9671 (N_9671,N_8901,N_8870);
nand U9672 (N_9672,N_8765,N_9265);
nor U9673 (N_9673,N_9005,N_8790);
or U9674 (N_9674,N_9342,N_9249);
nand U9675 (N_9675,N_9027,N_9278);
xnor U9676 (N_9676,N_9057,N_9047);
xnor U9677 (N_9677,N_8897,N_9328);
nand U9678 (N_9678,N_8920,N_8869);
nor U9679 (N_9679,N_8936,N_9144);
or U9680 (N_9680,N_9273,N_9271);
or U9681 (N_9681,N_9242,N_9096);
xnor U9682 (N_9682,N_8884,N_8907);
and U9683 (N_9683,N_9174,N_9009);
nor U9684 (N_9684,N_8910,N_9141);
nand U9685 (N_9685,N_9352,N_9314);
or U9686 (N_9686,N_9354,N_8944);
nand U9687 (N_9687,N_8837,N_8978);
or U9688 (N_9688,N_9297,N_8825);
nor U9689 (N_9689,N_9200,N_9004);
xor U9690 (N_9690,N_8801,N_9218);
and U9691 (N_9691,N_9315,N_8851);
and U9692 (N_9692,N_9070,N_9239);
or U9693 (N_9693,N_8916,N_9053);
or U9694 (N_9694,N_9116,N_9201);
nor U9695 (N_9695,N_9194,N_8899);
nand U9696 (N_9696,N_8907,N_9179);
xnor U9697 (N_9697,N_8820,N_9006);
nand U9698 (N_9698,N_9164,N_8786);
or U9699 (N_9699,N_9170,N_9209);
nor U9700 (N_9700,N_8906,N_8985);
nand U9701 (N_9701,N_8770,N_8920);
and U9702 (N_9702,N_9026,N_9203);
nand U9703 (N_9703,N_8896,N_8767);
xor U9704 (N_9704,N_8929,N_8875);
nor U9705 (N_9705,N_8861,N_9308);
and U9706 (N_9706,N_8793,N_9141);
nand U9707 (N_9707,N_8758,N_8982);
xnor U9708 (N_9708,N_9199,N_9186);
or U9709 (N_9709,N_8869,N_8940);
nor U9710 (N_9710,N_8919,N_9067);
nand U9711 (N_9711,N_8857,N_9044);
and U9712 (N_9712,N_9054,N_9128);
nor U9713 (N_9713,N_9226,N_9146);
nand U9714 (N_9714,N_9315,N_9370);
nor U9715 (N_9715,N_9105,N_9370);
nor U9716 (N_9716,N_8982,N_8768);
and U9717 (N_9717,N_8815,N_9373);
nand U9718 (N_9718,N_8962,N_8911);
and U9719 (N_9719,N_8809,N_9070);
nand U9720 (N_9720,N_9308,N_9265);
nor U9721 (N_9721,N_8925,N_9150);
nand U9722 (N_9722,N_8893,N_9188);
nor U9723 (N_9723,N_9233,N_8999);
and U9724 (N_9724,N_9347,N_9096);
and U9725 (N_9725,N_9246,N_9119);
or U9726 (N_9726,N_9298,N_9239);
nand U9727 (N_9727,N_9350,N_9157);
nor U9728 (N_9728,N_9103,N_9262);
or U9729 (N_9729,N_9360,N_8758);
nand U9730 (N_9730,N_9005,N_8822);
or U9731 (N_9731,N_9278,N_8827);
xnor U9732 (N_9732,N_9316,N_9297);
nor U9733 (N_9733,N_8806,N_9346);
nor U9734 (N_9734,N_8989,N_8934);
xor U9735 (N_9735,N_9202,N_8985);
xnor U9736 (N_9736,N_9215,N_8976);
nor U9737 (N_9737,N_8986,N_8860);
nor U9738 (N_9738,N_8780,N_8950);
xnor U9739 (N_9739,N_8971,N_8984);
and U9740 (N_9740,N_8834,N_9292);
or U9741 (N_9741,N_8799,N_8777);
or U9742 (N_9742,N_9137,N_9332);
nand U9743 (N_9743,N_8887,N_9033);
or U9744 (N_9744,N_8957,N_8904);
nor U9745 (N_9745,N_9346,N_9349);
and U9746 (N_9746,N_8915,N_9343);
xnor U9747 (N_9747,N_9286,N_8932);
nor U9748 (N_9748,N_9000,N_8797);
and U9749 (N_9749,N_9310,N_8987);
xor U9750 (N_9750,N_9143,N_8829);
or U9751 (N_9751,N_8832,N_9019);
or U9752 (N_9752,N_8827,N_9022);
nand U9753 (N_9753,N_9145,N_8798);
nand U9754 (N_9754,N_9138,N_9224);
nor U9755 (N_9755,N_9098,N_8968);
nor U9756 (N_9756,N_8983,N_8932);
nor U9757 (N_9757,N_8854,N_9229);
nor U9758 (N_9758,N_9028,N_9043);
xnor U9759 (N_9759,N_9198,N_8751);
xnor U9760 (N_9760,N_9311,N_9270);
and U9761 (N_9761,N_8769,N_9208);
nor U9762 (N_9762,N_9007,N_8936);
xor U9763 (N_9763,N_9286,N_9256);
or U9764 (N_9764,N_9248,N_9094);
or U9765 (N_9765,N_9167,N_9297);
nand U9766 (N_9766,N_9325,N_9202);
nor U9767 (N_9767,N_9353,N_8810);
nand U9768 (N_9768,N_9009,N_8903);
nand U9769 (N_9769,N_8968,N_9134);
nor U9770 (N_9770,N_9333,N_8838);
nand U9771 (N_9771,N_9157,N_9368);
and U9772 (N_9772,N_8963,N_8756);
or U9773 (N_9773,N_8918,N_9034);
and U9774 (N_9774,N_9337,N_9226);
nor U9775 (N_9775,N_9034,N_9178);
and U9776 (N_9776,N_8973,N_9190);
or U9777 (N_9777,N_9296,N_9197);
and U9778 (N_9778,N_8986,N_9370);
and U9779 (N_9779,N_9321,N_8923);
xnor U9780 (N_9780,N_9192,N_8797);
nor U9781 (N_9781,N_9195,N_8950);
or U9782 (N_9782,N_8904,N_8963);
and U9783 (N_9783,N_8829,N_9015);
xor U9784 (N_9784,N_9373,N_9366);
nand U9785 (N_9785,N_8948,N_8764);
and U9786 (N_9786,N_8812,N_9155);
and U9787 (N_9787,N_9100,N_9216);
and U9788 (N_9788,N_9315,N_9179);
and U9789 (N_9789,N_8914,N_9092);
or U9790 (N_9790,N_9090,N_9288);
and U9791 (N_9791,N_8789,N_8824);
or U9792 (N_9792,N_9184,N_9015);
or U9793 (N_9793,N_9051,N_8924);
and U9794 (N_9794,N_9153,N_9241);
or U9795 (N_9795,N_8756,N_9192);
or U9796 (N_9796,N_9145,N_9015);
xor U9797 (N_9797,N_9354,N_8959);
and U9798 (N_9798,N_9127,N_9038);
and U9799 (N_9799,N_8878,N_9221);
and U9800 (N_9800,N_9273,N_9043);
nand U9801 (N_9801,N_9241,N_8976);
nor U9802 (N_9802,N_8932,N_9019);
or U9803 (N_9803,N_9072,N_9160);
or U9804 (N_9804,N_8952,N_9357);
and U9805 (N_9805,N_9055,N_8824);
nor U9806 (N_9806,N_9153,N_8920);
and U9807 (N_9807,N_8830,N_9023);
xor U9808 (N_9808,N_8797,N_9233);
or U9809 (N_9809,N_8787,N_9098);
or U9810 (N_9810,N_8993,N_9257);
and U9811 (N_9811,N_9327,N_9054);
or U9812 (N_9812,N_8833,N_9146);
xnor U9813 (N_9813,N_8982,N_9054);
and U9814 (N_9814,N_9032,N_8955);
and U9815 (N_9815,N_8760,N_9353);
xor U9816 (N_9816,N_9211,N_9158);
nor U9817 (N_9817,N_8780,N_9022);
and U9818 (N_9818,N_8851,N_9078);
or U9819 (N_9819,N_9000,N_8763);
nand U9820 (N_9820,N_9218,N_9123);
nand U9821 (N_9821,N_9254,N_9287);
and U9822 (N_9822,N_8867,N_9242);
nor U9823 (N_9823,N_8838,N_8976);
xor U9824 (N_9824,N_8852,N_9220);
and U9825 (N_9825,N_8786,N_9283);
or U9826 (N_9826,N_9020,N_9110);
nor U9827 (N_9827,N_8801,N_8803);
nor U9828 (N_9828,N_8791,N_8801);
or U9829 (N_9829,N_9119,N_8963);
nand U9830 (N_9830,N_9252,N_9196);
xor U9831 (N_9831,N_9000,N_8912);
nand U9832 (N_9832,N_8924,N_8977);
or U9833 (N_9833,N_9251,N_8897);
xnor U9834 (N_9834,N_9101,N_8876);
and U9835 (N_9835,N_9348,N_9364);
nor U9836 (N_9836,N_9280,N_9158);
and U9837 (N_9837,N_9279,N_8755);
and U9838 (N_9838,N_8859,N_8910);
nor U9839 (N_9839,N_9149,N_8753);
nor U9840 (N_9840,N_9018,N_9120);
nor U9841 (N_9841,N_9371,N_9252);
nor U9842 (N_9842,N_9289,N_9094);
and U9843 (N_9843,N_9100,N_9266);
xor U9844 (N_9844,N_8969,N_8763);
nor U9845 (N_9845,N_9371,N_8824);
or U9846 (N_9846,N_9304,N_8752);
and U9847 (N_9847,N_8945,N_8918);
or U9848 (N_9848,N_8780,N_8834);
nand U9849 (N_9849,N_8990,N_8898);
nor U9850 (N_9850,N_9249,N_8805);
nor U9851 (N_9851,N_9203,N_9045);
or U9852 (N_9852,N_9184,N_9187);
nand U9853 (N_9853,N_9067,N_9059);
or U9854 (N_9854,N_9028,N_9066);
nand U9855 (N_9855,N_8761,N_8835);
nor U9856 (N_9856,N_8972,N_8875);
xor U9857 (N_9857,N_9081,N_8945);
or U9858 (N_9858,N_9159,N_8944);
nor U9859 (N_9859,N_8818,N_9176);
and U9860 (N_9860,N_9178,N_9113);
nand U9861 (N_9861,N_8845,N_9092);
or U9862 (N_9862,N_9139,N_9224);
or U9863 (N_9863,N_9125,N_8885);
and U9864 (N_9864,N_9154,N_9341);
and U9865 (N_9865,N_9316,N_9046);
nor U9866 (N_9866,N_8903,N_9195);
and U9867 (N_9867,N_9304,N_8965);
nand U9868 (N_9868,N_9199,N_9373);
nor U9869 (N_9869,N_9326,N_9099);
and U9870 (N_9870,N_9208,N_9066);
nor U9871 (N_9871,N_9107,N_8934);
or U9872 (N_9872,N_9232,N_9034);
nand U9873 (N_9873,N_9070,N_8952);
nor U9874 (N_9874,N_9126,N_9357);
nand U9875 (N_9875,N_9217,N_9337);
nor U9876 (N_9876,N_9241,N_8822);
and U9877 (N_9877,N_8922,N_9301);
nor U9878 (N_9878,N_9019,N_8920);
nor U9879 (N_9879,N_9268,N_9049);
and U9880 (N_9880,N_8907,N_8951);
or U9881 (N_9881,N_8772,N_9187);
nor U9882 (N_9882,N_9322,N_8893);
nand U9883 (N_9883,N_9172,N_9353);
nand U9884 (N_9884,N_8970,N_9186);
or U9885 (N_9885,N_8961,N_8839);
and U9886 (N_9886,N_8978,N_9133);
nand U9887 (N_9887,N_9110,N_8984);
nor U9888 (N_9888,N_9118,N_9021);
nor U9889 (N_9889,N_9187,N_9225);
nor U9890 (N_9890,N_8908,N_9137);
and U9891 (N_9891,N_9314,N_9264);
nor U9892 (N_9892,N_9170,N_9094);
nor U9893 (N_9893,N_8955,N_9313);
and U9894 (N_9894,N_8858,N_9364);
nor U9895 (N_9895,N_9128,N_8872);
nand U9896 (N_9896,N_9284,N_9097);
and U9897 (N_9897,N_9179,N_8756);
nor U9898 (N_9898,N_9350,N_9213);
or U9899 (N_9899,N_8906,N_9198);
nand U9900 (N_9900,N_9119,N_9025);
xnor U9901 (N_9901,N_8922,N_9027);
nor U9902 (N_9902,N_9177,N_8988);
and U9903 (N_9903,N_9085,N_9334);
and U9904 (N_9904,N_9204,N_8807);
and U9905 (N_9905,N_8831,N_9356);
nand U9906 (N_9906,N_8810,N_9216);
or U9907 (N_9907,N_8964,N_9046);
nand U9908 (N_9908,N_9285,N_8765);
and U9909 (N_9909,N_9208,N_9133);
and U9910 (N_9910,N_9288,N_8895);
nand U9911 (N_9911,N_9220,N_8768);
or U9912 (N_9912,N_9021,N_9105);
nor U9913 (N_9913,N_8792,N_9196);
or U9914 (N_9914,N_9020,N_8957);
nand U9915 (N_9915,N_9367,N_9306);
nor U9916 (N_9916,N_9348,N_9185);
or U9917 (N_9917,N_8823,N_8989);
nor U9918 (N_9918,N_8862,N_9045);
nand U9919 (N_9919,N_9008,N_8903);
and U9920 (N_9920,N_8825,N_9068);
nor U9921 (N_9921,N_8754,N_8755);
nand U9922 (N_9922,N_9246,N_9156);
nand U9923 (N_9923,N_9140,N_8929);
xor U9924 (N_9924,N_9354,N_9248);
or U9925 (N_9925,N_9215,N_9127);
and U9926 (N_9926,N_9247,N_9173);
and U9927 (N_9927,N_9035,N_9070);
nor U9928 (N_9928,N_9189,N_8827);
and U9929 (N_9929,N_9136,N_9337);
nor U9930 (N_9930,N_8788,N_9211);
or U9931 (N_9931,N_9265,N_9195);
and U9932 (N_9932,N_9206,N_8969);
nand U9933 (N_9933,N_9133,N_8843);
nand U9934 (N_9934,N_8974,N_9210);
and U9935 (N_9935,N_9107,N_8933);
nand U9936 (N_9936,N_9172,N_9240);
nand U9937 (N_9937,N_8870,N_9308);
and U9938 (N_9938,N_8879,N_9140);
xor U9939 (N_9939,N_8808,N_8929);
nor U9940 (N_9940,N_9108,N_9242);
and U9941 (N_9941,N_8790,N_8782);
and U9942 (N_9942,N_9227,N_9193);
xnor U9943 (N_9943,N_9309,N_8847);
or U9944 (N_9944,N_9062,N_9146);
xnor U9945 (N_9945,N_9141,N_9197);
nand U9946 (N_9946,N_9352,N_9014);
nor U9947 (N_9947,N_8918,N_9286);
xor U9948 (N_9948,N_9151,N_9233);
nor U9949 (N_9949,N_9001,N_8999);
and U9950 (N_9950,N_9164,N_9316);
nand U9951 (N_9951,N_9117,N_9077);
nor U9952 (N_9952,N_9227,N_9047);
or U9953 (N_9953,N_8927,N_9175);
xnor U9954 (N_9954,N_8817,N_9350);
xor U9955 (N_9955,N_8870,N_8945);
xor U9956 (N_9956,N_9128,N_9011);
nor U9957 (N_9957,N_8964,N_9060);
and U9958 (N_9958,N_9065,N_9200);
nor U9959 (N_9959,N_9053,N_8894);
nor U9960 (N_9960,N_9098,N_9311);
nor U9961 (N_9961,N_9143,N_8988);
or U9962 (N_9962,N_8952,N_8829);
and U9963 (N_9963,N_9114,N_9310);
or U9964 (N_9964,N_9354,N_9241);
and U9965 (N_9965,N_9150,N_9371);
nand U9966 (N_9966,N_9324,N_9074);
and U9967 (N_9967,N_9207,N_9128);
nor U9968 (N_9968,N_9327,N_9068);
nand U9969 (N_9969,N_9156,N_9110);
xor U9970 (N_9970,N_8931,N_9358);
nand U9971 (N_9971,N_8891,N_9319);
and U9972 (N_9972,N_8819,N_9312);
and U9973 (N_9973,N_9269,N_8787);
or U9974 (N_9974,N_9032,N_9166);
and U9975 (N_9975,N_9173,N_8859);
or U9976 (N_9976,N_8849,N_9093);
and U9977 (N_9977,N_9179,N_8953);
or U9978 (N_9978,N_9207,N_9269);
and U9979 (N_9979,N_9196,N_9108);
nor U9980 (N_9980,N_9262,N_8945);
nor U9981 (N_9981,N_9009,N_8863);
nor U9982 (N_9982,N_9177,N_9099);
nand U9983 (N_9983,N_8981,N_9265);
and U9984 (N_9984,N_9261,N_9192);
or U9985 (N_9985,N_9351,N_9365);
nand U9986 (N_9986,N_9070,N_9312);
nand U9987 (N_9987,N_9145,N_8861);
nand U9988 (N_9988,N_9311,N_8771);
xnor U9989 (N_9989,N_9221,N_9194);
nand U9990 (N_9990,N_9303,N_9363);
nand U9991 (N_9991,N_9140,N_8987);
and U9992 (N_9992,N_9042,N_9186);
and U9993 (N_9993,N_9137,N_9221);
nor U9994 (N_9994,N_8776,N_8792);
and U9995 (N_9995,N_8840,N_8810);
nand U9996 (N_9996,N_8979,N_9116);
nor U9997 (N_9997,N_9222,N_8920);
and U9998 (N_9998,N_9304,N_9187);
and U9999 (N_9999,N_9083,N_9230);
and U10000 (N_10000,N_9529,N_9685);
and U10001 (N_10001,N_9780,N_9583);
and U10002 (N_10002,N_9625,N_9810);
and U10003 (N_10003,N_9480,N_9944);
nand U10004 (N_10004,N_9858,N_9989);
nand U10005 (N_10005,N_9672,N_9574);
nor U10006 (N_10006,N_9702,N_9855);
and U10007 (N_10007,N_9669,N_9468);
nor U10008 (N_10008,N_9449,N_9748);
and U10009 (N_10009,N_9687,N_9700);
nand U10010 (N_10010,N_9710,N_9666);
nor U10011 (N_10011,N_9592,N_9661);
and U10012 (N_10012,N_9891,N_9376);
and U10013 (N_10013,N_9960,N_9949);
or U10014 (N_10014,N_9423,N_9504);
and U10015 (N_10015,N_9548,N_9851);
xor U10016 (N_10016,N_9857,N_9508);
and U10017 (N_10017,N_9751,N_9834);
nor U10018 (N_10018,N_9671,N_9564);
or U10019 (N_10019,N_9817,N_9405);
or U10020 (N_10020,N_9422,N_9615);
or U10021 (N_10021,N_9873,N_9448);
and U10022 (N_10022,N_9414,N_9756);
nor U10023 (N_10023,N_9708,N_9435);
or U10024 (N_10024,N_9519,N_9733);
nand U10025 (N_10025,N_9993,N_9840);
and U10026 (N_10026,N_9698,N_9550);
and U10027 (N_10027,N_9954,N_9491);
nand U10028 (N_10028,N_9838,N_9525);
xor U10029 (N_10029,N_9706,N_9815);
nand U10030 (N_10030,N_9852,N_9599);
xnor U10031 (N_10031,N_9743,N_9853);
nor U10032 (N_10032,N_9678,N_9663);
and U10033 (N_10033,N_9919,N_9938);
and U10034 (N_10034,N_9485,N_9575);
or U10035 (N_10035,N_9561,N_9772);
or U10036 (N_10036,N_9910,N_9464);
nor U10037 (N_10037,N_9498,N_9704);
xnor U10038 (N_10038,N_9439,N_9505);
nand U10039 (N_10039,N_9797,N_9579);
nand U10040 (N_10040,N_9653,N_9909);
or U10041 (N_10041,N_9454,N_9559);
or U10042 (N_10042,N_9479,N_9725);
or U10043 (N_10043,N_9676,N_9681);
or U10044 (N_10044,N_9903,N_9822);
or U10045 (N_10045,N_9682,N_9925);
xor U10046 (N_10046,N_9431,N_9864);
and U10047 (N_10047,N_9610,N_9621);
nor U10048 (N_10048,N_9406,N_9632);
or U10049 (N_10049,N_9601,N_9494);
nand U10050 (N_10050,N_9771,N_9667);
and U10051 (N_10051,N_9842,N_9399);
nand U10052 (N_10052,N_9979,N_9713);
nand U10053 (N_10053,N_9908,N_9495);
nor U10054 (N_10054,N_9729,N_9568);
or U10055 (N_10055,N_9641,N_9898);
or U10056 (N_10056,N_9546,N_9501);
and U10057 (N_10057,N_9695,N_9573);
nor U10058 (N_10058,N_9683,N_9850);
or U10059 (N_10059,N_9458,N_9869);
and U10060 (N_10060,N_9586,N_9524);
nor U10061 (N_10061,N_9897,N_9986);
and U10062 (N_10062,N_9432,N_9392);
or U10063 (N_10063,N_9389,N_9688);
nand U10064 (N_10064,N_9861,N_9745);
nand U10065 (N_10065,N_9947,N_9788);
nand U10066 (N_10066,N_9722,N_9848);
nand U10067 (N_10067,N_9488,N_9597);
nand U10068 (N_10068,N_9967,N_9400);
and U10069 (N_10069,N_9718,N_9441);
and U10070 (N_10070,N_9646,N_9930);
nor U10071 (N_10071,N_9415,N_9805);
nand U10072 (N_10072,N_9933,N_9477);
nand U10073 (N_10073,N_9746,N_9877);
nor U10074 (N_10074,N_9830,N_9383);
nor U10075 (N_10075,N_9821,N_9972);
nor U10076 (N_10076,N_9635,N_9530);
or U10077 (N_10077,N_9503,N_9499);
xnor U10078 (N_10078,N_9965,N_9553);
and U10079 (N_10079,N_9860,N_9715);
xnor U10080 (N_10080,N_9731,N_9680);
and U10081 (N_10081,N_9557,N_9964);
nor U10082 (N_10082,N_9462,N_9734);
nor U10083 (N_10083,N_9684,N_9995);
and U10084 (N_10084,N_9627,N_9447);
or U10085 (N_10085,N_9816,N_9926);
xor U10086 (N_10086,N_9460,N_9542);
and U10087 (N_10087,N_9915,N_9923);
and U10088 (N_10088,N_9461,N_9973);
nand U10089 (N_10089,N_9723,N_9711);
nor U10090 (N_10090,N_9657,N_9679);
nor U10091 (N_10091,N_9724,N_9847);
or U10092 (N_10092,N_9630,N_9781);
and U10093 (N_10093,N_9904,N_9662);
and U10094 (N_10094,N_9833,N_9963);
and U10095 (N_10095,N_9691,N_9975);
xor U10096 (N_10096,N_9803,N_9806);
or U10097 (N_10097,N_9388,N_9660);
nor U10098 (N_10098,N_9623,N_9841);
and U10099 (N_10099,N_9754,N_9878);
or U10100 (N_10100,N_9845,N_9712);
nand U10101 (N_10101,N_9379,N_9411);
nand U10102 (N_10102,N_9812,N_9612);
xnor U10103 (N_10103,N_9471,N_9570);
nand U10104 (N_10104,N_9808,N_9569);
nor U10105 (N_10105,N_9892,N_9436);
and U10106 (N_10106,N_9397,N_9478);
or U10107 (N_10107,N_9738,N_9918);
nand U10108 (N_10108,N_9976,N_9831);
and U10109 (N_10109,N_9467,N_9800);
nor U10110 (N_10110,N_9899,N_9636);
nor U10111 (N_10111,N_9577,N_9871);
and U10112 (N_10112,N_9854,N_9409);
nor U10113 (N_10113,N_9961,N_9560);
and U10114 (N_10114,N_9402,N_9759);
nor U10115 (N_10115,N_9451,N_9790);
nor U10116 (N_10116,N_9893,N_9887);
or U10117 (N_10117,N_9764,N_9894);
xnor U10118 (N_10118,N_9450,N_9533);
and U10119 (N_10119,N_9407,N_9613);
or U10120 (N_10120,N_9443,N_9554);
xor U10121 (N_10121,N_9532,N_9387);
nand U10122 (N_10122,N_9801,N_9493);
nand U10123 (N_10123,N_9928,N_9785);
nor U10124 (N_10124,N_9622,N_9496);
xnor U10125 (N_10125,N_9523,N_9673);
nor U10126 (N_10126,N_9827,N_9585);
nand U10127 (N_10127,N_9665,N_9483);
xor U10128 (N_10128,N_9728,N_9670);
or U10129 (N_10129,N_9403,N_9603);
and U10130 (N_10130,N_9658,N_9849);
nor U10131 (N_10131,N_9798,N_9437);
xnor U10132 (N_10132,N_9463,N_9936);
or U10133 (N_10133,N_9747,N_9825);
or U10134 (N_10134,N_9769,N_9652);
nor U10135 (N_10135,N_9880,N_9626);
nor U10136 (N_10136,N_9481,N_9418);
nor U10137 (N_10137,N_9521,N_9774);
nand U10138 (N_10138,N_9421,N_9526);
and U10139 (N_10139,N_9786,N_9955);
nand U10140 (N_10140,N_9633,N_9427);
nor U10141 (N_10141,N_9609,N_9582);
nand U10142 (N_10142,N_9901,N_9794);
nand U10143 (N_10143,N_9469,N_9647);
nor U10144 (N_10144,N_9590,N_9737);
and U10145 (N_10145,N_9719,N_9884);
or U10146 (N_10146,N_9643,N_9429);
nor U10147 (N_10147,N_9446,N_9377);
and U10148 (N_10148,N_9433,N_9430);
nor U10149 (N_10149,N_9921,N_9863);
nor U10150 (N_10150,N_9951,N_9907);
xor U10151 (N_10151,N_9572,N_9629);
nor U10152 (N_10152,N_9391,N_9757);
or U10153 (N_10153,N_9739,N_9958);
or U10154 (N_10154,N_9424,N_9701);
nor U10155 (N_10155,N_9466,N_9514);
or U10156 (N_10156,N_9549,N_9528);
or U10157 (N_10157,N_9924,N_9522);
nand U10158 (N_10158,N_9419,N_9656);
xnor U10159 (N_10159,N_9457,N_9992);
or U10160 (N_10160,N_9581,N_9902);
or U10161 (N_10161,N_9604,N_9645);
nor U10162 (N_10162,N_9917,N_9628);
xnor U10163 (N_10163,N_9796,N_9927);
nor U10164 (N_10164,N_9888,N_9942);
nand U10165 (N_10165,N_9906,N_9513);
and U10166 (N_10166,N_9968,N_9999);
or U10167 (N_10167,N_9616,N_9507);
nand U10168 (N_10168,N_9879,N_9882);
or U10169 (N_10169,N_9814,N_9948);
and U10170 (N_10170,N_9783,N_9937);
or U10171 (N_10171,N_9567,N_9386);
xor U10172 (N_10172,N_9982,N_9434);
or U10173 (N_10173,N_9889,N_9648);
xor U10174 (N_10174,N_9762,N_9516);
xnor U10175 (N_10175,N_9813,N_9766);
or U10176 (N_10176,N_9974,N_9594);
nand U10177 (N_10177,N_9998,N_9473);
and U10178 (N_10178,N_9922,N_9966);
nand U10179 (N_10179,N_9753,N_9375);
nand U10180 (N_10180,N_9544,N_9607);
or U10181 (N_10181,N_9872,N_9404);
nor U10182 (N_10182,N_9799,N_9789);
and U10183 (N_10183,N_9776,N_9588);
or U10184 (N_10184,N_9515,N_9792);
xnor U10185 (N_10185,N_9566,N_9939);
nor U10186 (N_10186,N_9654,N_9837);
or U10187 (N_10187,N_9941,N_9624);
nand U10188 (N_10188,N_9791,N_9677);
nor U10189 (N_10189,N_9905,N_9489);
or U10190 (N_10190,N_9959,N_9506);
and U10191 (N_10191,N_9517,N_9956);
nor U10192 (N_10192,N_9856,N_9868);
and U10193 (N_10193,N_9651,N_9482);
and U10194 (N_10194,N_9895,N_9390);
and U10195 (N_10195,N_9823,N_9824);
xnor U10196 (N_10196,N_9445,N_9385);
nand U10197 (N_10197,N_9578,N_9535);
nor U10198 (N_10198,N_9730,N_9587);
nor U10199 (N_10199,N_9401,N_9650);
and U10200 (N_10200,N_9876,N_9589);
xor U10201 (N_10201,N_9394,N_9620);
and U10202 (N_10202,N_9970,N_9608);
and U10203 (N_10203,N_9511,N_9977);
nor U10204 (N_10204,N_9758,N_9984);
nand U10205 (N_10205,N_9744,N_9770);
nand U10206 (N_10206,N_9484,N_9997);
nor U10207 (N_10207,N_9637,N_9969);
nor U10208 (N_10208,N_9735,N_9866);
and U10209 (N_10209,N_9664,N_9618);
and U10210 (N_10210,N_9846,N_9697);
and U10211 (N_10211,N_9512,N_9689);
nor U10212 (N_10212,N_9444,N_9765);
or U10213 (N_10213,N_9716,N_9865);
nor U10214 (N_10214,N_9777,N_9943);
nand U10215 (N_10215,N_9802,N_9721);
or U10216 (N_10216,N_9741,N_9520);
or U10217 (N_10217,N_9883,N_9382);
and U10218 (N_10218,N_9470,N_9487);
nor U10219 (N_10219,N_9717,N_9412);
xor U10220 (N_10220,N_9605,N_9558);
or U10221 (N_10221,N_9787,N_9552);
nand U10222 (N_10222,N_9809,N_9994);
nand U10223 (N_10223,N_9638,N_9659);
nand U10224 (N_10224,N_9900,N_9562);
nor U10225 (N_10225,N_9475,N_9571);
nor U10226 (N_10226,N_9699,N_9538);
and U10227 (N_10227,N_9752,N_9426);
and U10228 (N_10228,N_9875,N_9761);
and U10229 (N_10229,N_9991,N_9490);
or U10230 (N_10230,N_9886,N_9726);
nand U10231 (N_10231,N_9640,N_9912);
or U10232 (N_10232,N_9935,N_9606);
nand U10233 (N_10233,N_9600,N_9835);
or U10234 (N_10234,N_9536,N_9408);
nor U10235 (N_10235,N_9913,N_9619);
nor U10236 (N_10236,N_9502,N_9911);
xnor U10237 (N_10237,N_9410,N_9779);
xnor U10238 (N_10238,N_9547,N_9819);
nand U10239 (N_10239,N_9580,N_9983);
and U10240 (N_10240,N_9988,N_9413);
or U10241 (N_10241,N_9740,N_9459);
or U10242 (N_10242,N_9384,N_9393);
nand U10243 (N_10243,N_9811,N_9396);
xor U10244 (N_10244,N_9675,N_9693);
nand U10245 (N_10245,N_9844,N_9828);
or U10246 (N_10246,N_9655,N_9709);
or U10247 (N_10247,N_9438,N_9456);
or U10248 (N_10248,N_9634,N_9767);
and U10249 (N_10249,N_9420,N_9694);
and U10250 (N_10250,N_9920,N_9914);
xor U10251 (N_10251,N_9453,N_9795);
nand U10252 (N_10252,N_9820,N_9957);
nand U10253 (N_10253,N_9755,N_9707);
and U10254 (N_10254,N_9476,N_9696);
nor U10255 (N_10255,N_9642,N_9416);
nand U10256 (N_10256,N_9807,N_9596);
and U10257 (N_10257,N_9398,N_9531);
nor U10258 (N_10258,N_9953,N_9534);
and U10259 (N_10259,N_9639,N_9591);
and U10260 (N_10260,N_9563,N_9931);
nor U10261 (N_10261,N_9452,N_9425);
and U10262 (N_10262,N_9545,N_9395);
nor U10263 (N_10263,N_9946,N_9736);
or U10264 (N_10264,N_9556,N_9952);
nand U10265 (N_10265,N_9843,N_9826);
nand U10266 (N_10266,N_9782,N_9602);
xor U10267 (N_10267,N_9631,N_9978);
and U10268 (N_10268,N_9692,N_9668);
xnor U10269 (N_10269,N_9829,N_9465);
nand U10270 (N_10270,N_9551,N_9378);
nand U10271 (N_10271,N_9649,N_9742);
xor U10272 (N_10272,N_9870,N_9540);
nand U10273 (N_10273,N_9763,N_9539);
and U10274 (N_10274,N_9839,N_9760);
nand U10275 (N_10275,N_9950,N_9727);
xor U10276 (N_10276,N_9775,N_9555);
or U10277 (N_10277,N_9874,N_9380);
nor U10278 (N_10278,N_9541,N_9985);
xor U10279 (N_10279,N_9990,N_9543);
or U10280 (N_10280,N_9885,N_9862);
and U10281 (N_10281,N_9614,N_9510);
and U10282 (N_10282,N_9749,N_9674);
nand U10283 (N_10283,N_9576,N_9486);
or U10284 (N_10284,N_9934,N_9598);
xor U10285 (N_10285,N_9881,N_9455);
or U10286 (N_10286,N_9773,N_9859);
or U10287 (N_10287,N_9690,N_9440);
and U10288 (N_10288,N_9720,N_9750);
and U10289 (N_10289,N_9732,N_9644);
or U10290 (N_10290,N_9617,N_9971);
or U10291 (N_10291,N_9940,N_9593);
or U10292 (N_10292,N_9981,N_9714);
or U10293 (N_10293,N_9784,N_9987);
or U10294 (N_10294,N_9497,N_9611);
nor U10295 (N_10295,N_9472,N_9595);
nor U10296 (N_10296,N_9945,N_9381);
and U10297 (N_10297,N_9686,N_9832);
nor U10298 (N_10298,N_9996,N_9890);
nor U10299 (N_10299,N_9980,N_9428);
and U10300 (N_10300,N_9778,N_9584);
xnor U10301 (N_10301,N_9509,N_9929);
and U10302 (N_10302,N_9417,N_9818);
or U10303 (N_10303,N_9500,N_9705);
nor U10304 (N_10304,N_9836,N_9932);
and U10305 (N_10305,N_9867,N_9565);
nand U10306 (N_10306,N_9896,N_9804);
xor U10307 (N_10307,N_9537,N_9492);
nand U10308 (N_10308,N_9474,N_9442);
or U10309 (N_10309,N_9527,N_9703);
nor U10310 (N_10310,N_9518,N_9793);
and U10311 (N_10311,N_9916,N_9768);
or U10312 (N_10312,N_9962,N_9652);
xor U10313 (N_10313,N_9707,N_9956);
and U10314 (N_10314,N_9467,N_9992);
and U10315 (N_10315,N_9511,N_9514);
nor U10316 (N_10316,N_9391,N_9761);
and U10317 (N_10317,N_9410,N_9697);
nand U10318 (N_10318,N_9780,N_9980);
xor U10319 (N_10319,N_9882,N_9811);
or U10320 (N_10320,N_9938,N_9391);
or U10321 (N_10321,N_9839,N_9777);
and U10322 (N_10322,N_9409,N_9746);
or U10323 (N_10323,N_9718,N_9596);
nor U10324 (N_10324,N_9469,N_9653);
xor U10325 (N_10325,N_9602,N_9751);
nor U10326 (N_10326,N_9625,N_9462);
xnor U10327 (N_10327,N_9538,N_9560);
xnor U10328 (N_10328,N_9550,N_9943);
nand U10329 (N_10329,N_9724,N_9912);
nor U10330 (N_10330,N_9446,N_9882);
nand U10331 (N_10331,N_9428,N_9460);
or U10332 (N_10332,N_9908,N_9991);
nand U10333 (N_10333,N_9659,N_9764);
nor U10334 (N_10334,N_9504,N_9510);
nand U10335 (N_10335,N_9617,N_9709);
or U10336 (N_10336,N_9870,N_9552);
xor U10337 (N_10337,N_9449,N_9521);
and U10338 (N_10338,N_9914,N_9410);
nor U10339 (N_10339,N_9943,N_9497);
and U10340 (N_10340,N_9837,N_9375);
and U10341 (N_10341,N_9489,N_9953);
nor U10342 (N_10342,N_9749,N_9520);
and U10343 (N_10343,N_9413,N_9452);
nor U10344 (N_10344,N_9754,N_9604);
nand U10345 (N_10345,N_9692,N_9580);
nand U10346 (N_10346,N_9751,N_9562);
nand U10347 (N_10347,N_9664,N_9520);
xnor U10348 (N_10348,N_9564,N_9461);
nor U10349 (N_10349,N_9743,N_9884);
and U10350 (N_10350,N_9633,N_9789);
or U10351 (N_10351,N_9517,N_9954);
or U10352 (N_10352,N_9998,N_9846);
or U10353 (N_10353,N_9420,N_9532);
nand U10354 (N_10354,N_9796,N_9728);
nor U10355 (N_10355,N_9706,N_9619);
and U10356 (N_10356,N_9754,N_9545);
nand U10357 (N_10357,N_9654,N_9702);
nor U10358 (N_10358,N_9913,N_9723);
or U10359 (N_10359,N_9803,N_9986);
or U10360 (N_10360,N_9971,N_9475);
nor U10361 (N_10361,N_9657,N_9992);
nor U10362 (N_10362,N_9460,N_9759);
or U10363 (N_10363,N_9789,N_9384);
or U10364 (N_10364,N_9952,N_9642);
nand U10365 (N_10365,N_9506,N_9543);
nor U10366 (N_10366,N_9780,N_9505);
xnor U10367 (N_10367,N_9534,N_9768);
and U10368 (N_10368,N_9801,N_9856);
and U10369 (N_10369,N_9734,N_9532);
nand U10370 (N_10370,N_9493,N_9506);
nor U10371 (N_10371,N_9760,N_9792);
and U10372 (N_10372,N_9763,N_9541);
and U10373 (N_10373,N_9955,N_9505);
nand U10374 (N_10374,N_9409,N_9456);
xor U10375 (N_10375,N_9419,N_9986);
xnor U10376 (N_10376,N_9712,N_9699);
nand U10377 (N_10377,N_9847,N_9872);
nor U10378 (N_10378,N_9536,N_9490);
nand U10379 (N_10379,N_9819,N_9808);
and U10380 (N_10380,N_9488,N_9457);
xor U10381 (N_10381,N_9713,N_9907);
or U10382 (N_10382,N_9381,N_9605);
and U10383 (N_10383,N_9667,N_9889);
or U10384 (N_10384,N_9573,N_9660);
nor U10385 (N_10385,N_9441,N_9489);
and U10386 (N_10386,N_9727,N_9927);
and U10387 (N_10387,N_9857,N_9772);
nand U10388 (N_10388,N_9601,N_9512);
nand U10389 (N_10389,N_9739,N_9982);
or U10390 (N_10390,N_9394,N_9381);
or U10391 (N_10391,N_9406,N_9396);
nand U10392 (N_10392,N_9685,N_9936);
xnor U10393 (N_10393,N_9819,N_9811);
nand U10394 (N_10394,N_9898,N_9522);
nor U10395 (N_10395,N_9563,N_9431);
xnor U10396 (N_10396,N_9635,N_9533);
xor U10397 (N_10397,N_9382,N_9800);
nand U10398 (N_10398,N_9513,N_9860);
or U10399 (N_10399,N_9798,N_9563);
nor U10400 (N_10400,N_9644,N_9411);
nor U10401 (N_10401,N_9479,N_9636);
or U10402 (N_10402,N_9465,N_9964);
or U10403 (N_10403,N_9730,N_9418);
nor U10404 (N_10404,N_9616,N_9990);
or U10405 (N_10405,N_9857,N_9523);
or U10406 (N_10406,N_9766,N_9821);
nor U10407 (N_10407,N_9969,N_9427);
or U10408 (N_10408,N_9467,N_9836);
nand U10409 (N_10409,N_9817,N_9569);
xnor U10410 (N_10410,N_9623,N_9411);
and U10411 (N_10411,N_9686,N_9753);
xor U10412 (N_10412,N_9548,N_9521);
or U10413 (N_10413,N_9589,N_9735);
nor U10414 (N_10414,N_9899,N_9827);
and U10415 (N_10415,N_9547,N_9421);
nand U10416 (N_10416,N_9999,N_9583);
xor U10417 (N_10417,N_9619,N_9558);
nor U10418 (N_10418,N_9417,N_9725);
xnor U10419 (N_10419,N_9928,N_9649);
nor U10420 (N_10420,N_9627,N_9523);
or U10421 (N_10421,N_9520,N_9448);
or U10422 (N_10422,N_9480,N_9407);
and U10423 (N_10423,N_9805,N_9405);
nor U10424 (N_10424,N_9907,N_9973);
or U10425 (N_10425,N_9393,N_9880);
nand U10426 (N_10426,N_9742,N_9859);
nand U10427 (N_10427,N_9414,N_9550);
nor U10428 (N_10428,N_9427,N_9593);
or U10429 (N_10429,N_9658,N_9624);
xnor U10430 (N_10430,N_9829,N_9790);
nand U10431 (N_10431,N_9977,N_9935);
and U10432 (N_10432,N_9665,N_9920);
xor U10433 (N_10433,N_9398,N_9569);
nand U10434 (N_10434,N_9982,N_9485);
or U10435 (N_10435,N_9488,N_9953);
or U10436 (N_10436,N_9653,N_9652);
or U10437 (N_10437,N_9908,N_9794);
nor U10438 (N_10438,N_9553,N_9550);
nor U10439 (N_10439,N_9610,N_9581);
or U10440 (N_10440,N_9579,N_9557);
or U10441 (N_10441,N_9581,N_9964);
nor U10442 (N_10442,N_9607,N_9492);
and U10443 (N_10443,N_9949,N_9941);
nand U10444 (N_10444,N_9525,N_9593);
and U10445 (N_10445,N_9487,N_9747);
and U10446 (N_10446,N_9656,N_9765);
or U10447 (N_10447,N_9621,N_9807);
or U10448 (N_10448,N_9725,N_9702);
or U10449 (N_10449,N_9421,N_9874);
xnor U10450 (N_10450,N_9999,N_9788);
or U10451 (N_10451,N_9621,N_9710);
and U10452 (N_10452,N_9696,N_9750);
nor U10453 (N_10453,N_9603,N_9609);
or U10454 (N_10454,N_9412,N_9886);
xor U10455 (N_10455,N_9384,N_9601);
nand U10456 (N_10456,N_9767,N_9745);
nor U10457 (N_10457,N_9443,N_9407);
nor U10458 (N_10458,N_9663,N_9388);
nand U10459 (N_10459,N_9899,N_9943);
or U10460 (N_10460,N_9983,N_9393);
or U10461 (N_10461,N_9600,N_9541);
nor U10462 (N_10462,N_9778,N_9781);
nand U10463 (N_10463,N_9735,N_9858);
nor U10464 (N_10464,N_9643,N_9513);
xnor U10465 (N_10465,N_9541,N_9902);
and U10466 (N_10466,N_9743,N_9629);
nand U10467 (N_10467,N_9422,N_9850);
or U10468 (N_10468,N_9411,N_9897);
nor U10469 (N_10469,N_9829,N_9638);
xor U10470 (N_10470,N_9692,N_9610);
xor U10471 (N_10471,N_9508,N_9788);
or U10472 (N_10472,N_9721,N_9533);
or U10473 (N_10473,N_9384,N_9413);
nor U10474 (N_10474,N_9643,N_9932);
and U10475 (N_10475,N_9575,N_9629);
xnor U10476 (N_10476,N_9538,N_9517);
and U10477 (N_10477,N_9527,N_9972);
xor U10478 (N_10478,N_9550,N_9923);
and U10479 (N_10479,N_9640,N_9698);
nand U10480 (N_10480,N_9613,N_9885);
or U10481 (N_10481,N_9387,N_9996);
and U10482 (N_10482,N_9571,N_9646);
or U10483 (N_10483,N_9459,N_9478);
or U10484 (N_10484,N_9514,N_9789);
nor U10485 (N_10485,N_9667,N_9726);
nand U10486 (N_10486,N_9982,N_9863);
xor U10487 (N_10487,N_9903,N_9580);
and U10488 (N_10488,N_9615,N_9641);
and U10489 (N_10489,N_9430,N_9961);
nand U10490 (N_10490,N_9490,N_9482);
or U10491 (N_10491,N_9579,N_9551);
nand U10492 (N_10492,N_9702,N_9809);
and U10493 (N_10493,N_9923,N_9555);
or U10494 (N_10494,N_9982,N_9774);
and U10495 (N_10495,N_9406,N_9827);
and U10496 (N_10496,N_9822,N_9408);
and U10497 (N_10497,N_9492,N_9481);
or U10498 (N_10498,N_9428,N_9934);
xnor U10499 (N_10499,N_9811,N_9901);
nor U10500 (N_10500,N_9812,N_9701);
nand U10501 (N_10501,N_9685,N_9382);
nand U10502 (N_10502,N_9493,N_9912);
nor U10503 (N_10503,N_9600,N_9771);
xnor U10504 (N_10504,N_9631,N_9382);
nand U10505 (N_10505,N_9723,N_9891);
nand U10506 (N_10506,N_9635,N_9483);
nor U10507 (N_10507,N_9533,N_9784);
or U10508 (N_10508,N_9760,N_9388);
nor U10509 (N_10509,N_9452,N_9847);
nand U10510 (N_10510,N_9413,N_9573);
or U10511 (N_10511,N_9498,N_9500);
or U10512 (N_10512,N_9649,N_9701);
and U10513 (N_10513,N_9688,N_9691);
or U10514 (N_10514,N_9477,N_9672);
or U10515 (N_10515,N_9436,N_9772);
and U10516 (N_10516,N_9446,N_9832);
nand U10517 (N_10517,N_9728,N_9944);
nor U10518 (N_10518,N_9520,N_9401);
and U10519 (N_10519,N_9655,N_9479);
or U10520 (N_10520,N_9958,N_9859);
nor U10521 (N_10521,N_9511,N_9438);
or U10522 (N_10522,N_9520,N_9834);
and U10523 (N_10523,N_9775,N_9624);
and U10524 (N_10524,N_9817,N_9585);
xor U10525 (N_10525,N_9605,N_9763);
xor U10526 (N_10526,N_9730,N_9716);
or U10527 (N_10527,N_9469,N_9815);
or U10528 (N_10528,N_9952,N_9820);
and U10529 (N_10529,N_9511,N_9556);
nand U10530 (N_10530,N_9929,N_9633);
and U10531 (N_10531,N_9575,N_9498);
xor U10532 (N_10532,N_9402,N_9587);
nor U10533 (N_10533,N_9892,N_9810);
nand U10534 (N_10534,N_9748,N_9679);
nor U10535 (N_10535,N_9462,N_9419);
or U10536 (N_10536,N_9988,N_9891);
or U10537 (N_10537,N_9667,N_9624);
nor U10538 (N_10538,N_9510,N_9472);
or U10539 (N_10539,N_9620,N_9726);
nor U10540 (N_10540,N_9737,N_9478);
nand U10541 (N_10541,N_9814,N_9737);
and U10542 (N_10542,N_9757,N_9708);
and U10543 (N_10543,N_9768,N_9745);
and U10544 (N_10544,N_9820,N_9469);
nor U10545 (N_10545,N_9735,N_9476);
nand U10546 (N_10546,N_9945,N_9752);
nand U10547 (N_10547,N_9917,N_9462);
and U10548 (N_10548,N_9380,N_9650);
nor U10549 (N_10549,N_9755,N_9491);
nand U10550 (N_10550,N_9427,N_9553);
or U10551 (N_10551,N_9404,N_9997);
nor U10552 (N_10552,N_9873,N_9401);
nand U10553 (N_10553,N_9924,N_9933);
xnor U10554 (N_10554,N_9891,N_9982);
xnor U10555 (N_10555,N_9485,N_9691);
nand U10556 (N_10556,N_9381,N_9659);
nor U10557 (N_10557,N_9452,N_9897);
xnor U10558 (N_10558,N_9949,N_9987);
and U10559 (N_10559,N_9737,N_9486);
and U10560 (N_10560,N_9612,N_9779);
and U10561 (N_10561,N_9379,N_9921);
nand U10562 (N_10562,N_9972,N_9962);
and U10563 (N_10563,N_9969,N_9599);
or U10564 (N_10564,N_9451,N_9775);
or U10565 (N_10565,N_9633,N_9812);
nand U10566 (N_10566,N_9658,N_9873);
nor U10567 (N_10567,N_9836,N_9542);
and U10568 (N_10568,N_9768,N_9530);
or U10569 (N_10569,N_9511,N_9518);
and U10570 (N_10570,N_9950,N_9601);
nor U10571 (N_10571,N_9427,N_9671);
xnor U10572 (N_10572,N_9876,N_9443);
nor U10573 (N_10573,N_9378,N_9492);
xor U10574 (N_10574,N_9471,N_9941);
and U10575 (N_10575,N_9947,N_9682);
nor U10576 (N_10576,N_9901,N_9716);
xnor U10577 (N_10577,N_9873,N_9496);
or U10578 (N_10578,N_9991,N_9412);
or U10579 (N_10579,N_9384,N_9689);
or U10580 (N_10580,N_9398,N_9867);
and U10581 (N_10581,N_9679,N_9904);
nand U10582 (N_10582,N_9860,N_9382);
or U10583 (N_10583,N_9929,N_9932);
and U10584 (N_10584,N_9722,N_9779);
nor U10585 (N_10585,N_9654,N_9833);
and U10586 (N_10586,N_9482,N_9956);
nor U10587 (N_10587,N_9438,N_9682);
and U10588 (N_10588,N_9474,N_9991);
xor U10589 (N_10589,N_9719,N_9863);
and U10590 (N_10590,N_9978,N_9758);
nor U10591 (N_10591,N_9621,N_9889);
or U10592 (N_10592,N_9377,N_9894);
nand U10593 (N_10593,N_9712,N_9894);
nand U10594 (N_10594,N_9737,N_9988);
xnor U10595 (N_10595,N_9399,N_9803);
nand U10596 (N_10596,N_9892,N_9805);
nand U10597 (N_10597,N_9987,N_9772);
or U10598 (N_10598,N_9674,N_9443);
nand U10599 (N_10599,N_9761,N_9383);
nand U10600 (N_10600,N_9880,N_9877);
nand U10601 (N_10601,N_9448,N_9568);
nand U10602 (N_10602,N_9761,N_9836);
nand U10603 (N_10603,N_9785,N_9854);
nor U10604 (N_10604,N_9471,N_9748);
nor U10605 (N_10605,N_9539,N_9536);
xor U10606 (N_10606,N_9985,N_9381);
or U10607 (N_10607,N_9722,N_9951);
nand U10608 (N_10608,N_9583,N_9966);
nand U10609 (N_10609,N_9981,N_9635);
nand U10610 (N_10610,N_9798,N_9622);
and U10611 (N_10611,N_9510,N_9387);
or U10612 (N_10612,N_9573,N_9421);
nor U10613 (N_10613,N_9675,N_9626);
xnor U10614 (N_10614,N_9421,N_9454);
xor U10615 (N_10615,N_9760,N_9495);
and U10616 (N_10616,N_9524,N_9816);
nor U10617 (N_10617,N_9533,N_9432);
nor U10618 (N_10618,N_9525,N_9894);
nand U10619 (N_10619,N_9826,N_9519);
or U10620 (N_10620,N_9930,N_9987);
and U10621 (N_10621,N_9942,N_9388);
nor U10622 (N_10622,N_9420,N_9844);
or U10623 (N_10623,N_9817,N_9950);
nor U10624 (N_10624,N_9720,N_9846);
xor U10625 (N_10625,N_10569,N_10175);
nand U10626 (N_10626,N_10516,N_10238);
or U10627 (N_10627,N_10479,N_10024);
nand U10628 (N_10628,N_10139,N_10581);
nor U10629 (N_10629,N_10346,N_10452);
and U10630 (N_10630,N_10129,N_10058);
or U10631 (N_10631,N_10230,N_10324);
nor U10632 (N_10632,N_10561,N_10620);
nor U10633 (N_10633,N_10166,N_10467);
nand U10634 (N_10634,N_10353,N_10182);
and U10635 (N_10635,N_10536,N_10414);
nand U10636 (N_10636,N_10320,N_10586);
and U10637 (N_10637,N_10379,N_10174);
xnor U10638 (N_10638,N_10003,N_10065);
or U10639 (N_10639,N_10328,N_10015);
xnor U10640 (N_10640,N_10224,N_10270);
nor U10641 (N_10641,N_10053,N_10215);
or U10642 (N_10642,N_10391,N_10472);
or U10643 (N_10643,N_10564,N_10136);
or U10644 (N_10644,N_10153,N_10493);
and U10645 (N_10645,N_10432,N_10613);
nand U10646 (N_10646,N_10044,N_10462);
nor U10647 (N_10647,N_10524,N_10465);
xnor U10648 (N_10648,N_10026,N_10204);
nor U10649 (N_10649,N_10112,N_10510);
or U10650 (N_10650,N_10043,N_10411);
and U10651 (N_10651,N_10214,N_10241);
nor U10652 (N_10652,N_10508,N_10590);
nor U10653 (N_10653,N_10375,N_10016);
nand U10654 (N_10654,N_10611,N_10622);
and U10655 (N_10655,N_10056,N_10585);
and U10656 (N_10656,N_10192,N_10037);
and U10657 (N_10657,N_10009,N_10331);
or U10658 (N_10658,N_10080,N_10440);
nor U10659 (N_10659,N_10371,N_10064);
nand U10660 (N_10660,N_10595,N_10596);
or U10661 (N_10661,N_10374,N_10489);
and U10662 (N_10662,N_10228,N_10399);
nor U10663 (N_10663,N_10231,N_10504);
nand U10664 (N_10664,N_10202,N_10264);
nor U10665 (N_10665,N_10004,N_10030);
nor U10666 (N_10666,N_10351,N_10035);
and U10667 (N_10667,N_10394,N_10059);
and U10668 (N_10668,N_10071,N_10495);
or U10669 (N_10669,N_10439,N_10236);
and U10670 (N_10670,N_10535,N_10385);
and U10671 (N_10671,N_10521,N_10121);
nor U10672 (N_10672,N_10333,N_10225);
or U10673 (N_10673,N_10021,N_10617);
nor U10674 (N_10674,N_10522,N_10587);
nand U10675 (N_10675,N_10475,N_10171);
nor U10676 (N_10676,N_10213,N_10046);
nand U10677 (N_10677,N_10235,N_10575);
nand U10678 (N_10678,N_10151,N_10566);
or U10679 (N_10679,N_10459,N_10001);
nand U10680 (N_10680,N_10530,N_10081);
and U10681 (N_10681,N_10078,N_10152);
or U10682 (N_10682,N_10117,N_10261);
nand U10683 (N_10683,N_10332,N_10051);
or U10684 (N_10684,N_10477,N_10102);
and U10685 (N_10685,N_10570,N_10284);
nor U10686 (N_10686,N_10249,N_10578);
xor U10687 (N_10687,N_10050,N_10403);
and U10688 (N_10688,N_10386,N_10289);
nor U10689 (N_10689,N_10384,N_10122);
nor U10690 (N_10690,N_10589,N_10147);
or U10691 (N_10691,N_10062,N_10370);
nor U10692 (N_10692,N_10023,N_10106);
nor U10693 (N_10693,N_10594,N_10274);
nor U10694 (N_10694,N_10268,N_10551);
or U10695 (N_10695,N_10123,N_10142);
xnor U10696 (N_10696,N_10255,N_10216);
and U10697 (N_10697,N_10304,N_10098);
and U10698 (N_10698,N_10110,N_10275);
nor U10699 (N_10699,N_10156,N_10287);
nor U10700 (N_10700,N_10453,N_10031);
nand U10701 (N_10701,N_10093,N_10437);
nor U10702 (N_10702,N_10597,N_10515);
or U10703 (N_10703,N_10244,N_10203);
nand U10704 (N_10704,N_10036,N_10061);
and U10705 (N_10705,N_10278,N_10448);
xnor U10706 (N_10706,N_10464,N_10606);
nand U10707 (N_10707,N_10197,N_10226);
or U10708 (N_10708,N_10201,N_10612);
xor U10709 (N_10709,N_10257,N_10433);
or U10710 (N_10710,N_10115,N_10087);
xnor U10711 (N_10711,N_10267,N_10157);
or U10712 (N_10712,N_10045,N_10169);
or U10713 (N_10713,N_10429,N_10208);
or U10714 (N_10714,N_10577,N_10400);
xor U10715 (N_10715,N_10428,N_10588);
xor U10716 (N_10716,N_10471,N_10207);
nor U10717 (N_10717,N_10406,N_10259);
nand U10718 (N_10718,N_10438,N_10130);
or U10719 (N_10719,N_10150,N_10040);
nor U10720 (N_10720,N_10513,N_10316);
and U10721 (N_10721,N_10486,N_10181);
and U10722 (N_10722,N_10396,N_10000);
and U10723 (N_10723,N_10020,N_10014);
and U10724 (N_10724,N_10222,N_10425);
nand U10725 (N_10725,N_10246,N_10435);
xnor U10726 (N_10726,N_10105,N_10167);
and U10727 (N_10727,N_10283,N_10256);
nor U10728 (N_10728,N_10445,N_10017);
nand U10729 (N_10729,N_10481,N_10311);
and U10730 (N_10730,N_10325,N_10279);
or U10731 (N_10731,N_10184,N_10079);
nor U10732 (N_10732,N_10245,N_10434);
nor U10733 (N_10733,N_10327,N_10610);
or U10734 (N_10734,N_10473,N_10534);
nor U10735 (N_10735,N_10592,N_10041);
or U10736 (N_10736,N_10444,N_10321);
or U10737 (N_10737,N_10511,N_10178);
or U10738 (N_10738,N_10143,N_10196);
or U10739 (N_10739,N_10579,N_10373);
and U10740 (N_10740,N_10034,N_10565);
and U10741 (N_10741,N_10584,N_10544);
and U10742 (N_10742,N_10543,N_10463);
nand U10743 (N_10743,N_10159,N_10199);
nor U10744 (N_10744,N_10308,N_10146);
nand U10745 (N_10745,N_10563,N_10109);
nor U10746 (N_10746,N_10365,N_10296);
and U10747 (N_10747,N_10350,N_10126);
nor U10748 (N_10748,N_10048,N_10103);
or U10749 (N_10749,N_10312,N_10299);
nor U10750 (N_10750,N_10006,N_10125);
nor U10751 (N_10751,N_10600,N_10060);
or U10752 (N_10752,N_10421,N_10075);
nand U10753 (N_10753,N_10314,N_10148);
and U10754 (N_10754,N_10134,N_10393);
nor U10755 (N_10755,N_10198,N_10363);
xnor U10756 (N_10756,N_10357,N_10179);
and U10757 (N_10757,N_10388,N_10492);
nand U10758 (N_10758,N_10094,N_10395);
nand U10759 (N_10759,N_10605,N_10500);
and U10760 (N_10760,N_10286,N_10008);
and U10761 (N_10761,N_10621,N_10033);
or U10762 (N_10762,N_10029,N_10424);
nand U10763 (N_10763,N_10269,N_10276);
or U10764 (N_10764,N_10342,N_10319);
or U10765 (N_10765,N_10537,N_10413);
xor U10766 (N_10766,N_10392,N_10300);
and U10767 (N_10767,N_10533,N_10212);
and U10768 (N_10768,N_10624,N_10505);
nand U10769 (N_10769,N_10468,N_10458);
and U10770 (N_10770,N_10233,N_10221);
and U10771 (N_10771,N_10277,N_10329);
and U10772 (N_10772,N_10483,N_10525);
nor U10773 (N_10773,N_10366,N_10195);
nor U10774 (N_10774,N_10076,N_10054);
nand U10775 (N_10775,N_10022,N_10361);
nor U10776 (N_10776,N_10293,N_10108);
nand U10777 (N_10777,N_10084,N_10217);
or U10778 (N_10778,N_10042,N_10120);
xnor U10779 (N_10779,N_10091,N_10608);
and U10780 (N_10780,N_10191,N_10502);
nor U10781 (N_10781,N_10367,N_10019);
xnor U10782 (N_10782,N_10190,N_10252);
nor U10783 (N_10783,N_10177,N_10369);
nand U10784 (N_10784,N_10356,N_10083);
xnor U10785 (N_10785,N_10518,N_10514);
and U10786 (N_10786,N_10484,N_10262);
nand U10787 (N_10787,N_10441,N_10339);
or U10788 (N_10788,N_10598,N_10306);
or U10789 (N_10789,N_10101,N_10360);
nand U10790 (N_10790,N_10187,N_10368);
nand U10791 (N_10791,N_10422,N_10135);
and U10792 (N_10792,N_10007,N_10027);
xor U10793 (N_10793,N_10402,N_10461);
xnor U10794 (N_10794,N_10503,N_10302);
xnor U10795 (N_10795,N_10404,N_10412);
and U10796 (N_10796,N_10474,N_10086);
nand U10797 (N_10797,N_10055,N_10359);
and U10798 (N_10798,N_10457,N_10442);
nor U10799 (N_10799,N_10012,N_10280);
or U10800 (N_10800,N_10377,N_10100);
and U10801 (N_10801,N_10185,N_10431);
xnor U10802 (N_10802,N_10124,N_10310);
and U10803 (N_10803,N_10488,N_10172);
xor U10804 (N_10804,N_10128,N_10409);
nor U10805 (N_10805,N_10601,N_10025);
or U10806 (N_10806,N_10410,N_10200);
or U10807 (N_10807,N_10407,N_10193);
or U10808 (N_10808,N_10206,N_10095);
nand U10809 (N_10809,N_10160,N_10583);
nand U10810 (N_10810,N_10164,N_10313);
or U10811 (N_10811,N_10318,N_10390);
or U10812 (N_10812,N_10528,N_10451);
and U10813 (N_10813,N_10389,N_10506);
and U10814 (N_10814,N_10144,N_10419);
xnor U10815 (N_10815,N_10104,N_10573);
or U10816 (N_10816,N_10436,N_10554);
and U10817 (N_10817,N_10408,N_10116);
nand U10818 (N_10818,N_10415,N_10180);
nor U10819 (N_10819,N_10298,N_10427);
and U10820 (N_10820,N_10591,N_10540);
nand U10821 (N_10821,N_10247,N_10170);
xor U10822 (N_10822,N_10282,N_10232);
nor U10823 (N_10823,N_10599,N_10114);
or U10824 (N_10824,N_10227,N_10496);
and U10825 (N_10825,N_10345,N_10450);
or U10826 (N_10826,N_10607,N_10476);
and U10827 (N_10827,N_10265,N_10580);
or U10828 (N_10828,N_10301,N_10364);
or U10829 (N_10829,N_10501,N_10154);
or U10830 (N_10830,N_10616,N_10541);
and U10831 (N_10831,N_10548,N_10538);
xnor U10832 (N_10832,N_10049,N_10447);
xor U10833 (N_10833,N_10555,N_10138);
and U10834 (N_10834,N_10089,N_10295);
and U10835 (N_10835,N_10039,N_10571);
and U10836 (N_10836,N_10309,N_10322);
or U10837 (N_10837,N_10176,N_10290);
nor U10838 (N_10838,N_10531,N_10140);
nand U10839 (N_10839,N_10348,N_10376);
and U10840 (N_10840,N_10466,N_10099);
or U10841 (N_10841,N_10281,N_10066);
nor U10842 (N_10842,N_10420,N_10210);
and U10843 (N_10843,N_10323,N_10297);
and U10844 (N_10844,N_10085,N_10380);
xor U10845 (N_10845,N_10005,N_10082);
or U10846 (N_10846,N_10337,N_10010);
nor U10847 (N_10847,N_10512,N_10582);
nor U10848 (N_10848,N_10343,N_10494);
xnor U10849 (N_10849,N_10107,N_10341);
nand U10850 (N_10850,N_10416,N_10161);
nor U10851 (N_10851,N_10011,N_10478);
and U10852 (N_10852,N_10119,N_10335);
and U10853 (N_10853,N_10383,N_10443);
nand U10854 (N_10854,N_10326,N_10509);
nor U10855 (N_10855,N_10271,N_10545);
or U10856 (N_10856,N_10381,N_10446);
nand U10857 (N_10857,N_10547,N_10405);
nor U10858 (N_10858,N_10088,N_10307);
xnor U10859 (N_10859,N_10229,N_10552);
nand U10860 (N_10860,N_10372,N_10096);
or U10861 (N_10861,N_10338,N_10490);
nor U10862 (N_10862,N_10070,N_10189);
nand U10863 (N_10863,N_10188,N_10523);
and U10864 (N_10864,N_10194,N_10546);
and U10865 (N_10865,N_10315,N_10397);
or U10866 (N_10866,N_10572,N_10239);
nand U10867 (N_10867,N_10550,N_10334);
or U10868 (N_10868,N_10032,N_10223);
nor U10869 (N_10869,N_10568,N_10118);
or U10870 (N_10870,N_10567,N_10251);
nand U10871 (N_10871,N_10285,N_10354);
nand U10872 (N_10872,N_10173,N_10113);
nor U10873 (N_10873,N_10183,N_10340);
nor U10874 (N_10874,N_10097,N_10186);
and U10875 (N_10875,N_10219,N_10242);
nand U10876 (N_10876,N_10090,N_10382);
nand U10877 (N_10877,N_10234,N_10243);
nand U10878 (N_10878,N_10272,N_10292);
or U10879 (N_10879,N_10028,N_10344);
nand U10880 (N_10880,N_10067,N_10358);
nor U10881 (N_10881,N_10491,N_10253);
or U10882 (N_10882,N_10542,N_10254);
nor U10883 (N_10883,N_10602,N_10460);
nor U10884 (N_10884,N_10619,N_10218);
and U10885 (N_10885,N_10013,N_10291);
nand U10886 (N_10886,N_10336,N_10454);
and U10887 (N_10887,N_10347,N_10398);
and U10888 (N_10888,N_10556,N_10057);
nor U10889 (N_10889,N_10263,N_10539);
nor U10890 (N_10890,N_10387,N_10220);
nand U10891 (N_10891,N_10155,N_10073);
and U10892 (N_10892,N_10480,N_10258);
and U10893 (N_10893,N_10520,N_10482);
or U10894 (N_10894,N_10131,N_10378);
xnor U10895 (N_10895,N_10560,N_10162);
nor U10896 (N_10896,N_10052,N_10303);
nor U10897 (N_10897,N_10248,N_10426);
nor U10898 (N_10898,N_10470,N_10288);
and U10899 (N_10899,N_10266,N_10562);
nand U10900 (N_10900,N_10168,N_10092);
or U10901 (N_10901,N_10487,N_10576);
nand U10902 (N_10902,N_10352,N_10260);
or U10903 (N_10903,N_10519,N_10209);
nor U10904 (N_10904,N_10163,N_10526);
or U10905 (N_10905,N_10623,N_10559);
xnor U10906 (N_10906,N_10165,N_10132);
or U10907 (N_10907,N_10574,N_10593);
nor U10908 (N_10908,N_10240,N_10133);
nand U10909 (N_10909,N_10423,N_10469);
nor U10910 (N_10910,N_10069,N_10205);
nand U10911 (N_10911,N_10614,N_10615);
nor U10912 (N_10912,N_10330,N_10557);
nor U10913 (N_10913,N_10063,N_10517);
and U10914 (N_10914,N_10349,N_10074);
nor U10915 (N_10915,N_10507,N_10111);
nor U10916 (N_10916,N_10047,N_10529);
and U10917 (N_10917,N_10498,N_10145);
or U10918 (N_10918,N_10141,N_10355);
nand U10919 (N_10919,N_10273,N_10077);
nand U10920 (N_10920,N_10250,N_10068);
and U10921 (N_10921,N_10558,N_10149);
or U10922 (N_10922,N_10549,N_10158);
nor U10923 (N_10923,N_10485,N_10497);
and U10924 (N_10924,N_10430,N_10553);
or U10925 (N_10925,N_10317,N_10294);
or U10926 (N_10926,N_10002,N_10127);
xor U10927 (N_10927,N_10072,N_10401);
nor U10928 (N_10928,N_10449,N_10618);
and U10929 (N_10929,N_10211,N_10603);
nor U10930 (N_10930,N_10499,N_10038);
nor U10931 (N_10931,N_10362,N_10018);
nand U10932 (N_10932,N_10305,N_10456);
nor U10933 (N_10933,N_10418,N_10417);
or U10934 (N_10934,N_10609,N_10137);
xor U10935 (N_10935,N_10237,N_10527);
and U10936 (N_10936,N_10604,N_10532);
or U10937 (N_10937,N_10455,N_10599);
and U10938 (N_10938,N_10086,N_10447);
or U10939 (N_10939,N_10153,N_10233);
and U10940 (N_10940,N_10363,N_10360);
nor U10941 (N_10941,N_10203,N_10309);
nor U10942 (N_10942,N_10409,N_10568);
nor U10943 (N_10943,N_10170,N_10224);
xnor U10944 (N_10944,N_10622,N_10202);
and U10945 (N_10945,N_10195,N_10280);
or U10946 (N_10946,N_10215,N_10598);
and U10947 (N_10947,N_10506,N_10112);
or U10948 (N_10948,N_10309,N_10217);
nand U10949 (N_10949,N_10497,N_10541);
nor U10950 (N_10950,N_10359,N_10380);
nor U10951 (N_10951,N_10349,N_10229);
and U10952 (N_10952,N_10178,N_10156);
nand U10953 (N_10953,N_10577,N_10046);
or U10954 (N_10954,N_10440,N_10120);
or U10955 (N_10955,N_10408,N_10597);
nand U10956 (N_10956,N_10302,N_10615);
nand U10957 (N_10957,N_10085,N_10181);
nand U10958 (N_10958,N_10019,N_10621);
and U10959 (N_10959,N_10167,N_10039);
or U10960 (N_10960,N_10463,N_10521);
nand U10961 (N_10961,N_10492,N_10120);
or U10962 (N_10962,N_10176,N_10221);
nor U10963 (N_10963,N_10167,N_10605);
nand U10964 (N_10964,N_10125,N_10121);
and U10965 (N_10965,N_10006,N_10453);
nor U10966 (N_10966,N_10540,N_10566);
nor U10967 (N_10967,N_10075,N_10323);
xnor U10968 (N_10968,N_10393,N_10178);
or U10969 (N_10969,N_10613,N_10123);
nor U10970 (N_10970,N_10368,N_10374);
nor U10971 (N_10971,N_10270,N_10351);
and U10972 (N_10972,N_10218,N_10252);
and U10973 (N_10973,N_10075,N_10055);
nor U10974 (N_10974,N_10247,N_10443);
nor U10975 (N_10975,N_10255,N_10546);
nand U10976 (N_10976,N_10301,N_10116);
and U10977 (N_10977,N_10124,N_10035);
and U10978 (N_10978,N_10303,N_10445);
nor U10979 (N_10979,N_10485,N_10498);
nand U10980 (N_10980,N_10579,N_10498);
and U10981 (N_10981,N_10358,N_10601);
nand U10982 (N_10982,N_10203,N_10365);
nor U10983 (N_10983,N_10062,N_10136);
nand U10984 (N_10984,N_10041,N_10391);
and U10985 (N_10985,N_10038,N_10090);
nor U10986 (N_10986,N_10420,N_10452);
and U10987 (N_10987,N_10547,N_10233);
and U10988 (N_10988,N_10496,N_10422);
nor U10989 (N_10989,N_10071,N_10314);
and U10990 (N_10990,N_10260,N_10419);
nor U10991 (N_10991,N_10489,N_10456);
or U10992 (N_10992,N_10119,N_10585);
nand U10993 (N_10993,N_10492,N_10491);
nand U10994 (N_10994,N_10335,N_10377);
or U10995 (N_10995,N_10416,N_10206);
nor U10996 (N_10996,N_10217,N_10112);
or U10997 (N_10997,N_10545,N_10153);
nand U10998 (N_10998,N_10174,N_10583);
nor U10999 (N_10999,N_10495,N_10446);
nand U11000 (N_11000,N_10162,N_10308);
and U11001 (N_11001,N_10163,N_10395);
or U11002 (N_11002,N_10265,N_10335);
nand U11003 (N_11003,N_10111,N_10256);
or U11004 (N_11004,N_10033,N_10611);
nor U11005 (N_11005,N_10475,N_10225);
nand U11006 (N_11006,N_10076,N_10319);
nor U11007 (N_11007,N_10475,N_10586);
or U11008 (N_11008,N_10061,N_10283);
xor U11009 (N_11009,N_10525,N_10005);
xor U11010 (N_11010,N_10111,N_10301);
and U11011 (N_11011,N_10611,N_10009);
and U11012 (N_11012,N_10620,N_10449);
xor U11013 (N_11013,N_10503,N_10251);
and U11014 (N_11014,N_10413,N_10621);
or U11015 (N_11015,N_10354,N_10103);
and U11016 (N_11016,N_10548,N_10229);
nand U11017 (N_11017,N_10106,N_10038);
xnor U11018 (N_11018,N_10263,N_10256);
nand U11019 (N_11019,N_10394,N_10503);
and U11020 (N_11020,N_10175,N_10485);
and U11021 (N_11021,N_10200,N_10292);
or U11022 (N_11022,N_10623,N_10067);
nand U11023 (N_11023,N_10503,N_10208);
and U11024 (N_11024,N_10577,N_10090);
nand U11025 (N_11025,N_10007,N_10607);
and U11026 (N_11026,N_10075,N_10522);
nand U11027 (N_11027,N_10280,N_10461);
nor U11028 (N_11028,N_10101,N_10503);
xnor U11029 (N_11029,N_10161,N_10176);
nand U11030 (N_11030,N_10469,N_10584);
nand U11031 (N_11031,N_10028,N_10318);
nand U11032 (N_11032,N_10391,N_10387);
and U11033 (N_11033,N_10126,N_10599);
nor U11034 (N_11034,N_10363,N_10442);
and U11035 (N_11035,N_10027,N_10550);
or U11036 (N_11036,N_10474,N_10142);
and U11037 (N_11037,N_10576,N_10007);
xnor U11038 (N_11038,N_10278,N_10350);
nand U11039 (N_11039,N_10385,N_10592);
xor U11040 (N_11040,N_10371,N_10075);
nor U11041 (N_11041,N_10519,N_10557);
and U11042 (N_11042,N_10039,N_10057);
and U11043 (N_11043,N_10240,N_10590);
or U11044 (N_11044,N_10535,N_10543);
and U11045 (N_11045,N_10110,N_10420);
nor U11046 (N_11046,N_10214,N_10346);
nor U11047 (N_11047,N_10014,N_10076);
or U11048 (N_11048,N_10094,N_10352);
nor U11049 (N_11049,N_10097,N_10434);
nand U11050 (N_11050,N_10175,N_10232);
xnor U11051 (N_11051,N_10058,N_10253);
nand U11052 (N_11052,N_10108,N_10047);
nand U11053 (N_11053,N_10442,N_10008);
nand U11054 (N_11054,N_10605,N_10315);
or U11055 (N_11055,N_10504,N_10057);
or U11056 (N_11056,N_10145,N_10539);
or U11057 (N_11057,N_10019,N_10391);
nand U11058 (N_11058,N_10572,N_10093);
and U11059 (N_11059,N_10581,N_10459);
nor U11060 (N_11060,N_10533,N_10519);
nand U11061 (N_11061,N_10218,N_10163);
xnor U11062 (N_11062,N_10345,N_10034);
nor U11063 (N_11063,N_10226,N_10217);
and U11064 (N_11064,N_10305,N_10371);
nand U11065 (N_11065,N_10140,N_10230);
nor U11066 (N_11066,N_10302,N_10517);
and U11067 (N_11067,N_10442,N_10193);
nor U11068 (N_11068,N_10165,N_10535);
nor U11069 (N_11069,N_10565,N_10129);
nand U11070 (N_11070,N_10585,N_10275);
or U11071 (N_11071,N_10024,N_10617);
and U11072 (N_11072,N_10450,N_10200);
xor U11073 (N_11073,N_10079,N_10268);
nor U11074 (N_11074,N_10021,N_10580);
and U11075 (N_11075,N_10611,N_10472);
and U11076 (N_11076,N_10103,N_10373);
and U11077 (N_11077,N_10057,N_10353);
or U11078 (N_11078,N_10548,N_10219);
or U11079 (N_11079,N_10029,N_10203);
nor U11080 (N_11080,N_10280,N_10116);
nand U11081 (N_11081,N_10602,N_10243);
nor U11082 (N_11082,N_10535,N_10423);
and U11083 (N_11083,N_10561,N_10058);
nor U11084 (N_11084,N_10299,N_10551);
nor U11085 (N_11085,N_10458,N_10215);
and U11086 (N_11086,N_10151,N_10405);
nor U11087 (N_11087,N_10460,N_10410);
xor U11088 (N_11088,N_10494,N_10421);
or U11089 (N_11089,N_10504,N_10211);
nor U11090 (N_11090,N_10372,N_10277);
or U11091 (N_11091,N_10380,N_10088);
or U11092 (N_11092,N_10438,N_10049);
xnor U11093 (N_11093,N_10354,N_10477);
nand U11094 (N_11094,N_10345,N_10257);
or U11095 (N_11095,N_10467,N_10303);
or U11096 (N_11096,N_10019,N_10472);
and U11097 (N_11097,N_10554,N_10239);
or U11098 (N_11098,N_10149,N_10328);
nor U11099 (N_11099,N_10441,N_10594);
and U11100 (N_11100,N_10282,N_10295);
and U11101 (N_11101,N_10554,N_10463);
or U11102 (N_11102,N_10370,N_10035);
nand U11103 (N_11103,N_10471,N_10477);
nand U11104 (N_11104,N_10060,N_10419);
xnor U11105 (N_11105,N_10468,N_10366);
or U11106 (N_11106,N_10477,N_10016);
nor U11107 (N_11107,N_10032,N_10084);
nor U11108 (N_11108,N_10227,N_10102);
nor U11109 (N_11109,N_10590,N_10376);
nand U11110 (N_11110,N_10163,N_10015);
or U11111 (N_11111,N_10183,N_10455);
or U11112 (N_11112,N_10156,N_10140);
nand U11113 (N_11113,N_10047,N_10306);
xor U11114 (N_11114,N_10240,N_10090);
and U11115 (N_11115,N_10230,N_10483);
nor U11116 (N_11116,N_10223,N_10458);
nand U11117 (N_11117,N_10215,N_10155);
and U11118 (N_11118,N_10598,N_10305);
and U11119 (N_11119,N_10079,N_10556);
nand U11120 (N_11120,N_10391,N_10097);
or U11121 (N_11121,N_10380,N_10456);
nand U11122 (N_11122,N_10206,N_10085);
nand U11123 (N_11123,N_10238,N_10284);
or U11124 (N_11124,N_10164,N_10316);
nor U11125 (N_11125,N_10503,N_10122);
nand U11126 (N_11126,N_10093,N_10275);
and U11127 (N_11127,N_10281,N_10147);
nor U11128 (N_11128,N_10522,N_10380);
and U11129 (N_11129,N_10612,N_10220);
or U11130 (N_11130,N_10484,N_10511);
nor U11131 (N_11131,N_10127,N_10240);
or U11132 (N_11132,N_10233,N_10610);
nand U11133 (N_11133,N_10108,N_10454);
nand U11134 (N_11134,N_10101,N_10537);
nor U11135 (N_11135,N_10493,N_10328);
or U11136 (N_11136,N_10403,N_10383);
and U11137 (N_11137,N_10557,N_10595);
or U11138 (N_11138,N_10375,N_10616);
or U11139 (N_11139,N_10290,N_10362);
xnor U11140 (N_11140,N_10436,N_10479);
and U11141 (N_11141,N_10380,N_10394);
or U11142 (N_11142,N_10490,N_10548);
and U11143 (N_11143,N_10598,N_10381);
or U11144 (N_11144,N_10224,N_10197);
nand U11145 (N_11145,N_10102,N_10610);
nor U11146 (N_11146,N_10065,N_10473);
or U11147 (N_11147,N_10232,N_10365);
or U11148 (N_11148,N_10131,N_10078);
or U11149 (N_11149,N_10568,N_10470);
or U11150 (N_11150,N_10439,N_10043);
nand U11151 (N_11151,N_10356,N_10186);
nor U11152 (N_11152,N_10559,N_10377);
nand U11153 (N_11153,N_10159,N_10620);
nand U11154 (N_11154,N_10208,N_10047);
xor U11155 (N_11155,N_10145,N_10071);
nand U11156 (N_11156,N_10436,N_10138);
and U11157 (N_11157,N_10437,N_10039);
xor U11158 (N_11158,N_10463,N_10181);
nor U11159 (N_11159,N_10223,N_10231);
nor U11160 (N_11160,N_10434,N_10521);
nand U11161 (N_11161,N_10099,N_10103);
and U11162 (N_11162,N_10264,N_10112);
nor U11163 (N_11163,N_10464,N_10210);
nand U11164 (N_11164,N_10456,N_10118);
or U11165 (N_11165,N_10207,N_10182);
nand U11166 (N_11166,N_10515,N_10004);
and U11167 (N_11167,N_10494,N_10131);
nand U11168 (N_11168,N_10371,N_10171);
xor U11169 (N_11169,N_10187,N_10254);
xor U11170 (N_11170,N_10374,N_10613);
and U11171 (N_11171,N_10191,N_10119);
or U11172 (N_11172,N_10493,N_10531);
xor U11173 (N_11173,N_10189,N_10225);
nand U11174 (N_11174,N_10391,N_10213);
nor U11175 (N_11175,N_10180,N_10114);
nor U11176 (N_11176,N_10497,N_10614);
nand U11177 (N_11177,N_10265,N_10188);
or U11178 (N_11178,N_10528,N_10607);
or U11179 (N_11179,N_10031,N_10504);
or U11180 (N_11180,N_10138,N_10124);
or U11181 (N_11181,N_10517,N_10165);
xnor U11182 (N_11182,N_10602,N_10499);
or U11183 (N_11183,N_10064,N_10270);
nor U11184 (N_11184,N_10169,N_10111);
or U11185 (N_11185,N_10029,N_10570);
nand U11186 (N_11186,N_10160,N_10522);
and U11187 (N_11187,N_10368,N_10109);
or U11188 (N_11188,N_10019,N_10531);
nand U11189 (N_11189,N_10114,N_10571);
and U11190 (N_11190,N_10548,N_10335);
nand U11191 (N_11191,N_10262,N_10610);
or U11192 (N_11192,N_10459,N_10141);
nor U11193 (N_11193,N_10381,N_10094);
nand U11194 (N_11194,N_10081,N_10147);
or U11195 (N_11195,N_10064,N_10058);
and U11196 (N_11196,N_10012,N_10514);
nand U11197 (N_11197,N_10395,N_10128);
or U11198 (N_11198,N_10338,N_10213);
nor U11199 (N_11199,N_10498,N_10316);
nand U11200 (N_11200,N_10102,N_10336);
and U11201 (N_11201,N_10011,N_10144);
xor U11202 (N_11202,N_10377,N_10483);
or U11203 (N_11203,N_10624,N_10147);
and U11204 (N_11204,N_10084,N_10571);
or U11205 (N_11205,N_10290,N_10032);
and U11206 (N_11206,N_10601,N_10252);
and U11207 (N_11207,N_10358,N_10268);
nand U11208 (N_11208,N_10241,N_10425);
nor U11209 (N_11209,N_10518,N_10372);
and U11210 (N_11210,N_10390,N_10014);
nand U11211 (N_11211,N_10225,N_10038);
or U11212 (N_11212,N_10057,N_10344);
nand U11213 (N_11213,N_10098,N_10447);
nor U11214 (N_11214,N_10500,N_10340);
nand U11215 (N_11215,N_10454,N_10328);
nand U11216 (N_11216,N_10387,N_10112);
nand U11217 (N_11217,N_10541,N_10576);
nand U11218 (N_11218,N_10335,N_10346);
nor U11219 (N_11219,N_10138,N_10603);
and U11220 (N_11220,N_10132,N_10303);
nand U11221 (N_11221,N_10455,N_10423);
and U11222 (N_11222,N_10377,N_10435);
nand U11223 (N_11223,N_10323,N_10381);
and U11224 (N_11224,N_10552,N_10559);
and U11225 (N_11225,N_10147,N_10504);
nand U11226 (N_11226,N_10252,N_10276);
xor U11227 (N_11227,N_10488,N_10183);
xor U11228 (N_11228,N_10323,N_10029);
and U11229 (N_11229,N_10030,N_10024);
nor U11230 (N_11230,N_10389,N_10604);
or U11231 (N_11231,N_10462,N_10250);
nor U11232 (N_11232,N_10338,N_10525);
nand U11233 (N_11233,N_10270,N_10506);
nand U11234 (N_11234,N_10344,N_10313);
nand U11235 (N_11235,N_10402,N_10409);
nor U11236 (N_11236,N_10213,N_10327);
nor U11237 (N_11237,N_10263,N_10050);
nor U11238 (N_11238,N_10269,N_10539);
nor U11239 (N_11239,N_10532,N_10495);
and U11240 (N_11240,N_10470,N_10164);
nand U11241 (N_11241,N_10005,N_10058);
nand U11242 (N_11242,N_10194,N_10337);
nor U11243 (N_11243,N_10459,N_10137);
or U11244 (N_11244,N_10328,N_10339);
or U11245 (N_11245,N_10262,N_10401);
nor U11246 (N_11246,N_10612,N_10101);
nor U11247 (N_11247,N_10134,N_10098);
and U11248 (N_11248,N_10040,N_10288);
or U11249 (N_11249,N_10367,N_10613);
or U11250 (N_11250,N_11080,N_11159);
nor U11251 (N_11251,N_11086,N_10987);
xnor U11252 (N_11252,N_10939,N_11206);
or U11253 (N_11253,N_10967,N_11130);
xor U11254 (N_11254,N_10791,N_10677);
nand U11255 (N_11255,N_10798,N_11095);
or U11256 (N_11256,N_10644,N_10970);
nand U11257 (N_11257,N_10670,N_11032);
nor U11258 (N_11258,N_11045,N_11197);
nor U11259 (N_11259,N_10663,N_10876);
and U11260 (N_11260,N_10933,N_10897);
and U11261 (N_11261,N_10981,N_11015);
and U11262 (N_11262,N_10836,N_11220);
xnor U11263 (N_11263,N_11034,N_10942);
and U11264 (N_11264,N_11136,N_10658);
nand U11265 (N_11265,N_10999,N_11096);
and U11266 (N_11266,N_10772,N_10782);
or U11267 (N_11267,N_10764,N_11191);
xor U11268 (N_11268,N_10694,N_11066);
or U11269 (N_11269,N_10890,N_11177);
nand U11270 (N_11270,N_10880,N_10647);
or U11271 (N_11271,N_10683,N_10965);
nand U11272 (N_11272,N_10913,N_11128);
and U11273 (N_11273,N_11023,N_10918);
xor U11274 (N_11274,N_10912,N_10959);
or U11275 (N_11275,N_11214,N_11028);
nor U11276 (N_11276,N_11210,N_11043);
or U11277 (N_11277,N_11133,N_11085);
nor U11278 (N_11278,N_11005,N_11019);
nor U11279 (N_11279,N_10757,N_10727);
nand U11280 (N_11280,N_11147,N_11042);
and U11281 (N_11281,N_11030,N_11051);
and U11282 (N_11282,N_11190,N_10688);
or U11283 (N_11283,N_11169,N_10884);
and U11284 (N_11284,N_10674,N_10796);
xor U11285 (N_11285,N_11061,N_10947);
xor U11286 (N_11286,N_10927,N_10753);
or U11287 (N_11287,N_10926,N_11037);
nor U11288 (N_11288,N_10667,N_10758);
or U11289 (N_11289,N_11195,N_11004);
or U11290 (N_11290,N_10781,N_11204);
xor U11291 (N_11291,N_11074,N_10735);
nand U11292 (N_11292,N_10635,N_11044);
nand U11293 (N_11293,N_10633,N_10958);
nand U11294 (N_11294,N_10626,N_11104);
or U11295 (N_11295,N_10759,N_10669);
nand U11296 (N_11296,N_10818,N_11202);
nand U11297 (N_11297,N_10750,N_10744);
nand U11298 (N_11298,N_11065,N_10975);
nor U11299 (N_11299,N_10969,N_11137);
nor U11300 (N_11300,N_10696,N_11006);
and U11301 (N_11301,N_11231,N_10627);
or U11302 (N_11302,N_11027,N_10807);
xnor U11303 (N_11303,N_10861,N_11194);
nor U11304 (N_11304,N_10661,N_10769);
and U11305 (N_11305,N_10973,N_10976);
xnor U11306 (N_11306,N_10891,N_10954);
or U11307 (N_11307,N_11050,N_11064);
and U11308 (N_11308,N_10741,N_10808);
and U11309 (N_11309,N_10980,N_11236);
or U11310 (N_11310,N_10733,N_11154);
nand U11311 (N_11311,N_11225,N_10672);
nor U11312 (N_11312,N_11017,N_10809);
nand U11313 (N_11313,N_11033,N_11209);
or U11314 (N_11314,N_11091,N_11158);
or U11315 (N_11315,N_11014,N_10909);
or U11316 (N_11316,N_10883,N_10734);
or U11317 (N_11317,N_11180,N_11108);
nand U11318 (N_11318,N_10834,N_10638);
and U11319 (N_11319,N_10893,N_10863);
nand U11320 (N_11320,N_11162,N_11230);
and U11321 (N_11321,N_10665,N_11026);
xnor U11322 (N_11322,N_11000,N_11008);
and U11323 (N_11323,N_10774,N_10961);
nor U11324 (N_11324,N_10702,N_10841);
nor U11325 (N_11325,N_11172,N_10673);
nand U11326 (N_11326,N_10904,N_10823);
nor U11327 (N_11327,N_10820,N_11079);
and U11328 (N_11328,N_10656,N_10936);
nand U11329 (N_11329,N_10889,N_10868);
nor U11330 (N_11330,N_11122,N_10817);
xor U11331 (N_11331,N_11182,N_10697);
and U11332 (N_11332,N_10745,N_10920);
nand U11333 (N_11333,N_10625,N_10819);
nand U11334 (N_11334,N_10978,N_11148);
nand U11335 (N_11335,N_10642,N_11058);
nand U11336 (N_11336,N_10684,N_10680);
and U11337 (N_11337,N_10700,N_11179);
nor U11338 (N_11338,N_11041,N_10849);
and U11339 (N_11339,N_10873,N_10716);
and U11340 (N_11340,N_10768,N_10636);
nand U11341 (N_11341,N_10848,N_11139);
nor U11342 (N_11342,N_10941,N_10790);
nand U11343 (N_11343,N_10666,N_10832);
and U11344 (N_11344,N_10874,N_10968);
nand U11345 (N_11345,N_11078,N_10977);
and U11346 (N_11346,N_11114,N_10925);
nor U11347 (N_11347,N_10846,N_10945);
nor U11348 (N_11348,N_11208,N_11181);
or U11349 (N_11349,N_11161,N_11212);
and U11350 (N_11350,N_10655,N_10793);
and U11351 (N_11351,N_10944,N_10983);
nor U11352 (N_11352,N_10810,N_11235);
nand U11353 (N_11353,N_10915,N_11163);
nor U11354 (N_11354,N_10730,N_11121);
nand U11355 (N_11355,N_10989,N_10847);
and U11356 (N_11356,N_10997,N_10877);
nor U11357 (N_11357,N_10888,N_11056);
nor U11358 (N_11358,N_11116,N_10689);
xor U11359 (N_11359,N_10882,N_11146);
nand U11360 (N_11360,N_11092,N_10643);
and U11361 (N_11361,N_10708,N_11222);
or U11362 (N_11362,N_11036,N_10695);
nand U11363 (N_11363,N_11127,N_10984);
or U11364 (N_11364,N_10826,N_10824);
nor U11365 (N_11365,N_10776,N_11070);
xnor U11366 (N_11366,N_11089,N_10901);
xor U11367 (N_11367,N_11087,N_11048);
and U11368 (N_11368,N_10723,N_10634);
nor U11369 (N_11369,N_11010,N_10903);
nor U11370 (N_11370,N_11155,N_10726);
nand U11371 (N_11371,N_11075,N_10719);
nor U11372 (N_11372,N_11112,N_10935);
and U11373 (N_11373,N_10765,N_11141);
nand U11374 (N_11374,N_10761,N_11068);
nor U11375 (N_11375,N_11057,N_10738);
nand U11376 (N_11376,N_11219,N_10922);
nor U11377 (N_11377,N_10871,N_10825);
nor U11378 (N_11378,N_11203,N_10827);
nand U11379 (N_11379,N_11072,N_10844);
nor U11380 (N_11380,N_10657,N_10713);
or U11381 (N_11381,N_10923,N_11184);
and U11382 (N_11382,N_10906,N_11012);
nand U11383 (N_11383,N_11189,N_11054);
xnor U11384 (N_11384,N_11076,N_10870);
or U11385 (N_11385,N_11152,N_10664);
xnor U11386 (N_11386,N_10654,N_10682);
nor U11387 (N_11387,N_11150,N_10845);
nand U11388 (N_11388,N_11103,N_11186);
nor U11389 (N_11389,N_10932,N_11031);
or U11390 (N_11390,N_10878,N_11242);
and U11391 (N_11391,N_11187,N_11113);
nand U11392 (N_11392,N_11107,N_11165);
or U11393 (N_11393,N_10993,N_10875);
or U11394 (N_11394,N_10681,N_10632);
nor U11395 (N_11395,N_10899,N_11249);
nand U11396 (N_11396,N_10930,N_10749);
nor U11397 (N_11397,N_10950,N_10948);
and U11398 (N_11398,N_10706,N_10957);
and U11399 (N_11399,N_11025,N_10739);
and U11400 (N_11400,N_10966,N_11047);
nor U11401 (N_11401,N_10924,N_10946);
nor U11402 (N_11402,N_11218,N_10815);
or U11403 (N_11403,N_10857,N_11109);
nand U11404 (N_11404,N_10707,N_10865);
or U11405 (N_11405,N_11247,N_11105);
and U11406 (N_11406,N_10979,N_10699);
nor U11407 (N_11407,N_11088,N_10885);
and U11408 (N_11408,N_10686,N_11125);
nand U11409 (N_11409,N_11098,N_10703);
and U11410 (N_11410,N_11016,N_11223);
nor U11411 (N_11411,N_11248,N_10971);
nor U11412 (N_11412,N_10928,N_10653);
xor U11413 (N_11413,N_11166,N_10755);
nor U11414 (N_11414,N_11175,N_10770);
xor U11415 (N_11415,N_10717,N_10676);
nand U11416 (N_11416,N_10675,N_11062);
nand U11417 (N_11417,N_10692,N_11160);
or U11418 (N_11418,N_10828,N_10860);
nand U11419 (N_11419,N_10710,N_10729);
nor U11420 (N_11420,N_10640,N_11002);
or U11421 (N_11421,N_10974,N_11233);
nor U11422 (N_11422,N_11221,N_10900);
or U11423 (N_11423,N_10990,N_11007);
and U11424 (N_11424,N_10872,N_11021);
xor U11425 (N_11425,N_11193,N_11196);
nand U11426 (N_11426,N_10646,N_10982);
nor U11427 (N_11427,N_10940,N_10917);
nand U11428 (N_11428,N_10802,N_10775);
nand U11429 (N_11429,N_11153,N_10754);
and U11430 (N_11430,N_10631,N_11035);
nor U11431 (N_11431,N_10964,N_10822);
nor U11432 (N_11432,N_10869,N_11207);
or U11433 (N_11433,N_10756,N_10721);
xor U11434 (N_11434,N_10972,N_11001);
xnor U11435 (N_11435,N_10691,N_10859);
nor U11436 (N_11436,N_10777,N_10678);
and U11437 (N_11437,N_11145,N_11063);
nand U11438 (N_11438,N_11238,N_10910);
or U11439 (N_11439,N_11123,N_11240);
and U11440 (N_11440,N_10685,N_11111);
or U11441 (N_11441,N_10816,N_10722);
nand U11442 (N_11442,N_11084,N_10783);
or U11443 (N_11443,N_11135,N_10985);
nand U11444 (N_11444,N_10839,N_10795);
and U11445 (N_11445,N_10714,N_10931);
nand U11446 (N_11446,N_10712,N_10902);
or U11447 (N_11447,N_10830,N_10831);
nor U11448 (N_11448,N_10780,N_10850);
or U11449 (N_11449,N_11183,N_11241);
or U11450 (N_11450,N_10854,N_10881);
or U11451 (N_11451,N_11011,N_10701);
nor U11452 (N_11452,N_10956,N_11093);
nand U11453 (N_11453,N_11126,N_10760);
or U11454 (N_11454,N_10651,N_10806);
nand U11455 (N_11455,N_11022,N_11059);
and U11456 (N_11456,N_10914,N_11120);
nand U11457 (N_11457,N_10679,N_10879);
nor U11458 (N_11458,N_10892,N_10938);
and U11459 (N_11459,N_10737,N_10693);
nor U11460 (N_11460,N_10934,N_10766);
nor U11461 (N_11461,N_11174,N_10650);
nand U11462 (N_11462,N_10840,N_10887);
nand U11463 (N_11463,N_10929,N_11178);
nand U11464 (N_11464,N_10814,N_10728);
or U11465 (N_11465,N_10786,N_11060);
nand U11466 (N_11466,N_10629,N_11156);
and U11467 (N_11467,N_11213,N_11020);
nand U11468 (N_11468,N_11102,N_10898);
xor U11469 (N_11469,N_11046,N_10645);
and U11470 (N_11470,N_11167,N_10953);
and U11471 (N_11471,N_10630,N_10718);
nand U11472 (N_11472,N_10704,N_10963);
nand U11473 (N_11473,N_10799,N_10751);
nor U11474 (N_11474,N_11211,N_11185);
nand U11475 (N_11475,N_11118,N_10812);
and U11476 (N_11476,N_11227,N_10852);
and U11477 (N_11477,N_10762,N_11201);
xnor U11478 (N_11478,N_11115,N_11049);
or U11479 (N_11479,N_11040,N_10800);
and U11480 (N_11480,N_10628,N_10855);
or U11481 (N_11481,N_10687,N_10867);
xnor U11482 (N_11482,N_11229,N_10952);
xor U11483 (N_11483,N_11149,N_10778);
nor U11484 (N_11484,N_11038,N_11164);
and U11485 (N_11485,N_11244,N_11140);
nor U11486 (N_11486,N_11232,N_11168);
nand U11487 (N_11487,N_11117,N_11101);
nand U11488 (N_11488,N_10955,N_10988);
or U11489 (N_11489,N_10767,N_10905);
or U11490 (N_11490,N_10911,N_11237);
nor U11491 (N_11491,N_11055,N_11003);
nor U11492 (N_11492,N_10787,N_10851);
xor U11493 (N_11493,N_10732,N_11053);
nor U11494 (N_11494,N_11205,N_10736);
and U11495 (N_11495,N_10837,N_10864);
nor U11496 (N_11496,N_11069,N_10907);
or U11497 (N_11497,N_11246,N_11082);
or U11498 (N_11498,N_10801,N_11029);
or U11499 (N_11499,N_11110,N_10835);
and U11500 (N_11500,N_10919,N_10838);
or U11501 (N_11501,N_10937,N_11217);
or U11502 (N_11502,N_10949,N_11099);
xor U11503 (N_11503,N_11067,N_10842);
nor U11504 (N_11504,N_11124,N_11157);
xnor U11505 (N_11505,N_10856,N_10784);
or U11506 (N_11506,N_11018,N_10803);
and U11507 (N_11507,N_10804,N_10794);
or U11508 (N_11508,N_11199,N_10752);
or U11509 (N_11509,N_10731,N_10715);
and U11510 (N_11510,N_10996,N_11009);
and U11511 (N_11511,N_10998,N_11097);
nor U11512 (N_11512,N_11245,N_10962);
nand U11513 (N_11513,N_10671,N_10921);
and U11514 (N_11514,N_10858,N_10639);
nor U11515 (N_11515,N_11173,N_10811);
nand U11516 (N_11516,N_10690,N_11132);
and U11517 (N_11517,N_10709,N_10763);
xor U11518 (N_11518,N_10652,N_11171);
and U11519 (N_11519,N_10821,N_10705);
xor U11520 (N_11520,N_11119,N_10843);
nor U11521 (N_11521,N_11077,N_10813);
xor U11522 (N_11522,N_11243,N_10637);
and U11523 (N_11523,N_10742,N_11081);
nand U11524 (N_11524,N_11094,N_10668);
and U11525 (N_11525,N_11013,N_10785);
xnor U11526 (N_11526,N_10805,N_10894);
xnor U11527 (N_11527,N_11024,N_10833);
xor U11528 (N_11528,N_10725,N_11134);
nor U11529 (N_11529,N_10829,N_10746);
nand U11530 (N_11530,N_11188,N_11039);
nand U11531 (N_11531,N_11073,N_10797);
nor U11532 (N_11532,N_11216,N_10743);
and U11533 (N_11533,N_11143,N_11226);
and U11534 (N_11534,N_10748,N_11144);
xnor U11535 (N_11535,N_11151,N_10711);
nand U11536 (N_11536,N_11234,N_10853);
or U11537 (N_11537,N_11200,N_11198);
or U11538 (N_11538,N_11170,N_11142);
and U11539 (N_11539,N_11192,N_10951);
nand U11540 (N_11540,N_10771,N_11215);
nor U11541 (N_11541,N_11071,N_10641);
nand U11542 (N_11542,N_10788,N_10659);
nor U11543 (N_11543,N_10943,N_10649);
nor U11544 (N_11544,N_11090,N_10995);
nand U11545 (N_11545,N_10886,N_10773);
xor U11546 (N_11546,N_11083,N_10698);
nand U11547 (N_11547,N_10991,N_11176);
nand U11548 (N_11548,N_10740,N_11052);
nor U11549 (N_11549,N_10994,N_11224);
xor U11550 (N_11550,N_10862,N_10792);
or U11551 (N_11551,N_11239,N_10986);
xnor U11552 (N_11552,N_10648,N_10908);
nor U11553 (N_11553,N_10662,N_11106);
nand U11554 (N_11554,N_10916,N_10789);
nor U11555 (N_11555,N_10724,N_10660);
or U11556 (N_11556,N_11131,N_11228);
nand U11557 (N_11557,N_10779,N_11100);
nand U11558 (N_11558,N_10895,N_11138);
nand U11559 (N_11559,N_11129,N_10960);
nand U11560 (N_11560,N_10720,N_10747);
nor U11561 (N_11561,N_10992,N_10866);
and U11562 (N_11562,N_10896,N_11243);
xor U11563 (N_11563,N_10862,N_10999);
nor U11564 (N_11564,N_11204,N_10844);
or U11565 (N_11565,N_11124,N_10656);
and U11566 (N_11566,N_10942,N_11127);
and U11567 (N_11567,N_10894,N_11006);
nand U11568 (N_11568,N_11213,N_10675);
or U11569 (N_11569,N_11023,N_10829);
and U11570 (N_11570,N_11113,N_11226);
nand U11571 (N_11571,N_11137,N_11208);
xnor U11572 (N_11572,N_10985,N_10958);
xnor U11573 (N_11573,N_10882,N_10872);
nand U11574 (N_11574,N_11167,N_10794);
nor U11575 (N_11575,N_10954,N_10829);
and U11576 (N_11576,N_11206,N_10630);
nand U11577 (N_11577,N_11181,N_10917);
or U11578 (N_11578,N_10836,N_11203);
xor U11579 (N_11579,N_10825,N_10782);
nor U11580 (N_11580,N_10751,N_11096);
nor U11581 (N_11581,N_10770,N_11142);
nand U11582 (N_11582,N_10753,N_10894);
xor U11583 (N_11583,N_10826,N_10989);
nor U11584 (N_11584,N_10829,N_11127);
xor U11585 (N_11585,N_11024,N_10885);
and U11586 (N_11586,N_10920,N_11159);
or U11587 (N_11587,N_10646,N_10660);
or U11588 (N_11588,N_10710,N_10725);
and U11589 (N_11589,N_10700,N_10628);
xor U11590 (N_11590,N_10783,N_10931);
xnor U11591 (N_11591,N_11157,N_11061);
nor U11592 (N_11592,N_10988,N_11129);
and U11593 (N_11593,N_11213,N_10978);
nand U11594 (N_11594,N_11235,N_10780);
or U11595 (N_11595,N_10642,N_11074);
or U11596 (N_11596,N_10781,N_10722);
or U11597 (N_11597,N_10709,N_10916);
nand U11598 (N_11598,N_11175,N_11219);
or U11599 (N_11599,N_10992,N_10657);
or U11600 (N_11600,N_10754,N_11240);
xnor U11601 (N_11601,N_11242,N_11201);
or U11602 (N_11602,N_10862,N_10852);
and U11603 (N_11603,N_10827,N_11118);
or U11604 (N_11604,N_11141,N_10820);
or U11605 (N_11605,N_10721,N_10973);
or U11606 (N_11606,N_10706,N_10920);
nand U11607 (N_11607,N_11083,N_10757);
nor U11608 (N_11608,N_11164,N_10941);
and U11609 (N_11609,N_11233,N_10864);
or U11610 (N_11610,N_11128,N_10825);
and U11611 (N_11611,N_11206,N_11248);
nand U11612 (N_11612,N_10794,N_10934);
nor U11613 (N_11613,N_10642,N_11211);
and U11614 (N_11614,N_11236,N_10712);
or U11615 (N_11615,N_10960,N_10847);
or U11616 (N_11616,N_11143,N_11232);
nand U11617 (N_11617,N_10680,N_10989);
or U11618 (N_11618,N_10739,N_10876);
nor U11619 (N_11619,N_11033,N_10688);
and U11620 (N_11620,N_11181,N_11116);
xor U11621 (N_11621,N_11111,N_11186);
and U11622 (N_11622,N_11144,N_10887);
xor U11623 (N_11623,N_10777,N_11033);
and U11624 (N_11624,N_11098,N_10770);
and U11625 (N_11625,N_11143,N_10725);
nor U11626 (N_11626,N_10988,N_10786);
and U11627 (N_11627,N_10697,N_11027);
xnor U11628 (N_11628,N_10677,N_10946);
nor U11629 (N_11629,N_11108,N_11243);
nand U11630 (N_11630,N_10910,N_10708);
nand U11631 (N_11631,N_10739,N_10930);
nor U11632 (N_11632,N_11232,N_10863);
or U11633 (N_11633,N_10783,N_10920);
nand U11634 (N_11634,N_10870,N_10635);
or U11635 (N_11635,N_11170,N_11040);
nor U11636 (N_11636,N_10719,N_11105);
or U11637 (N_11637,N_10869,N_10802);
xor U11638 (N_11638,N_11036,N_11199);
nand U11639 (N_11639,N_10841,N_11118);
and U11640 (N_11640,N_10637,N_10772);
nand U11641 (N_11641,N_11045,N_10988);
and U11642 (N_11642,N_10869,N_10879);
and U11643 (N_11643,N_11189,N_10992);
nor U11644 (N_11644,N_10815,N_10767);
xor U11645 (N_11645,N_11217,N_10941);
nand U11646 (N_11646,N_10888,N_10880);
or U11647 (N_11647,N_11018,N_11228);
nor U11648 (N_11648,N_11136,N_10899);
nor U11649 (N_11649,N_11024,N_10628);
nand U11650 (N_11650,N_10679,N_11176);
xor U11651 (N_11651,N_11163,N_11154);
nand U11652 (N_11652,N_11230,N_11018);
and U11653 (N_11653,N_10693,N_11200);
xor U11654 (N_11654,N_11103,N_10737);
nor U11655 (N_11655,N_10633,N_11122);
or U11656 (N_11656,N_10730,N_10684);
and U11657 (N_11657,N_11226,N_10707);
and U11658 (N_11658,N_11151,N_11188);
and U11659 (N_11659,N_11141,N_10755);
nor U11660 (N_11660,N_10646,N_11000);
nor U11661 (N_11661,N_10893,N_10788);
or U11662 (N_11662,N_11130,N_11096);
nor U11663 (N_11663,N_10789,N_11186);
xnor U11664 (N_11664,N_10955,N_10634);
nand U11665 (N_11665,N_11045,N_11186);
and U11666 (N_11666,N_11214,N_11050);
and U11667 (N_11667,N_11031,N_11157);
nand U11668 (N_11668,N_10957,N_11167);
nand U11669 (N_11669,N_10944,N_10762);
or U11670 (N_11670,N_11238,N_10816);
nand U11671 (N_11671,N_11172,N_10997);
and U11672 (N_11672,N_10694,N_11120);
and U11673 (N_11673,N_10971,N_10826);
nor U11674 (N_11674,N_10800,N_10784);
nand U11675 (N_11675,N_10989,N_10648);
or U11676 (N_11676,N_10660,N_11091);
nand U11677 (N_11677,N_10655,N_11050);
nand U11678 (N_11678,N_10960,N_11020);
xor U11679 (N_11679,N_10630,N_10952);
nand U11680 (N_11680,N_10888,N_10839);
or U11681 (N_11681,N_11052,N_11196);
or U11682 (N_11682,N_10967,N_11117);
or U11683 (N_11683,N_10910,N_11181);
and U11684 (N_11684,N_11174,N_10802);
and U11685 (N_11685,N_10822,N_10848);
or U11686 (N_11686,N_10640,N_11131);
nand U11687 (N_11687,N_10866,N_11057);
and U11688 (N_11688,N_11183,N_10798);
xnor U11689 (N_11689,N_11093,N_11072);
nor U11690 (N_11690,N_10730,N_11197);
nand U11691 (N_11691,N_10707,N_11203);
and U11692 (N_11692,N_11046,N_10708);
or U11693 (N_11693,N_10666,N_10926);
xor U11694 (N_11694,N_10919,N_10763);
nand U11695 (N_11695,N_10693,N_10799);
nand U11696 (N_11696,N_11094,N_11038);
or U11697 (N_11697,N_11231,N_10998);
and U11698 (N_11698,N_10693,N_11236);
nand U11699 (N_11699,N_10984,N_11202);
or U11700 (N_11700,N_11159,N_10762);
and U11701 (N_11701,N_10900,N_11006);
nand U11702 (N_11702,N_11168,N_11239);
or U11703 (N_11703,N_10811,N_10858);
and U11704 (N_11704,N_10876,N_11045);
nor U11705 (N_11705,N_11066,N_10950);
xor U11706 (N_11706,N_10755,N_10847);
or U11707 (N_11707,N_11226,N_11146);
nor U11708 (N_11708,N_10756,N_11225);
nand U11709 (N_11709,N_11145,N_11147);
and U11710 (N_11710,N_11129,N_10684);
and U11711 (N_11711,N_11120,N_10880);
nor U11712 (N_11712,N_10869,N_10631);
and U11713 (N_11713,N_10729,N_10751);
or U11714 (N_11714,N_10746,N_10952);
and U11715 (N_11715,N_11047,N_11194);
and U11716 (N_11716,N_10765,N_10776);
nand U11717 (N_11717,N_10883,N_11094);
or U11718 (N_11718,N_10924,N_10781);
nor U11719 (N_11719,N_11176,N_11137);
nor U11720 (N_11720,N_11215,N_11152);
nor U11721 (N_11721,N_11025,N_11204);
and U11722 (N_11722,N_11026,N_11092);
xor U11723 (N_11723,N_11218,N_10791);
nand U11724 (N_11724,N_11194,N_10645);
nand U11725 (N_11725,N_11109,N_10753);
or U11726 (N_11726,N_11100,N_10973);
or U11727 (N_11727,N_10787,N_10706);
nor U11728 (N_11728,N_11161,N_10885);
and U11729 (N_11729,N_11107,N_10946);
xor U11730 (N_11730,N_11201,N_10721);
and U11731 (N_11731,N_10649,N_10627);
nor U11732 (N_11732,N_10731,N_10784);
or U11733 (N_11733,N_11096,N_10719);
or U11734 (N_11734,N_10922,N_11150);
nand U11735 (N_11735,N_10870,N_11128);
nand U11736 (N_11736,N_11095,N_11088);
and U11737 (N_11737,N_11151,N_10724);
nand U11738 (N_11738,N_10798,N_11191);
xnor U11739 (N_11739,N_10635,N_11228);
and U11740 (N_11740,N_11222,N_11163);
nor U11741 (N_11741,N_11160,N_11201);
and U11742 (N_11742,N_10638,N_11172);
nand U11743 (N_11743,N_10855,N_11032);
nor U11744 (N_11744,N_10950,N_10723);
nor U11745 (N_11745,N_11060,N_10958);
xor U11746 (N_11746,N_10850,N_11004);
or U11747 (N_11747,N_10868,N_10939);
xnor U11748 (N_11748,N_10686,N_11140);
nor U11749 (N_11749,N_10727,N_10703);
and U11750 (N_11750,N_10948,N_11196);
nand U11751 (N_11751,N_10941,N_11135);
and U11752 (N_11752,N_11169,N_10640);
xor U11753 (N_11753,N_11236,N_10724);
nor U11754 (N_11754,N_11201,N_10988);
and U11755 (N_11755,N_11031,N_11177);
nand U11756 (N_11756,N_10728,N_10856);
nor U11757 (N_11757,N_10860,N_10811);
nand U11758 (N_11758,N_10641,N_11125);
nand U11759 (N_11759,N_10931,N_10879);
or U11760 (N_11760,N_11051,N_10916);
nand U11761 (N_11761,N_11023,N_10874);
nand U11762 (N_11762,N_10956,N_10769);
xnor U11763 (N_11763,N_11067,N_10921);
and U11764 (N_11764,N_11123,N_10775);
nor U11765 (N_11765,N_11004,N_10935);
nand U11766 (N_11766,N_10672,N_10691);
and U11767 (N_11767,N_10700,N_11036);
and U11768 (N_11768,N_10661,N_10838);
nor U11769 (N_11769,N_10984,N_11135);
or U11770 (N_11770,N_11150,N_10770);
and U11771 (N_11771,N_11127,N_10704);
or U11772 (N_11772,N_10636,N_10786);
nand U11773 (N_11773,N_10633,N_11227);
nor U11774 (N_11774,N_11210,N_10751);
and U11775 (N_11775,N_10919,N_10718);
and U11776 (N_11776,N_11023,N_10933);
nand U11777 (N_11777,N_10865,N_10641);
nand U11778 (N_11778,N_10904,N_11116);
nor U11779 (N_11779,N_10675,N_10932);
or U11780 (N_11780,N_11167,N_10993);
nor U11781 (N_11781,N_11054,N_10894);
nor U11782 (N_11782,N_10850,N_10981);
nor U11783 (N_11783,N_11075,N_10678);
nor U11784 (N_11784,N_11008,N_11047);
nor U11785 (N_11785,N_10658,N_10815);
or U11786 (N_11786,N_11240,N_11100);
nand U11787 (N_11787,N_10642,N_11198);
nand U11788 (N_11788,N_11179,N_11058);
and U11789 (N_11789,N_11062,N_10716);
nor U11790 (N_11790,N_10827,N_10651);
or U11791 (N_11791,N_10874,N_10938);
and U11792 (N_11792,N_11226,N_10738);
xnor U11793 (N_11793,N_10991,N_11111);
nand U11794 (N_11794,N_10636,N_10687);
nor U11795 (N_11795,N_10627,N_10847);
nand U11796 (N_11796,N_10657,N_11077);
or U11797 (N_11797,N_11039,N_11154);
or U11798 (N_11798,N_10961,N_10978);
nand U11799 (N_11799,N_10969,N_10904);
and U11800 (N_11800,N_10874,N_10948);
nand U11801 (N_11801,N_11069,N_10675);
or U11802 (N_11802,N_10808,N_10626);
or U11803 (N_11803,N_10694,N_11103);
nor U11804 (N_11804,N_10805,N_10727);
or U11805 (N_11805,N_10772,N_11188);
nor U11806 (N_11806,N_11052,N_11117);
and U11807 (N_11807,N_10756,N_11118);
nand U11808 (N_11808,N_10667,N_10707);
nand U11809 (N_11809,N_10979,N_11066);
nand U11810 (N_11810,N_10805,N_11128);
nor U11811 (N_11811,N_10975,N_11219);
nor U11812 (N_11812,N_10898,N_11039);
nor U11813 (N_11813,N_10731,N_11235);
or U11814 (N_11814,N_10641,N_11066);
or U11815 (N_11815,N_11137,N_11188);
and U11816 (N_11816,N_11136,N_11110);
nand U11817 (N_11817,N_11221,N_10780);
and U11818 (N_11818,N_11072,N_11223);
nor U11819 (N_11819,N_10894,N_10682);
or U11820 (N_11820,N_10852,N_10973);
and U11821 (N_11821,N_11050,N_10883);
or U11822 (N_11822,N_10640,N_11027);
nor U11823 (N_11823,N_10641,N_10772);
xor U11824 (N_11824,N_10741,N_10782);
nand U11825 (N_11825,N_10708,N_10908);
nor U11826 (N_11826,N_11141,N_11215);
or U11827 (N_11827,N_11249,N_11042);
nor U11828 (N_11828,N_10656,N_11013);
nor U11829 (N_11829,N_10845,N_10653);
nor U11830 (N_11830,N_10714,N_10818);
or U11831 (N_11831,N_10724,N_10792);
xor U11832 (N_11832,N_10806,N_10690);
nand U11833 (N_11833,N_10908,N_11064);
or U11834 (N_11834,N_11008,N_11233);
and U11835 (N_11835,N_10919,N_10836);
or U11836 (N_11836,N_10923,N_11201);
nand U11837 (N_11837,N_10642,N_11066);
nor U11838 (N_11838,N_11204,N_10829);
or U11839 (N_11839,N_10994,N_11025);
xnor U11840 (N_11840,N_10853,N_10977);
nand U11841 (N_11841,N_10679,N_10638);
and U11842 (N_11842,N_11163,N_10879);
and U11843 (N_11843,N_10739,N_10685);
and U11844 (N_11844,N_11248,N_10744);
and U11845 (N_11845,N_10702,N_11145);
and U11846 (N_11846,N_11208,N_10912);
xor U11847 (N_11847,N_10999,N_11166);
nor U11848 (N_11848,N_11035,N_10857);
nor U11849 (N_11849,N_11057,N_10917);
nand U11850 (N_11850,N_10847,N_10698);
nand U11851 (N_11851,N_10835,N_10919);
nor U11852 (N_11852,N_10961,N_11031);
and U11853 (N_11853,N_10961,N_10673);
nand U11854 (N_11854,N_11109,N_11154);
nand U11855 (N_11855,N_10983,N_10727);
xor U11856 (N_11856,N_10681,N_10933);
xnor U11857 (N_11857,N_11243,N_11080);
nor U11858 (N_11858,N_10773,N_10687);
nor U11859 (N_11859,N_11048,N_11024);
or U11860 (N_11860,N_11232,N_10907);
and U11861 (N_11861,N_11018,N_10707);
or U11862 (N_11862,N_11130,N_11127);
nand U11863 (N_11863,N_10666,N_10875);
nand U11864 (N_11864,N_11069,N_11131);
nand U11865 (N_11865,N_10747,N_10691);
nand U11866 (N_11866,N_11230,N_10932);
nor U11867 (N_11867,N_11138,N_11038);
or U11868 (N_11868,N_10704,N_11084);
nor U11869 (N_11869,N_10646,N_10814);
nand U11870 (N_11870,N_10745,N_11145);
nand U11871 (N_11871,N_11198,N_11178);
or U11872 (N_11872,N_11148,N_11064);
nand U11873 (N_11873,N_11006,N_10867);
nand U11874 (N_11874,N_11077,N_11032);
and U11875 (N_11875,N_11277,N_11664);
and U11876 (N_11876,N_11324,N_11697);
xnor U11877 (N_11877,N_11714,N_11653);
nand U11878 (N_11878,N_11650,N_11546);
or U11879 (N_11879,N_11423,N_11281);
nor U11880 (N_11880,N_11402,N_11547);
nand U11881 (N_11881,N_11731,N_11774);
nand U11882 (N_11882,N_11723,N_11303);
and U11883 (N_11883,N_11317,N_11472);
and U11884 (N_11884,N_11651,N_11390);
or U11885 (N_11885,N_11506,N_11765);
nor U11886 (N_11886,N_11291,N_11753);
nand U11887 (N_11887,N_11795,N_11749);
nand U11888 (N_11888,N_11386,N_11777);
nand U11889 (N_11889,N_11853,N_11412);
and U11890 (N_11890,N_11453,N_11449);
xnor U11891 (N_11891,N_11778,N_11310);
and U11892 (N_11892,N_11670,N_11789);
nand U11893 (N_11893,N_11262,N_11334);
or U11894 (N_11894,N_11866,N_11603);
and U11895 (N_11895,N_11786,N_11422);
nand U11896 (N_11896,N_11411,N_11759);
xor U11897 (N_11897,N_11814,N_11843);
or U11898 (N_11898,N_11829,N_11838);
and U11899 (N_11899,N_11288,N_11632);
or U11900 (N_11900,N_11683,N_11699);
nor U11901 (N_11901,N_11286,N_11859);
nor U11902 (N_11902,N_11691,N_11542);
xnor U11903 (N_11903,N_11461,N_11358);
and U11904 (N_11904,N_11393,N_11710);
nand U11905 (N_11905,N_11821,N_11473);
nor U11906 (N_11906,N_11620,N_11576);
nor U11907 (N_11907,N_11515,N_11308);
nand U11908 (N_11908,N_11381,N_11490);
nand U11909 (N_11909,N_11374,N_11611);
or U11910 (N_11910,N_11595,N_11823);
nand U11911 (N_11911,N_11637,N_11251);
or U11912 (N_11912,N_11503,N_11619);
nor U11913 (N_11913,N_11689,N_11478);
and U11914 (N_11914,N_11252,N_11445);
or U11915 (N_11915,N_11690,N_11351);
nor U11916 (N_11916,N_11475,N_11533);
or U11917 (N_11917,N_11356,N_11682);
nor U11918 (N_11918,N_11497,N_11278);
nand U11919 (N_11919,N_11600,N_11773);
nor U11920 (N_11920,N_11638,N_11842);
and U11921 (N_11921,N_11874,N_11631);
nand U11922 (N_11922,N_11250,N_11703);
and U11923 (N_11923,N_11741,N_11819);
nor U11924 (N_11924,N_11695,N_11345);
nand U11925 (N_11925,N_11323,N_11815);
nand U11926 (N_11926,N_11481,N_11387);
and U11927 (N_11927,N_11719,N_11809);
nand U11928 (N_11928,N_11810,N_11450);
nand U11929 (N_11929,N_11455,N_11452);
nand U11930 (N_11930,N_11696,N_11626);
nand U11931 (N_11931,N_11663,N_11624);
and U11932 (N_11932,N_11764,N_11294);
and U11933 (N_11933,N_11369,N_11654);
or U11934 (N_11934,N_11325,N_11550);
and U11935 (N_11935,N_11768,N_11568);
and U11936 (N_11936,N_11344,N_11656);
and U11937 (N_11937,N_11767,N_11614);
and U11938 (N_11938,N_11556,N_11256);
and U11939 (N_11939,N_11672,N_11280);
and U11940 (N_11940,N_11382,N_11841);
nand U11941 (N_11941,N_11857,N_11808);
nor U11942 (N_11942,N_11426,N_11509);
nand U11943 (N_11943,N_11331,N_11312);
or U11944 (N_11944,N_11845,N_11712);
nor U11945 (N_11945,N_11391,N_11856);
nor U11946 (N_11946,N_11791,N_11313);
and U11947 (N_11947,N_11639,N_11319);
nand U11948 (N_11948,N_11359,N_11636);
or U11949 (N_11949,N_11667,N_11744);
nand U11950 (N_11950,N_11368,N_11514);
and U11951 (N_11951,N_11572,N_11378);
xor U11952 (N_11952,N_11813,N_11410);
nand U11953 (N_11953,N_11554,N_11725);
or U11954 (N_11954,N_11464,N_11543);
nor U11955 (N_11955,N_11282,N_11496);
and U11956 (N_11956,N_11427,N_11400);
nor U11957 (N_11957,N_11862,N_11660);
and U11958 (N_11958,N_11437,N_11716);
and U11959 (N_11959,N_11704,N_11812);
and U11960 (N_11960,N_11482,N_11362);
and U11961 (N_11961,N_11531,N_11567);
nor U11962 (N_11962,N_11357,N_11575);
or U11963 (N_11963,N_11558,N_11760);
or U11964 (N_11964,N_11476,N_11601);
or U11965 (N_11965,N_11536,N_11458);
or U11966 (N_11966,N_11775,N_11609);
or U11967 (N_11967,N_11755,N_11350);
or U11968 (N_11968,N_11817,N_11860);
nand U11969 (N_11969,N_11610,N_11442);
and U11970 (N_11970,N_11646,N_11621);
and U11971 (N_11971,N_11408,N_11618);
nand U11972 (N_11972,N_11720,N_11537);
and U11973 (N_11973,N_11526,N_11762);
nand U11974 (N_11974,N_11462,N_11848);
and U11975 (N_11975,N_11335,N_11589);
xnor U11976 (N_11976,N_11622,N_11258);
nor U11977 (N_11977,N_11519,N_11500);
nor U11978 (N_11978,N_11598,N_11394);
xor U11979 (N_11979,N_11499,N_11534);
or U11980 (N_11980,N_11295,N_11267);
or U11981 (N_11981,N_11512,N_11707);
nor U11982 (N_11982,N_11647,N_11306);
nor U11983 (N_11983,N_11435,N_11721);
nand U11984 (N_11984,N_11375,N_11852);
nor U11985 (N_11985,N_11265,N_11292);
nor U11986 (N_11986,N_11287,N_11376);
xnor U11987 (N_11987,N_11459,N_11388);
or U11988 (N_11988,N_11846,N_11474);
xnor U11989 (N_11989,N_11798,N_11365);
xnor U11990 (N_11990,N_11340,N_11428);
nor U11991 (N_11991,N_11831,N_11715);
xnor U11992 (N_11992,N_11806,N_11433);
nand U11993 (N_11993,N_11456,N_11513);
or U11994 (N_11994,N_11574,N_11865);
or U11995 (N_11995,N_11257,N_11772);
and U11996 (N_11996,N_11671,N_11676);
or U11997 (N_11997,N_11669,N_11599);
nor U11998 (N_11998,N_11782,N_11466);
and U11999 (N_11999,N_11439,N_11827);
nand U12000 (N_12000,N_11835,N_11854);
xor U12001 (N_12001,N_11726,N_11872);
nor U12002 (N_12002,N_11364,N_11487);
and U12003 (N_12003,N_11529,N_11327);
nand U12004 (N_12004,N_11805,N_11839);
and U12005 (N_12005,N_11858,N_11528);
nand U12006 (N_12006,N_11398,N_11718);
and U12007 (N_12007,N_11395,N_11826);
nand U12008 (N_12008,N_11561,N_11301);
and U12009 (N_12009,N_11465,N_11665);
and U12010 (N_12010,N_11800,N_11661);
nor U12011 (N_12011,N_11738,N_11830);
or U12012 (N_12012,N_11343,N_11489);
or U12013 (N_12013,N_11396,N_11684);
and U12014 (N_12014,N_11758,N_11743);
nand U12015 (N_12015,N_11700,N_11863);
or U12016 (N_12016,N_11493,N_11734);
or U12017 (N_12017,N_11592,N_11341);
and U12018 (N_12018,N_11436,N_11784);
or U12019 (N_12019,N_11263,N_11405);
or U12020 (N_12020,N_11771,N_11510);
and U12021 (N_12021,N_11285,N_11309);
nand U12022 (N_12022,N_11687,N_11776);
or U12023 (N_12023,N_11270,N_11380);
nand U12024 (N_12024,N_11328,N_11740);
and U12025 (N_12025,N_11747,N_11677);
nor U12026 (N_12026,N_11674,N_11480);
nor U12027 (N_12027,N_11491,N_11403);
or U12028 (N_12028,N_11494,N_11807);
and U12029 (N_12029,N_11315,N_11754);
and U12030 (N_12030,N_11421,N_11787);
nand U12031 (N_12031,N_11330,N_11460);
xor U12032 (N_12032,N_11652,N_11593);
nand U12033 (N_12033,N_11607,N_11516);
or U12034 (N_12034,N_11385,N_11802);
and U12035 (N_12035,N_11613,N_11641);
xor U12036 (N_12036,N_11794,N_11645);
xor U12037 (N_12037,N_11616,N_11602);
or U12038 (N_12038,N_11454,N_11431);
and U12039 (N_12039,N_11705,N_11785);
xnor U12040 (N_12040,N_11416,N_11290);
nor U12041 (N_12041,N_11255,N_11300);
nor U12042 (N_12042,N_11730,N_11584);
nand U12043 (N_12043,N_11681,N_11275);
nor U12044 (N_12044,N_11565,N_11520);
and U12045 (N_12045,N_11644,N_11634);
and U12046 (N_12046,N_11316,N_11658);
or U12047 (N_12047,N_11527,N_11483);
and U12048 (N_12048,N_11399,N_11837);
or U12049 (N_12049,N_11850,N_11861);
or U12050 (N_12050,N_11630,N_11430);
nor U12051 (N_12051,N_11864,N_11662);
nand U12052 (N_12052,N_11276,N_11596);
or U12053 (N_12053,N_11745,N_11505);
nand U12054 (N_12054,N_11836,N_11322);
or U12055 (N_12055,N_11659,N_11296);
nor U12056 (N_12056,N_11648,N_11264);
xor U12057 (N_12057,N_11492,N_11855);
and U12058 (N_12058,N_11457,N_11311);
xnor U12059 (N_12059,N_11606,N_11517);
nand U12060 (N_12060,N_11724,N_11790);
nand U12061 (N_12061,N_11305,N_11283);
nor U12062 (N_12062,N_11711,N_11686);
xnor U12063 (N_12063,N_11588,N_11642);
nand U12064 (N_12064,N_11511,N_11409);
nand U12065 (N_12065,N_11495,N_11337);
nand U12066 (N_12066,N_11261,N_11298);
or U12067 (N_12067,N_11441,N_11541);
nand U12068 (N_12068,N_11346,N_11870);
nand U12069 (N_12069,N_11419,N_11360);
nand U12070 (N_12070,N_11498,N_11816);
nor U12071 (N_12071,N_11549,N_11502);
and U12072 (N_12072,N_11587,N_11867);
or U12073 (N_12073,N_11293,N_11518);
nor U12074 (N_12074,N_11414,N_11297);
xnor U12075 (N_12075,N_11279,N_11544);
nand U12076 (N_12076,N_11389,N_11417);
nor U12077 (N_12077,N_11737,N_11443);
nor U12078 (N_12078,N_11748,N_11728);
nand U12079 (N_12079,N_11332,N_11424);
nor U12080 (N_12080,N_11418,N_11673);
nor U12081 (N_12081,N_11467,N_11451);
nor U12082 (N_12082,N_11627,N_11566);
and U12083 (N_12083,N_11643,N_11339);
xnor U12084 (N_12084,N_11629,N_11666);
and U12085 (N_12085,N_11635,N_11779);
xor U12086 (N_12086,N_11582,N_11254);
and U12087 (N_12087,N_11769,N_11307);
and U12088 (N_12088,N_11569,N_11851);
and U12089 (N_12089,N_11273,N_11548);
nor U12090 (N_12090,N_11625,N_11585);
nor U12091 (N_12091,N_11559,N_11367);
or U12092 (N_12092,N_11538,N_11605);
and U12093 (N_12093,N_11342,N_11253);
and U12094 (N_12094,N_11373,N_11871);
xor U12095 (N_12095,N_11463,N_11788);
nor U12096 (N_12096,N_11501,N_11352);
and U12097 (N_12097,N_11553,N_11525);
or U12098 (N_12098,N_11678,N_11633);
nand U12099 (N_12099,N_11742,N_11372);
xor U12100 (N_12100,N_11591,N_11680);
or U12101 (N_12101,N_11440,N_11688);
nand U12102 (N_12102,N_11384,N_11377);
nor U12103 (N_12103,N_11397,N_11326);
nand U12104 (N_12104,N_11523,N_11485);
nor U12105 (N_12105,N_11766,N_11628);
xor U12106 (N_12106,N_11338,N_11825);
nor U12107 (N_12107,N_11321,N_11545);
nor U12108 (N_12108,N_11425,N_11336);
nand U12109 (N_12109,N_11438,N_11302);
nor U12110 (N_12110,N_11522,N_11824);
and U12111 (N_12111,N_11552,N_11532);
and U12112 (N_12112,N_11822,N_11404);
or U12113 (N_12113,N_11706,N_11801);
and U12114 (N_12114,N_11353,N_11371);
xor U12115 (N_12115,N_11268,N_11479);
and U12116 (N_12116,N_11484,N_11694);
nor U12117 (N_12117,N_11318,N_11578);
and U12118 (N_12118,N_11780,N_11847);
nand U12119 (N_12119,N_11717,N_11803);
nor U12120 (N_12120,N_11597,N_11570);
and U12121 (N_12121,N_11849,N_11761);
or U12122 (N_12122,N_11354,N_11429);
and U12123 (N_12123,N_11655,N_11379);
or U12124 (N_12124,N_11733,N_11792);
or U12125 (N_12125,N_11521,N_11562);
or U12126 (N_12126,N_11530,N_11590);
nand U12127 (N_12127,N_11551,N_11469);
nor U12128 (N_12128,N_11868,N_11383);
nor U12129 (N_12129,N_11407,N_11709);
and U12130 (N_12130,N_11811,N_11756);
and U12131 (N_12131,N_11535,N_11693);
nor U12132 (N_12132,N_11299,N_11615);
and U12133 (N_12133,N_11415,N_11844);
and U12134 (N_12134,N_11752,N_11508);
nand U12135 (N_12135,N_11260,N_11833);
or U12136 (N_12136,N_11657,N_11729);
nor U12137 (N_12137,N_11580,N_11668);
nand U12138 (N_12138,N_11586,N_11746);
nand U12139 (N_12139,N_11675,N_11564);
nand U12140 (N_12140,N_11692,N_11763);
or U12141 (N_12141,N_11555,N_11722);
nor U12142 (N_12142,N_11732,N_11392);
or U12143 (N_12143,N_11649,N_11488);
nor U12144 (N_12144,N_11507,N_11750);
nor U12145 (N_12145,N_11617,N_11583);
nand U12146 (N_12146,N_11804,N_11470);
or U12147 (N_12147,N_11797,N_11573);
nand U12148 (N_12148,N_11799,N_11739);
and U12149 (N_12149,N_11370,N_11540);
or U12150 (N_12150,N_11640,N_11832);
or U12151 (N_12151,N_11736,N_11333);
nand U12152 (N_12152,N_11363,N_11366);
nand U12153 (N_12153,N_11577,N_11444);
or U12154 (N_12154,N_11713,N_11702);
nor U12155 (N_12155,N_11266,N_11560);
nand U12156 (N_12156,N_11468,N_11348);
nand U12157 (N_12157,N_11434,N_11781);
nand U12158 (N_12158,N_11581,N_11869);
and U12159 (N_12159,N_11361,N_11284);
or U12160 (N_12160,N_11557,N_11783);
nand U12161 (N_12161,N_11347,N_11679);
or U12162 (N_12162,N_11539,N_11432);
nand U12163 (N_12163,N_11698,N_11820);
nor U12164 (N_12164,N_11471,N_11259);
or U12165 (N_12165,N_11834,N_11793);
nand U12166 (N_12166,N_11571,N_11304);
and U12167 (N_12167,N_11701,N_11796);
nor U12168 (N_12168,N_11735,N_11349);
nor U12169 (N_12169,N_11274,N_11271);
nor U12170 (N_12170,N_11623,N_11524);
nor U12171 (N_12171,N_11355,N_11604);
nand U12172 (N_12172,N_11477,N_11563);
or U12173 (N_12173,N_11840,N_11420);
nand U12174 (N_12174,N_11446,N_11608);
xor U12175 (N_12175,N_11757,N_11314);
or U12176 (N_12176,N_11329,N_11818);
nor U12177 (N_12177,N_11272,N_11579);
nor U12178 (N_12178,N_11828,N_11448);
or U12179 (N_12179,N_11486,N_11594);
xor U12180 (N_12180,N_11401,N_11269);
nor U12181 (N_12181,N_11413,N_11320);
and U12182 (N_12182,N_11289,N_11708);
nor U12183 (N_12183,N_11447,N_11873);
nor U12184 (N_12184,N_11770,N_11504);
or U12185 (N_12185,N_11612,N_11751);
xnor U12186 (N_12186,N_11727,N_11406);
xnor U12187 (N_12187,N_11685,N_11647);
and U12188 (N_12188,N_11407,N_11558);
nor U12189 (N_12189,N_11833,N_11376);
nand U12190 (N_12190,N_11552,N_11706);
nand U12191 (N_12191,N_11346,N_11494);
nor U12192 (N_12192,N_11402,N_11720);
and U12193 (N_12193,N_11868,N_11530);
nor U12194 (N_12194,N_11350,N_11868);
nand U12195 (N_12195,N_11649,N_11726);
nor U12196 (N_12196,N_11625,N_11396);
nand U12197 (N_12197,N_11492,N_11591);
nor U12198 (N_12198,N_11792,N_11538);
nor U12199 (N_12199,N_11791,N_11479);
nand U12200 (N_12200,N_11409,N_11605);
or U12201 (N_12201,N_11665,N_11682);
or U12202 (N_12202,N_11488,N_11425);
nand U12203 (N_12203,N_11873,N_11602);
or U12204 (N_12204,N_11463,N_11405);
nor U12205 (N_12205,N_11780,N_11868);
or U12206 (N_12206,N_11483,N_11662);
nor U12207 (N_12207,N_11368,N_11720);
and U12208 (N_12208,N_11845,N_11817);
or U12209 (N_12209,N_11309,N_11347);
nand U12210 (N_12210,N_11364,N_11396);
nand U12211 (N_12211,N_11253,N_11827);
or U12212 (N_12212,N_11619,N_11659);
and U12213 (N_12213,N_11693,N_11474);
or U12214 (N_12214,N_11692,N_11717);
xnor U12215 (N_12215,N_11293,N_11345);
and U12216 (N_12216,N_11377,N_11398);
nand U12217 (N_12217,N_11375,N_11656);
nor U12218 (N_12218,N_11345,N_11463);
or U12219 (N_12219,N_11414,N_11258);
nor U12220 (N_12220,N_11849,N_11637);
or U12221 (N_12221,N_11469,N_11581);
nor U12222 (N_12222,N_11819,N_11548);
or U12223 (N_12223,N_11338,N_11683);
and U12224 (N_12224,N_11640,N_11545);
xnor U12225 (N_12225,N_11369,N_11469);
nand U12226 (N_12226,N_11810,N_11558);
nand U12227 (N_12227,N_11763,N_11752);
or U12228 (N_12228,N_11356,N_11422);
and U12229 (N_12229,N_11543,N_11548);
nor U12230 (N_12230,N_11874,N_11367);
or U12231 (N_12231,N_11587,N_11428);
and U12232 (N_12232,N_11326,N_11622);
and U12233 (N_12233,N_11313,N_11720);
xor U12234 (N_12234,N_11398,N_11499);
xnor U12235 (N_12235,N_11722,N_11781);
nand U12236 (N_12236,N_11292,N_11634);
nor U12237 (N_12237,N_11463,N_11832);
xor U12238 (N_12238,N_11528,N_11601);
nand U12239 (N_12239,N_11528,N_11801);
nand U12240 (N_12240,N_11294,N_11405);
nor U12241 (N_12241,N_11730,N_11804);
nor U12242 (N_12242,N_11459,N_11307);
or U12243 (N_12243,N_11417,N_11642);
nand U12244 (N_12244,N_11537,N_11291);
xor U12245 (N_12245,N_11870,N_11786);
nand U12246 (N_12246,N_11622,N_11364);
or U12247 (N_12247,N_11660,N_11769);
nor U12248 (N_12248,N_11501,N_11710);
nand U12249 (N_12249,N_11720,N_11254);
nor U12250 (N_12250,N_11279,N_11609);
or U12251 (N_12251,N_11613,N_11738);
xor U12252 (N_12252,N_11639,N_11398);
nor U12253 (N_12253,N_11626,N_11350);
and U12254 (N_12254,N_11808,N_11632);
nor U12255 (N_12255,N_11592,N_11869);
and U12256 (N_12256,N_11403,N_11767);
and U12257 (N_12257,N_11788,N_11869);
and U12258 (N_12258,N_11698,N_11375);
and U12259 (N_12259,N_11261,N_11464);
or U12260 (N_12260,N_11415,N_11516);
or U12261 (N_12261,N_11558,N_11459);
nand U12262 (N_12262,N_11578,N_11477);
nor U12263 (N_12263,N_11389,N_11324);
nor U12264 (N_12264,N_11589,N_11496);
or U12265 (N_12265,N_11697,N_11512);
and U12266 (N_12266,N_11405,N_11266);
and U12267 (N_12267,N_11334,N_11465);
nor U12268 (N_12268,N_11722,N_11359);
nand U12269 (N_12269,N_11398,N_11259);
nor U12270 (N_12270,N_11384,N_11347);
nand U12271 (N_12271,N_11414,N_11754);
nand U12272 (N_12272,N_11596,N_11511);
nor U12273 (N_12273,N_11869,N_11736);
nor U12274 (N_12274,N_11389,N_11372);
or U12275 (N_12275,N_11521,N_11648);
and U12276 (N_12276,N_11418,N_11433);
or U12277 (N_12277,N_11370,N_11867);
and U12278 (N_12278,N_11393,N_11365);
and U12279 (N_12279,N_11565,N_11473);
or U12280 (N_12280,N_11313,N_11563);
or U12281 (N_12281,N_11553,N_11725);
xnor U12282 (N_12282,N_11689,N_11581);
nor U12283 (N_12283,N_11769,N_11640);
xnor U12284 (N_12284,N_11456,N_11272);
nand U12285 (N_12285,N_11540,N_11746);
or U12286 (N_12286,N_11519,N_11773);
nor U12287 (N_12287,N_11826,N_11599);
nor U12288 (N_12288,N_11276,N_11680);
nor U12289 (N_12289,N_11683,N_11755);
or U12290 (N_12290,N_11299,N_11599);
and U12291 (N_12291,N_11432,N_11292);
and U12292 (N_12292,N_11420,N_11717);
or U12293 (N_12293,N_11648,N_11693);
nand U12294 (N_12294,N_11545,N_11567);
nor U12295 (N_12295,N_11564,N_11668);
xor U12296 (N_12296,N_11392,N_11298);
nand U12297 (N_12297,N_11517,N_11285);
nor U12298 (N_12298,N_11254,N_11451);
nor U12299 (N_12299,N_11675,N_11548);
nor U12300 (N_12300,N_11509,N_11815);
or U12301 (N_12301,N_11489,N_11459);
xor U12302 (N_12302,N_11361,N_11461);
nor U12303 (N_12303,N_11735,N_11279);
and U12304 (N_12304,N_11682,N_11469);
nor U12305 (N_12305,N_11759,N_11847);
and U12306 (N_12306,N_11671,N_11489);
and U12307 (N_12307,N_11667,N_11333);
nand U12308 (N_12308,N_11395,N_11415);
and U12309 (N_12309,N_11840,N_11256);
nor U12310 (N_12310,N_11529,N_11515);
nand U12311 (N_12311,N_11457,N_11394);
nand U12312 (N_12312,N_11570,N_11656);
nor U12313 (N_12313,N_11577,N_11850);
nor U12314 (N_12314,N_11513,N_11701);
or U12315 (N_12315,N_11766,N_11319);
nor U12316 (N_12316,N_11344,N_11724);
nand U12317 (N_12317,N_11721,N_11429);
nand U12318 (N_12318,N_11254,N_11305);
or U12319 (N_12319,N_11790,N_11499);
and U12320 (N_12320,N_11316,N_11747);
nor U12321 (N_12321,N_11360,N_11667);
nor U12322 (N_12322,N_11636,N_11803);
nand U12323 (N_12323,N_11862,N_11478);
nand U12324 (N_12324,N_11715,N_11772);
nor U12325 (N_12325,N_11848,N_11365);
and U12326 (N_12326,N_11836,N_11673);
nand U12327 (N_12327,N_11575,N_11323);
nor U12328 (N_12328,N_11600,N_11316);
and U12329 (N_12329,N_11720,N_11667);
and U12330 (N_12330,N_11441,N_11767);
nor U12331 (N_12331,N_11752,N_11606);
xnor U12332 (N_12332,N_11374,N_11844);
and U12333 (N_12333,N_11827,N_11513);
nand U12334 (N_12334,N_11814,N_11492);
nand U12335 (N_12335,N_11500,N_11540);
nor U12336 (N_12336,N_11692,N_11595);
nor U12337 (N_12337,N_11481,N_11529);
and U12338 (N_12338,N_11273,N_11547);
xnor U12339 (N_12339,N_11421,N_11629);
and U12340 (N_12340,N_11665,N_11263);
and U12341 (N_12341,N_11358,N_11261);
and U12342 (N_12342,N_11685,N_11397);
and U12343 (N_12343,N_11442,N_11810);
nor U12344 (N_12344,N_11383,N_11547);
or U12345 (N_12345,N_11867,N_11421);
nor U12346 (N_12346,N_11842,N_11663);
nand U12347 (N_12347,N_11312,N_11595);
and U12348 (N_12348,N_11580,N_11264);
or U12349 (N_12349,N_11597,N_11555);
or U12350 (N_12350,N_11273,N_11352);
xnor U12351 (N_12351,N_11845,N_11621);
xnor U12352 (N_12352,N_11350,N_11320);
nor U12353 (N_12353,N_11626,N_11431);
nor U12354 (N_12354,N_11832,N_11288);
nor U12355 (N_12355,N_11446,N_11781);
or U12356 (N_12356,N_11476,N_11365);
nand U12357 (N_12357,N_11507,N_11796);
and U12358 (N_12358,N_11377,N_11340);
nor U12359 (N_12359,N_11817,N_11519);
nand U12360 (N_12360,N_11637,N_11618);
xor U12361 (N_12361,N_11302,N_11768);
and U12362 (N_12362,N_11831,N_11508);
or U12363 (N_12363,N_11484,N_11567);
and U12364 (N_12364,N_11672,N_11376);
or U12365 (N_12365,N_11615,N_11853);
xor U12366 (N_12366,N_11655,N_11848);
or U12367 (N_12367,N_11580,N_11635);
and U12368 (N_12368,N_11293,N_11532);
and U12369 (N_12369,N_11693,N_11686);
or U12370 (N_12370,N_11624,N_11323);
and U12371 (N_12371,N_11316,N_11591);
or U12372 (N_12372,N_11855,N_11673);
nor U12373 (N_12373,N_11435,N_11818);
nand U12374 (N_12374,N_11436,N_11621);
and U12375 (N_12375,N_11869,N_11358);
xnor U12376 (N_12376,N_11788,N_11312);
nand U12377 (N_12377,N_11738,N_11583);
or U12378 (N_12378,N_11725,N_11870);
or U12379 (N_12379,N_11466,N_11438);
and U12380 (N_12380,N_11267,N_11325);
nand U12381 (N_12381,N_11425,N_11528);
xnor U12382 (N_12382,N_11406,N_11549);
nand U12383 (N_12383,N_11322,N_11377);
or U12384 (N_12384,N_11740,N_11330);
xnor U12385 (N_12385,N_11550,N_11384);
nand U12386 (N_12386,N_11822,N_11472);
nor U12387 (N_12387,N_11635,N_11835);
xor U12388 (N_12388,N_11637,N_11630);
nand U12389 (N_12389,N_11773,N_11428);
nor U12390 (N_12390,N_11862,N_11589);
nand U12391 (N_12391,N_11566,N_11761);
nand U12392 (N_12392,N_11613,N_11273);
and U12393 (N_12393,N_11463,N_11458);
or U12394 (N_12394,N_11268,N_11609);
nor U12395 (N_12395,N_11409,N_11523);
nor U12396 (N_12396,N_11336,N_11468);
xnor U12397 (N_12397,N_11585,N_11794);
nor U12398 (N_12398,N_11464,N_11751);
and U12399 (N_12399,N_11862,N_11787);
nand U12400 (N_12400,N_11375,N_11740);
and U12401 (N_12401,N_11442,N_11850);
xor U12402 (N_12402,N_11362,N_11741);
nand U12403 (N_12403,N_11562,N_11252);
nand U12404 (N_12404,N_11867,N_11787);
nor U12405 (N_12405,N_11400,N_11491);
and U12406 (N_12406,N_11462,N_11437);
nor U12407 (N_12407,N_11615,N_11865);
nand U12408 (N_12408,N_11439,N_11410);
nor U12409 (N_12409,N_11843,N_11664);
nor U12410 (N_12410,N_11346,N_11270);
xor U12411 (N_12411,N_11486,N_11616);
nand U12412 (N_12412,N_11766,N_11638);
nand U12413 (N_12413,N_11396,N_11516);
nand U12414 (N_12414,N_11553,N_11782);
nor U12415 (N_12415,N_11462,N_11749);
nor U12416 (N_12416,N_11562,N_11561);
nand U12417 (N_12417,N_11303,N_11583);
nor U12418 (N_12418,N_11481,N_11869);
nor U12419 (N_12419,N_11805,N_11339);
xor U12420 (N_12420,N_11290,N_11643);
or U12421 (N_12421,N_11725,N_11272);
or U12422 (N_12422,N_11665,N_11284);
nand U12423 (N_12423,N_11506,N_11752);
nand U12424 (N_12424,N_11568,N_11593);
or U12425 (N_12425,N_11837,N_11416);
or U12426 (N_12426,N_11359,N_11300);
nor U12427 (N_12427,N_11378,N_11556);
and U12428 (N_12428,N_11739,N_11584);
nor U12429 (N_12429,N_11352,N_11461);
nand U12430 (N_12430,N_11422,N_11447);
nor U12431 (N_12431,N_11670,N_11604);
nor U12432 (N_12432,N_11520,N_11651);
nor U12433 (N_12433,N_11564,N_11586);
or U12434 (N_12434,N_11572,N_11447);
or U12435 (N_12435,N_11544,N_11548);
or U12436 (N_12436,N_11782,N_11539);
or U12437 (N_12437,N_11827,N_11422);
nor U12438 (N_12438,N_11773,N_11654);
nor U12439 (N_12439,N_11465,N_11252);
nand U12440 (N_12440,N_11518,N_11341);
and U12441 (N_12441,N_11592,N_11863);
xor U12442 (N_12442,N_11737,N_11565);
or U12443 (N_12443,N_11335,N_11664);
nor U12444 (N_12444,N_11796,N_11346);
nand U12445 (N_12445,N_11786,N_11616);
and U12446 (N_12446,N_11509,N_11530);
nand U12447 (N_12447,N_11479,N_11347);
nor U12448 (N_12448,N_11586,N_11733);
nand U12449 (N_12449,N_11515,N_11282);
nor U12450 (N_12450,N_11450,N_11378);
or U12451 (N_12451,N_11784,N_11515);
nor U12452 (N_12452,N_11721,N_11419);
nor U12453 (N_12453,N_11338,N_11541);
xor U12454 (N_12454,N_11636,N_11752);
nand U12455 (N_12455,N_11452,N_11664);
xor U12456 (N_12456,N_11849,N_11513);
and U12457 (N_12457,N_11721,N_11516);
and U12458 (N_12458,N_11837,N_11287);
and U12459 (N_12459,N_11647,N_11638);
and U12460 (N_12460,N_11809,N_11670);
and U12461 (N_12461,N_11692,N_11784);
or U12462 (N_12462,N_11464,N_11479);
nor U12463 (N_12463,N_11372,N_11587);
and U12464 (N_12464,N_11853,N_11669);
nor U12465 (N_12465,N_11314,N_11386);
nand U12466 (N_12466,N_11749,N_11411);
nand U12467 (N_12467,N_11630,N_11705);
nand U12468 (N_12468,N_11820,N_11455);
and U12469 (N_12469,N_11520,N_11581);
or U12470 (N_12470,N_11309,N_11664);
nand U12471 (N_12471,N_11301,N_11446);
and U12472 (N_12472,N_11402,N_11597);
nand U12473 (N_12473,N_11478,N_11790);
nand U12474 (N_12474,N_11558,N_11826);
and U12475 (N_12475,N_11744,N_11493);
nor U12476 (N_12476,N_11476,N_11750);
or U12477 (N_12477,N_11490,N_11274);
or U12478 (N_12478,N_11850,N_11540);
xnor U12479 (N_12479,N_11658,N_11370);
xnor U12480 (N_12480,N_11284,N_11752);
or U12481 (N_12481,N_11267,N_11825);
nor U12482 (N_12482,N_11818,N_11688);
xor U12483 (N_12483,N_11734,N_11565);
or U12484 (N_12484,N_11608,N_11672);
xnor U12485 (N_12485,N_11458,N_11654);
nand U12486 (N_12486,N_11601,N_11506);
xnor U12487 (N_12487,N_11427,N_11254);
nand U12488 (N_12488,N_11493,N_11602);
or U12489 (N_12489,N_11759,N_11668);
and U12490 (N_12490,N_11831,N_11686);
nand U12491 (N_12491,N_11852,N_11670);
nor U12492 (N_12492,N_11815,N_11326);
or U12493 (N_12493,N_11816,N_11268);
and U12494 (N_12494,N_11790,N_11335);
and U12495 (N_12495,N_11253,N_11697);
nor U12496 (N_12496,N_11570,N_11414);
nor U12497 (N_12497,N_11505,N_11555);
nand U12498 (N_12498,N_11393,N_11861);
xnor U12499 (N_12499,N_11416,N_11669);
nand U12500 (N_12500,N_12150,N_12023);
xor U12501 (N_12501,N_12381,N_12018);
and U12502 (N_12502,N_12144,N_11926);
nand U12503 (N_12503,N_12186,N_11913);
nor U12504 (N_12504,N_12413,N_12232);
nand U12505 (N_12505,N_12180,N_12184);
or U12506 (N_12506,N_12099,N_12455);
nand U12507 (N_12507,N_12187,N_12147);
nand U12508 (N_12508,N_11877,N_12353);
and U12509 (N_12509,N_12448,N_11948);
nor U12510 (N_12510,N_11876,N_12121);
or U12511 (N_12511,N_11960,N_12272);
nand U12512 (N_12512,N_11957,N_12400);
xor U12513 (N_12513,N_12211,N_12071);
or U12514 (N_12514,N_12252,N_12346);
nand U12515 (N_12515,N_12473,N_12468);
and U12516 (N_12516,N_12243,N_12214);
nand U12517 (N_12517,N_12484,N_11944);
or U12518 (N_12518,N_12410,N_12287);
or U12519 (N_12519,N_11911,N_12225);
nand U12520 (N_12520,N_12055,N_12148);
nor U12521 (N_12521,N_12335,N_12409);
and U12522 (N_12522,N_12193,N_12207);
or U12523 (N_12523,N_11924,N_11943);
xor U12524 (N_12524,N_12034,N_12212);
nor U12525 (N_12525,N_11880,N_12163);
xor U12526 (N_12526,N_12160,N_12191);
xnor U12527 (N_12527,N_12117,N_12269);
or U12528 (N_12528,N_12462,N_12161);
or U12529 (N_12529,N_12192,N_12495);
xor U12530 (N_12530,N_11975,N_12472);
and U12531 (N_12531,N_12258,N_11942);
nand U12532 (N_12532,N_12102,N_12320);
nor U12533 (N_12533,N_12053,N_12376);
nand U12534 (N_12534,N_12299,N_12303);
xor U12535 (N_12535,N_12266,N_11965);
or U12536 (N_12536,N_12218,N_12429);
or U12537 (N_12537,N_11908,N_12227);
nor U12538 (N_12538,N_12097,N_12137);
or U12539 (N_12539,N_11983,N_12329);
or U12540 (N_12540,N_11879,N_12242);
nand U12541 (N_12541,N_12190,N_11995);
and U12542 (N_12542,N_12419,N_11930);
nand U12543 (N_12543,N_12444,N_12103);
and U12544 (N_12544,N_12426,N_12246);
nand U12545 (N_12545,N_11976,N_12222);
and U12546 (N_12546,N_12255,N_12306);
nor U12547 (N_12547,N_12067,N_11999);
or U12548 (N_12548,N_12321,N_12402);
nand U12549 (N_12549,N_12364,N_12213);
and U12550 (N_12550,N_12088,N_12136);
and U12551 (N_12551,N_11977,N_12465);
xnor U12552 (N_12552,N_11900,N_12479);
nand U12553 (N_12553,N_11917,N_12074);
or U12554 (N_12554,N_12307,N_12334);
nor U12555 (N_12555,N_12384,N_12058);
xnor U12556 (N_12556,N_12296,N_12267);
and U12557 (N_12557,N_12302,N_12134);
nor U12558 (N_12558,N_12265,N_11914);
or U12559 (N_12559,N_12205,N_12133);
nand U12560 (N_12560,N_12124,N_12156);
or U12561 (N_12561,N_12342,N_11988);
and U12562 (N_12562,N_11893,N_11909);
and U12563 (N_12563,N_12268,N_12172);
nor U12564 (N_12564,N_12003,N_12069);
nor U12565 (N_12565,N_12285,N_12417);
and U12566 (N_12566,N_12349,N_12217);
and U12567 (N_12567,N_12141,N_12322);
or U12568 (N_12568,N_11969,N_12026);
nand U12569 (N_12569,N_12399,N_12151);
nor U12570 (N_12570,N_12294,N_12254);
nor U12571 (N_12571,N_12263,N_12314);
and U12572 (N_12572,N_12092,N_11918);
or U12573 (N_12573,N_12203,N_12244);
nand U12574 (N_12574,N_12100,N_12290);
or U12575 (N_12575,N_12230,N_11994);
or U12576 (N_12576,N_12079,N_12408);
and U12577 (N_12577,N_12139,N_12024);
nor U12578 (N_12578,N_12428,N_12486);
or U12579 (N_12579,N_12378,N_12389);
or U12580 (N_12580,N_12273,N_12446);
or U12581 (N_12581,N_12293,N_12499);
nand U12582 (N_12582,N_12339,N_12105);
nand U12583 (N_12583,N_12206,N_12281);
nand U12584 (N_12584,N_11937,N_11940);
nand U12585 (N_12585,N_12131,N_12166);
nand U12586 (N_12586,N_12391,N_12220);
or U12587 (N_12587,N_12398,N_12453);
and U12588 (N_12588,N_12138,N_12310);
and U12589 (N_12589,N_11993,N_12330);
nand U12590 (N_12590,N_12326,N_12075);
nand U12591 (N_12591,N_12096,N_12280);
or U12592 (N_12592,N_11952,N_12009);
or U12593 (N_12593,N_12028,N_11915);
nand U12594 (N_12594,N_12475,N_12056);
and U12595 (N_12595,N_12210,N_11898);
xor U12596 (N_12596,N_11916,N_12171);
nand U12597 (N_12597,N_12070,N_12279);
nor U12598 (N_12598,N_12081,N_11963);
nor U12599 (N_12599,N_11936,N_12177);
and U12600 (N_12600,N_12434,N_12316);
and U12601 (N_12601,N_12292,N_11949);
and U12602 (N_12602,N_12372,N_11885);
nor U12603 (N_12603,N_12460,N_12315);
nand U12604 (N_12604,N_11902,N_12140);
nand U12605 (N_12605,N_12392,N_12328);
and U12606 (N_12606,N_12345,N_12343);
nor U12607 (N_12607,N_11928,N_11888);
and U12608 (N_12608,N_11984,N_12149);
nor U12609 (N_12609,N_11886,N_12135);
xnor U12610 (N_12610,N_12275,N_12062);
or U12611 (N_12611,N_12492,N_11989);
nand U12612 (N_12612,N_12078,N_12439);
xor U12613 (N_12613,N_12411,N_12032);
and U12614 (N_12614,N_12194,N_12235);
nand U12615 (N_12615,N_12170,N_12017);
and U12616 (N_12616,N_11979,N_12437);
and U12617 (N_12617,N_12371,N_12282);
nand U12618 (N_12618,N_12189,N_11951);
xor U12619 (N_12619,N_12311,N_12167);
and U12620 (N_12620,N_12481,N_12174);
nand U12621 (N_12621,N_12489,N_11891);
nor U12622 (N_12622,N_12030,N_12424);
or U12623 (N_12623,N_12083,N_12301);
nand U12624 (N_12624,N_12035,N_12241);
xnor U12625 (N_12625,N_12388,N_12435);
nand U12626 (N_12626,N_12297,N_12498);
and U12627 (N_12627,N_12188,N_12236);
nor U12628 (N_12628,N_11882,N_11933);
nand U12629 (N_12629,N_12129,N_12120);
nand U12630 (N_12630,N_12060,N_11892);
nor U12631 (N_12631,N_12383,N_12000);
and U12632 (N_12632,N_11967,N_11887);
nor U12633 (N_12633,N_12045,N_12040);
nand U12634 (N_12634,N_12277,N_12362);
nor U12635 (N_12635,N_12039,N_11987);
nand U12636 (N_12636,N_12101,N_12029);
nand U12637 (N_12637,N_11927,N_12332);
and U12638 (N_12638,N_12317,N_12354);
and U12639 (N_12639,N_12065,N_11910);
and U12640 (N_12640,N_12262,N_12361);
nor U12641 (N_12641,N_12229,N_12366);
xor U12642 (N_12642,N_11945,N_12084);
xor U12643 (N_12643,N_11932,N_12404);
and U12644 (N_12644,N_11990,N_12260);
nor U12645 (N_12645,N_12369,N_12360);
and U12646 (N_12646,N_12432,N_12431);
nor U12647 (N_12647,N_12393,N_12031);
or U12648 (N_12648,N_11878,N_12365);
nand U12649 (N_12649,N_12022,N_12179);
or U12650 (N_12650,N_12412,N_12086);
nor U12651 (N_12651,N_12142,N_12005);
or U12652 (N_12652,N_11929,N_12198);
nor U12653 (N_12653,N_12082,N_12199);
nor U12654 (N_12654,N_11923,N_12430);
nand U12655 (N_12655,N_11890,N_12041);
nand U12656 (N_12656,N_11946,N_12452);
nand U12657 (N_12657,N_11959,N_12123);
xnor U12658 (N_12658,N_12348,N_12467);
nand U12659 (N_12659,N_12112,N_12338);
nand U12660 (N_12660,N_12340,N_12350);
and U12661 (N_12661,N_12458,N_11935);
and U12662 (N_12662,N_12415,N_12368);
or U12663 (N_12663,N_11980,N_12333);
and U12664 (N_12664,N_12356,N_12471);
nand U12665 (N_12665,N_12158,N_12497);
or U12666 (N_12666,N_12020,N_12228);
and U12667 (N_12667,N_12438,N_11972);
or U12668 (N_12668,N_12216,N_12487);
nand U12669 (N_12669,N_11991,N_12363);
nor U12670 (N_12670,N_12049,N_12089);
nor U12671 (N_12671,N_12323,N_12401);
nor U12672 (N_12672,N_12164,N_12196);
nand U12673 (N_12673,N_12240,N_12226);
nor U12674 (N_12674,N_12488,N_12178);
nand U12675 (N_12675,N_12480,N_11922);
or U12676 (N_12676,N_12113,N_12386);
nor U12677 (N_12677,N_11903,N_12450);
nor U12678 (N_12678,N_12331,N_12173);
or U12679 (N_12679,N_11964,N_12204);
xnor U12680 (N_12680,N_12093,N_12390);
or U12681 (N_12681,N_12110,N_12238);
and U12682 (N_12682,N_12042,N_12445);
nand U12683 (N_12683,N_12491,N_12048);
nand U12684 (N_12684,N_12394,N_12051);
nor U12685 (N_12685,N_11919,N_12490);
or U12686 (N_12686,N_12341,N_12066);
and U12687 (N_12687,N_11875,N_11889);
and U12688 (N_12688,N_12397,N_12012);
and U12689 (N_12689,N_11997,N_12143);
xor U12690 (N_12690,N_11974,N_12200);
and U12691 (N_12691,N_12256,N_12385);
nor U12692 (N_12692,N_12403,N_12441);
nor U12693 (N_12693,N_11941,N_12251);
nor U12694 (N_12694,N_12168,N_11962);
or U12695 (N_12695,N_12010,N_12037);
nor U12696 (N_12696,N_12312,N_12118);
nand U12697 (N_12697,N_11897,N_12483);
xnor U12698 (N_12698,N_11934,N_12061);
or U12699 (N_12699,N_12215,N_12091);
or U12700 (N_12700,N_12406,N_12059);
or U12701 (N_12701,N_12208,N_12283);
or U12702 (N_12702,N_12063,N_12237);
xnor U12703 (N_12703,N_12496,N_12457);
nand U12704 (N_12704,N_12057,N_11998);
or U12705 (N_12705,N_12154,N_12440);
or U12706 (N_12706,N_11953,N_12153);
or U12707 (N_12707,N_11961,N_11966);
nor U12708 (N_12708,N_12033,N_12318);
nor U12709 (N_12709,N_12182,N_12347);
nand U12710 (N_12710,N_12375,N_12351);
xnor U12711 (N_12711,N_12344,N_12248);
and U12712 (N_12712,N_12370,N_12423);
or U12713 (N_12713,N_12261,N_12264);
xnor U12714 (N_12714,N_12016,N_12373);
and U12715 (N_12715,N_12271,N_12485);
and U12716 (N_12716,N_12175,N_12427);
nor U12717 (N_12717,N_12231,N_12132);
nand U12718 (N_12718,N_11985,N_12197);
and U12719 (N_12719,N_12108,N_12374);
nand U12720 (N_12720,N_12305,N_12433);
nor U12721 (N_12721,N_12352,N_12477);
and U12722 (N_12722,N_12414,N_12098);
and U12723 (N_12723,N_11938,N_12195);
nand U12724 (N_12724,N_12224,N_12127);
xnor U12725 (N_12725,N_12202,N_12044);
nand U12726 (N_12726,N_12476,N_12052);
and U12727 (N_12727,N_12126,N_12181);
nand U12728 (N_12728,N_11920,N_12001);
nand U12729 (N_12729,N_11986,N_12221);
nor U12730 (N_12730,N_12270,N_12289);
and U12731 (N_12731,N_12219,N_12185);
nand U12732 (N_12732,N_11896,N_12077);
nand U12733 (N_12733,N_11912,N_12159);
xnor U12734 (N_12734,N_11905,N_12443);
nor U12735 (N_12735,N_12464,N_12257);
and U12736 (N_12736,N_11992,N_12358);
nand U12737 (N_12737,N_12493,N_12116);
nand U12738 (N_12738,N_12245,N_12380);
xnor U12739 (N_12739,N_12111,N_12064);
xor U12740 (N_12740,N_12122,N_12407);
or U12741 (N_12741,N_12395,N_11947);
nand U12742 (N_12742,N_12157,N_12463);
nand U12743 (N_12743,N_12313,N_12019);
nor U12744 (N_12744,N_12309,N_12233);
or U12745 (N_12745,N_11899,N_12085);
nand U12746 (N_12746,N_12359,N_11981);
nand U12747 (N_12747,N_12405,N_11895);
or U12748 (N_12748,N_12253,N_12014);
nand U12749 (N_12749,N_12046,N_12308);
and U12750 (N_12750,N_12119,N_12461);
nor U12751 (N_12751,N_12336,N_11958);
and U12752 (N_12752,N_12259,N_12201);
nor U12753 (N_12753,N_12021,N_12145);
and U12754 (N_12754,N_12416,N_12087);
nand U12755 (N_12755,N_12274,N_12288);
nor U12756 (N_12756,N_12165,N_12325);
and U12757 (N_12757,N_12436,N_12209);
and U12758 (N_12758,N_12109,N_12276);
nand U12759 (N_12759,N_12454,N_12013);
or U12760 (N_12760,N_11968,N_11955);
nor U12761 (N_12761,N_12470,N_12080);
and U12762 (N_12762,N_11894,N_12011);
and U12763 (N_12763,N_12025,N_12015);
nor U12764 (N_12764,N_12146,N_12449);
xnor U12765 (N_12765,N_12456,N_11907);
nor U12766 (N_12766,N_12298,N_12447);
xnor U12767 (N_12767,N_12115,N_12291);
xnor U12768 (N_12768,N_12073,N_12072);
nor U12769 (N_12769,N_12278,N_12043);
or U12770 (N_12770,N_11925,N_12425);
nor U12771 (N_12771,N_11921,N_11956);
and U12772 (N_12772,N_12008,N_12169);
xnor U12773 (N_12773,N_12054,N_12076);
nor U12774 (N_12774,N_12300,N_11931);
or U12775 (N_12775,N_11904,N_11954);
nand U12776 (N_12776,N_12068,N_11901);
or U12777 (N_12777,N_12295,N_12387);
nand U12778 (N_12778,N_12234,N_11939);
nand U12779 (N_12779,N_12250,N_12442);
xnor U12780 (N_12780,N_12130,N_12451);
or U12781 (N_12781,N_12036,N_11906);
nor U12782 (N_12782,N_12478,N_12247);
and U12783 (N_12783,N_12337,N_12367);
nor U12784 (N_12784,N_12382,N_12104);
and U12785 (N_12785,N_12494,N_12038);
and U12786 (N_12786,N_11970,N_12357);
and U12787 (N_12787,N_12162,N_12466);
nor U12788 (N_12788,N_11973,N_12286);
nand U12789 (N_12789,N_12094,N_12155);
nand U12790 (N_12790,N_12421,N_12418);
nand U12791 (N_12791,N_12125,N_12183);
nor U12792 (N_12792,N_12324,N_12007);
nor U12793 (N_12793,N_11971,N_12469);
xnor U12794 (N_12794,N_12249,N_11883);
nand U12795 (N_12795,N_12004,N_12006);
and U12796 (N_12796,N_12050,N_12152);
nor U12797 (N_12797,N_12319,N_12047);
and U12798 (N_12798,N_11996,N_12304);
nand U12799 (N_12799,N_12095,N_12027);
and U12800 (N_12800,N_11884,N_12459);
nor U12801 (N_12801,N_12107,N_12128);
nor U12802 (N_12802,N_12422,N_12474);
and U12803 (N_12803,N_12106,N_12396);
xnor U12804 (N_12804,N_12002,N_12090);
nand U12805 (N_12805,N_12284,N_12114);
or U12806 (N_12806,N_12377,N_12223);
xnor U12807 (N_12807,N_12420,N_11950);
and U12808 (N_12808,N_11881,N_12239);
nand U12809 (N_12809,N_12327,N_11978);
xor U12810 (N_12810,N_11982,N_12379);
nor U12811 (N_12811,N_12355,N_12482);
nor U12812 (N_12812,N_12176,N_12389);
and U12813 (N_12813,N_12198,N_12363);
nand U12814 (N_12814,N_12467,N_12119);
xor U12815 (N_12815,N_12035,N_12406);
nor U12816 (N_12816,N_11920,N_12351);
and U12817 (N_12817,N_11971,N_12139);
nand U12818 (N_12818,N_12122,N_12038);
nor U12819 (N_12819,N_12121,N_12227);
nand U12820 (N_12820,N_12031,N_12046);
and U12821 (N_12821,N_11911,N_12155);
and U12822 (N_12822,N_11990,N_11979);
or U12823 (N_12823,N_12312,N_12026);
nand U12824 (N_12824,N_12394,N_12085);
nand U12825 (N_12825,N_11881,N_12344);
nor U12826 (N_12826,N_12340,N_12087);
and U12827 (N_12827,N_12474,N_12314);
and U12828 (N_12828,N_12305,N_11884);
or U12829 (N_12829,N_12049,N_12221);
and U12830 (N_12830,N_12212,N_12487);
and U12831 (N_12831,N_11945,N_12174);
nor U12832 (N_12832,N_12353,N_12181);
or U12833 (N_12833,N_12145,N_12361);
and U12834 (N_12834,N_12177,N_12119);
or U12835 (N_12835,N_12477,N_12094);
xor U12836 (N_12836,N_12160,N_11935);
xor U12837 (N_12837,N_12131,N_12221);
or U12838 (N_12838,N_12282,N_12219);
and U12839 (N_12839,N_12428,N_12463);
nand U12840 (N_12840,N_12070,N_12003);
or U12841 (N_12841,N_12071,N_12095);
and U12842 (N_12842,N_12471,N_12476);
nor U12843 (N_12843,N_11987,N_12276);
and U12844 (N_12844,N_12038,N_12076);
nand U12845 (N_12845,N_11883,N_12267);
and U12846 (N_12846,N_11929,N_12138);
or U12847 (N_12847,N_12420,N_12136);
xor U12848 (N_12848,N_12072,N_12247);
nand U12849 (N_12849,N_12256,N_12280);
or U12850 (N_12850,N_12313,N_12138);
nor U12851 (N_12851,N_11890,N_12103);
nand U12852 (N_12852,N_11933,N_12209);
nand U12853 (N_12853,N_12140,N_12424);
and U12854 (N_12854,N_12089,N_11988);
or U12855 (N_12855,N_12404,N_12489);
nor U12856 (N_12856,N_12009,N_12431);
nand U12857 (N_12857,N_12353,N_12362);
or U12858 (N_12858,N_12446,N_11906);
or U12859 (N_12859,N_11902,N_12316);
and U12860 (N_12860,N_12230,N_12065);
nand U12861 (N_12861,N_12490,N_12015);
nor U12862 (N_12862,N_12035,N_12390);
xor U12863 (N_12863,N_12346,N_12051);
or U12864 (N_12864,N_12031,N_12112);
xnor U12865 (N_12865,N_12225,N_12250);
and U12866 (N_12866,N_12102,N_11992);
nor U12867 (N_12867,N_12280,N_12473);
nand U12868 (N_12868,N_12000,N_12488);
or U12869 (N_12869,N_12297,N_12448);
nand U12870 (N_12870,N_12365,N_12130);
nor U12871 (N_12871,N_12258,N_12397);
and U12872 (N_12872,N_12372,N_12222);
and U12873 (N_12873,N_11998,N_12410);
and U12874 (N_12874,N_12060,N_12232);
xor U12875 (N_12875,N_12466,N_12416);
nor U12876 (N_12876,N_12201,N_11949);
xnor U12877 (N_12877,N_12477,N_12155);
and U12878 (N_12878,N_11914,N_12060);
and U12879 (N_12879,N_11973,N_12406);
nor U12880 (N_12880,N_12213,N_12417);
and U12881 (N_12881,N_12336,N_12467);
nor U12882 (N_12882,N_11998,N_12252);
nand U12883 (N_12883,N_11891,N_12491);
nand U12884 (N_12884,N_12069,N_12214);
nor U12885 (N_12885,N_12138,N_11951);
nand U12886 (N_12886,N_12301,N_12297);
or U12887 (N_12887,N_12034,N_12303);
xnor U12888 (N_12888,N_12353,N_12338);
and U12889 (N_12889,N_12442,N_12294);
or U12890 (N_12890,N_12061,N_12365);
nand U12891 (N_12891,N_11923,N_11877);
nor U12892 (N_12892,N_12455,N_12162);
and U12893 (N_12893,N_12366,N_12321);
and U12894 (N_12894,N_12035,N_11877);
and U12895 (N_12895,N_12284,N_12257);
or U12896 (N_12896,N_12263,N_12358);
xnor U12897 (N_12897,N_12085,N_11981);
and U12898 (N_12898,N_12304,N_12325);
xor U12899 (N_12899,N_12411,N_11938);
nand U12900 (N_12900,N_12280,N_11951);
nand U12901 (N_12901,N_12338,N_12160);
or U12902 (N_12902,N_12356,N_12064);
or U12903 (N_12903,N_12388,N_12403);
nor U12904 (N_12904,N_12020,N_12176);
or U12905 (N_12905,N_11936,N_12462);
nand U12906 (N_12906,N_12356,N_12095);
and U12907 (N_12907,N_11956,N_12334);
and U12908 (N_12908,N_11937,N_12456);
and U12909 (N_12909,N_11965,N_12457);
xor U12910 (N_12910,N_12440,N_12077);
and U12911 (N_12911,N_12006,N_12270);
nand U12912 (N_12912,N_12027,N_11894);
xor U12913 (N_12913,N_12064,N_12152);
nor U12914 (N_12914,N_12433,N_12065);
xor U12915 (N_12915,N_12462,N_12309);
nor U12916 (N_12916,N_12461,N_12274);
and U12917 (N_12917,N_12483,N_12052);
and U12918 (N_12918,N_12496,N_12210);
nand U12919 (N_12919,N_12320,N_12383);
and U12920 (N_12920,N_12214,N_11884);
nor U12921 (N_12921,N_11966,N_12275);
and U12922 (N_12922,N_12440,N_12366);
xnor U12923 (N_12923,N_12186,N_12275);
nor U12924 (N_12924,N_12060,N_12369);
nand U12925 (N_12925,N_12006,N_12441);
or U12926 (N_12926,N_12495,N_11897);
and U12927 (N_12927,N_12248,N_12063);
nor U12928 (N_12928,N_12265,N_12120);
nor U12929 (N_12929,N_12437,N_11917);
or U12930 (N_12930,N_11966,N_12423);
nand U12931 (N_12931,N_12084,N_12090);
nor U12932 (N_12932,N_11921,N_12260);
nand U12933 (N_12933,N_11932,N_11968);
nand U12934 (N_12934,N_12177,N_12434);
nor U12935 (N_12935,N_12277,N_12198);
nand U12936 (N_12936,N_12054,N_11976);
nand U12937 (N_12937,N_12335,N_12282);
or U12938 (N_12938,N_12095,N_11985);
and U12939 (N_12939,N_12174,N_12479);
and U12940 (N_12940,N_12031,N_11970);
nor U12941 (N_12941,N_11967,N_11981);
nand U12942 (N_12942,N_12415,N_12212);
or U12943 (N_12943,N_11937,N_12277);
or U12944 (N_12944,N_11993,N_12344);
and U12945 (N_12945,N_12438,N_12236);
nor U12946 (N_12946,N_11937,N_12353);
and U12947 (N_12947,N_12373,N_12236);
or U12948 (N_12948,N_12102,N_12449);
nand U12949 (N_12949,N_11966,N_12042);
nor U12950 (N_12950,N_11932,N_11940);
nor U12951 (N_12951,N_12122,N_12328);
and U12952 (N_12952,N_12334,N_12102);
or U12953 (N_12953,N_11942,N_12128);
xnor U12954 (N_12954,N_12129,N_11939);
and U12955 (N_12955,N_12402,N_12156);
or U12956 (N_12956,N_12387,N_12228);
nand U12957 (N_12957,N_12250,N_12430);
or U12958 (N_12958,N_12446,N_12022);
and U12959 (N_12959,N_12365,N_11879);
nor U12960 (N_12960,N_11946,N_12493);
nor U12961 (N_12961,N_12338,N_11971);
nor U12962 (N_12962,N_12273,N_12471);
nand U12963 (N_12963,N_12143,N_12176);
nand U12964 (N_12964,N_12457,N_12260);
xor U12965 (N_12965,N_12223,N_12369);
nor U12966 (N_12966,N_12090,N_12495);
xnor U12967 (N_12967,N_12455,N_12065);
xor U12968 (N_12968,N_12141,N_12116);
or U12969 (N_12969,N_12238,N_12282);
or U12970 (N_12970,N_12367,N_12437);
or U12971 (N_12971,N_12337,N_12146);
nand U12972 (N_12972,N_12324,N_11970);
and U12973 (N_12973,N_12322,N_11941);
and U12974 (N_12974,N_11989,N_12185);
and U12975 (N_12975,N_12027,N_12127);
nand U12976 (N_12976,N_11888,N_12065);
nand U12977 (N_12977,N_12210,N_12498);
xor U12978 (N_12978,N_12163,N_12369);
xor U12979 (N_12979,N_12436,N_11898);
nor U12980 (N_12980,N_11974,N_12286);
or U12981 (N_12981,N_12166,N_12051);
nor U12982 (N_12982,N_12485,N_12216);
or U12983 (N_12983,N_12237,N_11881);
xnor U12984 (N_12984,N_12006,N_12230);
nand U12985 (N_12985,N_11893,N_11892);
xor U12986 (N_12986,N_12075,N_12113);
nor U12987 (N_12987,N_12113,N_12480);
nor U12988 (N_12988,N_12146,N_12410);
and U12989 (N_12989,N_12481,N_12262);
nand U12990 (N_12990,N_12298,N_11939);
nor U12991 (N_12991,N_11883,N_12215);
or U12992 (N_12992,N_12192,N_12029);
and U12993 (N_12993,N_11884,N_12027);
nand U12994 (N_12994,N_12031,N_12213);
or U12995 (N_12995,N_11965,N_11905);
nand U12996 (N_12996,N_11886,N_12088);
nand U12997 (N_12997,N_12113,N_11900);
or U12998 (N_12998,N_12422,N_12010);
nor U12999 (N_12999,N_11938,N_12159);
nand U13000 (N_13000,N_12264,N_12217);
and U13001 (N_13001,N_12450,N_12427);
nor U13002 (N_13002,N_12312,N_11949);
nor U13003 (N_13003,N_12210,N_11951);
nor U13004 (N_13004,N_11983,N_11956);
nor U13005 (N_13005,N_11980,N_11979);
and U13006 (N_13006,N_12267,N_11915);
nand U13007 (N_13007,N_12474,N_12224);
nand U13008 (N_13008,N_12220,N_12056);
or U13009 (N_13009,N_11890,N_11904);
and U13010 (N_13010,N_12243,N_12306);
or U13011 (N_13011,N_12053,N_11906);
or U13012 (N_13012,N_12327,N_12201);
nor U13013 (N_13013,N_11999,N_12339);
nor U13014 (N_13014,N_12209,N_12131);
nand U13015 (N_13015,N_11887,N_12357);
nor U13016 (N_13016,N_11979,N_12302);
or U13017 (N_13017,N_12477,N_12466);
or U13018 (N_13018,N_12275,N_12430);
nand U13019 (N_13019,N_12446,N_12314);
nand U13020 (N_13020,N_11975,N_12449);
or U13021 (N_13021,N_12450,N_12364);
and U13022 (N_13022,N_12138,N_12373);
xnor U13023 (N_13023,N_12099,N_12463);
and U13024 (N_13024,N_12206,N_12335);
and U13025 (N_13025,N_12432,N_11885);
and U13026 (N_13026,N_12041,N_12305);
nand U13027 (N_13027,N_12317,N_12051);
and U13028 (N_13028,N_11945,N_11925);
nor U13029 (N_13029,N_12375,N_12472);
or U13030 (N_13030,N_12126,N_12098);
and U13031 (N_13031,N_12253,N_12243);
or U13032 (N_13032,N_12415,N_11905);
and U13033 (N_13033,N_12125,N_12289);
or U13034 (N_13034,N_12037,N_12185);
or U13035 (N_13035,N_12455,N_12051);
nand U13036 (N_13036,N_12069,N_12368);
and U13037 (N_13037,N_12239,N_11939);
xnor U13038 (N_13038,N_12093,N_12312);
or U13039 (N_13039,N_12121,N_12337);
nand U13040 (N_13040,N_12202,N_12109);
or U13041 (N_13041,N_12082,N_12069);
nor U13042 (N_13042,N_11968,N_12350);
nor U13043 (N_13043,N_12079,N_11999);
nand U13044 (N_13044,N_12340,N_12111);
nand U13045 (N_13045,N_12246,N_12183);
nand U13046 (N_13046,N_12466,N_12168);
nand U13047 (N_13047,N_12452,N_12403);
or U13048 (N_13048,N_12164,N_12363);
or U13049 (N_13049,N_12298,N_12401);
nand U13050 (N_13050,N_12439,N_11994);
or U13051 (N_13051,N_12379,N_11998);
nor U13052 (N_13052,N_11943,N_12267);
nor U13053 (N_13053,N_12065,N_12480);
nor U13054 (N_13054,N_12225,N_12448);
or U13055 (N_13055,N_12161,N_12063);
nand U13056 (N_13056,N_12341,N_12240);
nor U13057 (N_13057,N_12228,N_11893);
nor U13058 (N_13058,N_11885,N_12495);
nand U13059 (N_13059,N_12059,N_12429);
or U13060 (N_13060,N_12328,N_12189);
and U13061 (N_13061,N_12166,N_12161);
nor U13062 (N_13062,N_12252,N_11982);
or U13063 (N_13063,N_12484,N_12089);
nor U13064 (N_13064,N_12410,N_11887);
nor U13065 (N_13065,N_12160,N_12431);
nand U13066 (N_13066,N_12177,N_12343);
nor U13067 (N_13067,N_12099,N_12242);
or U13068 (N_13068,N_11946,N_12307);
nand U13069 (N_13069,N_12464,N_12173);
or U13070 (N_13070,N_12038,N_11957);
or U13071 (N_13071,N_12271,N_12278);
nor U13072 (N_13072,N_12243,N_12166);
or U13073 (N_13073,N_12382,N_12486);
and U13074 (N_13074,N_12308,N_12085);
or U13075 (N_13075,N_12286,N_12300);
or U13076 (N_13076,N_11954,N_12418);
nand U13077 (N_13077,N_12254,N_12337);
or U13078 (N_13078,N_12014,N_12056);
and U13079 (N_13079,N_12051,N_12407);
and U13080 (N_13080,N_12377,N_12200);
nand U13081 (N_13081,N_12194,N_12403);
nand U13082 (N_13082,N_12483,N_12010);
or U13083 (N_13083,N_11928,N_12144);
nor U13084 (N_13084,N_12201,N_12036);
and U13085 (N_13085,N_12197,N_12230);
xnor U13086 (N_13086,N_12094,N_12340);
nand U13087 (N_13087,N_11986,N_12351);
or U13088 (N_13088,N_12326,N_12422);
or U13089 (N_13089,N_12443,N_12112);
nand U13090 (N_13090,N_12123,N_12259);
nor U13091 (N_13091,N_12044,N_12367);
nand U13092 (N_13092,N_12092,N_12053);
or U13093 (N_13093,N_12426,N_11986);
xor U13094 (N_13094,N_12395,N_11883);
nor U13095 (N_13095,N_11877,N_12326);
xnor U13096 (N_13096,N_12224,N_12290);
xor U13097 (N_13097,N_12452,N_12278);
nand U13098 (N_13098,N_12276,N_12094);
nor U13099 (N_13099,N_12175,N_12182);
nand U13100 (N_13100,N_12367,N_12257);
or U13101 (N_13101,N_12271,N_12163);
or U13102 (N_13102,N_11892,N_12180);
or U13103 (N_13103,N_12387,N_12150);
or U13104 (N_13104,N_11877,N_12161);
nor U13105 (N_13105,N_12296,N_12482);
nand U13106 (N_13106,N_11953,N_12402);
xor U13107 (N_13107,N_12244,N_12161);
or U13108 (N_13108,N_12044,N_12305);
nor U13109 (N_13109,N_12013,N_12050);
or U13110 (N_13110,N_11900,N_11890);
xnor U13111 (N_13111,N_11987,N_12452);
nor U13112 (N_13112,N_12238,N_11918);
nor U13113 (N_13113,N_11955,N_12145);
xor U13114 (N_13114,N_12335,N_11945);
nor U13115 (N_13115,N_11956,N_12341);
nor U13116 (N_13116,N_12248,N_12360);
and U13117 (N_13117,N_11960,N_11948);
nor U13118 (N_13118,N_12017,N_12118);
nor U13119 (N_13119,N_12285,N_12233);
nand U13120 (N_13120,N_11892,N_12360);
nand U13121 (N_13121,N_12449,N_12376);
nor U13122 (N_13122,N_12095,N_12322);
nor U13123 (N_13123,N_12372,N_11891);
and U13124 (N_13124,N_11898,N_12028);
or U13125 (N_13125,N_12844,N_12794);
and U13126 (N_13126,N_13073,N_12701);
nor U13127 (N_13127,N_13091,N_12698);
or U13128 (N_13128,N_12569,N_13040);
xnor U13129 (N_13129,N_13028,N_12929);
and U13130 (N_13130,N_12741,N_13048);
or U13131 (N_13131,N_12774,N_12849);
or U13132 (N_13132,N_12557,N_12946);
and U13133 (N_13133,N_12727,N_13099);
or U13134 (N_13134,N_12678,N_12918);
nand U13135 (N_13135,N_12944,N_12853);
nor U13136 (N_13136,N_12745,N_12642);
and U13137 (N_13137,N_13019,N_12668);
or U13138 (N_13138,N_12768,N_12775);
xnor U13139 (N_13139,N_12759,N_12872);
nand U13140 (N_13140,N_13076,N_12613);
or U13141 (N_13141,N_12987,N_13055);
nand U13142 (N_13142,N_12817,N_12735);
nor U13143 (N_13143,N_13121,N_12742);
or U13144 (N_13144,N_12978,N_12605);
or U13145 (N_13145,N_12704,N_13086);
or U13146 (N_13146,N_13089,N_12910);
nand U13147 (N_13147,N_13120,N_12841);
nor U13148 (N_13148,N_12663,N_12680);
and U13149 (N_13149,N_13006,N_12916);
nor U13150 (N_13150,N_12705,N_12536);
or U13151 (N_13151,N_12537,N_12691);
and U13152 (N_13152,N_12512,N_12956);
and U13153 (N_13153,N_13057,N_12685);
and U13154 (N_13154,N_13097,N_13085);
nand U13155 (N_13155,N_12810,N_12693);
nor U13156 (N_13156,N_12554,N_12639);
nor U13157 (N_13157,N_12731,N_12878);
or U13158 (N_13158,N_13066,N_12934);
or U13159 (N_13159,N_12508,N_12836);
nor U13160 (N_13160,N_13020,N_12848);
and U13161 (N_13161,N_13045,N_12711);
and U13162 (N_13162,N_12957,N_13052);
xor U13163 (N_13163,N_12779,N_12656);
nor U13164 (N_13164,N_12764,N_12733);
xor U13165 (N_13165,N_12976,N_12545);
nand U13166 (N_13166,N_13093,N_12912);
or U13167 (N_13167,N_12730,N_12596);
and U13168 (N_13168,N_12887,N_12631);
and U13169 (N_13169,N_12796,N_12591);
or U13170 (N_13170,N_12542,N_12973);
or U13171 (N_13171,N_12869,N_12683);
and U13172 (N_13172,N_12552,N_12861);
or U13173 (N_13173,N_12615,N_12863);
xor U13174 (N_13174,N_13079,N_13000);
nand U13175 (N_13175,N_12833,N_12658);
nand U13176 (N_13176,N_12959,N_12590);
and U13177 (N_13177,N_13050,N_12805);
and U13178 (N_13178,N_12716,N_12576);
or U13179 (N_13179,N_12626,N_12634);
xor U13180 (N_13180,N_12564,N_12824);
or U13181 (N_13181,N_12945,N_12958);
or U13182 (N_13182,N_12669,N_12516);
nand U13183 (N_13183,N_12850,N_12897);
nor U13184 (N_13184,N_12518,N_13108);
nor U13185 (N_13185,N_12773,N_13116);
or U13186 (N_13186,N_12795,N_12769);
and U13187 (N_13187,N_12927,N_12643);
nand U13188 (N_13188,N_13013,N_12835);
nand U13189 (N_13189,N_12601,N_13034);
nor U13190 (N_13190,N_12575,N_13077);
or U13191 (N_13191,N_12780,N_12965);
nand U13192 (N_13192,N_12619,N_12889);
nand U13193 (N_13193,N_12664,N_12837);
nor U13194 (N_13194,N_12649,N_12748);
nand U13195 (N_13195,N_12567,N_12538);
and U13196 (N_13196,N_12938,N_12717);
or U13197 (N_13197,N_12798,N_12936);
and U13198 (N_13198,N_12600,N_13119);
or U13199 (N_13199,N_12931,N_12706);
and U13200 (N_13200,N_12900,N_12988);
nand U13201 (N_13201,N_12722,N_12886);
nand U13202 (N_13202,N_13053,N_13021);
nor U13203 (N_13203,N_12992,N_12939);
nand U13204 (N_13204,N_12905,N_12699);
and U13205 (N_13205,N_12563,N_12829);
nor U13206 (N_13206,N_12989,N_12868);
and U13207 (N_13207,N_12559,N_12708);
nor U13208 (N_13208,N_12790,N_12654);
nand U13209 (N_13209,N_13058,N_12899);
and U13210 (N_13210,N_12804,N_12800);
or U13211 (N_13211,N_12504,N_12502);
nor U13212 (N_13212,N_12550,N_12793);
nor U13213 (N_13213,N_12876,N_12909);
nor U13214 (N_13214,N_12766,N_12855);
or U13215 (N_13215,N_12703,N_12712);
or U13216 (N_13216,N_12879,N_12527);
nor U13217 (N_13217,N_12834,N_12884);
nand U13218 (N_13218,N_12993,N_12534);
or U13219 (N_13219,N_13054,N_12515);
or U13220 (N_13220,N_13035,N_12644);
nand U13221 (N_13221,N_12894,N_12921);
or U13222 (N_13222,N_12924,N_12819);
nand U13223 (N_13223,N_13017,N_13038);
nand U13224 (N_13224,N_12763,N_12906);
or U13225 (N_13225,N_13075,N_12547);
and U13226 (N_13226,N_12581,N_12877);
or U13227 (N_13227,N_13088,N_12867);
nor U13228 (N_13228,N_13025,N_12751);
nand U13229 (N_13229,N_12592,N_13113);
nor U13230 (N_13230,N_12700,N_12635);
nand U13231 (N_13231,N_12568,N_13068);
or U13232 (N_13232,N_12941,N_12570);
and U13233 (N_13233,N_12787,N_12604);
nand U13234 (N_13234,N_13070,N_12666);
nand U13235 (N_13235,N_12714,N_12771);
nor U13236 (N_13236,N_12791,N_12673);
nand U13237 (N_13237,N_12767,N_12636);
and U13238 (N_13238,N_12503,N_12803);
and U13239 (N_13239,N_13015,N_13074);
and U13240 (N_13240,N_12839,N_12828);
nand U13241 (N_13241,N_12566,N_12676);
or U13242 (N_13242,N_12858,N_12937);
or U13243 (N_13243,N_12611,N_12528);
and U13244 (N_13244,N_12873,N_13117);
nand U13245 (N_13245,N_12971,N_13016);
nor U13246 (N_13246,N_13061,N_12648);
nand U13247 (N_13247,N_12926,N_12859);
nor U13248 (N_13248,N_12962,N_12757);
or U13249 (N_13249,N_13063,N_12851);
nand U13250 (N_13250,N_12917,N_12902);
and U13251 (N_13251,N_12792,N_12728);
nor U13252 (N_13252,N_13082,N_12572);
nor U13253 (N_13253,N_13105,N_13112);
nor U13254 (N_13254,N_12770,N_12997);
nand U13255 (N_13255,N_12684,N_12734);
nor U13256 (N_13256,N_12674,N_12895);
nor U13257 (N_13257,N_12786,N_12752);
nand U13258 (N_13258,N_12535,N_12920);
and U13259 (N_13259,N_12638,N_12585);
and U13260 (N_13260,N_12506,N_13114);
and U13261 (N_13261,N_13106,N_12624);
and U13262 (N_13262,N_12651,N_12864);
nor U13263 (N_13263,N_12632,N_12551);
nand U13264 (N_13264,N_12736,N_12577);
and U13265 (N_13265,N_12765,N_12919);
and U13266 (N_13266,N_12726,N_12784);
or U13267 (N_13267,N_12637,N_12583);
nand U13268 (N_13268,N_12911,N_12862);
and U13269 (N_13269,N_12732,N_13011);
nand U13270 (N_13270,N_12820,N_12808);
or U13271 (N_13271,N_12866,N_12578);
nand U13272 (N_13272,N_12606,N_12832);
xor U13273 (N_13273,N_12947,N_13109);
and U13274 (N_13274,N_13004,N_13118);
nor U13275 (N_13275,N_12740,N_12995);
and U13276 (N_13276,N_12645,N_12519);
and U13277 (N_13277,N_12854,N_13030);
and U13278 (N_13278,N_12998,N_12513);
nor U13279 (N_13279,N_13010,N_12620);
nand U13280 (N_13280,N_12826,N_12500);
nor U13281 (N_13281,N_13022,N_12729);
or U13282 (N_13282,N_12893,N_12975);
nor U13283 (N_13283,N_12560,N_12781);
xor U13284 (N_13284,N_12598,N_13051);
or U13285 (N_13285,N_12709,N_12514);
and U13286 (N_13286,N_12687,N_12907);
nand U13287 (N_13287,N_12874,N_12621);
nand U13288 (N_13288,N_12799,N_12540);
or U13289 (N_13289,N_12818,N_12589);
xor U13290 (N_13290,N_12749,N_12614);
or U13291 (N_13291,N_12969,N_12935);
or U13292 (N_13292,N_12718,N_13003);
nor U13293 (N_13293,N_12580,N_12607);
nor U13294 (N_13294,N_12857,N_12949);
nor U13295 (N_13295,N_12772,N_12692);
xor U13296 (N_13296,N_12524,N_12555);
or U13297 (N_13297,N_12558,N_12890);
nor U13298 (N_13298,N_12640,N_12821);
nor U13299 (N_13299,N_12814,N_13012);
xor U13300 (N_13300,N_12659,N_12922);
nor U13301 (N_13301,N_12758,N_12530);
nand U13302 (N_13302,N_13060,N_12677);
nor U13303 (N_13303,N_13027,N_12756);
and U13304 (N_13304,N_13014,N_12831);
or U13305 (N_13305,N_12845,N_12885);
or U13306 (N_13306,N_12671,N_13095);
nand U13307 (N_13307,N_12622,N_12562);
xnor U13308 (N_13308,N_12933,N_12582);
nor U13309 (N_13309,N_12892,N_12737);
nor U13310 (N_13310,N_13026,N_12616);
or U13311 (N_13311,N_13102,N_12594);
or U13312 (N_13312,N_13123,N_12746);
nor U13313 (N_13313,N_12702,N_13092);
nor U13314 (N_13314,N_12517,N_12754);
or U13315 (N_13315,N_12882,N_13065);
or U13316 (N_13316,N_13009,N_12972);
nor U13317 (N_13317,N_13023,N_13072);
nor U13318 (N_13318,N_13107,N_12843);
nor U13319 (N_13319,N_12891,N_12925);
and U13320 (N_13320,N_12608,N_13024);
and U13321 (N_13321,N_12521,N_12801);
and U13322 (N_13322,N_12908,N_12719);
xor U13323 (N_13323,N_12595,N_13033);
or U13324 (N_13324,N_13084,N_13039);
nand U13325 (N_13325,N_12963,N_12830);
and U13326 (N_13326,N_12968,N_12707);
and U13327 (N_13327,N_13056,N_12721);
and U13328 (N_13328,N_12682,N_12695);
or U13329 (N_13329,N_12599,N_12553);
and U13330 (N_13330,N_12541,N_12511);
nor U13331 (N_13331,N_12686,N_12825);
nand U13332 (N_13332,N_12696,N_12915);
xor U13333 (N_13333,N_12549,N_12507);
or U13334 (N_13334,N_12523,N_13115);
or U13335 (N_13335,N_12531,N_12990);
xor U13336 (N_13336,N_12544,N_12565);
nand U13337 (N_13337,N_13044,N_12672);
xnor U13338 (N_13338,N_12739,N_13101);
xor U13339 (N_13339,N_12548,N_12865);
nand U13340 (N_13340,N_12617,N_12623);
nand U13341 (N_13341,N_12667,N_12930);
nor U13342 (N_13342,N_12522,N_12713);
nand U13343 (N_13343,N_13002,N_12710);
nor U13344 (N_13344,N_12625,N_12846);
and U13345 (N_13345,N_12744,N_12966);
nor U13346 (N_13346,N_12602,N_12871);
xnor U13347 (N_13347,N_12657,N_12743);
and U13348 (N_13348,N_13080,N_12630);
or U13349 (N_13349,N_13098,N_12967);
and U13350 (N_13350,N_12982,N_12986);
xor U13351 (N_13351,N_12561,N_12661);
and U13352 (N_13352,N_12812,N_12960);
xnor U13353 (N_13353,N_12951,N_13069);
nand U13354 (N_13354,N_12525,N_12646);
and U13355 (N_13355,N_12755,N_12904);
and U13356 (N_13356,N_12533,N_12943);
nor U13357 (N_13357,N_12655,N_12689);
and U13358 (N_13358,N_12760,N_12778);
or U13359 (N_13359,N_12586,N_12970);
xor U13360 (N_13360,N_12627,N_12579);
or U13361 (N_13361,N_12954,N_12688);
or U13362 (N_13362,N_12815,N_12501);
and U13363 (N_13363,N_12647,N_12520);
nand U13364 (N_13364,N_12811,N_12526);
or U13365 (N_13365,N_12913,N_12928);
and U13366 (N_13366,N_13005,N_12977);
nand U13367 (N_13367,N_13007,N_12964);
or U13368 (N_13368,N_12603,N_13064);
xor U13369 (N_13369,N_12797,N_12510);
nand U13370 (N_13370,N_12984,N_12593);
nor U13371 (N_13371,N_12675,N_12980);
and U13372 (N_13372,N_13041,N_12983);
xor U13373 (N_13373,N_13047,N_13071);
or U13374 (N_13374,N_12783,N_12961);
nor U13375 (N_13375,N_12888,N_12679);
nor U13376 (N_13376,N_12856,N_12923);
and U13377 (N_13377,N_12901,N_12762);
nand U13378 (N_13378,N_12597,N_13046);
or U13379 (N_13379,N_13090,N_12556);
nand U13380 (N_13380,N_12914,N_12694);
nand U13381 (N_13381,N_12952,N_12999);
and U13382 (N_13382,N_12838,N_12785);
and U13383 (N_13383,N_13081,N_12809);
or U13384 (N_13384,N_12653,N_12633);
nor U13385 (N_13385,N_12681,N_12641);
and U13386 (N_13386,N_12822,N_12991);
nand U13387 (N_13387,N_13032,N_13037);
or U13388 (N_13388,N_12628,N_12670);
nor U13389 (N_13389,N_12652,N_12842);
nand U13390 (N_13390,N_12896,N_13049);
nand U13391 (N_13391,N_12573,N_12789);
or U13392 (N_13392,N_13110,N_13036);
or U13393 (N_13393,N_12985,N_13094);
nor U13394 (N_13394,N_12612,N_12932);
or U13395 (N_13395,N_12883,N_13083);
and U13396 (N_13396,N_12750,N_12609);
nand U13397 (N_13397,N_12788,N_12940);
or U13398 (N_13398,N_13111,N_13087);
or U13399 (N_13399,N_13078,N_12584);
nor U13400 (N_13400,N_12546,N_12860);
nor U13401 (N_13401,N_12880,N_13062);
xnor U13402 (N_13402,N_13100,N_12827);
and U13403 (N_13403,N_13103,N_12697);
xor U13404 (N_13404,N_12955,N_12618);
xnor U13405 (N_13405,N_12870,N_12847);
nand U13406 (N_13406,N_12840,N_13104);
nand U13407 (N_13407,N_12996,N_13096);
nor U13408 (N_13408,N_12715,N_12813);
and U13409 (N_13409,N_12807,N_12662);
or U13410 (N_13410,N_12875,N_12881);
and U13411 (N_13411,N_12738,N_12571);
nor U13412 (N_13412,N_12782,N_12660);
nor U13413 (N_13413,N_12505,N_12650);
or U13414 (N_13414,N_13043,N_12950);
nor U13415 (N_13415,N_12974,N_12587);
nand U13416 (N_13416,N_13042,N_12776);
and U13417 (N_13417,N_12747,N_12724);
and U13418 (N_13418,N_12979,N_12725);
nand U13419 (N_13419,N_12610,N_12529);
nor U13420 (N_13420,N_12665,N_12903);
and U13421 (N_13421,N_12948,N_12539);
and U13422 (N_13422,N_12720,N_12690);
nand U13423 (N_13423,N_13067,N_13018);
or U13424 (N_13424,N_13029,N_13008);
nor U13425 (N_13425,N_12802,N_12532);
xnor U13426 (N_13426,N_12574,N_13122);
nand U13427 (N_13427,N_12723,N_12994);
xor U13428 (N_13428,N_13001,N_12543);
nand U13429 (N_13429,N_12777,N_12898);
nor U13430 (N_13430,N_12953,N_12852);
nor U13431 (N_13431,N_12753,N_12509);
xor U13432 (N_13432,N_12981,N_13059);
or U13433 (N_13433,N_13124,N_12942);
and U13434 (N_13434,N_12761,N_12588);
or U13435 (N_13435,N_13031,N_12629);
nor U13436 (N_13436,N_12806,N_12823);
nand U13437 (N_13437,N_12816,N_13058);
nor U13438 (N_13438,N_12976,N_12983);
or U13439 (N_13439,N_12727,N_12805);
or U13440 (N_13440,N_12916,N_12740);
and U13441 (N_13441,N_12669,N_13030);
nor U13442 (N_13442,N_12593,N_12934);
nand U13443 (N_13443,N_12835,N_13028);
and U13444 (N_13444,N_13114,N_12754);
nand U13445 (N_13445,N_12984,N_12881);
or U13446 (N_13446,N_13046,N_12523);
and U13447 (N_13447,N_12558,N_13069);
nand U13448 (N_13448,N_13067,N_12687);
nor U13449 (N_13449,N_12736,N_12727);
nor U13450 (N_13450,N_12772,N_12817);
nand U13451 (N_13451,N_12602,N_12630);
or U13452 (N_13452,N_12513,N_12545);
or U13453 (N_13453,N_13086,N_13030);
xnor U13454 (N_13454,N_12740,N_13120);
nand U13455 (N_13455,N_12612,N_13100);
and U13456 (N_13456,N_12803,N_12700);
and U13457 (N_13457,N_12621,N_12780);
xnor U13458 (N_13458,N_12522,N_12799);
and U13459 (N_13459,N_12950,N_12510);
nor U13460 (N_13460,N_12689,N_12991);
xnor U13461 (N_13461,N_12751,N_12790);
xnor U13462 (N_13462,N_13034,N_12964);
nor U13463 (N_13463,N_12568,N_12949);
or U13464 (N_13464,N_12639,N_12895);
or U13465 (N_13465,N_12878,N_13080);
nand U13466 (N_13466,N_12823,N_12905);
or U13467 (N_13467,N_12573,N_13013);
or U13468 (N_13468,N_13000,N_12520);
nor U13469 (N_13469,N_12974,N_12867);
and U13470 (N_13470,N_12574,N_13081);
nand U13471 (N_13471,N_13011,N_12789);
or U13472 (N_13472,N_12882,N_13083);
nand U13473 (N_13473,N_12964,N_12900);
and U13474 (N_13474,N_12696,N_12899);
or U13475 (N_13475,N_13113,N_12913);
nand U13476 (N_13476,N_13034,N_13006);
nand U13477 (N_13477,N_12625,N_13079);
nand U13478 (N_13478,N_13030,N_12529);
and U13479 (N_13479,N_12963,N_12638);
and U13480 (N_13480,N_12854,N_12780);
nor U13481 (N_13481,N_12960,N_12878);
or U13482 (N_13482,N_12895,N_13070);
xor U13483 (N_13483,N_13094,N_12596);
and U13484 (N_13484,N_12723,N_12753);
or U13485 (N_13485,N_12668,N_12647);
xor U13486 (N_13486,N_12603,N_12737);
and U13487 (N_13487,N_12668,N_12987);
and U13488 (N_13488,N_12712,N_12670);
or U13489 (N_13489,N_12977,N_12617);
and U13490 (N_13490,N_12528,N_12879);
or U13491 (N_13491,N_12981,N_13100);
and U13492 (N_13492,N_12570,N_12546);
nor U13493 (N_13493,N_12805,N_12881);
and U13494 (N_13494,N_12991,N_12922);
or U13495 (N_13495,N_13040,N_12879);
and U13496 (N_13496,N_12734,N_12598);
nand U13497 (N_13497,N_12904,N_13033);
or U13498 (N_13498,N_12657,N_12648);
or U13499 (N_13499,N_13033,N_12991);
and U13500 (N_13500,N_12689,N_12726);
nand U13501 (N_13501,N_13116,N_12758);
and U13502 (N_13502,N_12832,N_12752);
and U13503 (N_13503,N_12585,N_12880);
nand U13504 (N_13504,N_12594,N_13117);
nand U13505 (N_13505,N_12987,N_13038);
nor U13506 (N_13506,N_12850,N_13018);
and U13507 (N_13507,N_13031,N_12819);
or U13508 (N_13508,N_12752,N_12589);
and U13509 (N_13509,N_12507,N_12602);
nor U13510 (N_13510,N_12962,N_13013);
and U13511 (N_13511,N_12827,N_12696);
nor U13512 (N_13512,N_12748,N_12899);
nand U13513 (N_13513,N_12653,N_12955);
or U13514 (N_13514,N_12882,N_12551);
and U13515 (N_13515,N_12518,N_12627);
or U13516 (N_13516,N_12997,N_12524);
nor U13517 (N_13517,N_12531,N_12525);
nor U13518 (N_13518,N_13073,N_12661);
nand U13519 (N_13519,N_12606,N_12609);
xnor U13520 (N_13520,N_12551,N_13042);
nor U13521 (N_13521,N_12526,N_12949);
and U13522 (N_13522,N_12540,N_12703);
nor U13523 (N_13523,N_12732,N_12705);
nor U13524 (N_13524,N_12662,N_12948);
or U13525 (N_13525,N_13072,N_12670);
nor U13526 (N_13526,N_12932,N_12632);
or U13527 (N_13527,N_12610,N_12954);
nand U13528 (N_13528,N_13026,N_12669);
or U13529 (N_13529,N_12950,N_13026);
or U13530 (N_13530,N_12832,N_12939);
nand U13531 (N_13531,N_12619,N_12770);
and U13532 (N_13532,N_12577,N_12728);
and U13533 (N_13533,N_12539,N_13106);
or U13534 (N_13534,N_12952,N_12688);
nand U13535 (N_13535,N_12877,N_12509);
and U13536 (N_13536,N_12983,N_12764);
nor U13537 (N_13537,N_12901,N_12937);
nor U13538 (N_13538,N_12903,N_12598);
and U13539 (N_13539,N_12723,N_12646);
nand U13540 (N_13540,N_12883,N_12991);
or U13541 (N_13541,N_12665,N_12893);
and U13542 (N_13542,N_12978,N_12850);
nand U13543 (N_13543,N_12773,N_12876);
nand U13544 (N_13544,N_12978,N_12759);
nor U13545 (N_13545,N_12841,N_13062);
and U13546 (N_13546,N_13059,N_12755);
or U13547 (N_13547,N_12580,N_12918);
nor U13548 (N_13548,N_12655,N_12750);
or U13549 (N_13549,N_13056,N_12676);
and U13550 (N_13550,N_12881,N_12910);
or U13551 (N_13551,N_12732,N_12742);
nor U13552 (N_13552,N_13029,N_12980);
or U13553 (N_13553,N_12875,N_12851);
nor U13554 (N_13554,N_12879,N_12907);
or U13555 (N_13555,N_12791,N_12948);
or U13556 (N_13556,N_12783,N_12975);
nor U13557 (N_13557,N_12982,N_12929);
and U13558 (N_13558,N_12829,N_12865);
or U13559 (N_13559,N_12955,N_12640);
nand U13560 (N_13560,N_12907,N_12974);
and U13561 (N_13561,N_13124,N_12809);
nor U13562 (N_13562,N_12678,N_12854);
and U13563 (N_13563,N_12713,N_12840);
and U13564 (N_13564,N_12790,N_12780);
and U13565 (N_13565,N_12851,N_12907);
xor U13566 (N_13566,N_13027,N_12842);
nor U13567 (N_13567,N_13077,N_13016);
xnor U13568 (N_13568,N_12930,N_12994);
nor U13569 (N_13569,N_12748,N_13115);
or U13570 (N_13570,N_13051,N_12869);
nand U13571 (N_13571,N_12783,N_13115);
or U13572 (N_13572,N_12790,N_12529);
nand U13573 (N_13573,N_12501,N_12740);
nand U13574 (N_13574,N_12514,N_12775);
nand U13575 (N_13575,N_12551,N_12555);
or U13576 (N_13576,N_12576,N_12949);
nor U13577 (N_13577,N_12881,N_12517);
nor U13578 (N_13578,N_12588,N_12911);
and U13579 (N_13579,N_12546,N_12867);
and U13580 (N_13580,N_13075,N_12874);
nand U13581 (N_13581,N_13065,N_12684);
or U13582 (N_13582,N_12754,N_12883);
nand U13583 (N_13583,N_12638,N_12783);
or U13584 (N_13584,N_12934,N_13004);
nand U13585 (N_13585,N_12670,N_12826);
nand U13586 (N_13586,N_12912,N_12632);
nor U13587 (N_13587,N_12823,N_12602);
nor U13588 (N_13588,N_12836,N_12936);
nor U13589 (N_13589,N_12901,N_12642);
and U13590 (N_13590,N_12541,N_12575);
nand U13591 (N_13591,N_12941,N_13106);
nand U13592 (N_13592,N_13082,N_12809);
or U13593 (N_13593,N_12588,N_12695);
nor U13594 (N_13594,N_13026,N_12576);
nor U13595 (N_13595,N_12703,N_12964);
and U13596 (N_13596,N_12902,N_12711);
nand U13597 (N_13597,N_12673,N_12559);
or U13598 (N_13598,N_12656,N_12595);
and U13599 (N_13599,N_12923,N_12989);
or U13600 (N_13600,N_13031,N_12803);
or U13601 (N_13601,N_12915,N_12528);
nor U13602 (N_13602,N_12705,N_12511);
or U13603 (N_13603,N_12674,N_12858);
nor U13604 (N_13604,N_13038,N_13121);
nor U13605 (N_13605,N_12696,N_12838);
nand U13606 (N_13606,N_12980,N_12775);
nor U13607 (N_13607,N_12545,N_12987);
nor U13608 (N_13608,N_12898,N_12554);
nor U13609 (N_13609,N_13056,N_12556);
and U13610 (N_13610,N_12577,N_12860);
and U13611 (N_13611,N_12816,N_13048);
xnor U13612 (N_13612,N_12673,N_12904);
and U13613 (N_13613,N_12888,N_12775);
xnor U13614 (N_13614,N_13094,N_12620);
or U13615 (N_13615,N_12510,N_13059);
nor U13616 (N_13616,N_12865,N_12725);
nand U13617 (N_13617,N_12793,N_13078);
or U13618 (N_13618,N_12557,N_13079);
and U13619 (N_13619,N_12625,N_12525);
nor U13620 (N_13620,N_13049,N_12527);
nor U13621 (N_13621,N_12607,N_12842);
nor U13622 (N_13622,N_12837,N_12929);
xor U13623 (N_13623,N_12618,N_12956);
nand U13624 (N_13624,N_12991,N_12837);
or U13625 (N_13625,N_12705,N_12528);
or U13626 (N_13626,N_12767,N_12960);
nand U13627 (N_13627,N_12925,N_12644);
or U13628 (N_13628,N_12516,N_12653);
and U13629 (N_13629,N_12729,N_12507);
or U13630 (N_13630,N_13093,N_12835);
and U13631 (N_13631,N_12616,N_12823);
xor U13632 (N_13632,N_13056,N_12577);
nor U13633 (N_13633,N_12983,N_12560);
nand U13634 (N_13634,N_12887,N_12849);
or U13635 (N_13635,N_12898,N_12802);
and U13636 (N_13636,N_12975,N_12614);
and U13637 (N_13637,N_12657,N_12812);
xnor U13638 (N_13638,N_12627,N_12672);
xnor U13639 (N_13639,N_13017,N_12898);
nor U13640 (N_13640,N_13091,N_12893);
or U13641 (N_13641,N_12753,N_12521);
and U13642 (N_13642,N_12882,N_12982);
nor U13643 (N_13643,N_12506,N_13100);
or U13644 (N_13644,N_12888,N_13042);
or U13645 (N_13645,N_12530,N_12991);
or U13646 (N_13646,N_13072,N_13096);
and U13647 (N_13647,N_12984,N_12995);
and U13648 (N_13648,N_13060,N_13071);
nand U13649 (N_13649,N_13120,N_12548);
nand U13650 (N_13650,N_12884,N_12703);
nand U13651 (N_13651,N_13101,N_13078);
nor U13652 (N_13652,N_12877,N_12999);
or U13653 (N_13653,N_12896,N_12709);
and U13654 (N_13654,N_12625,N_12762);
xor U13655 (N_13655,N_13009,N_12501);
nor U13656 (N_13656,N_12867,N_12823);
nor U13657 (N_13657,N_12519,N_12571);
nand U13658 (N_13658,N_12907,N_12503);
xor U13659 (N_13659,N_12761,N_12792);
or U13660 (N_13660,N_12556,N_12801);
nor U13661 (N_13661,N_12903,N_12736);
nand U13662 (N_13662,N_12886,N_13021);
or U13663 (N_13663,N_12829,N_12520);
and U13664 (N_13664,N_13048,N_12673);
nand U13665 (N_13665,N_12950,N_12500);
nand U13666 (N_13666,N_12596,N_13000);
and U13667 (N_13667,N_12552,N_13023);
or U13668 (N_13668,N_13037,N_12598);
or U13669 (N_13669,N_12627,N_12904);
nand U13670 (N_13670,N_12637,N_13000);
nand U13671 (N_13671,N_12847,N_12524);
nor U13672 (N_13672,N_12754,N_12857);
or U13673 (N_13673,N_12650,N_12822);
xnor U13674 (N_13674,N_12939,N_13116);
or U13675 (N_13675,N_13018,N_12598);
xor U13676 (N_13676,N_13017,N_12914);
and U13677 (N_13677,N_12583,N_12815);
nor U13678 (N_13678,N_12562,N_13123);
nor U13679 (N_13679,N_12921,N_12895);
nor U13680 (N_13680,N_12633,N_12608);
or U13681 (N_13681,N_12997,N_12709);
nor U13682 (N_13682,N_13019,N_12754);
and U13683 (N_13683,N_12712,N_12983);
nor U13684 (N_13684,N_12902,N_12573);
nand U13685 (N_13685,N_12927,N_12952);
nand U13686 (N_13686,N_12959,N_12503);
or U13687 (N_13687,N_12752,N_12557);
and U13688 (N_13688,N_12871,N_12961);
and U13689 (N_13689,N_12917,N_12704);
nor U13690 (N_13690,N_12977,N_12578);
or U13691 (N_13691,N_12962,N_12770);
nor U13692 (N_13692,N_12823,N_12675);
nand U13693 (N_13693,N_12988,N_12987);
nor U13694 (N_13694,N_12870,N_13079);
or U13695 (N_13695,N_13055,N_12556);
or U13696 (N_13696,N_12746,N_12512);
or U13697 (N_13697,N_12537,N_12662);
nand U13698 (N_13698,N_12688,N_13071);
nand U13699 (N_13699,N_13057,N_12551);
or U13700 (N_13700,N_12944,N_12713);
nand U13701 (N_13701,N_12809,N_12612);
nand U13702 (N_13702,N_12578,N_13111);
nor U13703 (N_13703,N_12989,N_12573);
and U13704 (N_13704,N_12682,N_12629);
or U13705 (N_13705,N_12522,N_12548);
nand U13706 (N_13706,N_12722,N_12788);
xor U13707 (N_13707,N_13106,N_12546);
or U13708 (N_13708,N_12776,N_12755);
nand U13709 (N_13709,N_12574,N_13096);
nor U13710 (N_13710,N_12794,N_12962);
nand U13711 (N_13711,N_13066,N_12799);
nor U13712 (N_13712,N_12539,N_12887);
nor U13713 (N_13713,N_12568,N_12869);
and U13714 (N_13714,N_12725,N_12704);
nand U13715 (N_13715,N_12919,N_12909);
nor U13716 (N_13716,N_12932,N_12847);
and U13717 (N_13717,N_12880,N_12764);
nor U13718 (N_13718,N_12967,N_12581);
xor U13719 (N_13719,N_12515,N_12858);
and U13720 (N_13720,N_12857,N_12954);
and U13721 (N_13721,N_12609,N_12670);
and U13722 (N_13722,N_13097,N_12688);
or U13723 (N_13723,N_12977,N_12646);
and U13724 (N_13724,N_13101,N_12941);
nand U13725 (N_13725,N_12751,N_12724);
nor U13726 (N_13726,N_12914,N_12705);
nor U13727 (N_13727,N_12724,N_12848);
nor U13728 (N_13728,N_12546,N_12803);
and U13729 (N_13729,N_13048,N_12924);
or U13730 (N_13730,N_12509,N_13079);
xor U13731 (N_13731,N_12620,N_12715);
nor U13732 (N_13732,N_12630,N_13016);
or U13733 (N_13733,N_12903,N_12548);
nand U13734 (N_13734,N_12660,N_12637);
or U13735 (N_13735,N_12567,N_12526);
or U13736 (N_13736,N_13092,N_12803);
nor U13737 (N_13737,N_12582,N_13114);
nor U13738 (N_13738,N_12547,N_12518);
nor U13739 (N_13739,N_12747,N_12570);
nand U13740 (N_13740,N_12793,N_12781);
or U13741 (N_13741,N_12932,N_13038);
nand U13742 (N_13742,N_12614,N_13045);
xor U13743 (N_13743,N_12630,N_12853);
nand U13744 (N_13744,N_12940,N_13056);
or U13745 (N_13745,N_12860,N_12514);
nor U13746 (N_13746,N_12824,N_13031);
nor U13747 (N_13747,N_12533,N_12945);
and U13748 (N_13748,N_12969,N_12798);
and U13749 (N_13749,N_12645,N_12839);
nor U13750 (N_13750,N_13254,N_13154);
nor U13751 (N_13751,N_13234,N_13406);
xor U13752 (N_13752,N_13170,N_13262);
xor U13753 (N_13753,N_13471,N_13683);
or U13754 (N_13754,N_13668,N_13616);
nand U13755 (N_13755,N_13129,N_13309);
nand U13756 (N_13756,N_13670,N_13724);
nand U13757 (N_13757,N_13520,N_13171);
nand U13758 (N_13758,N_13594,N_13696);
nor U13759 (N_13759,N_13585,N_13175);
and U13760 (N_13760,N_13613,N_13287);
nor U13761 (N_13761,N_13235,N_13715);
nand U13762 (N_13762,N_13513,N_13629);
xor U13763 (N_13763,N_13178,N_13223);
nor U13764 (N_13764,N_13230,N_13656);
nor U13765 (N_13765,N_13623,N_13222);
and U13766 (N_13766,N_13172,N_13450);
xnor U13767 (N_13767,N_13276,N_13540);
nand U13768 (N_13768,N_13151,N_13738);
or U13769 (N_13769,N_13425,N_13625);
nand U13770 (N_13770,N_13719,N_13577);
nand U13771 (N_13771,N_13144,N_13675);
nand U13772 (N_13772,N_13581,N_13542);
nor U13773 (N_13773,N_13249,N_13680);
nand U13774 (N_13774,N_13311,N_13664);
xor U13775 (N_13775,N_13229,N_13159);
and U13776 (N_13776,N_13499,N_13631);
or U13777 (N_13777,N_13486,N_13502);
xor U13778 (N_13778,N_13575,N_13663);
nand U13779 (N_13779,N_13231,N_13268);
nand U13780 (N_13780,N_13252,N_13624);
or U13781 (N_13781,N_13557,N_13443);
and U13782 (N_13782,N_13457,N_13560);
nand U13783 (N_13783,N_13605,N_13173);
nor U13784 (N_13784,N_13697,N_13195);
nand U13785 (N_13785,N_13676,N_13487);
nand U13786 (N_13786,N_13459,N_13237);
nor U13787 (N_13787,N_13401,N_13449);
xnor U13788 (N_13788,N_13693,N_13367);
nor U13789 (N_13789,N_13298,N_13387);
nor U13790 (N_13790,N_13704,N_13570);
and U13791 (N_13791,N_13511,N_13141);
nand U13792 (N_13792,N_13305,N_13568);
and U13793 (N_13793,N_13546,N_13208);
or U13794 (N_13794,N_13745,N_13167);
or U13795 (N_13795,N_13211,N_13277);
nor U13796 (N_13796,N_13165,N_13346);
nand U13797 (N_13797,N_13528,N_13140);
nand U13798 (N_13798,N_13348,N_13359);
and U13799 (N_13799,N_13431,N_13498);
nand U13800 (N_13800,N_13391,N_13588);
nand U13801 (N_13801,N_13349,N_13324);
nor U13802 (N_13802,N_13242,N_13283);
nand U13803 (N_13803,N_13727,N_13150);
nor U13804 (N_13804,N_13204,N_13429);
and U13805 (N_13805,N_13410,N_13477);
and U13806 (N_13806,N_13174,N_13257);
and U13807 (N_13807,N_13723,N_13399);
and U13808 (N_13808,N_13317,N_13721);
or U13809 (N_13809,N_13645,N_13294);
nand U13810 (N_13810,N_13428,N_13186);
nor U13811 (N_13811,N_13691,N_13126);
nand U13812 (N_13812,N_13419,N_13571);
and U13813 (N_13813,N_13271,N_13488);
nand U13814 (N_13814,N_13341,N_13319);
nor U13815 (N_13815,N_13344,N_13168);
nor U13816 (N_13816,N_13489,N_13279);
and U13817 (N_13817,N_13632,N_13411);
and U13818 (N_13818,N_13491,N_13325);
or U13819 (N_13819,N_13306,N_13659);
xor U13820 (N_13820,N_13274,N_13197);
nor U13821 (N_13821,N_13470,N_13439);
nand U13822 (N_13822,N_13689,N_13701);
nand U13823 (N_13823,N_13636,N_13381);
nor U13824 (N_13824,N_13127,N_13200);
nor U13825 (N_13825,N_13515,N_13579);
nand U13826 (N_13826,N_13467,N_13203);
nor U13827 (N_13827,N_13650,N_13610);
or U13828 (N_13828,N_13490,N_13558);
or U13829 (N_13829,N_13370,N_13352);
or U13830 (N_13830,N_13238,N_13331);
nor U13831 (N_13831,N_13734,N_13464);
or U13832 (N_13832,N_13576,N_13148);
nor U13833 (N_13833,N_13593,N_13639);
nor U13834 (N_13834,N_13247,N_13420);
nor U13835 (N_13835,N_13627,N_13472);
or U13836 (N_13836,N_13648,N_13493);
and U13837 (N_13837,N_13240,N_13444);
nor U13838 (N_13838,N_13651,N_13714);
nor U13839 (N_13839,N_13149,N_13617);
nor U13840 (N_13840,N_13452,N_13496);
and U13841 (N_13841,N_13382,N_13350);
nor U13842 (N_13842,N_13157,N_13481);
or U13843 (N_13843,N_13469,N_13398);
or U13844 (N_13844,N_13389,N_13649);
nor U13845 (N_13845,N_13363,N_13412);
xor U13846 (N_13846,N_13720,N_13255);
nor U13847 (N_13847,N_13441,N_13674);
or U13848 (N_13848,N_13602,N_13426);
nor U13849 (N_13849,N_13364,N_13404);
nor U13850 (N_13850,N_13531,N_13620);
xor U13851 (N_13851,N_13316,N_13741);
nand U13852 (N_13852,N_13708,N_13589);
xnor U13853 (N_13853,N_13694,N_13518);
nor U13854 (N_13854,N_13226,N_13711);
nand U13855 (N_13855,N_13749,N_13633);
or U13856 (N_13856,N_13534,N_13660);
and U13857 (N_13857,N_13742,N_13156);
or U13858 (N_13858,N_13597,N_13508);
or U13859 (N_13859,N_13574,N_13461);
and U13860 (N_13860,N_13160,N_13747);
and U13861 (N_13861,N_13525,N_13626);
nand U13862 (N_13862,N_13228,N_13572);
nand U13863 (N_13863,N_13296,N_13530);
or U13864 (N_13864,N_13586,N_13308);
or U13865 (N_13865,N_13545,N_13286);
nor U13866 (N_13866,N_13218,N_13686);
nand U13867 (N_13867,N_13604,N_13466);
xor U13868 (N_13868,N_13265,N_13590);
or U13869 (N_13869,N_13512,N_13408);
or U13870 (N_13870,N_13678,N_13264);
or U13871 (N_13871,N_13495,N_13259);
nor U13872 (N_13872,N_13637,N_13563);
or U13873 (N_13873,N_13136,N_13373);
nand U13874 (N_13874,N_13733,N_13462);
nor U13875 (N_13875,N_13554,N_13147);
or U13876 (N_13876,N_13524,N_13288);
nor U13877 (N_13877,N_13374,N_13519);
or U13878 (N_13878,N_13451,N_13722);
or U13879 (N_13879,N_13267,N_13413);
or U13880 (N_13880,N_13337,N_13700);
nand U13881 (N_13881,N_13421,N_13392);
xnor U13882 (N_13882,N_13388,N_13216);
nor U13883 (N_13883,N_13169,N_13740);
or U13884 (N_13884,N_13500,N_13517);
or U13885 (N_13885,N_13281,N_13134);
nor U13886 (N_13886,N_13427,N_13227);
and U13887 (N_13887,N_13282,N_13474);
xnor U13888 (N_13888,N_13698,N_13516);
nor U13889 (N_13889,N_13260,N_13293);
nand U13890 (N_13890,N_13202,N_13166);
nand U13891 (N_13891,N_13125,N_13385);
and U13892 (N_13892,N_13638,N_13552);
nand U13893 (N_13893,N_13191,N_13379);
nand U13894 (N_13894,N_13320,N_13644);
and U13895 (N_13895,N_13333,N_13177);
nand U13896 (N_13896,N_13566,N_13607);
xnor U13897 (N_13897,N_13354,N_13329);
or U13898 (N_13898,N_13403,N_13261);
nand U13899 (N_13899,N_13190,N_13210);
or U13900 (N_13900,N_13556,N_13601);
or U13901 (N_13901,N_13301,N_13395);
xnor U13902 (N_13902,N_13430,N_13330);
nand U13903 (N_13903,N_13219,N_13578);
nand U13904 (N_13904,N_13315,N_13386);
and U13905 (N_13905,N_13608,N_13506);
nand U13906 (N_13906,N_13334,N_13256);
or U13907 (N_13907,N_13299,N_13248);
and U13908 (N_13908,N_13340,N_13304);
and U13909 (N_13909,N_13414,N_13661);
and U13910 (N_13910,N_13244,N_13384);
nor U13911 (N_13911,N_13193,N_13322);
and U13912 (N_13912,N_13327,N_13569);
nand U13913 (N_13913,N_13258,N_13143);
or U13914 (N_13914,N_13250,N_13713);
or U13915 (N_13915,N_13416,N_13194);
nand U13916 (N_13916,N_13746,N_13446);
or U13917 (N_13917,N_13243,N_13215);
nor U13918 (N_13918,N_13236,N_13241);
xor U13919 (N_13919,N_13640,N_13454);
and U13920 (N_13920,N_13744,N_13339);
or U13921 (N_13921,N_13437,N_13278);
nor U13922 (N_13922,N_13679,N_13145);
and U13923 (N_13923,N_13358,N_13189);
nand U13924 (N_13924,N_13463,N_13269);
or U13925 (N_13925,N_13310,N_13188);
nand U13926 (N_13926,N_13728,N_13297);
and U13927 (N_13927,N_13538,N_13669);
nor U13928 (N_13928,N_13183,N_13702);
xnor U13929 (N_13929,N_13532,N_13690);
and U13930 (N_13930,N_13338,N_13533);
nand U13931 (N_13931,N_13290,N_13647);
and U13932 (N_13932,N_13369,N_13402);
and U13933 (N_13933,N_13688,N_13666);
xor U13934 (N_13934,N_13335,N_13323);
nor U13935 (N_13935,N_13537,N_13492);
nor U13936 (N_13936,N_13523,N_13507);
or U13937 (N_13937,N_13209,N_13280);
nor U13938 (N_13938,N_13351,N_13158);
nand U13939 (N_13939,N_13187,N_13564);
or U13940 (N_13940,N_13232,N_13442);
xor U13941 (N_13941,N_13584,N_13362);
or U13942 (N_13942,N_13251,N_13641);
nor U13943 (N_13943,N_13559,N_13662);
and U13944 (N_13944,N_13729,N_13609);
nand U13945 (N_13945,N_13326,N_13380);
and U13946 (N_13946,N_13553,N_13405);
nand U13947 (N_13947,N_13181,N_13549);
or U13948 (N_13948,N_13709,N_13447);
and U13949 (N_13949,N_13565,N_13284);
xor U13950 (N_13950,N_13685,N_13684);
or U13951 (N_13951,N_13184,N_13424);
or U13952 (N_13952,N_13460,N_13551);
xor U13953 (N_13953,N_13292,N_13510);
nand U13954 (N_13954,N_13635,N_13361);
or U13955 (N_13955,N_13699,N_13573);
nor U13956 (N_13956,N_13478,N_13435);
or U13957 (N_13957,N_13473,N_13436);
nor U13958 (N_13958,N_13422,N_13703);
and U13959 (N_13959,N_13548,N_13527);
xnor U13960 (N_13960,N_13434,N_13376);
xnor U13961 (N_13961,N_13595,N_13494);
and U13962 (N_13962,N_13302,N_13618);
nand U13963 (N_13963,N_13706,N_13225);
and U13964 (N_13964,N_13164,N_13342);
or U13965 (N_13965,N_13163,N_13418);
nor U13966 (N_13966,N_13619,N_13476);
nand U13967 (N_13967,N_13614,N_13205);
and U13968 (N_13968,N_13142,N_13383);
or U13969 (N_13969,N_13562,N_13482);
xnor U13970 (N_13970,N_13509,N_13677);
nor U13971 (N_13971,N_13654,N_13139);
nor U13972 (N_13972,N_13375,N_13396);
nor U13973 (N_13973,N_13212,N_13529);
nor U13974 (N_13974,N_13522,N_13213);
nand U13975 (N_13975,N_13567,N_13291);
nor U13976 (N_13976,N_13355,N_13390);
nor U13977 (N_13977,N_13253,N_13133);
or U13978 (N_13978,N_13735,N_13521);
nand U13979 (N_13979,N_13465,N_13539);
nor U13980 (N_13980,N_13409,N_13514);
nor U13981 (N_13981,N_13185,N_13198);
and U13982 (N_13982,N_13128,N_13611);
nand U13983 (N_13983,N_13415,N_13131);
and U13984 (N_13984,N_13199,N_13712);
and U13985 (N_13985,N_13397,N_13221);
xnor U13986 (N_13986,N_13407,N_13162);
nor U13987 (N_13987,N_13657,N_13592);
xnor U13988 (N_13988,N_13345,N_13161);
nand U13989 (N_13989,N_13497,N_13423);
nand U13990 (N_13990,N_13692,N_13155);
nand U13991 (N_13991,N_13152,N_13132);
xor U13992 (N_13992,N_13456,N_13366);
xnor U13993 (N_13993,N_13591,N_13646);
nor U13994 (N_13994,N_13718,N_13653);
and U13995 (N_13995,N_13289,N_13321);
xor U13996 (N_13996,N_13598,N_13146);
xnor U13997 (N_13997,N_13458,N_13480);
or U13998 (N_13998,N_13541,N_13318);
nor U13999 (N_13999,N_13313,N_13214);
nor U14000 (N_14000,N_13716,N_13673);
nor U14001 (N_14001,N_13737,N_13137);
nand U14002 (N_14002,N_13135,N_13206);
or U14003 (N_14003,N_13365,N_13196);
nand U14004 (N_14004,N_13535,N_13138);
nand U14005 (N_14005,N_13503,N_13432);
nand U14006 (N_14006,N_13440,N_13353);
xnor U14007 (N_14007,N_13455,N_13182);
xnor U14008 (N_14008,N_13372,N_13642);
nor U14009 (N_14009,N_13634,N_13587);
nor U14010 (N_14010,N_13479,N_13233);
and U14011 (N_14011,N_13736,N_13483);
nor U14012 (N_14012,N_13484,N_13731);
or U14013 (N_14013,N_13600,N_13615);
nand U14014 (N_14014,N_13717,N_13201);
or U14015 (N_14015,N_13246,N_13176);
and U14016 (N_14016,N_13504,N_13314);
or U14017 (N_14017,N_13695,N_13501);
nor U14018 (N_14018,N_13378,N_13266);
nand U14019 (N_14019,N_13347,N_13153);
or U14020 (N_14020,N_13582,N_13393);
or U14021 (N_14021,N_13433,N_13606);
or U14022 (N_14022,N_13739,N_13705);
nor U14023 (N_14023,N_13732,N_13599);
and U14024 (N_14024,N_13628,N_13303);
or U14025 (N_14025,N_13307,N_13312);
nor U14026 (N_14026,N_13748,N_13224);
and U14027 (N_14027,N_13445,N_13332);
nor U14028 (N_14028,N_13179,N_13300);
or U14029 (N_14029,N_13357,N_13485);
and U14030 (N_14030,N_13468,N_13273);
xor U14031 (N_14031,N_13360,N_13622);
and U14032 (N_14032,N_13400,N_13336);
nor U14033 (N_14033,N_13687,N_13356);
nor U14034 (N_14034,N_13263,N_13526);
nor U14035 (N_14035,N_13596,N_13180);
nand U14036 (N_14036,N_13547,N_13658);
and U14037 (N_14037,N_13275,N_13417);
xnor U14038 (N_14038,N_13730,N_13438);
or U14039 (N_14039,N_13743,N_13343);
nor U14040 (N_14040,N_13394,N_13665);
or U14041 (N_14041,N_13207,N_13655);
and U14042 (N_14042,N_13328,N_13543);
nor U14043 (N_14043,N_13612,N_13725);
or U14044 (N_14044,N_13371,N_13295);
and U14045 (N_14045,N_13285,N_13368);
xnor U14046 (N_14046,N_13536,N_13505);
and U14047 (N_14047,N_13475,N_13272);
nor U14048 (N_14048,N_13583,N_13453);
or U14049 (N_14049,N_13220,N_13544);
nand U14050 (N_14050,N_13580,N_13561);
nor U14051 (N_14051,N_13707,N_13192);
or U14052 (N_14052,N_13710,N_13130);
or U14053 (N_14053,N_13603,N_13448);
nor U14054 (N_14054,N_13270,N_13239);
nand U14055 (N_14055,N_13555,N_13630);
nand U14056 (N_14056,N_13550,N_13671);
nor U14057 (N_14057,N_13217,N_13621);
xor U14058 (N_14058,N_13643,N_13377);
nand U14059 (N_14059,N_13652,N_13681);
nor U14060 (N_14060,N_13667,N_13245);
nand U14061 (N_14061,N_13672,N_13726);
and U14062 (N_14062,N_13682,N_13388);
xnor U14063 (N_14063,N_13425,N_13157);
xnor U14064 (N_14064,N_13667,N_13295);
or U14065 (N_14065,N_13493,N_13514);
and U14066 (N_14066,N_13138,N_13548);
or U14067 (N_14067,N_13154,N_13445);
and U14068 (N_14068,N_13227,N_13715);
nor U14069 (N_14069,N_13705,N_13125);
and U14070 (N_14070,N_13590,N_13498);
nor U14071 (N_14071,N_13721,N_13726);
and U14072 (N_14072,N_13128,N_13392);
or U14073 (N_14073,N_13360,N_13288);
xor U14074 (N_14074,N_13469,N_13304);
xor U14075 (N_14075,N_13220,N_13704);
nand U14076 (N_14076,N_13587,N_13493);
nor U14077 (N_14077,N_13183,N_13499);
and U14078 (N_14078,N_13195,N_13395);
or U14079 (N_14079,N_13189,N_13152);
nand U14080 (N_14080,N_13470,N_13264);
or U14081 (N_14081,N_13390,N_13741);
or U14082 (N_14082,N_13313,N_13446);
and U14083 (N_14083,N_13277,N_13557);
or U14084 (N_14084,N_13451,N_13425);
or U14085 (N_14085,N_13323,N_13217);
and U14086 (N_14086,N_13351,N_13188);
or U14087 (N_14087,N_13163,N_13649);
nor U14088 (N_14088,N_13518,N_13484);
nor U14089 (N_14089,N_13294,N_13344);
nor U14090 (N_14090,N_13434,N_13654);
nor U14091 (N_14091,N_13661,N_13617);
nor U14092 (N_14092,N_13702,N_13270);
and U14093 (N_14093,N_13186,N_13214);
or U14094 (N_14094,N_13362,N_13209);
nor U14095 (N_14095,N_13219,N_13666);
nor U14096 (N_14096,N_13348,N_13621);
nand U14097 (N_14097,N_13451,N_13240);
or U14098 (N_14098,N_13396,N_13369);
nand U14099 (N_14099,N_13718,N_13397);
and U14100 (N_14100,N_13181,N_13480);
nor U14101 (N_14101,N_13560,N_13472);
and U14102 (N_14102,N_13264,N_13732);
or U14103 (N_14103,N_13280,N_13371);
nand U14104 (N_14104,N_13345,N_13563);
xor U14105 (N_14105,N_13146,N_13580);
nor U14106 (N_14106,N_13450,N_13477);
nand U14107 (N_14107,N_13703,N_13275);
nand U14108 (N_14108,N_13254,N_13727);
nand U14109 (N_14109,N_13133,N_13244);
or U14110 (N_14110,N_13435,N_13222);
xnor U14111 (N_14111,N_13611,N_13162);
nor U14112 (N_14112,N_13218,N_13531);
nand U14113 (N_14113,N_13534,N_13524);
nand U14114 (N_14114,N_13303,N_13341);
and U14115 (N_14115,N_13617,N_13480);
or U14116 (N_14116,N_13153,N_13476);
xor U14117 (N_14117,N_13249,N_13171);
nand U14118 (N_14118,N_13149,N_13215);
xor U14119 (N_14119,N_13141,N_13168);
nand U14120 (N_14120,N_13581,N_13701);
and U14121 (N_14121,N_13586,N_13744);
and U14122 (N_14122,N_13254,N_13643);
and U14123 (N_14123,N_13220,N_13533);
and U14124 (N_14124,N_13531,N_13367);
and U14125 (N_14125,N_13304,N_13536);
nor U14126 (N_14126,N_13230,N_13498);
or U14127 (N_14127,N_13128,N_13593);
nand U14128 (N_14128,N_13205,N_13596);
and U14129 (N_14129,N_13540,N_13621);
or U14130 (N_14130,N_13444,N_13436);
or U14131 (N_14131,N_13681,N_13327);
or U14132 (N_14132,N_13598,N_13484);
or U14133 (N_14133,N_13322,N_13394);
and U14134 (N_14134,N_13693,N_13223);
nor U14135 (N_14135,N_13145,N_13436);
xnor U14136 (N_14136,N_13157,N_13352);
nor U14137 (N_14137,N_13526,N_13705);
xnor U14138 (N_14138,N_13335,N_13183);
nor U14139 (N_14139,N_13715,N_13181);
or U14140 (N_14140,N_13709,N_13416);
xnor U14141 (N_14141,N_13133,N_13450);
nor U14142 (N_14142,N_13430,N_13446);
nor U14143 (N_14143,N_13219,N_13501);
or U14144 (N_14144,N_13578,N_13369);
and U14145 (N_14145,N_13321,N_13197);
nor U14146 (N_14146,N_13296,N_13642);
nor U14147 (N_14147,N_13255,N_13329);
nor U14148 (N_14148,N_13169,N_13666);
and U14149 (N_14149,N_13395,N_13142);
nand U14150 (N_14150,N_13462,N_13696);
nand U14151 (N_14151,N_13378,N_13667);
or U14152 (N_14152,N_13722,N_13207);
nand U14153 (N_14153,N_13388,N_13337);
nand U14154 (N_14154,N_13470,N_13500);
nor U14155 (N_14155,N_13510,N_13362);
and U14156 (N_14156,N_13189,N_13169);
nor U14157 (N_14157,N_13412,N_13229);
and U14158 (N_14158,N_13740,N_13266);
nand U14159 (N_14159,N_13455,N_13745);
nor U14160 (N_14160,N_13532,N_13149);
nand U14161 (N_14161,N_13349,N_13485);
xnor U14162 (N_14162,N_13535,N_13739);
nand U14163 (N_14163,N_13376,N_13530);
or U14164 (N_14164,N_13351,N_13376);
xnor U14165 (N_14165,N_13164,N_13425);
nand U14166 (N_14166,N_13476,N_13392);
or U14167 (N_14167,N_13681,N_13293);
nand U14168 (N_14168,N_13304,N_13339);
xnor U14169 (N_14169,N_13382,N_13244);
nand U14170 (N_14170,N_13650,N_13240);
xor U14171 (N_14171,N_13384,N_13248);
or U14172 (N_14172,N_13529,N_13579);
nand U14173 (N_14173,N_13478,N_13523);
and U14174 (N_14174,N_13229,N_13508);
nand U14175 (N_14175,N_13291,N_13481);
xor U14176 (N_14176,N_13166,N_13268);
nor U14177 (N_14177,N_13358,N_13636);
and U14178 (N_14178,N_13450,N_13624);
or U14179 (N_14179,N_13481,N_13730);
nor U14180 (N_14180,N_13391,N_13620);
and U14181 (N_14181,N_13433,N_13496);
nand U14182 (N_14182,N_13606,N_13649);
nand U14183 (N_14183,N_13669,N_13245);
or U14184 (N_14184,N_13249,N_13435);
nand U14185 (N_14185,N_13382,N_13257);
nand U14186 (N_14186,N_13617,N_13317);
or U14187 (N_14187,N_13606,N_13362);
and U14188 (N_14188,N_13228,N_13433);
or U14189 (N_14189,N_13335,N_13740);
and U14190 (N_14190,N_13528,N_13353);
nand U14191 (N_14191,N_13607,N_13168);
nor U14192 (N_14192,N_13686,N_13495);
xnor U14193 (N_14193,N_13146,N_13362);
xnor U14194 (N_14194,N_13490,N_13488);
nor U14195 (N_14195,N_13651,N_13198);
or U14196 (N_14196,N_13690,N_13595);
or U14197 (N_14197,N_13195,N_13554);
nor U14198 (N_14198,N_13211,N_13744);
nor U14199 (N_14199,N_13493,N_13180);
nor U14200 (N_14200,N_13641,N_13358);
xor U14201 (N_14201,N_13614,N_13716);
and U14202 (N_14202,N_13721,N_13160);
nand U14203 (N_14203,N_13513,N_13663);
nor U14204 (N_14204,N_13483,N_13156);
and U14205 (N_14205,N_13224,N_13182);
and U14206 (N_14206,N_13695,N_13340);
or U14207 (N_14207,N_13350,N_13379);
or U14208 (N_14208,N_13481,N_13394);
nor U14209 (N_14209,N_13534,N_13206);
or U14210 (N_14210,N_13569,N_13559);
or U14211 (N_14211,N_13160,N_13579);
nand U14212 (N_14212,N_13269,N_13564);
and U14213 (N_14213,N_13273,N_13242);
and U14214 (N_14214,N_13404,N_13527);
and U14215 (N_14215,N_13240,N_13468);
nor U14216 (N_14216,N_13183,N_13738);
and U14217 (N_14217,N_13332,N_13426);
and U14218 (N_14218,N_13595,N_13370);
xnor U14219 (N_14219,N_13699,N_13575);
nor U14220 (N_14220,N_13734,N_13676);
nor U14221 (N_14221,N_13591,N_13195);
nor U14222 (N_14222,N_13383,N_13391);
xnor U14223 (N_14223,N_13527,N_13346);
nand U14224 (N_14224,N_13155,N_13217);
and U14225 (N_14225,N_13386,N_13441);
and U14226 (N_14226,N_13409,N_13488);
nand U14227 (N_14227,N_13185,N_13236);
nand U14228 (N_14228,N_13656,N_13319);
nor U14229 (N_14229,N_13428,N_13396);
xor U14230 (N_14230,N_13518,N_13387);
xor U14231 (N_14231,N_13281,N_13178);
or U14232 (N_14232,N_13315,N_13622);
and U14233 (N_14233,N_13582,N_13374);
nor U14234 (N_14234,N_13516,N_13227);
nor U14235 (N_14235,N_13437,N_13643);
or U14236 (N_14236,N_13499,N_13719);
and U14237 (N_14237,N_13654,N_13601);
nand U14238 (N_14238,N_13468,N_13578);
nor U14239 (N_14239,N_13626,N_13483);
or U14240 (N_14240,N_13603,N_13715);
nor U14241 (N_14241,N_13426,N_13654);
and U14242 (N_14242,N_13436,N_13413);
or U14243 (N_14243,N_13272,N_13151);
or U14244 (N_14244,N_13440,N_13697);
nor U14245 (N_14245,N_13595,N_13217);
nand U14246 (N_14246,N_13367,N_13515);
or U14247 (N_14247,N_13200,N_13385);
or U14248 (N_14248,N_13627,N_13561);
nor U14249 (N_14249,N_13577,N_13386);
nor U14250 (N_14250,N_13443,N_13475);
nor U14251 (N_14251,N_13364,N_13169);
and U14252 (N_14252,N_13490,N_13315);
or U14253 (N_14253,N_13608,N_13212);
or U14254 (N_14254,N_13237,N_13575);
and U14255 (N_14255,N_13661,N_13627);
or U14256 (N_14256,N_13528,N_13381);
and U14257 (N_14257,N_13547,N_13536);
nand U14258 (N_14258,N_13475,N_13657);
xnor U14259 (N_14259,N_13342,N_13670);
xor U14260 (N_14260,N_13729,N_13182);
nor U14261 (N_14261,N_13316,N_13628);
nor U14262 (N_14262,N_13482,N_13716);
nor U14263 (N_14263,N_13237,N_13557);
or U14264 (N_14264,N_13371,N_13199);
and U14265 (N_14265,N_13140,N_13531);
nand U14266 (N_14266,N_13668,N_13443);
nand U14267 (N_14267,N_13512,N_13497);
nand U14268 (N_14268,N_13611,N_13518);
or U14269 (N_14269,N_13738,N_13643);
or U14270 (N_14270,N_13128,N_13579);
or U14271 (N_14271,N_13260,N_13337);
nor U14272 (N_14272,N_13512,N_13676);
and U14273 (N_14273,N_13331,N_13475);
or U14274 (N_14274,N_13398,N_13575);
or U14275 (N_14275,N_13301,N_13216);
or U14276 (N_14276,N_13173,N_13341);
or U14277 (N_14277,N_13510,N_13466);
nand U14278 (N_14278,N_13330,N_13196);
or U14279 (N_14279,N_13718,N_13406);
or U14280 (N_14280,N_13442,N_13321);
and U14281 (N_14281,N_13386,N_13408);
xnor U14282 (N_14282,N_13596,N_13339);
xor U14283 (N_14283,N_13318,N_13172);
nor U14284 (N_14284,N_13409,N_13226);
and U14285 (N_14285,N_13492,N_13244);
nand U14286 (N_14286,N_13617,N_13421);
or U14287 (N_14287,N_13254,N_13286);
or U14288 (N_14288,N_13666,N_13476);
nor U14289 (N_14289,N_13237,N_13529);
and U14290 (N_14290,N_13295,N_13716);
nor U14291 (N_14291,N_13300,N_13666);
xor U14292 (N_14292,N_13275,N_13366);
and U14293 (N_14293,N_13708,N_13399);
xor U14294 (N_14294,N_13205,N_13310);
nand U14295 (N_14295,N_13664,N_13568);
nand U14296 (N_14296,N_13512,N_13468);
and U14297 (N_14297,N_13321,N_13393);
nand U14298 (N_14298,N_13333,N_13146);
or U14299 (N_14299,N_13309,N_13389);
nand U14300 (N_14300,N_13274,N_13324);
nor U14301 (N_14301,N_13217,N_13639);
or U14302 (N_14302,N_13372,N_13616);
nor U14303 (N_14303,N_13257,N_13711);
and U14304 (N_14304,N_13742,N_13427);
and U14305 (N_14305,N_13492,N_13310);
nor U14306 (N_14306,N_13517,N_13484);
and U14307 (N_14307,N_13744,N_13163);
or U14308 (N_14308,N_13170,N_13144);
nor U14309 (N_14309,N_13724,N_13583);
and U14310 (N_14310,N_13393,N_13548);
nor U14311 (N_14311,N_13153,N_13504);
or U14312 (N_14312,N_13348,N_13467);
xnor U14313 (N_14313,N_13498,N_13602);
xnor U14314 (N_14314,N_13218,N_13193);
nand U14315 (N_14315,N_13423,N_13645);
nand U14316 (N_14316,N_13610,N_13581);
and U14317 (N_14317,N_13396,N_13216);
or U14318 (N_14318,N_13586,N_13222);
nand U14319 (N_14319,N_13458,N_13431);
nor U14320 (N_14320,N_13688,N_13542);
or U14321 (N_14321,N_13151,N_13653);
nor U14322 (N_14322,N_13576,N_13353);
xor U14323 (N_14323,N_13419,N_13343);
xnor U14324 (N_14324,N_13508,N_13487);
and U14325 (N_14325,N_13512,N_13473);
or U14326 (N_14326,N_13576,N_13493);
nand U14327 (N_14327,N_13479,N_13627);
nor U14328 (N_14328,N_13381,N_13543);
nor U14329 (N_14329,N_13144,N_13515);
nor U14330 (N_14330,N_13741,N_13199);
xor U14331 (N_14331,N_13232,N_13386);
or U14332 (N_14332,N_13313,N_13697);
nand U14333 (N_14333,N_13451,N_13158);
or U14334 (N_14334,N_13305,N_13209);
and U14335 (N_14335,N_13350,N_13591);
nand U14336 (N_14336,N_13487,N_13140);
nand U14337 (N_14337,N_13397,N_13464);
nand U14338 (N_14338,N_13639,N_13592);
nand U14339 (N_14339,N_13464,N_13514);
nand U14340 (N_14340,N_13697,N_13333);
nand U14341 (N_14341,N_13263,N_13570);
xor U14342 (N_14342,N_13281,N_13286);
and U14343 (N_14343,N_13738,N_13165);
nand U14344 (N_14344,N_13426,N_13304);
or U14345 (N_14345,N_13200,N_13542);
or U14346 (N_14346,N_13619,N_13284);
nor U14347 (N_14347,N_13197,N_13500);
nand U14348 (N_14348,N_13485,N_13244);
or U14349 (N_14349,N_13674,N_13226);
nor U14350 (N_14350,N_13340,N_13134);
nor U14351 (N_14351,N_13529,N_13556);
xnor U14352 (N_14352,N_13168,N_13177);
and U14353 (N_14353,N_13375,N_13147);
nor U14354 (N_14354,N_13505,N_13702);
and U14355 (N_14355,N_13208,N_13679);
or U14356 (N_14356,N_13480,N_13510);
nor U14357 (N_14357,N_13647,N_13662);
or U14358 (N_14358,N_13351,N_13613);
and U14359 (N_14359,N_13462,N_13425);
or U14360 (N_14360,N_13138,N_13609);
nand U14361 (N_14361,N_13237,N_13396);
nor U14362 (N_14362,N_13536,N_13401);
nand U14363 (N_14363,N_13701,N_13532);
nand U14364 (N_14364,N_13680,N_13158);
and U14365 (N_14365,N_13700,N_13252);
xor U14366 (N_14366,N_13189,N_13323);
or U14367 (N_14367,N_13341,N_13513);
nor U14368 (N_14368,N_13640,N_13191);
nor U14369 (N_14369,N_13552,N_13159);
or U14370 (N_14370,N_13308,N_13257);
xor U14371 (N_14371,N_13157,N_13428);
or U14372 (N_14372,N_13626,N_13719);
and U14373 (N_14373,N_13241,N_13538);
nand U14374 (N_14374,N_13310,N_13181);
nand U14375 (N_14375,N_14304,N_14129);
and U14376 (N_14376,N_13873,N_13954);
nor U14377 (N_14377,N_14124,N_14121);
or U14378 (N_14378,N_14007,N_14148);
nand U14379 (N_14379,N_13958,N_14293);
xor U14380 (N_14380,N_14239,N_14101);
nand U14381 (N_14381,N_14335,N_13939);
xnor U14382 (N_14382,N_14256,N_13844);
nor U14383 (N_14383,N_14282,N_13962);
nand U14384 (N_14384,N_14050,N_14104);
or U14385 (N_14385,N_14296,N_13922);
nand U14386 (N_14386,N_14230,N_14283);
nand U14387 (N_14387,N_14057,N_14082);
and U14388 (N_14388,N_13854,N_14126);
and U14389 (N_14389,N_13918,N_13864);
and U14390 (N_14390,N_13911,N_13879);
and U14391 (N_14391,N_14180,N_13969);
nand U14392 (N_14392,N_14088,N_14317);
and U14393 (N_14393,N_13915,N_14292);
nor U14394 (N_14394,N_13941,N_13995);
or U14395 (N_14395,N_13838,N_13887);
nor U14396 (N_14396,N_13874,N_14300);
nand U14397 (N_14397,N_14345,N_14172);
xnor U14398 (N_14398,N_13779,N_13920);
and U14399 (N_14399,N_14078,N_13999);
nand U14400 (N_14400,N_14095,N_13947);
nor U14401 (N_14401,N_13866,N_13908);
or U14402 (N_14402,N_14086,N_13778);
or U14403 (N_14403,N_14175,N_14374);
and U14404 (N_14404,N_13896,N_14331);
xor U14405 (N_14405,N_14062,N_14307);
nor U14406 (N_14406,N_14333,N_13913);
nand U14407 (N_14407,N_13974,N_13897);
nor U14408 (N_14408,N_13830,N_13891);
nand U14409 (N_14409,N_14272,N_14193);
and U14410 (N_14410,N_14259,N_14246);
nand U14411 (N_14411,N_14368,N_14211);
nor U14412 (N_14412,N_13878,N_14109);
or U14413 (N_14413,N_14102,N_13968);
or U14414 (N_14414,N_14045,N_14092);
or U14415 (N_14415,N_14264,N_14159);
and U14416 (N_14416,N_13814,N_14116);
nand U14417 (N_14417,N_14155,N_13919);
and U14418 (N_14418,N_14027,N_14228);
nand U14419 (N_14419,N_13867,N_14357);
or U14420 (N_14420,N_14332,N_14015);
nand U14421 (N_14421,N_13776,N_14318);
xnor U14422 (N_14422,N_14373,N_14360);
nor U14423 (N_14423,N_14367,N_14218);
xnor U14424 (N_14424,N_13817,N_14067);
xnor U14425 (N_14425,N_14149,N_14139);
xnor U14426 (N_14426,N_13893,N_14217);
nor U14427 (N_14427,N_14053,N_14080);
and U14428 (N_14428,N_14182,N_14079);
and U14429 (N_14429,N_14094,N_14163);
nor U14430 (N_14430,N_14351,N_13860);
nor U14431 (N_14431,N_14209,N_13957);
xnor U14432 (N_14432,N_14023,N_13925);
and U14433 (N_14433,N_14251,N_14359);
nor U14434 (N_14434,N_13934,N_13903);
or U14435 (N_14435,N_14096,N_14236);
and U14436 (N_14436,N_14261,N_13890);
and U14437 (N_14437,N_14347,N_14018);
nand U14438 (N_14438,N_14137,N_13805);
nand U14439 (N_14439,N_14036,N_13886);
nand U14440 (N_14440,N_14299,N_14042);
or U14441 (N_14441,N_13998,N_13952);
nand U14442 (N_14442,N_14221,N_13754);
xnor U14443 (N_14443,N_13950,N_13948);
nor U14444 (N_14444,N_14321,N_13807);
nor U14445 (N_14445,N_13985,N_14074);
and U14446 (N_14446,N_14201,N_14103);
nor U14447 (N_14447,N_13983,N_14302);
nand U14448 (N_14448,N_14028,N_13956);
nor U14449 (N_14449,N_14213,N_13976);
xor U14450 (N_14450,N_13883,N_13964);
or U14451 (N_14451,N_13765,N_14242);
and U14452 (N_14452,N_14122,N_13912);
or U14453 (N_14453,N_14111,N_13764);
nand U14454 (N_14454,N_14198,N_13872);
and U14455 (N_14455,N_14058,N_13851);
nand U14456 (N_14456,N_14108,N_14268);
xnor U14457 (N_14457,N_13986,N_14248);
or U14458 (N_14458,N_14269,N_13882);
or U14459 (N_14459,N_13822,N_13837);
nand U14460 (N_14460,N_13780,N_13823);
nand U14461 (N_14461,N_13931,N_13933);
nor U14462 (N_14462,N_13752,N_13810);
and U14463 (N_14463,N_14176,N_13877);
nor U14464 (N_14464,N_13953,N_13875);
nand U14465 (N_14465,N_14305,N_13800);
xnor U14466 (N_14466,N_13813,N_14289);
xor U14467 (N_14467,N_14140,N_13768);
nand U14468 (N_14468,N_14056,N_14308);
nand U14469 (N_14469,N_13771,N_13761);
or U14470 (N_14470,N_14195,N_14255);
and U14471 (N_14471,N_14219,N_14278);
nand U14472 (N_14472,N_14224,N_14090);
nand U14473 (N_14473,N_13816,N_14130);
and U14474 (N_14474,N_13812,N_14098);
nand U14475 (N_14475,N_14136,N_14310);
or U14476 (N_14476,N_14047,N_14273);
or U14477 (N_14477,N_13781,N_13782);
nand U14478 (N_14478,N_13892,N_14006);
or U14479 (N_14479,N_13839,N_14105);
nand U14480 (N_14480,N_14110,N_14059);
nand U14481 (N_14481,N_13898,N_13824);
xnor U14482 (N_14482,N_13905,N_13990);
nor U14483 (N_14483,N_14004,N_14340);
nand U14484 (N_14484,N_14014,N_13929);
and U14485 (N_14485,N_14189,N_13930);
or U14486 (N_14486,N_13856,N_14235);
and U14487 (N_14487,N_13815,N_13750);
and U14488 (N_14488,N_13785,N_14324);
xnor U14489 (N_14489,N_14348,N_14026);
nand U14490 (N_14490,N_14156,N_14019);
or U14491 (N_14491,N_13993,N_14069);
xnor U14492 (N_14492,N_13804,N_14052);
or U14493 (N_14493,N_14084,N_14190);
xnor U14494 (N_14494,N_13827,N_13869);
nand U14495 (N_14495,N_13787,N_14133);
nand U14496 (N_14496,N_14070,N_14257);
nor U14497 (N_14497,N_13861,N_13806);
or U14498 (N_14498,N_14303,N_13840);
or U14499 (N_14499,N_14134,N_13858);
nor U14500 (N_14500,N_14097,N_13826);
nor U14501 (N_14501,N_14187,N_13820);
nor U14502 (N_14502,N_14112,N_13944);
nor U14503 (N_14503,N_14286,N_14337);
nor U14504 (N_14504,N_14055,N_13759);
nor U14505 (N_14505,N_14280,N_13819);
or U14506 (N_14506,N_13794,N_13799);
and U14507 (N_14507,N_14284,N_13997);
or U14508 (N_14508,N_13862,N_13756);
nand U14509 (N_14509,N_13849,N_14087);
xnor U14510 (N_14510,N_14362,N_14358);
nand U14511 (N_14511,N_14154,N_13783);
and U14512 (N_14512,N_13901,N_13921);
or U14513 (N_14513,N_14035,N_14285);
nand U14514 (N_14514,N_14295,N_14234);
nor U14515 (N_14515,N_13766,N_14250);
nand U14516 (N_14516,N_14263,N_13841);
or U14517 (N_14517,N_13889,N_13899);
or U14518 (N_14518,N_14326,N_14008);
nand U14519 (N_14519,N_14244,N_14115);
nor U14520 (N_14520,N_13751,N_13885);
and U14521 (N_14521,N_14290,N_14147);
and U14522 (N_14522,N_14298,N_14165);
or U14523 (N_14523,N_13763,N_13834);
and U14524 (N_14524,N_14204,N_13907);
nand U14525 (N_14525,N_14071,N_13963);
and U14526 (N_14526,N_14085,N_14021);
or U14527 (N_14527,N_14162,N_14060);
nand U14528 (N_14528,N_13973,N_14150);
or U14529 (N_14529,N_14033,N_14229);
nand U14530 (N_14530,N_14031,N_13792);
or U14531 (N_14531,N_13847,N_14089);
nand U14532 (N_14532,N_14314,N_14107);
or U14533 (N_14533,N_14178,N_14081);
and U14534 (N_14534,N_14334,N_14046);
nand U14535 (N_14535,N_13857,N_13972);
nor U14536 (N_14536,N_14179,N_13788);
or U14537 (N_14537,N_14000,N_14157);
and U14538 (N_14538,N_13829,N_13888);
nor U14539 (N_14539,N_13832,N_13987);
nand U14540 (N_14540,N_14312,N_13960);
nand U14541 (N_14541,N_14322,N_14048);
and U14542 (N_14542,N_14186,N_13865);
and U14543 (N_14543,N_13965,N_14016);
xor U14544 (N_14544,N_14181,N_14311);
and U14545 (N_14545,N_14350,N_13977);
nand U14546 (N_14546,N_14044,N_13932);
and U14547 (N_14547,N_14313,N_14301);
nand U14548 (N_14548,N_14241,N_14315);
or U14549 (N_14549,N_14353,N_14005);
and U14550 (N_14550,N_14215,N_13846);
or U14551 (N_14551,N_13876,N_14169);
and U14552 (N_14552,N_14316,N_14275);
nand U14553 (N_14553,N_13916,N_14338);
or U14554 (N_14554,N_14151,N_13845);
and U14555 (N_14555,N_14200,N_14064);
and U14556 (N_14556,N_14166,N_13828);
or U14557 (N_14557,N_14063,N_13762);
and U14558 (N_14558,N_13802,N_13809);
and U14559 (N_14559,N_13786,N_14135);
or U14560 (N_14560,N_14002,N_13970);
nand U14561 (N_14561,N_13818,N_14131);
or U14562 (N_14562,N_14168,N_14363);
nand U14563 (N_14563,N_14142,N_14127);
nor U14564 (N_14564,N_14223,N_14254);
xnor U14565 (N_14565,N_14065,N_13910);
and U14566 (N_14566,N_13902,N_14011);
nor U14567 (N_14567,N_14017,N_13803);
and U14568 (N_14568,N_13961,N_13852);
or U14569 (N_14569,N_13855,N_14029);
nor U14570 (N_14570,N_14329,N_13955);
or U14571 (N_14571,N_14106,N_14153);
nor U14572 (N_14572,N_14207,N_13784);
or U14573 (N_14573,N_14197,N_13774);
and U14574 (N_14574,N_13797,N_14212);
or U14575 (N_14575,N_14328,N_14342);
xor U14576 (N_14576,N_13757,N_13940);
nor U14577 (N_14577,N_14076,N_14346);
nand U14578 (N_14578,N_14114,N_13789);
nand U14579 (N_14579,N_13831,N_14274);
and U14580 (N_14580,N_13917,N_14253);
nor U14581 (N_14581,N_14199,N_13909);
and U14582 (N_14582,N_14262,N_14291);
or U14583 (N_14583,N_14245,N_13796);
and U14584 (N_14584,N_14012,N_14355);
and U14585 (N_14585,N_14309,N_13980);
nand U14586 (N_14586,N_13880,N_14267);
xor U14587 (N_14587,N_13871,N_13906);
and U14588 (N_14588,N_13870,N_14352);
nor U14589 (N_14589,N_13791,N_14206);
nor U14590 (N_14590,N_13801,N_14222);
and U14591 (N_14591,N_14361,N_14349);
or U14592 (N_14592,N_14024,N_14191);
nand U14593 (N_14593,N_13811,N_14184);
nand U14594 (N_14594,N_13975,N_14039);
or U14595 (N_14595,N_14226,N_14160);
xnor U14596 (N_14596,N_14073,N_13863);
or U14597 (N_14597,N_14225,N_14123);
nand U14598 (N_14598,N_14049,N_14339);
nand U14599 (N_14599,N_14022,N_13971);
nor U14600 (N_14600,N_13966,N_14161);
and U14601 (N_14601,N_14214,N_13842);
xor U14602 (N_14602,N_14306,N_14077);
and U14603 (N_14603,N_14054,N_14281);
or U14604 (N_14604,N_14118,N_14192);
xnor U14605 (N_14605,N_14132,N_14243);
xnor U14606 (N_14606,N_14158,N_13798);
nand U14607 (N_14607,N_14287,N_14010);
or U14608 (N_14608,N_14091,N_14227);
nand U14609 (N_14609,N_14083,N_14037);
xor U14610 (N_14610,N_14003,N_13914);
nand U14611 (N_14611,N_13937,N_13758);
nand U14612 (N_14612,N_14075,N_14117);
nand U14613 (N_14613,N_13943,N_14113);
nand U14614 (N_14614,N_14320,N_13978);
and U14615 (N_14615,N_13949,N_14194);
nor U14616 (N_14616,N_14277,N_14068);
or U14617 (N_14617,N_14143,N_14266);
nor U14618 (N_14618,N_13760,N_14208);
nor U14619 (N_14619,N_13996,N_13992);
nor U14620 (N_14620,N_14258,N_14043);
nand U14621 (N_14621,N_14041,N_13859);
and U14622 (N_14622,N_14040,N_14120);
nand U14623 (N_14623,N_14001,N_13843);
or U14624 (N_14624,N_13923,N_14364);
and U14625 (N_14625,N_14119,N_14174);
nand U14626 (N_14626,N_13848,N_14188);
nor U14627 (N_14627,N_13994,N_14128);
or U14628 (N_14628,N_13755,N_14249);
nand U14629 (N_14629,N_13790,N_14330);
and U14630 (N_14630,N_13772,N_13770);
nand U14631 (N_14631,N_14196,N_13926);
xnor U14632 (N_14632,N_13938,N_14270);
xor U14633 (N_14633,N_14252,N_13981);
nand U14634 (N_14634,N_13989,N_13900);
nand U14635 (N_14635,N_14323,N_14297);
or U14636 (N_14636,N_13825,N_14237);
or U14637 (N_14637,N_13894,N_14288);
nor U14638 (N_14638,N_13821,N_14051);
nor U14639 (N_14639,N_13936,N_13753);
or U14640 (N_14640,N_13904,N_14372);
nand U14641 (N_14641,N_14185,N_14173);
nor U14642 (N_14642,N_14265,N_14240);
or U14643 (N_14643,N_14205,N_14232);
xor U14644 (N_14644,N_14145,N_14276);
nor U14645 (N_14645,N_13988,N_14325);
or U14646 (N_14646,N_14152,N_13850);
nand U14647 (N_14647,N_14013,N_14370);
nor U14648 (N_14648,N_14354,N_13984);
and U14649 (N_14649,N_13775,N_14009);
or U14650 (N_14650,N_14167,N_14341);
or U14651 (N_14651,N_13979,N_14260);
and U14652 (N_14652,N_13945,N_14099);
xnor U14653 (N_14653,N_13927,N_14279);
nand U14654 (N_14654,N_14170,N_14327);
nor U14655 (N_14655,N_14138,N_13959);
or U14656 (N_14656,N_14038,N_14141);
nor U14657 (N_14657,N_13793,N_14210);
or U14658 (N_14658,N_13777,N_14343);
or U14659 (N_14659,N_14025,N_14072);
xnor U14660 (N_14660,N_13895,N_14032);
nand U14661 (N_14661,N_13836,N_14271);
nor U14662 (N_14662,N_13769,N_13808);
and U14663 (N_14663,N_13773,N_13924);
and U14664 (N_14664,N_14231,N_14164);
nor U14665 (N_14665,N_14177,N_14203);
nor U14666 (N_14666,N_14146,N_14220);
and U14667 (N_14667,N_14202,N_14066);
nor U14668 (N_14668,N_14366,N_13928);
or U14669 (N_14669,N_13884,N_13946);
nor U14670 (N_14670,N_13951,N_14247);
xor U14671 (N_14671,N_13967,N_14125);
and U14672 (N_14672,N_13942,N_14319);
nor U14673 (N_14673,N_14144,N_14030);
nand U14674 (N_14674,N_13795,N_14356);
nor U14675 (N_14675,N_14369,N_14034);
nand U14676 (N_14676,N_14100,N_14061);
or U14677 (N_14677,N_14238,N_14371);
xnor U14678 (N_14678,N_14365,N_13991);
nand U14679 (N_14679,N_13982,N_13935);
nand U14680 (N_14680,N_14294,N_14020);
and U14681 (N_14681,N_14336,N_13835);
nand U14682 (N_14682,N_13833,N_14233);
and U14683 (N_14683,N_14216,N_13881);
nor U14684 (N_14684,N_13853,N_14183);
nor U14685 (N_14685,N_13868,N_14344);
nand U14686 (N_14686,N_13767,N_14093);
and U14687 (N_14687,N_14171,N_14137);
xnor U14688 (N_14688,N_13831,N_13882);
or U14689 (N_14689,N_14059,N_14347);
and U14690 (N_14690,N_14172,N_14043);
xor U14691 (N_14691,N_13922,N_13992);
and U14692 (N_14692,N_13796,N_13913);
or U14693 (N_14693,N_14240,N_13878);
or U14694 (N_14694,N_14100,N_14373);
nand U14695 (N_14695,N_14037,N_14103);
nand U14696 (N_14696,N_13756,N_14353);
or U14697 (N_14697,N_14057,N_13940);
nor U14698 (N_14698,N_13870,N_14235);
and U14699 (N_14699,N_13841,N_14311);
and U14700 (N_14700,N_13759,N_13783);
or U14701 (N_14701,N_13948,N_13791);
xor U14702 (N_14702,N_13833,N_14125);
or U14703 (N_14703,N_14272,N_13794);
nor U14704 (N_14704,N_14340,N_13983);
or U14705 (N_14705,N_13943,N_14288);
xnor U14706 (N_14706,N_14065,N_13886);
and U14707 (N_14707,N_13871,N_13916);
nor U14708 (N_14708,N_14119,N_13928);
nor U14709 (N_14709,N_14286,N_14238);
and U14710 (N_14710,N_14017,N_14374);
nor U14711 (N_14711,N_14271,N_14145);
and U14712 (N_14712,N_13977,N_14052);
or U14713 (N_14713,N_14175,N_14030);
and U14714 (N_14714,N_13861,N_13820);
or U14715 (N_14715,N_14307,N_13848);
or U14716 (N_14716,N_13869,N_13844);
nand U14717 (N_14717,N_13833,N_14187);
nor U14718 (N_14718,N_13953,N_14220);
xor U14719 (N_14719,N_14274,N_14120);
xnor U14720 (N_14720,N_13992,N_14095);
nand U14721 (N_14721,N_13896,N_14239);
nand U14722 (N_14722,N_14194,N_14028);
nor U14723 (N_14723,N_13934,N_14029);
nor U14724 (N_14724,N_13817,N_14113);
nor U14725 (N_14725,N_14337,N_14016);
and U14726 (N_14726,N_13983,N_13997);
nor U14727 (N_14727,N_14315,N_14000);
and U14728 (N_14728,N_13759,N_13875);
nand U14729 (N_14729,N_14370,N_13820);
nand U14730 (N_14730,N_14172,N_14341);
xnor U14731 (N_14731,N_13949,N_14343);
and U14732 (N_14732,N_14251,N_13917);
xor U14733 (N_14733,N_14355,N_13774);
and U14734 (N_14734,N_14070,N_13839);
nand U14735 (N_14735,N_14238,N_13779);
nor U14736 (N_14736,N_13832,N_13984);
nand U14737 (N_14737,N_14061,N_13937);
nand U14738 (N_14738,N_13933,N_14258);
nor U14739 (N_14739,N_13795,N_13781);
nand U14740 (N_14740,N_13956,N_14371);
nand U14741 (N_14741,N_14105,N_14083);
and U14742 (N_14742,N_13855,N_14301);
nand U14743 (N_14743,N_14037,N_14260);
or U14744 (N_14744,N_14159,N_13826);
nand U14745 (N_14745,N_13929,N_13785);
and U14746 (N_14746,N_14088,N_14120);
xor U14747 (N_14747,N_13900,N_14086);
nand U14748 (N_14748,N_14185,N_14099);
nand U14749 (N_14749,N_14210,N_14203);
or U14750 (N_14750,N_13990,N_13892);
nor U14751 (N_14751,N_14149,N_14278);
or U14752 (N_14752,N_13856,N_13807);
xor U14753 (N_14753,N_13804,N_13928);
xor U14754 (N_14754,N_13926,N_13869);
nand U14755 (N_14755,N_13903,N_14038);
or U14756 (N_14756,N_13895,N_13795);
xnor U14757 (N_14757,N_13952,N_14270);
or U14758 (N_14758,N_14290,N_13783);
nor U14759 (N_14759,N_14006,N_14299);
nand U14760 (N_14760,N_14291,N_14252);
or U14761 (N_14761,N_14176,N_14340);
and U14762 (N_14762,N_14186,N_13921);
and U14763 (N_14763,N_14324,N_14219);
or U14764 (N_14764,N_14217,N_13900);
nand U14765 (N_14765,N_13917,N_13926);
and U14766 (N_14766,N_13884,N_14362);
xor U14767 (N_14767,N_14080,N_14099);
or U14768 (N_14768,N_13862,N_14117);
or U14769 (N_14769,N_14066,N_14369);
nor U14770 (N_14770,N_14048,N_14141);
or U14771 (N_14771,N_13927,N_14086);
nor U14772 (N_14772,N_14196,N_13783);
nand U14773 (N_14773,N_14229,N_14058);
nand U14774 (N_14774,N_14029,N_13757);
and U14775 (N_14775,N_13939,N_14229);
and U14776 (N_14776,N_14021,N_14263);
and U14777 (N_14777,N_14150,N_13964);
or U14778 (N_14778,N_13945,N_14259);
or U14779 (N_14779,N_14153,N_14146);
or U14780 (N_14780,N_14222,N_14048);
nand U14781 (N_14781,N_13930,N_14159);
xnor U14782 (N_14782,N_14257,N_14044);
nor U14783 (N_14783,N_14226,N_13865);
or U14784 (N_14784,N_14334,N_14277);
and U14785 (N_14785,N_13889,N_14200);
xor U14786 (N_14786,N_13948,N_14213);
and U14787 (N_14787,N_13879,N_13787);
and U14788 (N_14788,N_14274,N_13938);
nor U14789 (N_14789,N_13897,N_14132);
nand U14790 (N_14790,N_13956,N_14200);
nor U14791 (N_14791,N_13861,N_14007);
or U14792 (N_14792,N_14092,N_13932);
and U14793 (N_14793,N_14108,N_14010);
nand U14794 (N_14794,N_13786,N_14174);
nand U14795 (N_14795,N_13805,N_14028);
nand U14796 (N_14796,N_14128,N_14268);
nor U14797 (N_14797,N_14059,N_14267);
nor U14798 (N_14798,N_14205,N_14272);
xnor U14799 (N_14799,N_13947,N_14109);
nand U14800 (N_14800,N_13956,N_13921);
nor U14801 (N_14801,N_13805,N_14325);
or U14802 (N_14802,N_14179,N_13899);
or U14803 (N_14803,N_14011,N_13828);
xnor U14804 (N_14804,N_14290,N_14106);
or U14805 (N_14805,N_13842,N_14210);
and U14806 (N_14806,N_14088,N_14069);
nand U14807 (N_14807,N_14239,N_14123);
or U14808 (N_14808,N_14182,N_14333);
and U14809 (N_14809,N_14374,N_14077);
nor U14810 (N_14810,N_14300,N_14273);
nor U14811 (N_14811,N_13756,N_14277);
or U14812 (N_14812,N_13859,N_13908);
or U14813 (N_14813,N_14347,N_14071);
and U14814 (N_14814,N_14245,N_14303);
and U14815 (N_14815,N_14183,N_13872);
or U14816 (N_14816,N_13857,N_14253);
nand U14817 (N_14817,N_13752,N_13800);
nor U14818 (N_14818,N_14060,N_14017);
xnor U14819 (N_14819,N_14113,N_13956);
nor U14820 (N_14820,N_13987,N_14258);
nor U14821 (N_14821,N_14072,N_14214);
and U14822 (N_14822,N_14116,N_14283);
and U14823 (N_14823,N_14135,N_14232);
nand U14824 (N_14824,N_14311,N_14178);
nor U14825 (N_14825,N_14225,N_14199);
nand U14826 (N_14826,N_14165,N_13944);
or U14827 (N_14827,N_13771,N_14193);
and U14828 (N_14828,N_14040,N_14316);
nand U14829 (N_14829,N_13924,N_13838);
and U14830 (N_14830,N_14332,N_13978);
and U14831 (N_14831,N_14255,N_13970);
xnor U14832 (N_14832,N_13949,N_14132);
nand U14833 (N_14833,N_14110,N_13911);
and U14834 (N_14834,N_14283,N_13902);
nand U14835 (N_14835,N_14239,N_14181);
nor U14836 (N_14836,N_14139,N_14162);
nand U14837 (N_14837,N_13848,N_14257);
xnor U14838 (N_14838,N_14006,N_13772);
nand U14839 (N_14839,N_14152,N_13953);
and U14840 (N_14840,N_14031,N_13977);
nand U14841 (N_14841,N_14181,N_14039);
nand U14842 (N_14842,N_13842,N_14147);
or U14843 (N_14843,N_13856,N_14298);
nand U14844 (N_14844,N_14149,N_14147);
nor U14845 (N_14845,N_13752,N_13957);
and U14846 (N_14846,N_14325,N_14135);
nand U14847 (N_14847,N_14256,N_13803);
xnor U14848 (N_14848,N_14031,N_13803);
nand U14849 (N_14849,N_13812,N_14368);
nor U14850 (N_14850,N_14100,N_13875);
nor U14851 (N_14851,N_14075,N_14344);
nand U14852 (N_14852,N_14354,N_14112);
or U14853 (N_14853,N_14316,N_14134);
nand U14854 (N_14854,N_14214,N_13763);
or U14855 (N_14855,N_14169,N_13936);
xnor U14856 (N_14856,N_13851,N_14239);
nand U14857 (N_14857,N_14063,N_13956);
nor U14858 (N_14858,N_14113,N_14374);
nand U14859 (N_14859,N_13774,N_14280);
or U14860 (N_14860,N_14239,N_13799);
nor U14861 (N_14861,N_14090,N_14284);
and U14862 (N_14862,N_14143,N_14362);
or U14863 (N_14863,N_13799,N_14301);
or U14864 (N_14864,N_14313,N_14040);
or U14865 (N_14865,N_14015,N_14158);
and U14866 (N_14866,N_14184,N_13819);
nor U14867 (N_14867,N_14268,N_13984);
nor U14868 (N_14868,N_13752,N_13903);
and U14869 (N_14869,N_14167,N_14266);
nor U14870 (N_14870,N_14223,N_13957);
xnor U14871 (N_14871,N_13931,N_14029);
nand U14872 (N_14872,N_14283,N_13849);
and U14873 (N_14873,N_14073,N_14254);
or U14874 (N_14874,N_14198,N_13986);
and U14875 (N_14875,N_14244,N_13913);
nand U14876 (N_14876,N_14330,N_14015);
nand U14877 (N_14877,N_14013,N_14161);
or U14878 (N_14878,N_13888,N_13991);
nand U14879 (N_14879,N_14236,N_14266);
xor U14880 (N_14880,N_14285,N_14106);
nor U14881 (N_14881,N_13791,N_13912);
nand U14882 (N_14882,N_14250,N_14066);
xnor U14883 (N_14883,N_14310,N_13925);
nor U14884 (N_14884,N_14063,N_14057);
nor U14885 (N_14885,N_14257,N_14187);
nand U14886 (N_14886,N_14355,N_13869);
nor U14887 (N_14887,N_14113,N_14035);
nor U14888 (N_14888,N_13910,N_14124);
or U14889 (N_14889,N_14048,N_13812);
or U14890 (N_14890,N_13814,N_14194);
nand U14891 (N_14891,N_14205,N_14099);
nand U14892 (N_14892,N_14296,N_14244);
or U14893 (N_14893,N_14246,N_13795);
nor U14894 (N_14894,N_13888,N_14246);
nor U14895 (N_14895,N_14286,N_13782);
nand U14896 (N_14896,N_14176,N_13809);
nand U14897 (N_14897,N_13988,N_13970);
nor U14898 (N_14898,N_13840,N_13811);
nor U14899 (N_14899,N_13817,N_13931);
nor U14900 (N_14900,N_14103,N_13989);
xnor U14901 (N_14901,N_13837,N_14165);
and U14902 (N_14902,N_14287,N_13880);
and U14903 (N_14903,N_14369,N_13859);
and U14904 (N_14904,N_14374,N_14237);
and U14905 (N_14905,N_14293,N_13925);
or U14906 (N_14906,N_14252,N_13985);
nor U14907 (N_14907,N_13808,N_14290);
nand U14908 (N_14908,N_14212,N_13986);
or U14909 (N_14909,N_14318,N_13881);
xnor U14910 (N_14910,N_14282,N_13778);
or U14911 (N_14911,N_14340,N_13787);
or U14912 (N_14912,N_14014,N_13835);
nor U14913 (N_14913,N_14332,N_14079);
or U14914 (N_14914,N_13952,N_13813);
and U14915 (N_14915,N_13995,N_13782);
nor U14916 (N_14916,N_14165,N_14202);
or U14917 (N_14917,N_13996,N_13948);
and U14918 (N_14918,N_14056,N_14143);
nand U14919 (N_14919,N_14056,N_14359);
and U14920 (N_14920,N_14032,N_14201);
nor U14921 (N_14921,N_14272,N_14356);
nand U14922 (N_14922,N_14346,N_14203);
nand U14923 (N_14923,N_14355,N_13911);
nor U14924 (N_14924,N_14044,N_14237);
nand U14925 (N_14925,N_14246,N_13773);
xnor U14926 (N_14926,N_14100,N_14234);
nand U14927 (N_14927,N_14230,N_14365);
xor U14928 (N_14928,N_14181,N_14141);
or U14929 (N_14929,N_13898,N_14063);
and U14930 (N_14930,N_14029,N_14091);
nor U14931 (N_14931,N_14331,N_14340);
nor U14932 (N_14932,N_14004,N_14224);
nor U14933 (N_14933,N_13794,N_14014);
nor U14934 (N_14934,N_13951,N_14072);
xor U14935 (N_14935,N_14312,N_14077);
and U14936 (N_14936,N_14065,N_13902);
xor U14937 (N_14937,N_14209,N_14301);
nand U14938 (N_14938,N_14008,N_14203);
and U14939 (N_14939,N_14339,N_14105);
nand U14940 (N_14940,N_14113,N_14059);
nand U14941 (N_14941,N_14204,N_14360);
nor U14942 (N_14942,N_13967,N_14093);
nor U14943 (N_14943,N_14183,N_14107);
and U14944 (N_14944,N_14021,N_14046);
xnor U14945 (N_14945,N_14114,N_14044);
nand U14946 (N_14946,N_14237,N_14201);
nand U14947 (N_14947,N_14247,N_14017);
or U14948 (N_14948,N_13978,N_14288);
nand U14949 (N_14949,N_13933,N_14020);
or U14950 (N_14950,N_14070,N_14038);
and U14951 (N_14951,N_14363,N_14366);
or U14952 (N_14952,N_13834,N_13913);
nor U14953 (N_14953,N_14219,N_14322);
nand U14954 (N_14954,N_14284,N_13886);
nand U14955 (N_14955,N_14251,N_13866);
nor U14956 (N_14956,N_13800,N_14041);
and U14957 (N_14957,N_14233,N_14017);
xor U14958 (N_14958,N_14146,N_14168);
xnor U14959 (N_14959,N_13908,N_14257);
xor U14960 (N_14960,N_14014,N_14224);
xnor U14961 (N_14961,N_14209,N_14157);
or U14962 (N_14962,N_14295,N_13788);
nor U14963 (N_14963,N_14341,N_13889);
and U14964 (N_14964,N_13786,N_14214);
and U14965 (N_14965,N_14372,N_13970);
or U14966 (N_14966,N_14330,N_13892);
and U14967 (N_14967,N_13995,N_14300);
nor U14968 (N_14968,N_14276,N_13763);
or U14969 (N_14969,N_14222,N_13955);
xor U14970 (N_14970,N_13913,N_13837);
or U14971 (N_14971,N_14342,N_13923);
and U14972 (N_14972,N_14052,N_14058);
nor U14973 (N_14973,N_14015,N_14093);
or U14974 (N_14974,N_13997,N_13989);
nor U14975 (N_14975,N_13853,N_13904);
and U14976 (N_14976,N_14374,N_14116);
nor U14977 (N_14977,N_13961,N_14005);
nand U14978 (N_14978,N_13801,N_14347);
xor U14979 (N_14979,N_14115,N_13756);
or U14980 (N_14980,N_14243,N_14113);
and U14981 (N_14981,N_13794,N_13815);
and U14982 (N_14982,N_13770,N_14014);
xnor U14983 (N_14983,N_14213,N_14252);
xnor U14984 (N_14984,N_14079,N_13930);
nand U14985 (N_14985,N_14009,N_14253);
or U14986 (N_14986,N_13977,N_14109);
nand U14987 (N_14987,N_14074,N_13963);
xor U14988 (N_14988,N_14236,N_14212);
or U14989 (N_14989,N_14246,N_13979);
or U14990 (N_14990,N_14049,N_14175);
xnor U14991 (N_14991,N_13978,N_13966);
and U14992 (N_14992,N_13885,N_13771);
nor U14993 (N_14993,N_13866,N_14135);
or U14994 (N_14994,N_13794,N_14080);
xnor U14995 (N_14995,N_14241,N_14207);
nand U14996 (N_14996,N_13971,N_14011);
and U14997 (N_14997,N_14030,N_13978);
or U14998 (N_14998,N_14209,N_14159);
nor U14999 (N_14999,N_14308,N_14140);
and U15000 (N_15000,N_14844,N_14635);
nor U15001 (N_15001,N_14587,N_14814);
or U15002 (N_15002,N_14644,N_14861);
nor U15003 (N_15003,N_14738,N_14399);
nand U15004 (N_15004,N_14490,N_14522);
nand U15005 (N_15005,N_14904,N_14655);
nor U15006 (N_15006,N_14556,N_14726);
or U15007 (N_15007,N_14531,N_14873);
and U15008 (N_15008,N_14643,N_14764);
nor U15009 (N_15009,N_14530,N_14460);
or U15010 (N_15010,N_14827,N_14629);
and U15011 (N_15011,N_14456,N_14408);
or U15012 (N_15012,N_14618,N_14687);
nand U15013 (N_15013,N_14616,N_14778);
and U15014 (N_15014,N_14513,N_14736);
nand U15015 (N_15015,N_14458,N_14463);
nor U15016 (N_15016,N_14588,N_14877);
or U15017 (N_15017,N_14808,N_14582);
or U15018 (N_15018,N_14951,N_14999);
nor U15019 (N_15019,N_14989,N_14659);
or U15020 (N_15020,N_14622,N_14452);
nand U15021 (N_15021,N_14979,N_14426);
nand U15022 (N_15022,N_14545,N_14943);
xor U15023 (N_15023,N_14416,N_14699);
and U15024 (N_15024,N_14613,N_14594);
xor U15025 (N_15025,N_14538,N_14880);
or U15026 (N_15026,N_14684,N_14983);
nand U15027 (N_15027,N_14473,N_14624);
nor U15028 (N_15028,N_14892,N_14902);
nor U15029 (N_15029,N_14995,N_14383);
nand U15030 (N_15030,N_14905,N_14822);
nand U15031 (N_15031,N_14568,N_14579);
nor U15032 (N_15032,N_14879,N_14917);
nor U15033 (N_15033,N_14443,N_14719);
nand U15034 (N_15034,N_14851,N_14605);
nand U15035 (N_15035,N_14955,N_14679);
and U15036 (N_15036,N_14832,N_14535);
and U15037 (N_15037,N_14550,N_14639);
nand U15038 (N_15038,N_14547,N_14481);
nand U15039 (N_15039,N_14413,N_14649);
and U15040 (N_15040,N_14876,N_14920);
xor U15041 (N_15041,N_14772,N_14666);
or U15042 (N_15042,N_14509,N_14576);
or U15043 (N_15043,N_14821,N_14710);
nand U15044 (N_15044,N_14698,N_14669);
xor U15045 (N_15045,N_14985,N_14656);
and U15046 (N_15046,N_14966,N_14852);
or U15047 (N_15047,N_14391,N_14394);
nand U15048 (N_15048,N_14503,N_14665);
nand U15049 (N_15049,N_14575,N_14615);
nor U15050 (N_15050,N_14801,N_14878);
or U15051 (N_15051,N_14646,N_14753);
and U15052 (N_15052,N_14382,N_14725);
nor U15053 (N_15053,N_14381,N_14933);
and U15054 (N_15054,N_14889,N_14514);
or U15055 (N_15055,N_14454,N_14406);
nand U15056 (N_15056,N_14405,N_14584);
nand U15057 (N_15057,N_14922,N_14578);
or U15058 (N_15058,N_14745,N_14768);
nor U15059 (N_15059,N_14591,N_14968);
nand U15060 (N_15060,N_14941,N_14981);
nor U15061 (N_15061,N_14479,N_14818);
nand U15062 (N_15062,N_14694,N_14987);
nand U15063 (N_15063,N_14988,N_14478);
and U15064 (N_15064,N_14537,N_14396);
or U15065 (N_15065,N_14692,N_14900);
or U15066 (N_15066,N_14676,N_14414);
or U15067 (N_15067,N_14862,N_14846);
nor U15068 (N_15068,N_14491,N_14502);
or U15069 (N_15069,N_14740,N_14492);
nor U15070 (N_15070,N_14404,N_14543);
and U15071 (N_15071,N_14883,N_14901);
nor U15072 (N_15072,N_14984,N_14440);
xor U15073 (N_15073,N_14907,N_14602);
nand U15074 (N_15074,N_14668,N_14724);
or U15075 (N_15075,N_14886,N_14507);
or U15076 (N_15076,N_14449,N_14388);
nor U15077 (N_15077,N_14817,N_14779);
nor U15078 (N_15078,N_14563,N_14612);
nand U15079 (N_15079,N_14586,N_14841);
nor U15080 (N_15080,N_14558,N_14657);
nand U15081 (N_15081,N_14422,N_14908);
nor U15082 (N_15082,N_14662,N_14720);
nand U15083 (N_15083,N_14896,N_14378);
xnor U15084 (N_15084,N_14882,N_14885);
xor U15085 (N_15085,N_14804,N_14609);
nand U15086 (N_15086,N_14592,N_14658);
nand U15087 (N_15087,N_14627,N_14957);
nor U15088 (N_15088,N_14748,N_14648);
nor U15089 (N_15089,N_14527,N_14833);
xnor U15090 (N_15090,N_14867,N_14386);
nor U15091 (N_15091,N_14465,N_14916);
nand U15092 (N_15092,N_14810,N_14400);
and U15093 (N_15093,N_14675,N_14683);
or U15094 (N_15094,N_14718,N_14737);
or U15095 (N_15095,N_14500,N_14777);
and U15096 (N_15096,N_14897,N_14802);
nor U15097 (N_15097,N_14435,N_14497);
nand U15098 (N_15098,N_14775,N_14806);
nand U15099 (N_15099,N_14633,N_14891);
nor U15100 (N_15100,N_14993,N_14632);
nand U15101 (N_15101,N_14638,N_14825);
xnor U15102 (N_15102,N_14599,N_14474);
nor U15103 (N_15103,N_14570,N_14533);
or U15104 (N_15104,N_14704,N_14577);
nand U15105 (N_15105,N_14467,N_14919);
and U15106 (N_15106,N_14845,N_14762);
nand U15107 (N_15107,N_14721,N_14975);
xnor U15108 (N_15108,N_14485,N_14420);
and U15109 (N_15109,N_14767,N_14480);
xor U15110 (N_15110,N_14536,N_14826);
nor U15111 (N_15111,N_14785,N_14690);
nand U15112 (N_15112,N_14505,N_14793);
xor U15113 (N_15113,N_14604,N_14758);
xor U15114 (N_15114,N_14837,N_14540);
or U15115 (N_15115,N_14739,N_14411);
or U15116 (N_15116,N_14385,N_14702);
nor U15117 (N_15117,N_14663,N_14760);
nand U15118 (N_15118,N_14483,N_14800);
or U15119 (N_15119,N_14515,N_14723);
and U15120 (N_15120,N_14561,N_14432);
nor U15121 (N_15121,N_14567,N_14963);
nand U15122 (N_15122,N_14789,N_14766);
nor U15123 (N_15123,N_14645,N_14850);
nor U15124 (N_15124,N_14462,N_14595);
and U15125 (N_15125,N_14560,N_14512);
nor U15126 (N_15126,N_14392,N_14991);
or U15127 (N_15127,N_14598,N_14996);
or U15128 (N_15128,N_14534,N_14562);
nand U15129 (N_15129,N_14954,N_14744);
nand U15130 (N_15130,N_14998,N_14791);
and U15131 (N_15131,N_14436,N_14652);
and U15132 (N_15132,N_14823,N_14788);
and U15133 (N_15133,N_14375,N_14402);
nand U15134 (N_15134,N_14972,N_14664);
and U15135 (N_15135,N_14461,N_14630);
or U15136 (N_15136,N_14820,N_14994);
and U15137 (N_15137,N_14784,N_14417);
nand U15138 (N_15138,N_14847,N_14870);
nand U15139 (N_15139,N_14703,N_14783);
nor U15140 (N_15140,N_14819,N_14967);
nor U15141 (N_15141,N_14746,N_14978);
and U15142 (N_15142,N_14854,N_14924);
nand U15143 (N_15143,N_14839,N_14680);
nor U15144 (N_15144,N_14442,N_14596);
or U15145 (N_15145,N_14705,N_14672);
or U15146 (N_15146,N_14523,N_14494);
or U15147 (N_15147,N_14403,N_14696);
and U15148 (N_15148,N_14713,N_14600);
and U15149 (N_15149,N_14947,N_14830);
nor U15150 (N_15150,N_14464,N_14489);
and U15151 (N_15151,N_14795,N_14756);
and U15152 (N_15152,N_14812,N_14541);
nand U15153 (N_15153,N_14376,N_14487);
or U15154 (N_15154,N_14660,N_14903);
nand U15155 (N_15155,N_14637,N_14899);
nor U15156 (N_15156,N_14939,N_14603);
nand U15157 (N_15157,N_14695,N_14455);
and U15158 (N_15158,N_14722,N_14921);
nor U15159 (N_15159,N_14667,N_14387);
or U15160 (N_15160,N_14453,N_14792);
nand U15161 (N_15161,N_14790,N_14750);
or U15162 (N_15162,N_14593,N_14379);
or U15163 (N_15163,N_14625,N_14734);
or U15164 (N_15164,N_14755,N_14499);
nand U15165 (N_15165,N_14843,N_14834);
and U15166 (N_15166,N_14524,N_14642);
nor U15167 (N_15167,N_14516,N_14752);
and U15168 (N_15168,N_14958,N_14913);
nor U15169 (N_15169,N_14647,N_14773);
nand U15170 (N_15170,N_14759,N_14496);
or U15171 (N_15171,N_14807,N_14931);
and U15172 (N_15172,N_14433,N_14945);
or U15173 (N_15173,N_14621,N_14786);
or U15174 (N_15174,N_14743,N_14971);
nand U15175 (N_15175,N_14796,N_14770);
nand U15176 (N_15176,N_14636,N_14677);
nor U15177 (N_15177,N_14398,N_14787);
and U15178 (N_15178,N_14735,N_14765);
nor U15179 (N_15179,N_14559,N_14393);
nand U15180 (N_15180,N_14691,N_14554);
nand U15181 (N_15181,N_14869,N_14508);
nand U15182 (N_15182,N_14553,N_14868);
nor U15183 (N_15183,N_14428,N_14693);
nor U15184 (N_15184,N_14937,N_14729);
nor U15185 (N_15185,N_14776,N_14551);
nand U15186 (N_15186,N_14678,N_14395);
or U15187 (N_15187,N_14557,N_14674);
xnor U15188 (N_15188,N_14970,N_14888);
and U15189 (N_15189,N_14701,N_14544);
and U15190 (N_15190,N_14439,N_14976);
nor U15191 (N_15191,N_14871,N_14620);
or U15192 (N_15192,N_14751,N_14427);
and U15193 (N_15193,N_14451,N_14938);
or U15194 (N_15194,N_14617,N_14472);
and U15195 (N_15195,N_14589,N_14708);
and U15196 (N_15196,N_14741,N_14434);
or U15197 (N_15197,N_14798,N_14520);
nor U15198 (N_15198,N_14488,N_14377);
or U15199 (N_15199,N_14401,N_14504);
or U15200 (N_15200,N_14840,N_14641);
nand U15201 (N_15201,N_14730,N_14842);
nand U15202 (N_15202,N_14688,N_14856);
nor U15203 (N_15203,N_14528,N_14510);
xnor U15204 (N_15204,N_14815,N_14619);
and U15205 (N_15205,N_14486,N_14857);
nand U15206 (N_15206,N_14910,N_14511);
and U15207 (N_15207,N_14742,N_14495);
nand U15208 (N_15208,N_14813,N_14781);
xor U15209 (N_15209,N_14441,N_14893);
or U15210 (N_15210,N_14731,N_14585);
xnor U15211 (N_15211,N_14969,N_14623);
nor U15212 (N_15212,N_14757,N_14608);
and U15213 (N_15213,N_14997,N_14733);
and U15214 (N_15214,N_14960,N_14912);
nand U15215 (N_15215,N_14949,N_14709);
nand U15216 (N_15216,N_14761,N_14574);
nand U15217 (N_15217,N_14858,N_14525);
nand U15218 (N_15218,N_14606,N_14909);
nor U15219 (N_15219,N_14824,N_14895);
and U15220 (N_15220,N_14874,N_14727);
nand U15221 (N_15221,N_14884,N_14390);
xor U15222 (N_15222,N_14389,N_14468);
and U15223 (N_15223,N_14835,N_14681);
or U15224 (N_15224,N_14477,N_14650);
nor U15225 (N_15225,N_14447,N_14894);
nor U15226 (N_15226,N_14601,N_14711);
nand U15227 (N_15227,N_14935,N_14973);
and U15228 (N_15228,N_14457,N_14532);
nand U15229 (N_15229,N_14397,N_14546);
nor U15230 (N_15230,N_14934,N_14864);
and U15231 (N_15231,N_14446,N_14927);
or U15232 (N_15232,N_14566,N_14419);
xor U15233 (N_15233,N_14425,N_14469);
nand U15234 (N_15234,N_14542,N_14805);
nand U15235 (N_15235,N_14626,N_14831);
xor U15236 (N_15236,N_14671,N_14860);
or U15237 (N_15237,N_14670,N_14572);
xnor U15238 (N_15238,N_14610,N_14521);
nor U15239 (N_15239,N_14848,N_14717);
or U15240 (N_15240,N_14849,N_14926);
or U15241 (N_15241,N_14942,N_14407);
and U15242 (N_15242,N_14986,N_14549);
or U15243 (N_15243,N_14580,N_14747);
or U15244 (N_15244,N_14929,N_14948);
xnor U15245 (N_15245,N_14707,N_14881);
nor U15246 (N_15246,N_14529,N_14686);
nor U15247 (N_15247,N_14809,N_14782);
xor U15248 (N_15248,N_14590,N_14838);
nand U15249 (N_15249,N_14769,N_14863);
nor U15250 (N_15250,N_14424,N_14431);
or U15251 (N_15251,N_14906,N_14493);
nand U15252 (N_15252,N_14429,N_14853);
or U15253 (N_15253,N_14715,N_14459);
nor U15254 (N_15254,N_14614,N_14423);
nor U15255 (N_15255,N_14548,N_14816);
or U15256 (N_15256,N_14977,N_14475);
nor U15257 (N_15257,N_14539,N_14571);
or U15258 (N_15258,N_14962,N_14859);
nor U15259 (N_15259,N_14654,N_14990);
or U15260 (N_15260,N_14811,N_14866);
or U15261 (N_15261,N_14506,N_14923);
or U15262 (N_15262,N_14925,N_14682);
or U15263 (N_15263,N_14438,N_14961);
nor U15264 (N_15264,N_14898,N_14697);
nor U15265 (N_15265,N_14430,N_14384);
nand U15266 (N_15266,N_14890,N_14872);
and U15267 (N_15267,N_14875,N_14466);
nor U15268 (N_15268,N_14953,N_14661);
or U15269 (N_15269,N_14940,N_14640);
nor U15270 (N_15270,N_14569,N_14484);
and U15271 (N_15271,N_14911,N_14936);
nand U15272 (N_15272,N_14771,N_14445);
or U15273 (N_15273,N_14628,N_14980);
xor U15274 (N_15274,N_14749,N_14418);
xor U15275 (N_15275,N_14476,N_14611);
or U15276 (N_15276,N_14415,N_14930);
or U15277 (N_15277,N_14555,N_14448);
nand U15278 (N_15278,N_14865,N_14573);
or U15279 (N_15279,N_14410,N_14797);
nand U15280 (N_15280,N_14828,N_14728);
and U15281 (N_15281,N_14928,N_14689);
nand U15282 (N_15282,N_14498,N_14565);
nor U15283 (N_15283,N_14409,N_14780);
nand U15284 (N_15284,N_14803,N_14918);
and U15285 (N_15285,N_14774,N_14982);
and U15286 (N_15286,N_14915,N_14564);
or U15287 (N_15287,N_14673,N_14716);
and U15288 (N_15288,N_14794,N_14685);
and U15289 (N_15289,N_14517,N_14950);
nand U15290 (N_15290,N_14829,N_14754);
and U15291 (N_15291,N_14471,N_14700);
and U15292 (N_15292,N_14714,N_14946);
and U15293 (N_15293,N_14552,N_14763);
nand U15294 (N_15294,N_14583,N_14952);
nor U15295 (N_15295,N_14712,N_14482);
or U15296 (N_15296,N_14470,N_14932);
nand U15297 (N_15297,N_14799,N_14887);
nor U15298 (N_15298,N_14956,N_14597);
and U15299 (N_15299,N_14581,N_14450);
and U15300 (N_15300,N_14634,N_14974);
and U15301 (N_15301,N_14412,N_14519);
and U15302 (N_15302,N_14444,N_14965);
nor U15303 (N_15303,N_14421,N_14653);
nand U15304 (N_15304,N_14501,N_14992);
or U15305 (N_15305,N_14964,N_14959);
or U15306 (N_15306,N_14526,N_14944);
and U15307 (N_15307,N_14631,N_14706);
or U15308 (N_15308,N_14732,N_14437);
and U15309 (N_15309,N_14380,N_14651);
nand U15310 (N_15310,N_14607,N_14914);
xnor U15311 (N_15311,N_14518,N_14836);
nand U15312 (N_15312,N_14855,N_14410);
xnor U15313 (N_15313,N_14612,N_14447);
nand U15314 (N_15314,N_14743,N_14938);
xor U15315 (N_15315,N_14862,N_14602);
xor U15316 (N_15316,N_14441,N_14382);
xnor U15317 (N_15317,N_14773,N_14700);
nor U15318 (N_15318,N_14538,N_14521);
and U15319 (N_15319,N_14891,N_14814);
and U15320 (N_15320,N_14453,N_14491);
nand U15321 (N_15321,N_14756,N_14995);
and U15322 (N_15322,N_14813,N_14403);
xnor U15323 (N_15323,N_14375,N_14494);
or U15324 (N_15324,N_14536,N_14890);
nor U15325 (N_15325,N_14919,N_14676);
or U15326 (N_15326,N_14838,N_14552);
nor U15327 (N_15327,N_14688,N_14583);
nand U15328 (N_15328,N_14809,N_14670);
nor U15329 (N_15329,N_14769,N_14966);
and U15330 (N_15330,N_14382,N_14761);
and U15331 (N_15331,N_14683,N_14858);
nor U15332 (N_15332,N_14589,N_14878);
or U15333 (N_15333,N_14722,N_14541);
nor U15334 (N_15334,N_14405,N_14675);
nor U15335 (N_15335,N_14695,N_14991);
nor U15336 (N_15336,N_14970,N_14847);
and U15337 (N_15337,N_14605,N_14619);
nor U15338 (N_15338,N_14733,N_14730);
and U15339 (N_15339,N_14583,N_14714);
and U15340 (N_15340,N_14632,N_14574);
or U15341 (N_15341,N_14655,N_14566);
nand U15342 (N_15342,N_14448,N_14777);
nand U15343 (N_15343,N_14417,N_14925);
nor U15344 (N_15344,N_14571,N_14495);
nor U15345 (N_15345,N_14422,N_14981);
nor U15346 (N_15346,N_14906,N_14546);
nand U15347 (N_15347,N_14922,N_14387);
xnor U15348 (N_15348,N_14579,N_14585);
nand U15349 (N_15349,N_14378,N_14905);
and U15350 (N_15350,N_14999,N_14845);
or U15351 (N_15351,N_14709,N_14676);
and U15352 (N_15352,N_14612,N_14533);
and U15353 (N_15353,N_14701,N_14945);
nand U15354 (N_15354,N_14847,N_14594);
nor U15355 (N_15355,N_14719,N_14668);
nor U15356 (N_15356,N_14660,N_14515);
or U15357 (N_15357,N_14993,N_14919);
nand U15358 (N_15358,N_14709,N_14712);
nand U15359 (N_15359,N_14745,N_14639);
and U15360 (N_15360,N_14672,N_14478);
nand U15361 (N_15361,N_14479,N_14395);
nor U15362 (N_15362,N_14673,N_14672);
xor U15363 (N_15363,N_14829,N_14669);
nor U15364 (N_15364,N_14620,N_14847);
and U15365 (N_15365,N_14789,N_14908);
nand U15366 (N_15366,N_14438,N_14386);
and U15367 (N_15367,N_14994,N_14826);
nor U15368 (N_15368,N_14755,N_14715);
and U15369 (N_15369,N_14647,N_14991);
nor U15370 (N_15370,N_14975,N_14932);
xnor U15371 (N_15371,N_14776,N_14377);
and U15372 (N_15372,N_14492,N_14504);
and U15373 (N_15373,N_14464,N_14928);
or U15374 (N_15374,N_14750,N_14448);
xor U15375 (N_15375,N_14521,N_14632);
or U15376 (N_15376,N_14470,N_14456);
or U15377 (N_15377,N_14408,N_14423);
nor U15378 (N_15378,N_14731,N_14557);
nor U15379 (N_15379,N_14625,N_14708);
or U15380 (N_15380,N_14669,N_14725);
or U15381 (N_15381,N_14405,N_14610);
and U15382 (N_15382,N_14744,N_14487);
and U15383 (N_15383,N_14701,N_14663);
and U15384 (N_15384,N_14706,N_14932);
and U15385 (N_15385,N_14950,N_14828);
nor U15386 (N_15386,N_14702,N_14953);
nor U15387 (N_15387,N_14690,N_14943);
nand U15388 (N_15388,N_14881,N_14816);
nor U15389 (N_15389,N_14719,N_14616);
nor U15390 (N_15390,N_14821,N_14965);
nor U15391 (N_15391,N_14904,N_14638);
nor U15392 (N_15392,N_14723,N_14629);
nand U15393 (N_15393,N_14809,N_14496);
nor U15394 (N_15394,N_14586,N_14874);
nor U15395 (N_15395,N_14530,N_14727);
nor U15396 (N_15396,N_14744,N_14914);
and U15397 (N_15397,N_14844,N_14670);
or U15398 (N_15398,N_14435,N_14773);
or U15399 (N_15399,N_14820,N_14763);
and U15400 (N_15400,N_14554,N_14457);
or U15401 (N_15401,N_14959,N_14766);
nor U15402 (N_15402,N_14393,N_14795);
xor U15403 (N_15403,N_14989,N_14572);
or U15404 (N_15404,N_14655,N_14636);
and U15405 (N_15405,N_14516,N_14910);
and U15406 (N_15406,N_14412,N_14876);
or U15407 (N_15407,N_14637,N_14701);
nor U15408 (N_15408,N_14418,N_14530);
xnor U15409 (N_15409,N_14988,N_14812);
nand U15410 (N_15410,N_14624,N_14450);
and U15411 (N_15411,N_14979,N_14983);
or U15412 (N_15412,N_14696,N_14830);
or U15413 (N_15413,N_14927,N_14934);
or U15414 (N_15414,N_14699,N_14410);
nor U15415 (N_15415,N_14839,N_14901);
nand U15416 (N_15416,N_14977,N_14384);
xor U15417 (N_15417,N_14416,N_14527);
nor U15418 (N_15418,N_14694,N_14631);
and U15419 (N_15419,N_14768,N_14790);
xnor U15420 (N_15420,N_14666,N_14574);
and U15421 (N_15421,N_14440,N_14894);
nand U15422 (N_15422,N_14733,N_14605);
or U15423 (N_15423,N_14909,N_14458);
nand U15424 (N_15424,N_14993,N_14795);
and U15425 (N_15425,N_14715,N_14593);
and U15426 (N_15426,N_14494,N_14475);
or U15427 (N_15427,N_14634,N_14598);
nor U15428 (N_15428,N_14428,N_14612);
nor U15429 (N_15429,N_14968,N_14747);
or U15430 (N_15430,N_14945,N_14942);
xnor U15431 (N_15431,N_14982,N_14412);
and U15432 (N_15432,N_14440,N_14854);
and U15433 (N_15433,N_14877,N_14443);
and U15434 (N_15434,N_14631,N_14626);
nand U15435 (N_15435,N_14733,N_14575);
or U15436 (N_15436,N_14727,N_14416);
or U15437 (N_15437,N_14679,N_14419);
or U15438 (N_15438,N_14531,N_14397);
xor U15439 (N_15439,N_14479,N_14909);
or U15440 (N_15440,N_14872,N_14396);
or U15441 (N_15441,N_14661,N_14671);
nand U15442 (N_15442,N_14976,N_14484);
and U15443 (N_15443,N_14412,N_14520);
or U15444 (N_15444,N_14899,N_14420);
or U15445 (N_15445,N_14500,N_14650);
nor U15446 (N_15446,N_14725,N_14638);
nor U15447 (N_15447,N_14422,N_14603);
nor U15448 (N_15448,N_14610,N_14917);
and U15449 (N_15449,N_14818,N_14393);
nor U15450 (N_15450,N_14816,N_14474);
xnor U15451 (N_15451,N_14490,N_14842);
and U15452 (N_15452,N_14549,N_14820);
nand U15453 (N_15453,N_14605,N_14436);
nor U15454 (N_15454,N_14764,N_14625);
and U15455 (N_15455,N_14862,N_14482);
nand U15456 (N_15456,N_14659,N_14618);
or U15457 (N_15457,N_14496,N_14487);
xor U15458 (N_15458,N_14562,N_14620);
or U15459 (N_15459,N_14493,N_14605);
or U15460 (N_15460,N_14911,N_14978);
or U15461 (N_15461,N_14531,N_14400);
nor U15462 (N_15462,N_14618,N_14600);
nand U15463 (N_15463,N_14638,N_14780);
or U15464 (N_15464,N_14641,N_14681);
and U15465 (N_15465,N_14759,N_14890);
or U15466 (N_15466,N_14963,N_14786);
nor U15467 (N_15467,N_14760,N_14457);
or U15468 (N_15468,N_14469,N_14662);
nor U15469 (N_15469,N_14655,N_14494);
nand U15470 (N_15470,N_14413,N_14805);
or U15471 (N_15471,N_14984,N_14873);
nand U15472 (N_15472,N_14677,N_14475);
nor U15473 (N_15473,N_14746,N_14975);
or U15474 (N_15474,N_14587,N_14482);
and U15475 (N_15475,N_14704,N_14946);
and U15476 (N_15476,N_14428,N_14511);
or U15477 (N_15477,N_14412,N_14561);
nor U15478 (N_15478,N_14442,N_14478);
xor U15479 (N_15479,N_14802,N_14764);
and U15480 (N_15480,N_14770,N_14443);
xor U15481 (N_15481,N_14874,N_14686);
and U15482 (N_15482,N_14967,N_14436);
xnor U15483 (N_15483,N_14867,N_14483);
nand U15484 (N_15484,N_14461,N_14468);
nand U15485 (N_15485,N_14403,N_14760);
nand U15486 (N_15486,N_14673,N_14933);
or U15487 (N_15487,N_14753,N_14744);
nand U15488 (N_15488,N_14939,N_14734);
and U15489 (N_15489,N_14471,N_14568);
nand U15490 (N_15490,N_14843,N_14572);
nor U15491 (N_15491,N_14569,N_14423);
nand U15492 (N_15492,N_14807,N_14830);
nand U15493 (N_15493,N_14636,N_14483);
nand U15494 (N_15494,N_14584,N_14720);
and U15495 (N_15495,N_14441,N_14865);
and U15496 (N_15496,N_14888,N_14618);
nand U15497 (N_15497,N_14905,N_14681);
nor U15498 (N_15498,N_14520,N_14511);
or U15499 (N_15499,N_14822,N_14951);
nand U15500 (N_15500,N_14509,N_14958);
nor U15501 (N_15501,N_14598,N_14496);
nand U15502 (N_15502,N_14607,N_14875);
xor U15503 (N_15503,N_14684,N_14652);
or U15504 (N_15504,N_14512,N_14410);
nand U15505 (N_15505,N_14444,N_14566);
and U15506 (N_15506,N_14649,N_14552);
nor U15507 (N_15507,N_14568,N_14401);
nand U15508 (N_15508,N_14743,N_14752);
xor U15509 (N_15509,N_14779,N_14746);
and U15510 (N_15510,N_14674,N_14631);
and U15511 (N_15511,N_14495,N_14398);
nor U15512 (N_15512,N_14606,N_14693);
nor U15513 (N_15513,N_14385,N_14688);
nand U15514 (N_15514,N_14458,N_14791);
nand U15515 (N_15515,N_14726,N_14937);
nand U15516 (N_15516,N_14690,N_14691);
and U15517 (N_15517,N_14476,N_14804);
and U15518 (N_15518,N_14752,N_14674);
and U15519 (N_15519,N_14414,N_14794);
and U15520 (N_15520,N_14463,N_14476);
nand U15521 (N_15521,N_14543,N_14546);
or U15522 (N_15522,N_14579,N_14644);
nand U15523 (N_15523,N_14705,N_14484);
or U15524 (N_15524,N_14563,N_14694);
and U15525 (N_15525,N_14646,N_14494);
nand U15526 (N_15526,N_14761,N_14434);
nand U15527 (N_15527,N_14565,N_14603);
nor U15528 (N_15528,N_14900,N_14410);
and U15529 (N_15529,N_14795,N_14846);
nand U15530 (N_15530,N_14422,N_14518);
or U15531 (N_15531,N_14949,N_14692);
nand U15532 (N_15532,N_14830,N_14825);
nand U15533 (N_15533,N_14575,N_14839);
or U15534 (N_15534,N_14941,N_14949);
nor U15535 (N_15535,N_14443,N_14908);
xor U15536 (N_15536,N_14740,N_14624);
or U15537 (N_15537,N_14690,N_14642);
nand U15538 (N_15538,N_14936,N_14653);
or U15539 (N_15539,N_14789,N_14971);
or U15540 (N_15540,N_14778,N_14595);
and U15541 (N_15541,N_14656,N_14733);
nor U15542 (N_15542,N_14809,N_14428);
nand U15543 (N_15543,N_14510,N_14752);
nor U15544 (N_15544,N_14465,N_14862);
nand U15545 (N_15545,N_14589,N_14502);
and U15546 (N_15546,N_14513,N_14844);
nor U15547 (N_15547,N_14606,N_14950);
nand U15548 (N_15548,N_14820,N_14928);
or U15549 (N_15549,N_14885,N_14918);
xnor U15550 (N_15550,N_14482,N_14458);
and U15551 (N_15551,N_14567,N_14558);
and U15552 (N_15552,N_14380,N_14435);
and U15553 (N_15553,N_14650,N_14475);
nand U15554 (N_15554,N_14559,N_14610);
nor U15555 (N_15555,N_14512,N_14799);
nor U15556 (N_15556,N_14939,N_14893);
or U15557 (N_15557,N_14461,N_14746);
and U15558 (N_15558,N_14950,N_14667);
nor U15559 (N_15559,N_14648,N_14965);
or U15560 (N_15560,N_14966,N_14725);
nand U15561 (N_15561,N_14821,N_14439);
nand U15562 (N_15562,N_14673,N_14948);
nor U15563 (N_15563,N_14663,N_14941);
and U15564 (N_15564,N_14494,N_14927);
and U15565 (N_15565,N_14587,N_14604);
and U15566 (N_15566,N_14603,N_14636);
nand U15567 (N_15567,N_14824,N_14777);
nand U15568 (N_15568,N_14883,N_14762);
nand U15569 (N_15569,N_14815,N_14840);
nor U15570 (N_15570,N_14413,N_14916);
nor U15571 (N_15571,N_14836,N_14386);
and U15572 (N_15572,N_14891,N_14771);
or U15573 (N_15573,N_14651,N_14667);
nor U15574 (N_15574,N_14995,N_14867);
nor U15575 (N_15575,N_14752,N_14976);
and U15576 (N_15576,N_14939,N_14834);
nor U15577 (N_15577,N_14838,N_14487);
or U15578 (N_15578,N_14428,N_14851);
nor U15579 (N_15579,N_14934,N_14923);
or U15580 (N_15580,N_14509,N_14794);
nor U15581 (N_15581,N_14526,N_14841);
and U15582 (N_15582,N_14676,N_14640);
or U15583 (N_15583,N_14442,N_14522);
nor U15584 (N_15584,N_14892,N_14395);
or U15585 (N_15585,N_14402,N_14764);
xor U15586 (N_15586,N_14543,N_14902);
nand U15587 (N_15587,N_14658,N_14561);
nand U15588 (N_15588,N_14501,N_14639);
and U15589 (N_15589,N_14906,N_14603);
nor U15590 (N_15590,N_14608,N_14614);
and U15591 (N_15591,N_14489,N_14432);
nand U15592 (N_15592,N_14990,N_14564);
or U15593 (N_15593,N_14960,N_14796);
or U15594 (N_15594,N_14839,N_14395);
and U15595 (N_15595,N_14881,N_14413);
nand U15596 (N_15596,N_14704,N_14967);
nand U15597 (N_15597,N_14642,N_14503);
xor U15598 (N_15598,N_14415,N_14946);
nand U15599 (N_15599,N_14987,N_14421);
and U15600 (N_15600,N_14825,N_14916);
nor U15601 (N_15601,N_14600,N_14570);
nor U15602 (N_15602,N_14942,N_14685);
xnor U15603 (N_15603,N_14421,N_14743);
xnor U15604 (N_15604,N_14714,N_14866);
xnor U15605 (N_15605,N_14778,N_14605);
nor U15606 (N_15606,N_14641,N_14759);
or U15607 (N_15607,N_14497,N_14628);
xnor U15608 (N_15608,N_14684,N_14728);
nor U15609 (N_15609,N_14654,N_14389);
and U15610 (N_15610,N_14803,N_14890);
and U15611 (N_15611,N_14612,N_14569);
nand U15612 (N_15612,N_14841,N_14378);
nor U15613 (N_15613,N_14925,N_14663);
or U15614 (N_15614,N_14981,N_14785);
or U15615 (N_15615,N_14809,N_14446);
and U15616 (N_15616,N_14531,N_14643);
nand U15617 (N_15617,N_14819,N_14914);
xor U15618 (N_15618,N_14450,N_14616);
and U15619 (N_15619,N_14826,N_14631);
nand U15620 (N_15620,N_14711,N_14389);
nor U15621 (N_15621,N_14420,N_14907);
xnor U15622 (N_15622,N_14785,N_14587);
nor U15623 (N_15623,N_14697,N_14986);
xor U15624 (N_15624,N_14527,N_14737);
and U15625 (N_15625,N_15438,N_15383);
or U15626 (N_15626,N_15172,N_15111);
nor U15627 (N_15627,N_15454,N_15305);
nand U15628 (N_15628,N_15162,N_15423);
nand U15629 (N_15629,N_15098,N_15518);
nor U15630 (N_15630,N_15060,N_15363);
and U15631 (N_15631,N_15067,N_15319);
or U15632 (N_15632,N_15266,N_15011);
or U15633 (N_15633,N_15347,N_15083);
nand U15634 (N_15634,N_15493,N_15047);
nor U15635 (N_15635,N_15291,N_15257);
and U15636 (N_15636,N_15290,N_15317);
and U15637 (N_15637,N_15124,N_15270);
xor U15638 (N_15638,N_15443,N_15262);
and U15639 (N_15639,N_15497,N_15404);
nor U15640 (N_15640,N_15128,N_15148);
nand U15641 (N_15641,N_15224,N_15177);
nor U15642 (N_15642,N_15178,N_15594);
nand U15643 (N_15643,N_15514,N_15409);
or U15644 (N_15644,N_15254,N_15462);
and U15645 (N_15645,N_15055,N_15314);
nand U15646 (N_15646,N_15492,N_15231);
or U15647 (N_15647,N_15465,N_15010);
and U15648 (N_15648,N_15031,N_15420);
or U15649 (N_15649,N_15209,N_15250);
or U15650 (N_15650,N_15119,N_15338);
and U15651 (N_15651,N_15592,N_15308);
nor U15652 (N_15652,N_15132,N_15088);
or U15653 (N_15653,N_15028,N_15073);
xnor U15654 (N_15654,N_15244,N_15623);
or U15655 (N_15655,N_15237,N_15134);
and U15656 (N_15656,N_15442,N_15439);
nor U15657 (N_15657,N_15387,N_15612);
or U15658 (N_15658,N_15546,N_15100);
and U15659 (N_15659,N_15530,N_15551);
xnor U15660 (N_15660,N_15488,N_15105);
or U15661 (N_15661,N_15273,N_15045);
nor U15662 (N_15662,N_15416,N_15240);
nand U15663 (N_15663,N_15371,N_15152);
nor U15664 (N_15664,N_15298,N_15188);
xor U15665 (N_15665,N_15142,N_15212);
xor U15666 (N_15666,N_15446,N_15115);
or U15667 (N_15667,N_15059,N_15522);
and U15668 (N_15668,N_15200,N_15141);
nor U15669 (N_15669,N_15515,N_15012);
nand U15670 (N_15670,N_15025,N_15198);
and U15671 (N_15671,N_15410,N_15516);
nand U15672 (N_15672,N_15620,N_15364);
nor U15673 (N_15673,N_15099,N_15334);
and U15674 (N_15674,N_15597,N_15390);
and U15675 (N_15675,N_15370,N_15455);
and U15676 (N_15676,N_15258,N_15274);
or U15677 (N_15677,N_15158,N_15386);
or U15678 (N_15678,N_15357,N_15474);
or U15679 (N_15679,N_15304,N_15121);
nand U15680 (N_15680,N_15016,N_15260);
nor U15681 (N_15681,N_15211,N_15373);
nor U15682 (N_15682,N_15384,N_15160);
nor U15683 (N_15683,N_15603,N_15261);
nand U15684 (N_15684,N_15513,N_15070);
nand U15685 (N_15685,N_15379,N_15502);
and U15686 (N_15686,N_15399,N_15206);
or U15687 (N_15687,N_15496,N_15295);
nand U15688 (N_15688,N_15131,N_15065);
and U15689 (N_15689,N_15227,N_15569);
or U15690 (N_15690,N_15368,N_15577);
or U15691 (N_15691,N_15269,N_15267);
and U15692 (N_15692,N_15264,N_15579);
xor U15693 (N_15693,N_15071,N_15208);
or U15694 (N_15694,N_15351,N_15453);
and U15695 (N_15695,N_15552,N_15478);
nand U15696 (N_15696,N_15043,N_15299);
and U15697 (N_15697,N_15604,N_15582);
or U15698 (N_15698,N_15234,N_15150);
xnor U15699 (N_15699,N_15221,N_15553);
and U15700 (N_15700,N_15035,N_15157);
and U15701 (N_15701,N_15598,N_15210);
nand U15702 (N_15702,N_15600,N_15168);
nand U15703 (N_15703,N_15560,N_15102);
xnor U15704 (N_15704,N_15116,N_15170);
and U15705 (N_15705,N_15617,N_15312);
nand U15706 (N_15706,N_15459,N_15380);
nor U15707 (N_15707,N_15547,N_15203);
nor U15708 (N_15708,N_15507,N_15500);
nand U15709 (N_15709,N_15356,N_15108);
xnor U15710 (N_15710,N_15041,N_15126);
xnor U15711 (N_15711,N_15343,N_15434);
xnor U15712 (N_15712,N_15220,N_15335);
or U15713 (N_15713,N_15532,N_15483);
and U15714 (N_15714,N_15614,N_15535);
or U15715 (N_15715,N_15315,N_15584);
nand U15716 (N_15716,N_15398,N_15097);
xor U15717 (N_15717,N_15214,N_15018);
xnor U15718 (N_15718,N_15329,N_15447);
or U15719 (N_15719,N_15174,N_15293);
nor U15720 (N_15720,N_15036,N_15498);
nor U15721 (N_15721,N_15359,N_15136);
nand U15722 (N_15722,N_15327,N_15183);
nor U15723 (N_15723,N_15272,N_15505);
nand U15724 (N_15724,N_15280,N_15068);
nor U15725 (N_15725,N_15281,N_15382);
xnor U15726 (N_15726,N_15138,N_15189);
xor U15727 (N_15727,N_15355,N_15217);
and U15728 (N_15728,N_15029,N_15089);
nor U15729 (N_15729,N_15246,N_15524);
nand U15730 (N_15730,N_15169,N_15512);
nand U15731 (N_15731,N_15292,N_15086);
nand U15732 (N_15732,N_15540,N_15021);
nand U15733 (N_15733,N_15185,N_15079);
nor U15734 (N_15734,N_15143,N_15531);
and U15735 (N_15735,N_15557,N_15448);
and U15736 (N_15736,N_15618,N_15032);
and U15737 (N_15737,N_15601,N_15320);
and U15738 (N_15738,N_15048,N_15468);
and U15739 (N_15739,N_15288,N_15568);
nand U15740 (N_15740,N_15107,N_15092);
nand U15741 (N_15741,N_15578,N_15187);
or U15742 (N_15742,N_15415,N_15595);
nor U15743 (N_15743,N_15616,N_15133);
and U15744 (N_15744,N_15477,N_15606);
and U15745 (N_15745,N_15407,N_15590);
nand U15746 (N_15746,N_15374,N_15112);
nor U15747 (N_15747,N_15457,N_15147);
xor U15748 (N_15748,N_15511,N_15326);
xnor U15749 (N_15749,N_15276,N_15622);
nand U15750 (N_15750,N_15182,N_15085);
or U15751 (N_15751,N_15378,N_15309);
and U15752 (N_15752,N_15425,N_15440);
nor U15753 (N_15753,N_15419,N_15243);
nor U15754 (N_15754,N_15332,N_15122);
nor U15755 (N_15755,N_15003,N_15389);
nor U15756 (N_15756,N_15545,N_15275);
nor U15757 (N_15757,N_15471,N_15554);
nand U15758 (N_15758,N_15323,N_15619);
or U15759 (N_15759,N_15395,N_15000);
nand U15760 (N_15760,N_15192,N_15228);
and U15761 (N_15761,N_15113,N_15479);
and U15762 (N_15762,N_15422,N_15023);
and U15763 (N_15763,N_15521,N_15322);
and U15764 (N_15764,N_15367,N_15296);
nor U15765 (N_15765,N_15608,N_15585);
nand U15766 (N_15766,N_15570,N_15181);
and U15767 (N_15767,N_15544,N_15624);
and U15768 (N_15768,N_15044,N_15485);
and U15769 (N_15769,N_15056,N_15583);
or U15770 (N_15770,N_15233,N_15615);
and U15771 (N_15771,N_15534,N_15104);
or U15772 (N_15772,N_15571,N_15196);
nor U15773 (N_15773,N_15341,N_15194);
or U15774 (N_15774,N_15596,N_15084);
or U15775 (N_15775,N_15171,N_15490);
nor U15776 (N_15776,N_15241,N_15561);
or U15777 (N_15777,N_15421,N_15451);
nor U15778 (N_15778,N_15253,N_15247);
xor U15779 (N_15779,N_15350,N_15205);
nor U15780 (N_15780,N_15572,N_15392);
xnor U15781 (N_15781,N_15548,N_15473);
and U15782 (N_15782,N_15489,N_15316);
nand U15783 (N_15783,N_15197,N_15175);
and U15784 (N_15784,N_15081,N_15051);
and U15785 (N_15785,N_15216,N_15057);
and U15786 (N_15786,N_15366,N_15005);
nor U15787 (N_15787,N_15445,N_15580);
and U15788 (N_15788,N_15400,N_15263);
nor U15789 (N_15789,N_15574,N_15426);
nor U15790 (N_15790,N_15340,N_15542);
and U15791 (N_15791,N_15388,N_15218);
nand U15792 (N_15792,N_15159,N_15487);
nand U15793 (N_15793,N_15501,N_15480);
and U15794 (N_15794,N_15195,N_15215);
xnor U15795 (N_15795,N_15167,N_15476);
nand U15796 (N_15796,N_15467,N_15180);
or U15797 (N_15797,N_15325,N_15082);
nor U15798 (N_15798,N_15565,N_15433);
xnor U15799 (N_15799,N_15144,N_15255);
nor U15800 (N_15800,N_15394,N_15526);
and U15801 (N_15801,N_15300,N_15009);
nor U15802 (N_15802,N_15344,N_15484);
or U15803 (N_15803,N_15232,N_15061);
nand U15804 (N_15804,N_15176,N_15127);
xnor U15805 (N_15805,N_15405,N_15017);
or U15806 (N_15806,N_15236,N_15278);
nor U15807 (N_15807,N_15245,N_15239);
and U15808 (N_15808,N_15015,N_15014);
and U15809 (N_15809,N_15581,N_15284);
nand U15810 (N_15810,N_15053,N_15069);
and U15811 (N_15811,N_15223,N_15184);
nor U15812 (N_15812,N_15091,N_15406);
nand U15813 (N_15813,N_15001,N_15106);
nor U15814 (N_15814,N_15452,N_15049);
or U15815 (N_15815,N_15130,N_15613);
or U15816 (N_15816,N_15529,N_15103);
nand U15817 (N_15817,N_15006,N_15567);
and U15818 (N_15818,N_15525,N_15607);
nand U15819 (N_15819,N_15372,N_15564);
or U15820 (N_15820,N_15078,N_15376);
or U15821 (N_15821,N_15271,N_15418);
xnor U15822 (N_15822,N_15431,N_15153);
or U15823 (N_15823,N_15466,N_15002);
nor U15824 (N_15824,N_15283,N_15249);
nand U15825 (N_15825,N_15336,N_15039);
nand U15826 (N_15826,N_15556,N_15412);
and U15827 (N_15827,N_15441,N_15251);
or U15828 (N_15828,N_15589,N_15311);
nand U15829 (N_15829,N_15310,N_15034);
nor U15830 (N_15830,N_15328,N_15424);
nor U15831 (N_15831,N_15075,N_15137);
or U15832 (N_15832,N_15587,N_15156);
and U15833 (N_15833,N_15428,N_15605);
or U15834 (N_15834,N_15118,N_15353);
or U15835 (N_15835,N_15062,N_15040);
nor U15836 (N_15836,N_15599,N_15621);
nand U15837 (N_15837,N_15302,N_15077);
nand U15838 (N_15838,N_15164,N_15307);
xnor U15839 (N_15839,N_15007,N_15191);
nor U15840 (N_15840,N_15125,N_15279);
and U15841 (N_15841,N_15019,N_15238);
xnor U15842 (N_15842,N_15321,N_15093);
nor U15843 (N_15843,N_15401,N_15555);
or U15844 (N_15844,N_15052,N_15145);
and U15845 (N_15845,N_15285,N_15414);
or U15846 (N_15846,N_15411,N_15054);
or U15847 (N_15847,N_15576,N_15109);
nor U15848 (N_15848,N_15226,N_15360);
or U15849 (N_15849,N_15430,N_15461);
or U15850 (N_15850,N_15222,N_15611);
nor U15851 (N_15851,N_15163,N_15361);
or U15852 (N_15852,N_15499,N_15199);
and U15853 (N_15853,N_15472,N_15469);
nor U15854 (N_15854,N_15339,N_15008);
and U15855 (N_15855,N_15166,N_15602);
nand U15856 (N_15856,N_15566,N_15277);
nand U15857 (N_15857,N_15074,N_15123);
nand U15858 (N_15858,N_15139,N_15463);
and U15859 (N_15859,N_15033,N_15179);
xnor U15860 (N_15860,N_15348,N_15509);
nor U15861 (N_15861,N_15064,N_15550);
and U15862 (N_15862,N_15591,N_15573);
nand U15863 (N_15863,N_15482,N_15225);
or U15864 (N_15864,N_15369,N_15193);
and U15865 (N_15865,N_15202,N_15449);
and U15866 (N_15866,N_15460,N_15094);
nor U15867 (N_15867,N_15201,N_15173);
nor U15868 (N_15868,N_15190,N_15265);
or U15869 (N_15869,N_15358,N_15080);
nand U15870 (N_15870,N_15397,N_15385);
nand U15871 (N_15871,N_15235,N_15301);
nor U15872 (N_15872,N_15318,N_15432);
nor U15873 (N_15873,N_15110,N_15004);
nand U15874 (N_15874,N_15146,N_15345);
nor U15875 (N_15875,N_15562,N_15539);
nand U15876 (N_15876,N_15095,N_15349);
nand U15877 (N_15877,N_15519,N_15186);
nor U15878 (N_15878,N_15337,N_15527);
and U15879 (N_15879,N_15346,N_15559);
nand U15880 (N_15880,N_15213,N_15333);
or U15881 (N_15881,N_15354,N_15475);
xnor U15882 (N_15882,N_15096,N_15204);
xor U15883 (N_15883,N_15362,N_15342);
nand U15884 (N_15884,N_15090,N_15437);
nand U15885 (N_15885,N_15149,N_15377);
xnor U15886 (N_15886,N_15549,N_15117);
and U15887 (N_15887,N_15129,N_15391);
or U15888 (N_15888,N_15456,N_15508);
nor U15889 (N_15889,N_15486,N_15161);
nand U15890 (N_15890,N_15038,N_15252);
nor U15891 (N_15891,N_15427,N_15429);
nor U15892 (N_15892,N_15523,N_15609);
and U15893 (N_15893,N_15536,N_15219);
nand U15894 (N_15894,N_15066,N_15393);
nor U15895 (N_15895,N_15026,N_15037);
nor U15896 (N_15896,N_15537,N_15030);
and U15897 (N_15897,N_15408,N_15331);
nor U15898 (N_15898,N_15470,N_15294);
or U15899 (N_15899,N_15558,N_15533);
or U15900 (N_15900,N_15396,N_15207);
nand U15901 (N_15901,N_15072,N_15229);
and U15902 (N_15902,N_15436,N_15510);
and U15903 (N_15903,N_15324,N_15027);
and U15904 (N_15904,N_15444,N_15503);
xor U15905 (N_15905,N_15154,N_15063);
nor U15906 (N_15906,N_15248,N_15042);
or U15907 (N_15907,N_15268,N_15114);
nand U15908 (N_15908,N_15046,N_15435);
nor U15909 (N_15909,N_15151,N_15365);
nor U15910 (N_15910,N_15495,N_15543);
or U15911 (N_15911,N_15541,N_15259);
and U15912 (N_15912,N_15013,N_15242);
and U15913 (N_15913,N_15165,N_15417);
nand U15914 (N_15914,N_15303,N_15450);
or U15915 (N_15915,N_15087,N_15101);
xor U15916 (N_15916,N_15058,N_15506);
nor U15917 (N_15917,N_15491,N_15256);
and U15918 (N_15918,N_15481,N_15135);
nor U15919 (N_15919,N_15610,N_15297);
nor U15920 (N_15920,N_15563,N_15155);
nand U15921 (N_15921,N_15289,N_15306);
xor U15922 (N_15922,N_15282,N_15375);
or U15923 (N_15923,N_15588,N_15286);
nor U15924 (N_15924,N_15230,N_15020);
nand U15925 (N_15925,N_15022,N_15287);
nand U15926 (N_15926,N_15575,N_15538);
nand U15927 (N_15927,N_15050,N_15413);
nand U15928 (N_15928,N_15381,N_15403);
and U15929 (N_15929,N_15517,N_15593);
nand U15930 (N_15930,N_15120,N_15586);
nand U15931 (N_15931,N_15140,N_15076);
nor U15932 (N_15932,N_15528,N_15402);
nor U15933 (N_15933,N_15330,N_15504);
nand U15934 (N_15934,N_15352,N_15464);
and U15935 (N_15935,N_15458,N_15494);
nor U15936 (N_15936,N_15520,N_15024);
xnor U15937 (N_15937,N_15313,N_15276);
nand U15938 (N_15938,N_15345,N_15606);
nor U15939 (N_15939,N_15064,N_15518);
or U15940 (N_15940,N_15568,N_15443);
nand U15941 (N_15941,N_15476,N_15234);
xor U15942 (N_15942,N_15452,N_15092);
xor U15943 (N_15943,N_15376,N_15440);
nand U15944 (N_15944,N_15177,N_15550);
and U15945 (N_15945,N_15170,N_15209);
nand U15946 (N_15946,N_15104,N_15457);
xor U15947 (N_15947,N_15019,N_15489);
and U15948 (N_15948,N_15451,N_15088);
or U15949 (N_15949,N_15062,N_15350);
nand U15950 (N_15950,N_15456,N_15067);
nand U15951 (N_15951,N_15171,N_15448);
and U15952 (N_15952,N_15018,N_15329);
nor U15953 (N_15953,N_15503,N_15162);
nand U15954 (N_15954,N_15364,N_15160);
nand U15955 (N_15955,N_15052,N_15233);
or U15956 (N_15956,N_15241,N_15252);
xnor U15957 (N_15957,N_15505,N_15349);
or U15958 (N_15958,N_15308,N_15510);
and U15959 (N_15959,N_15600,N_15375);
or U15960 (N_15960,N_15274,N_15325);
or U15961 (N_15961,N_15066,N_15173);
nand U15962 (N_15962,N_15614,N_15266);
or U15963 (N_15963,N_15577,N_15239);
nand U15964 (N_15964,N_15591,N_15105);
or U15965 (N_15965,N_15362,N_15144);
xnor U15966 (N_15966,N_15192,N_15090);
xnor U15967 (N_15967,N_15431,N_15492);
nand U15968 (N_15968,N_15250,N_15291);
and U15969 (N_15969,N_15570,N_15590);
and U15970 (N_15970,N_15035,N_15427);
nand U15971 (N_15971,N_15120,N_15485);
nor U15972 (N_15972,N_15605,N_15017);
nor U15973 (N_15973,N_15444,N_15054);
or U15974 (N_15974,N_15098,N_15029);
nor U15975 (N_15975,N_15350,N_15166);
and U15976 (N_15976,N_15534,N_15015);
or U15977 (N_15977,N_15494,N_15296);
and U15978 (N_15978,N_15085,N_15297);
xor U15979 (N_15979,N_15108,N_15051);
nor U15980 (N_15980,N_15027,N_15059);
nand U15981 (N_15981,N_15344,N_15115);
nor U15982 (N_15982,N_15262,N_15534);
xnor U15983 (N_15983,N_15394,N_15044);
nor U15984 (N_15984,N_15170,N_15364);
nor U15985 (N_15985,N_15385,N_15594);
nor U15986 (N_15986,N_15298,N_15238);
nor U15987 (N_15987,N_15143,N_15517);
xor U15988 (N_15988,N_15097,N_15395);
or U15989 (N_15989,N_15420,N_15167);
or U15990 (N_15990,N_15503,N_15332);
nand U15991 (N_15991,N_15359,N_15617);
nand U15992 (N_15992,N_15619,N_15551);
nand U15993 (N_15993,N_15270,N_15191);
and U15994 (N_15994,N_15365,N_15441);
xnor U15995 (N_15995,N_15340,N_15321);
nor U15996 (N_15996,N_15461,N_15121);
nor U15997 (N_15997,N_15178,N_15164);
xnor U15998 (N_15998,N_15322,N_15622);
nor U15999 (N_15999,N_15488,N_15598);
nor U16000 (N_16000,N_15162,N_15426);
nand U16001 (N_16001,N_15311,N_15197);
nand U16002 (N_16002,N_15513,N_15202);
nor U16003 (N_16003,N_15006,N_15163);
nand U16004 (N_16004,N_15095,N_15226);
and U16005 (N_16005,N_15121,N_15460);
and U16006 (N_16006,N_15502,N_15498);
nand U16007 (N_16007,N_15490,N_15137);
or U16008 (N_16008,N_15095,N_15599);
nor U16009 (N_16009,N_15269,N_15233);
or U16010 (N_16010,N_15160,N_15298);
nand U16011 (N_16011,N_15173,N_15083);
or U16012 (N_16012,N_15565,N_15548);
nand U16013 (N_16013,N_15059,N_15294);
xor U16014 (N_16014,N_15516,N_15618);
and U16015 (N_16015,N_15476,N_15132);
nor U16016 (N_16016,N_15089,N_15085);
and U16017 (N_16017,N_15359,N_15189);
nor U16018 (N_16018,N_15134,N_15014);
or U16019 (N_16019,N_15212,N_15452);
nor U16020 (N_16020,N_15623,N_15600);
nor U16021 (N_16021,N_15238,N_15046);
nand U16022 (N_16022,N_15365,N_15535);
xor U16023 (N_16023,N_15425,N_15381);
or U16024 (N_16024,N_15425,N_15608);
or U16025 (N_16025,N_15431,N_15132);
nand U16026 (N_16026,N_15111,N_15281);
nand U16027 (N_16027,N_15481,N_15408);
and U16028 (N_16028,N_15064,N_15285);
nand U16029 (N_16029,N_15008,N_15524);
or U16030 (N_16030,N_15384,N_15428);
or U16031 (N_16031,N_15487,N_15362);
nor U16032 (N_16032,N_15389,N_15383);
and U16033 (N_16033,N_15575,N_15076);
nand U16034 (N_16034,N_15304,N_15226);
nor U16035 (N_16035,N_15296,N_15282);
or U16036 (N_16036,N_15053,N_15476);
xnor U16037 (N_16037,N_15334,N_15129);
and U16038 (N_16038,N_15465,N_15101);
nand U16039 (N_16039,N_15398,N_15531);
nand U16040 (N_16040,N_15591,N_15482);
nand U16041 (N_16041,N_15479,N_15449);
or U16042 (N_16042,N_15569,N_15454);
nor U16043 (N_16043,N_15092,N_15300);
nand U16044 (N_16044,N_15328,N_15364);
nor U16045 (N_16045,N_15023,N_15528);
or U16046 (N_16046,N_15176,N_15295);
xnor U16047 (N_16047,N_15162,N_15160);
xor U16048 (N_16048,N_15074,N_15169);
nor U16049 (N_16049,N_15176,N_15045);
nand U16050 (N_16050,N_15242,N_15540);
and U16051 (N_16051,N_15193,N_15447);
or U16052 (N_16052,N_15136,N_15117);
nand U16053 (N_16053,N_15347,N_15516);
nor U16054 (N_16054,N_15182,N_15609);
nand U16055 (N_16055,N_15426,N_15590);
or U16056 (N_16056,N_15414,N_15401);
nor U16057 (N_16057,N_15617,N_15143);
nor U16058 (N_16058,N_15209,N_15457);
nor U16059 (N_16059,N_15298,N_15215);
nor U16060 (N_16060,N_15266,N_15000);
nand U16061 (N_16061,N_15574,N_15373);
nand U16062 (N_16062,N_15015,N_15433);
or U16063 (N_16063,N_15048,N_15582);
or U16064 (N_16064,N_15533,N_15211);
nand U16065 (N_16065,N_15333,N_15288);
nand U16066 (N_16066,N_15010,N_15241);
and U16067 (N_16067,N_15302,N_15622);
nand U16068 (N_16068,N_15481,N_15177);
nand U16069 (N_16069,N_15365,N_15113);
or U16070 (N_16070,N_15274,N_15429);
and U16071 (N_16071,N_15014,N_15313);
nand U16072 (N_16072,N_15312,N_15440);
or U16073 (N_16073,N_15298,N_15025);
or U16074 (N_16074,N_15127,N_15479);
nand U16075 (N_16075,N_15490,N_15232);
and U16076 (N_16076,N_15301,N_15537);
or U16077 (N_16077,N_15221,N_15064);
nand U16078 (N_16078,N_15180,N_15326);
or U16079 (N_16079,N_15007,N_15017);
and U16080 (N_16080,N_15018,N_15317);
and U16081 (N_16081,N_15433,N_15027);
nor U16082 (N_16082,N_15035,N_15552);
nand U16083 (N_16083,N_15580,N_15541);
and U16084 (N_16084,N_15509,N_15469);
nand U16085 (N_16085,N_15585,N_15309);
and U16086 (N_16086,N_15421,N_15019);
nand U16087 (N_16087,N_15451,N_15464);
xnor U16088 (N_16088,N_15080,N_15273);
nor U16089 (N_16089,N_15034,N_15000);
and U16090 (N_16090,N_15225,N_15058);
and U16091 (N_16091,N_15082,N_15543);
nor U16092 (N_16092,N_15264,N_15562);
or U16093 (N_16093,N_15446,N_15182);
xor U16094 (N_16094,N_15186,N_15497);
nor U16095 (N_16095,N_15082,N_15406);
nor U16096 (N_16096,N_15341,N_15423);
nor U16097 (N_16097,N_15408,N_15227);
nor U16098 (N_16098,N_15391,N_15331);
and U16099 (N_16099,N_15100,N_15446);
nor U16100 (N_16100,N_15190,N_15536);
or U16101 (N_16101,N_15546,N_15187);
or U16102 (N_16102,N_15117,N_15023);
nor U16103 (N_16103,N_15497,N_15200);
nand U16104 (N_16104,N_15414,N_15399);
or U16105 (N_16105,N_15531,N_15307);
xor U16106 (N_16106,N_15482,N_15558);
nor U16107 (N_16107,N_15017,N_15332);
nand U16108 (N_16108,N_15230,N_15539);
and U16109 (N_16109,N_15417,N_15476);
nor U16110 (N_16110,N_15302,N_15135);
and U16111 (N_16111,N_15399,N_15154);
and U16112 (N_16112,N_15454,N_15206);
or U16113 (N_16113,N_15227,N_15138);
and U16114 (N_16114,N_15400,N_15353);
and U16115 (N_16115,N_15300,N_15374);
xor U16116 (N_16116,N_15602,N_15208);
nor U16117 (N_16117,N_15551,N_15022);
nor U16118 (N_16118,N_15327,N_15339);
nor U16119 (N_16119,N_15032,N_15440);
xnor U16120 (N_16120,N_15296,N_15406);
or U16121 (N_16121,N_15466,N_15359);
or U16122 (N_16122,N_15447,N_15569);
nor U16123 (N_16123,N_15353,N_15361);
or U16124 (N_16124,N_15021,N_15354);
nand U16125 (N_16125,N_15117,N_15267);
nand U16126 (N_16126,N_15001,N_15502);
and U16127 (N_16127,N_15524,N_15198);
and U16128 (N_16128,N_15461,N_15359);
nor U16129 (N_16129,N_15223,N_15285);
and U16130 (N_16130,N_15454,N_15539);
or U16131 (N_16131,N_15539,N_15102);
xor U16132 (N_16132,N_15262,N_15238);
or U16133 (N_16133,N_15174,N_15605);
or U16134 (N_16134,N_15162,N_15306);
and U16135 (N_16135,N_15136,N_15554);
nor U16136 (N_16136,N_15316,N_15598);
and U16137 (N_16137,N_15226,N_15402);
and U16138 (N_16138,N_15579,N_15467);
nand U16139 (N_16139,N_15473,N_15464);
nor U16140 (N_16140,N_15134,N_15613);
and U16141 (N_16141,N_15084,N_15434);
or U16142 (N_16142,N_15504,N_15160);
nor U16143 (N_16143,N_15113,N_15408);
nor U16144 (N_16144,N_15402,N_15612);
nand U16145 (N_16145,N_15414,N_15148);
nor U16146 (N_16146,N_15204,N_15399);
nand U16147 (N_16147,N_15100,N_15371);
nor U16148 (N_16148,N_15227,N_15494);
or U16149 (N_16149,N_15295,N_15593);
and U16150 (N_16150,N_15494,N_15243);
and U16151 (N_16151,N_15160,N_15143);
nand U16152 (N_16152,N_15521,N_15063);
and U16153 (N_16153,N_15591,N_15107);
and U16154 (N_16154,N_15328,N_15075);
nor U16155 (N_16155,N_15523,N_15455);
and U16156 (N_16156,N_15320,N_15342);
and U16157 (N_16157,N_15432,N_15168);
and U16158 (N_16158,N_15066,N_15563);
nor U16159 (N_16159,N_15154,N_15064);
xnor U16160 (N_16160,N_15142,N_15149);
nand U16161 (N_16161,N_15351,N_15212);
and U16162 (N_16162,N_15317,N_15273);
and U16163 (N_16163,N_15503,N_15401);
and U16164 (N_16164,N_15293,N_15153);
nand U16165 (N_16165,N_15277,N_15537);
nand U16166 (N_16166,N_15296,N_15027);
or U16167 (N_16167,N_15460,N_15020);
and U16168 (N_16168,N_15262,N_15572);
nor U16169 (N_16169,N_15407,N_15396);
or U16170 (N_16170,N_15125,N_15365);
and U16171 (N_16171,N_15114,N_15063);
or U16172 (N_16172,N_15312,N_15063);
nor U16173 (N_16173,N_15453,N_15358);
nor U16174 (N_16174,N_15005,N_15309);
nor U16175 (N_16175,N_15403,N_15460);
or U16176 (N_16176,N_15213,N_15214);
nand U16177 (N_16177,N_15514,N_15179);
nand U16178 (N_16178,N_15369,N_15387);
and U16179 (N_16179,N_15343,N_15131);
nor U16180 (N_16180,N_15242,N_15081);
xnor U16181 (N_16181,N_15118,N_15369);
or U16182 (N_16182,N_15141,N_15172);
and U16183 (N_16183,N_15444,N_15226);
nor U16184 (N_16184,N_15516,N_15435);
xnor U16185 (N_16185,N_15607,N_15441);
nand U16186 (N_16186,N_15587,N_15134);
nor U16187 (N_16187,N_15389,N_15147);
nand U16188 (N_16188,N_15247,N_15407);
nand U16189 (N_16189,N_15229,N_15359);
or U16190 (N_16190,N_15431,N_15310);
and U16191 (N_16191,N_15142,N_15150);
nand U16192 (N_16192,N_15490,N_15277);
xor U16193 (N_16193,N_15611,N_15246);
nand U16194 (N_16194,N_15162,N_15226);
and U16195 (N_16195,N_15431,N_15064);
and U16196 (N_16196,N_15152,N_15248);
or U16197 (N_16197,N_15480,N_15091);
xnor U16198 (N_16198,N_15282,N_15194);
and U16199 (N_16199,N_15040,N_15082);
and U16200 (N_16200,N_15249,N_15030);
xor U16201 (N_16201,N_15449,N_15089);
and U16202 (N_16202,N_15304,N_15079);
or U16203 (N_16203,N_15451,N_15216);
or U16204 (N_16204,N_15343,N_15203);
nor U16205 (N_16205,N_15365,N_15526);
or U16206 (N_16206,N_15447,N_15553);
nand U16207 (N_16207,N_15516,N_15025);
and U16208 (N_16208,N_15440,N_15439);
nand U16209 (N_16209,N_15473,N_15492);
nand U16210 (N_16210,N_15135,N_15227);
nor U16211 (N_16211,N_15495,N_15385);
nand U16212 (N_16212,N_15159,N_15275);
and U16213 (N_16213,N_15620,N_15148);
nand U16214 (N_16214,N_15059,N_15221);
or U16215 (N_16215,N_15013,N_15272);
and U16216 (N_16216,N_15476,N_15126);
nand U16217 (N_16217,N_15020,N_15488);
and U16218 (N_16218,N_15062,N_15494);
nor U16219 (N_16219,N_15236,N_15177);
xor U16220 (N_16220,N_15351,N_15603);
and U16221 (N_16221,N_15373,N_15559);
xor U16222 (N_16222,N_15412,N_15580);
nand U16223 (N_16223,N_15216,N_15000);
nand U16224 (N_16224,N_15154,N_15153);
and U16225 (N_16225,N_15152,N_15120);
and U16226 (N_16226,N_15243,N_15302);
or U16227 (N_16227,N_15122,N_15423);
or U16228 (N_16228,N_15435,N_15595);
nor U16229 (N_16229,N_15095,N_15207);
or U16230 (N_16230,N_15611,N_15056);
nor U16231 (N_16231,N_15369,N_15417);
nor U16232 (N_16232,N_15148,N_15065);
and U16233 (N_16233,N_15368,N_15360);
nand U16234 (N_16234,N_15041,N_15499);
or U16235 (N_16235,N_15387,N_15197);
nand U16236 (N_16236,N_15455,N_15245);
nand U16237 (N_16237,N_15275,N_15368);
nor U16238 (N_16238,N_15136,N_15482);
nor U16239 (N_16239,N_15263,N_15016);
and U16240 (N_16240,N_15253,N_15275);
and U16241 (N_16241,N_15161,N_15032);
nor U16242 (N_16242,N_15324,N_15171);
and U16243 (N_16243,N_15573,N_15297);
nand U16244 (N_16244,N_15181,N_15521);
xnor U16245 (N_16245,N_15316,N_15511);
nand U16246 (N_16246,N_15209,N_15355);
or U16247 (N_16247,N_15374,N_15452);
or U16248 (N_16248,N_15294,N_15408);
nor U16249 (N_16249,N_15113,N_15586);
nand U16250 (N_16250,N_15896,N_15841);
nor U16251 (N_16251,N_16042,N_15850);
or U16252 (N_16252,N_15752,N_16019);
nor U16253 (N_16253,N_15744,N_16211);
nand U16254 (N_16254,N_15871,N_15929);
nand U16255 (N_16255,N_15989,N_15703);
nor U16256 (N_16256,N_15666,N_15658);
xor U16257 (N_16257,N_15971,N_16061);
nor U16258 (N_16258,N_16141,N_15980);
nand U16259 (N_16259,N_16164,N_16009);
nor U16260 (N_16260,N_15751,N_16246);
nand U16261 (N_16261,N_16007,N_15722);
or U16262 (N_16262,N_16182,N_15735);
and U16263 (N_16263,N_15996,N_16068);
or U16264 (N_16264,N_16233,N_16113);
and U16265 (N_16265,N_15922,N_16112);
and U16266 (N_16266,N_15970,N_15713);
and U16267 (N_16267,N_15978,N_15808);
nor U16268 (N_16268,N_16193,N_15824);
xor U16269 (N_16269,N_15910,N_16088);
or U16270 (N_16270,N_15914,N_16210);
and U16271 (N_16271,N_15801,N_16011);
or U16272 (N_16272,N_15899,N_15763);
xor U16273 (N_16273,N_15927,N_15721);
or U16274 (N_16274,N_15845,N_15687);
and U16275 (N_16275,N_16216,N_15738);
or U16276 (N_16276,N_16067,N_15962);
and U16277 (N_16277,N_15895,N_16109);
xor U16278 (N_16278,N_15965,N_15985);
or U16279 (N_16279,N_15657,N_16097);
or U16280 (N_16280,N_15844,N_16077);
xor U16281 (N_16281,N_16179,N_15660);
and U16282 (N_16282,N_15832,N_15955);
and U16283 (N_16283,N_16059,N_15884);
nor U16284 (N_16284,N_15685,N_15973);
nand U16285 (N_16285,N_16010,N_15785);
or U16286 (N_16286,N_15644,N_16188);
nand U16287 (N_16287,N_15793,N_15692);
or U16288 (N_16288,N_15662,N_16227);
or U16289 (N_16289,N_15696,N_15786);
and U16290 (N_16290,N_16021,N_16041);
and U16291 (N_16291,N_15982,N_15745);
xnor U16292 (N_16292,N_15717,N_16015);
and U16293 (N_16293,N_16121,N_15648);
and U16294 (N_16294,N_15689,N_16118);
nor U16295 (N_16295,N_15716,N_15736);
nand U16296 (N_16296,N_15676,N_15972);
nor U16297 (N_16297,N_16034,N_15647);
and U16298 (N_16298,N_15931,N_15852);
and U16299 (N_16299,N_16214,N_16157);
and U16300 (N_16300,N_16129,N_16110);
and U16301 (N_16301,N_15788,N_15942);
nor U16302 (N_16302,N_16160,N_16050);
nand U16303 (N_16303,N_16238,N_15774);
nand U16304 (N_16304,N_15649,N_16000);
or U16305 (N_16305,N_15748,N_15819);
xnor U16306 (N_16306,N_16151,N_16229);
nand U16307 (N_16307,N_15946,N_16114);
or U16308 (N_16308,N_15723,N_16090);
nor U16309 (N_16309,N_16092,N_15809);
xnor U16310 (N_16310,N_16140,N_15961);
or U16311 (N_16311,N_16029,N_15963);
nor U16312 (N_16312,N_15878,N_16071);
nand U16313 (N_16313,N_16069,N_16087);
nor U16314 (N_16314,N_15737,N_15883);
nand U16315 (N_16315,N_16091,N_15995);
nor U16316 (N_16316,N_16076,N_15664);
nor U16317 (N_16317,N_15901,N_16155);
or U16318 (N_16318,N_16190,N_16247);
nor U16319 (N_16319,N_15755,N_16014);
or U16320 (N_16320,N_15756,N_15966);
or U16321 (N_16321,N_15759,N_16181);
and U16322 (N_16322,N_15853,N_16171);
nand U16323 (N_16323,N_16205,N_15794);
nor U16324 (N_16324,N_15939,N_15903);
and U16325 (N_16325,N_16230,N_15943);
or U16326 (N_16326,N_15925,N_15694);
or U16327 (N_16327,N_15987,N_16082);
nor U16328 (N_16328,N_16107,N_15829);
or U16329 (N_16329,N_15906,N_16184);
nand U16330 (N_16330,N_15765,N_16131);
and U16331 (N_16331,N_16146,N_16116);
nor U16332 (N_16332,N_15706,N_16200);
nor U16333 (N_16333,N_15754,N_15678);
nand U16334 (N_16334,N_15947,N_16203);
or U16335 (N_16335,N_16186,N_16167);
nor U16336 (N_16336,N_15673,N_15761);
nand U16337 (N_16337,N_15650,N_16185);
nor U16338 (N_16338,N_16183,N_15839);
and U16339 (N_16339,N_16150,N_15792);
or U16340 (N_16340,N_16040,N_16108);
and U16341 (N_16341,N_15731,N_16066);
and U16342 (N_16342,N_16248,N_16224);
nor U16343 (N_16343,N_15861,N_16045);
xor U16344 (N_16344,N_15799,N_16030);
and U16345 (N_16345,N_16031,N_15826);
nand U16346 (N_16346,N_15636,N_15770);
nand U16347 (N_16347,N_15710,N_15767);
and U16348 (N_16348,N_15828,N_15905);
nand U16349 (N_16349,N_16051,N_16174);
or U16350 (N_16350,N_15881,N_15870);
and U16351 (N_16351,N_15697,N_15979);
or U16352 (N_16352,N_16176,N_15741);
or U16353 (N_16353,N_15693,N_15628);
xor U16354 (N_16354,N_15892,N_15632);
nor U16355 (N_16355,N_15709,N_16168);
or U16356 (N_16356,N_15969,N_15814);
nor U16357 (N_16357,N_15669,N_16062);
nor U16358 (N_16358,N_15976,N_15967);
nand U16359 (N_16359,N_16012,N_15911);
and U16360 (N_16360,N_15919,N_16145);
or U16361 (N_16361,N_16212,N_15886);
nand U16362 (N_16362,N_15997,N_16132);
nand U16363 (N_16363,N_16208,N_15683);
or U16364 (N_16364,N_16104,N_15672);
nand U16365 (N_16365,N_15728,N_15775);
or U16366 (N_16366,N_15633,N_15798);
or U16367 (N_16367,N_15642,N_15981);
nand U16368 (N_16368,N_16102,N_15827);
or U16369 (N_16369,N_15749,N_15637);
nand U16370 (N_16370,N_16004,N_15912);
nor U16371 (N_16371,N_15806,N_15695);
nor U16372 (N_16372,N_15780,N_15953);
xor U16373 (N_16373,N_15783,N_15900);
xor U16374 (N_16374,N_15958,N_16197);
nor U16375 (N_16375,N_16024,N_15708);
or U16376 (N_16376,N_15630,N_15830);
nor U16377 (N_16377,N_15791,N_16046);
xnor U16378 (N_16378,N_15872,N_15629);
nand U16379 (N_16379,N_16038,N_15859);
nand U16380 (N_16380,N_16119,N_16135);
or U16381 (N_16381,N_16003,N_15908);
or U16382 (N_16382,N_15818,N_15860);
and U16383 (N_16383,N_15627,N_15864);
and U16384 (N_16384,N_15994,N_15638);
or U16385 (N_16385,N_15777,N_15807);
nand U16386 (N_16386,N_15984,N_15877);
xnor U16387 (N_16387,N_15890,N_16219);
or U16388 (N_16388,N_16133,N_15952);
nor U16389 (N_16389,N_16232,N_15889);
nand U16390 (N_16390,N_15677,N_16234);
xor U16391 (N_16391,N_16039,N_15804);
nand U16392 (N_16392,N_16023,N_15940);
nor U16393 (N_16393,N_15838,N_16178);
or U16394 (N_16394,N_15885,N_15837);
and U16395 (N_16395,N_16189,N_15945);
or U16396 (N_16396,N_16101,N_15776);
or U16397 (N_16397,N_16032,N_16073);
nor U16398 (N_16398,N_15724,N_15817);
or U16399 (N_16399,N_15702,N_15730);
and U16400 (N_16400,N_15897,N_16242);
or U16401 (N_16401,N_15862,N_16228);
nand U16402 (N_16402,N_15941,N_15773);
and U16403 (N_16403,N_15974,N_15848);
nor U16404 (N_16404,N_15868,N_15812);
or U16405 (N_16405,N_16147,N_15949);
or U16406 (N_16406,N_16134,N_16136);
nand U16407 (N_16407,N_15986,N_15951);
nor U16408 (N_16408,N_16037,N_16152);
nor U16409 (N_16409,N_16165,N_15671);
nand U16410 (N_16410,N_15691,N_16064);
xor U16411 (N_16411,N_16063,N_15879);
or U16412 (N_16412,N_15968,N_15656);
and U16413 (N_16413,N_15880,N_15831);
nand U16414 (N_16414,N_15909,N_15936);
or U16415 (N_16415,N_15932,N_15681);
and U16416 (N_16416,N_15990,N_15639);
and U16417 (N_16417,N_15787,N_16047);
or U16418 (N_16418,N_16222,N_16106);
nor U16419 (N_16419,N_16244,N_15813);
nor U16420 (N_16420,N_15651,N_15757);
or U16421 (N_16421,N_16079,N_16142);
nand U16422 (N_16422,N_15934,N_16033);
and U16423 (N_16423,N_16055,N_16199);
nand U16424 (N_16424,N_15954,N_16156);
or U16425 (N_16425,N_16093,N_16209);
nand U16426 (N_16426,N_16060,N_16139);
nor U16427 (N_16427,N_15840,N_15805);
nor U16428 (N_16428,N_15933,N_15999);
or U16429 (N_16429,N_15641,N_16169);
and U16430 (N_16430,N_15904,N_16043);
or U16431 (N_16431,N_15668,N_16100);
nor U16432 (N_16432,N_15779,N_16235);
xor U16433 (N_16433,N_15843,N_15882);
nor U16434 (N_16434,N_16008,N_15790);
nor U16435 (N_16435,N_15680,N_15816);
or U16436 (N_16436,N_15898,N_16125);
nor U16437 (N_16437,N_15873,N_15795);
and U16438 (N_16438,N_16163,N_15729);
nor U16439 (N_16439,N_15869,N_16245);
nand U16440 (N_16440,N_15701,N_16027);
or U16441 (N_16441,N_16220,N_15825);
xnor U16442 (N_16442,N_16215,N_15907);
and U16443 (N_16443,N_16127,N_15916);
nand U16444 (N_16444,N_16162,N_15854);
nor U16445 (N_16445,N_15863,N_15836);
and U16446 (N_16446,N_16124,N_15928);
and U16447 (N_16447,N_16005,N_15921);
or U16448 (N_16448,N_15867,N_16138);
nor U16449 (N_16449,N_16198,N_15690);
or U16450 (N_16450,N_16149,N_15772);
or U16451 (N_16451,N_16013,N_15714);
nor U16452 (N_16452,N_15874,N_16099);
and U16453 (N_16453,N_15959,N_15930);
xor U16454 (N_16454,N_15727,N_15719);
and U16455 (N_16455,N_16196,N_16207);
nand U16456 (N_16456,N_15802,N_15888);
and U16457 (N_16457,N_16172,N_15822);
or U16458 (N_16458,N_15771,N_15766);
xnor U16459 (N_16459,N_15700,N_15712);
nor U16460 (N_16460,N_15998,N_15920);
or U16461 (N_16461,N_16187,N_16239);
nor U16462 (N_16462,N_15820,N_16158);
nor U16463 (N_16463,N_15846,N_16217);
nor U16464 (N_16464,N_16001,N_15768);
or U16465 (N_16465,N_16225,N_15758);
xnor U16466 (N_16466,N_15688,N_15635);
or U16467 (N_16467,N_15674,N_15699);
or U16468 (N_16468,N_16115,N_15815);
or U16469 (N_16469,N_15704,N_15789);
nand U16470 (N_16470,N_15742,N_16249);
nand U16471 (N_16471,N_16006,N_15725);
or U16472 (N_16472,N_15993,N_16085);
and U16473 (N_16473,N_15856,N_15705);
nand U16474 (N_16474,N_16074,N_15964);
nor U16475 (N_16475,N_15891,N_15734);
nor U16476 (N_16476,N_15653,N_15893);
nand U16477 (N_16477,N_15800,N_16052);
and U16478 (N_16478,N_16223,N_16231);
or U16479 (N_16479,N_16170,N_15796);
xnor U16480 (N_16480,N_15740,N_16086);
nand U16481 (N_16481,N_16002,N_15847);
or U16482 (N_16482,N_16022,N_16148);
nand U16483 (N_16483,N_16128,N_16161);
nor U16484 (N_16484,N_15849,N_16080);
and U16485 (N_16485,N_16083,N_15944);
nor U16486 (N_16486,N_16123,N_15894);
nand U16487 (N_16487,N_15753,N_15926);
nand U16488 (N_16488,N_15887,N_15902);
nor U16489 (N_16489,N_16221,N_15626);
nor U16490 (N_16490,N_15631,N_16105);
and U16491 (N_16491,N_15956,N_15698);
xnor U16492 (N_16492,N_16175,N_16236);
or U16493 (N_16493,N_15917,N_16177);
and U16494 (N_16494,N_15640,N_16026);
xor U16495 (N_16495,N_16237,N_15855);
nor U16496 (N_16496,N_15983,N_15764);
xnor U16497 (N_16497,N_15747,N_15975);
xnor U16498 (N_16498,N_16194,N_15762);
nand U16499 (N_16499,N_16191,N_15937);
xor U16500 (N_16500,N_16240,N_16094);
and U16501 (N_16501,N_16057,N_15634);
nand U16502 (N_16502,N_16098,N_16078);
nor U16503 (N_16503,N_16016,N_15726);
or U16504 (N_16504,N_15865,N_16084);
or U16505 (N_16505,N_16065,N_16180);
and U16506 (N_16506,N_15643,N_15663);
or U16507 (N_16507,N_16020,N_15866);
nor U16508 (N_16508,N_16201,N_15821);
nor U16509 (N_16509,N_15733,N_15957);
xor U16510 (N_16510,N_15875,N_16025);
nand U16511 (N_16511,N_15675,N_16054);
nand U16512 (N_16512,N_15842,N_15746);
nand U16513 (N_16513,N_15670,N_16154);
nand U16514 (N_16514,N_15823,N_16120);
nor U16515 (N_16515,N_15743,N_15739);
or U16516 (N_16516,N_15778,N_16111);
nand U16517 (N_16517,N_16056,N_16058);
nor U16518 (N_16518,N_16072,N_16192);
nor U16519 (N_16519,N_16153,N_16159);
nor U16520 (N_16520,N_15991,N_16166);
nor U16521 (N_16521,N_15834,N_15718);
nor U16522 (N_16522,N_15667,N_16204);
nor U16523 (N_16523,N_15833,N_15781);
and U16524 (N_16524,N_16206,N_15858);
and U16525 (N_16525,N_16144,N_15851);
and U16526 (N_16526,N_15665,N_16089);
xor U16527 (N_16527,N_16028,N_15679);
nand U16528 (N_16528,N_15682,N_16195);
nor U16529 (N_16529,N_16143,N_16048);
or U16530 (N_16530,N_15655,N_15732);
xnor U16531 (N_16531,N_16117,N_15769);
nand U16532 (N_16532,N_15782,N_16018);
or U16533 (N_16533,N_15950,N_16218);
xnor U16534 (N_16534,N_15645,N_16137);
nor U16535 (N_16535,N_16017,N_16035);
nand U16536 (N_16536,N_15835,N_16243);
nor U16537 (N_16537,N_16095,N_16036);
nor U16538 (N_16538,N_15686,N_15988);
and U16539 (N_16539,N_16241,N_16213);
nand U16540 (N_16540,N_15810,N_16122);
or U16541 (N_16541,N_15811,N_16096);
nor U16542 (N_16542,N_15923,N_15652);
and U16543 (N_16543,N_16053,N_15857);
nor U16544 (N_16544,N_15915,N_16226);
or U16545 (N_16545,N_16202,N_16103);
nor U16546 (N_16546,N_15646,N_15992);
and U16547 (N_16547,N_15918,N_15625);
nor U16548 (N_16548,N_15720,N_15654);
or U16549 (N_16549,N_16070,N_15661);
nor U16550 (N_16550,N_16126,N_15760);
nand U16551 (N_16551,N_16049,N_16075);
and U16552 (N_16552,N_15684,N_15977);
nor U16553 (N_16553,N_15797,N_15707);
nor U16554 (N_16554,N_15711,N_15935);
xnor U16555 (N_16555,N_16081,N_15876);
nor U16556 (N_16556,N_15715,N_15784);
and U16557 (N_16557,N_15803,N_15750);
nor U16558 (N_16558,N_15960,N_16130);
and U16559 (N_16559,N_15659,N_15938);
nand U16560 (N_16560,N_15924,N_15948);
nand U16561 (N_16561,N_16044,N_16173);
nor U16562 (N_16562,N_15913,N_15889);
or U16563 (N_16563,N_15812,N_16129);
and U16564 (N_16564,N_15658,N_15716);
nand U16565 (N_16565,N_16163,N_15914);
nor U16566 (N_16566,N_15890,N_15732);
and U16567 (N_16567,N_15683,N_16089);
and U16568 (N_16568,N_15945,N_15725);
nand U16569 (N_16569,N_15994,N_16207);
and U16570 (N_16570,N_16134,N_15804);
nand U16571 (N_16571,N_15915,N_15665);
and U16572 (N_16572,N_16029,N_15798);
or U16573 (N_16573,N_16028,N_15785);
nand U16574 (N_16574,N_15989,N_16196);
nand U16575 (N_16575,N_15935,N_16094);
nor U16576 (N_16576,N_16182,N_15627);
and U16577 (N_16577,N_15667,N_15681);
or U16578 (N_16578,N_15986,N_16107);
xnor U16579 (N_16579,N_15683,N_15627);
nor U16580 (N_16580,N_16116,N_15916);
nand U16581 (N_16581,N_15832,N_16003);
and U16582 (N_16582,N_15812,N_16057);
nor U16583 (N_16583,N_15633,N_15879);
nor U16584 (N_16584,N_16186,N_15663);
or U16585 (N_16585,N_15952,N_16078);
or U16586 (N_16586,N_16055,N_15759);
or U16587 (N_16587,N_15958,N_16068);
nor U16588 (N_16588,N_15840,N_15933);
and U16589 (N_16589,N_16056,N_15851);
xor U16590 (N_16590,N_15887,N_15994);
and U16591 (N_16591,N_15668,N_15973);
xnor U16592 (N_16592,N_15762,N_15780);
nor U16593 (N_16593,N_16200,N_15757);
nand U16594 (N_16594,N_15882,N_15643);
nor U16595 (N_16595,N_15855,N_15796);
and U16596 (N_16596,N_16085,N_16127);
nand U16597 (N_16597,N_16032,N_15958);
or U16598 (N_16598,N_15692,N_15924);
xnor U16599 (N_16599,N_15669,N_16184);
or U16600 (N_16600,N_15832,N_15867);
or U16601 (N_16601,N_15900,N_15772);
or U16602 (N_16602,N_15850,N_16046);
nor U16603 (N_16603,N_15890,N_16222);
and U16604 (N_16604,N_16187,N_15861);
xor U16605 (N_16605,N_15804,N_16138);
nand U16606 (N_16606,N_15942,N_15789);
nand U16607 (N_16607,N_15724,N_15956);
nand U16608 (N_16608,N_15763,N_15706);
or U16609 (N_16609,N_16011,N_15809);
nand U16610 (N_16610,N_15941,N_16087);
nand U16611 (N_16611,N_15903,N_15732);
xor U16612 (N_16612,N_15959,N_15738);
nor U16613 (N_16613,N_15743,N_16120);
nand U16614 (N_16614,N_15709,N_16188);
nand U16615 (N_16615,N_16228,N_16069);
or U16616 (N_16616,N_16041,N_15678);
or U16617 (N_16617,N_15968,N_16236);
and U16618 (N_16618,N_16151,N_15919);
or U16619 (N_16619,N_16014,N_15659);
and U16620 (N_16620,N_16148,N_15697);
nor U16621 (N_16621,N_15742,N_15770);
nand U16622 (N_16622,N_15843,N_16164);
nand U16623 (N_16623,N_15897,N_16018);
xor U16624 (N_16624,N_15828,N_16174);
and U16625 (N_16625,N_15994,N_16170);
xor U16626 (N_16626,N_15898,N_15632);
and U16627 (N_16627,N_15735,N_15919);
nor U16628 (N_16628,N_16215,N_16019);
or U16629 (N_16629,N_16091,N_15907);
nand U16630 (N_16630,N_15833,N_16065);
or U16631 (N_16631,N_16195,N_15761);
nand U16632 (N_16632,N_16054,N_16110);
nand U16633 (N_16633,N_16032,N_16069);
or U16634 (N_16634,N_15675,N_15844);
or U16635 (N_16635,N_16240,N_16203);
xor U16636 (N_16636,N_16151,N_15953);
nor U16637 (N_16637,N_15853,N_15756);
nand U16638 (N_16638,N_16143,N_16038);
and U16639 (N_16639,N_16083,N_16175);
xnor U16640 (N_16640,N_16019,N_15929);
nand U16641 (N_16641,N_16147,N_15745);
or U16642 (N_16642,N_16158,N_15896);
and U16643 (N_16643,N_15910,N_15981);
nand U16644 (N_16644,N_15846,N_15793);
nand U16645 (N_16645,N_15983,N_16128);
nand U16646 (N_16646,N_16195,N_15964);
nor U16647 (N_16647,N_15670,N_16060);
and U16648 (N_16648,N_16207,N_15641);
nand U16649 (N_16649,N_15652,N_15744);
nor U16650 (N_16650,N_15749,N_16228);
or U16651 (N_16651,N_15965,N_16018);
and U16652 (N_16652,N_15909,N_15873);
nor U16653 (N_16653,N_16076,N_15752);
xnor U16654 (N_16654,N_16140,N_15883);
or U16655 (N_16655,N_15822,N_16114);
and U16656 (N_16656,N_15641,N_16156);
or U16657 (N_16657,N_15745,N_15802);
or U16658 (N_16658,N_16023,N_15679);
nand U16659 (N_16659,N_15688,N_16174);
and U16660 (N_16660,N_15674,N_15936);
and U16661 (N_16661,N_15875,N_16074);
or U16662 (N_16662,N_15931,N_16200);
or U16663 (N_16663,N_16112,N_15862);
and U16664 (N_16664,N_15631,N_15893);
or U16665 (N_16665,N_16205,N_15709);
or U16666 (N_16666,N_15668,N_16173);
nand U16667 (N_16667,N_15783,N_15841);
or U16668 (N_16668,N_16095,N_16122);
nand U16669 (N_16669,N_16119,N_15698);
or U16670 (N_16670,N_16084,N_16063);
xor U16671 (N_16671,N_15654,N_15903);
nor U16672 (N_16672,N_16159,N_15956);
nor U16673 (N_16673,N_16128,N_16051);
nand U16674 (N_16674,N_16249,N_16013);
or U16675 (N_16675,N_15806,N_16166);
nand U16676 (N_16676,N_15808,N_16240);
and U16677 (N_16677,N_15880,N_15994);
nand U16678 (N_16678,N_15792,N_15956);
xor U16679 (N_16679,N_15626,N_16096);
nand U16680 (N_16680,N_15710,N_16191);
nand U16681 (N_16681,N_16160,N_15814);
and U16682 (N_16682,N_15644,N_15739);
xnor U16683 (N_16683,N_16031,N_16032);
and U16684 (N_16684,N_15724,N_15984);
nand U16685 (N_16685,N_15703,N_15877);
nor U16686 (N_16686,N_15628,N_16041);
or U16687 (N_16687,N_15885,N_16057);
or U16688 (N_16688,N_16128,N_15794);
or U16689 (N_16689,N_15845,N_16146);
nand U16690 (N_16690,N_16124,N_16055);
nor U16691 (N_16691,N_16210,N_16230);
and U16692 (N_16692,N_16216,N_15884);
nand U16693 (N_16693,N_16232,N_16000);
nor U16694 (N_16694,N_15657,N_16103);
and U16695 (N_16695,N_15760,N_15866);
and U16696 (N_16696,N_15845,N_16009);
and U16697 (N_16697,N_15968,N_15956);
or U16698 (N_16698,N_15977,N_15922);
xnor U16699 (N_16699,N_16233,N_15958);
or U16700 (N_16700,N_16221,N_15914);
nor U16701 (N_16701,N_15866,N_16072);
nand U16702 (N_16702,N_15733,N_15726);
or U16703 (N_16703,N_15658,N_15949);
and U16704 (N_16704,N_15981,N_16187);
or U16705 (N_16705,N_15625,N_15626);
or U16706 (N_16706,N_15872,N_15941);
or U16707 (N_16707,N_15868,N_15796);
and U16708 (N_16708,N_16004,N_15780);
xnor U16709 (N_16709,N_16167,N_16157);
nand U16710 (N_16710,N_16151,N_15853);
or U16711 (N_16711,N_15864,N_16241);
nand U16712 (N_16712,N_15713,N_15712);
or U16713 (N_16713,N_16198,N_16062);
or U16714 (N_16714,N_15732,N_15710);
and U16715 (N_16715,N_15957,N_15911);
and U16716 (N_16716,N_15884,N_15950);
xor U16717 (N_16717,N_16208,N_15857);
and U16718 (N_16718,N_16071,N_15769);
xnor U16719 (N_16719,N_15864,N_16105);
or U16720 (N_16720,N_15743,N_16118);
xor U16721 (N_16721,N_15989,N_16226);
xor U16722 (N_16722,N_16007,N_16240);
and U16723 (N_16723,N_16099,N_15707);
xnor U16724 (N_16724,N_15964,N_15690);
nor U16725 (N_16725,N_16004,N_16077);
or U16726 (N_16726,N_16089,N_15707);
nor U16727 (N_16727,N_15733,N_15811);
nor U16728 (N_16728,N_15888,N_15659);
or U16729 (N_16729,N_15874,N_16197);
nand U16730 (N_16730,N_16040,N_15830);
and U16731 (N_16731,N_15942,N_15871);
nor U16732 (N_16732,N_15726,N_16027);
or U16733 (N_16733,N_16033,N_16046);
or U16734 (N_16734,N_15960,N_15831);
nand U16735 (N_16735,N_15854,N_15785);
nand U16736 (N_16736,N_16103,N_15776);
nor U16737 (N_16737,N_16078,N_15801);
nor U16738 (N_16738,N_15703,N_15820);
nand U16739 (N_16739,N_15820,N_15738);
nor U16740 (N_16740,N_15788,N_15697);
nor U16741 (N_16741,N_16198,N_16095);
nor U16742 (N_16742,N_16103,N_15956);
xnor U16743 (N_16743,N_15816,N_16165);
or U16744 (N_16744,N_16001,N_15987);
or U16745 (N_16745,N_16222,N_16128);
nor U16746 (N_16746,N_15814,N_15707);
nor U16747 (N_16747,N_15992,N_15944);
or U16748 (N_16748,N_16150,N_15975);
and U16749 (N_16749,N_16083,N_15989);
and U16750 (N_16750,N_15641,N_16184);
nor U16751 (N_16751,N_15740,N_15723);
and U16752 (N_16752,N_16224,N_16129);
xor U16753 (N_16753,N_16090,N_15817);
nor U16754 (N_16754,N_15666,N_15708);
nor U16755 (N_16755,N_15763,N_16148);
or U16756 (N_16756,N_16186,N_15998);
nor U16757 (N_16757,N_15756,N_15702);
or U16758 (N_16758,N_16184,N_15842);
or U16759 (N_16759,N_16211,N_15634);
and U16760 (N_16760,N_16156,N_15678);
or U16761 (N_16761,N_16197,N_16228);
and U16762 (N_16762,N_15912,N_15678);
or U16763 (N_16763,N_16125,N_15907);
xnor U16764 (N_16764,N_15909,N_15731);
nand U16765 (N_16765,N_15854,N_16147);
and U16766 (N_16766,N_15659,N_15767);
or U16767 (N_16767,N_16149,N_15708);
nor U16768 (N_16768,N_16018,N_15645);
and U16769 (N_16769,N_16088,N_15743);
nand U16770 (N_16770,N_15894,N_16062);
or U16771 (N_16771,N_16118,N_15712);
or U16772 (N_16772,N_16023,N_15853);
or U16773 (N_16773,N_15933,N_15910);
xor U16774 (N_16774,N_15718,N_15961);
or U16775 (N_16775,N_15726,N_15988);
and U16776 (N_16776,N_15646,N_16152);
nand U16777 (N_16777,N_15820,N_15968);
xnor U16778 (N_16778,N_15973,N_15967);
or U16779 (N_16779,N_15952,N_15794);
nor U16780 (N_16780,N_16226,N_15802);
nor U16781 (N_16781,N_15931,N_16197);
nor U16782 (N_16782,N_15895,N_16174);
nand U16783 (N_16783,N_15971,N_15800);
nand U16784 (N_16784,N_16244,N_15878);
or U16785 (N_16785,N_16130,N_15682);
nor U16786 (N_16786,N_16243,N_16241);
xnor U16787 (N_16787,N_15844,N_15628);
nand U16788 (N_16788,N_15767,N_15816);
nand U16789 (N_16789,N_15773,N_15995);
or U16790 (N_16790,N_16081,N_15696);
nand U16791 (N_16791,N_16235,N_15703);
or U16792 (N_16792,N_15880,N_15858);
nor U16793 (N_16793,N_16063,N_16213);
nand U16794 (N_16794,N_15806,N_15761);
or U16795 (N_16795,N_15868,N_15640);
or U16796 (N_16796,N_15870,N_15863);
nor U16797 (N_16797,N_15968,N_15851);
nor U16798 (N_16798,N_16007,N_16058);
or U16799 (N_16799,N_16193,N_15835);
nand U16800 (N_16800,N_15968,N_16019);
and U16801 (N_16801,N_15945,N_15646);
nor U16802 (N_16802,N_15647,N_16150);
nand U16803 (N_16803,N_15643,N_15972);
nand U16804 (N_16804,N_15744,N_15985);
nor U16805 (N_16805,N_15893,N_16154);
or U16806 (N_16806,N_16135,N_15685);
nor U16807 (N_16807,N_15752,N_16112);
or U16808 (N_16808,N_15753,N_15693);
nand U16809 (N_16809,N_15690,N_16097);
nor U16810 (N_16810,N_15957,N_15759);
or U16811 (N_16811,N_16232,N_15688);
or U16812 (N_16812,N_15909,N_16193);
nand U16813 (N_16813,N_15852,N_16198);
nor U16814 (N_16814,N_16062,N_16022);
xnor U16815 (N_16815,N_15903,N_15870);
and U16816 (N_16816,N_15690,N_16042);
xnor U16817 (N_16817,N_15698,N_15750);
nand U16818 (N_16818,N_15815,N_16165);
and U16819 (N_16819,N_16007,N_15816);
and U16820 (N_16820,N_15798,N_16014);
and U16821 (N_16821,N_15660,N_15994);
and U16822 (N_16822,N_16138,N_15839);
and U16823 (N_16823,N_15798,N_16073);
nand U16824 (N_16824,N_15682,N_15678);
xor U16825 (N_16825,N_15705,N_15963);
or U16826 (N_16826,N_16151,N_15799);
or U16827 (N_16827,N_16169,N_15939);
and U16828 (N_16828,N_16027,N_15671);
or U16829 (N_16829,N_15847,N_15962);
nor U16830 (N_16830,N_15910,N_15756);
or U16831 (N_16831,N_16124,N_16160);
nor U16832 (N_16832,N_16076,N_15749);
and U16833 (N_16833,N_16206,N_16179);
or U16834 (N_16834,N_15800,N_15765);
or U16835 (N_16835,N_15895,N_15938);
or U16836 (N_16836,N_15999,N_15863);
nand U16837 (N_16837,N_15873,N_16217);
nand U16838 (N_16838,N_16112,N_16161);
and U16839 (N_16839,N_16038,N_15632);
nor U16840 (N_16840,N_15814,N_16213);
and U16841 (N_16841,N_15629,N_15685);
nand U16842 (N_16842,N_15756,N_15684);
or U16843 (N_16843,N_15693,N_16080);
xor U16844 (N_16844,N_15834,N_15792);
and U16845 (N_16845,N_15942,N_15783);
xor U16846 (N_16846,N_15808,N_15691);
nor U16847 (N_16847,N_15691,N_15662);
nor U16848 (N_16848,N_15951,N_15714);
xnor U16849 (N_16849,N_15858,N_15841);
nor U16850 (N_16850,N_15932,N_15897);
and U16851 (N_16851,N_16247,N_16105);
nand U16852 (N_16852,N_15861,N_15828);
and U16853 (N_16853,N_16126,N_15825);
or U16854 (N_16854,N_16087,N_15930);
xnor U16855 (N_16855,N_15821,N_15996);
and U16856 (N_16856,N_15835,N_16202);
or U16857 (N_16857,N_15746,N_16191);
nand U16858 (N_16858,N_15918,N_15670);
nor U16859 (N_16859,N_15981,N_16012);
or U16860 (N_16860,N_16082,N_15934);
nand U16861 (N_16861,N_15937,N_15730);
nor U16862 (N_16862,N_15853,N_15988);
nor U16863 (N_16863,N_16200,N_16096);
nor U16864 (N_16864,N_15848,N_16123);
nand U16865 (N_16865,N_15659,N_15690);
or U16866 (N_16866,N_16011,N_16171);
nor U16867 (N_16867,N_16198,N_16223);
nor U16868 (N_16868,N_15681,N_16233);
and U16869 (N_16869,N_16039,N_15657);
nand U16870 (N_16870,N_15794,N_15706);
and U16871 (N_16871,N_16185,N_15822);
or U16872 (N_16872,N_16126,N_16233);
nand U16873 (N_16873,N_15721,N_15679);
or U16874 (N_16874,N_16111,N_15885);
and U16875 (N_16875,N_16612,N_16474);
nand U16876 (N_16876,N_16476,N_16757);
or U16877 (N_16877,N_16815,N_16847);
nor U16878 (N_16878,N_16710,N_16342);
or U16879 (N_16879,N_16574,N_16546);
or U16880 (N_16880,N_16775,N_16427);
nor U16881 (N_16881,N_16550,N_16782);
or U16882 (N_16882,N_16841,N_16631);
nor U16883 (N_16883,N_16842,N_16452);
nand U16884 (N_16884,N_16515,N_16378);
or U16885 (N_16885,N_16516,N_16251);
nor U16886 (N_16886,N_16656,N_16596);
nand U16887 (N_16887,N_16716,N_16362);
nand U16888 (N_16888,N_16393,N_16691);
and U16889 (N_16889,N_16412,N_16661);
and U16890 (N_16890,N_16492,N_16318);
nand U16891 (N_16891,N_16717,N_16762);
nor U16892 (N_16892,N_16824,N_16781);
and U16893 (N_16893,N_16754,N_16403);
nand U16894 (N_16894,N_16576,N_16486);
and U16895 (N_16895,N_16314,N_16750);
xor U16896 (N_16896,N_16537,N_16281);
xor U16897 (N_16897,N_16471,N_16798);
nor U16898 (N_16898,N_16709,N_16786);
and U16899 (N_16899,N_16418,N_16852);
and U16900 (N_16900,N_16681,N_16644);
or U16901 (N_16901,N_16529,N_16316);
and U16902 (N_16902,N_16862,N_16769);
nand U16903 (N_16903,N_16706,N_16466);
nand U16904 (N_16904,N_16745,N_16264);
nand U16905 (N_16905,N_16291,N_16547);
and U16906 (N_16906,N_16791,N_16505);
xnor U16907 (N_16907,N_16873,N_16273);
nand U16908 (N_16908,N_16366,N_16541);
or U16909 (N_16909,N_16563,N_16851);
or U16910 (N_16910,N_16329,N_16472);
and U16911 (N_16911,N_16677,N_16693);
nor U16912 (N_16912,N_16272,N_16692);
nand U16913 (N_16913,N_16475,N_16712);
nand U16914 (N_16914,N_16614,N_16768);
or U16915 (N_16915,N_16835,N_16483);
and U16916 (N_16916,N_16761,N_16860);
nand U16917 (N_16917,N_16334,N_16501);
nor U16918 (N_16918,N_16578,N_16313);
nor U16919 (N_16919,N_16404,N_16635);
nand U16920 (N_16920,N_16360,N_16784);
nor U16921 (N_16921,N_16751,N_16361);
nor U16922 (N_16922,N_16737,N_16871);
and U16923 (N_16923,N_16494,N_16863);
or U16924 (N_16924,N_16726,N_16715);
or U16925 (N_16925,N_16419,N_16694);
and U16926 (N_16926,N_16363,N_16479);
nand U16927 (N_16927,N_16305,N_16292);
nor U16928 (N_16928,N_16290,N_16430);
xor U16929 (N_16929,N_16338,N_16662);
and U16930 (N_16930,N_16487,N_16640);
and U16931 (N_16931,N_16810,N_16438);
and U16932 (N_16932,N_16280,N_16489);
and U16933 (N_16933,N_16506,N_16748);
nand U16934 (N_16934,N_16323,N_16428);
nand U16935 (N_16935,N_16671,N_16389);
and U16936 (N_16936,N_16268,N_16702);
or U16937 (N_16937,N_16713,N_16434);
and U16938 (N_16938,N_16705,N_16857);
and U16939 (N_16939,N_16295,N_16255);
and U16940 (N_16940,N_16566,N_16267);
or U16941 (N_16941,N_16499,N_16813);
and U16942 (N_16942,N_16374,N_16573);
and U16943 (N_16943,N_16834,N_16535);
or U16944 (N_16944,N_16773,N_16846);
and U16945 (N_16945,N_16869,N_16509);
nand U16946 (N_16946,N_16561,N_16669);
and U16947 (N_16947,N_16420,N_16667);
or U16948 (N_16948,N_16413,N_16649);
and U16949 (N_16949,N_16260,N_16792);
nand U16950 (N_16950,N_16534,N_16375);
nor U16951 (N_16951,N_16437,N_16594);
and U16952 (N_16952,N_16687,N_16504);
nor U16953 (N_16953,N_16304,N_16302);
nor U16954 (N_16954,N_16779,N_16368);
or U16955 (N_16955,N_16819,N_16733);
xnor U16956 (N_16956,N_16743,N_16530);
and U16957 (N_16957,N_16785,N_16340);
or U16958 (N_16958,N_16580,N_16511);
nand U16959 (N_16959,N_16488,N_16480);
nor U16960 (N_16960,N_16558,N_16611);
nand U16961 (N_16961,N_16337,N_16325);
nor U16962 (N_16962,N_16676,N_16645);
and U16963 (N_16963,N_16440,N_16777);
nor U16964 (N_16964,N_16630,N_16606);
xor U16965 (N_16965,N_16592,N_16829);
nand U16966 (N_16966,N_16348,N_16600);
nor U16967 (N_16967,N_16738,N_16559);
nand U16968 (N_16968,N_16840,N_16758);
nand U16969 (N_16969,N_16582,N_16523);
and U16970 (N_16970,N_16454,N_16357);
nor U16971 (N_16971,N_16849,N_16394);
or U16972 (N_16972,N_16807,N_16827);
and U16973 (N_16973,N_16446,N_16690);
and U16974 (N_16974,N_16411,N_16753);
nand U16975 (N_16975,N_16482,N_16727);
or U16976 (N_16976,N_16823,N_16657);
and U16977 (N_16977,N_16684,N_16557);
or U16978 (N_16978,N_16700,N_16520);
and U16979 (N_16979,N_16821,N_16364);
and U16980 (N_16980,N_16533,N_16283);
and U16981 (N_16981,N_16457,N_16682);
nor U16982 (N_16982,N_16759,N_16579);
nor U16983 (N_16983,N_16435,N_16310);
or U16984 (N_16984,N_16774,N_16639);
nor U16985 (N_16985,N_16828,N_16674);
and U16986 (N_16986,N_16512,N_16287);
and U16987 (N_16987,N_16556,N_16730);
or U16988 (N_16988,N_16593,N_16736);
nor U16989 (N_16989,N_16409,N_16262);
or U16990 (N_16990,N_16335,N_16376);
xnor U16991 (N_16991,N_16806,N_16542);
or U16992 (N_16992,N_16392,N_16383);
nand U16993 (N_16993,N_16500,N_16618);
and U16994 (N_16994,N_16652,N_16586);
nand U16995 (N_16995,N_16755,N_16455);
nand U16996 (N_16996,N_16861,N_16818);
and U16997 (N_16997,N_16814,N_16633);
nor U16998 (N_16998,N_16493,N_16636);
nand U16999 (N_16999,N_16524,N_16299);
or U17000 (N_17000,N_16298,N_16679);
nand U17001 (N_17001,N_16385,N_16655);
xor U17002 (N_17002,N_16551,N_16503);
or U17003 (N_17003,N_16598,N_16648);
or U17004 (N_17004,N_16327,N_16695);
or U17005 (N_17005,N_16321,N_16417);
or U17006 (N_17006,N_16589,N_16303);
and U17007 (N_17007,N_16306,N_16402);
and U17008 (N_17008,N_16372,N_16742);
or U17009 (N_17009,N_16845,N_16508);
and U17010 (N_17010,N_16653,N_16444);
or U17011 (N_17011,N_16469,N_16347);
and U17012 (N_17012,N_16560,N_16549);
xnor U17013 (N_17013,N_16432,N_16673);
or U17014 (N_17014,N_16270,N_16461);
and U17015 (N_17015,N_16450,N_16590);
and U17016 (N_17016,N_16628,N_16658);
nand U17017 (N_17017,N_16353,N_16805);
and U17018 (N_17018,N_16689,N_16458);
and U17019 (N_17019,N_16767,N_16554);
and U17020 (N_17020,N_16351,N_16591);
or U17021 (N_17021,N_16540,N_16485);
and U17022 (N_17022,N_16790,N_16837);
and U17023 (N_17023,N_16367,N_16783);
xor U17024 (N_17024,N_16266,N_16756);
or U17025 (N_17025,N_16296,N_16464);
or U17026 (N_17026,N_16544,N_16607);
or U17027 (N_17027,N_16619,N_16473);
nor U17028 (N_17028,N_16780,N_16269);
and U17029 (N_17029,N_16634,N_16445);
nand U17030 (N_17030,N_16620,N_16514);
nand U17031 (N_17031,N_16701,N_16562);
nand U17032 (N_17032,N_16626,N_16646);
nor U17033 (N_17033,N_16804,N_16519);
or U17034 (N_17034,N_16604,N_16627);
nand U17035 (N_17035,N_16453,N_16406);
nand U17036 (N_17036,N_16465,N_16746);
or U17037 (N_17037,N_16250,N_16369);
xnor U17038 (N_17038,N_16431,N_16355);
nor U17039 (N_17039,N_16498,N_16872);
xnor U17040 (N_17040,N_16564,N_16567);
or U17041 (N_17041,N_16808,N_16311);
nor U17042 (N_17042,N_16258,N_16495);
nor U17043 (N_17043,N_16345,N_16405);
nand U17044 (N_17044,N_16532,N_16809);
or U17045 (N_17045,N_16300,N_16396);
nor U17046 (N_17046,N_16731,N_16531);
and U17047 (N_17047,N_16795,N_16497);
nor U17048 (N_17048,N_16772,N_16421);
nor U17049 (N_17049,N_16387,N_16714);
and U17050 (N_17050,N_16525,N_16339);
nand U17051 (N_17051,N_16443,N_16796);
nand U17052 (N_17052,N_16859,N_16831);
nand U17053 (N_17053,N_16722,N_16449);
or U17054 (N_17054,N_16408,N_16324);
nor U17055 (N_17055,N_16518,N_16349);
xnor U17056 (N_17056,N_16552,N_16553);
nand U17057 (N_17057,N_16401,N_16642);
nand U17058 (N_17058,N_16484,N_16253);
and U17059 (N_17059,N_16800,N_16838);
and U17060 (N_17060,N_16297,N_16568);
nand U17061 (N_17061,N_16858,N_16616);
nand U17062 (N_17062,N_16641,N_16548);
nand U17063 (N_17063,N_16665,N_16584);
nand U17064 (N_17064,N_16670,N_16666);
and U17065 (N_17065,N_16447,N_16650);
nand U17066 (N_17066,N_16856,N_16343);
nor U17067 (N_17067,N_16624,N_16254);
and U17068 (N_17068,N_16771,N_16336);
nand U17069 (N_17069,N_16341,N_16416);
and U17070 (N_17070,N_16587,N_16734);
nand U17071 (N_17071,N_16707,N_16536);
and U17072 (N_17072,N_16812,N_16422);
or U17073 (N_17073,N_16799,N_16629);
nand U17074 (N_17074,N_16732,N_16312);
nor U17075 (N_17075,N_16718,N_16721);
nor U17076 (N_17076,N_16704,N_16259);
nor U17077 (N_17077,N_16720,N_16678);
nor U17078 (N_17078,N_16870,N_16424);
nand U17079 (N_17079,N_16462,N_16326);
nand U17080 (N_17080,N_16328,N_16728);
or U17081 (N_17081,N_16448,N_16333);
nor U17082 (N_17082,N_16848,N_16803);
and U17083 (N_17083,N_16659,N_16853);
nor U17084 (N_17084,N_16315,N_16330);
nand U17085 (N_17085,N_16688,N_16766);
and U17086 (N_17086,N_16617,N_16289);
and U17087 (N_17087,N_16816,N_16460);
or U17088 (N_17088,N_16577,N_16850);
nor U17089 (N_17089,N_16293,N_16256);
and U17090 (N_17090,N_16836,N_16844);
xor U17091 (N_17091,N_16346,N_16344);
nand U17092 (N_17092,N_16274,N_16571);
or U17093 (N_17093,N_16735,N_16384);
or U17094 (N_17094,N_16703,N_16708);
and U17095 (N_17095,N_16654,N_16764);
nand U17096 (N_17096,N_16276,N_16252);
or U17097 (N_17097,N_16277,N_16386);
nor U17098 (N_17098,N_16356,N_16686);
and U17099 (N_17099,N_16866,N_16569);
nand U17100 (N_17100,N_16407,N_16522);
nor U17101 (N_17101,N_16599,N_16468);
nor U17102 (N_17102,N_16825,N_16663);
nor U17103 (N_17103,N_16414,N_16371);
nor U17104 (N_17104,N_16660,N_16601);
and U17105 (N_17105,N_16725,N_16388);
xnor U17106 (N_17106,N_16789,N_16770);
or U17107 (N_17107,N_16605,N_16855);
xor U17108 (N_17108,N_16491,N_16284);
xor U17109 (N_17109,N_16583,N_16822);
nand U17110 (N_17110,N_16271,N_16615);
and U17111 (N_17111,N_16826,N_16352);
or U17112 (N_17112,N_16729,N_16502);
nand U17113 (N_17113,N_16470,N_16651);
nand U17114 (N_17114,N_16477,N_16257);
or U17115 (N_17115,N_16797,N_16747);
or U17116 (N_17116,N_16623,N_16358);
nand U17117 (N_17117,N_16697,N_16545);
and U17118 (N_17118,N_16680,N_16320);
nor U17119 (N_17119,N_16811,N_16839);
or U17120 (N_17120,N_16638,N_16397);
nor U17121 (N_17121,N_16380,N_16467);
nand U17122 (N_17122,N_16539,N_16613);
or U17123 (N_17123,N_16581,N_16575);
and U17124 (N_17124,N_16282,N_16776);
nand U17125 (N_17125,N_16609,N_16740);
nor U17126 (N_17126,N_16830,N_16278);
nand U17127 (N_17127,N_16672,N_16426);
or U17128 (N_17128,N_16572,N_16741);
or U17129 (N_17129,N_16429,N_16749);
and U17130 (N_17130,N_16664,N_16399);
and U17131 (N_17131,N_16622,N_16867);
nor U17132 (N_17132,N_16864,N_16865);
nor U17133 (N_17133,N_16513,N_16719);
nand U17134 (N_17134,N_16365,N_16595);
and U17135 (N_17135,N_16279,N_16543);
nand U17136 (N_17136,N_16456,N_16832);
nand U17137 (N_17137,N_16793,N_16332);
nor U17138 (N_17138,N_16379,N_16763);
xnor U17139 (N_17139,N_16752,N_16265);
and U17140 (N_17140,N_16527,N_16787);
nand U17141 (N_17141,N_16382,N_16565);
nand U17142 (N_17142,N_16410,N_16538);
nand U17143 (N_17143,N_16490,N_16621);
nand U17144 (N_17144,N_16854,N_16442);
and U17145 (N_17145,N_16391,N_16436);
or U17146 (N_17146,N_16370,N_16698);
nor U17147 (N_17147,N_16381,N_16390);
or U17148 (N_17148,N_16322,N_16647);
and U17149 (N_17149,N_16843,N_16668);
or U17150 (N_17150,N_16377,N_16597);
nor U17151 (N_17151,N_16395,N_16788);
xnor U17152 (N_17152,N_16585,N_16496);
and U17153 (N_17153,N_16354,N_16625);
nor U17154 (N_17154,N_16570,N_16309);
nand U17155 (N_17155,N_16603,N_16685);
and U17156 (N_17156,N_16459,N_16528);
xnor U17157 (N_17157,N_16433,N_16555);
or U17158 (N_17158,N_16261,N_16331);
xnor U17159 (N_17159,N_16526,N_16373);
and U17160 (N_17160,N_16425,N_16833);
or U17161 (N_17161,N_16683,N_16874);
nor U17162 (N_17162,N_16675,N_16820);
or U17163 (N_17163,N_16602,N_16463);
nand U17164 (N_17164,N_16643,N_16760);
and U17165 (N_17165,N_16286,N_16507);
nand U17166 (N_17166,N_16317,N_16739);
and U17167 (N_17167,N_16794,N_16632);
xor U17168 (N_17168,N_16801,N_16307);
nor U17169 (N_17169,N_16588,N_16521);
nand U17170 (N_17170,N_16637,N_16608);
xor U17171 (N_17171,N_16359,N_16294);
or U17172 (N_17172,N_16400,N_16610);
and U17173 (N_17173,N_16439,N_16285);
nand U17174 (N_17174,N_16765,N_16451);
or U17175 (N_17175,N_16478,N_16288);
or U17176 (N_17176,N_16724,N_16263);
nand U17177 (N_17177,N_16510,N_16481);
and U17178 (N_17178,N_16723,N_16517);
nand U17179 (N_17179,N_16301,N_16817);
or U17180 (N_17180,N_16802,N_16699);
nand U17181 (N_17181,N_16868,N_16319);
nor U17182 (N_17182,N_16423,N_16744);
or U17183 (N_17183,N_16275,N_16415);
nand U17184 (N_17184,N_16778,N_16711);
xnor U17185 (N_17185,N_16350,N_16308);
and U17186 (N_17186,N_16398,N_16441);
nor U17187 (N_17187,N_16696,N_16373);
or U17188 (N_17188,N_16564,N_16404);
and U17189 (N_17189,N_16477,N_16321);
nor U17190 (N_17190,N_16867,N_16698);
nor U17191 (N_17191,N_16317,N_16320);
nor U17192 (N_17192,N_16585,N_16760);
and U17193 (N_17193,N_16486,N_16619);
and U17194 (N_17194,N_16704,N_16535);
or U17195 (N_17195,N_16543,N_16323);
xor U17196 (N_17196,N_16688,N_16305);
xnor U17197 (N_17197,N_16350,N_16271);
nor U17198 (N_17198,N_16266,N_16832);
and U17199 (N_17199,N_16386,N_16646);
and U17200 (N_17200,N_16332,N_16448);
and U17201 (N_17201,N_16752,N_16431);
nor U17202 (N_17202,N_16605,N_16603);
and U17203 (N_17203,N_16779,N_16491);
and U17204 (N_17204,N_16816,N_16423);
nor U17205 (N_17205,N_16652,N_16467);
and U17206 (N_17206,N_16846,N_16795);
nand U17207 (N_17207,N_16275,N_16250);
nor U17208 (N_17208,N_16729,N_16671);
nand U17209 (N_17209,N_16804,N_16526);
xnor U17210 (N_17210,N_16632,N_16843);
or U17211 (N_17211,N_16738,N_16560);
and U17212 (N_17212,N_16613,N_16445);
xnor U17213 (N_17213,N_16610,N_16497);
or U17214 (N_17214,N_16334,N_16716);
and U17215 (N_17215,N_16468,N_16273);
nand U17216 (N_17216,N_16276,N_16606);
nor U17217 (N_17217,N_16391,N_16383);
nor U17218 (N_17218,N_16584,N_16326);
or U17219 (N_17219,N_16349,N_16702);
nor U17220 (N_17220,N_16323,N_16358);
or U17221 (N_17221,N_16732,N_16420);
or U17222 (N_17222,N_16786,N_16404);
and U17223 (N_17223,N_16552,N_16277);
or U17224 (N_17224,N_16745,N_16610);
and U17225 (N_17225,N_16462,N_16690);
nand U17226 (N_17226,N_16602,N_16633);
nor U17227 (N_17227,N_16581,N_16700);
xor U17228 (N_17228,N_16790,N_16330);
nor U17229 (N_17229,N_16735,N_16323);
nor U17230 (N_17230,N_16266,N_16774);
and U17231 (N_17231,N_16505,N_16621);
and U17232 (N_17232,N_16387,N_16251);
or U17233 (N_17233,N_16824,N_16754);
nand U17234 (N_17234,N_16625,N_16837);
xor U17235 (N_17235,N_16677,N_16337);
nor U17236 (N_17236,N_16333,N_16308);
and U17237 (N_17237,N_16671,N_16734);
or U17238 (N_17238,N_16680,N_16867);
nand U17239 (N_17239,N_16733,N_16479);
xor U17240 (N_17240,N_16519,N_16787);
nand U17241 (N_17241,N_16765,N_16861);
and U17242 (N_17242,N_16555,N_16639);
xnor U17243 (N_17243,N_16654,N_16784);
xor U17244 (N_17244,N_16635,N_16324);
nor U17245 (N_17245,N_16835,N_16457);
and U17246 (N_17246,N_16290,N_16602);
and U17247 (N_17247,N_16397,N_16598);
or U17248 (N_17248,N_16382,N_16855);
nor U17249 (N_17249,N_16415,N_16620);
and U17250 (N_17250,N_16489,N_16705);
or U17251 (N_17251,N_16798,N_16543);
nor U17252 (N_17252,N_16817,N_16779);
or U17253 (N_17253,N_16666,N_16252);
nor U17254 (N_17254,N_16555,N_16478);
xor U17255 (N_17255,N_16487,N_16309);
nor U17256 (N_17256,N_16518,N_16698);
nand U17257 (N_17257,N_16810,N_16502);
nor U17258 (N_17258,N_16871,N_16293);
xnor U17259 (N_17259,N_16569,N_16562);
or U17260 (N_17260,N_16339,N_16527);
or U17261 (N_17261,N_16865,N_16600);
and U17262 (N_17262,N_16837,N_16600);
or U17263 (N_17263,N_16285,N_16263);
nand U17264 (N_17264,N_16625,N_16559);
and U17265 (N_17265,N_16372,N_16276);
nand U17266 (N_17266,N_16260,N_16327);
nor U17267 (N_17267,N_16462,N_16471);
and U17268 (N_17268,N_16444,N_16362);
nor U17269 (N_17269,N_16383,N_16364);
xor U17270 (N_17270,N_16432,N_16289);
and U17271 (N_17271,N_16362,N_16859);
nor U17272 (N_17272,N_16425,N_16387);
nor U17273 (N_17273,N_16527,N_16803);
and U17274 (N_17274,N_16313,N_16446);
nor U17275 (N_17275,N_16468,N_16485);
nand U17276 (N_17276,N_16562,N_16365);
nor U17277 (N_17277,N_16814,N_16332);
and U17278 (N_17278,N_16668,N_16541);
and U17279 (N_17279,N_16381,N_16683);
nor U17280 (N_17280,N_16781,N_16682);
nor U17281 (N_17281,N_16288,N_16518);
or U17282 (N_17282,N_16640,N_16326);
nor U17283 (N_17283,N_16332,N_16625);
or U17284 (N_17284,N_16844,N_16568);
or U17285 (N_17285,N_16681,N_16709);
xnor U17286 (N_17286,N_16368,N_16549);
nor U17287 (N_17287,N_16424,N_16446);
or U17288 (N_17288,N_16861,N_16522);
or U17289 (N_17289,N_16370,N_16631);
xor U17290 (N_17290,N_16351,N_16530);
nor U17291 (N_17291,N_16501,N_16784);
nand U17292 (N_17292,N_16716,N_16538);
and U17293 (N_17293,N_16819,N_16648);
and U17294 (N_17294,N_16729,N_16482);
nand U17295 (N_17295,N_16310,N_16252);
xor U17296 (N_17296,N_16374,N_16819);
nand U17297 (N_17297,N_16734,N_16251);
or U17298 (N_17298,N_16615,N_16667);
or U17299 (N_17299,N_16510,N_16528);
nor U17300 (N_17300,N_16789,N_16587);
nor U17301 (N_17301,N_16351,N_16440);
nand U17302 (N_17302,N_16786,N_16851);
xor U17303 (N_17303,N_16457,N_16757);
and U17304 (N_17304,N_16752,N_16733);
nand U17305 (N_17305,N_16655,N_16801);
or U17306 (N_17306,N_16660,N_16330);
nand U17307 (N_17307,N_16663,N_16399);
or U17308 (N_17308,N_16536,N_16813);
nor U17309 (N_17309,N_16572,N_16737);
xnor U17310 (N_17310,N_16391,N_16787);
nand U17311 (N_17311,N_16431,N_16701);
nor U17312 (N_17312,N_16326,N_16839);
nor U17313 (N_17313,N_16692,N_16420);
or U17314 (N_17314,N_16296,N_16620);
nand U17315 (N_17315,N_16617,N_16471);
nor U17316 (N_17316,N_16388,N_16362);
nor U17317 (N_17317,N_16624,N_16420);
or U17318 (N_17318,N_16675,N_16346);
or U17319 (N_17319,N_16292,N_16545);
or U17320 (N_17320,N_16630,N_16386);
nand U17321 (N_17321,N_16376,N_16587);
nand U17322 (N_17322,N_16825,N_16728);
or U17323 (N_17323,N_16280,N_16406);
xor U17324 (N_17324,N_16764,N_16294);
or U17325 (N_17325,N_16301,N_16262);
or U17326 (N_17326,N_16293,N_16554);
or U17327 (N_17327,N_16604,N_16862);
and U17328 (N_17328,N_16546,N_16759);
nand U17329 (N_17329,N_16365,N_16430);
or U17330 (N_17330,N_16305,N_16709);
nand U17331 (N_17331,N_16299,N_16641);
or U17332 (N_17332,N_16747,N_16422);
nand U17333 (N_17333,N_16562,N_16760);
xor U17334 (N_17334,N_16814,N_16376);
nand U17335 (N_17335,N_16805,N_16284);
or U17336 (N_17336,N_16620,N_16553);
nand U17337 (N_17337,N_16462,N_16597);
nor U17338 (N_17338,N_16867,N_16761);
nand U17339 (N_17339,N_16327,N_16496);
nor U17340 (N_17340,N_16703,N_16546);
nor U17341 (N_17341,N_16473,N_16594);
nand U17342 (N_17342,N_16308,N_16353);
nor U17343 (N_17343,N_16583,N_16813);
xor U17344 (N_17344,N_16479,N_16435);
or U17345 (N_17345,N_16684,N_16633);
and U17346 (N_17346,N_16572,N_16678);
or U17347 (N_17347,N_16752,N_16696);
and U17348 (N_17348,N_16293,N_16305);
nand U17349 (N_17349,N_16489,N_16546);
nor U17350 (N_17350,N_16815,N_16579);
and U17351 (N_17351,N_16445,N_16376);
or U17352 (N_17352,N_16549,N_16789);
nand U17353 (N_17353,N_16432,N_16657);
nand U17354 (N_17354,N_16375,N_16649);
nand U17355 (N_17355,N_16801,N_16493);
or U17356 (N_17356,N_16482,N_16300);
nand U17357 (N_17357,N_16518,N_16787);
or U17358 (N_17358,N_16785,N_16646);
or U17359 (N_17359,N_16829,N_16858);
nand U17360 (N_17360,N_16655,N_16645);
xor U17361 (N_17361,N_16557,N_16368);
or U17362 (N_17362,N_16603,N_16698);
and U17363 (N_17363,N_16540,N_16380);
and U17364 (N_17364,N_16683,N_16618);
nand U17365 (N_17365,N_16873,N_16443);
nor U17366 (N_17366,N_16869,N_16527);
nor U17367 (N_17367,N_16293,N_16641);
or U17368 (N_17368,N_16488,N_16540);
nor U17369 (N_17369,N_16559,N_16327);
and U17370 (N_17370,N_16340,N_16413);
and U17371 (N_17371,N_16382,N_16720);
xor U17372 (N_17372,N_16585,N_16394);
xor U17373 (N_17373,N_16530,N_16288);
or U17374 (N_17374,N_16741,N_16623);
or U17375 (N_17375,N_16843,N_16539);
or U17376 (N_17376,N_16624,N_16701);
nand U17377 (N_17377,N_16324,N_16631);
xor U17378 (N_17378,N_16273,N_16616);
nand U17379 (N_17379,N_16512,N_16829);
nor U17380 (N_17380,N_16853,N_16360);
or U17381 (N_17381,N_16754,N_16728);
nor U17382 (N_17382,N_16416,N_16666);
and U17383 (N_17383,N_16510,N_16411);
nor U17384 (N_17384,N_16845,N_16591);
or U17385 (N_17385,N_16398,N_16528);
nand U17386 (N_17386,N_16414,N_16837);
or U17387 (N_17387,N_16679,N_16698);
and U17388 (N_17388,N_16388,N_16438);
nand U17389 (N_17389,N_16740,N_16855);
nand U17390 (N_17390,N_16331,N_16602);
and U17391 (N_17391,N_16426,N_16754);
or U17392 (N_17392,N_16252,N_16565);
and U17393 (N_17393,N_16733,N_16549);
and U17394 (N_17394,N_16659,N_16584);
or U17395 (N_17395,N_16856,N_16655);
nand U17396 (N_17396,N_16490,N_16658);
and U17397 (N_17397,N_16778,N_16663);
nor U17398 (N_17398,N_16828,N_16520);
nand U17399 (N_17399,N_16366,N_16766);
xnor U17400 (N_17400,N_16441,N_16813);
nor U17401 (N_17401,N_16457,N_16319);
xor U17402 (N_17402,N_16790,N_16488);
xor U17403 (N_17403,N_16712,N_16703);
nand U17404 (N_17404,N_16359,N_16749);
nor U17405 (N_17405,N_16358,N_16516);
and U17406 (N_17406,N_16522,N_16718);
nor U17407 (N_17407,N_16444,N_16779);
or U17408 (N_17408,N_16265,N_16434);
nor U17409 (N_17409,N_16527,N_16480);
or U17410 (N_17410,N_16489,N_16265);
or U17411 (N_17411,N_16389,N_16817);
xor U17412 (N_17412,N_16628,N_16536);
and U17413 (N_17413,N_16256,N_16826);
nor U17414 (N_17414,N_16521,N_16375);
nand U17415 (N_17415,N_16252,N_16655);
and U17416 (N_17416,N_16727,N_16837);
and U17417 (N_17417,N_16543,N_16289);
nand U17418 (N_17418,N_16291,N_16259);
nand U17419 (N_17419,N_16562,N_16639);
nand U17420 (N_17420,N_16375,N_16343);
or U17421 (N_17421,N_16559,N_16372);
nor U17422 (N_17422,N_16347,N_16582);
or U17423 (N_17423,N_16382,N_16396);
or U17424 (N_17424,N_16513,N_16409);
nand U17425 (N_17425,N_16288,N_16874);
xnor U17426 (N_17426,N_16642,N_16680);
and U17427 (N_17427,N_16744,N_16543);
and U17428 (N_17428,N_16705,N_16429);
xor U17429 (N_17429,N_16349,N_16305);
nand U17430 (N_17430,N_16266,N_16614);
nor U17431 (N_17431,N_16733,N_16622);
nor U17432 (N_17432,N_16479,N_16617);
and U17433 (N_17433,N_16695,N_16861);
nand U17434 (N_17434,N_16732,N_16568);
or U17435 (N_17435,N_16511,N_16684);
or U17436 (N_17436,N_16613,N_16621);
nor U17437 (N_17437,N_16683,N_16502);
or U17438 (N_17438,N_16411,N_16492);
xor U17439 (N_17439,N_16755,N_16772);
and U17440 (N_17440,N_16603,N_16388);
nand U17441 (N_17441,N_16602,N_16533);
nand U17442 (N_17442,N_16451,N_16696);
nor U17443 (N_17443,N_16471,N_16775);
or U17444 (N_17444,N_16295,N_16829);
nor U17445 (N_17445,N_16561,N_16828);
xor U17446 (N_17446,N_16493,N_16788);
nand U17447 (N_17447,N_16582,N_16572);
nand U17448 (N_17448,N_16812,N_16758);
nand U17449 (N_17449,N_16253,N_16461);
xor U17450 (N_17450,N_16360,N_16859);
nand U17451 (N_17451,N_16590,N_16307);
or U17452 (N_17452,N_16791,N_16841);
or U17453 (N_17453,N_16395,N_16721);
and U17454 (N_17454,N_16680,N_16816);
and U17455 (N_17455,N_16291,N_16455);
xor U17456 (N_17456,N_16817,N_16371);
nor U17457 (N_17457,N_16587,N_16394);
nor U17458 (N_17458,N_16809,N_16332);
and U17459 (N_17459,N_16761,N_16557);
nand U17460 (N_17460,N_16832,N_16721);
and U17461 (N_17461,N_16433,N_16514);
and U17462 (N_17462,N_16256,N_16629);
nand U17463 (N_17463,N_16651,N_16461);
and U17464 (N_17464,N_16708,N_16281);
nand U17465 (N_17465,N_16546,N_16299);
or U17466 (N_17466,N_16346,N_16787);
nand U17467 (N_17467,N_16440,N_16361);
nor U17468 (N_17468,N_16728,N_16785);
nand U17469 (N_17469,N_16428,N_16426);
and U17470 (N_17470,N_16475,N_16337);
or U17471 (N_17471,N_16774,N_16475);
or U17472 (N_17472,N_16410,N_16643);
and U17473 (N_17473,N_16412,N_16530);
nand U17474 (N_17474,N_16639,N_16816);
or U17475 (N_17475,N_16483,N_16667);
nand U17476 (N_17476,N_16438,N_16401);
and U17477 (N_17477,N_16252,N_16720);
nor U17478 (N_17478,N_16533,N_16872);
nor U17479 (N_17479,N_16509,N_16366);
or U17480 (N_17480,N_16838,N_16429);
nor U17481 (N_17481,N_16810,N_16550);
nand U17482 (N_17482,N_16758,N_16532);
nand U17483 (N_17483,N_16413,N_16596);
and U17484 (N_17484,N_16353,N_16749);
nand U17485 (N_17485,N_16673,N_16439);
or U17486 (N_17486,N_16416,N_16678);
and U17487 (N_17487,N_16442,N_16568);
nand U17488 (N_17488,N_16633,N_16474);
and U17489 (N_17489,N_16288,N_16433);
nor U17490 (N_17490,N_16327,N_16572);
nand U17491 (N_17491,N_16869,N_16502);
nor U17492 (N_17492,N_16342,N_16547);
nor U17493 (N_17493,N_16378,N_16533);
nand U17494 (N_17494,N_16327,N_16289);
and U17495 (N_17495,N_16369,N_16667);
xor U17496 (N_17496,N_16794,N_16781);
nand U17497 (N_17497,N_16261,N_16484);
nand U17498 (N_17498,N_16375,N_16444);
or U17499 (N_17499,N_16400,N_16318);
or U17500 (N_17500,N_17406,N_17205);
nor U17501 (N_17501,N_17105,N_17222);
nand U17502 (N_17502,N_17334,N_17193);
and U17503 (N_17503,N_16989,N_17249);
nand U17504 (N_17504,N_17322,N_17375);
nor U17505 (N_17505,N_17066,N_17012);
nor U17506 (N_17506,N_17359,N_16954);
or U17507 (N_17507,N_17332,N_17153);
nor U17508 (N_17508,N_16957,N_17290);
xnor U17509 (N_17509,N_16917,N_17043);
nor U17510 (N_17510,N_16985,N_17433);
nor U17511 (N_17511,N_17420,N_17013);
xnor U17512 (N_17512,N_17469,N_17472);
nand U17513 (N_17513,N_16958,N_16993);
and U17514 (N_17514,N_17197,N_17301);
nand U17515 (N_17515,N_17095,N_17115);
or U17516 (N_17516,N_17045,N_16945);
nor U17517 (N_17517,N_17201,N_17461);
or U17518 (N_17518,N_16905,N_17267);
or U17519 (N_17519,N_16935,N_17340);
xor U17520 (N_17520,N_17055,N_17454);
nand U17521 (N_17521,N_17260,N_17304);
or U17522 (N_17522,N_17208,N_17402);
nor U17523 (N_17523,N_16894,N_17492);
nor U17524 (N_17524,N_16994,N_17282);
nand U17525 (N_17525,N_17067,N_17320);
nor U17526 (N_17526,N_17146,N_17302);
and U17527 (N_17527,N_16931,N_17457);
nand U17528 (N_17528,N_17215,N_17064);
nor U17529 (N_17529,N_16979,N_17382);
nand U17530 (N_17530,N_17463,N_16943);
nand U17531 (N_17531,N_17030,N_17243);
nand U17532 (N_17532,N_17148,N_17385);
or U17533 (N_17533,N_16984,N_17104);
and U17534 (N_17534,N_17180,N_17430);
nor U17535 (N_17535,N_17174,N_17210);
nand U17536 (N_17536,N_17296,N_17220);
nand U17537 (N_17537,N_16912,N_17379);
and U17538 (N_17538,N_17179,N_16995);
or U17539 (N_17539,N_16930,N_17116);
or U17540 (N_17540,N_16952,N_17170);
nand U17541 (N_17541,N_16987,N_17265);
or U17542 (N_17542,N_17086,N_16900);
nand U17543 (N_17543,N_17446,N_17311);
nor U17544 (N_17544,N_17156,N_17256);
nand U17545 (N_17545,N_17278,N_17005);
and U17546 (N_17546,N_16896,N_17008);
xor U17547 (N_17547,N_17400,N_17032);
nand U17548 (N_17548,N_17294,N_17052);
nand U17549 (N_17549,N_17368,N_17031);
nor U17550 (N_17550,N_17289,N_17303);
or U17551 (N_17551,N_16884,N_17337);
nand U17552 (N_17552,N_17245,N_17333);
or U17553 (N_17553,N_17074,N_16923);
or U17554 (N_17554,N_16882,N_16961);
nor U17555 (N_17555,N_17076,N_17452);
and U17556 (N_17556,N_17060,N_17422);
or U17557 (N_17557,N_17355,N_17440);
or U17558 (N_17558,N_16901,N_16950);
nor U17559 (N_17559,N_17135,N_17364);
or U17560 (N_17560,N_17324,N_17234);
nor U17561 (N_17561,N_16955,N_17435);
or U17562 (N_17562,N_17439,N_17152);
nand U17563 (N_17563,N_17130,N_17258);
xnor U17564 (N_17564,N_17285,N_16890);
nor U17565 (N_17565,N_16951,N_16953);
nand U17566 (N_17566,N_17183,N_16990);
xnor U17567 (N_17567,N_17128,N_17474);
and U17568 (N_17568,N_17218,N_17036);
nor U17569 (N_17569,N_17229,N_17438);
and U17570 (N_17570,N_17247,N_17058);
nor U17571 (N_17571,N_17407,N_17001);
nand U17572 (N_17572,N_17255,N_17122);
nor U17573 (N_17573,N_17214,N_16891);
or U17574 (N_17574,N_17161,N_16988);
nor U17575 (N_17575,N_17004,N_17150);
and U17576 (N_17576,N_17056,N_17139);
nand U17577 (N_17577,N_17022,N_17317);
nand U17578 (N_17578,N_16929,N_17313);
and U17579 (N_17579,N_17342,N_16926);
nand U17580 (N_17580,N_16965,N_17347);
xnor U17581 (N_17581,N_17073,N_17014);
or U17582 (N_17582,N_17119,N_17389);
nand U17583 (N_17583,N_17354,N_16910);
nand U17584 (N_17584,N_17266,N_16970);
nor U17585 (N_17585,N_17353,N_16933);
or U17586 (N_17586,N_17292,N_17112);
nor U17587 (N_17587,N_17419,N_17033);
nand U17588 (N_17588,N_17371,N_17336);
or U17589 (N_17589,N_17381,N_17274);
nand U17590 (N_17590,N_17018,N_17445);
or U17591 (N_17591,N_17000,N_17464);
or U17592 (N_17592,N_17221,N_17273);
nand U17593 (N_17593,N_17228,N_17498);
or U17594 (N_17594,N_17493,N_17037);
xor U17595 (N_17595,N_17137,N_17281);
nand U17596 (N_17596,N_17141,N_16940);
nand U17597 (N_17597,N_16977,N_16897);
nand U17598 (N_17598,N_16983,N_17028);
or U17599 (N_17599,N_17094,N_17190);
or U17600 (N_17600,N_16949,N_17168);
nor U17601 (N_17601,N_17203,N_17275);
and U17602 (N_17602,N_17189,N_16963);
xnor U17603 (N_17603,N_16932,N_17216);
and U17604 (N_17604,N_17209,N_17227);
and U17605 (N_17605,N_17329,N_17328);
or U17606 (N_17606,N_17306,N_17127);
nor U17607 (N_17607,N_17449,N_17065);
and U17608 (N_17608,N_16934,N_17416);
and U17609 (N_17609,N_17075,N_17102);
nor U17610 (N_17610,N_17039,N_17162);
or U17611 (N_17611,N_17478,N_17388);
or U17612 (N_17612,N_17432,N_17434);
xnor U17613 (N_17613,N_16925,N_17090);
nand U17614 (N_17614,N_17259,N_17191);
or U17615 (N_17615,N_17237,N_17113);
or U17616 (N_17616,N_16919,N_17300);
or U17617 (N_17617,N_16982,N_16974);
or U17618 (N_17618,N_17269,N_16876);
nor U17619 (N_17619,N_17479,N_17428);
xor U17620 (N_17620,N_17424,N_17133);
and U17621 (N_17621,N_17466,N_17029);
nand U17622 (N_17622,N_17473,N_17108);
nor U17623 (N_17623,N_17323,N_17142);
nor U17624 (N_17624,N_17326,N_17476);
or U17625 (N_17625,N_17475,N_17040);
xor U17626 (N_17626,N_16972,N_17341);
nor U17627 (N_17627,N_17070,N_17471);
xor U17628 (N_17628,N_17280,N_17054);
nand U17629 (N_17629,N_17253,N_17426);
nor U17630 (N_17630,N_17405,N_17182);
nand U17631 (N_17631,N_17360,N_17077);
nand U17632 (N_17632,N_17268,N_17305);
and U17633 (N_17633,N_17376,N_17468);
nand U17634 (N_17634,N_17423,N_16973);
and U17635 (N_17635,N_17129,N_17158);
nand U17636 (N_17636,N_17362,N_17240);
xor U17637 (N_17637,N_16886,N_17431);
nor U17638 (N_17638,N_17017,N_16903);
nor U17639 (N_17639,N_17194,N_17458);
and U17640 (N_17640,N_17436,N_17262);
nand U17641 (N_17641,N_16885,N_17042);
nor U17642 (N_17642,N_17176,N_16889);
nand U17643 (N_17643,N_17490,N_17465);
nand U17644 (N_17644,N_17188,N_17496);
and U17645 (N_17645,N_17025,N_16975);
nand U17646 (N_17646,N_17338,N_17034);
or U17647 (N_17647,N_17175,N_16893);
nor U17648 (N_17648,N_17134,N_17101);
or U17649 (N_17649,N_17069,N_17003);
or U17650 (N_17650,N_16967,N_17319);
nand U17651 (N_17651,N_17109,N_17386);
nand U17652 (N_17652,N_17261,N_17235);
nand U17653 (N_17653,N_17287,N_17299);
or U17654 (N_17654,N_17023,N_16927);
nand U17655 (N_17655,N_17225,N_17250);
and U17656 (N_17656,N_17011,N_17467);
and U17657 (N_17657,N_17114,N_17395);
nand U17658 (N_17658,N_17082,N_17448);
and U17659 (N_17659,N_17110,N_17339);
nor U17660 (N_17660,N_17233,N_16962);
or U17661 (N_17661,N_17357,N_17230);
nor U17662 (N_17662,N_17173,N_17450);
xnor U17663 (N_17663,N_16907,N_17213);
nand U17664 (N_17664,N_17038,N_16956);
nor U17665 (N_17665,N_17295,N_17316);
nor U17666 (N_17666,N_17041,N_17021);
xnor U17667 (N_17667,N_17126,N_17373);
or U17668 (N_17668,N_17482,N_17314);
nand U17669 (N_17669,N_16960,N_17470);
xnor U17670 (N_17670,N_17283,N_17051);
or U17671 (N_17671,N_17096,N_17124);
nor U17672 (N_17672,N_17160,N_17263);
nor U17673 (N_17673,N_17413,N_16942);
nand U17674 (N_17674,N_17047,N_16899);
nor U17675 (N_17675,N_17120,N_17186);
nor U17676 (N_17676,N_17231,N_16898);
or U17677 (N_17677,N_17459,N_17192);
nand U17678 (N_17678,N_17370,N_16906);
nor U17679 (N_17679,N_17421,N_17195);
nand U17680 (N_17680,N_16920,N_17318);
nand U17681 (N_17681,N_17200,N_17167);
xor U17682 (N_17682,N_17123,N_16980);
or U17683 (N_17683,N_16913,N_17393);
nor U17684 (N_17684,N_17427,N_17151);
or U17685 (N_17685,N_17044,N_16928);
or U17686 (N_17686,N_17121,N_17270);
nand U17687 (N_17687,N_17050,N_17199);
and U17688 (N_17688,N_17089,N_17027);
nand U17689 (N_17689,N_17335,N_16879);
nor U17690 (N_17690,N_17272,N_17140);
nand U17691 (N_17691,N_16880,N_17091);
or U17692 (N_17692,N_16978,N_17418);
and U17693 (N_17693,N_17369,N_17020);
and U17694 (N_17694,N_17083,N_17226);
or U17695 (N_17695,N_17125,N_17410);
nand U17696 (N_17696,N_17092,N_16887);
nor U17697 (N_17697,N_17138,N_17396);
nand U17698 (N_17698,N_17107,N_17223);
nor U17699 (N_17699,N_17079,N_17172);
or U17700 (N_17700,N_17164,N_17015);
or U17701 (N_17701,N_17085,N_17411);
nand U17702 (N_17702,N_16992,N_16991);
nor U17703 (N_17703,N_16914,N_17063);
and U17704 (N_17704,N_17048,N_17309);
and U17705 (N_17705,N_16986,N_17232);
or U17706 (N_17706,N_17163,N_17497);
nand U17707 (N_17707,N_17325,N_17293);
and U17708 (N_17708,N_17071,N_16911);
nand U17709 (N_17709,N_17387,N_17437);
nor U17710 (N_17710,N_17211,N_17248);
nand U17711 (N_17711,N_17351,N_17481);
nor U17712 (N_17712,N_17352,N_16968);
or U17713 (N_17713,N_16916,N_17307);
and U17714 (N_17714,N_17392,N_16939);
nor U17715 (N_17715,N_17157,N_17111);
xnor U17716 (N_17716,N_17310,N_17219);
nand U17717 (N_17717,N_16959,N_16996);
and U17718 (N_17718,N_17315,N_16908);
nand U17719 (N_17719,N_17046,N_17425);
or U17720 (N_17720,N_17429,N_17276);
or U17721 (N_17721,N_17477,N_17346);
or U17722 (N_17722,N_16999,N_17099);
and U17723 (N_17723,N_17378,N_17016);
and U17724 (N_17724,N_16915,N_17365);
nor U17725 (N_17725,N_17257,N_17344);
or U17726 (N_17726,N_17312,N_17297);
and U17727 (N_17727,N_17007,N_17026);
xor U17728 (N_17728,N_17495,N_17035);
and U17729 (N_17729,N_17131,N_17455);
nand U17730 (N_17730,N_16875,N_17072);
xnor U17731 (N_17731,N_17499,N_17377);
or U17732 (N_17732,N_17155,N_17059);
or U17733 (N_17733,N_16918,N_16878);
and U17734 (N_17734,N_17356,N_17217);
xnor U17735 (N_17735,N_17279,N_17483);
nand U17736 (N_17736,N_17291,N_17453);
and U17737 (N_17737,N_17308,N_16971);
nand U17738 (N_17738,N_17145,N_17383);
xnor U17739 (N_17739,N_17277,N_16944);
xor U17740 (N_17740,N_17100,N_17408);
and U17741 (N_17741,N_17238,N_17202);
and U17742 (N_17742,N_17103,N_17391);
and U17743 (N_17743,N_17489,N_17264);
nor U17744 (N_17744,N_17132,N_17321);
or U17745 (N_17745,N_16881,N_17204);
nand U17746 (N_17746,N_17441,N_16938);
and U17747 (N_17747,N_16969,N_17159);
xor U17748 (N_17748,N_17480,N_17397);
nand U17749 (N_17749,N_17185,N_16936);
xor U17750 (N_17750,N_17349,N_17398);
xnor U17751 (N_17751,N_17078,N_17363);
nor U17752 (N_17752,N_17358,N_16976);
nand U17753 (N_17753,N_17178,N_17187);
or U17754 (N_17754,N_17380,N_17184);
or U17755 (N_17755,N_17403,N_17198);
nand U17756 (N_17756,N_16966,N_17374);
or U17757 (N_17757,N_17331,N_16922);
and U17758 (N_17758,N_17062,N_17444);
nand U17759 (N_17759,N_17149,N_17118);
nand U17760 (N_17760,N_17081,N_17068);
or U17761 (N_17761,N_16909,N_17053);
nand U17762 (N_17762,N_17361,N_17241);
and U17763 (N_17763,N_16883,N_17447);
and U17764 (N_17764,N_17087,N_16904);
and U17765 (N_17765,N_17394,N_17491);
and U17766 (N_17766,N_16964,N_16895);
or U17767 (N_17767,N_17080,N_17414);
nor U17768 (N_17768,N_17417,N_17399);
nand U17769 (N_17769,N_17284,N_17485);
xnor U17770 (N_17770,N_17390,N_17098);
or U17771 (N_17771,N_17181,N_16937);
or U17772 (N_17772,N_17212,N_17244);
and U17773 (N_17773,N_17484,N_17147);
xnor U17774 (N_17774,N_17144,N_17487);
nand U17775 (N_17775,N_17196,N_17288);
or U17776 (N_17776,N_17494,N_16941);
nand U17777 (N_17777,N_17236,N_16877);
nor U17778 (N_17778,N_16947,N_16888);
nor U17779 (N_17779,N_17143,N_17343);
or U17780 (N_17780,N_17061,N_17366);
nor U17781 (N_17781,N_16892,N_16902);
nor U17782 (N_17782,N_17460,N_17372);
nor U17783 (N_17783,N_17330,N_17224);
nor U17784 (N_17784,N_17488,N_16948);
nand U17785 (N_17785,N_17486,N_17327);
nor U17786 (N_17786,N_17207,N_17271);
and U17787 (N_17787,N_16981,N_17415);
xor U17788 (N_17788,N_17002,N_17088);
or U17789 (N_17789,N_17348,N_17286);
xnor U17790 (N_17790,N_16997,N_17404);
nor U17791 (N_17791,N_16921,N_17165);
nor U17792 (N_17792,N_17252,N_17462);
and U17793 (N_17793,N_17049,N_17239);
and U17794 (N_17794,N_17024,N_17106);
nand U17795 (N_17795,N_17350,N_17298);
nand U17796 (N_17796,N_17009,N_17010);
and U17797 (N_17797,N_17206,N_17136);
nand U17798 (N_17798,N_17117,N_16946);
nor U17799 (N_17799,N_17057,N_17006);
nor U17800 (N_17800,N_17084,N_17169);
nand U17801 (N_17801,N_17254,N_17451);
or U17802 (N_17802,N_17171,N_17242);
nand U17803 (N_17803,N_17401,N_16998);
or U17804 (N_17804,N_17456,N_17412);
nand U17805 (N_17805,N_17384,N_17443);
and U17806 (N_17806,N_17019,N_17166);
nor U17807 (N_17807,N_17093,N_17097);
xor U17808 (N_17808,N_17251,N_17246);
nand U17809 (N_17809,N_17409,N_17345);
nor U17810 (N_17810,N_17442,N_17367);
or U17811 (N_17811,N_17177,N_17154);
or U17812 (N_17812,N_16924,N_17251);
nor U17813 (N_17813,N_17181,N_16903);
and U17814 (N_17814,N_17447,N_16896);
and U17815 (N_17815,N_17320,N_17222);
nor U17816 (N_17816,N_17480,N_16934);
nor U17817 (N_17817,N_17490,N_16944);
xnor U17818 (N_17818,N_17218,N_16996);
nand U17819 (N_17819,N_17496,N_17092);
xnor U17820 (N_17820,N_16890,N_17467);
nor U17821 (N_17821,N_17308,N_17030);
and U17822 (N_17822,N_17315,N_17174);
and U17823 (N_17823,N_17472,N_17433);
nand U17824 (N_17824,N_17075,N_16902);
xor U17825 (N_17825,N_17155,N_16909);
xor U17826 (N_17826,N_16974,N_17105);
nand U17827 (N_17827,N_17470,N_17241);
nand U17828 (N_17828,N_17320,N_17272);
or U17829 (N_17829,N_16996,N_17386);
or U17830 (N_17830,N_17461,N_17061);
nand U17831 (N_17831,N_17205,N_17425);
or U17832 (N_17832,N_17374,N_17430);
and U17833 (N_17833,N_17389,N_17460);
or U17834 (N_17834,N_17107,N_17321);
and U17835 (N_17835,N_16980,N_17081);
xnor U17836 (N_17836,N_17075,N_17215);
or U17837 (N_17837,N_16912,N_17295);
and U17838 (N_17838,N_17288,N_17459);
or U17839 (N_17839,N_17074,N_17045);
nor U17840 (N_17840,N_16951,N_17098);
nor U17841 (N_17841,N_17305,N_17261);
nand U17842 (N_17842,N_17108,N_17316);
or U17843 (N_17843,N_17122,N_17478);
and U17844 (N_17844,N_16900,N_17269);
and U17845 (N_17845,N_17076,N_17062);
nor U17846 (N_17846,N_17489,N_17214);
or U17847 (N_17847,N_17294,N_17173);
nor U17848 (N_17848,N_16942,N_17192);
and U17849 (N_17849,N_16934,N_17217);
or U17850 (N_17850,N_17006,N_17318);
nor U17851 (N_17851,N_17037,N_16927);
or U17852 (N_17852,N_17208,N_16916);
and U17853 (N_17853,N_16900,N_17344);
nor U17854 (N_17854,N_17250,N_17321);
or U17855 (N_17855,N_16982,N_17337);
nor U17856 (N_17856,N_17239,N_16893);
nand U17857 (N_17857,N_16911,N_17132);
nor U17858 (N_17858,N_17451,N_17461);
xnor U17859 (N_17859,N_17106,N_16978);
nand U17860 (N_17860,N_17182,N_17459);
nor U17861 (N_17861,N_16914,N_16997);
or U17862 (N_17862,N_16943,N_17200);
and U17863 (N_17863,N_17251,N_17017);
nor U17864 (N_17864,N_16897,N_16998);
or U17865 (N_17865,N_17444,N_17074);
nor U17866 (N_17866,N_17040,N_17213);
or U17867 (N_17867,N_17410,N_17241);
nand U17868 (N_17868,N_17205,N_17276);
and U17869 (N_17869,N_17109,N_17392);
nor U17870 (N_17870,N_17291,N_17074);
nand U17871 (N_17871,N_17309,N_17104);
nor U17872 (N_17872,N_16883,N_17034);
nand U17873 (N_17873,N_17249,N_16911);
or U17874 (N_17874,N_17420,N_17072);
nand U17875 (N_17875,N_16920,N_17277);
or U17876 (N_17876,N_17043,N_17401);
and U17877 (N_17877,N_17459,N_17217);
nand U17878 (N_17878,N_17127,N_17315);
nand U17879 (N_17879,N_16967,N_17122);
and U17880 (N_17880,N_17063,N_17336);
and U17881 (N_17881,N_17327,N_17487);
or U17882 (N_17882,N_17285,N_17183);
xnor U17883 (N_17883,N_17276,N_17399);
nor U17884 (N_17884,N_17225,N_17139);
nand U17885 (N_17885,N_17197,N_17491);
nor U17886 (N_17886,N_17205,N_16948);
nor U17887 (N_17887,N_17281,N_17170);
xor U17888 (N_17888,N_17464,N_17402);
nor U17889 (N_17889,N_17386,N_17141);
or U17890 (N_17890,N_17213,N_17402);
and U17891 (N_17891,N_17089,N_17374);
or U17892 (N_17892,N_17370,N_17372);
or U17893 (N_17893,N_17093,N_17264);
or U17894 (N_17894,N_17004,N_17486);
nor U17895 (N_17895,N_17166,N_17236);
or U17896 (N_17896,N_17113,N_16902);
or U17897 (N_17897,N_17080,N_17045);
or U17898 (N_17898,N_17405,N_16946);
or U17899 (N_17899,N_17092,N_17483);
nor U17900 (N_17900,N_17010,N_16921);
nand U17901 (N_17901,N_17385,N_17355);
and U17902 (N_17902,N_16967,N_17063);
xor U17903 (N_17903,N_17094,N_17437);
nor U17904 (N_17904,N_17120,N_17144);
or U17905 (N_17905,N_17251,N_17235);
nor U17906 (N_17906,N_17369,N_17425);
nand U17907 (N_17907,N_17372,N_17064);
nand U17908 (N_17908,N_17467,N_17060);
and U17909 (N_17909,N_17133,N_17178);
nor U17910 (N_17910,N_17246,N_17298);
or U17911 (N_17911,N_17076,N_16935);
or U17912 (N_17912,N_17177,N_17083);
and U17913 (N_17913,N_17472,N_17425);
or U17914 (N_17914,N_17100,N_16962);
and U17915 (N_17915,N_17053,N_17383);
nand U17916 (N_17916,N_17332,N_17133);
nand U17917 (N_17917,N_17422,N_17105);
and U17918 (N_17918,N_17210,N_17324);
and U17919 (N_17919,N_17241,N_17467);
or U17920 (N_17920,N_17475,N_17283);
or U17921 (N_17921,N_17121,N_17068);
nor U17922 (N_17922,N_17113,N_17088);
and U17923 (N_17923,N_17457,N_17138);
and U17924 (N_17924,N_16924,N_17008);
nand U17925 (N_17925,N_17089,N_17366);
xnor U17926 (N_17926,N_16934,N_17330);
xor U17927 (N_17927,N_17226,N_17463);
nand U17928 (N_17928,N_17467,N_17258);
or U17929 (N_17929,N_16897,N_17366);
and U17930 (N_17930,N_16904,N_16988);
xnor U17931 (N_17931,N_17491,N_17024);
nor U17932 (N_17932,N_17344,N_17115);
nand U17933 (N_17933,N_17492,N_17288);
nor U17934 (N_17934,N_17449,N_17371);
nor U17935 (N_17935,N_17326,N_17167);
and U17936 (N_17936,N_17289,N_17037);
nand U17937 (N_17937,N_17121,N_17050);
or U17938 (N_17938,N_16980,N_17134);
nor U17939 (N_17939,N_17034,N_17246);
or U17940 (N_17940,N_16979,N_17429);
nor U17941 (N_17941,N_17494,N_17484);
nor U17942 (N_17942,N_16926,N_17188);
nand U17943 (N_17943,N_16895,N_17499);
xnor U17944 (N_17944,N_17350,N_16892);
and U17945 (N_17945,N_17161,N_17026);
xnor U17946 (N_17946,N_17425,N_17279);
or U17947 (N_17947,N_17255,N_17179);
and U17948 (N_17948,N_17443,N_17042);
and U17949 (N_17949,N_17496,N_17250);
nor U17950 (N_17950,N_17017,N_17478);
and U17951 (N_17951,N_16878,N_17427);
or U17952 (N_17952,N_16941,N_17493);
nor U17953 (N_17953,N_16876,N_17093);
nand U17954 (N_17954,N_16943,N_17376);
and U17955 (N_17955,N_16880,N_16963);
nand U17956 (N_17956,N_17479,N_17246);
nand U17957 (N_17957,N_17330,N_17192);
and U17958 (N_17958,N_17125,N_17187);
nand U17959 (N_17959,N_17438,N_17347);
nand U17960 (N_17960,N_17242,N_17004);
and U17961 (N_17961,N_17237,N_16932);
nand U17962 (N_17962,N_17198,N_17378);
or U17963 (N_17963,N_17429,N_17365);
and U17964 (N_17964,N_17277,N_16930);
nor U17965 (N_17965,N_17048,N_17070);
xor U17966 (N_17966,N_16919,N_17005);
and U17967 (N_17967,N_17493,N_17496);
and U17968 (N_17968,N_17100,N_17361);
and U17969 (N_17969,N_17290,N_16944);
nand U17970 (N_17970,N_17322,N_17091);
nor U17971 (N_17971,N_17182,N_17279);
xor U17972 (N_17972,N_17002,N_17019);
nor U17973 (N_17973,N_17478,N_17052);
nor U17974 (N_17974,N_17428,N_17203);
xnor U17975 (N_17975,N_16912,N_17235);
or U17976 (N_17976,N_17012,N_17218);
and U17977 (N_17977,N_17173,N_17019);
or U17978 (N_17978,N_17056,N_17357);
nand U17979 (N_17979,N_17083,N_16888);
and U17980 (N_17980,N_17300,N_17107);
or U17981 (N_17981,N_17074,N_17434);
xor U17982 (N_17982,N_17355,N_17201);
nor U17983 (N_17983,N_16907,N_17342);
nand U17984 (N_17984,N_17448,N_17339);
nor U17985 (N_17985,N_17128,N_17324);
or U17986 (N_17986,N_17097,N_16970);
and U17987 (N_17987,N_17374,N_17487);
nor U17988 (N_17988,N_16899,N_17214);
nand U17989 (N_17989,N_17200,N_17366);
or U17990 (N_17990,N_17177,N_17441);
xor U17991 (N_17991,N_17112,N_17310);
nand U17992 (N_17992,N_17036,N_16878);
nor U17993 (N_17993,N_16939,N_17180);
nand U17994 (N_17994,N_17062,N_17201);
or U17995 (N_17995,N_17288,N_17497);
nor U17996 (N_17996,N_16875,N_17314);
and U17997 (N_17997,N_17447,N_17432);
nor U17998 (N_17998,N_17432,N_16946);
and U17999 (N_17999,N_17331,N_17358);
and U18000 (N_18000,N_17375,N_17377);
nand U18001 (N_18001,N_17455,N_17043);
and U18002 (N_18002,N_16975,N_17096);
and U18003 (N_18003,N_17484,N_16919);
nor U18004 (N_18004,N_17217,N_17285);
nand U18005 (N_18005,N_17436,N_17416);
xor U18006 (N_18006,N_16938,N_17043);
nand U18007 (N_18007,N_17465,N_17459);
nor U18008 (N_18008,N_17336,N_17485);
nand U18009 (N_18009,N_17149,N_16958);
nand U18010 (N_18010,N_17032,N_17004);
nor U18011 (N_18011,N_17037,N_17042);
or U18012 (N_18012,N_17430,N_17238);
and U18013 (N_18013,N_16951,N_17429);
or U18014 (N_18014,N_17224,N_17262);
or U18015 (N_18015,N_17457,N_17052);
and U18016 (N_18016,N_17215,N_17223);
xor U18017 (N_18017,N_17254,N_17072);
and U18018 (N_18018,N_17172,N_17211);
and U18019 (N_18019,N_17422,N_17397);
and U18020 (N_18020,N_16992,N_17099);
and U18021 (N_18021,N_16988,N_17339);
or U18022 (N_18022,N_17202,N_17047);
nand U18023 (N_18023,N_17066,N_17185);
and U18024 (N_18024,N_17150,N_16993);
and U18025 (N_18025,N_17310,N_16907);
xor U18026 (N_18026,N_17256,N_17077);
nand U18027 (N_18027,N_17487,N_17110);
or U18028 (N_18028,N_17045,N_17178);
nand U18029 (N_18029,N_16895,N_17235);
xnor U18030 (N_18030,N_17297,N_17371);
nor U18031 (N_18031,N_17356,N_17120);
nor U18032 (N_18032,N_17229,N_17235);
nand U18033 (N_18033,N_17017,N_17098);
or U18034 (N_18034,N_17116,N_17368);
and U18035 (N_18035,N_17422,N_17190);
and U18036 (N_18036,N_16967,N_17268);
nor U18037 (N_18037,N_17329,N_17094);
nand U18038 (N_18038,N_17315,N_17042);
or U18039 (N_18039,N_17072,N_17276);
nor U18040 (N_18040,N_17082,N_17243);
or U18041 (N_18041,N_17217,N_17353);
nand U18042 (N_18042,N_17178,N_16902);
and U18043 (N_18043,N_17476,N_17312);
nor U18044 (N_18044,N_17346,N_17017);
nor U18045 (N_18045,N_17162,N_17256);
and U18046 (N_18046,N_17406,N_17457);
nand U18047 (N_18047,N_17186,N_17416);
nor U18048 (N_18048,N_17308,N_17032);
nand U18049 (N_18049,N_17286,N_17496);
xnor U18050 (N_18050,N_17471,N_17305);
xnor U18051 (N_18051,N_17358,N_17102);
nand U18052 (N_18052,N_17281,N_17457);
and U18053 (N_18053,N_17386,N_17382);
or U18054 (N_18054,N_17358,N_16966);
or U18055 (N_18055,N_17499,N_17199);
and U18056 (N_18056,N_17070,N_17448);
or U18057 (N_18057,N_17237,N_17483);
or U18058 (N_18058,N_16988,N_17069);
or U18059 (N_18059,N_17137,N_17315);
nor U18060 (N_18060,N_17230,N_17141);
and U18061 (N_18061,N_16970,N_16921);
nor U18062 (N_18062,N_17361,N_17000);
nor U18063 (N_18063,N_16963,N_16917);
nor U18064 (N_18064,N_17315,N_17480);
nand U18065 (N_18065,N_16990,N_17402);
nand U18066 (N_18066,N_16966,N_17439);
nand U18067 (N_18067,N_17488,N_17413);
and U18068 (N_18068,N_17219,N_17182);
or U18069 (N_18069,N_17394,N_17449);
and U18070 (N_18070,N_17144,N_17036);
nor U18071 (N_18071,N_17077,N_17053);
nand U18072 (N_18072,N_17314,N_17367);
nor U18073 (N_18073,N_17278,N_17314);
nand U18074 (N_18074,N_17086,N_17069);
nor U18075 (N_18075,N_17248,N_17097);
xnor U18076 (N_18076,N_16924,N_17401);
nand U18077 (N_18077,N_17225,N_17186);
nand U18078 (N_18078,N_17260,N_16989);
or U18079 (N_18079,N_17201,N_17272);
or U18080 (N_18080,N_17267,N_17451);
or U18081 (N_18081,N_17386,N_16911);
and U18082 (N_18082,N_17431,N_16959);
xnor U18083 (N_18083,N_16898,N_16998);
nor U18084 (N_18084,N_17179,N_17345);
and U18085 (N_18085,N_16913,N_16957);
nand U18086 (N_18086,N_17113,N_17057);
nand U18087 (N_18087,N_17053,N_17215);
or U18088 (N_18088,N_17188,N_17115);
nand U18089 (N_18089,N_17055,N_17232);
nand U18090 (N_18090,N_17408,N_16950);
or U18091 (N_18091,N_17232,N_17479);
or U18092 (N_18092,N_17273,N_17083);
and U18093 (N_18093,N_17205,N_17481);
nand U18094 (N_18094,N_16969,N_17047);
nor U18095 (N_18095,N_17258,N_17278);
or U18096 (N_18096,N_17329,N_17212);
nor U18097 (N_18097,N_16879,N_17323);
or U18098 (N_18098,N_17030,N_17027);
nor U18099 (N_18099,N_17285,N_17450);
and U18100 (N_18100,N_16935,N_17308);
and U18101 (N_18101,N_17101,N_17030);
nor U18102 (N_18102,N_17343,N_17383);
nand U18103 (N_18103,N_17428,N_17492);
nor U18104 (N_18104,N_17011,N_17452);
and U18105 (N_18105,N_17353,N_17485);
or U18106 (N_18106,N_17123,N_17049);
nand U18107 (N_18107,N_17000,N_17498);
xor U18108 (N_18108,N_16995,N_17209);
xnor U18109 (N_18109,N_17400,N_16974);
nor U18110 (N_18110,N_17225,N_17365);
xnor U18111 (N_18111,N_17199,N_16971);
nor U18112 (N_18112,N_16990,N_17209);
or U18113 (N_18113,N_16944,N_17305);
nor U18114 (N_18114,N_16941,N_17358);
nor U18115 (N_18115,N_17002,N_16988);
xor U18116 (N_18116,N_17141,N_17209);
and U18117 (N_18117,N_17313,N_17284);
xnor U18118 (N_18118,N_17211,N_17160);
or U18119 (N_18119,N_16969,N_17200);
or U18120 (N_18120,N_16909,N_17207);
nor U18121 (N_18121,N_17381,N_16930);
nor U18122 (N_18122,N_16914,N_16920);
or U18123 (N_18123,N_17037,N_16883);
nand U18124 (N_18124,N_17337,N_17397);
and U18125 (N_18125,N_17756,N_17559);
nor U18126 (N_18126,N_17708,N_17686);
nand U18127 (N_18127,N_17579,N_17969);
nand U18128 (N_18128,N_17507,N_17654);
nand U18129 (N_18129,N_17752,N_17778);
nand U18130 (N_18130,N_17548,N_17854);
or U18131 (N_18131,N_18086,N_17881);
or U18132 (N_18132,N_17744,N_18055);
and U18133 (N_18133,N_17924,N_17672);
or U18134 (N_18134,N_17605,N_17642);
or U18135 (N_18135,N_17821,N_17758);
or U18136 (N_18136,N_17864,N_18075);
or U18137 (N_18137,N_17814,N_17954);
xor U18138 (N_18138,N_17721,N_17733);
and U18139 (N_18139,N_17957,N_17989);
nor U18140 (N_18140,N_17658,N_17594);
nand U18141 (N_18141,N_17953,N_17618);
and U18142 (N_18142,N_18056,N_17998);
nand U18143 (N_18143,N_17556,N_17676);
or U18144 (N_18144,N_17608,N_17857);
or U18145 (N_18145,N_17921,N_18046);
nand U18146 (N_18146,N_17941,N_17757);
or U18147 (N_18147,N_17952,N_18044);
nand U18148 (N_18148,N_17662,N_18053);
or U18149 (N_18149,N_17585,N_17689);
or U18150 (N_18150,N_18094,N_17684);
nor U18151 (N_18151,N_17877,N_17976);
and U18152 (N_18152,N_18040,N_18028);
and U18153 (N_18153,N_17745,N_17697);
and U18154 (N_18154,N_17502,N_17932);
and U18155 (N_18155,N_17902,N_17996);
or U18156 (N_18156,N_17698,N_17865);
nor U18157 (N_18157,N_17533,N_17500);
or U18158 (N_18158,N_17732,N_18101);
or U18159 (N_18159,N_17804,N_17798);
and U18160 (N_18160,N_17611,N_17616);
nor U18161 (N_18161,N_17771,N_17833);
nor U18162 (N_18162,N_17977,N_17550);
and U18163 (N_18163,N_17925,N_18084);
nor U18164 (N_18164,N_17772,N_18027);
nor U18165 (N_18165,N_17781,N_17888);
nand U18166 (N_18166,N_17918,N_17527);
and U18167 (N_18167,N_17828,N_17809);
nand U18168 (N_18168,N_17631,N_17589);
xor U18169 (N_18169,N_17749,N_18010);
nand U18170 (N_18170,N_17838,N_17841);
nand U18171 (N_18171,N_18079,N_17903);
nor U18172 (N_18172,N_17670,N_17719);
and U18173 (N_18173,N_17806,N_18004);
or U18174 (N_18174,N_17907,N_17629);
xor U18175 (N_18175,N_17805,N_17819);
and U18176 (N_18176,N_17965,N_17598);
nor U18177 (N_18177,N_18097,N_18018);
and U18178 (N_18178,N_17650,N_17935);
or U18179 (N_18179,N_17609,N_17825);
or U18180 (N_18180,N_18108,N_17648);
xnor U18181 (N_18181,N_17788,N_17984);
xnor U18182 (N_18182,N_17722,N_17766);
nor U18183 (N_18183,N_17999,N_18090);
or U18184 (N_18184,N_17547,N_18005);
or U18185 (N_18185,N_17668,N_17940);
and U18186 (N_18186,N_17955,N_17807);
and U18187 (N_18187,N_17554,N_17621);
and U18188 (N_18188,N_17920,N_17718);
and U18189 (N_18189,N_17612,N_17937);
xor U18190 (N_18190,N_17770,N_17894);
xor U18191 (N_18191,N_17826,N_17529);
nand U18192 (N_18192,N_17704,N_17649);
nand U18193 (N_18193,N_17614,N_18045);
xnor U18194 (N_18194,N_17970,N_18054);
nand U18195 (N_18195,N_17678,N_17567);
or U18196 (N_18196,N_17593,N_17961);
and U18197 (N_18197,N_17503,N_17905);
nor U18198 (N_18198,N_17730,N_17523);
and U18199 (N_18199,N_17768,N_18059);
and U18200 (N_18200,N_18074,N_18122);
nor U18201 (N_18201,N_18111,N_17844);
nand U18202 (N_18202,N_17876,N_17873);
or U18203 (N_18203,N_17975,N_17724);
or U18204 (N_18204,N_17812,N_17521);
or U18205 (N_18205,N_17510,N_18070);
nor U18206 (N_18206,N_17960,N_17696);
or U18207 (N_18207,N_18106,N_18049);
nor U18208 (N_18208,N_17640,N_18008);
nand U18209 (N_18209,N_17701,N_17728);
nor U18210 (N_18210,N_17705,N_17536);
or U18211 (N_18211,N_17762,N_17799);
or U18212 (N_18212,N_17685,N_17513);
nor U18213 (N_18213,N_17851,N_17600);
nor U18214 (N_18214,N_17586,N_18093);
xnor U18215 (N_18215,N_17775,N_18073);
or U18216 (N_18216,N_17540,N_17963);
xor U18217 (N_18217,N_18117,N_17761);
or U18218 (N_18218,N_17584,N_17610);
xor U18219 (N_18219,N_17982,N_17546);
and U18220 (N_18220,N_17782,N_17707);
xor U18221 (N_18221,N_17561,N_18007);
nor U18222 (N_18222,N_17945,N_18031);
xnor U18223 (N_18223,N_17747,N_17638);
nor U18224 (N_18224,N_17994,N_17580);
or U18225 (N_18225,N_17874,N_17769);
nand U18226 (N_18226,N_17964,N_17538);
or U18227 (N_18227,N_17832,N_17843);
nand U18228 (N_18228,N_18113,N_17987);
or U18229 (N_18229,N_17870,N_18114);
nand U18230 (N_18230,N_17751,N_18095);
nor U18231 (N_18231,N_17802,N_17635);
xnor U18232 (N_18232,N_17531,N_17632);
xor U18233 (N_18233,N_17690,N_18051);
or U18234 (N_18234,N_17607,N_18047);
nor U18235 (N_18235,N_17777,N_17665);
nor U18236 (N_18236,N_17817,N_17947);
or U18237 (N_18237,N_17726,N_17505);
or U18238 (N_18238,N_17501,N_18064);
or U18239 (N_18239,N_17880,N_17655);
xnor U18240 (N_18240,N_17716,N_17700);
nand U18241 (N_18241,N_17891,N_17801);
nor U18242 (N_18242,N_18060,N_17958);
and U18243 (N_18243,N_17581,N_17552);
nor U18244 (N_18244,N_17675,N_17951);
or U18245 (N_18245,N_18082,N_17934);
and U18246 (N_18246,N_17897,N_17827);
nand U18247 (N_18247,N_17741,N_18042);
nand U18248 (N_18248,N_17995,N_17712);
nand U18249 (N_18249,N_17816,N_17985);
and U18250 (N_18250,N_18015,N_17750);
nor U18251 (N_18251,N_17783,N_17646);
nand U18252 (N_18252,N_17717,N_17867);
nor U18253 (N_18253,N_17911,N_18119);
and U18254 (N_18254,N_17626,N_17709);
nand U18255 (N_18255,N_17908,N_17639);
nor U18256 (N_18256,N_17822,N_17810);
nor U18257 (N_18257,N_18072,N_17524);
or U18258 (N_18258,N_18038,N_18071);
and U18259 (N_18259,N_17660,N_18061);
xor U18260 (N_18260,N_17780,N_17659);
or U18261 (N_18261,N_18034,N_17691);
nor U18262 (N_18262,N_18002,N_17846);
and U18263 (N_18263,N_17915,N_17791);
nor U18264 (N_18264,N_17919,N_17590);
or U18265 (N_18265,N_18088,N_18012);
xnor U18266 (N_18266,N_17837,N_17517);
or U18267 (N_18267,N_17560,N_18091);
nand U18268 (N_18268,N_17574,N_17991);
or U18269 (N_18269,N_18033,N_17742);
or U18270 (N_18270,N_17656,N_18096);
nand U18271 (N_18271,N_17636,N_17884);
nand U18272 (N_18272,N_17959,N_17988);
nor U18273 (N_18273,N_18120,N_17606);
nand U18274 (N_18274,N_18016,N_17850);
or U18275 (N_18275,N_17504,N_17723);
nand U18276 (N_18276,N_18115,N_17519);
or U18277 (N_18277,N_17784,N_17889);
nor U18278 (N_18278,N_18116,N_17759);
nor U18279 (N_18279,N_18087,N_18069);
xor U18280 (N_18280,N_17644,N_17542);
nor U18281 (N_18281,N_17871,N_17647);
or U18282 (N_18282,N_18026,N_18036);
and U18283 (N_18283,N_18021,N_18067);
nor U18284 (N_18284,N_17683,N_17949);
and U18285 (N_18285,N_17824,N_17910);
and U18286 (N_18286,N_17901,N_17736);
or U18287 (N_18287,N_17673,N_17859);
nand U18288 (N_18288,N_17620,N_17776);
xor U18289 (N_18289,N_17852,N_17922);
or U18290 (N_18290,N_17702,N_18104);
nand U18291 (N_18291,N_18019,N_17792);
and U18292 (N_18292,N_17823,N_17514);
or U18293 (N_18293,N_18078,N_17667);
and U18294 (N_18294,N_17653,N_17595);
or U18295 (N_18295,N_17558,N_18098);
or U18296 (N_18296,N_17830,N_17652);
nand U18297 (N_18297,N_17848,N_17875);
nand U18298 (N_18298,N_18014,N_17680);
nand U18299 (N_18299,N_17928,N_17890);
nand U18300 (N_18300,N_17914,N_17624);
nor U18301 (N_18301,N_17617,N_17882);
and U18302 (N_18302,N_17737,N_17643);
nor U18303 (N_18303,N_17666,N_17734);
nor U18304 (N_18304,N_17516,N_17604);
or U18305 (N_18305,N_17509,N_17869);
nor U18306 (N_18306,N_17633,N_17714);
nor U18307 (N_18307,N_17811,N_17980);
or U18308 (N_18308,N_17909,N_18013);
nand U18309 (N_18309,N_17535,N_17856);
nor U18310 (N_18310,N_17829,N_17942);
and U18311 (N_18311,N_17973,N_18011);
nand U18312 (N_18312,N_17571,N_17966);
nand U18313 (N_18313,N_18035,N_18066);
or U18314 (N_18314,N_17615,N_18025);
xor U18315 (N_18315,N_17883,N_18085);
xor U18316 (N_18316,N_17743,N_18058);
nand U18317 (N_18317,N_17948,N_17863);
and U18318 (N_18318,N_17855,N_17886);
nand U18319 (N_18319,N_17622,N_17834);
or U18320 (N_18320,N_17979,N_17862);
nand U18321 (N_18321,N_17895,N_17564);
nand U18322 (N_18322,N_17511,N_17602);
nor U18323 (N_18323,N_17603,N_17860);
and U18324 (N_18324,N_17694,N_17840);
nor U18325 (N_18325,N_18077,N_17861);
nand U18326 (N_18326,N_17893,N_17986);
xnor U18327 (N_18327,N_18043,N_17568);
and U18328 (N_18328,N_17849,N_17787);
xnor U18329 (N_18329,N_17779,N_17657);
or U18330 (N_18330,N_17773,N_17713);
and U18331 (N_18331,N_17900,N_17926);
nor U18332 (N_18332,N_18112,N_17695);
or U18333 (N_18333,N_17572,N_18032);
nor U18334 (N_18334,N_18068,N_17518);
and U18335 (N_18335,N_17687,N_17931);
or U18336 (N_18336,N_17577,N_17727);
nor U18337 (N_18337,N_17930,N_17813);
or U18338 (N_18338,N_17936,N_17929);
nor U18339 (N_18339,N_17946,N_17663);
or U18340 (N_18340,N_17836,N_17754);
nor U18341 (N_18341,N_17767,N_18118);
or U18342 (N_18342,N_17575,N_17619);
or U18343 (N_18343,N_17566,N_17790);
nand U18344 (N_18344,N_17868,N_17710);
and U18345 (N_18345,N_17537,N_18076);
and U18346 (N_18346,N_18039,N_18022);
nand U18347 (N_18347,N_17753,N_17699);
and U18348 (N_18348,N_17508,N_18057);
nor U18349 (N_18349,N_17587,N_17847);
nor U18350 (N_18350,N_17725,N_17715);
nand U18351 (N_18351,N_17576,N_17944);
or U18352 (N_18352,N_17968,N_17927);
and U18353 (N_18353,N_18089,N_17962);
nand U18354 (N_18354,N_18121,N_17532);
nand U18355 (N_18355,N_17755,N_17591);
xnor U18356 (N_18356,N_17746,N_17800);
or U18357 (N_18357,N_17565,N_17764);
xnor U18358 (N_18358,N_17793,N_17740);
nor U18359 (N_18359,N_18123,N_17872);
nand U18360 (N_18360,N_17879,N_17627);
nand U18361 (N_18361,N_17526,N_18110);
nand U18362 (N_18362,N_17534,N_18023);
nand U18363 (N_18363,N_17628,N_17543);
nor U18364 (N_18364,N_17917,N_17803);
nand U18365 (N_18365,N_18020,N_18080);
xnor U18366 (N_18366,N_17645,N_18006);
nand U18367 (N_18367,N_17735,N_17679);
and U18368 (N_18368,N_17731,N_17899);
xnor U18369 (N_18369,N_17553,N_17703);
nand U18370 (N_18370,N_17938,N_18009);
xnor U18371 (N_18371,N_17520,N_18083);
and U18372 (N_18372,N_17858,N_17885);
nor U18373 (N_18373,N_17866,N_17916);
and U18374 (N_18374,N_17739,N_17981);
nor U18375 (N_18375,N_17669,N_17748);
or U18376 (N_18376,N_17923,N_17671);
and U18377 (N_18377,N_18062,N_18065);
or U18378 (N_18378,N_18037,N_17878);
nor U18379 (N_18379,N_17797,N_17651);
or U18380 (N_18380,N_17613,N_18063);
nand U18381 (N_18381,N_17528,N_17939);
and U18382 (N_18382,N_18050,N_17637);
xor U18383 (N_18383,N_17990,N_17539);
nand U18384 (N_18384,N_17786,N_17692);
or U18385 (N_18385,N_17842,N_17625);
and U18386 (N_18386,N_17808,N_17570);
nor U18387 (N_18387,N_18099,N_17818);
nor U18388 (N_18388,N_17515,N_17892);
and U18389 (N_18389,N_17592,N_17898);
nand U18390 (N_18390,N_18103,N_17688);
xnor U18391 (N_18391,N_17738,N_17555);
and U18392 (N_18392,N_17630,N_17912);
and U18393 (N_18393,N_17729,N_17763);
nor U18394 (N_18394,N_17972,N_17997);
and U18395 (N_18395,N_17795,N_17971);
nor U18396 (N_18396,N_17682,N_17943);
and U18397 (N_18397,N_17563,N_17796);
and U18398 (N_18398,N_17588,N_17760);
nor U18399 (N_18399,N_18092,N_17569);
nor U18400 (N_18400,N_17544,N_17506);
nor U18401 (N_18401,N_17839,N_17557);
or U18402 (N_18402,N_17512,N_17794);
nor U18403 (N_18403,N_17674,N_17820);
or U18404 (N_18404,N_17582,N_18001);
nand U18405 (N_18405,N_17573,N_18124);
nor U18406 (N_18406,N_17983,N_17765);
nor U18407 (N_18407,N_18017,N_17597);
nand U18408 (N_18408,N_17677,N_17693);
and U18409 (N_18409,N_17541,N_17774);
nor U18410 (N_18410,N_17562,N_18000);
or U18411 (N_18411,N_17596,N_17661);
nor U18412 (N_18412,N_18041,N_18048);
nand U18413 (N_18413,N_18003,N_17545);
nor U18414 (N_18414,N_17720,N_17525);
nor U18415 (N_18415,N_17992,N_17789);
nor U18416 (N_18416,N_17601,N_18081);
or U18417 (N_18417,N_17950,N_17578);
and U18418 (N_18418,N_17835,N_17711);
nor U18419 (N_18419,N_18029,N_17623);
nand U18420 (N_18420,N_18030,N_17974);
nand U18421 (N_18421,N_18102,N_17583);
nor U18422 (N_18422,N_17634,N_17530);
nand U18423 (N_18423,N_17785,N_17815);
xnor U18424 (N_18424,N_17896,N_18100);
or U18425 (N_18425,N_17956,N_18109);
nor U18426 (N_18426,N_17993,N_17641);
or U18427 (N_18427,N_17551,N_18107);
nand U18428 (N_18428,N_17904,N_17706);
or U18429 (N_18429,N_17978,N_17522);
nor U18430 (N_18430,N_17906,N_17845);
nand U18431 (N_18431,N_17664,N_18024);
and U18432 (N_18432,N_17887,N_18105);
nor U18433 (N_18433,N_17933,N_17681);
or U18434 (N_18434,N_17967,N_17549);
nand U18435 (N_18435,N_17853,N_17831);
nor U18436 (N_18436,N_17913,N_17599);
or U18437 (N_18437,N_18052,N_17924);
and U18438 (N_18438,N_17879,N_17934);
xnor U18439 (N_18439,N_17965,N_17690);
nand U18440 (N_18440,N_17901,N_18081);
or U18441 (N_18441,N_17936,N_17669);
nand U18442 (N_18442,N_17886,N_18053);
nand U18443 (N_18443,N_17690,N_17504);
nor U18444 (N_18444,N_17675,N_17636);
nand U18445 (N_18445,N_18067,N_17691);
nor U18446 (N_18446,N_17756,N_17637);
or U18447 (N_18447,N_17584,N_17866);
or U18448 (N_18448,N_17657,N_18033);
nand U18449 (N_18449,N_17675,N_17595);
and U18450 (N_18450,N_18064,N_18010);
and U18451 (N_18451,N_18056,N_17869);
nor U18452 (N_18452,N_17520,N_17864);
xnor U18453 (N_18453,N_17586,N_17692);
and U18454 (N_18454,N_18072,N_17837);
nand U18455 (N_18455,N_18048,N_17821);
nor U18456 (N_18456,N_18004,N_17622);
nor U18457 (N_18457,N_17889,N_17677);
nand U18458 (N_18458,N_17662,N_18029);
nor U18459 (N_18459,N_17684,N_17693);
or U18460 (N_18460,N_17885,N_17953);
nor U18461 (N_18461,N_18099,N_17887);
and U18462 (N_18462,N_17941,N_17800);
or U18463 (N_18463,N_17619,N_18052);
xnor U18464 (N_18464,N_17886,N_17913);
xor U18465 (N_18465,N_17590,N_17527);
or U18466 (N_18466,N_18115,N_18054);
and U18467 (N_18467,N_17859,N_17885);
or U18468 (N_18468,N_17740,N_17577);
and U18469 (N_18469,N_18070,N_18008);
or U18470 (N_18470,N_17794,N_17723);
xnor U18471 (N_18471,N_17540,N_17739);
and U18472 (N_18472,N_17616,N_18023);
nand U18473 (N_18473,N_17979,N_17619);
nand U18474 (N_18474,N_17600,N_17631);
or U18475 (N_18475,N_17520,N_18026);
nand U18476 (N_18476,N_17552,N_17510);
nand U18477 (N_18477,N_17794,N_18047);
xnor U18478 (N_18478,N_18121,N_17901);
nand U18479 (N_18479,N_18074,N_17680);
and U18480 (N_18480,N_17527,N_17753);
nor U18481 (N_18481,N_17715,N_17693);
or U18482 (N_18482,N_17794,N_17709);
or U18483 (N_18483,N_17949,N_17522);
and U18484 (N_18484,N_17868,N_17605);
or U18485 (N_18485,N_17792,N_17995);
nand U18486 (N_18486,N_18001,N_17774);
xor U18487 (N_18487,N_17897,N_18116);
and U18488 (N_18488,N_17533,N_17930);
nor U18489 (N_18489,N_18100,N_17973);
xnor U18490 (N_18490,N_17526,N_17782);
nor U18491 (N_18491,N_18047,N_17812);
and U18492 (N_18492,N_17875,N_17500);
nand U18493 (N_18493,N_17682,N_17597);
nand U18494 (N_18494,N_17813,N_17810);
and U18495 (N_18495,N_17528,N_18026);
nand U18496 (N_18496,N_18090,N_18030);
and U18497 (N_18497,N_17637,N_17881);
nand U18498 (N_18498,N_18048,N_17744);
nand U18499 (N_18499,N_17935,N_18018);
and U18500 (N_18500,N_17955,N_17967);
or U18501 (N_18501,N_17540,N_17775);
nand U18502 (N_18502,N_17768,N_17526);
nand U18503 (N_18503,N_17538,N_17531);
nor U18504 (N_18504,N_17509,N_18013);
nor U18505 (N_18505,N_17986,N_17932);
nand U18506 (N_18506,N_18044,N_17853);
xor U18507 (N_18507,N_17592,N_17859);
nor U18508 (N_18508,N_17947,N_17502);
or U18509 (N_18509,N_17920,N_17872);
xnor U18510 (N_18510,N_17755,N_17935);
nor U18511 (N_18511,N_17506,N_17754);
or U18512 (N_18512,N_17807,N_17681);
nor U18513 (N_18513,N_17580,N_17503);
nor U18514 (N_18514,N_17575,N_18097);
or U18515 (N_18515,N_17528,N_18086);
and U18516 (N_18516,N_17897,N_17787);
xor U18517 (N_18517,N_17597,N_17633);
nand U18518 (N_18518,N_17889,N_17625);
nand U18519 (N_18519,N_18060,N_18016);
xor U18520 (N_18520,N_17579,N_17506);
or U18521 (N_18521,N_17603,N_17716);
nand U18522 (N_18522,N_17724,N_17636);
and U18523 (N_18523,N_17681,N_17806);
nand U18524 (N_18524,N_17776,N_17767);
nor U18525 (N_18525,N_17513,N_18087);
nor U18526 (N_18526,N_17785,N_17888);
and U18527 (N_18527,N_17908,N_17920);
nor U18528 (N_18528,N_17518,N_17779);
xnor U18529 (N_18529,N_17551,N_17918);
nor U18530 (N_18530,N_17699,N_17636);
and U18531 (N_18531,N_17670,N_17857);
nand U18532 (N_18532,N_17832,N_17568);
nor U18533 (N_18533,N_17707,N_18110);
and U18534 (N_18534,N_17949,N_17850);
nand U18535 (N_18535,N_17774,N_18045);
nor U18536 (N_18536,N_18004,N_17633);
or U18537 (N_18537,N_17790,N_17924);
and U18538 (N_18538,N_17931,N_17766);
or U18539 (N_18539,N_18008,N_17899);
nand U18540 (N_18540,N_18076,N_18018);
nand U18541 (N_18541,N_18038,N_17777);
nand U18542 (N_18542,N_17955,N_17617);
xnor U18543 (N_18543,N_17803,N_17975);
or U18544 (N_18544,N_17525,N_17627);
or U18545 (N_18545,N_18015,N_17691);
nand U18546 (N_18546,N_17751,N_17507);
or U18547 (N_18547,N_17941,N_17678);
nand U18548 (N_18548,N_17748,N_17520);
nor U18549 (N_18549,N_18100,N_17909);
and U18550 (N_18550,N_18052,N_17593);
and U18551 (N_18551,N_18058,N_17505);
or U18552 (N_18552,N_17792,N_17530);
or U18553 (N_18553,N_18030,N_18114);
nand U18554 (N_18554,N_17662,N_18086);
nor U18555 (N_18555,N_17802,N_17863);
or U18556 (N_18556,N_17605,N_17520);
or U18557 (N_18557,N_17889,N_17548);
nor U18558 (N_18558,N_17579,N_17680);
nor U18559 (N_18559,N_17933,N_17742);
or U18560 (N_18560,N_17821,N_17646);
nand U18561 (N_18561,N_17929,N_18046);
and U18562 (N_18562,N_17559,N_17552);
or U18563 (N_18563,N_18013,N_17968);
or U18564 (N_18564,N_17634,N_17697);
and U18565 (N_18565,N_17751,N_17593);
xnor U18566 (N_18566,N_17858,N_17823);
nand U18567 (N_18567,N_17988,N_17586);
and U18568 (N_18568,N_18099,N_17674);
and U18569 (N_18569,N_17870,N_17843);
or U18570 (N_18570,N_18022,N_18041);
xnor U18571 (N_18571,N_17658,N_17834);
or U18572 (N_18572,N_17797,N_18038);
and U18573 (N_18573,N_17791,N_17742);
nor U18574 (N_18574,N_17644,N_17908);
nor U18575 (N_18575,N_17830,N_17667);
nand U18576 (N_18576,N_17655,N_17903);
nand U18577 (N_18577,N_17579,N_18045);
or U18578 (N_18578,N_17867,N_17732);
and U18579 (N_18579,N_17670,N_18079);
or U18580 (N_18580,N_17940,N_17560);
and U18581 (N_18581,N_17591,N_18063);
or U18582 (N_18582,N_17626,N_17515);
nand U18583 (N_18583,N_17706,N_17576);
and U18584 (N_18584,N_17539,N_17771);
or U18585 (N_18585,N_17801,N_17663);
xnor U18586 (N_18586,N_17618,N_17599);
and U18587 (N_18587,N_17986,N_18065);
and U18588 (N_18588,N_17927,N_17863);
or U18589 (N_18589,N_17772,N_17889);
or U18590 (N_18590,N_17505,N_18093);
nor U18591 (N_18591,N_17895,N_17874);
and U18592 (N_18592,N_17881,N_17908);
nor U18593 (N_18593,N_17848,N_18117);
or U18594 (N_18594,N_17663,N_17624);
nor U18595 (N_18595,N_17644,N_17506);
or U18596 (N_18596,N_18032,N_17995);
and U18597 (N_18597,N_17947,N_17825);
or U18598 (N_18598,N_17506,N_17610);
nor U18599 (N_18599,N_17588,N_17772);
nand U18600 (N_18600,N_17550,N_17604);
or U18601 (N_18601,N_17626,N_17896);
or U18602 (N_18602,N_17631,N_17595);
or U18603 (N_18603,N_17868,N_17714);
and U18604 (N_18604,N_17872,N_17550);
nand U18605 (N_18605,N_17708,N_18076);
nand U18606 (N_18606,N_17523,N_17605);
nand U18607 (N_18607,N_17621,N_17675);
or U18608 (N_18608,N_18088,N_17779);
or U18609 (N_18609,N_18069,N_17558);
xnor U18610 (N_18610,N_17638,N_17840);
or U18611 (N_18611,N_17656,N_17903);
nor U18612 (N_18612,N_17655,N_17904);
nand U18613 (N_18613,N_17514,N_17840);
or U18614 (N_18614,N_17881,N_17594);
or U18615 (N_18615,N_17831,N_17755);
xor U18616 (N_18616,N_17587,N_17581);
nor U18617 (N_18617,N_17693,N_17575);
and U18618 (N_18618,N_17831,N_17577);
nand U18619 (N_18619,N_17802,N_17561);
nor U18620 (N_18620,N_18014,N_18074);
and U18621 (N_18621,N_17507,N_17781);
and U18622 (N_18622,N_18108,N_18055);
nor U18623 (N_18623,N_18054,N_18098);
nand U18624 (N_18624,N_17914,N_17875);
and U18625 (N_18625,N_17642,N_18003);
nor U18626 (N_18626,N_17827,N_17798);
or U18627 (N_18627,N_18061,N_18014);
nor U18628 (N_18628,N_17795,N_17902);
nand U18629 (N_18629,N_18121,N_17754);
nand U18630 (N_18630,N_17939,N_18010);
and U18631 (N_18631,N_17798,N_17812);
nand U18632 (N_18632,N_18114,N_17970);
nand U18633 (N_18633,N_17650,N_17881);
nor U18634 (N_18634,N_17711,N_17725);
nor U18635 (N_18635,N_17647,N_17874);
xor U18636 (N_18636,N_17629,N_17546);
nand U18637 (N_18637,N_17639,N_17809);
nand U18638 (N_18638,N_18103,N_17593);
nor U18639 (N_18639,N_17828,N_17501);
nor U18640 (N_18640,N_18028,N_17737);
nand U18641 (N_18641,N_17649,N_17593);
nand U18642 (N_18642,N_17821,N_18061);
nor U18643 (N_18643,N_17977,N_17988);
nand U18644 (N_18644,N_17733,N_17540);
nor U18645 (N_18645,N_17945,N_17515);
and U18646 (N_18646,N_17658,N_17560);
nand U18647 (N_18647,N_17673,N_17530);
nor U18648 (N_18648,N_17646,N_18075);
nor U18649 (N_18649,N_17825,N_17655);
nand U18650 (N_18650,N_17559,N_17527);
or U18651 (N_18651,N_18072,N_18085);
nand U18652 (N_18652,N_17620,N_17804);
or U18653 (N_18653,N_17608,N_17597);
or U18654 (N_18654,N_17880,N_17693);
or U18655 (N_18655,N_17781,N_18051);
and U18656 (N_18656,N_17684,N_17947);
and U18657 (N_18657,N_17735,N_18010);
nor U18658 (N_18658,N_17943,N_17815);
and U18659 (N_18659,N_17872,N_17710);
or U18660 (N_18660,N_17986,N_17658);
or U18661 (N_18661,N_17860,N_17830);
and U18662 (N_18662,N_17745,N_18022);
nand U18663 (N_18663,N_17654,N_17669);
xor U18664 (N_18664,N_17820,N_17885);
nor U18665 (N_18665,N_18090,N_17937);
or U18666 (N_18666,N_17945,N_17514);
nand U18667 (N_18667,N_18054,N_18112);
or U18668 (N_18668,N_17848,N_17682);
xnor U18669 (N_18669,N_17757,N_18097);
xor U18670 (N_18670,N_18116,N_18050);
or U18671 (N_18671,N_17795,N_18004);
xnor U18672 (N_18672,N_17890,N_17626);
nand U18673 (N_18673,N_18013,N_17855);
nand U18674 (N_18674,N_17986,N_18113);
or U18675 (N_18675,N_17642,N_17558);
nor U18676 (N_18676,N_18032,N_18079);
and U18677 (N_18677,N_17840,N_18051);
and U18678 (N_18678,N_18028,N_17712);
xor U18679 (N_18679,N_17914,N_17923);
nor U18680 (N_18680,N_17649,N_17923);
nand U18681 (N_18681,N_17624,N_17904);
nor U18682 (N_18682,N_18080,N_17637);
nor U18683 (N_18683,N_17698,N_17618);
and U18684 (N_18684,N_17838,N_18079);
or U18685 (N_18685,N_17618,N_17753);
nand U18686 (N_18686,N_17981,N_18117);
nor U18687 (N_18687,N_17985,N_17992);
nor U18688 (N_18688,N_17667,N_18096);
or U18689 (N_18689,N_17633,N_17683);
and U18690 (N_18690,N_17864,N_17509);
or U18691 (N_18691,N_17724,N_17685);
and U18692 (N_18692,N_17671,N_17651);
nand U18693 (N_18693,N_17910,N_17980);
nand U18694 (N_18694,N_17771,N_17816);
nor U18695 (N_18695,N_17781,N_17568);
nand U18696 (N_18696,N_17954,N_17572);
and U18697 (N_18697,N_17769,N_17570);
xnor U18698 (N_18698,N_18105,N_17601);
nor U18699 (N_18699,N_18042,N_17540);
or U18700 (N_18700,N_18062,N_18073);
or U18701 (N_18701,N_17824,N_17583);
nand U18702 (N_18702,N_17662,N_17532);
and U18703 (N_18703,N_17606,N_18096);
and U18704 (N_18704,N_17952,N_17521);
nand U18705 (N_18705,N_17554,N_17808);
nand U18706 (N_18706,N_17995,N_17707);
and U18707 (N_18707,N_17935,N_17711);
and U18708 (N_18708,N_17927,N_17978);
nor U18709 (N_18709,N_17883,N_17892);
nand U18710 (N_18710,N_17806,N_17608);
and U18711 (N_18711,N_17774,N_17963);
nor U18712 (N_18712,N_18070,N_17970);
or U18713 (N_18713,N_17665,N_17945);
or U18714 (N_18714,N_17621,N_17705);
nand U18715 (N_18715,N_17649,N_17912);
nor U18716 (N_18716,N_17792,N_17551);
nor U18717 (N_18717,N_17819,N_17555);
or U18718 (N_18718,N_17922,N_17505);
nand U18719 (N_18719,N_17824,N_17648);
xnor U18720 (N_18720,N_17702,N_17604);
nor U18721 (N_18721,N_17957,N_17583);
xnor U18722 (N_18722,N_17799,N_17582);
xor U18723 (N_18723,N_17608,N_17925);
nor U18724 (N_18724,N_18067,N_17502);
and U18725 (N_18725,N_18087,N_17572);
or U18726 (N_18726,N_17675,N_17604);
xor U18727 (N_18727,N_17616,N_17846);
or U18728 (N_18728,N_17817,N_17557);
and U18729 (N_18729,N_18031,N_17576);
nand U18730 (N_18730,N_18044,N_17775);
and U18731 (N_18731,N_17946,N_17990);
and U18732 (N_18732,N_17822,N_17654);
and U18733 (N_18733,N_17517,N_17882);
or U18734 (N_18734,N_17724,N_17526);
or U18735 (N_18735,N_17525,N_17973);
or U18736 (N_18736,N_17594,N_18107);
xnor U18737 (N_18737,N_17935,N_17747);
nand U18738 (N_18738,N_17787,N_17623);
nand U18739 (N_18739,N_17984,N_17500);
nor U18740 (N_18740,N_17652,N_17956);
nor U18741 (N_18741,N_18106,N_17839);
xnor U18742 (N_18742,N_18109,N_17544);
nand U18743 (N_18743,N_17530,N_17707);
or U18744 (N_18744,N_17852,N_17552);
nor U18745 (N_18745,N_18122,N_17930);
and U18746 (N_18746,N_17568,N_17739);
and U18747 (N_18747,N_18074,N_17651);
nor U18748 (N_18748,N_17822,N_17639);
xor U18749 (N_18749,N_18094,N_17833);
or U18750 (N_18750,N_18582,N_18173);
and U18751 (N_18751,N_18509,N_18706);
or U18752 (N_18752,N_18231,N_18278);
and U18753 (N_18753,N_18674,N_18483);
nor U18754 (N_18754,N_18647,N_18634);
or U18755 (N_18755,N_18283,N_18346);
nor U18756 (N_18756,N_18748,N_18485);
and U18757 (N_18757,N_18540,N_18343);
and U18758 (N_18758,N_18664,N_18377);
or U18759 (N_18759,N_18251,N_18630);
and U18760 (N_18760,N_18252,N_18613);
and U18761 (N_18761,N_18361,N_18450);
and U18762 (N_18762,N_18274,N_18288);
nor U18763 (N_18763,N_18736,N_18575);
and U18764 (N_18764,N_18516,N_18682);
nand U18765 (N_18765,N_18280,N_18461);
nor U18766 (N_18766,N_18224,N_18271);
or U18767 (N_18767,N_18368,N_18693);
xnor U18768 (N_18768,N_18642,N_18220);
or U18769 (N_18769,N_18621,N_18718);
nor U18770 (N_18770,N_18431,N_18383);
or U18771 (N_18771,N_18667,N_18260);
or U18772 (N_18772,N_18716,N_18386);
xnor U18773 (N_18773,N_18728,N_18448);
or U18774 (N_18774,N_18396,N_18645);
xor U18775 (N_18775,N_18465,N_18519);
or U18776 (N_18776,N_18671,N_18347);
and U18777 (N_18777,N_18189,N_18155);
and U18778 (N_18778,N_18496,N_18282);
and U18779 (N_18779,N_18458,N_18417);
nand U18780 (N_18780,N_18545,N_18380);
xor U18781 (N_18781,N_18734,N_18363);
and U18782 (N_18782,N_18565,N_18602);
or U18783 (N_18783,N_18619,N_18307);
nand U18784 (N_18784,N_18241,N_18385);
or U18785 (N_18785,N_18196,N_18273);
and U18786 (N_18786,N_18709,N_18354);
nor U18787 (N_18787,N_18317,N_18356);
nor U18788 (N_18788,N_18321,N_18256);
nand U18789 (N_18789,N_18344,N_18358);
nand U18790 (N_18790,N_18585,N_18410);
nand U18791 (N_18791,N_18408,N_18503);
nand U18792 (N_18792,N_18146,N_18434);
nand U18793 (N_18793,N_18133,N_18436);
xor U18794 (N_18794,N_18330,N_18334);
or U18795 (N_18795,N_18319,N_18167);
nand U18796 (N_18796,N_18699,N_18250);
or U18797 (N_18797,N_18400,N_18232);
or U18798 (N_18798,N_18178,N_18229);
or U18799 (N_18799,N_18429,N_18290);
nand U18800 (N_18800,N_18394,N_18524);
nor U18801 (N_18801,N_18745,N_18275);
and U18802 (N_18802,N_18158,N_18180);
nand U18803 (N_18803,N_18705,N_18292);
nor U18804 (N_18804,N_18309,N_18562);
and U18805 (N_18805,N_18299,N_18494);
nor U18806 (N_18806,N_18353,N_18153);
nor U18807 (N_18807,N_18481,N_18639);
nor U18808 (N_18808,N_18176,N_18614);
nand U18809 (N_18809,N_18201,N_18515);
and U18810 (N_18810,N_18217,N_18659);
or U18811 (N_18811,N_18154,N_18142);
and U18812 (N_18812,N_18574,N_18175);
and U18813 (N_18813,N_18308,N_18744);
xnor U18814 (N_18814,N_18533,N_18596);
nor U18815 (N_18815,N_18402,N_18738);
nand U18816 (N_18816,N_18650,N_18589);
or U18817 (N_18817,N_18723,N_18199);
nand U18818 (N_18818,N_18156,N_18473);
and U18819 (N_18819,N_18631,N_18187);
nor U18820 (N_18820,N_18493,N_18542);
nand U18821 (N_18821,N_18277,N_18507);
nor U18822 (N_18822,N_18610,N_18471);
or U18823 (N_18823,N_18612,N_18710);
or U18824 (N_18824,N_18295,N_18336);
and U18825 (N_18825,N_18214,N_18615);
or U18826 (N_18826,N_18412,N_18580);
xor U18827 (N_18827,N_18703,N_18419);
nor U18828 (N_18828,N_18409,N_18502);
nor U18829 (N_18829,N_18457,N_18676);
and U18830 (N_18830,N_18418,N_18237);
or U18831 (N_18831,N_18428,N_18677);
xor U18832 (N_18832,N_18238,N_18543);
nand U18833 (N_18833,N_18143,N_18658);
nand U18834 (N_18834,N_18670,N_18310);
or U18835 (N_18835,N_18648,N_18666);
nand U18836 (N_18836,N_18351,N_18495);
nand U18837 (N_18837,N_18576,N_18573);
nand U18838 (N_18838,N_18510,N_18269);
nor U18839 (N_18839,N_18215,N_18695);
or U18840 (N_18840,N_18297,N_18242);
and U18841 (N_18841,N_18160,N_18643);
nand U18842 (N_18842,N_18475,N_18314);
or U18843 (N_18843,N_18595,N_18304);
and U18844 (N_18844,N_18328,N_18726);
nor U18845 (N_18845,N_18372,N_18511);
nor U18846 (N_18846,N_18590,N_18253);
or U18847 (N_18847,N_18629,N_18443);
nand U18848 (N_18848,N_18255,N_18732);
nor U18849 (N_18849,N_18512,N_18139);
xor U18850 (N_18850,N_18185,N_18239);
and U18851 (N_18851,N_18742,N_18287);
nand U18852 (N_18852,N_18460,N_18374);
xor U18853 (N_18853,N_18130,N_18147);
nor U18854 (N_18854,N_18478,N_18668);
or U18855 (N_18855,N_18535,N_18449);
nor U18856 (N_18856,N_18636,N_18192);
and U18857 (N_18857,N_18135,N_18479);
or U18858 (N_18858,N_18195,N_18737);
and U18859 (N_18859,N_18568,N_18561);
and U18860 (N_18860,N_18714,N_18451);
and U18861 (N_18861,N_18704,N_18349);
xnor U18862 (N_18862,N_18379,N_18741);
nor U18863 (N_18863,N_18365,N_18675);
xnor U18864 (N_18864,N_18456,N_18236);
nand U18865 (N_18865,N_18712,N_18414);
and U18866 (N_18866,N_18708,N_18687);
nand U18867 (N_18867,N_18541,N_18322);
nor U18868 (N_18868,N_18184,N_18247);
and U18869 (N_18869,N_18174,N_18551);
or U18870 (N_18870,N_18606,N_18504);
nand U18871 (N_18871,N_18729,N_18286);
nand U18872 (N_18872,N_18134,N_18508);
and U18873 (N_18873,N_18598,N_18455);
or U18874 (N_18874,N_18702,N_18454);
and U18875 (N_18875,N_18244,N_18222);
nand U18876 (N_18876,N_18207,N_18392);
nand U18877 (N_18877,N_18165,N_18149);
nand U18878 (N_18878,N_18550,N_18583);
or U18879 (N_18879,N_18326,N_18557);
or U18880 (N_18880,N_18416,N_18554);
nand U18881 (N_18881,N_18381,N_18259);
nand U18882 (N_18882,N_18168,N_18216);
nand U18883 (N_18883,N_18513,N_18281);
or U18884 (N_18884,N_18452,N_18388);
and U18885 (N_18885,N_18616,N_18506);
and U18886 (N_18886,N_18657,N_18268);
nor U18887 (N_18887,N_18679,N_18691);
xor U18888 (N_18888,N_18638,N_18469);
and U18889 (N_18889,N_18532,N_18164);
and U18890 (N_18890,N_18663,N_18651);
nand U18891 (N_18891,N_18673,N_18713);
nor U18892 (N_18892,N_18206,N_18570);
or U18893 (N_18893,N_18571,N_18186);
nor U18894 (N_18894,N_18652,N_18246);
nand U18895 (N_18895,N_18422,N_18411);
or U18896 (N_18896,N_18291,N_18492);
nor U18897 (N_18897,N_18624,N_18538);
and U18898 (N_18898,N_18161,N_18254);
nand U18899 (N_18899,N_18440,N_18279);
or U18900 (N_18900,N_18625,N_18618);
and U18901 (N_18901,N_18592,N_18749);
nand U18902 (N_18902,N_18521,N_18727);
nor U18903 (N_18903,N_18453,N_18403);
or U18904 (N_18904,N_18267,N_18528);
nand U18905 (N_18905,N_18438,N_18439);
and U18906 (N_18906,N_18644,N_18371);
nand U18907 (N_18907,N_18669,N_18531);
nor U18908 (N_18908,N_18566,N_18219);
nand U18909 (N_18909,N_18484,N_18662);
and U18910 (N_18910,N_18633,N_18132);
nand U18911 (N_18911,N_18743,N_18205);
and U18912 (N_18912,N_18325,N_18293);
or U18913 (N_18913,N_18415,N_18261);
or U18914 (N_18914,N_18405,N_18223);
xor U18915 (N_18915,N_18157,N_18637);
or U18916 (N_18916,N_18315,N_18337);
nand U18917 (N_18917,N_18477,N_18359);
nor U18918 (N_18918,N_18686,N_18387);
and U18919 (N_18919,N_18721,N_18193);
nor U18920 (N_18920,N_18746,N_18678);
and U18921 (N_18921,N_18498,N_18563);
and U18922 (N_18922,N_18225,N_18525);
nor U18923 (N_18923,N_18649,N_18435);
or U18924 (N_18924,N_18620,N_18311);
nand U18925 (N_18925,N_18560,N_18426);
nand U18926 (N_18926,N_18382,N_18144);
nor U18927 (N_18927,N_18437,N_18301);
or U18928 (N_18928,N_18198,N_18127);
nand U18929 (N_18929,N_18601,N_18316);
nand U18930 (N_18930,N_18430,N_18378);
or U18931 (N_18931,N_18213,N_18169);
or U18932 (N_18932,N_18586,N_18536);
or U18933 (N_18933,N_18623,N_18672);
nor U18934 (N_18934,N_18424,N_18318);
nand U18935 (N_18935,N_18302,N_18162);
or U18936 (N_18936,N_18406,N_18298);
nor U18937 (N_18937,N_18427,N_18526);
and U18938 (N_18938,N_18480,N_18170);
xor U18939 (N_18939,N_18603,N_18534);
and U18940 (N_18940,N_18725,N_18505);
or U18941 (N_18941,N_18499,N_18599);
nand U18942 (N_18942,N_18514,N_18593);
and U18943 (N_18943,N_18235,N_18497);
nand U18944 (N_18944,N_18464,N_18537);
and U18945 (N_18945,N_18635,N_18445);
or U18946 (N_18946,N_18722,N_18587);
nor U18947 (N_18947,N_18628,N_18681);
nand U18948 (N_18948,N_18689,N_18553);
xnor U18949 (N_18949,N_18398,N_18352);
or U18950 (N_18950,N_18569,N_18640);
nor U18951 (N_18951,N_18257,N_18204);
or U18952 (N_18952,N_18605,N_18501);
and U18953 (N_18953,N_18350,N_18329);
xnor U18954 (N_18954,N_18340,N_18547);
xor U18955 (N_18955,N_18357,N_18463);
nand U18956 (N_18956,N_18539,N_18183);
or U18957 (N_18957,N_18369,N_18468);
and U18958 (N_18958,N_18303,N_18230);
and U18959 (N_18959,N_18611,N_18730);
and U18960 (N_18960,N_18470,N_18572);
nor U18961 (N_18961,N_18420,N_18720);
or U18962 (N_18962,N_18622,N_18202);
nand U18963 (N_18963,N_18366,N_18240);
and U18964 (N_18964,N_18700,N_18641);
and U18965 (N_18965,N_18270,N_18320);
nor U18966 (N_18966,N_18362,N_18442);
nor U18967 (N_18967,N_18735,N_18444);
and U18968 (N_18968,N_18128,N_18653);
or U18969 (N_18969,N_18433,N_18399);
and U18970 (N_18970,N_18129,N_18276);
or U18971 (N_18971,N_18548,N_18384);
nand U18972 (N_18972,N_18530,N_18740);
and U18973 (N_18973,N_18243,N_18393);
and U18974 (N_18974,N_18266,N_18182);
or U18975 (N_18975,N_18367,N_18552);
xor U18976 (N_18976,N_18264,N_18306);
or U18977 (N_18977,N_18421,N_18577);
or U18978 (N_18978,N_18375,N_18476);
or U18979 (N_18979,N_18262,N_18467);
or U18980 (N_18980,N_18459,N_18294);
nor U18981 (N_18981,N_18159,N_18660);
xnor U18982 (N_18982,N_18285,N_18263);
or U18983 (N_18983,N_18345,N_18627);
nor U18984 (N_18984,N_18177,N_18342);
and U18985 (N_18985,N_18698,N_18209);
or U18986 (N_18986,N_18441,N_18701);
nor U18987 (N_18987,N_18523,N_18407);
nor U18988 (N_18988,N_18685,N_18690);
nand U18989 (N_18989,N_18594,N_18338);
and U18990 (N_18990,N_18172,N_18697);
nand U18991 (N_18991,N_18212,N_18210);
and U18992 (N_18992,N_18323,N_18688);
nor U18993 (N_18993,N_18446,N_18696);
or U18994 (N_18994,N_18683,N_18425);
and U18995 (N_18995,N_18607,N_18137);
nor U18996 (N_18996,N_18188,N_18360);
nand U18997 (N_18997,N_18684,N_18739);
or U18998 (N_18998,N_18151,N_18488);
and U18999 (N_18999,N_18138,N_18556);
and U19000 (N_19000,N_18482,N_18715);
nor U19001 (N_19001,N_18474,N_18227);
and U19002 (N_19002,N_18131,N_18284);
and U19003 (N_19003,N_18401,N_18194);
and U19004 (N_19004,N_18233,N_18218);
and U19005 (N_19005,N_18355,N_18339);
nand U19006 (N_19006,N_18272,N_18717);
nor U19007 (N_19007,N_18567,N_18517);
or U19008 (N_19008,N_18376,N_18707);
or U19009 (N_19009,N_18564,N_18208);
and U19010 (N_19010,N_18163,N_18462);
nand U19011 (N_19011,N_18141,N_18520);
or U19012 (N_19012,N_18265,N_18711);
xor U19013 (N_19013,N_18617,N_18348);
xnor U19014 (N_19014,N_18609,N_18680);
nand U19015 (N_19015,N_18692,N_18312);
nor U19016 (N_19016,N_18486,N_18136);
nor U19017 (N_19017,N_18370,N_18518);
nor U19018 (N_19018,N_18390,N_18608);
or U19019 (N_19019,N_18190,N_18364);
nor U19020 (N_19020,N_18581,N_18656);
or U19021 (N_19021,N_18203,N_18211);
and U19022 (N_19022,N_18733,N_18221);
nor U19023 (N_19023,N_18588,N_18335);
and U19024 (N_19024,N_18171,N_18591);
nand U19025 (N_19025,N_18179,N_18491);
nor U19026 (N_19026,N_18489,N_18305);
or U19027 (N_19027,N_18719,N_18258);
xor U19028 (N_19028,N_18604,N_18432);
nand U19029 (N_19029,N_18145,N_18397);
and U19030 (N_19030,N_18500,N_18584);
nand U19031 (N_19031,N_18166,N_18395);
nor U19032 (N_19032,N_18200,N_18391);
or U19033 (N_19033,N_18125,N_18327);
or U19034 (N_19034,N_18333,N_18447);
or U19035 (N_19035,N_18423,N_18626);
nand U19036 (N_19036,N_18373,N_18296);
nor U19037 (N_19037,N_18152,N_18245);
and U19038 (N_19038,N_18555,N_18661);
nor U19039 (N_19039,N_18527,N_18731);
nand U19040 (N_19040,N_18597,N_18490);
or U19041 (N_19041,N_18466,N_18228);
nor U19042 (N_19042,N_18234,N_18546);
nor U19043 (N_19043,N_18646,N_18558);
and U19044 (N_19044,N_18191,N_18140);
and U19045 (N_19045,N_18300,N_18150);
and U19046 (N_19046,N_18578,N_18579);
nand U19047 (N_19047,N_18197,N_18313);
nor U19048 (N_19048,N_18529,N_18181);
nand U19049 (N_19049,N_18331,N_18487);
or U19050 (N_19050,N_18724,N_18289);
nand U19051 (N_19051,N_18549,N_18249);
or U19052 (N_19052,N_18654,N_18655);
or U19053 (N_19053,N_18324,N_18472);
and U19054 (N_19054,N_18413,N_18694);
nor U19055 (N_19055,N_18600,N_18665);
xnor U19056 (N_19056,N_18148,N_18522);
nand U19057 (N_19057,N_18404,N_18559);
nand U19058 (N_19058,N_18226,N_18389);
nor U19059 (N_19059,N_18126,N_18747);
or U19060 (N_19060,N_18332,N_18341);
or U19061 (N_19061,N_18632,N_18248);
nand U19062 (N_19062,N_18544,N_18469);
and U19063 (N_19063,N_18194,N_18632);
or U19064 (N_19064,N_18484,N_18531);
and U19065 (N_19065,N_18324,N_18153);
and U19066 (N_19066,N_18591,N_18326);
and U19067 (N_19067,N_18168,N_18219);
nor U19068 (N_19068,N_18204,N_18450);
nor U19069 (N_19069,N_18434,N_18542);
nand U19070 (N_19070,N_18683,N_18198);
xor U19071 (N_19071,N_18249,N_18689);
nand U19072 (N_19072,N_18180,N_18681);
nand U19073 (N_19073,N_18308,N_18483);
xnor U19074 (N_19074,N_18588,N_18441);
nand U19075 (N_19075,N_18516,N_18603);
nor U19076 (N_19076,N_18225,N_18552);
nor U19077 (N_19077,N_18654,N_18579);
or U19078 (N_19078,N_18457,N_18499);
or U19079 (N_19079,N_18600,N_18291);
and U19080 (N_19080,N_18318,N_18279);
nor U19081 (N_19081,N_18376,N_18354);
and U19082 (N_19082,N_18343,N_18516);
nor U19083 (N_19083,N_18166,N_18341);
nor U19084 (N_19084,N_18415,N_18231);
and U19085 (N_19085,N_18449,N_18629);
nand U19086 (N_19086,N_18748,N_18649);
or U19087 (N_19087,N_18318,N_18464);
or U19088 (N_19088,N_18225,N_18411);
and U19089 (N_19089,N_18484,N_18369);
and U19090 (N_19090,N_18186,N_18323);
or U19091 (N_19091,N_18447,N_18551);
or U19092 (N_19092,N_18137,N_18588);
nor U19093 (N_19093,N_18421,N_18320);
nand U19094 (N_19094,N_18390,N_18148);
and U19095 (N_19095,N_18455,N_18651);
nand U19096 (N_19096,N_18405,N_18301);
and U19097 (N_19097,N_18579,N_18550);
or U19098 (N_19098,N_18398,N_18381);
nor U19099 (N_19099,N_18321,N_18601);
nor U19100 (N_19100,N_18665,N_18173);
and U19101 (N_19101,N_18464,N_18161);
xor U19102 (N_19102,N_18628,N_18531);
nor U19103 (N_19103,N_18577,N_18303);
xnor U19104 (N_19104,N_18186,N_18474);
and U19105 (N_19105,N_18591,N_18725);
nor U19106 (N_19106,N_18231,N_18445);
nand U19107 (N_19107,N_18536,N_18684);
and U19108 (N_19108,N_18715,N_18367);
nor U19109 (N_19109,N_18675,N_18236);
or U19110 (N_19110,N_18641,N_18741);
or U19111 (N_19111,N_18739,N_18416);
or U19112 (N_19112,N_18554,N_18144);
nor U19113 (N_19113,N_18746,N_18570);
or U19114 (N_19114,N_18656,N_18665);
and U19115 (N_19115,N_18142,N_18471);
and U19116 (N_19116,N_18290,N_18298);
nand U19117 (N_19117,N_18392,N_18251);
nor U19118 (N_19118,N_18616,N_18704);
or U19119 (N_19119,N_18626,N_18253);
nor U19120 (N_19120,N_18593,N_18503);
and U19121 (N_19121,N_18167,N_18632);
nor U19122 (N_19122,N_18321,N_18397);
nand U19123 (N_19123,N_18674,N_18621);
or U19124 (N_19124,N_18306,N_18247);
nor U19125 (N_19125,N_18340,N_18303);
and U19126 (N_19126,N_18495,N_18188);
and U19127 (N_19127,N_18580,N_18667);
or U19128 (N_19128,N_18349,N_18507);
nand U19129 (N_19129,N_18197,N_18247);
nor U19130 (N_19130,N_18297,N_18509);
nor U19131 (N_19131,N_18665,N_18215);
nor U19132 (N_19132,N_18519,N_18339);
nor U19133 (N_19133,N_18178,N_18184);
nand U19134 (N_19134,N_18202,N_18522);
or U19135 (N_19135,N_18239,N_18658);
or U19136 (N_19136,N_18308,N_18160);
or U19137 (N_19137,N_18258,N_18298);
nand U19138 (N_19138,N_18193,N_18617);
and U19139 (N_19139,N_18496,N_18386);
nor U19140 (N_19140,N_18171,N_18246);
nor U19141 (N_19141,N_18161,N_18437);
and U19142 (N_19142,N_18531,N_18549);
and U19143 (N_19143,N_18704,N_18677);
nor U19144 (N_19144,N_18517,N_18315);
nor U19145 (N_19145,N_18154,N_18293);
and U19146 (N_19146,N_18550,N_18308);
xor U19147 (N_19147,N_18192,N_18350);
nand U19148 (N_19148,N_18721,N_18236);
and U19149 (N_19149,N_18211,N_18503);
or U19150 (N_19150,N_18182,N_18412);
and U19151 (N_19151,N_18219,N_18297);
and U19152 (N_19152,N_18746,N_18274);
and U19153 (N_19153,N_18156,N_18219);
nand U19154 (N_19154,N_18652,N_18423);
or U19155 (N_19155,N_18489,N_18662);
or U19156 (N_19156,N_18589,N_18625);
nor U19157 (N_19157,N_18137,N_18508);
and U19158 (N_19158,N_18137,N_18171);
and U19159 (N_19159,N_18250,N_18599);
and U19160 (N_19160,N_18632,N_18386);
nand U19161 (N_19161,N_18478,N_18481);
nor U19162 (N_19162,N_18567,N_18535);
nor U19163 (N_19163,N_18385,N_18552);
nor U19164 (N_19164,N_18219,N_18611);
and U19165 (N_19165,N_18506,N_18560);
nor U19166 (N_19166,N_18284,N_18472);
xor U19167 (N_19167,N_18448,N_18186);
nor U19168 (N_19168,N_18687,N_18590);
nand U19169 (N_19169,N_18170,N_18273);
or U19170 (N_19170,N_18234,N_18606);
xnor U19171 (N_19171,N_18648,N_18458);
xnor U19172 (N_19172,N_18559,N_18434);
nor U19173 (N_19173,N_18410,N_18704);
xor U19174 (N_19174,N_18226,N_18692);
nor U19175 (N_19175,N_18426,N_18156);
nand U19176 (N_19176,N_18192,N_18384);
xnor U19177 (N_19177,N_18708,N_18343);
or U19178 (N_19178,N_18544,N_18437);
and U19179 (N_19179,N_18615,N_18313);
xnor U19180 (N_19180,N_18147,N_18478);
and U19181 (N_19181,N_18363,N_18246);
nor U19182 (N_19182,N_18494,N_18207);
or U19183 (N_19183,N_18453,N_18149);
nor U19184 (N_19184,N_18582,N_18558);
or U19185 (N_19185,N_18217,N_18294);
xor U19186 (N_19186,N_18538,N_18477);
nand U19187 (N_19187,N_18514,N_18359);
or U19188 (N_19188,N_18480,N_18462);
or U19189 (N_19189,N_18727,N_18346);
or U19190 (N_19190,N_18321,N_18685);
and U19191 (N_19191,N_18530,N_18711);
or U19192 (N_19192,N_18535,N_18668);
nor U19193 (N_19193,N_18435,N_18686);
nand U19194 (N_19194,N_18744,N_18204);
nor U19195 (N_19195,N_18507,N_18138);
and U19196 (N_19196,N_18180,N_18659);
or U19197 (N_19197,N_18318,N_18218);
nand U19198 (N_19198,N_18342,N_18348);
nor U19199 (N_19199,N_18741,N_18586);
nor U19200 (N_19200,N_18482,N_18532);
nor U19201 (N_19201,N_18712,N_18399);
and U19202 (N_19202,N_18563,N_18668);
nor U19203 (N_19203,N_18136,N_18577);
xnor U19204 (N_19204,N_18231,N_18572);
or U19205 (N_19205,N_18333,N_18564);
nand U19206 (N_19206,N_18172,N_18605);
nand U19207 (N_19207,N_18627,N_18309);
and U19208 (N_19208,N_18152,N_18204);
and U19209 (N_19209,N_18674,N_18658);
nor U19210 (N_19210,N_18215,N_18635);
or U19211 (N_19211,N_18419,N_18475);
or U19212 (N_19212,N_18738,N_18732);
xnor U19213 (N_19213,N_18393,N_18513);
and U19214 (N_19214,N_18165,N_18196);
nand U19215 (N_19215,N_18708,N_18373);
xnor U19216 (N_19216,N_18699,N_18493);
and U19217 (N_19217,N_18587,N_18566);
and U19218 (N_19218,N_18455,N_18224);
nor U19219 (N_19219,N_18226,N_18738);
or U19220 (N_19220,N_18615,N_18476);
nor U19221 (N_19221,N_18474,N_18241);
nand U19222 (N_19222,N_18367,N_18214);
xor U19223 (N_19223,N_18608,N_18262);
nor U19224 (N_19224,N_18626,N_18168);
xnor U19225 (N_19225,N_18382,N_18452);
xor U19226 (N_19226,N_18237,N_18260);
nor U19227 (N_19227,N_18241,N_18576);
nor U19228 (N_19228,N_18149,N_18407);
or U19229 (N_19229,N_18462,N_18229);
or U19230 (N_19230,N_18423,N_18560);
nor U19231 (N_19231,N_18722,N_18337);
nand U19232 (N_19232,N_18266,N_18276);
nor U19233 (N_19233,N_18528,N_18690);
nor U19234 (N_19234,N_18297,N_18195);
xor U19235 (N_19235,N_18163,N_18322);
nor U19236 (N_19236,N_18128,N_18481);
xnor U19237 (N_19237,N_18351,N_18336);
nor U19238 (N_19238,N_18607,N_18390);
nand U19239 (N_19239,N_18618,N_18279);
nand U19240 (N_19240,N_18647,N_18670);
xnor U19241 (N_19241,N_18389,N_18732);
xnor U19242 (N_19242,N_18422,N_18554);
nor U19243 (N_19243,N_18550,N_18370);
nor U19244 (N_19244,N_18196,N_18296);
nor U19245 (N_19245,N_18138,N_18325);
and U19246 (N_19246,N_18267,N_18243);
nand U19247 (N_19247,N_18421,N_18209);
or U19248 (N_19248,N_18238,N_18295);
and U19249 (N_19249,N_18635,N_18678);
nor U19250 (N_19250,N_18445,N_18466);
nand U19251 (N_19251,N_18533,N_18563);
nand U19252 (N_19252,N_18464,N_18621);
and U19253 (N_19253,N_18133,N_18163);
nor U19254 (N_19254,N_18706,N_18410);
nand U19255 (N_19255,N_18229,N_18364);
nor U19256 (N_19256,N_18370,N_18681);
xor U19257 (N_19257,N_18502,N_18195);
or U19258 (N_19258,N_18509,N_18558);
nand U19259 (N_19259,N_18492,N_18225);
and U19260 (N_19260,N_18568,N_18276);
nand U19261 (N_19261,N_18224,N_18693);
nor U19262 (N_19262,N_18448,N_18262);
and U19263 (N_19263,N_18490,N_18445);
or U19264 (N_19264,N_18642,N_18441);
and U19265 (N_19265,N_18461,N_18414);
nand U19266 (N_19266,N_18147,N_18465);
or U19267 (N_19267,N_18442,N_18136);
or U19268 (N_19268,N_18244,N_18613);
and U19269 (N_19269,N_18235,N_18635);
or U19270 (N_19270,N_18250,N_18658);
nand U19271 (N_19271,N_18438,N_18375);
nand U19272 (N_19272,N_18153,N_18699);
nor U19273 (N_19273,N_18601,N_18481);
nor U19274 (N_19274,N_18647,N_18632);
and U19275 (N_19275,N_18701,N_18475);
and U19276 (N_19276,N_18591,N_18181);
or U19277 (N_19277,N_18546,N_18155);
and U19278 (N_19278,N_18581,N_18576);
nor U19279 (N_19279,N_18443,N_18199);
nor U19280 (N_19280,N_18341,N_18210);
and U19281 (N_19281,N_18450,N_18183);
and U19282 (N_19282,N_18705,N_18230);
nor U19283 (N_19283,N_18150,N_18584);
xnor U19284 (N_19284,N_18234,N_18598);
nor U19285 (N_19285,N_18231,N_18455);
or U19286 (N_19286,N_18182,N_18373);
or U19287 (N_19287,N_18190,N_18709);
and U19288 (N_19288,N_18597,N_18639);
nand U19289 (N_19289,N_18527,N_18518);
and U19290 (N_19290,N_18441,N_18186);
or U19291 (N_19291,N_18516,N_18365);
and U19292 (N_19292,N_18551,N_18372);
nand U19293 (N_19293,N_18273,N_18690);
nand U19294 (N_19294,N_18241,N_18378);
or U19295 (N_19295,N_18631,N_18715);
nor U19296 (N_19296,N_18233,N_18655);
nor U19297 (N_19297,N_18488,N_18149);
nand U19298 (N_19298,N_18419,N_18537);
nand U19299 (N_19299,N_18532,N_18620);
or U19300 (N_19300,N_18634,N_18274);
xor U19301 (N_19301,N_18163,N_18349);
nor U19302 (N_19302,N_18708,N_18527);
nor U19303 (N_19303,N_18644,N_18612);
or U19304 (N_19304,N_18256,N_18741);
xor U19305 (N_19305,N_18321,N_18233);
nor U19306 (N_19306,N_18238,N_18621);
nor U19307 (N_19307,N_18394,N_18506);
nand U19308 (N_19308,N_18207,N_18234);
nand U19309 (N_19309,N_18410,N_18571);
nor U19310 (N_19310,N_18443,N_18483);
nor U19311 (N_19311,N_18638,N_18537);
nand U19312 (N_19312,N_18407,N_18211);
or U19313 (N_19313,N_18722,N_18232);
xor U19314 (N_19314,N_18634,N_18289);
or U19315 (N_19315,N_18632,N_18200);
xnor U19316 (N_19316,N_18671,N_18484);
xor U19317 (N_19317,N_18328,N_18674);
xnor U19318 (N_19318,N_18445,N_18566);
and U19319 (N_19319,N_18169,N_18483);
or U19320 (N_19320,N_18579,N_18747);
and U19321 (N_19321,N_18673,N_18456);
or U19322 (N_19322,N_18150,N_18424);
or U19323 (N_19323,N_18464,N_18374);
nor U19324 (N_19324,N_18305,N_18641);
or U19325 (N_19325,N_18415,N_18283);
or U19326 (N_19326,N_18478,N_18448);
nand U19327 (N_19327,N_18572,N_18243);
nor U19328 (N_19328,N_18533,N_18395);
or U19329 (N_19329,N_18281,N_18715);
xor U19330 (N_19330,N_18166,N_18508);
xnor U19331 (N_19331,N_18295,N_18204);
and U19332 (N_19332,N_18522,N_18608);
or U19333 (N_19333,N_18345,N_18472);
or U19334 (N_19334,N_18265,N_18211);
or U19335 (N_19335,N_18411,N_18715);
nor U19336 (N_19336,N_18585,N_18228);
or U19337 (N_19337,N_18416,N_18312);
and U19338 (N_19338,N_18570,N_18536);
and U19339 (N_19339,N_18255,N_18209);
nor U19340 (N_19340,N_18171,N_18445);
or U19341 (N_19341,N_18705,N_18713);
or U19342 (N_19342,N_18125,N_18357);
nor U19343 (N_19343,N_18264,N_18136);
and U19344 (N_19344,N_18188,N_18542);
nand U19345 (N_19345,N_18373,N_18143);
or U19346 (N_19346,N_18316,N_18391);
and U19347 (N_19347,N_18525,N_18145);
and U19348 (N_19348,N_18302,N_18307);
nand U19349 (N_19349,N_18584,N_18499);
and U19350 (N_19350,N_18718,N_18680);
nor U19351 (N_19351,N_18438,N_18416);
nor U19352 (N_19352,N_18441,N_18584);
nand U19353 (N_19353,N_18639,N_18416);
and U19354 (N_19354,N_18746,N_18721);
nand U19355 (N_19355,N_18144,N_18546);
nor U19356 (N_19356,N_18358,N_18209);
or U19357 (N_19357,N_18438,N_18566);
and U19358 (N_19358,N_18203,N_18147);
nand U19359 (N_19359,N_18635,N_18397);
nor U19360 (N_19360,N_18692,N_18470);
xnor U19361 (N_19361,N_18287,N_18682);
xor U19362 (N_19362,N_18628,N_18659);
nand U19363 (N_19363,N_18553,N_18389);
nand U19364 (N_19364,N_18262,N_18380);
and U19365 (N_19365,N_18611,N_18201);
nand U19366 (N_19366,N_18394,N_18654);
or U19367 (N_19367,N_18254,N_18677);
nor U19368 (N_19368,N_18462,N_18630);
nand U19369 (N_19369,N_18578,N_18480);
nor U19370 (N_19370,N_18497,N_18617);
xnor U19371 (N_19371,N_18512,N_18703);
nor U19372 (N_19372,N_18345,N_18636);
or U19373 (N_19373,N_18266,N_18454);
xnor U19374 (N_19374,N_18652,N_18344);
nor U19375 (N_19375,N_18875,N_18814);
and U19376 (N_19376,N_19192,N_19314);
nand U19377 (N_19377,N_19270,N_19305);
nor U19378 (N_19378,N_19140,N_18937);
or U19379 (N_19379,N_19208,N_19260);
nand U19380 (N_19380,N_18780,N_19173);
and U19381 (N_19381,N_19363,N_19042);
and U19382 (N_19382,N_18840,N_19009);
nand U19383 (N_19383,N_19135,N_19052);
or U19384 (N_19384,N_19133,N_18792);
or U19385 (N_19385,N_19327,N_19287);
nor U19386 (N_19386,N_19157,N_18862);
nor U19387 (N_19387,N_19209,N_18815);
and U19388 (N_19388,N_19152,N_19085);
or U19389 (N_19389,N_19016,N_19190);
or U19390 (N_19390,N_19269,N_19291);
xnor U19391 (N_19391,N_19244,N_18867);
or U19392 (N_19392,N_18813,N_18935);
xor U19393 (N_19393,N_18931,N_19337);
nor U19394 (N_19394,N_18972,N_19206);
nand U19395 (N_19395,N_19268,N_19350);
nand U19396 (N_19396,N_19321,N_19089);
and U19397 (N_19397,N_18873,N_18828);
nor U19398 (N_19398,N_19195,N_18760);
nor U19399 (N_19399,N_19188,N_19194);
and U19400 (N_19400,N_18899,N_19356);
nand U19401 (N_19401,N_19351,N_18806);
nand U19402 (N_19402,N_18766,N_19347);
nand U19403 (N_19403,N_19171,N_18857);
or U19404 (N_19404,N_19116,N_19143);
nand U19405 (N_19405,N_19340,N_19086);
nor U19406 (N_19406,N_19285,N_18791);
nor U19407 (N_19407,N_18753,N_19020);
xor U19408 (N_19408,N_19373,N_18881);
and U19409 (N_19409,N_18933,N_18771);
nor U19410 (N_19410,N_18893,N_19183);
xnor U19411 (N_19411,N_18966,N_19145);
or U19412 (N_19412,N_18779,N_19141);
and U19413 (N_19413,N_18955,N_19300);
nor U19414 (N_19414,N_19304,N_19237);
or U19415 (N_19415,N_19370,N_18913);
and U19416 (N_19416,N_18889,N_19047);
or U19417 (N_19417,N_18863,N_19144);
or U19418 (N_19418,N_19082,N_18936);
or U19419 (N_19419,N_18823,N_18951);
nor U19420 (N_19420,N_18874,N_19202);
nor U19421 (N_19421,N_19094,N_19036);
nand U19422 (N_19422,N_19367,N_19003);
xor U19423 (N_19423,N_18856,N_18953);
nand U19424 (N_19424,N_19056,N_19187);
nand U19425 (N_19425,N_18923,N_18910);
or U19426 (N_19426,N_18905,N_18860);
or U19427 (N_19427,N_19250,N_19101);
xor U19428 (N_19428,N_18793,N_18908);
xor U19429 (N_19429,N_19332,N_18825);
or U19430 (N_19430,N_18979,N_18961);
nand U19431 (N_19431,N_18775,N_19000);
xnor U19432 (N_19432,N_18880,N_19158);
or U19433 (N_19433,N_18892,N_18981);
nand U19434 (N_19434,N_18767,N_19127);
and U19435 (N_19435,N_19212,N_18830);
nor U19436 (N_19436,N_19091,N_18888);
and U19437 (N_19437,N_19197,N_19067);
or U19438 (N_19438,N_19092,N_19164);
xnor U19439 (N_19439,N_18820,N_19177);
nor U19440 (N_19440,N_19069,N_19100);
and U19441 (N_19441,N_19057,N_18963);
and U19442 (N_19442,N_18801,N_19031);
and U19443 (N_19443,N_19245,N_19303);
nand U19444 (N_19444,N_19231,N_19315);
nand U19445 (N_19445,N_19199,N_18934);
or U19446 (N_19446,N_19162,N_18783);
nand U19447 (N_19447,N_18940,N_19252);
nor U19448 (N_19448,N_19153,N_18831);
or U19449 (N_19449,N_19040,N_19239);
xor U19450 (N_19450,N_18900,N_19193);
or U19451 (N_19451,N_19362,N_18802);
and U19452 (N_19452,N_19115,N_18788);
nor U19453 (N_19453,N_18808,N_18773);
nand U19454 (N_19454,N_19147,N_19324);
or U19455 (N_19455,N_19018,N_18759);
nor U19456 (N_19456,N_19038,N_18784);
or U19457 (N_19457,N_18973,N_19130);
or U19458 (N_19458,N_18958,N_19084);
and U19459 (N_19459,N_19150,N_19166);
and U19460 (N_19460,N_18975,N_19265);
xnor U19461 (N_19461,N_19186,N_19023);
nand U19462 (N_19462,N_18970,N_19293);
and U19463 (N_19463,N_19159,N_19241);
and U19464 (N_19464,N_19064,N_19182);
and U19465 (N_19465,N_18890,N_18757);
or U19466 (N_19466,N_19170,N_19322);
nor U19467 (N_19467,N_19323,N_18948);
xnor U19468 (N_19468,N_19176,N_18751);
or U19469 (N_19469,N_19275,N_18996);
and U19470 (N_19470,N_18841,N_19032);
nand U19471 (N_19471,N_18998,N_19219);
and U19472 (N_19472,N_18897,N_18997);
and U19473 (N_19473,N_18962,N_18985);
nand U19474 (N_19474,N_19142,N_18837);
or U19475 (N_19475,N_18916,N_19129);
and U19476 (N_19476,N_19369,N_19372);
and U19477 (N_19477,N_18822,N_18844);
nor U19478 (N_19478,N_19181,N_18778);
and U19479 (N_19479,N_18906,N_19077);
and U19480 (N_19480,N_18918,N_19027);
or U19481 (N_19481,N_19246,N_19251);
nor U19482 (N_19482,N_19290,N_19341);
xnor U19483 (N_19483,N_18922,N_19215);
nand U19484 (N_19484,N_19048,N_18790);
nor U19485 (N_19485,N_18971,N_19336);
nand U19486 (N_19486,N_18817,N_19149);
and U19487 (N_19487,N_19119,N_18843);
and U19488 (N_19488,N_19294,N_18879);
nor U19489 (N_19489,N_18764,N_18870);
xor U19490 (N_19490,N_19041,N_18839);
nand U19491 (N_19491,N_19223,N_19165);
and U19492 (N_19492,N_18989,N_19062);
nand U19493 (N_19493,N_18827,N_19081);
and U19494 (N_19494,N_18804,N_19360);
nand U19495 (N_19495,N_19277,N_19346);
or U19496 (N_19496,N_19095,N_18903);
or U19497 (N_19497,N_19232,N_19266);
xor U19498 (N_19498,N_19026,N_19110);
or U19499 (N_19499,N_19179,N_19112);
and U19500 (N_19500,N_18786,N_18852);
and U19501 (N_19501,N_18920,N_19284);
or U19502 (N_19502,N_18904,N_19228);
nor U19503 (N_19503,N_18782,N_19214);
nand U19504 (N_19504,N_19236,N_18758);
xnor U19505 (N_19505,N_19205,N_19167);
nand U19506 (N_19506,N_19161,N_19055);
xor U19507 (N_19507,N_19121,N_19216);
or U19508 (N_19508,N_19156,N_19124);
nor U19509 (N_19509,N_19050,N_18924);
or U19510 (N_19510,N_19282,N_19146);
or U19511 (N_19511,N_19238,N_19151);
and U19512 (N_19512,N_19028,N_19087);
nand U19513 (N_19513,N_19316,N_19189);
or U19514 (N_19514,N_18886,N_19310);
xnor U19515 (N_19515,N_18858,N_19333);
nand U19516 (N_19516,N_19024,N_18845);
nand U19517 (N_19517,N_19271,N_18947);
nor U19518 (N_19518,N_18978,N_19201);
nand U19519 (N_19519,N_18868,N_19178);
nor U19520 (N_19520,N_19348,N_18969);
or U19521 (N_19521,N_19235,N_19279);
xnor U19522 (N_19522,N_19169,N_19014);
or U19523 (N_19523,N_18912,N_19203);
nand U19524 (N_19524,N_18974,N_19043);
nand U19525 (N_19525,N_19120,N_19218);
xor U19526 (N_19526,N_18950,N_18756);
xnor U19527 (N_19527,N_19353,N_19045);
xnor U19528 (N_19528,N_18838,N_19059);
and U19529 (N_19529,N_19334,N_18930);
nand U19530 (N_19530,N_19292,N_19051);
nand U19531 (N_19531,N_19163,N_18891);
or U19532 (N_19532,N_19273,N_19025);
or U19533 (N_19533,N_19037,N_19261);
or U19534 (N_19534,N_18777,N_18928);
or U19535 (N_19535,N_19256,N_19078);
nor U19536 (N_19536,N_18800,N_18959);
nand U19537 (N_19537,N_18787,N_18945);
or U19538 (N_19538,N_18987,N_18943);
nor U19539 (N_19539,N_19075,N_19317);
xor U19540 (N_19540,N_18929,N_18750);
and U19541 (N_19541,N_18770,N_19058);
xnor U19542 (N_19542,N_19102,N_19011);
nor U19543 (N_19543,N_18849,N_19262);
or U19544 (N_19544,N_18864,N_19286);
nor U19545 (N_19545,N_19008,N_19006);
or U19546 (N_19546,N_19359,N_18762);
and U19547 (N_19547,N_18854,N_19184);
or U19548 (N_19548,N_19005,N_19111);
and U19549 (N_19549,N_19233,N_19076);
nand U19550 (N_19550,N_19301,N_19331);
and U19551 (N_19551,N_18865,N_19012);
or U19552 (N_19552,N_19065,N_19079);
nand U19553 (N_19553,N_18907,N_19320);
or U19554 (N_19554,N_18861,N_18809);
nor U19555 (N_19555,N_19318,N_19103);
and U19556 (N_19556,N_19308,N_19044);
or U19557 (N_19557,N_19221,N_18859);
nor U19558 (N_19558,N_19295,N_18810);
xnor U19559 (N_19559,N_19312,N_18988);
xor U19560 (N_19560,N_18803,N_18772);
and U19561 (N_19561,N_19004,N_19220);
nor U19562 (N_19562,N_18994,N_19148);
or U19563 (N_19563,N_18914,N_19276);
and U19564 (N_19564,N_18965,N_19240);
nand U19565 (N_19565,N_19174,N_18811);
nand U19566 (N_19566,N_19364,N_18896);
and U19567 (N_19567,N_18768,N_18765);
nor U19568 (N_19568,N_18842,N_19243);
and U19569 (N_19569,N_19361,N_19343);
nand U19570 (N_19570,N_18833,N_18774);
and U19571 (N_19571,N_18915,N_18986);
nand U19572 (N_19572,N_18884,N_19210);
and U19573 (N_19573,N_18926,N_18826);
or U19574 (N_19574,N_18993,N_19039);
nand U19575 (N_19575,N_19083,N_19342);
nor U19576 (N_19576,N_19267,N_19108);
xnor U19577 (N_19577,N_18992,N_19309);
xnor U19578 (N_19578,N_19010,N_18967);
nor U19579 (N_19579,N_18853,N_19234);
and U19580 (N_19580,N_18789,N_18902);
nor U19581 (N_19581,N_19154,N_18983);
or U19582 (N_19582,N_18944,N_18816);
or U19583 (N_19583,N_19125,N_18871);
nor U19584 (N_19584,N_19299,N_19097);
nand U19585 (N_19585,N_19128,N_18869);
or U19586 (N_19586,N_18829,N_19107);
nor U19587 (N_19587,N_19306,N_18872);
or U19588 (N_19588,N_19296,N_18901);
nor U19589 (N_19589,N_19017,N_19217);
and U19590 (N_19590,N_18932,N_18885);
nor U19591 (N_19591,N_18834,N_19272);
and U19592 (N_19592,N_18807,N_18909);
nor U19593 (N_19593,N_19106,N_18761);
nand U19594 (N_19594,N_18991,N_19175);
or U19595 (N_19595,N_19222,N_19049);
and U19596 (N_19596,N_19068,N_18836);
and U19597 (N_19597,N_19073,N_19123);
and U19598 (N_19598,N_19330,N_19328);
or U19599 (N_19599,N_19227,N_19109);
nor U19600 (N_19600,N_18847,N_19259);
nor U19601 (N_19601,N_18855,N_18984);
and U19602 (N_19602,N_18964,N_18832);
nand U19603 (N_19603,N_19326,N_18960);
nand U19604 (N_19604,N_19139,N_19242);
nand U19605 (N_19605,N_19113,N_19002);
nand U19606 (N_19606,N_19019,N_18763);
nand U19607 (N_19607,N_19207,N_19180);
xor U19608 (N_19608,N_18824,N_19371);
or U19609 (N_19609,N_18980,N_19224);
nor U19610 (N_19610,N_18898,N_18925);
and U19611 (N_19611,N_18878,N_18946);
or U19612 (N_19612,N_18799,N_19253);
or U19613 (N_19613,N_19200,N_19104);
or U19614 (N_19614,N_18921,N_18785);
and U19615 (N_19615,N_19090,N_19211);
nor U19616 (N_19616,N_19021,N_18805);
nor U19617 (N_19617,N_19365,N_18942);
or U19618 (N_19618,N_19344,N_19263);
nor U19619 (N_19619,N_18835,N_19325);
and U19620 (N_19620,N_19247,N_19329);
and U19621 (N_19621,N_18894,N_18977);
nand U19622 (N_19622,N_19035,N_19264);
nand U19623 (N_19623,N_19374,N_19054);
nand U19624 (N_19624,N_19288,N_19196);
nor U19625 (N_19625,N_18819,N_19033);
or U19626 (N_19626,N_19280,N_19071);
or U19627 (N_19627,N_18949,N_19298);
and U19628 (N_19628,N_19117,N_19099);
nor U19629 (N_19629,N_19278,N_19134);
xnor U19630 (N_19630,N_19155,N_19160);
xor U19631 (N_19631,N_18752,N_19226);
nor U19632 (N_19632,N_18954,N_19230);
and U19633 (N_19633,N_19096,N_19302);
nand U19634 (N_19634,N_19126,N_18755);
nor U19635 (N_19635,N_19198,N_18877);
and U19636 (N_19636,N_18990,N_19063);
nand U19637 (N_19637,N_19213,N_19357);
nor U19638 (N_19638,N_19136,N_19339);
or U19639 (N_19639,N_19185,N_18850);
nor U19640 (N_19640,N_19022,N_19254);
and U19641 (N_19641,N_19366,N_18957);
and U19642 (N_19642,N_19053,N_19007);
nor U19643 (N_19643,N_19274,N_19137);
and U19644 (N_19644,N_18846,N_19249);
nor U19645 (N_19645,N_19191,N_18976);
or U19646 (N_19646,N_19255,N_19105);
or U19647 (N_19647,N_19168,N_19258);
or U19648 (N_19648,N_18812,N_18887);
or U19649 (N_19649,N_19289,N_18968);
or U19650 (N_19650,N_19080,N_18982);
nor U19651 (N_19651,N_19013,N_19060);
nor U19652 (N_19652,N_19172,N_19307);
nand U19653 (N_19653,N_19074,N_18882);
nor U19654 (N_19654,N_18895,N_19355);
or U19655 (N_19655,N_18919,N_18927);
and U19656 (N_19656,N_18938,N_18851);
or U19657 (N_19657,N_19358,N_18952);
and U19658 (N_19658,N_18818,N_18995);
nor U19659 (N_19659,N_19352,N_19297);
and U19660 (N_19660,N_18769,N_19061);
xnor U19661 (N_19661,N_18781,N_19070);
or U19662 (N_19662,N_19030,N_19066);
and U19663 (N_19663,N_19034,N_19114);
nand U19664 (N_19664,N_19335,N_18821);
and U19665 (N_19665,N_18883,N_18798);
nand U19666 (N_19666,N_19118,N_19072);
and U19667 (N_19667,N_19138,N_19122);
nor U19668 (N_19668,N_19093,N_18794);
nand U19669 (N_19669,N_19132,N_18795);
or U19670 (N_19670,N_18754,N_18876);
and U19671 (N_19671,N_18911,N_19368);
or U19672 (N_19672,N_19349,N_19338);
and U19673 (N_19673,N_19281,N_18941);
xor U19674 (N_19674,N_19098,N_18796);
nor U19675 (N_19675,N_19313,N_19029);
nor U19676 (N_19676,N_19257,N_19319);
and U19677 (N_19677,N_19088,N_19046);
nand U19678 (N_19678,N_18917,N_19131);
or U19679 (N_19679,N_19015,N_18999);
or U19680 (N_19680,N_18797,N_19311);
or U19681 (N_19681,N_18956,N_19001);
xor U19682 (N_19682,N_19354,N_19229);
nor U19683 (N_19683,N_19204,N_18848);
and U19684 (N_19684,N_18866,N_19225);
nand U19685 (N_19685,N_19248,N_19283);
or U19686 (N_19686,N_18776,N_19345);
nor U19687 (N_19687,N_18939,N_18817);
xnor U19688 (N_19688,N_18894,N_19337);
and U19689 (N_19689,N_19272,N_19142);
nand U19690 (N_19690,N_19097,N_19139);
nand U19691 (N_19691,N_18806,N_19139);
nand U19692 (N_19692,N_19361,N_18825);
and U19693 (N_19693,N_19223,N_18958);
and U19694 (N_19694,N_18949,N_19262);
and U19695 (N_19695,N_18774,N_19355);
or U19696 (N_19696,N_19336,N_18767);
nor U19697 (N_19697,N_19193,N_18872);
and U19698 (N_19698,N_19095,N_18762);
and U19699 (N_19699,N_18852,N_19252);
or U19700 (N_19700,N_19021,N_19178);
nor U19701 (N_19701,N_18949,N_19218);
and U19702 (N_19702,N_19254,N_19153);
or U19703 (N_19703,N_18845,N_18909);
xnor U19704 (N_19704,N_19359,N_19213);
xnor U19705 (N_19705,N_18978,N_18929);
nor U19706 (N_19706,N_19001,N_18759);
nor U19707 (N_19707,N_19320,N_19370);
or U19708 (N_19708,N_19098,N_18806);
nor U19709 (N_19709,N_18877,N_18869);
or U19710 (N_19710,N_18758,N_18817);
nand U19711 (N_19711,N_19172,N_19005);
and U19712 (N_19712,N_18984,N_19160);
and U19713 (N_19713,N_19187,N_18892);
nand U19714 (N_19714,N_19109,N_18984);
or U19715 (N_19715,N_18983,N_19327);
nand U19716 (N_19716,N_19147,N_19085);
nor U19717 (N_19717,N_18988,N_18986);
and U19718 (N_19718,N_18826,N_19322);
nor U19719 (N_19719,N_19264,N_19041);
nand U19720 (N_19720,N_18897,N_19359);
nand U19721 (N_19721,N_18944,N_19183);
nand U19722 (N_19722,N_18868,N_18819);
nand U19723 (N_19723,N_19120,N_19115);
nor U19724 (N_19724,N_18816,N_18975);
nor U19725 (N_19725,N_19068,N_19171);
nor U19726 (N_19726,N_19162,N_18753);
or U19727 (N_19727,N_18952,N_18766);
and U19728 (N_19728,N_19028,N_19312);
or U19729 (N_19729,N_18957,N_18949);
or U19730 (N_19730,N_18879,N_18758);
and U19731 (N_19731,N_19025,N_18769);
nor U19732 (N_19732,N_19212,N_18789);
nor U19733 (N_19733,N_18803,N_18847);
nand U19734 (N_19734,N_19329,N_19291);
nor U19735 (N_19735,N_19178,N_18855);
nand U19736 (N_19736,N_19065,N_18970);
nand U19737 (N_19737,N_18965,N_19036);
or U19738 (N_19738,N_19238,N_19306);
and U19739 (N_19739,N_19226,N_18943);
nand U19740 (N_19740,N_19016,N_19005);
and U19741 (N_19741,N_18994,N_18874);
nor U19742 (N_19742,N_19131,N_18982);
nor U19743 (N_19743,N_19073,N_18902);
nand U19744 (N_19744,N_19325,N_19076);
nor U19745 (N_19745,N_18752,N_19026);
and U19746 (N_19746,N_19371,N_19352);
nand U19747 (N_19747,N_18794,N_18925);
nand U19748 (N_19748,N_19263,N_19175);
nor U19749 (N_19749,N_18857,N_19127);
nor U19750 (N_19750,N_19293,N_19264);
and U19751 (N_19751,N_19264,N_19170);
and U19752 (N_19752,N_19139,N_18804);
nand U19753 (N_19753,N_19150,N_19066);
and U19754 (N_19754,N_18976,N_19005);
or U19755 (N_19755,N_18894,N_19374);
nor U19756 (N_19756,N_18832,N_19290);
nor U19757 (N_19757,N_18779,N_19361);
xnor U19758 (N_19758,N_19127,N_19120);
nor U19759 (N_19759,N_19132,N_18864);
nor U19760 (N_19760,N_19345,N_19167);
and U19761 (N_19761,N_18761,N_19336);
nand U19762 (N_19762,N_19364,N_19047);
and U19763 (N_19763,N_18789,N_18975);
and U19764 (N_19764,N_19035,N_18845);
nor U19765 (N_19765,N_18866,N_19144);
nor U19766 (N_19766,N_19004,N_18842);
nand U19767 (N_19767,N_18875,N_19187);
and U19768 (N_19768,N_18884,N_18837);
nand U19769 (N_19769,N_19066,N_18970);
nand U19770 (N_19770,N_19079,N_18870);
nand U19771 (N_19771,N_19265,N_18996);
and U19772 (N_19772,N_19118,N_18766);
or U19773 (N_19773,N_19248,N_19185);
xor U19774 (N_19774,N_19201,N_18968);
nor U19775 (N_19775,N_19238,N_19054);
nor U19776 (N_19776,N_19352,N_18865);
xor U19777 (N_19777,N_19016,N_18979);
xor U19778 (N_19778,N_18821,N_19193);
nand U19779 (N_19779,N_18907,N_19234);
nor U19780 (N_19780,N_19371,N_19316);
nand U19781 (N_19781,N_19106,N_19259);
or U19782 (N_19782,N_18767,N_19205);
nor U19783 (N_19783,N_19030,N_19019);
and U19784 (N_19784,N_19107,N_18969);
or U19785 (N_19785,N_19198,N_18942);
nor U19786 (N_19786,N_19355,N_19301);
nor U19787 (N_19787,N_18855,N_19229);
xnor U19788 (N_19788,N_19073,N_18841);
and U19789 (N_19789,N_19222,N_19365);
nand U19790 (N_19790,N_19020,N_19153);
nor U19791 (N_19791,N_18970,N_18792);
and U19792 (N_19792,N_19222,N_19251);
or U19793 (N_19793,N_18981,N_18924);
or U19794 (N_19794,N_19237,N_19316);
nor U19795 (N_19795,N_18895,N_19064);
and U19796 (N_19796,N_19133,N_19203);
nor U19797 (N_19797,N_18781,N_18905);
xnor U19798 (N_19798,N_19011,N_19277);
or U19799 (N_19799,N_19189,N_18993);
or U19800 (N_19800,N_18849,N_19091);
and U19801 (N_19801,N_19213,N_19247);
and U19802 (N_19802,N_19368,N_18765);
nor U19803 (N_19803,N_19157,N_19245);
nand U19804 (N_19804,N_19038,N_19143);
nand U19805 (N_19805,N_18849,N_18912);
xor U19806 (N_19806,N_18987,N_19280);
or U19807 (N_19807,N_19031,N_19005);
nand U19808 (N_19808,N_19279,N_18896);
and U19809 (N_19809,N_18981,N_18973);
or U19810 (N_19810,N_18845,N_19195);
nor U19811 (N_19811,N_19138,N_19211);
nor U19812 (N_19812,N_19030,N_19276);
or U19813 (N_19813,N_18811,N_18832);
nor U19814 (N_19814,N_19225,N_19103);
xor U19815 (N_19815,N_19342,N_19356);
nor U19816 (N_19816,N_18838,N_18839);
or U19817 (N_19817,N_19062,N_18828);
nor U19818 (N_19818,N_19345,N_19042);
xor U19819 (N_19819,N_19129,N_19167);
or U19820 (N_19820,N_19239,N_19119);
nand U19821 (N_19821,N_18916,N_19009);
nand U19822 (N_19822,N_19200,N_19046);
or U19823 (N_19823,N_18902,N_18856);
or U19824 (N_19824,N_19348,N_19051);
nor U19825 (N_19825,N_18914,N_18819);
or U19826 (N_19826,N_18989,N_18921);
or U19827 (N_19827,N_18960,N_18914);
nand U19828 (N_19828,N_18811,N_18829);
or U19829 (N_19829,N_19176,N_19323);
xor U19830 (N_19830,N_19114,N_18924);
or U19831 (N_19831,N_19299,N_19212);
or U19832 (N_19832,N_19202,N_18890);
nand U19833 (N_19833,N_19301,N_19047);
and U19834 (N_19834,N_19189,N_18785);
and U19835 (N_19835,N_19092,N_19243);
nor U19836 (N_19836,N_18908,N_19315);
and U19837 (N_19837,N_19059,N_19121);
or U19838 (N_19838,N_19165,N_18851);
xnor U19839 (N_19839,N_19083,N_19087);
nand U19840 (N_19840,N_19233,N_18873);
and U19841 (N_19841,N_19035,N_19237);
or U19842 (N_19842,N_19020,N_18970);
nand U19843 (N_19843,N_18836,N_18859);
and U19844 (N_19844,N_19059,N_19132);
nor U19845 (N_19845,N_18858,N_18868);
nor U19846 (N_19846,N_19095,N_19046);
or U19847 (N_19847,N_18797,N_18946);
or U19848 (N_19848,N_19327,N_18891);
xnor U19849 (N_19849,N_19126,N_19116);
or U19850 (N_19850,N_19065,N_19239);
nor U19851 (N_19851,N_18832,N_19201);
and U19852 (N_19852,N_19117,N_19331);
nor U19853 (N_19853,N_18993,N_19101);
or U19854 (N_19854,N_19068,N_19255);
or U19855 (N_19855,N_19007,N_19369);
nand U19856 (N_19856,N_19184,N_19342);
nand U19857 (N_19857,N_19195,N_19023);
nand U19858 (N_19858,N_18854,N_18913);
or U19859 (N_19859,N_19372,N_19061);
and U19860 (N_19860,N_18874,N_19149);
nor U19861 (N_19861,N_19105,N_18920);
and U19862 (N_19862,N_19003,N_19331);
or U19863 (N_19863,N_19002,N_18912);
or U19864 (N_19864,N_19186,N_19006);
xnor U19865 (N_19865,N_18973,N_18954);
or U19866 (N_19866,N_19096,N_18758);
or U19867 (N_19867,N_19338,N_19046);
nor U19868 (N_19868,N_19120,N_18896);
or U19869 (N_19869,N_19128,N_19219);
and U19870 (N_19870,N_19216,N_18900);
and U19871 (N_19871,N_19092,N_19269);
nand U19872 (N_19872,N_18779,N_18920);
nor U19873 (N_19873,N_18910,N_18882);
and U19874 (N_19874,N_18824,N_18779);
or U19875 (N_19875,N_18841,N_18952);
nand U19876 (N_19876,N_18994,N_18979);
nand U19877 (N_19877,N_18937,N_19351);
or U19878 (N_19878,N_19216,N_19153);
nor U19879 (N_19879,N_18803,N_19355);
xor U19880 (N_19880,N_19309,N_18808);
nor U19881 (N_19881,N_18762,N_19041);
and U19882 (N_19882,N_18834,N_19290);
nor U19883 (N_19883,N_18963,N_19138);
nor U19884 (N_19884,N_19063,N_19176);
or U19885 (N_19885,N_19267,N_18983);
and U19886 (N_19886,N_19215,N_19065);
nor U19887 (N_19887,N_19141,N_18891);
and U19888 (N_19888,N_19280,N_19011);
or U19889 (N_19889,N_19031,N_18767);
and U19890 (N_19890,N_19146,N_19319);
xor U19891 (N_19891,N_19132,N_18797);
and U19892 (N_19892,N_19320,N_18781);
and U19893 (N_19893,N_19266,N_19110);
nor U19894 (N_19894,N_18803,N_18842);
nand U19895 (N_19895,N_18977,N_19022);
nand U19896 (N_19896,N_19284,N_19350);
xnor U19897 (N_19897,N_19087,N_18788);
and U19898 (N_19898,N_19147,N_19008);
and U19899 (N_19899,N_19342,N_19258);
nor U19900 (N_19900,N_19326,N_19110);
and U19901 (N_19901,N_18796,N_18836);
nand U19902 (N_19902,N_19200,N_19265);
nor U19903 (N_19903,N_19028,N_18864);
and U19904 (N_19904,N_19321,N_19005);
nand U19905 (N_19905,N_19042,N_19011);
or U19906 (N_19906,N_18794,N_19028);
or U19907 (N_19907,N_19170,N_18845);
nand U19908 (N_19908,N_19157,N_18934);
xnor U19909 (N_19909,N_18968,N_19252);
and U19910 (N_19910,N_18982,N_19322);
and U19911 (N_19911,N_18946,N_19361);
nand U19912 (N_19912,N_19299,N_18949);
nor U19913 (N_19913,N_19074,N_18772);
nor U19914 (N_19914,N_18973,N_18791);
or U19915 (N_19915,N_19325,N_19254);
nand U19916 (N_19916,N_19025,N_19168);
nand U19917 (N_19917,N_18980,N_19325);
nor U19918 (N_19918,N_18875,N_19112);
xnor U19919 (N_19919,N_19050,N_18944);
xor U19920 (N_19920,N_18758,N_19001);
and U19921 (N_19921,N_19028,N_19140);
nand U19922 (N_19922,N_19316,N_18813);
xnor U19923 (N_19923,N_19043,N_19089);
or U19924 (N_19924,N_18970,N_18917);
nor U19925 (N_19925,N_19360,N_19188);
nor U19926 (N_19926,N_18971,N_18956);
nand U19927 (N_19927,N_18790,N_18769);
nor U19928 (N_19928,N_19062,N_18926);
and U19929 (N_19929,N_18812,N_19337);
or U19930 (N_19930,N_19060,N_19033);
xnor U19931 (N_19931,N_19120,N_18832);
or U19932 (N_19932,N_19160,N_19029);
and U19933 (N_19933,N_19269,N_18779);
or U19934 (N_19934,N_19212,N_18847);
and U19935 (N_19935,N_18914,N_19309);
nor U19936 (N_19936,N_18844,N_19345);
xnor U19937 (N_19937,N_18993,N_19334);
or U19938 (N_19938,N_19149,N_18885);
or U19939 (N_19939,N_19231,N_18786);
or U19940 (N_19940,N_19009,N_18760);
or U19941 (N_19941,N_18915,N_19130);
xnor U19942 (N_19942,N_19145,N_18893);
and U19943 (N_19943,N_19290,N_18948);
nand U19944 (N_19944,N_19203,N_19147);
xor U19945 (N_19945,N_19209,N_18980);
and U19946 (N_19946,N_19372,N_18828);
and U19947 (N_19947,N_18804,N_18865);
or U19948 (N_19948,N_18818,N_19130);
nand U19949 (N_19949,N_18988,N_19270);
and U19950 (N_19950,N_19096,N_18879);
xor U19951 (N_19951,N_18812,N_18788);
nor U19952 (N_19952,N_19315,N_18877);
xnor U19953 (N_19953,N_18871,N_18915);
nand U19954 (N_19954,N_18774,N_18810);
xor U19955 (N_19955,N_19343,N_19316);
xnor U19956 (N_19956,N_19183,N_19250);
nand U19957 (N_19957,N_18968,N_19358);
or U19958 (N_19958,N_18912,N_19218);
nand U19959 (N_19959,N_18850,N_19110);
nor U19960 (N_19960,N_19043,N_19103);
or U19961 (N_19961,N_19236,N_18797);
or U19962 (N_19962,N_19253,N_18966);
nand U19963 (N_19963,N_19234,N_19140);
xor U19964 (N_19964,N_19183,N_19275);
and U19965 (N_19965,N_19290,N_19025);
or U19966 (N_19966,N_18788,N_18769);
nor U19967 (N_19967,N_18782,N_19368);
and U19968 (N_19968,N_19230,N_19072);
nand U19969 (N_19969,N_19050,N_19013);
and U19970 (N_19970,N_18792,N_19197);
and U19971 (N_19971,N_19183,N_19205);
or U19972 (N_19972,N_19161,N_18879);
xor U19973 (N_19973,N_19103,N_19313);
and U19974 (N_19974,N_19141,N_19029);
and U19975 (N_19975,N_19125,N_19146);
nor U19976 (N_19976,N_18762,N_19302);
nor U19977 (N_19977,N_19255,N_18975);
or U19978 (N_19978,N_19357,N_19261);
nor U19979 (N_19979,N_19111,N_18824);
or U19980 (N_19980,N_19028,N_19036);
nand U19981 (N_19981,N_19130,N_18919);
or U19982 (N_19982,N_19217,N_18776);
nor U19983 (N_19983,N_19064,N_19030);
xor U19984 (N_19984,N_19290,N_18757);
nor U19985 (N_19985,N_19137,N_18763);
and U19986 (N_19986,N_18867,N_19137);
or U19987 (N_19987,N_19034,N_18875);
xor U19988 (N_19988,N_19371,N_19148);
or U19989 (N_19989,N_19326,N_18971);
and U19990 (N_19990,N_19369,N_18843);
nand U19991 (N_19991,N_19161,N_18776);
nor U19992 (N_19992,N_19238,N_19268);
xor U19993 (N_19993,N_19281,N_19097);
or U19994 (N_19994,N_18898,N_18890);
and U19995 (N_19995,N_18902,N_18932);
and U19996 (N_19996,N_18871,N_19118);
nand U19997 (N_19997,N_18762,N_19352);
nand U19998 (N_19998,N_19230,N_19369);
nor U19999 (N_19999,N_19054,N_19167);
and U20000 (N_20000,N_19557,N_19488);
or U20001 (N_20001,N_19762,N_19925);
and U20002 (N_20002,N_19969,N_19394);
nor U20003 (N_20003,N_19595,N_19763);
or U20004 (N_20004,N_19566,N_19503);
nand U20005 (N_20005,N_19842,N_19779);
and U20006 (N_20006,N_19849,N_19623);
and U20007 (N_20007,N_19630,N_19568);
or U20008 (N_20008,N_19543,N_19975);
and U20009 (N_20009,N_19793,N_19482);
or U20010 (N_20010,N_19963,N_19855);
nor U20011 (N_20011,N_19902,N_19754);
or U20012 (N_20012,N_19714,N_19713);
nand U20013 (N_20013,N_19625,N_19863);
or U20014 (N_20014,N_19706,N_19947);
or U20015 (N_20015,N_19799,N_19388);
nand U20016 (N_20016,N_19632,N_19689);
nand U20017 (N_20017,N_19945,N_19476);
nand U20018 (N_20018,N_19585,N_19679);
and U20019 (N_20019,N_19937,N_19845);
and U20020 (N_20020,N_19796,N_19742);
nor U20021 (N_20021,N_19724,N_19446);
nand U20022 (N_20022,N_19577,N_19899);
xnor U20023 (N_20023,N_19429,N_19660);
nor U20024 (N_20024,N_19470,N_19750);
and U20025 (N_20025,N_19997,N_19616);
nor U20026 (N_20026,N_19390,N_19594);
nand U20027 (N_20027,N_19564,N_19588);
or U20028 (N_20028,N_19707,N_19556);
nor U20029 (N_20029,N_19619,N_19574);
or U20030 (N_20030,N_19560,N_19930);
and U20031 (N_20031,N_19803,N_19752);
or U20032 (N_20032,N_19927,N_19965);
or U20033 (N_20033,N_19719,N_19434);
and U20034 (N_20034,N_19549,N_19650);
and U20035 (N_20035,N_19596,N_19696);
nand U20036 (N_20036,N_19573,N_19634);
and U20037 (N_20037,N_19960,N_19858);
xor U20038 (N_20038,N_19904,N_19738);
nor U20039 (N_20039,N_19915,N_19721);
nand U20040 (N_20040,N_19415,N_19489);
and U20041 (N_20041,N_19726,N_19532);
or U20042 (N_20042,N_19479,N_19455);
nor U20043 (N_20043,N_19946,N_19758);
and U20044 (N_20044,N_19867,N_19493);
nand U20045 (N_20045,N_19962,N_19983);
nand U20046 (N_20046,N_19697,N_19545);
nor U20047 (N_20047,N_19398,N_19408);
nand U20048 (N_20048,N_19513,N_19467);
and U20049 (N_20049,N_19744,N_19993);
nand U20050 (N_20050,N_19686,N_19868);
nand U20051 (N_20051,N_19575,N_19458);
nand U20052 (N_20052,N_19943,N_19882);
and U20053 (N_20053,N_19454,N_19794);
xnor U20054 (N_20054,N_19741,N_19802);
and U20055 (N_20055,N_19501,N_19584);
xor U20056 (N_20056,N_19675,N_19773);
or U20057 (N_20057,N_19691,N_19959);
xnor U20058 (N_20058,N_19857,N_19729);
or U20059 (N_20059,N_19603,N_19693);
nand U20060 (N_20060,N_19774,N_19526);
and U20061 (N_20061,N_19643,N_19627);
nand U20062 (N_20062,N_19725,N_19905);
and U20063 (N_20063,N_19480,N_19912);
and U20064 (N_20064,N_19539,N_19417);
or U20065 (N_20065,N_19524,N_19816);
or U20066 (N_20066,N_19866,N_19984);
and U20067 (N_20067,N_19778,N_19921);
and U20068 (N_20068,N_19854,N_19777);
xor U20069 (N_20069,N_19880,N_19824);
or U20070 (N_20070,N_19391,N_19843);
xnor U20071 (N_20071,N_19807,N_19734);
and U20072 (N_20072,N_19544,N_19520);
nand U20073 (N_20073,N_19386,N_19471);
or U20074 (N_20074,N_19582,N_19720);
xnor U20075 (N_20075,N_19892,N_19887);
xor U20076 (N_20076,N_19635,N_19486);
nand U20077 (N_20077,N_19525,N_19615);
or U20078 (N_20078,N_19590,N_19812);
xor U20079 (N_20079,N_19604,N_19514);
nand U20080 (N_20080,N_19387,N_19555);
or U20081 (N_20081,N_19425,N_19497);
or U20082 (N_20082,N_19864,N_19416);
and U20083 (N_20083,N_19607,N_19620);
or U20084 (N_20084,N_19688,N_19547);
or U20085 (N_20085,N_19654,N_19835);
nor U20086 (N_20086,N_19700,N_19533);
nand U20087 (N_20087,N_19841,N_19920);
nand U20088 (N_20088,N_19780,N_19562);
or U20089 (N_20089,N_19669,N_19808);
and U20090 (N_20090,N_19929,N_19822);
or U20091 (N_20091,N_19468,N_19940);
or U20092 (N_20092,N_19901,N_19475);
and U20093 (N_20093,N_19678,N_19382);
nor U20094 (N_20094,N_19839,N_19976);
xor U20095 (N_20095,N_19487,N_19610);
nand U20096 (N_20096,N_19916,N_19601);
and U20097 (N_20097,N_19759,N_19834);
or U20098 (N_20098,N_19571,N_19606);
or U20099 (N_20099,N_19553,N_19837);
nand U20100 (N_20100,N_19414,N_19860);
nand U20101 (N_20101,N_19403,N_19847);
nand U20102 (N_20102,N_19853,N_19385);
or U20103 (N_20103,N_19889,N_19448);
xnor U20104 (N_20104,N_19612,N_19450);
nand U20105 (N_20105,N_19683,N_19576);
nor U20106 (N_20106,N_19551,N_19751);
nand U20107 (N_20107,N_19666,N_19756);
and U20108 (N_20108,N_19917,N_19626);
nor U20109 (N_20109,N_19891,N_19699);
xnor U20110 (N_20110,N_19953,N_19961);
nor U20111 (N_20111,N_19787,N_19609);
or U20112 (N_20112,N_19786,N_19465);
and U20113 (N_20113,N_19814,N_19770);
or U20114 (N_20114,N_19936,N_19733);
or U20115 (N_20115,N_19833,N_19636);
nand U20116 (N_20116,N_19859,N_19852);
or U20117 (N_20117,N_19405,N_19548);
or U20118 (N_20118,N_19851,N_19379);
and U20119 (N_20119,N_19954,N_19638);
xor U20120 (N_20120,N_19771,N_19376);
nor U20121 (N_20121,N_19844,N_19783);
nand U20122 (N_20122,N_19810,N_19979);
nor U20123 (N_20123,N_19667,N_19884);
and U20124 (N_20124,N_19830,N_19529);
and U20125 (N_20125,N_19437,N_19523);
nand U20126 (N_20126,N_19875,N_19519);
and U20127 (N_20127,N_19651,N_19587);
or U20128 (N_20128,N_19500,N_19644);
nand U20129 (N_20129,N_19765,N_19570);
nand U20130 (N_20130,N_19941,N_19591);
or U20131 (N_20131,N_19980,N_19420);
or U20132 (N_20132,N_19788,N_19723);
and U20133 (N_20133,N_19516,N_19443);
nand U20134 (N_20134,N_19978,N_19659);
xnor U20135 (N_20135,N_19813,N_19491);
xnor U20136 (N_20136,N_19994,N_19618);
nor U20137 (N_20137,N_19567,N_19730);
nor U20138 (N_20138,N_19861,N_19657);
nand U20139 (N_20139,N_19732,N_19641);
nand U20140 (N_20140,N_19749,N_19484);
and U20141 (N_20141,N_19970,N_19438);
nor U20142 (N_20142,N_19670,N_19422);
nand U20143 (N_20143,N_19809,N_19820);
xor U20144 (N_20144,N_19764,N_19561);
and U20145 (N_20145,N_19922,N_19435);
and U20146 (N_20146,N_19581,N_19512);
nand U20147 (N_20147,N_19890,N_19451);
or U20148 (N_20148,N_19938,N_19400);
or U20149 (N_20149,N_19614,N_19597);
xor U20150 (N_20150,N_19613,N_19428);
or U20151 (N_20151,N_19897,N_19459);
nand U20152 (N_20152,N_19888,N_19492);
and U20153 (N_20153,N_19554,N_19878);
or U20154 (N_20154,N_19506,N_19461);
nand U20155 (N_20155,N_19444,N_19541);
xor U20156 (N_20156,N_19998,N_19622);
or U20157 (N_20157,N_19537,N_19848);
nand U20158 (N_20158,N_19424,N_19407);
xnor U20159 (N_20159,N_19441,N_19818);
and U20160 (N_20160,N_19914,N_19456);
or U20161 (N_20161,N_19766,N_19846);
xnor U20162 (N_20162,N_19426,N_19410);
xor U20163 (N_20163,N_19474,N_19423);
nor U20164 (N_20164,N_19727,N_19578);
nand U20165 (N_20165,N_19563,N_19681);
xnor U20166 (N_20166,N_19982,N_19973);
and U20167 (N_20167,N_19692,N_19419);
or U20168 (N_20168,N_19785,N_19502);
nor U20169 (N_20169,N_19992,N_19649);
nand U20170 (N_20170,N_19457,N_19442);
nand U20171 (N_20171,N_19792,N_19781);
nor U20172 (N_20172,N_19886,N_19999);
and U20173 (N_20173,N_19495,N_19736);
nand U20174 (N_20174,N_19977,N_19430);
nand U20175 (N_20175,N_19894,N_19815);
nor U20176 (N_20176,N_19665,N_19447);
xor U20177 (N_20177,N_19440,N_19798);
and U20178 (N_20178,N_19522,N_19827);
nand U20179 (N_20179,N_19731,N_19392);
or U20180 (N_20180,N_19509,N_19821);
and U20181 (N_20181,N_19913,N_19510);
or U20182 (N_20182,N_19378,N_19462);
nand U20183 (N_20183,N_19988,N_19645);
nand U20184 (N_20184,N_19873,N_19381);
nand U20185 (N_20185,N_19935,N_19923);
nand U20186 (N_20186,N_19605,N_19629);
nand U20187 (N_20187,N_19735,N_19789);
and U20188 (N_20188,N_19705,N_19748);
or U20189 (N_20189,N_19755,N_19445);
and U20190 (N_20190,N_19710,N_19974);
nand U20191 (N_20191,N_19463,N_19530);
and U20192 (N_20192,N_19828,N_19986);
nor U20193 (N_20193,N_19949,N_19637);
nand U20194 (N_20194,N_19739,N_19608);
xor U20195 (N_20195,N_19987,N_19478);
or U20196 (N_20196,N_19599,N_19746);
nor U20197 (N_20197,N_19964,N_19896);
or U20198 (N_20198,N_19647,N_19850);
and U20199 (N_20199,N_19939,N_19804);
and U20200 (N_20200,N_19399,N_19377);
and U20201 (N_20201,N_19879,N_19690);
and U20202 (N_20202,N_19825,N_19682);
or U20203 (N_20203,N_19704,N_19611);
nand U20204 (N_20204,N_19421,N_19481);
nand U20205 (N_20205,N_19711,N_19684);
nand U20206 (N_20206,N_19586,N_19527);
or U20207 (N_20207,N_19743,N_19401);
nand U20208 (N_20208,N_19663,N_19671);
nor U20209 (N_20209,N_19900,N_19717);
and U20210 (N_20210,N_19473,N_19413);
nor U20211 (N_20211,N_19477,N_19996);
and U20212 (N_20212,N_19673,N_19593);
nand U20213 (N_20213,N_19972,N_19602);
and U20214 (N_20214,N_19862,N_19499);
and U20215 (N_20215,N_19956,N_19968);
nor U20216 (N_20216,N_19712,N_19811);
nor U20217 (N_20217,N_19715,N_19436);
and U20218 (N_20218,N_19515,N_19800);
nand U20219 (N_20219,N_19757,N_19652);
or U20220 (N_20220,N_19559,N_19709);
nor U20221 (N_20221,N_19542,N_19579);
nor U20222 (N_20222,N_19795,N_19589);
nand U20223 (N_20223,N_19661,N_19664);
xnor U20224 (N_20224,N_19791,N_19538);
or U20225 (N_20225,N_19942,N_19680);
and U20226 (N_20226,N_19640,N_19535);
and U20227 (N_20227,N_19952,N_19452);
nand U20228 (N_20228,N_19885,N_19832);
or U20229 (N_20229,N_19404,N_19883);
nor U20230 (N_20230,N_19919,N_19427);
nor U20231 (N_20231,N_19797,N_19469);
or U20232 (N_20232,N_19685,N_19817);
xnor U20233 (N_20233,N_19869,N_19775);
nor U20234 (N_20234,N_19865,N_19384);
or U20235 (N_20235,N_19881,N_19776);
or U20236 (N_20236,N_19950,N_19662);
xnor U20237 (N_20237,N_19874,N_19558);
nor U20238 (N_20238,N_19656,N_19870);
and U20239 (N_20239,N_19550,N_19985);
or U20240 (N_20240,N_19546,N_19910);
nand U20241 (N_20241,N_19698,N_19677);
nor U20242 (N_20242,N_19383,N_19831);
nand U20243 (N_20243,N_19967,N_19722);
or U20244 (N_20244,N_19989,N_19395);
and U20245 (N_20245,N_19624,N_19655);
nor U20246 (N_20246,N_19909,N_19871);
or U20247 (N_20247,N_19521,N_19406);
xnor U20248 (N_20248,N_19701,N_19536);
or U20249 (N_20249,N_19494,N_19876);
nand U20250 (N_20250,N_19453,N_19924);
nand U20251 (N_20251,N_19971,N_19639);
nor U20252 (N_20252,N_19621,N_19931);
xnor U20253 (N_20253,N_19995,N_19716);
or U20254 (N_20254,N_19432,N_19375);
or U20255 (N_20255,N_19397,N_19840);
or U20256 (N_20256,N_19958,N_19790);
nor U20257 (N_20257,N_19511,N_19402);
and U20258 (N_20258,N_19466,N_19806);
nor U20259 (N_20259,N_19668,N_19583);
or U20260 (N_20260,N_19653,N_19801);
or U20261 (N_20261,N_19768,N_19694);
nor U20262 (N_20262,N_19496,N_19507);
and U20263 (N_20263,N_19966,N_19418);
nand U20264 (N_20264,N_19838,N_19528);
nand U20265 (N_20265,N_19895,N_19926);
and U20266 (N_20266,N_19592,N_19598);
nor U20267 (N_20267,N_19893,N_19631);
nand U20268 (N_20268,N_19829,N_19753);
or U20269 (N_20269,N_19490,N_19819);
or U20270 (N_20270,N_19981,N_19918);
nand U20271 (N_20271,N_19951,N_19745);
or U20272 (N_20272,N_19540,N_19439);
nor U20273 (N_20273,N_19805,N_19648);
or U20274 (N_20274,N_19552,N_19464);
and U20275 (N_20275,N_19695,N_19856);
and U20276 (N_20276,N_19782,N_19460);
and U20277 (N_20277,N_19903,N_19504);
or U20278 (N_20278,N_19565,N_19580);
nand U20279 (N_20279,N_19955,N_19633);
or U20280 (N_20280,N_19642,N_19534);
nor U20281 (N_20281,N_19672,N_19784);
nand U20282 (N_20282,N_19411,N_19702);
and U20283 (N_20283,N_19396,N_19991);
xor U20284 (N_20284,N_19747,N_19737);
and U20285 (N_20285,N_19517,N_19767);
nor U20286 (N_20286,N_19728,N_19908);
or U20287 (N_20287,N_19472,N_19569);
nor U20288 (N_20288,N_19483,N_19628);
nor U20289 (N_20289,N_19934,N_19772);
nand U20290 (N_20290,N_19932,N_19948);
and U20291 (N_20291,N_19761,N_19531);
nor U20292 (N_20292,N_19877,N_19906);
nand U20293 (N_20293,N_19409,N_19836);
nor U20294 (N_20294,N_19907,N_19718);
or U20295 (N_20295,N_19823,N_19572);
and U20296 (N_20296,N_19760,N_19498);
nand U20297 (N_20297,N_19658,N_19389);
xnor U20298 (N_20298,N_19380,N_19990);
and U20299 (N_20299,N_19617,N_19518);
nand U20300 (N_20300,N_19933,N_19393);
xnor U20301 (N_20301,N_19646,N_19431);
and U20302 (N_20302,N_19703,N_19676);
nor U20303 (N_20303,N_19944,N_19687);
and U20304 (N_20304,N_19957,N_19740);
or U20305 (N_20305,N_19674,N_19898);
and U20306 (N_20306,N_19505,N_19508);
and U20307 (N_20307,N_19826,N_19485);
nand U20308 (N_20308,N_19708,N_19449);
or U20309 (N_20309,N_19433,N_19928);
nand U20310 (N_20310,N_19412,N_19769);
xnor U20311 (N_20311,N_19872,N_19600);
nor U20312 (N_20312,N_19911,N_19786);
and U20313 (N_20313,N_19803,N_19473);
nor U20314 (N_20314,N_19443,N_19890);
nor U20315 (N_20315,N_19584,N_19740);
nand U20316 (N_20316,N_19784,N_19499);
nand U20317 (N_20317,N_19697,N_19591);
and U20318 (N_20318,N_19630,N_19917);
or U20319 (N_20319,N_19854,N_19762);
or U20320 (N_20320,N_19678,N_19878);
nand U20321 (N_20321,N_19707,N_19848);
xnor U20322 (N_20322,N_19881,N_19728);
nor U20323 (N_20323,N_19698,N_19905);
nor U20324 (N_20324,N_19528,N_19755);
and U20325 (N_20325,N_19548,N_19868);
xor U20326 (N_20326,N_19473,N_19461);
nor U20327 (N_20327,N_19799,N_19508);
nand U20328 (N_20328,N_19733,N_19485);
or U20329 (N_20329,N_19874,N_19659);
or U20330 (N_20330,N_19541,N_19942);
nor U20331 (N_20331,N_19756,N_19411);
nor U20332 (N_20332,N_19818,N_19558);
nor U20333 (N_20333,N_19540,N_19971);
nand U20334 (N_20334,N_19477,N_19482);
xor U20335 (N_20335,N_19866,N_19520);
nand U20336 (N_20336,N_19702,N_19898);
xor U20337 (N_20337,N_19557,N_19853);
xnor U20338 (N_20338,N_19606,N_19721);
nor U20339 (N_20339,N_19911,N_19452);
and U20340 (N_20340,N_19985,N_19716);
nand U20341 (N_20341,N_19800,N_19661);
and U20342 (N_20342,N_19616,N_19646);
and U20343 (N_20343,N_19837,N_19796);
nor U20344 (N_20344,N_19575,N_19491);
nand U20345 (N_20345,N_19433,N_19473);
nor U20346 (N_20346,N_19716,N_19587);
or U20347 (N_20347,N_19805,N_19995);
xnor U20348 (N_20348,N_19495,N_19940);
and U20349 (N_20349,N_19993,N_19955);
and U20350 (N_20350,N_19689,N_19775);
and U20351 (N_20351,N_19937,N_19792);
nand U20352 (N_20352,N_19909,N_19453);
or U20353 (N_20353,N_19581,N_19993);
and U20354 (N_20354,N_19384,N_19593);
or U20355 (N_20355,N_19770,N_19680);
nor U20356 (N_20356,N_19904,N_19527);
and U20357 (N_20357,N_19711,N_19825);
nor U20358 (N_20358,N_19561,N_19861);
and U20359 (N_20359,N_19444,N_19641);
or U20360 (N_20360,N_19794,N_19491);
and U20361 (N_20361,N_19986,N_19588);
nor U20362 (N_20362,N_19574,N_19410);
or U20363 (N_20363,N_19585,N_19837);
xnor U20364 (N_20364,N_19870,N_19437);
or U20365 (N_20365,N_19740,N_19807);
nor U20366 (N_20366,N_19501,N_19641);
or U20367 (N_20367,N_19913,N_19838);
nor U20368 (N_20368,N_19716,N_19618);
nor U20369 (N_20369,N_19904,N_19587);
nor U20370 (N_20370,N_19802,N_19538);
or U20371 (N_20371,N_19803,N_19404);
and U20372 (N_20372,N_19763,N_19845);
nor U20373 (N_20373,N_19951,N_19888);
and U20374 (N_20374,N_19423,N_19645);
or U20375 (N_20375,N_19976,N_19527);
nor U20376 (N_20376,N_19694,N_19556);
nand U20377 (N_20377,N_19748,N_19519);
nand U20378 (N_20378,N_19468,N_19516);
nor U20379 (N_20379,N_19564,N_19969);
nor U20380 (N_20380,N_19740,N_19867);
xor U20381 (N_20381,N_19684,N_19809);
or U20382 (N_20382,N_19728,N_19688);
and U20383 (N_20383,N_19764,N_19998);
nor U20384 (N_20384,N_19843,N_19542);
nor U20385 (N_20385,N_19822,N_19495);
nand U20386 (N_20386,N_19797,N_19647);
xor U20387 (N_20387,N_19400,N_19391);
or U20388 (N_20388,N_19503,N_19632);
nor U20389 (N_20389,N_19777,N_19451);
nor U20390 (N_20390,N_19515,N_19414);
nor U20391 (N_20391,N_19550,N_19464);
nor U20392 (N_20392,N_19796,N_19937);
and U20393 (N_20393,N_19872,N_19686);
nor U20394 (N_20394,N_19452,N_19800);
nand U20395 (N_20395,N_19990,N_19948);
xor U20396 (N_20396,N_19457,N_19640);
nand U20397 (N_20397,N_19643,N_19991);
or U20398 (N_20398,N_19760,N_19535);
nand U20399 (N_20399,N_19537,N_19967);
nor U20400 (N_20400,N_19779,N_19826);
nor U20401 (N_20401,N_19686,N_19664);
nand U20402 (N_20402,N_19806,N_19723);
or U20403 (N_20403,N_19674,N_19817);
or U20404 (N_20404,N_19575,N_19677);
or U20405 (N_20405,N_19427,N_19694);
and U20406 (N_20406,N_19852,N_19926);
xnor U20407 (N_20407,N_19485,N_19487);
nand U20408 (N_20408,N_19375,N_19671);
or U20409 (N_20409,N_19806,N_19444);
and U20410 (N_20410,N_19803,N_19876);
or U20411 (N_20411,N_19631,N_19982);
or U20412 (N_20412,N_19748,N_19816);
xor U20413 (N_20413,N_19949,N_19888);
or U20414 (N_20414,N_19475,N_19955);
nand U20415 (N_20415,N_19636,N_19579);
nand U20416 (N_20416,N_19807,N_19551);
and U20417 (N_20417,N_19526,N_19609);
or U20418 (N_20418,N_19471,N_19394);
or U20419 (N_20419,N_19978,N_19468);
nand U20420 (N_20420,N_19679,N_19670);
nor U20421 (N_20421,N_19937,N_19965);
nand U20422 (N_20422,N_19406,N_19897);
or U20423 (N_20423,N_19830,N_19590);
nand U20424 (N_20424,N_19784,N_19539);
nand U20425 (N_20425,N_19472,N_19715);
nand U20426 (N_20426,N_19758,N_19503);
or U20427 (N_20427,N_19827,N_19472);
and U20428 (N_20428,N_19726,N_19706);
xnor U20429 (N_20429,N_19910,N_19990);
nor U20430 (N_20430,N_19989,N_19865);
nor U20431 (N_20431,N_19825,N_19391);
nor U20432 (N_20432,N_19820,N_19514);
nor U20433 (N_20433,N_19589,N_19737);
and U20434 (N_20434,N_19653,N_19517);
nand U20435 (N_20435,N_19671,N_19813);
nand U20436 (N_20436,N_19452,N_19892);
or U20437 (N_20437,N_19825,N_19897);
nor U20438 (N_20438,N_19419,N_19740);
or U20439 (N_20439,N_19629,N_19455);
nor U20440 (N_20440,N_19574,N_19539);
nand U20441 (N_20441,N_19988,N_19724);
and U20442 (N_20442,N_19426,N_19677);
nand U20443 (N_20443,N_19890,N_19482);
nor U20444 (N_20444,N_19649,N_19581);
or U20445 (N_20445,N_19841,N_19476);
or U20446 (N_20446,N_19854,N_19414);
and U20447 (N_20447,N_19382,N_19588);
xor U20448 (N_20448,N_19864,N_19992);
or U20449 (N_20449,N_19832,N_19863);
nand U20450 (N_20450,N_19965,N_19618);
nor U20451 (N_20451,N_19695,N_19983);
or U20452 (N_20452,N_19459,N_19932);
and U20453 (N_20453,N_19387,N_19958);
nor U20454 (N_20454,N_19390,N_19474);
and U20455 (N_20455,N_19727,N_19625);
and U20456 (N_20456,N_19539,N_19602);
and U20457 (N_20457,N_19753,N_19565);
nand U20458 (N_20458,N_19784,N_19972);
nand U20459 (N_20459,N_19718,N_19475);
nor U20460 (N_20460,N_19470,N_19887);
nand U20461 (N_20461,N_19659,N_19831);
nor U20462 (N_20462,N_19611,N_19755);
or U20463 (N_20463,N_19690,N_19849);
nor U20464 (N_20464,N_19610,N_19731);
nor U20465 (N_20465,N_19445,N_19468);
xnor U20466 (N_20466,N_19436,N_19831);
nor U20467 (N_20467,N_19966,N_19813);
or U20468 (N_20468,N_19580,N_19425);
nor U20469 (N_20469,N_19559,N_19407);
xnor U20470 (N_20470,N_19639,N_19861);
nand U20471 (N_20471,N_19965,N_19655);
nand U20472 (N_20472,N_19918,N_19382);
nor U20473 (N_20473,N_19715,N_19663);
nor U20474 (N_20474,N_19824,N_19873);
nand U20475 (N_20475,N_19904,N_19845);
nor U20476 (N_20476,N_19410,N_19455);
nand U20477 (N_20477,N_19740,N_19575);
and U20478 (N_20478,N_19601,N_19943);
xor U20479 (N_20479,N_19628,N_19479);
or U20480 (N_20480,N_19837,N_19501);
xnor U20481 (N_20481,N_19467,N_19519);
xnor U20482 (N_20482,N_19896,N_19818);
nor U20483 (N_20483,N_19720,N_19604);
xor U20484 (N_20484,N_19948,N_19410);
and U20485 (N_20485,N_19375,N_19906);
and U20486 (N_20486,N_19388,N_19390);
or U20487 (N_20487,N_19483,N_19836);
or U20488 (N_20488,N_19533,N_19991);
nand U20489 (N_20489,N_19667,N_19621);
xor U20490 (N_20490,N_19430,N_19925);
or U20491 (N_20491,N_19744,N_19708);
nor U20492 (N_20492,N_19593,N_19873);
nand U20493 (N_20493,N_19480,N_19651);
xnor U20494 (N_20494,N_19553,N_19725);
nor U20495 (N_20495,N_19411,N_19612);
nor U20496 (N_20496,N_19790,N_19454);
nor U20497 (N_20497,N_19452,N_19818);
nor U20498 (N_20498,N_19937,N_19919);
or U20499 (N_20499,N_19850,N_19691);
nor U20500 (N_20500,N_19825,N_19502);
or U20501 (N_20501,N_19650,N_19508);
nand U20502 (N_20502,N_19975,N_19950);
nand U20503 (N_20503,N_19672,N_19532);
nor U20504 (N_20504,N_19388,N_19959);
and U20505 (N_20505,N_19682,N_19557);
or U20506 (N_20506,N_19763,N_19750);
and U20507 (N_20507,N_19829,N_19982);
xnor U20508 (N_20508,N_19549,N_19626);
or U20509 (N_20509,N_19445,N_19572);
nand U20510 (N_20510,N_19913,N_19732);
nand U20511 (N_20511,N_19964,N_19653);
nand U20512 (N_20512,N_19446,N_19707);
nand U20513 (N_20513,N_19428,N_19735);
nor U20514 (N_20514,N_19639,N_19590);
and U20515 (N_20515,N_19822,N_19928);
or U20516 (N_20516,N_19782,N_19552);
nor U20517 (N_20517,N_19577,N_19460);
and U20518 (N_20518,N_19997,N_19795);
nor U20519 (N_20519,N_19437,N_19947);
and U20520 (N_20520,N_19576,N_19679);
and U20521 (N_20521,N_19665,N_19970);
or U20522 (N_20522,N_19711,N_19846);
xor U20523 (N_20523,N_19986,N_19505);
nand U20524 (N_20524,N_19916,N_19712);
nor U20525 (N_20525,N_19701,N_19780);
xnor U20526 (N_20526,N_19492,N_19734);
nand U20527 (N_20527,N_19527,N_19855);
or U20528 (N_20528,N_19687,N_19749);
nor U20529 (N_20529,N_19423,N_19675);
xnor U20530 (N_20530,N_19687,N_19710);
nor U20531 (N_20531,N_19660,N_19528);
nor U20532 (N_20532,N_19432,N_19424);
nand U20533 (N_20533,N_19473,N_19928);
xnor U20534 (N_20534,N_19567,N_19746);
xor U20535 (N_20535,N_19602,N_19408);
and U20536 (N_20536,N_19633,N_19412);
and U20537 (N_20537,N_19733,N_19511);
or U20538 (N_20538,N_19775,N_19941);
nor U20539 (N_20539,N_19761,N_19951);
nor U20540 (N_20540,N_19718,N_19620);
nand U20541 (N_20541,N_19877,N_19385);
nand U20542 (N_20542,N_19838,N_19999);
or U20543 (N_20543,N_19740,N_19782);
nand U20544 (N_20544,N_19488,N_19821);
xnor U20545 (N_20545,N_19641,N_19975);
or U20546 (N_20546,N_19470,N_19432);
or U20547 (N_20547,N_19890,N_19980);
or U20548 (N_20548,N_19520,N_19851);
or U20549 (N_20549,N_19546,N_19432);
and U20550 (N_20550,N_19997,N_19951);
nor U20551 (N_20551,N_19649,N_19744);
or U20552 (N_20552,N_19411,N_19523);
nor U20553 (N_20553,N_19923,N_19546);
or U20554 (N_20554,N_19696,N_19753);
or U20555 (N_20555,N_19658,N_19478);
or U20556 (N_20556,N_19723,N_19598);
or U20557 (N_20557,N_19743,N_19706);
xor U20558 (N_20558,N_19487,N_19601);
nor U20559 (N_20559,N_19569,N_19698);
or U20560 (N_20560,N_19636,N_19394);
and U20561 (N_20561,N_19412,N_19835);
nand U20562 (N_20562,N_19798,N_19910);
nand U20563 (N_20563,N_19553,N_19526);
nand U20564 (N_20564,N_19998,N_19531);
and U20565 (N_20565,N_19708,N_19701);
xor U20566 (N_20566,N_19406,N_19837);
nand U20567 (N_20567,N_19834,N_19477);
and U20568 (N_20568,N_19874,N_19429);
and U20569 (N_20569,N_19973,N_19844);
and U20570 (N_20570,N_19567,N_19627);
and U20571 (N_20571,N_19705,N_19409);
and U20572 (N_20572,N_19745,N_19532);
or U20573 (N_20573,N_19386,N_19773);
xnor U20574 (N_20574,N_19727,N_19499);
and U20575 (N_20575,N_19893,N_19864);
and U20576 (N_20576,N_19386,N_19589);
nor U20577 (N_20577,N_19921,N_19595);
nor U20578 (N_20578,N_19566,N_19641);
and U20579 (N_20579,N_19830,N_19885);
and U20580 (N_20580,N_19456,N_19822);
nand U20581 (N_20581,N_19774,N_19589);
and U20582 (N_20582,N_19966,N_19685);
nand U20583 (N_20583,N_19596,N_19704);
nor U20584 (N_20584,N_19607,N_19659);
nand U20585 (N_20585,N_19775,N_19424);
and U20586 (N_20586,N_19713,N_19773);
nor U20587 (N_20587,N_19684,N_19489);
and U20588 (N_20588,N_19585,N_19420);
nand U20589 (N_20589,N_19523,N_19481);
and U20590 (N_20590,N_19799,N_19641);
or U20591 (N_20591,N_19770,N_19529);
and U20592 (N_20592,N_19925,N_19766);
or U20593 (N_20593,N_19395,N_19430);
and U20594 (N_20594,N_19485,N_19685);
or U20595 (N_20595,N_19638,N_19836);
nor U20596 (N_20596,N_19750,N_19917);
nand U20597 (N_20597,N_19395,N_19798);
and U20598 (N_20598,N_19377,N_19699);
nor U20599 (N_20599,N_19640,N_19382);
and U20600 (N_20600,N_19695,N_19991);
and U20601 (N_20601,N_19761,N_19856);
nand U20602 (N_20602,N_19954,N_19599);
nand U20603 (N_20603,N_19643,N_19671);
nand U20604 (N_20604,N_19925,N_19931);
or U20605 (N_20605,N_19518,N_19911);
and U20606 (N_20606,N_19571,N_19605);
and U20607 (N_20607,N_19935,N_19815);
and U20608 (N_20608,N_19501,N_19444);
or U20609 (N_20609,N_19773,N_19436);
nand U20610 (N_20610,N_19522,N_19976);
nand U20611 (N_20611,N_19384,N_19944);
nand U20612 (N_20612,N_19890,N_19681);
xnor U20613 (N_20613,N_19611,N_19960);
nand U20614 (N_20614,N_19536,N_19831);
xnor U20615 (N_20615,N_19989,N_19497);
and U20616 (N_20616,N_19979,N_19526);
nor U20617 (N_20617,N_19505,N_19700);
nand U20618 (N_20618,N_19878,N_19483);
nor U20619 (N_20619,N_19598,N_19540);
nor U20620 (N_20620,N_19723,N_19962);
nand U20621 (N_20621,N_19741,N_19525);
nand U20622 (N_20622,N_19738,N_19510);
nor U20623 (N_20623,N_19453,N_19598);
nand U20624 (N_20624,N_19476,N_19932);
and U20625 (N_20625,N_20217,N_20559);
or U20626 (N_20626,N_20382,N_20482);
or U20627 (N_20627,N_20246,N_20289);
and U20628 (N_20628,N_20140,N_20132);
nand U20629 (N_20629,N_20238,N_20104);
and U20630 (N_20630,N_20001,N_20307);
and U20631 (N_20631,N_20254,N_20204);
nor U20632 (N_20632,N_20506,N_20274);
nor U20633 (N_20633,N_20038,N_20061);
or U20634 (N_20634,N_20519,N_20481);
xor U20635 (N_20635,N_20281,N_20549);
or U20636 (N_20636,N_20213,N_20265);
xor U20637 (N_20637,N_20521,N_20465);
and U20638 (N_20638,N_20545,N_20362);
nor U20639 (N_20639,N_20435,N_20497);
xor U20640 (N_20640,N_20157,N_20210);
or U20641 (N_20641,N_20496,N_20169);
xnor U20642 (N_20642,N_20242,N_20313);
nand U20643 (N_20643,N_20244,N_20224);
and U20644 (N_20644,N_20056,N_20294);
nand U20645 (N_20645,N_20308,N_20413);
nand U20646 (N_20646,N_20417,N_20615);
nand U20647 (N_20647,N_20309,N_20427);
nor U20648 (N_20648,N_20196,N_20145);
nand U20649 (N_20649,N_20415,N_20105);
nor U20650 (N_20650,N_20037,N_20245);
or U20651 (N_20651,N_20490,N_20152);
or U20652 (N_20652,N_20447,N_20315);
or U20653 (N_20653,N_20511,N_20151);
nor U20654 (N_20654,N_20555,N_20248);
and U20655 (N_20655,N_20174,N_20120);
nand U20656 (N_20656,N_20541,N_20453);
nor U20657 (N_20657,N_20408,N_20109);
xor U20658 (N_20658,N_20601,N_20259);
nand U20659 (N_20659,N_20445,N_20161);
xor U20660 (N_20660,N_20147,N_20434);
nor U20661 (N_20661,N_20030,N_20319);
or U20662 (N_20662,N_20581,N_20112);
and U20663 (N_20663,N_20525,N_20546);
and U20664 (N_20664,N_20304,N_20373);
nor U20665 (N_20665,N_20084,N_20488);
nor U20666 (N_20666,N_20070,N_20032);
nand U20667 (N_20667,N_20192,N_20341);
nor U20668 (N_20668,N_20428,N_20197);
nor U20669 (N_20669,N_20436,N_20438);
nand U20670 (N_20670,N_20252,N_20047);
nand U20671 (N_20671,N_20457,N_20522);
nor U20672 (N_20672,N_20303,N_20595);
or U20673 (N_20673,N_20097,N_20227);
nand U20674 (N_20674,N_20071,N_20214);
and U20675 (N_20675,N_20005,N_20396);
or U20676 (N_20676,N_20473,N_20237);
or U20677 (N_20677,N_20524,N_20321);
and U20678 (N_20678,N_20149,N_20311);
or U20679 (N_20679,N_20059,N_20574);
xnor U20680 (N_20680,N_20386,N_20069);
or U20681 (N_20681,N_20023,N_20166);
nor U20682 (N_20682,N_20229,N_20159);
nor U20683 (N_20683,N_20279,N_20552);
nor U20684 (N_20684,N_20374,N_20221);
or U20685 (N_20685,N_20528,N_20134);
or U20686 (N_20686,N_20062,N_20337);
nand U20687 (N_20687,N_20580,N_20006);
nand U20688 (N_20688,N_20195,N_20357);
nor U20689 (N_20689,N_20587,N_20225);
and U20690 (N_20690,N_20578,N_20532);
nand U20691 (N_20691,N_20586,N_20123);
nor U20692 (N_20692,N_20589,N_20489);
xor U20693 (N_20693,N_20012,N_20460);
and U20694 (N_20694,N_20098,N_20518);
or U20695 (N_20695,N_20461,N_20544);
or U20696 (N_20696,N_20010,N_20291);
nor U20697 (N_20697,N_20613,N_20472);
or U20698 (N_20698,N_20231,N_20573);
or U20699 (N_20699,N_20409,N_20218);
or U20700 (N_20700,N_20364,N_20397);
and U20701 (N_20701,N_20222,N_20464);
nor U20702 (N_20702,N_20422,N_20558);
nor U20703 (N_20703,N_20366,N_20385);
and U20704 (N_20704,N_20493,N_20329);
nor U20705 (N_20705,N_20085,N_20517);
and U20706 (N_20706,N_20407,N_20380);
nand U20707 (N_20707,N_20604,N_20264);
nand U20708 (N_20708,N_20015,N_20442);
nor U20709 (N_20709,N_20526,N_20475);
and U20710 (N_20710,N_20219,N_20534);
and U20711 (N_20711,N_20345,N_20563);
nand U20712 (N_20712,N_20441,N_20343);
or U20713 (N_20713,N_20096,N_20361);
and U20714 (N_20714,N_20561,N_20326);
or U20715 (N_20715,N_20505,N_20371);
nand U20716 (N_20716,N_20004,N_20448);
nor U20717 (N_20717,N_20250,N_20141);
xor U20718 (N_20718,N_20027,N_20236);
or U20719 (N_20719,N_20554,N_20451);
nor U20720 (N_20720,N_20124,N_20455);
and U20721 (N_20721,N_20216,N_20398);
nor U20722 (N_20722,N_20117,N_20597);
xor U20723 (N_20723,N_20256,N_20223);
or U20724 (N_20724,N_20606,N_20257);
xnor U20725 (N_20725,N_20175,N_20530);
nor U20726 (N_20726,N_20280,N_20111);
nor U20727 (N_20727,N_20463,N_20450);
nor U20728 (N_20728,N_20146,N_20179);
nand U20729 (N_20729,N_20094,N_20144);
or U20730 (N_20730,N_20351,N_20241);
nor U20731 (N_20731,N_20261,N_20235);
and U20732 (N_20732,N_20278,N_20619);
nor U20733 (N_20733,N_20116,N_20452);
and U20734 (N_20734,N_20154,N_20440);
nand U20735 (N_20735,N_20499,N_20390);
nor U20736 (N_20736,N_20103,N_20080);
nor U20737 (N_20737,N_20480,N_20082);
xor U20738 (N_20738,N_20042,N_20334);
or U20739 (N_20739,N_20287,N_20553);
and U20740 (N_20740,N_20599,N_20108);
and U20741 (N_20741,N_20429,N_20336);
and U20742 (N_20742,N_20058,N_20318);
and U20743 (N_20743,N_20421,N_20483);
xnor U20744 (N_20744,N_20317,N_20028);
or U20745 (N_20745,N_20286,N_20536);
xor U20746 (N_20746,N_20305,N_20439);
nand U20747 (N_20747,N_20026,N_20014);
or U20748 (N_20748,N_20076,N_20471);
and U20749 (N_20749,N_20158,N_20133);
or U20750 (N_20750,N_20168,N_20199);
or U20751 (N_20751,N_20583,N_20470);
or U20752 (N_20752,N_20310,N_20228);
or U20753 (N_20753,N_20618,N_20063);
nor U20754 (N_20754,N_20101,N_20614);
or U20755 (N_20755,N_20065,N_20127);
xor U20756 (N_20756,N_20412,N_20608);
nor U20757 (N_20757,N_20515,N_20255);
nor U20758 (N_20758,N_20295,N_20509);
nand U20759 (N_20759,N_20284,N_20090);
nand U20760 (N_20760,N_20234,N_20314);
and U20761 (N_20761,N_20469,N_20339);
and U20762 (N_20762,N_20399,N_20535);
xor U20763 (N_20763,N_20571,N_20359);
nor U20764 (N_20764,N_20567,N_20383);
or U20765 (N_20765,N_20239,N_20406);
nor U20766 (N_20766,N_20263,N_20495);
and U20767 (N_20767,N_20083,N_20122);
and U20768 (N_20768,N_20494,N_20538);
nor U20769 (N_20769,N_20403,N_20138);
nor U20770 (N_20770,N_20107,N_20388);
or U20771 (N_20771,N_20560,N_20142);
and U20772 (N_20772,N_20297,N_20548);
and U20773 (N_20773,N_20603,N_20332);
and U20774 (N_20774,N_20075,N_20054);
and U20775 (N_20775,N_20432,N_20277);
xnor U20776 (N_20776,N_20491,N_20593);
or U20777 (N_20777,N_20500,N_20520);
or U20778 (N_20778,N_20160,N_20596);
nor U20779 (N_20779,N_20365,N_20106);
nand U20780 (N_20780,N_20017,N_20089);
and U20781 (N_20781,N_20007,N_20272);
and U20782 (N_20782,N_20299,N_20610);
or U20783 (N_20783,N_20016,N_20379);
or U20784 (N_20784,N_20503,N_20135);
or U20785 (N_20785,N_20184,N_20346);
nor U20786 (N_20786,N_20207,N_20331);
nor U20787 (N_20787,N_20527,N_20323);
nand U20788 (N_20788,N_20095,N_20164);
nand U20789 (N_20789,N_20130,N_20600);
xor U20790 (N_20790,N_20565,N_20201);
and U20791 (N_20791,N_20300,N_20232);
nand U20792 (N_20792,N_20011,N_20301);
and U20793 (N_20793,N_20392,N_20024);
nor U20794 (N_20794,N_20173,N_20260);
or U20795 (N_20795,N_20582,N_20577);
or U20796 (N_20796,N_20121,N_20542);
and U20797 (N_20797,N_20276,N_20370);
and U20798 (N_20798,N_20352,N_20088);
and U20799 (N_20799,N_20044,N_20043);
nand U20800 (N_20800,N_20181,N_20302);
xor U20801 (N_20801,N_20414,N_20372);
nor U20802 (N_20802,N_20437,N_20285);
and U20803 (N_20803,N_20202,N_20191);
nand U20804 (N_20804,N_20325,N_20592);
nand U20805 (N_20805,N_20431,N_20347);
and U20806 (N_20806,N_20609,N_20607);
nor U20807 (N_20807,N_20150,N_20139);
and U20808 (N_20808,N_20008,N_20588);
nand U20809 (N_20809,N_20344,N_20510);
nor U20810 (N_20810,N_20153,N_20189);
or U20811 (N_20811,N_20208,N_20529);
and U20812 (N_20812,N_20267,N_20477);
nand U20813 (N_20813,N_20594,N_20029);
nand U20814 (N_20814,N_20622,N_20531);
nand U20815 (N_20815,N_20114,N_20226);
nor U20816 (N_20816,N_20020,N_20367);
nand U20817 (N_20817,N_20590,N_20046);
and U20818 (N_20818,N_20035,N_20576);
nand U20819 (N_20819,N_20355,N_20547);
and U20820 (N_20820,N_20376,N_20176);
xnor U20821 (N_20821,N_20262,N_20420);
nand U20822 (N_20822,N_20049,N_20353);
xor U20823 (N_20823,N_20551,N_20391);
or U20824 (N_20824,N_20087,N_20335);
or U20825 (N_20825,N_20591,N_20467);
nor U20826 (N_20826,N_20602,N_20411);
or U20827 (N_20827,N_20093,N_20220);
nor U20828 (N_20828,N_20312,N_20516);
or U20829 (N_20829,N_20419,N_20572);
and U20830 (N_20830,N_20324,N_20200);
nor U20831 (N_20831,N_20078,N_20557);
nor U20832 (N_20832,N_20079,N_20212);
xor U20833 (N_20833,N_20474,N_20404);
nor U20834 (N_20834,N_20570,N_20400);
nand U20835 (N_20835,N_20433,N_20290);
or U20836 (N_20836,N_20183,N_20129);
or U20837 (N_20837,N_20115,N_20350);
nor U20838 (N_20838,N_20584,N_20416);
and U20839 (N_20839,N_20206,N_20394);
nor U20840 (N_20840,N_20426,N_20501);
and U20841 (N_20841,N_20185,N_20378);
nor U20842 (N_20842,N_20193,N_20498);
xnor U20843 (N_20843,N_20479,N_20100);
or U20844 (N_20844,N_20623,N_20556);
or U20845 (N_20845,N_20136,N_20230);
or U20846 (N_20846,N_20025,N_20033);
nand U20847 (N_20847,N_20569,N_20036);
nand U20848 (N_20848,N_20045,N_20502);
and U20849 (N_20849,N_20233,N_20292);
nor U20850 (N_20850,N_20612,N_20209);
and U20851 (N_20851,N_20354,N_20395);
nor U20852 (N_20852,N_20333,N_20377);
and U20853 (N_20853,N_20002,N_20349);
nand U20854 (N_20854,N_20617,N_20266);
nor U20855 (N_20855,N_20102,N_20211);
xnor U20856 (N_20856,N_20031,N_20092);
nand U20857 (N_20857,N_20253,N_20268);
xor U20858 (N_20858,N_20050,N_20128);
nand U20859 (N_20859,N_20430,N_20198);
or U20860 (N_20860,N_20550,N_20454);
nor U20861 (N_20861,N_20073,N_20443);
and U20862 (N_20862,N_20459,N_20468);
nand U20863 (N_20863,N_20320,N_20533);
nand U20864 (N_20864,N_20180,N_20393);
nor U20865 (N_20865,N_20485,N_20249);
or U20866 (N_20866,N_20585,N_20539);
and U20867 (N_20867,N_20369,N_20171);
nor U20868 (N_20868,N_20476,N_20401);
nor U20869 (N_20869,N_20271,N_20446);
nor U20870 (N_20870,N_20039,N_20052);
xnor U20871 (N_20871,N_20003,N_20040);
nand U20872 (N_20872,N_20243,N_20456);
or U20873 (N_20873,N_20099,N_20188);
and U20874 (N_20874,N_20172,N_20537);
nor U20875 (N_20875,N_20186,N_20270);
nor U20876 (N_20876,N_20381,N_20621);
xnor U20877 (N_20877,N_20358,N_20484);
nand U20878 (N_20878,N_20616,N_20512);
and U20879 (N_20879,N_20620,N_20110);
or U20880 (N_20880,N_20247,N_20269);
and U20881 (N_20881,N_20118,N_20275);
nand U20882 (N_20882,N_20306,N_20148);
and U20883 (N_20883,N_20540,N_20055);
nor U20884 (N_20884,N_20338,N_20478);
nand U20885 (N_20885,N_20077,N_20330);
nor U20886 (N_20886,N_20282,N_20605);
and U20887 (N_20887,N_20203,N_20327);
or U20888 (N_20888,N_20126,N_20579);
xor U20889 (N_20889,N_20598,N_20187);
and U20890 (N_20890,N_20492,N_20298);
or U20891 (N_20891,N_20523,N_20156);
nand U20892 (N_20892,N_20125,N_20283);
nand U20893 (N_20893,N_20182,N_20064);
and U20894 (N_20894,N_20273,N_20424);
and U20895 (N_20895,N_20190,N_20205);
or U20896 (N_20896,N_20564,N_20562);
and U20897 (N_20897,N_20258,N_20177);
nor U20898 (N_20898,N_20387,N_20155);
or U20899 (N_20899,N_20018,N_20009);
nand U20900 (N_20900,N_20389,N_20514);
and U20901 (N_20901,N_20458,N_20170);
xnor U20902 (N_20902,N_20167,N_20402);
nand U20903 (N_20903,N_20425,N_20444);
nand U20904 (N_20904,N_20487,N_20322);
or U20905 (N_20905,N_20360,N_20066);
or U20906 (N_20906,N_20566,N_20328);
or U20907 (N_20907,N_20057,N_20081);
nor U20908 (N_20908,N_20178,N_20068);
nand U20909 (N_20909,N_20296,N_20067);
nor U20910 (N_20910,N_20363,N_20624);
nand U20911 (N_20911,N_20215,N_20060);
and U20912 (N_20912,N_20410,N_20507);
or U20913 (N_20913,N_20288,N_20513);
nor U20914 (N_20914,N_20074,N_20048);
nand U20915 (N_20915,N_20163,N_20143);
and U20916 (N_20916,N_20013,N_20486);
nand U20917 (N_20917,N_20568,N_20449);
nand U20918 (N_20918,N_20022,N_20356);
nor U20919 (N_20919,N_20131,N_20041);
and U20920 (N_20920,N_20405,N_20340);
and U20921 (N_20921,N_20113,N_20119);
and U20922 (N_20922,N_20368,N_20053);
nand U20923 (N_20923,N_20423,N_20034);
or U20924 (N_20924,N_20000,N_20251);
and U20925 (N_20925,N_20019,N_20316);
nand U20926 (N_20926,N_20021,N_20086);
nand U20927 (N_20927,N_20091,N_20342);
and U20928 (N_20928,N_20293,N_20543);
nor U20929 (N_20929,N_20508,N_20165);
nor U20930 (N_20930,N_20611,N_20194);
nor U20931 (N_20931,N_20072,N_20462);
and U20932 (N_20932,N_20240,N_20575);
or U20933 (N_20933,N_20348,N_20375);
xnor U20934 (N_20934,N_20051,N_20162);
nand U20935 (N_20935,N_20504,N_20466);
or U20936 (N_20936,N_20137,N_20418);
nor U20937 (N_20937,N_20384,N_20408);
or U20938 (N_20938,N_20425,N_20295);
nand U20939 (N_20939,N_20258,N_20573);
or U20940 (N_20940,N_20531,N_20511);
or U20941 (N_20941,N_20250,N_20108);
or U20942 (N_20942,N_20189,N_20043);
nand U20943 (N_20943,N_20515,N_20060);
nand U20944 (N_20944,N_20133,N_20202);
or U20945 (N_20945,N_20194,N_20313);
nor U20946 (N_20946,N_20468,N_20290);
nor U20947 (N_20947,N_20328,N_20331);
or U20948 (N_20948,N_20279,N_20381);
nand U20949 (N_20949,N_20619,N_20400);
or U20950 (N_20950,N_20147,N_20038);
or U20951 (N_20951,N_20269,N_20101);
xnor U20952 (N_20952,N_20238,N_20216);
and U20953 (N_20953,N_20410,N_20148);
nand U20954 (N_20954,N_20035,N_20131);
nand U20955 (N_20955,N_20134,N_20468);
xnor U20956 (N_20956,N_20092,N_20568);
nor U20957 (N_20957,N_20429,N_20500);
and U20958 (N_20958,N_20422,N_20098);
nor U20959 (N_20959,N_20430,N_20591);
nor U20960 (N_20960,N_20270,N_20132);
xor U20961 (N_20961,N_20433,N_20304);
nor U20962 (N_20962,N_20005,N_20203);
and U20963 (N_20963,N_20493,N_20135);
nand U20964 (N_20964,N_20512,N_20275);
nor U20965 (N_20965,N_20288,N_20417);
xor U20966 (N_20966,N_20055,N_20147);
or U20967 (N_20967,N_20171,N_20463);
nand U20968 (N_20968,N_20039,N_20473);
nand U20969 (N_20969,N_20071,N_20367);
xor U20970 (N_20970,N_20085,N_20098);
or U20971 (N_20971,N_20570,N_20616);
nor U20972 (N_20972,N_20006,N_20194);
and U20973 (N_20973,N_20021,N_20425);
and U20974 (N_20974,N_20619,N_20533);
or U20975 (N_20975,N_20379,N_20606);
xnor U20976 (N_20976,N_20322,N_20283);
xnor U20977 (N_20977,N_20280,N_20412);
xnor U20978 (N_20978,N_20525,N_20176);
or U20979 (N_20979,N_20462,N_20028);
and U20980 (N_20980,N_20151,N_20594);
or U20981 (N_20981,N_20456,N_20506);
xnor U20982 (N_20982,N_20527,N_20446);
nor U20983 (N_20983,N_20621,N_20239);
nand U20984 (N_20984,N_20406,N_20071);
or U20985 (N_20985,N_20415,N_20110);
nand U20986 (N_20986,N_20370,N_20620);
or U20987 (N_20987,N_20554,N_20281);
nor U20988 (N_20988,N_20425,N_20502);
or U20989 (N_20989,N_20447,N_20427);
and U20990 (N_20990,N_20259,N_20435);
or U20991 (N_20991,N_20319,N_20171);
nand U20992 (N_20992,N_20333,N_20116);
nor U20993 (N_20993,N_20087,N_20245);
and U20994 (N_20994,N_20014,N_20357);
nor U20995 (N_20995,N_20274,N_20416);
or U20996 (N_20996,N_20136,N_20444);
and U20997 (N_20997,N_20504,N_20253);
or U20998 (N_20998,N_20405,N_20503);
nor U20999 (N_20999,N_20053,N_20285);
nand U21000 (N_21000,N_20488,N_20549);
xor U21001 (N_21001,N_20220,N_20477);
or U21002 (N_21002,N_20376,N_20562);
nand U21003 (N_21003,N_20079,N_20570);
nand U21004 (N_21004,N_20402,N_20307);
xor U21005 (N_21005,N_20156,N_20493);
nor U21006 (N_21006,N_20185,N_20067);
nor U21007 (N_21007,N_20306,N_20106);
nor U21008 (N_21008,N_20569,N_20593);
and U21009 (N_21009,N_20101,N_20257);
and U21010 (N_21010,N_20002,N_20583);
nor U21011 (N_21011,N_20455,N_20081);
xnor U21012 (N_21012,N_20512,N_20012);
or U21013 (N_21013,N_20075,N_20515);
or U21014 (N_21014,N_20571,N_20072);
xor U21015 (N_21015,N_20599,N_20123);
nor U21016 (N_21016,N_20486,N_20498);
nand U21017 (N_21017,N_20114,N_20393);
nor U21018 (N_21018,N_20075,N_20525);
or U21019 (N_21019,N_20590,N_20415);
or U21020 (N_21020,N_20536,N_20482);
nor U21021 (N_21021,N_20162,N_20221);
and U21022 (N_21022,N_20354,N_20608);
nor U21023 (N_21023,N_20421,N_20197);
nand U21024 (N_21024,N_20248,N_20061);
nand U21025 (N_21025,N_20135,N_20069);
xor U21026 (N_21026,N_20245,N_20166);
nand U21027 (N_21027,N_20488,N_20241);
and U21028 (N_21028,N_20463,N_20558);
nand U21029 (N_21029,N_20264,N_20160);
and U21030 (N_21030,N_20586,N_20503);
and U21031 (N_21031,N_20127,N_20152);
and U21032 (N_21032,N_20204,N_20209);
or U21033 (N_21033,N_20405,N_20596);
xor U21034 (N_21034,N_20119,N_20050);
or U21035 (N_21035,N_20622,N_20146);
or U21036 (N_21036,N_20206,N_20336);
nor U21037 (N_21037,N_20592,N_20190);
nor U21038 (N_21038,N_20233,N_20317);
nand U21039 (N_21039,N_20212,N_20125);
or U21040 (N_21040,N_20240,N_20596);
nand U21041 (N_21041,N_20374,N_20231);
nand U21042 (N_21042,N_20151,N_20569);
nor U21043 (N_21043,N_20118,N_20060);
nand U21044 (N_21044,N_20061,N_20537);
nand U21045 (N_21045,N_20501,N_20399);
nor U21046 (N_21046,N_20270,N_20437);
xor U21047 (N_21047,N_20456,N_20071);
or U21048 (N_21048,N_20227,N_20090);
nor U21049 (N_21049,N_20309,N_20408);
xor U21050 (N_21050,N_20301,N_20117);
and U21051 (N_21051,N_20462,N_20113);
xnor U21052 (N_21052,N_20116,N_20038);
nor U21053 (N_21053,N_20422,N_20451);
nor U21054 (N_21054,N_20204,N_20494);
and U21055 (N_21055,N_20069,N_20227);
and U21056 (N_21056,N_20225,N_20488);
xnor U21057 (N_21057,N_20277,N_20040);
xnor U21058 (N_21058,N_20358,N_20146);
nor U21059 (N_21059,N_20122,N_20497);
nand U21060 (N_21060,N_20266,N_20535);
nand U21061 (N_21061,N_20300,N_20413);
nor U21062 (N_21062,N_20184,N_20442);
nor U21063 (N_21063,N_20039,N_20503);
nand U21064 (N_21064,N_20530,N_20270);
or U21065 (N_21065,N_20550,N_20028);
and U21066 (N_21066,N_20076,N_20138);
nor U21067 (N_21067,N_20366,N_20151);
or U21068 (N_21068,N_20124,N_20607);
or U21069 (N_21069,N_20423,N_20523);
and U21070 (N_21070,N_20395,N_20505);
and U21071 (N_21071,N_20500,N_20064);
and U21072 (N_21072,N_20465,N_20514);
nand U21073 (N_21073,N_20043,N_20127);
or U21074 (N_21074,N_20446,N_20177);
nor U21075 (N_21075,N_20023,N_20560);
or U21076 (N_21076,N_20003,N_20180);
nand U21077 (N_21077,N_20318,N_20169);
and U21078 (N_21078,N_20394,N_20465);
and U21079 (N_21079,N_20501,N_20447);
and U21080 (N_21080,N_20103,N_20548);
and U21081 (N_21081,N_20299,N_20543);
nand U21082 (N_21082,N_20455,N_20532);
and U21083 (N_21083,N_20080,N_20150);
and U21084 (N_21084,N_20170,N_20044);
nor U21085 (N_21085,N_20220,N_20058);
nor U21086 (N_21086,N_20460,N_20306);
xnor U21087 (N_21087,N_20193,N_20349);
and U21088 (N_21088,N_20549,N_20391);
and U21089 (N_21089,N_20495,N_20082);
nor U21090 (N_21090,N_20030,N_20365);
or U21091 (N_21091,N_20366,N_20063);
or U21092 (N_21092,N_20442,N_20406);
nand U21093 (N_21093,N_20587,N_20320);
or U21094 (N_21094,N_20484,N_20619);
and U21095 (N_21095,N_20519,N_20030);
nor U21096 (N_21096,N_20277,N_20455);
nand U21097 (N_21097,N_20208,N_20272);
and U21098 (N_21098,N_20202,N_20573);
xor U21099 (N_21099,N_20440,N_20362);
or U21100 (N_21100,N_20528,N_20261);
or U21101 (N_21101,N_20560,N_20121);
and U21102 (N_21102,N_20574,N_20021);
and U21103 (N_21103,N_20017,N_20040);
or U21104 (N_21104,N_20334,N_20223);
or U21105 (N_21105,N_20066,N_20093);
and U21106 (N_21106,N_20569,N_20279);
or U21107 (N_21107,N_20554,N_20254);
nand U21108 (N_21108,N_20325,N_20447);
nor U21109 (N_21109,N_20335,N_20570);
nor U21110 (N_21110,N_20292,N_20243);
and U21111 (N_21111,N_20088,N_20262);
and U21112 (N_21112,N_20181,N_20433);
nand U21113 (N_21113,N_20461,N_20538);
or U21114 (N_21114,N_20555,N_20338);
and U21115 (N_21115,N_20472,N_20306);
xor U21116 (N_21116,N_20296,N_20397);
and U21117 (N_21117,N_20611,N_20060);
and U21118 (N_21118,N_20290,N_20214);
and U21119 (N_21119,N_20244,N_20354);
nand U21120 (N_21120,N_20122,N_20594);
and U21121 (N_21121,N_20270,N_20197);
xor U21122 (N_21122,N_20061,N_20479);
or U21123 (N_21123,N_20242,N_20344);
nand U21124 (N_21124,N_20109,N_20397);
and U21125 (N_21125,N_20389,N_20252);
and U21126 (N_21126,N_20361,N_20597);
xor U21127 (N_21127,N_20441,N_20022);
nand U21128 (N_21128,N_20217,N_20103);
or U21129 (N_21129,N_20463,N_20179);
nor U21130 (N_21130,N_20498,N_20460);
and U21131 (N_21131,N_20498,N_20600);
nand U21132 (N_21132,N_20374,N_20081);
nor U21133 (N_21133,N_20029,N_20621);
nand U21134 (N_21134,N_20044,N_20234);
xnor U21135 (N_21135,N_20561,N_20282);
nor U21136 (N_21136,N_20231,N_20365);
or U21137 (N_21137,N_20512,N_20476);
and U21138 (N_21138,N_20113,N_20114);
nand U21139 (N_21139,N_20199,N_20130);
or U21140 (N_21140,N_20280,N_20404);
nand U21141 (N_21141,N_20587,N_20488);
nand U21142 (N_21142,N_20002,N_20298);
nor U21143 (N_21143,N_20515,N_20367);
or U21144 (N_21144,N_20562,N_20512);
nand U21145 (N_21145,N_20087,N_20197);
nor U21146 (N_21146,N_20393,N_20054);
nor U21147 (N_21147,N_20327,N_20223);
nand U21148 (N_21148,N_20035,N_20080);
or U21149 (N_21149,N_20453,N_20136);
nor U21150 (N_21150,N_20290,N_20330);
and U21151 (N_21151,N_20100,N_20528);
or U21152 (N_21152,N_20306,N_20261);
or U21153 (N_21153,N_20525,N_20486);
nor U21154 (N_21154,N_20394,N_20416);
and U21155 (N_21155,N_20551,N_20488);
nor U21156 (N_21156,N_20497,N_20281);
or U21157 (N_21157,N_20360,N_20329);
and U21158 (N_21158,N_20312,N_20081);
and U21159 (N_21159,N_20364,N_20620);
or U21160 (N_21160,N_20102,N_20532);
or U21161 (N_21161,N_20590,N_20459);
nand U21162 (N_21162,N_20246,N_20352);
and U21163 (N_21163,N_20548,N_20608);
and U21164 (N_21164,N_20455,N_20102);
and U21165 (N_21165,N_20601,N_20317);
nor U21166 (N_21166,N_20494,N_20318);
or U21167 (N_21167,N_20049,N_20537);
nand U21168 (N_21168,N_20003,N_20176);
nand U21169 (N_21169,N_20391,N_20472);
nor U21170 (N_21170,N_20255,N_20235);
xor U21171 (N_21171,N_20539,N_20180);
or U21172 (N_21172,N_20493,N_20208);
nor U21173 (N_21173,N_20171,N_20266);
nand U21174 (N_21174,N_20286,N_20237);
xnor U21175 (N_21175,N_20039,N_20161);
nor U21176 (N_21176,N_20422,N_20204);
nor U21177 (N_21177,N_20048,N_20160);
or U21178 (N_21178,N_20610,N_20213);
nand U21179 (N_21179,N_20101,N_20349);
and U21180 (N_21180,N_20382,N_20235);
and U21181 (N_21181,N_20398,N_20270);
nor U21182 (N_21182,N_20090,N_20253);
nand U21183 (N_21183,N_20249,N_20003);
nor U21184 (N_21184,N_20565,N_20280);
nor U21185 (N_21185,N_20068,N_20213);
nor U21186 (N_21186,N_20433,N_20442);
nor U21187 (N_21187,N_20541,N_20598);
nand U21188 (N_21188,N_20126,N_20191);
and U21189 (N_21189,N_20516,N_20425);
and U21190 (N_21190,N_20100,N_20037);
nand U21191 (N_21191,N_20137,N_20337);
or U21192 (N_21192,N_20194,N_20101);
nand U21193 (N_21193,N_20306,N_20567);
and U21194 (N_21194,N_20290,N_20220);
nor U21195 (N_21195,N_20459,N_20578);
nand U21196 (N_21196,N_20019,N_20107);
or U21197 (N_21197,N_20590,N_20621);
or U21198 (N_21198,N_20311,N_20278);
xor U21199 (N_21199,N_20066,N_20589);
and U21200 (N_21200,N_20491,N_20231);
and U21201 (N_21201,N_20566,N_20086);
nand U21202 (N_21202,N_20415,N_20157);
nor U21203 (N_21203,N_20137,N_20089);
nor U21204 (N_21204,N_20585,N_20589);
nand U21205 (N_21205,N_20000,N_20320);
or U21206 (N_21206,N_20269,N_20540);
or U21207 (N_21207,N_20162,N_20360);
nand U21208 (N_21208,N_20575,N_20329);
or U21209 (N_21209,N_20343,N_20277);
xor U21210 (N_21210,N_20436,N_20276);
or U21211 (N_21211,N_20256,N_20151);
and U21212 (N_21212,N_20180,N_20020);
or U21213 (N_21213,N_20062,N_20436);
or U21214 (N_21214,N_20514,N_20085);
or U21215 (N_21215,N_20421,N_20443);
and U21216 (N_21216,N_20504,N_20287);
or U21217 (N_21217,N_20440,N_20124);
nand U21218 (N_21218,N_20267,N_20513);
or U21219 (N_21219,N_20456,N_20452);
nor U21220 (N_21220,N_20410,N_20549);
nor U21221 (N_21221,N_20381,N_20116);
or U21222 (N_21222,N_20603,N_20221);
and U21223 (N_21223,N_20376,N_20171);
nand U21224 (N_21224,N_20537,N_20464);
nor U21225 (N_21225,N_20509,N_20350);
nor U21226 (N_21226,N_20026,N_20056);
and U21227 (N_21227,N_20426,N_20340);
nor U21228 (N_21228,N_20411,N_20261);
nor U21229 (N_21229,N_20386,N_20604);
nand U21230 (N_21230,N_20187,N_20518);
nor U21231 (N_21231,N_20517,N_20476);
xor U21232 (N_21232,N_20176,N_20182);
or U21233 (N_21233,N_20383,N_20352);
xnor U21234 (N_21234,N_20166,N_20021);
nor U21235 (N_21235,N_20182,N_20082);
nor U21236 (N_21236,N_20140,N_20287);
or U21237 (N_21237,N_20399,N_20586);
nor U21238 (N_21238,N_20618,N_20396);
nand U21239 (N_21239,N_20525,N_20433);
nor U21240 (N_21240,N_20300,N_20514);
or U21241 (N_21241,N_20074,N_20139);
and U21242 (N_21242,N_20290,N_20592);
nand U21243 (N_21243,N_20087,N_20175);
nand U21244 (N_21244,N_20614,N_20007);
nand U21245 (N_21245,N_20221,N_20192);
or U21246 (N_21246,N_20439,N_20263);
nor U21247 (N_21247,N_20210,N_20608);
or U21248 (N_21248,N_20566,N_20588);
nand U21249 (N_21249,N_20564,N_20038);
nand U21250 (N_21250,N_21036,N_20884);
or U21251 (N_21251,N_20808,N_20740);
xnor U21252 (N_21252,N_20661,N_21104);
nand U21253 (N_21253,N_20665,N_20919);
nor U21254 (N_21254,N_20763,N_20830);
nand U21255 (N_21255,N_21069,N_20681);
and U21256 (N_21256,N_21115,N_20805);
or U21257 (N_21257,N_20709,N_20952);
nor U21258 (N_21258,N_20839,N_20698);
or U21259 (N_21259,N_21113,N_21128);
nand U21260 (N_21260,N_20993,N_21004);
nand U21261 (N_21261,N_20925,N_20883);
nand U21262 (N_21262,N_20869,N_21162);
xor U21263 (N_21263,N_21074,N_20820);
or U21264 (N_21264,N_20652,N_20859);
and U21265 (N_21265,N_21080,N_20813);
or U21266 (N_21266,N_21138,N_20906);
nor U21267 (N_21267,N_20942,N_21220);
nor U21268 (N_21268,N_20890,N_20902);
nor U21269 (N_21269,N_21020,N_21103);
xor U21270 (N_21270,N_20880,N_20670);
nor U21271 (N_21271,N_20856,N_20785);
nand U21272 (N_21272,N_21105,N_21135);
and U21273 (N_21273,N_21034,N_20967);
nand U21274 (N_21274,N_21249,N_20987);
or U21275 (N_21275,N_20625,N_20928);
and U21276 (N_21276,N_20825,N_20804);
and U21277 (N_21277,N_20746,N_21017);
and U21278 (N_21278,N_21029,N_20640);
or U21279 (N_21279,N_20687,N_20806);
nor U21280 (N_21280,N_20650,N_21009);
or U21281 (N_21281,N_21170,N_20947);
or U21282 (N_21282,N_21235,N_20837);
and U21283 (N_21283,N_21018,N_20937);
or U21284 (N_21284,N_20719,N_21091);
xor U21285 (N_21285,N_21125,N_21070);
or U21286 (N_21286,N_20827,N_20848);
nor U21287 (N_21287,N_20770,N_21136);
or U21288 (N_21288,N_21176,N_21085);
nor U21289 (N_21289,N_20767,N_20730);
nand U21290 (N_21290,N_21071,N_20799);
and U21291 (N_21291,N_21043,N_20678);
and U21292 (N_21292,N_21047,N_20940);
nor U21293 (N_21293,N_20817,N_21243);
and U21294 (N_21294,N_21076,N_20929);
or U21295 (N_21295,N_20781,N_20841);
or U21296 (N_21296,N_20680,N_20823);
or U21297 (N_21297,N_21232,N_20751);
nor U21298 (N_21298,N_21062,N_20703);
or U21299 (N_21299,N_20668,N_20992);
or U21300 (N_21300,N_21155,N_21184);
nor U21301 (N_21301,N_21120,N_21233);
nor U21302 (N_21302,N_20803,N_20642);
nor U21303 (N_21303,N_20791,N_21003);
nor U21304 (N_21304,N_20860,N_20842);
nor U21305 (N_21305,N_21141,N_20733);
and U21306 (N_21306,N_21044,N_20855);
xnor U21307 (N_21307,N_21073,N_20801);
or U21308 (N_21308,N_20946,N_20714);
or U21309 (N_21309,N_20754,N_20677);
or U21310 (N_21310,N_20894,N_20838);
nor U21311 (N_21311,N_21021,N_20968);
nand U21312 (N_21312,N_21211,N_20829);
or U21313 (N_21313,N_21189,N_21035);
and U21314 (N_21314,N_20981,N_20818);
nor U21315 (N_21315,N_21122,N_21229);
and U21316 (N_21316,N_20983,N_21090);
nor U21317 (N_21317,N_20927,N_21078);
or U21318 (N_21318,N_20699,N_20912);
xnor U21319 (N_21319,N_20922,N_21234);
nand U21320 (N_21320,N_21041,N_21227);
and U21321 (N_21321,N_20851,N_21192);
xor U21322 (N_21322,N_20995,N_20760);
nand U21323 (N_21323,N_21168,N_21019);
or U21324 (N_21324,N_21228,N_20914);
and U21325 (N_21325,N_20702,N_21033);
nor U21326 (N_21326,N_20713,N_21007);
or U21327 (N_21327,N_20634,N_21181);
and U21328 (N_21328,N_21023,N_20792);
xor U21329 (N_21329,N_21077,N_20950);
or U21330 (N_21330,N_20982,N_20750);
or U21331 (N_21331,N_20951,N_20846);
nand U21332 (N_21332,N_20811,N_20908);
or U21333 (N_21333,N_21154,N_20718);
nand U21334 (N_21334,N_21193,N_20957);
or U21335 (N_21335,N_21101,N_20831);
and U21336 (N_21336,N_21165,N_21147);
and U21337 (N_21337,N_20654,N_20915);
nand U21338 (N_21338,N_20628,N_20828);
and U21339 (N_21339,N_21127,N_20978);
nor U21340 (N_21340,N_21027,N_21191);
or U21341 (N_21341,N_21025,N_20705);
or U21342 (N_21342,N_20786,N_20861);
nor U21343 (N_21343,N_20891,N_21140);
or U21344 (N_21344,N_20695,N_20826);
xor U21345 (N_21345,N_20787,N_20756);
and U21346 (N_21346,N_20753,N_20773);
nor U21347 (N_21347,N_20819,N_20941);
xor U21348 (N_21348,N_21012,N_20676);
or U21349 (N_21349,N_20874,N_21016);
xor U21350 (N_21350,N_20643,N_21067);
or U21351 (N_21351,N_20971,N_21221);
and U21352 (N_21352,N_20758,N_20994);
and U21353 (N_21353,N_21183,N_20669);
or U21354 (N_21354,N_20759,N_20966);
nor U21355 (N_21355,N_20736,N_20970);
or U21356 (N_21356,N_20660,N_20857);
nor U21357 (N_21357,N_20633,N_20782);
nor U21358 (N_21358,N_20933,N_20868);
or U21359 (N_21359,N_20706,N_20683);
or U21360 (N_21360,N_20778,N_21049);
or U21361 (N_21361,N_21039,N_21096);
or U21362 (N_21362,N_21028,N_21093);
and U21363 (N_21363,N_20885,N_20895);
xnor U21364 (N_21364,N_21087,N_20959);
and U21365 (N_21365,N_20744,N_21177);
and U21366 (N_21366,N_20795,N_21010);
or U21367 (N_21367,N_21201,N_20667);
nand U21368 (N_21368,N_21055,N_21095);
and U21369 (N_21369,N_20638,N_21110);
nand U21370 (N_21370,N_21015,N_20732);
and U21371 (N_21371,N_21245,N_21218);
xnor U21372 (N_21372,N_21005,N_20815);
nor U21373 (N_21373,N_20905,N_20696);
or U21374 (N_21374,N_20693,N_21143);
and U21375 (N_21375,N_20737,N_21180);
or U21376 (N_21376,N_21240,N_21088);
or U21377 (N_21377,N_20910,N_21040);
or U21378 (N_21378,N_20986,N_21118);
or U21379 (N_21379,N_21222,N_20641);
or U21380 (N_21380,N_20739,N_20936);
nand U21381 (N_21381,N_20635,N_21013);
nand U21382 (N_21382,N_20742,N_21150);
and U21383 (N_21383,N_20793,N_21030);
nor U21384 (N_21384,N_20892,N_21058);
nor U21385 (N_21385,N_21031,N_20631);
or U21386 (N_21386,N_20802,N_20704);
nor U21387 (N_21387,N_20844,N_21083);
and U21388 (N_21388,N_20916,N_20664);
xnor U21389 (N_21389,N_20889,N_20663);
and U21390 (N_21390,N_20822,N_21172);
and U21391 (N_21391,N_21084,N_21146);
nor U21392 (N_21392,N_21198,N_20666);
or U21393 (N_21393,N_21056,N_20707);
nor U21394 (N_21394,N_21107,N_20903);
nand U21395 (N_21395,N_20685,N_20783);
xor U21396 (N_21396,N_20988,N_21089);
or U21397 (N_21397,N_21171,N_21117);
and U21398 (N_21398,N_20887,N_20961);
and U21399 (N_21399,N_21152,N_20765);
nand U21400 (N_21400,N_20948,N_20990);
and U21401 (N_21401,N_20715,N_20794);
and U21402 (N_21402,N_20757,N_21068);
and U21403 (N_21403,N_21037,N_21203);
or U21404 (N_21404,N_20812,N_21075);
and U21405 (N_21405,N_21001,N_21022);
or U21406 (N_21406,N_21124,N_20735);
xor U21407 (N_21407,N_20866,N_20862);
nor U21408 (N_21408,N_21063,N_21239);
nand U21409 (N_21409,N_20870,N_20741);
nand U21410 (N_21410,N_20907,N_20913);
xor U21411 (N_21411,N_21046,N_20807);
or U21412 (N_21412,N_20694,N_21224);
nor U21413 (N_21413,N_20832,N_20899);
nor U21414 (N_21414,N_21179,N_21237);
and U21415 (N_21415,N_20720,N_21026);
and U21416 (N_21416,N_21116,N_20979);
nor U21417 (N_21417,N_21209,N_20717);
and U21418 (N_21418,N_21108,N_21208);
xnor U21419 (N_21419,N_20748,N_21210);
nand U21420 (N_21420,N_21045,N_20980);
xnor U21421 (N_21421,N_21064,N_21173);
or U21422 (N_21422,N_21188,N_20921);
and U21423 (N_21423,N_20658,N_20973);
nor U21424 (N_21424,N_21175,N_20931);
nor U21425 (N_21425,N_21163,N_20896);
nand U21426 (N_21426,N_21238,N_21212);
or U21427 (N_21427,N_21048,N_20647);
and U21428 (N_21428,N_20840,N_20656);
nand U21429 (N_21429,N_21157,N_20875);
nor U21430 (N_21430,N_20777,N_20873);
nor U21431 (N_21431,N_21161,N_20727);
and U21432 (N_21432,N_21151,N_21052);
nand U21433 (N_21433,N_20675,N_21106);
nor U21434 (N_21434,N_20984,N_21014);
nand U21435 (N_21435,N_20965,N_21137);
and U21436 (N_21436,N_21248,N_20878);
and U21437 (N_21437,N_20996,N_20689);
or U21438 (N_21438,N_20729,N_21159);
or U21439 (N_21439,N_21182,N_20833);
or U21440 (N_21440,N_21119,N_21223);
nand U21441 (N_21441,N_20843,N_21053);
nand U21442 (N_21442,N_20917,N_20836);
nor U21443 (N_21443,N_20886,N_20701);
nand U21444 (N_21444,N_20943,N_21131);
nor U21445 (N_21445,N_20645,N_21167);
and U21446 (N_21446,N_21086,N_20632);
and U21447 (N_21447,N_21242,N_20692);
xor U21448 (N_21448,N_20648,N_20821);
nand U21449 (N_21449,N_21134,N_21126);
or U21450 (N_21450,N_21072,N_20772);
or U21451 (N_21451,N_21079,N_20964);
nand U21452 (N_21452,N_20898,N_20725);
and U21453 (N_21453,N_20649,N_20918);
nor U21454 (N_21454,N_20845,N_21109);
and U21455 (N_21455,N_21097,N_21112);
and U21456 (N_21456,N_21129,N_21098);
and U21457 (N_21457,N_21002,N_20897);
xnor U21458 (N_21458,N_21100,N_21199);
nor U21459 (N_21459,N_20749,N_20769);
or U21460 (N_21460,N_20662,N_20901);
nand U21461 (N_21461,N_20998,N_20834);
xnor U21462 (N_21462,N_20651,N_20771);
nand U21463 (N_21463,N_20997,N_21169);
and U21464 (N_21464,N_20956,N_21065);
nand U21465 (N_21465,N_21213,N_21215);
nor U21466 (N_21466,N_20762,N_21241);
nor U21467 (N_21467,N_20731,N_21059);
xor U21468 (N_21468,N_20776,N_21133);
or U21469 (N_21469,N_21144,N_21236);
or U21470 (N_21470,N_20708,N_20882);
or U21471 (N_21471,N_20955,N_20682);
and U21472 (N_21472,N_20752,N_20939);
or U21473 (N_21473,N_20659,N_20867);
xnor U21474 (N_21474,N_21246,N_20944);
and U21475 (N_21475,N_20977,N_20796);
and U21476 (N_21476,N_20974,N_20888);
nand U21477 (N_21477,N_20626,N_20671);
and U21478 (N_21478,N_21050,N_21123);
xor U21479 (N_21479,N_20644,N_21214);
nor U21480 (N_21480,N_21185,N_20726);
nor U21481 (N_21481,N_20657,N_20688);
or U21482 (N_21482,N_21187,N_21130);
or U21483 (N_21483,N_20945,N_20900);
nand U21484 (N_21484,N_21174,N_20728);
nand U21485 (N_21485,N_21196,N_20653);
or U21486 (N_21486,N_21158,N_20800);
nand U21487 (N_21487,N_20847,N_20932);
and U21488 (N_21488,N_21206,N_20871);
or U21489 (N_21489,N_21038,N_20755);
and U21490 (N_21490,N_21178,N_21102);
nand U21491 (N_21491,N_21226,N_20711);
or U21492 (N_21492,N_21092,N_21166);
nor U21493 (N_21493,N_21032,N_20864);
nor U21494 (N_21494,N_20745,N_20850);
nand U21495 (N_21495,N_21099,N_20674);
nand U21496 (N_21496,N_20716,N_21156);
nor U21497 (N_21497,N_20747,N_20975);
and U21498 (N_21498,N_20969,N_21244);
nor U21499 (N_21499,N_21205,N_20930);
and U21500 (N_21500,N_20784,N_20679);
nand U21501 (N_21501,N_21061,N_20723);
or U21502 (N_21502,N_21024,N_20636);
and U21503 (N_21503,N_20985,N_20646);
or U21504 (N_21504,N_20630,N_21153);
nor U21505 (N_21505,N_21204,N_21011);
or U21506 (N_21506,N_20738,N_21197);
or U21507 (N_21507,N_20963,N_21000);
nand U21508 (N_21508,N_20909,N_20673);
nand U21509 (N_21509,N_20876,N_20768);
nand U21510 (N_21510,N_20637,N_21006);
nor U21511 (N_21511,N_20684,N_21230);
nor U21512 (N_21512,N_20690,N_20893);
or U21513 (N_21513,N_20686,N_21051);
nand U21514 (N_21514,N_20938,N_20989);
and U21515 (N_21515,N_21190,N_21008);
nand U21516 (N_21516,N_20797,N_20790);
or U21517 (N_21517,N_20734,N_21200);
nor U21518 (N_21518,N_20824,N_20999);
or U21519 (N_21519,N_20724,N_21231);
or U21520 (N_21520,N_21082,N_20629);
nand U21521 (N_21521,N_20854,N_20949);
nand U21522 (N_21522,N_21219,N_20672);
or U21523 (N_21523,N_20655,N_20761);
or U21524 (N_21524,N_20863,N_21145);
xor U21525 (N_21525,N_20775,N_20976);
xnor U21526 (N_21526,N_21142,N_20809);
nor U21527 (N_21527,N_21060,N_21114);
xnor U21528 (N_21528,N_20639,N_20991);
or U21529 (N_21529,N_20766,N_20877);
nor U21530 (N_21530,N_20810,N_20697);
and U21531 (N_21531,N_20764,N_20710);
or U21532 (N_21532,N_21160,N_21094);
or U21533 (N_21533,N_20691,N_20872);
nor U21534 (N_21534,N_20849,N_20852);
or U21535 (N_21535,N_20958,N_21217);
nand U21536 (N_21536,N_20814,N_21207);
nor U21537 (N_21537,N_20865,N_20722);
nor U21538 (N_21538,N_21132,N_20835);
or U21539 (N_21539,N_20627,N_21195);
and U21540 (N_21540,N_20798,N_20789);
nor U21541 (N_21541,N_20972,N_21042);
nor U21542 (N_21542,N_20879,N_21054);
and U21543 (N_21543,N_20700,N_20960);
xor U21544 (N_21544,N_20924,N_20858);
xor U21545 (N_21545,N_20926,N_21194);
nand U21546 (N_21546,N_21057,N_21164);
and U21547 (N_21547,N_20953,N_21148);
xnor U21548 (N_21548,N_20904,N_20954);
nor U21549 (N_21549,N_20911,N_20881);
nand U21550 (N_21550,N_21247,N_20774);
and U21551 (N_21551,N_21066,N_21202);
and U21552 (N_21552,N_20779,N_21216);
nor U21553 (N_21553,N_20780,N_20935);
and U21554 (N_21554,N_20923,N_20920);
nor U21555 (N_21555,N_21139,N_21111);
nand U21556 (N_21556,N_21149,N_20816);
nand U21557 (N_21557,N_21121,N_20788);
or U21558 (N_21558,N_20743,N_21186);
and U21559 (N_21559,N_20721,N_20934);
nand U21560 (N_21560,N_21225,N_21081);
xor U21561 (N_21561,N_20853,N_20712);
nand U21562 (N_21562,N_20962,N_20652);
or U21563 (N_21563,N_20682,N_20712);
nand U21564 (N_21564,N_21222,N_21158);
or U21565 (N_21565,N_20632,N_21183);
and U21566 (N_21566,N_20990,N_20664);
nor U21567 (N_21567,N_20815,N_20985);
nor U21568 (N_21568,N_20768,N_21232);
nor U21569 (N_21569,N_21111,N_20855);
nor U21570 (N_21570,N_21221,N_21103);
nor U21571 (N_21571,N_20905,N_21000);
and U21572 (N_21572,N_20701,N_21121);
nand U21573 (N_21573,N_20743,N_20733);
and U21574 (N_21574,N_21043,N_20684);
nand U21575 (N_21575,N_20737,N_20888);
and U21576 (N_21576,N_21127,N_21197);
or U21577 (N_21577,N_21146,N_21243);
or U21578 (N_21578,N_20741,N_20902);
nand U21579 (N_21579,N_20803,N_21110);
or U21580 (N_21580,N_21084,N_20637);
nor U21581 (N_21581,N_20696,N_20694);
and U21582 (N_21582,N_21003,N_20818);
xor U21583 (N_21583,N_20930,N_21222);
and U21584 (N_21584,N_20819,N_20625);
xor U21585 (N_21585,N_20993,N_21196);
or U21586 (N_21586,N_21234,N_20896);
nand U21587 (N_21587,N_20948,N_21211);
xor U21588 (N_21588,N_21043,N_20630);
nand U21589 (N_21589,N_20996,N_21249);
nor U21590 (N_21590,N_20861,N_20925);
xor U21591 (N_21591,N_20786,N_20763);
or U21592 (N_21592,N_20803,N_20626);
and U21593 (N_21593,N_21164,N_20632);
nand U21594 (N_21594,N_20748,N_20831);
and U21595 (N_21595,N_20906,N_21142);
nor U21596 (N_21596,N_20784,N_20668);
xnor U21597 (N_21597,N_20912,N_20844);
and U21598 (N_21598,N_21238,N_21184);
nand U21599 (N_21599,N_20825,N_21227);
nor U21600 (N_21600,N_21157,N_20869);
and U21601 (N_21601,N_20668,N_20857);
nand U21602 (N_21602,N_20663,N_20691);
and U21603 (N_21603,N_20908,N_21013);
nor U21604 (N_21604,N_20716,N_20730);
nand U21605 (N_21605,N_20884,N_21003);
nand U21606 (N_21606,N_21201,N_21023);
xnor U21607 (N_21607,N_20704,N_21058);
and U21608 (N_21608,N_20850,N_20773);
xor U21609 (N_21609,N_20950,N_20876);
nor U21610 (N_21610,N_21203,N_20765);
nor U21611 (N_21611,N_21112,N_20898);
nor U21612 (N_21612,N_20674,N_20953);
or U21613 (N_21613,N_20958,N_21134);
nor U21614 (N_21614,N_20914,N_21205);
nand U21615 (N_21615,N_20691,N_21122);
xor U21616 (N_21616,N_20939,N_21225);
nand U21617 (N_21617,N_21003,N_21185);
xor U21618 (N_21618,N_20790,N_20682);
nor U21619 (N_21619,N_20740,N_20719);
nand U21620 (N_21620,N_21111,N_20726);
nor U21621 (N_21621,N_21185,N_20647);
nor U21622 (N_21622,N_21102,N_20698);
or U21623 (N_21623,N_20678,N_20897);
nor U21624 (N_21624,N_21071,N_20743);
nor U21625 (N_21625,N_21049,N_20842);
and U21626 (N_21626,N_20690,N_21001);
nand U21627 (N_21627,N_20798,N_21188);
or U21628 (N_21628,N_20737,N_20869);
xor U21629 (N_21629,N_20894,N_20768);
and U21630 (N_21630,N_21171,N_20872);
nand U21631 (N_21631,N_20925,N_20705);
and U21632 (N_21632,N_21024,N_20809);
and U21633 (N_21633,N_21224,N_20876);
nor U21634 (N_21634,N_21104,N_21153);
xor U21635 (N_21635,N_21224,N_21153);
or U21636 (N_21636,N_20635,N_20896);
or U21637 (N_21637,N_20905,N_21179);
and U21638 (N_21638,N_20697,N_20964);
nor U21639 (N_21639,N_20967,N_20738);
and U21640 (N_21640,N_20791,N_20983);
and U21641 (N_21641,N_21244,N_21212);
and U21642 (N_21642,N_20885,N_20755);
nand U21643 (N_21643,N_20673,N_21145);
nor U21644 (N_21644,N_21006,N_20932);
nor U21645 (N_21645,N_21118,N_21056);
nand U21646 (N_21646,N_20661,N_20822);
and U21647 (N_21647,N_20855,N_21181);
and U21648 (N_21648,N_20917,N_20851);
or U21649 (N_21649,N_21062,N_20972);
or U21650 (N_21650,N_20708,N_20740);
and U21651 (N_21651,N_21069,N_20640);
or U21652 (N_21652,N_21239,N_20637);
and U21653 (N_21653,N_20642,N_21130);
and U21654 (N_21654,N_20978,N_21176);
nand U21655 (N_21655,N_21167,N_21166);
nor U21656 (N_21656,N_20710,N_21070);
nor U21657 (N_21657,N_20832,N_20902);
and U21658 (N_21658,N_20791,N_21029);
nor U21659 (N_21659,N_21211,N_20754);
nor U21660 (N_21660,N_20978,N_21244);
nand U21661 (N_21661,N_20774,N_20971);
xor U21662 (N_21662,N_20764,N_20940);
nand U21663 (N_21663,N_20984,N_20644);
or U21664 (N_21664,N_20952,N_21048);
nor U21665 (N_21665,N_21131,N_20636);
nand U21666 (N_21666,N_20754,N_20831);
nand U21667 (N_21667,N_20763,N_20777);
and U21668 (N_21668,N_20788,N_20842);
or U21669 (N_21669,N_21033,N_20741);
nor U21670 (N_21670,N_21124,N_21122);
or U21671 (N_21671,N_21141,N_20735);
nor U21672 (N_21672,N_20833,N_21231);
and U21673 (N_21673,N_20944,N_20850);
xnor U21674 (N_21674,N_20732,N_21237);
nand U21675 (N_21675,N_21004,N_20914);
xnor U21676 (N_21676,N_20860,N_21171);
or U21677 (N_21677,N_21125,N_21028);
nand U21678 (N_21678,N_21211,N_20903);
nand U21679 (N_21679,N_20675,N_20877);
nor U21680 (N_21680,N_20636,N_21106);
nand U21681 (N_21681,N_21086,N_20744);
nand U21682 (N_21682,N_20956,N_21011);
or U21683 (N_21683,N_21102,N_20991);
and U21684 (N_21684,N_21187,N_20976);
nand U21685 (N_21685,N_20935,N_20949);
nor U21686 (N_21686,N_21140,N_20967);
and U21687 (N_21687,N_20955,N_20868);
nand U21688 (N_21688,N_21109,N_20982);
xor U21689 (N_21689,N_20733,N_21188);
nand U21690 (N_21690,N_21011,N_21032);
and U21691 (N_21691,N_20665,N_20667);
nand U21692 (N_21692,N_20935,N_20660);
nand U21693 (N_21693,N_20953,N_21220);
or U21694 (N_21694,N_20667,N_21137);
nand U21695 (N_21695,N_21087,N_20708);
and U21696 (N_21696,N_21028,N_21148);
nor U21697 (N_21697,N_20835,N_20954);
or U21698 (N_21698,N_20927,N_21141);
xnor U21699 (N_21699,N_20734,N_20689);
or U21700 (N_21700,N_21198,N_21138);
and U21701 (N_21701,N_20793,N_21152);
and U21702 (N_21702,N_20826,N_21041);
xor U21703 (N_21703,N_21073,N_21038);
nand U21704 (N_21704,N_20972,N_20837);
nand U21705 (N_21705,N_20815,N_20973);
nor U21706 (N_21706,N_20689,N_21105);
nand U21707 (N_21707,N_20910,N_20760);
nand U21708 (N_21708,N_20998,N_21201);
or U21709 (N_21709,N_21204,N_21014);
or U21710 (N_21710,N_21031,N_20862);
nand U21711 (N_21711,N_20812,N_20872);
or U21712 (N_21712,N_20821,N_20642);
or U21713 (N_21713,N_21099,N_21111);
or U21714 (N_21714,N_21032,N_21045);
and U21715 (N_21715,N_21024,N_20775);
xor U21716 (N_21716,N_20719,N_20972);
nor U21717 (N_21717,N_21158,N_20955);
nand U21718 (N_21718,N_20805,N_20881);
or U21719 (N_21719,N_20667,N_20682);
and U21720 (N_21720,N_21051,N_21142);
nand U21721 (N_21721,N_21088,N_20625);
or U21722 (N_21722,N_21017,N_20721);
xor U21723 (N_21723,N_21016,N_21040);
or U21724 (N_21724,N_20727,N_20873);
or U21725 (N_21725,N_20980,N_21155);
and U21726 (N_21726,N_20982,N_20631);
or U21727 (N_21727,N_21027,N_20965);
nor U21728 (N_21728,N_20754,N_21000);
nand U21729 (N_21729,N_21200,N_21174);
nand U21730 (N_21730,N_20690,N_21217);
or U21731 (N_21731,N_21002,N_21037);
nand U21732 (N_21732,N_20779,N_20848);
and U21733 (N_21733,N_21201,N_21196);
nor U21734 (N_21734,N_21138,N_21088);
or U21735 (N_21735,N_21207,N_20914);
or U21736 (N_21736,N_21137,N_20990);
and U21737 (N_21737,N_21047,N_21148);
nor U21738 (N_21738,N_21040,N_20834);
or U21739 (N_21739,N_21224,N_21018);
or U21740 (N_21740,N_21010,N_20804);
nand U21741 (N_21741,N_20923,N_21048);
and U21742 (N_21742,N_20681,N_21187);
nand U21743 (N_21743,N_20719,N_21235);
or U21744 (N_21744,N_20673,N_21045);
and U21745 (N_21745,N_21009,N_20914);
xor U21746 (N_21746,N_21127,N_21146);
nand U21747 (N_21747,N_20922,N_20985);
nand U21748 (N_21748,N_21090,N_21082);
nor U21749 (N_21749,N_20879,N_20868);
or U21750 (N_21750,N_20634,N_20738);
nor U21751 (N_21751,N_20750,N_20990);
nor U21752 (N_21752,N_20802,N_20714);
nand U21753 (N_21753,N_21248,N_20996);
or U21754 (N_21754,N_20960,N_20706);
or U21755 (N_21755,N_20787,N_21166);
xnor U21756 (N_21756,N_21139,N_20861);
and U21757 (N_21757,N_21073,N_20638);
nand U21758 (N_21758,N_21192,N_20743);
xor U21759 (N_21759,N_20789,N_21094);
nor U21760 (N_21760,N_20685,N_21066);
nor U21761 (N_21761,N_20904,N_20956);
xnor U21762 (N_21762,N_21206,N_20763);
nand U21763 (N_21763,N_20741,N_20681);
nor U21764 (N_21764,N_21058,N_20742);
and U21765 (N_21765,N_21096,N_21232);
and U21766 (N_21766,N_20842,N_21141);
nor U21767 (N_21767,N_21016,N_20733);
or U21768 (N_21768,N_20753,N_21155);
and U21769 (N_21769,N_21127,N_20926);
nor U21770 (N_21770,N_20938,N_20781);
or U21771 (N_21771,N_21248,N_20968);
or U21772 (N_21772,N_21231,N_20643);
and U21773 (N_21773,N_21070,N_21085);
nand U21774 (N_21774,N_21100,N_20774);
nand U21775 (N_21775,N_20772,N_20929);
nand U21776 (N_21776,N_20993,N_21211);
nor U21777 (N_21777,N_20997,N_20890);
nor U21778 (N_21778,N_21217,N_20944);
nor U21779 (N_21779,N_20973,N_21120);
or U21780 (N_21780,N_21087,N_20942);
nand U21781 (N_21781,N_21088,N_20868);
or U21782 (N_21782,N_20952,N_21180);
xnor U21783 (N_21783,N_21005,N_20955);
nor U21784 (N_21784,N_21044,N_21079);
nand U21785 (N_21785,N_20889,N_21097);
nand U21786 (N_21786,N_21071,N_21247);
xor U21787 (N_21787,N_20809,N_21130);
xnor U21788 (N_21788,N_20871,N_20975);
nand U21789 (N_21789,N_21044,N_21135);
or U21790 (N_21790,N_21004,N_20653);
nor U21791 (N_21791,N_20641,N_21159);
nand U21792 (N_21792,N_20634,N_20869);
nand U21793 (N_21793,N_20635,N_20695);
nor U21794 (N_21794,N_20725,N_21240);
or U21795 (N_21795,N_21068,N_21023);
nor U21796 (N_21796,N_21105,N_20715);
or U21797 (N_21797,N_20733,N_21060);
nor U21798 (N_21798,N_20812,N_20997);
or U21799 (N_21799,N_20697,N_20756);
xor U21800 (N_21800,N_20905,N_21120);
nand U21801 (N_21801,N_20625,N_20995);
xnor U21802 (N_21802,N_20715,N_21028);
and U21803 (N_21803,N_20786,N_21248);
nor U21804 (N_21804,N_20899,N_21070);
nand U21805 (N_21805,N_20710,N_20847);
and U21806 (N_21806,N_20768,N_21106);
or U21807 (N_21807,N_20626,N_21055);
or U21808 (N_21808,N_21179,N_20711);
and U21809 (N_21809,N_20959,N_20683);
nand U21810 (N_21810,N_20942,N_20709);
nand U21811 (N_21811,N_20841,N_20664);
nor U21812 (N_21812,N_21070,N_21130);
nand U21813 (N_21813,N_20899,N_20699);
or U21814 (N_21814,N_20983,N_20953);
and U21815 (N_21815,N_20998,N_20898);
xnor U21816 (N_21816,N_20677,N_20857);
and U21817 (N_21817,N_20882,N_20860);
nand U21818 (N_21818,N_20665,N_20893);
nor U21819 (N_21819,N_20770,N_21238);
and U21820 (N_21820,N_20741,N_21164);
and U21821 (N_21821,N_21249,N_20917);
xor U21822 (N_21822,N_21148,N_20948);
or U21823 (N_21823,N_21079,N_21137);
and U21824 (N_21824,N_21001,N_20878);
nand U21825 (N_21825,N_20787,N_20845);
nand U21826 (N_21826,N_20969,N_20731);
or U21827 (N_21827,N_20917,N_20814);
and U21828 (N_21828,N_20881,N_20803);
nand U21829 (N_21829,N_21178,N_20998);
or U21830 (N_21830,N_20918,N_20853);
and U21831 (N_21831,N_20797,N_20872);
nor U21832 (N_21832,N_21080,N_20693);
nand U21833 (N_21833,N_20737,N_21137);
nor U21834 (N_21834,N_20886,N_21240);
and U21835 (N_21835,N_20962,N_20641);
xor U21836 (N_21836,N_20740,N_20983);
or U21837 (N_21837,N_21013,N_21111);
nor U21838 (N_21838,N_21024,N_20690);
nor U21839 (N_21839,N_21242,N_20861);
or U21840 (N_21840,N_21230,N_20977);
nor U21841 (N_21841,N_20674,N_20650);
or U21842 (N_21842,N_21162,N_20952);
nor U21843 (N_21843,N_20704,N_20821);
nor U21844 (N_21844,N_20809,N_21005);
or U21845 (N_21845,N_21011,N_20705);
or U21846 (N_21846,N_20700,N_20743);
or U21847 (N_21847,N_21246,N_21154);
nor U21848 (N_21848,N_20989,N_21052);
nand U21849 (N_21849,N_21022,N_21066);
nor U21850 (N_21850,N_20984,N_20829);
nor U21851 (N_21851,N_20791,N_20795);
or U21852 (N_21852,N_21058,N_21106);
nand U21853 (N_21853,N_20636,N_20934);
xor U21854 (N_21854,N_20837,N_21123);
xnor U21855 (N_21855,N_20856,N_20694);
and U21856 (N_21856,N_20647,N_21006);
nor U21857 (N_21857,N_20877,N_21142);
nand U21858 (N_21858,N_20899,N_21201);
and U21859 (N_21859,N_21175,N_21141);
and U21860 (N_21860,N_21079,N_20900);
nand U21861 (N_21861,N_20686,N_21027);
nor U21862 (N_21862,N_20743,N_21076);
or U21863 (N_21863,N_20974,N_20732);
xor U21864 (N_21864,N_20631,N_21166);
nand U21865 (N_21865,N_20798,N_20963);
or U21866 (N_21866,N_20815,N_20643);
xor U21867 (N_21867,N_20732,N_20949);
or U21868 (N_21868,N_21170,N_20710);
and U21869 (N_21869,N_20659,N_20868);
or U21870 (N_21870,N_20922,N_20750);
and U21871 (N_21871,N_20968,N_21011);
and U21872 (N_21872,N_20963,N_20639);
xnor U21873 (N_21873,N_21116,N_21114);
and U21874 (N_21874,N_20980,N_21024);
and U21875 (N_21875,N_21547,N_21355);
and U21876 (N_21876,N_21779,N_21801);
and U21877 (N_21877,N_21759,N_21544);
and U21878 (N_21878,N_21294,N_21467);
nor U21879 (N_21879,N_21439,N_21481);
nor U21880 (N_21880,N_21745,N_21386);
and U21881 (N_21881,N_21468,N_21560);
and U21882 (N_21882,N_21620,N_21354);
nor U21883 (N_21883,N_21316,N_21400);
or U21884 (N_21884,N_21507,N_21292);
nand U21885 (N_21885,N_21325,N_21819);
and U21886 (N_21886,N_21768,N_21852);
or U21887 (N_21887,N_21662,N_21697);
and U21888 (N_21888,N_21426,N_21712);
or U21889 (N_21889,N_21760,N_21539);
xor U21890 (N_21890,N_21252,N_21848);
and U21891 (N_21891,N_21731,N_21659);
nor U21892 (N_21892,N_21617,N_21633);
and U21893 (N_21893,N_21677,N_21710);
nor U21894 (N_21894,N_21775,N_21624);
nor U21895 (N_21895,N_21698,N_21519);
nor U21896 (N_21896,N_21326,N_21791);
nand U21897 (N_21897,N_21749,N_21510);
nand U21898 (N_21898,N_21684,N_21310);
and U21899 (N_21899,N_21838,N_21654);
nand U21900 (N_21900,N_21714,N_21524);
or U21901 (N_21901,N_21689,N_21847);
and U21902 (N_21902,N_21504,N_21328);
nor U21903 (N_21903,N_21757,N_21376);
nor U21904 (N_21904,N_21457,N_21776);
or U21905 (N_21905,N_21827,N_21360);
and U21906 (N_21906,N_21313,N_21844);
and U21907 (N_21907,N_21632,N_21564);
and U21908 (N_21908,N_21756,N_21339);
nor U21909 (N_21909,N_21713,N_21583);
or U21910 (N_21910,N_21482,N_21683);
or U21911 (N_21911,N_21259,N_21650);
or U21912 (N_21912,N_21676,N_21549);
and U21913 (N_21913,N_21611,N_21554);
and U21914 (N_21914,N_21771,N_21347);
and U21915 (N_21915,N_21614,N_21300);
nand U21916 (N_21916,N_21785,N_21484);
or U21917 (N_21917,N_21843,N_21857);
xnor U21918 (N_21918,N_21734,N_21271);
nor U21919 (N_21919,N_21730,N_21494);
xnor U21920 (N_21920,N_21580,N_21559);
nand U21921 (N_21921,N_21767,N_21441);
nand U21922 (N_21922,N_21696,N_21332);
nand U21923 (N_21923,N_21766,N_21378);
nor U21924 (N_21924,N_21609,N_21666);
or U21925 (N_21925,N_21588,N_21597);
or U21926 (N_21926,N_21485,N_21682);
or U21927 (N_21927,N_21809,N_21456);
and U21928 (N_21928,N_21331,N_21258);
nand U21929 (N_21929,N_21299,N_21585);
nor U21930 (N_21930,N_21266,N_21594);
and U21931 (N_21931,N_21639,N_21407);
nor U21932 (N_21932,N_21637,N_21579);
nor U21933 (N_21933,N_21470,N_21543);
nor U21934 (N_21934,N_21513,N_21829);
and U21935 (N_21935,N_21527,N_21402);
and U21936 (N_21936,N_21555,N_21808);
or U21937 (N_21937,N_21694,N_21389);
nor U21938 (N_21938,N_21590,N_21604);
or U21939 (N_21939,N_21334,N_21281);
and U21940 (N_21940,N_21872,N_21670);
nand U21941 (N_21941,N_21781,N_21416);
and U21942 (N_21942,N_21570,N_21511);
or U21943 (N_21943,N_21849,N_21799);
nand U21944 (N_21944,N_21502,N_21871);
nand U21945 (N_21945,N_21828,N_21551);
nor U21946 (N_21946,N_21520,N_21692);
or U21947 (N_21947,N_21303,N_21423);
and U21948 (N_21948,N_21647,N_21412);
xnor U21949 (N_21949,N_21802,N_21257);
and U21950 (N_21950,N_21593,N_21602);
and U21951 (N_21951,N_21516,N_21415);
and U21952 (N_21952,N_21653,N_21874);
and U21953 (N_21953,N_21702,N_21859);
and U21954 (N_21954,N_21794,N_21429);
nand U21955 (N_21955,N_21433,N_21797);
nor U21956 (N_21956,N_21391,N_21866);
xor U21957 (N_21957,N_21368,N_21664);
nand U21958 (N_21958,N_21351,N_21569);
and U21959 (N_21959,N_21419,N_21701);
nand U21960 (N_21960,N_21803,N_21601);
nand U21961 (N_21961,N_21740,N_21600);
nand U21962 (N_21962,N_21619,N_21338);
nand U21963 (N_21963,N_21846,N_21681);
xor U21964 (N_21964,N_21312,N_21317);
nor U21965 (N_21965,N_21306,N_21764);
or U21966 (N_21966,N_21474,N_21725);
and U21967 (N_21967,N_21518,N_21853);
or U21968 (N_21968,N_21792,N_21542);
nor U21969 (N_21969,N_21761,N_21384);
nand U21970 (N_21970,N_21301,N_21422);
nand U21971 (N_21971,N_21536,N_21751);
nand U21972 (N_21972,N_21302,N_21811);
nand U21973 (N_21973,N_21469,N_21733);
or U21974 (N_21974,N_21591,N_21371);
and U21975 (N_21975,N_21497,N_21625);
or U21976 (N_21976,N_21550,N_21421);
nand U21977 (N_21977,N_21443,N_21501);
or U21978 (N_21978,N_21820,N_21599);
nor U21979 (N_21979,N_21277,N_21298);
nor U21980 (N_21980,N_21483,N_21773);
xnor U21981 (N_21981,N_21658,N_21788);
nand U21982 (N_21982,N_21603,N_21635);
or U21983 (N_21983,N_21699,N_21262);
or U21984 (N_21984,N_21736,N_21854);
nor U21985 (N_21985,N_21275,N_21411);
xor U21986 (N_21986,N_21642,N_21521);
xnor U21987 (N_21987,N_21595,N_21668);
or U21988 (N_21988,N_21430,N_21674);
nor U21989 (N_21989,N_21406,N_21405);
nand U21990 (N_21990,N_21466,N_21370);
nor U21991 (N_21991,N_21529,N_21556);
nor U21992 (N_21992,N_21722,N_21623);
and U21993 (N_21993,N_21398,N_21765);
nor U21994 (N_21994,N_21750,N_21748);
xnor U21995 (N_21995,N_21345,N_21574);
nor U21996 (N_21996,N_21655,N_21571);
nor U21997 (N_21997,N_21295,N_21724);
nor U21998 (N_21998,N_21693,N_21489);
nand U21999 (N_21999,N_21287,N_21308);
xor U22000 (N_22000,N_21250,N_21762);
nor U22001 (N_22001,N_21533,N_21818);
nand U22002 (N_22002,N_21311,N_21867);
and U22003 (N_22003,N_21293,N_21414);
nor U22004 (N_22004,N_21831,N_21589);
nand U22005 (N_22005,N_21784,N_21758);
or U22006 (N_22006,N_21538,N_21873);
nor U22007 (N_22007,N_21297,N_21868);
or U22008 (N_22008,N_21735,N_21289);
and U22009 (N_22009,N_21274,N_21256);
or U22010 (N_22010,N_21621,N_21315);
and U22011 (N_22011,N_21522,N_21821);
nand U22012 (N_22012,N_21401,N_21488);
and U22013 (N_22013,N_21573,N_21272);
nor U22014 (N_22014,N_21390,N_21318);
nand U22015 (N_22015,N_21763,N_21596);
or U22016 (N_22016,N_21253,N_21778);
nor U22017 (N_22017,N_21329,N_21631);
or U22018 (N_22018,N_21700,N_21649);
and U22019 (N_22019,N_21616,N_21451);
nand U22020 (N_22020,N_21581,N_21431);
and U22021 (N_22021,N_21263,N_21324);
or U22022 (N_22022,N_21862,N_21517);
and U22023 (N_22023,N_21327,N_21814);
or U22024 (N_22024,N_21687,N_21629);
or U22025 (N_22025,N_21512,N_21335);
and U22026 (N_22026,N_21561,N_21656);
xor U22027 (N_22027,N_21691,N_21265);
or U22028 (N_22028,N_21486,N_21362);
nor U22029 (N_22029,N_21540,N_21806);
and U22030 (N_22030,N_21418,N_21336);
and U22031 (N_22031,N_21323,N_21496);
or U22032 (N_22032,N_21753,N_21665);
or U22033 (N_22033,N_21385,N_21833);
xor U22034 (N_22034,N_21672,N_21462);
or U22035 (N_22035,N_21851,N_21845);
or U22036 (N_22036,N_21744,N_21586);
or U22037 (N_22037,N_21680,N_21690);
nor U22038 (N_22038,N_21251,N_21365);
and U22039 (N_22039,N_21634,N_21491);
nand U22040 (N_22040,N_21839,N_21352);
nand U22041 (N_22041,N_21816,N_21787);
nor U22042 (N_22042,N_21812,N_21798);
xor U22043 (N_22043,N_21563,N_21627);
and U22044 (N_22044,N_21453,N_21707);
xnor U22045 (N_22045,N_21333,N_21545);
nor U22046 (N_22046,N_21841,N_21377);
and U22047 (N_22047,N_21557,N_21738);
nand U22048 (N_22048,N_21458,N_21514);
nor U22049 (N_22049,N_21471,N_21410);
nor U22050 (N_22050,N_21461,N_21372);
and U22051 (N_22051,N_21508,N_21780);
xor U22052 (N_22052,N_21706,N_21737);
or U22053 (N_22053,N_21537,N_21606);
and U22054 (N_22054,N_21836,N_21769);
and U22055 (N_22055,N_21445,N_21671);
or U22056 (N_22056,N_21472,N_21553);
xnor U22057 (N_22057,N_21427,N_21678);
nor U22058 (N_22058,N_21720,N_21492);
or U22059 (N_22059,N_21532,N_21661);
and U22060 (N_22060,N_21503,N_21282);
xnor U22061 (N_22061,N_21552,N_21777);
nand U22062 (N_22062,N_21436,N_21576);
or U22063 (N_22063,N_21379,N_21359);
and U22064 (N_22064,N_21358,N_21709);
nand U22065 (N_22065,N_21715,N_21754);
and U22066 (N_22066,N_21476,N_21346);
and U22067 (N_22067,N_21598,N_21645);
nand U22068 (N_22068,N_21273,N_21770);
nand U22069 (N_22069,N_21528,N_21449);
and U22070 (N_22070,N_21636,N_21782);
or U22071 (N_22071,N_21304,N_21450);
nor U22072 (N_22072,N_21452,N_21361);
and U22073 (N_22073,N_21344,N_21727);
or U22074 (N_22074,N_21864,N_21353);
nand U22075 (N_22075,N_21409,N_21279);
nand U22076 (N_22076,N_21269,N_21437);
nor U22077 (N_22077,N_21646,N_21837);
or U22078 (N_22078,N_21499,N_21319);
and U22079 (N_22079,N_21830,N_21626);
nand U22080 (N_22080,N_21343,N_21870);
nand U22081 (N_22081,N_21267,N_21442);
and U22082 (N_22082,N_21741,N_21506);
or U22083 (N_22083,N_21424,N_21622);
or U22084 (N_22084,N_21800,N_21286);
nand U22085 (N_22085,N_21348,N_21657);
nand U22086 (N_22086,N_21509,N_21505);
and U22087 (N_22087,N_21288,N_21703);
nand U22088 (N_22088,N_21739,N_21708);
and U22089 (N_22089,N_21610,N_21478);
nor U22090 (N_22090,N_21577,N_21607);
and U22091 (N_22091,N_21823,N_21825);
xor U22092 (N_22092,N_21322,N_21465);
and U22093 (N_22093,N_21826,N_21790);
and U22094 (N_22094,N_21732,N_21305);
nor U22095 (N_22095,N_21815,N_21395);
and U22096 (N_22096,N_21705,N_21397);
nor U22097 (N_22097,N_21546,N_21369);
and U22098 (N_22098,N_21455,N_21810);
nor U22099 (N_22099,N_21535,N_21565);
and U22100 (N_22100,N_21480,N_21541);
and U22101 (N_22101,N_21669,N_21381);
or U22102 (N_22102,N_21515,N_21793);
and U22103 (N_22103,N_21796,N_21789);
nand U22104 (N_22104,N_21432,N_21380);
or U22105 (N_22105,N_21349,N_21534);
or U22106 (N_22106,N_21575,N_21280);
xor U22107 (N_22107,N_21578,N_21742);
or U22108 (N_22108,N_21526,N_21382);
nand U22109 (N_22109,N_21718,N_21394);
or U22110 (N_22110,N_21321,N_21464);
xor U22111 (N_22111,N_21834,N_21493);
nand U22112 (N_22112,N_21861,N_21675);
and U22113 (N_22113,N_21630,N_21337);
nand U22114 (N_22114,N_21291,N_21747);
nand U22115 (N_22115,N_21587,N_21392);
and U22116 (N_22116,N_21366,N_21374);
nand U22117 (N_22117,N_21855,N_21572);
and U22118 (N_22118,N_21695,N_21723);
or U22119 (N_22119,N_21448,N_21268);
or U22120 (N_22120,N_21832,N_21804);
nand U22121 (N_22121,N_21805,N_21638);
xor U22122 (N_22122,N_21842,N_21270);
nor U22123 (N_22123,N_21673,N_21605);
and U22124 (N_22124,N_21446,N_21813);
and U22125 (N_22125,N_21644,N_21729);
or U22126 (N_22126,N_21425,N_21567);
nand U22127 (N_22127,N_21858,N_21869);
or U22128 (N_22128,N_21685,N_21479);
nor U22129 (N_22129,N_21717,N_21651);
nand U22130 (N_22130,N_21641,N_21373);
or U22131 (N_22131,N_21660,N_21615);
and U22132 (N_22132,N_21743,N_21417);
nand U22133 (N_22133,N_21640,N_21686);
and U22134 (N_22134,N_21850,N_21613);
nor U22135 (N_22135,N_21428,N_21396);
or U22136 (N_22136,N_21388,N_21679);
and U22137 (N_22137,N_21475,N_21435);
or U22138 (N_22138,N_21403,N_21663);
or U22139 (N_22139,N_21817,N_21824);
nand U22140 (N_22140,N_21568,N_21383);
nor U22141 (N_22141,N_21314,N_21477);
and U22142 (N_22142,N_21283,N_21296);
or U22143 (N_22143,N_21562,N_21835);
nor U22144 (N_22144,N_21774,N_21350);
nand U22145 (N_22145,N_21719,N_21618);
nand U22146 (N_22146,N_21582,N_21454);
nor U22147 (N_22147,N_21726,N_21255);
nor U22148 (N_22148,N_21783,N_21531);
nor U22149 (N_22149,N_21807,N_21490);
xnor U22150 (N_22150,N_21688,N_21364);
xor U22151 (N_22151,N_21608,N_21404);
and U22152 (N_22152,N_21612,N_21363);
nand U22153 (N_22153,N_21460,N_21822);
or U22154 (N_22154,N_21307,N_21420);
or U22155 (N_22155,N_21721,N_21260);
or U22156 (N_22156,N_21434,N_21444);
nand U22157 (N_22157,N_21309,N_21860);
nand U22158 (N_22158,N_21447,N_21856);
or U22159 (N_22159,N_21367,N_21558);
and U22160 (N_22160,N_21495,N_21340);
and U22161 (N_22161,N_21290,N_21704);
and U22162 (N_22162,N_21628,N_21648);
or U22163 (N_22163,N_21716,N_21525);
and U22164 (N_22164,N_21752,N_21356);
nor U22165 (N_22165,N_21463,N_21393);
nand U22166 (N_22166,N_21487,N_21840);
and U22167 (N_22167,N_21375,N_21440);
or U22168 (N_22168,N_21530,N_21566);
or U22169 (N_22169,N_21320,N_21459);
nand U22170 (N_22170,N_21284,N_21276);
nor U22171 (N_22171,N_21667,N_21772);
nand U22172 (N_22172,N_21500,N_21264);
and U22173 (N_22173,N_21342,N_21399);
and U22174 (N_22174,N_21357,N_21592);
or U22175 (N_22175,N_21755,N_21498);
nor U22176 (N_22176,N_21795,N_21643);
or U22177 (N_22177,N_21254,N_21438);
nor U22178 (N_22178,N_21652,N_21330);
or U22179 (N_22179,N_21473,N_21408);
xor U22180 (N_22180,N_21285,N_21746);
nand U22181 (N_22181,N_21413,N_21786);
xnor U22182 (N_22182,N_21278,N_21728);
or U22183 (N_22183,N_21584,N_21387);
nor U22184 (N_22184,N_21865,N_21261);
nand U22185 (N_22185,N_21548,N_21711);
or U22186 (N_22186,N_21341,N_21863);
xor U22187 (N_22187,N_21523,N_21850);
and U22188 (N_22188,N_21496,N_21751);
nand U22189 (N_22189,N_21780,N_21676);
and U22190 (N_22190,N_21693,N_21855);
or U22191 (N_22191,N_21623,N_21548);
nand U22192 (N_22192,N_21763,N_21672);
and U22193 (N_22193,N_21578,N_21530);
or U22194 (N_22194,N_21437,N_21611);
or U22195 (N_22195,N_21785,N_21586);
and U22196 (N_22196,N_21323,N_21801);
and U22197 (N_22197,N_21710,N_21341);
xor U22198 (N_22198,N_21592,N_21683);
nand U22199 (N_22199,N_21440,N_21422);
nand U22200 (N_22200,N_21516,N_21514);
nand U22201 (N_22201,N_21566,N_21531);
nor U22202 (N_22202,N_21298,N_21575);
or U22203 (N_22203,N_21600,N_21315);
nor U22204 (N_22204,N_21606,N_21593);
nand U22205 (N_22205,N_21870,N_21632);
and U22206 (N_22206,N_21866,N_21363);
nor U22207 (N_22207,N_21514,N_21357);
nand U22208 (N_22208,N_21317,N_21816);
nand U22209 (N_22209,N_21429,N_21531);
and U22210 (N_22210,N_21710,N_21812);
nor U22211 (N_22211,N_21637,N_21531);
nor U22212 (N_22212,N_21491,N_21547);
and U22213 (N_22213,N_21425,N_21733);
xor U22214 (N_22214,N_21537,N_21447);
or U22215 (N_22215,N_21696,N_21869);
or U22216 (N_22216,N_21396,N_21676);
nand U22217 (N_22217,N_21580,N_21448);
and U22218 (N_22218,N_21749,N_21835);
and U22219 (N_22219,N_21255,N_21301);
xnor U22220 (N_22220,N_21486,N_21422);
nor U22221 (N_22221,N_21430,N_21561);
nand U22222 (N_22222,N_21665,N_21775);
or U22223 (N_22223,N_21264,N_21836);
nor U22224 (N_22224,N_21666,N_21298);
nor U22225 (N_22225,N_21456,N_21682);
and U22226 (N_22226,N_21262,N_21747);
nor U22227 (N_22227,N_21521,N_21562);
or U22228 (N_22228,N_21423,N_21475);
and U22229 (N_22229,N_21784,N_21851);
nor U22230 (N_22230,N_21823,N_21301);
xor U22231 (N_22231,N_21547,N_21477);
nor U22232 (N_22232,N_21857,N_21417);
or U22233 (N_22233,N_21298,N_21561);
and U22234 (N_22234,N_21398,N_21817);
and U22235 (N_22235,N_21746,N_21485);
nor U22236 (N_22236,N_21757,N_21445);
or U22237 (N_22237,N_21359,N_21632);
or U22238 (N_22238,N_21460,N_21397);
or U22239 (N_22239,N_21488,N_21341);
nand U22240 (N_22240,N_21466,N_21759);
xor U22241 (N_22241,N_21583,N_21560);
nor U22242 (N_22242,N_21687,N_21786);
or U22243 (N_22243,N_21818,N_21869);
nand U22244 (N_22244,N_21470,N_21334);
nand U22245 (N_22245,N_21836,N_21713);
and U22246 (N_22246,N_21635,N_21467);
nor U22247 (N_22247,N_21847,N_21574);
and U22248 (N_22248,N_21564,N_21857);
or U22249 (N_22249,N_21660,N_21856);
and U22250 (N_22250,N_21324,N_21649);
or U22251 (N_22251,N_21405,N_21282);
xnor U22252 (N_22252,N_21846,N_21497);
xor U22253 (N_22253,N_21735,N_21676);
or U22254 (N_22254,N_21623,N_21730);
and U22255 (N_22255,N_21496,N_21680);
nor U22256 (N_22256,N_21571,N_21681);
or U22257 (N_22257,N_21673,N_21458);
xnor U22258 (N_22258,N_21664,N_21579);
nor U22259 (N_22259,N_21822,N_21288);
and U22260 (N_22260,N_21711,N_21874);
and U22261 (N_22261,N_21394,N_21551);
and U22262 (N_22262,N_21774,N_21728);
nor U22263 (N_22263,N_21441,N_21361);
and U22264 (N_22264,N_21705,N_21839);
xor U22265 (N_22265,N_21668,N_21567);
or U22266 (N_22266,N_21424,N_21310);
and U22267 (N_22267,N_21509,N_21678);
nor U22268 (N_22268,N_21635,N_21717);
or U22269 (N_22269,N_21758,N_21339);
or U22270 (N_22270,N_21673,N_21710);
or U22271 (N_22271,N_21569,N_21299);
nor U22272 (N_22272,N_21260,N_21849);
or U22273 (N_22273,N_21497,N_21392);
or U22274 (N_22274,N_21369,N_21725);
or U22275 (N_22275,N_21266,N_21846);
or U22276 (N_22276,N_21291,N_21662);
xor U22277 (N_22277,N_21719,N_21737);
or U22278 (N_22278,N_21660,N_21337);
xnor U22279 (N_22279,N_21602,N_21265);
and U22280 (N_22280,N_21866,N_21840);
nand U22281 (N_22281,N_21456,N_21808);
nor U22282 (N_22282,N_21534,N_21815);
or U22283 (N_22283,N_21447,N_21376);
and U22284 (N_22284,N_21310,N_21290);
xnor U22285 (N_22285,N_21740,N_21361);
or U22286 (N_22286,N_21338,N_21762);
or U22287 (N_22287,N_21459,N_21254);
and U22288 (N_22288,N_21372,N_21666);
nand U22289 (N_22289,N_21296,N_21403);
or U22290 (N_22290,N_21779,N_21376);
xnor U22291 (N_22291,N_21407,N_21759);
or U22292 (N_22292,N_21797,N_21585);
and U22293 (N_22293,N_21802,N_21345);
or U22294 (N_22294,N_21380,N_21440);
nor U22295 (N_22295,N_21616,N_21744);
xor U22296 (N_22296,N_21707,N_21551);
and U22297 (N_22297,N_21397,N_21699);
nand U22298 (N_22298,N_21277,N_21802);
nor U22299 (N_22299,N_21873,N_21574);
and U22300 (N_22300,N_21276,N_21432);
nand U22301 (N_22301,N_21517,N_21271);
or U22302 (N_22302,N_21629,N_21669);
and U22303 (N_22303,N_21811,N_21327);
xor U22304 (N_22304,N_21421,N_21292);
nor U22305 (N_22305,N_21361,N_21590);
or U22306 (N_22306,N_21326,N_21463);
nand U22307 (N_22307,N_21366,N_21566);
and U22308 (N_22308,N_21762,N_21267);
nand U22309 (N_22309,N_21697,N_21309);
and U22310 (N_22310,N_21429,N_21704);
and U22311 (N_22311,N_21285,N_21699);
and U22312 (N_22312,N_21839,N_21728);
or U22313 (N_22313,N_21290,N_21487);
nand U22314 (N_22314,N_21358,N_21408);
nor U22315 (N_22315,N_21471,N_21312);
nor U22316 (N_22316,N_21779,N_21822);
xnor U22317 (N_22317,N_21355,N_21626);
nor U22318 (N_22318,N_21463,N_21464);
nor U22319 (N_22319,N_21315,N_21400);
nor U22320 (N_22320,N_21404,N_21263);
nand U22321 (N_22321,N_21335,N_21539);
or U22322 (N_22322,N_21521,N_21667);
nor U22323 (N_22323,N_21470,N_21494);
and U22324 (N_22324,N_21720,N_21461);
xnor U22325 (N_22325,N_21370,N_21394);
or U22326 (N_22326,N_21762,N_21802);
nand U22327 (N_22327,N_21266,N_21263);
or U22328 (N_22328,N_21637,N_21862);
and U22329 (N_22329,N_21588,N_21395);
nand U22330 (N_22330,N_21743,N_21873);
nand U22331 (N_22331,N_21798,N_21508);
nor U22332 (N_22332,N_21594,N_21325);
nand U22333 (N_22333,N_21342,N_21483);
nand U22334 (N_22334,N_21338,N_21818);
nor U22335 (N_22335,N_21319,N_21305);
nor U22336 (N_22336,N_21735,N_21772);
nand U22337 (N_22337,N_21785,N_21417);
and U22338 (N_22338,N_21861,N_21594);
nand U22339 (N_22339,N_21686,N_21598);
nand U22340 (N_22340,N_21656,N_21568);
xnor U22341 (N_22341,N_21532,N_21775);
or U22342 (N_22342,N_21366,N_21537);
nor U22343 (N_22343,N_21514,N_21414);
or U22344 (N_22344,N_21330,N_21820);
nor U22345 (N_22345,N_21426,N_21579);
or U22346 (N_22346,N_21272,N_21585);
nor U22347 (N_22347,N_21701,N_21696);
or U22348 (N_22348,N_21467,N_21619);
or U22349 (N_22349,N_21323,N_21489);
and U22350 (N_22350,N_21447,N_21520);
xor U22351 (N_22351,N_21734,N_21640);
nand U22352 (N_22352,N_21527,N_21411);
or U22353 (N_22353,N_21477,N_21690);
nand U22354 (N_22354,N_21739,N_21606);
xor U22355 (N_22355,N_21326,N_21583);
nor U22356 (N_22356,N_21619,N_21330);
or U22357 (N_22357,N_21489,N_21763);
or U22358 (N_22358,N_21505,N_21822);
xor U22359 (N_22359,N_21342,N_21750);
xor U22360 (N_22360,N_21333,N_21654);
and U22361 (N_22361,N_21469,N_21717);
or U22362 (N_22362,N_21319,N_21520);
or U22363 (N_22363,N_21666,N_21335);
nand U22364 (N_22364,N_21389,N_21757);
or U22365 (N_22365,N_21440,N_21439);
or U22366 (N_22366,N_21612,N_21391);
nor U22367 (N_22367,N_21524,N_21676);
xor U22368 (N_22368,N_21794,N_21279);
or U22369 (N_22369,N_21492,N_21726);
xnor U22370 (N_22370,N_21435,N_21580);
and U22371 (N_22371,N_21468,N_21401);
and U22372 (N_22372,N_21866,N_21539);
or U22373 (N_22373,N_21484,N_21722);
nand U22374 (N_22374,N_21684,N_21603);
or U22375 (N_22375,N_21427,N_21523);
or U22376 (N_22376,N_21832,N_21723);
and U22377 (N_22377,N_21267,N_21315);
and U22378 (N_22378,N_21735,N_21724);
and U22379 (N_22379,N_21593,N_21575);
and U22380 (N_22380,N_21344,N_21722);
nor U22381 (N_22381,N_21459,N_21281);
nor U22382 (N_22382,N_21731,N_21546);
or U22383 (N_22383,N_21326,N_21307);
nand U22384 (N_22384,N_21728,N_21363);
nor U22385 (N_22385,N_21711,N_21573);
nor U22386 (N_22386,N_21623,N_21682);
nand U22387 (N_22387,N_21379,N_21444);
nor U22388 (N_22388,N_21532,N_21726);
or U22389 (N_22389,N_21669,N_21763);
or U22390 (N_22390,N_21715,N_21619);
xor U22391 (N_22391,N_21754,N_21610);
nand U22392 (N_22392,N_21297,N_21695);
nand U22393 (N_22393,N_21297,N_21590);
or U22394 (N_22394,N_21799,N_21254);
nor U22395 (N_22395,N_21679,N_21576);
xor U22396 (N_22396,N_21645,N_21458);
and U22397 (N_22397,N_21632,N_21636);
or U22398 (N_22398,N_21538,N_21638);
and U22399 (N_22399,N_21611,N_21389);
nor U22400 (N_22400,N_21380,N_21561);
nand U22401 (N_22401,N_21618,N_21522);
nor U22402 (N_22402,N_21480,N_21684);
nand U22403 (N_22403,N_21741,N_21334);
or U22404 (N_22404,N_21283,N_21622);
and U22405 (N_22405,N_21289,N_21265);
nor U22406 (N_22406,N_21475,N_21804);
nand U22407 (N_22407,N_21521,N_21761);
xnor U22408 (N_22408,N_21739,N_21348);
and U22409 (N_22409,N_21258,N_21839);
nand U22410 (N_22410,N_21457,N_21835);
nand U22411 (N_22411,N_21738,N_21599);
xor U22412 (N_22412,N_21374,N_21269);
nor U22413 (N_22413,N_21867,N_21518);
xnor U22414 (N_22414,N_21861,N_21390);
or U22415 (N_22415,N_21617,N_21672);
or U22416 (N_22416,N_21758,N_21627);
xnor U22417 (N_22417,N_21357,N_21530);
or U22418 (N_22418,N_21827,N_21528);
nor U22419 (N_22419,N_21488,N_21742);
and U22420 (N_22420,N_21629,N_21327);
nor U22421 (N_22421,N_21523,N_21380);
or U22422 (N_22422,N_21716,N_21535);
xor U22423 (N_22423,N_21709,N_21596);
and U22424 (N_22424,N_21867,N_21570);
nand U22425 (N_22425,N_21790,N_21772);
nor U22426 (N_22426,N_21721,N_21350);
or U22427 (N_22427,N_21355,N_21280);
or U22428 (N_22428,N_21309,N_21463);
nand U22429 (N_22429,N_21416,N_21405);
or U22430 (N_22430,N_21443,N_21326);
and U22431 (N_22431,N_21578,N_21874);
or U22432 (N_22432,N_21542,N_21253);
or U22433 (N_22433,N_21638,N_21271);
and U22434 (N_22434,N_21340,N_21540);
or U22435 (N_22435,N_21475,N_21690);
nand U22436 (N_22436,N_21657,N_21760);
nand U22437 (N_22437,N_21767,N_21693);
nor U22438 (N_22438,N_21327,N_21314);
nand U22439 (N_22439,N_21470,N_21562);
nand U22440 (N_22440,N_21622,N_21826);
and U22441 (N_22441,N_21313,N_21333);
nor U22442 (N_22442,N_21534,N_21500);
xor U22443 (N_22443,N_21331,N_21477);
or U22444 (N_22444,N_21348,N_21554);
nor U22445 (N_22445,N_21856,N_21272);
nor U22446 (N_22446,N_21748,N_21767);
and U22447 (N_22447,N_21269,N_21653);
and U22448 (N_22448,N_21690,N_21705);
nor U22449 (N_22449,N_21811,N_21297);
nor U22450 (N_22450,N_21846,N_21661);
and U22451 (N_22451,N_21618,N_21823);
nor U22452 (N_22452,N_21416,N_21815);
or U22453 (N_22453,N_21798,N_21607);
nand U22454 (N_22454,N_21313,N_21439);
and U22455 (N_22455,N_21382,N_21708);
xnor U22456 (N_22456,N_21692,N_21488);
nor U22457 (N_22457,N_21367,N_21510);
nor U22458 (N_22458,N_21589,N_21380);
nor U22459 (N_22459,N_21569,N_21474);
and U22460 (N_22460,N_21690,N_21653);
xnor U22461 (N_22461,N_21659,N_21664);
nor U22462 (N_22462,N_21549,N_21329);
nor U22463 (N_22463,N_21775,N_21377);
nor U22464 (N_22464,N_21626,N_21442);
xor U22465 (N_22465,N_21435,N_21634);
nor U22466 (N_22466,N_21542,N_21612);
nor U22467 (N_22467,N_21799,N_21532);
nor U22468 (N_22468,N_21620,N_21470);
or U22469 (N_22469,N_21698,N_21567);
or U22470 (N_22470,N_21317,N_21725);
nor U22471 (N_22471,N_21656,N_21254);
nand U22472 (N_22472,N_21674,N_21730);
xnor U22473 (N_22473,N_21299,N_21289);
xnor U22474 (N_22474,N_21250,N_21359);
or U22475 (N_22475,N_21269,N_21632);
nand U22476 (N_22476,N_21811,N_21873);
nor U22477 (N_22477,N_21806,N_21533);
xor U22478 (N_22478,N_21577,N_21772);
and U22479 (N_22479,N_21415,N_21638);
or U22480 (N_22480,N_21294,N_21660);
and U22481 (N_22481,N_21306,N_21316);
and U22482 (N_22482,N_21667,N_21751);
nand U22483 (N_22483,N_21749,N_21515);
and U22484 (N_22484,N_21457,N_21356);
nand U22485 (N_22485,N_21498,N_21840);
and U22486 (N_22486,N_21600,N_21414);
nand U22487 (N_22487,N_21558,N_21543);
nand U22488 (N_22488,N_21854,N_21749);
nor U22489 (N_22489,N_21449,N_21715);
nor U22490 (N_22490,N_21479,N_21823);
nand U22491 (N_22491,N_21271,N_21822);
nor U22492 (N_22492,N_21862,N_21520);
and U22493 (N_22493,N_21383,N_21363);
or U22494 (N_22494,N_21641,N_21677);
nor U22495 (N_22495,N_21833,N_21697);
xor U22496 (N_22496,N_21601,N_21411);
nand U22497 (N_22497,N_21660,N_21463);
or U22498 (N_22498,N_21650,N_21794);
xnor U22499 (N_22499,N_21866,N_21301);
and U22500 (N_22500,N_22121,N_22087);
nor U22501 (N_22501,N_22219,N_22295);
or U22502 (N_22502,N_22246,N_22028);
nand U22503 (N_22503,N_22381,N_22438);
xor U22504 (N_22504,N_22106,N_22138);
xor U22505 (N_22505,N_22092,N_22254);
nand U22506 (N_22506,N_22492,N_21883);
and U22507 (N_22507,N_21973,N_21927);
or U22508 (N_22508,N_21953,N_22238);
or U22509 (N_22509,N_22173,N_22032);
or U22510 (N_22510,N_21961,N_22355);
nand U22511 (N_22511,N_22080,N_22304);
nand U22512 (N_22512,N_21955,N_22296);
nor U22513 (N_22513,N_22021,N_22207);
nor U22514 (N_22514,N_22373,N_22039);
and U22515 (N_22515,N_22199,N_22435);
nand U22516 (N_22516,N_22306,N_21985);
and U22517 (N_22517,N_22198,N_22111);
and U22518 (N_22518,N_22382,N_22083);
and U22519 (N_22519,N_22142,N_22062);
nor U22520 (N_22520,N_21937,N_22241);
or U22521 (N_22521,N_22264,N_22461);
and U22522 (N_22522,N_22042,N_22345);
nor U22523 (N_22523,N_22495,N_21980);
or U22524 (N_22524,N_22401,N_22444);
nor U22525 (N_22525,N_22457,N_22251);
xor U22526 (N_22526,N_22068,N_22147);
and U22527 (N_22527,N_22011,N_22233);
nor U22528 (N_22528,N_22108,N_21960);
nor U22529 (N_22529,N_21981,N_22416);
nor U22530 (N_22530,N_22239,N_22353);
and U22531 (N_22531,N_21903,N_22483);
and U22532 (N_22532,N_22336,N_22144);
nor U22533 (N_22533,N_21877,N_22112);
or U22534 (N_22534,N_22486,N_22195);
nor U22535 (N_22535,N_22051,N_22115);
and U22536 (N_22536,N_21935,N_22452);
nor U22537 (N_22537,N_22300,N_22344);
nor U22538 (N_22538,N_22424,N_22427);
nand U22539 (N_22539,N_22110,N_22282);
nand U22540 (N_22540,N_21963,N_21896);
nand U22541 (N_22541,N_22456,N_22003);
nand U22542 (N_22542,N_22440,N_21881);
nand U22543 (N_22543,N_22078,N_22314);
nor U22544 (N_22544,N_21987,N_21879);
and U22545 (N_22545,N_22118,N_22046);
and U22546 (N_22546,N_21932,N_22349);
and U22547 (N_22547,N_22363,N_21956);
and U22548 (N_22548,N_22129,N_22482);
xor U22549 (N_22549,N_22160,N_22458);
and U22550 (N_22550,N_22367,N_21912);
or U22551 (N_22551,N_22259,N_22136);
or U22552 (N_22552,N_22037,N_22171);
and U22553 (N_22553,N_22311,N_22220);
nor U22554 (N_22554,N_22043,N_22002);
nor U22555 (N_22555,N_22408,N_22348);
xor U22556 (N_22556,N_22356,N_22499);
xnor U22557 (N_22557,N_22268,N_22075);
or U22558 (N_22558,N_22470,N_22232);
and U22559 (N_22559,N_22298,N_22474);
nand U22560 (N_22560,N_21999,N_22377);
or U22561 (N_22561,N_22030,N_22286);
or U22562 (N_22562,N_21967,N_22380);
nand U22563 (N_22563,N_22411,N_22479);
nand U22564 (N_22564,N_22359,N_22386);
and U22565 (N_22565,N_22364,N_22274);
and U22566 (N_22566,N_22006,N_21929);
and U22567 (N_22567,N_22124,N_22493);
nand U22568 (N_22568,N_22013,N_21957);
or U22569 (N_22569,N_21965,N_22064);
nand U22570 (N_22570,N_22392,N_22001);
nor U22571 (N_22571,N_22188,N_22409);
nand U22572 (N_22572,N_22229,N_22098);
and U22573 (N_22573,N_21942,N_22150);
or U22574 (N_22574,N_22225,N_22186);
and U22575 (N_22575,N_21888,N_22465);
nand U22576 (N_22576,N_22217,N_21890);
or U22577 (N_22577,N_22293,N_22489);
or U22578 (N_22578,N_21944,N_22404);
and U22579 (N_22579,N_22308,N_22091);
and U22580 (N_22580,N_21934,N_21892);
nor U22581 (N_22581,N_22278,N_22156);
nand U22582 (N_22582,N_21940,N_21966);
or U22583 (N_22583,N_22323,N_22339);
or U22584 (N_22584,N_22163,N_22387);
nor U22585 (N_22585,N_22463,N_22430);
nand U22586 (N_22586,N_22146,N_22284);
nor U22587 (N_22587,N_22369,N_22354);
nor U22588 (N_22588,N_22275,N_22454);
xnor U22589 (N_22589,N_22109,N_22012);
and U22590 (N_22590,N_22069,N_22405);
or U22591 (N_22591,N_21978,N_21899);
nor U22592 (N_22592,N_22168,N_22289);
nor U22593 (N_22593,N_22135,N_22291);
and U22594 (N_22594,N_22185,N_22089);
nand U22595 (N_22595,N_22335,N_22056);
nand U22596 (N_22596,N_21908,N_22179);
and U22597 (N_22597,N_21971,N_22297);
nor U22598 (N_22598,N_21996,N_22439);
nor U22599 (N_22599,N_22227,N_22172);
or U22600 (N_22600,N_22020,N_22352);
or U22601 (N_22601,N_21982,N_21950);
or U22602 (N_22602,N_22016,N_22317);
and U22603 (N_22603,N_22182,N_22368);
nor U22604 (N_22604,N_22266,N_22009);
or U22605 (N_22605,N_22299,N_22476);
nor U22606 (N_22606,N_22212,N_22017);
nand U22607 (N_22607,N_22361,N_22200);
or U22608 (N_22608,N_22162,N_22272);
and U22609 (N_22609,N_22191,N_22468);
nor U22610 (N_22610,N_22120,N_22370);
xnor U22611 (N_22611,N_22258,N_22022);
or U22612 (N_22612,N_22005,N_22175);
and U22613 (N_22613,N_22079,N_22215);
nor U22614 (N_22614,N_22366,N_22450);
nor U22615 (N_22615,N_22052,N_22464);
nand U22616 (N_22616,N_22252,N_22059);
and U22617 (N_22617,N_21951,N_22221);
and U22618 (N_22618,N_22332,N_22139);
xnor U22619 (N_22619,N_22161,N_22050);
xor U22620 (N_22620,N_22477,N_21914);
or U22621 (N_22621,N_22211,N_22174);
or U22622 (N_22622,N_22248,N_22036);
and U22623 (N_22623,N_22395,N_22434);
or U22624 (N_22624,N_22183,N_22360);
nand U22625 (N_22625,N_22234,N_22034);
and U22626 (N_22626,N_22031,N_22343);
or U22627 (N_22627,N_22460,N_22329);
nand U22628 (N_22628,N_22316,N_21891);
nand U22629 (N_22629,N_22393,N_22331);
and U22630 (N_22630,N_22255,N_21976);
nor U22631 (N_22631,N_22378,N_22473);
nor U22632 (N_22632,N_22431,N_22384);
or U22633 (N_22633,N_22128,N_22184);
and U22634 (N_22634,N_22469,N_22014);
nand U22635 (N_22635,N_22351,N_21958);
nand U22636 (N_22636,N_22204,N_21994);
and U22637 (N_22637,N_22257,N_22421);
or U22638 (N_22638,N_21933,N_21954);
nand U22639 (N_22639,N_22117,N_22243);
or U22640 (N_22640,N_22250,N_22410);
and U22641 (N_22641,N_22342,N_21986);
or U22642 (N_22642,N_22058,N_22165);
nor U22643 (N_22643,N_21979,N_22029);
and U22644 (N_22644,N_21972,N_22177);
and U22645 (N_22645,N_22226,N_22152);
and U22646 (N_22646,N_22350,N_21931);
nand U22647 (N_22647,N_22472,N_22223);
nand U22648 (N_22648,N_22023,N_22310);
nor U22649 (N_22649,N_22480,N_22490);
nand U22650 (N_22650,N_22292,N_22097);
nand U22651 (N_22651,N_22374,N_22385);
xnor U22652 (N_22652,N_22337,N_22280);
xor U22653 (N_22653,N_22467,N_22396);
nor U22654 (N_22654,N_21930,N_22498);
or U22655 (N_22655,N_22145,N_22245);
nand U22656 (N_22656,N_22389,N_22497);
and U22657 (N_22657,N_22273,N_22305);
and U22658 (N_22658,N_22203,N_21897);
nor U22659 (N_22659,N_22481,N_22445);
xnor U22660 (N_22660,N_22433,N_22063);
and U22661 (N_22661,N_21923,N_22442);
nor U22662 (N_22662,N_22169,N_22281);
and U22663 (N_22663,N_22277,N_21876);
and U22664 (N_22664,N_21924,N_21880);
xnor U22665 (N_22665,N_22082,N_22099);
or U22666 (N_22666,N_22073,N_22010);
nor U22667 (N_22667,N_22055,N_22302);
nand U22668 (N_22668,N_22287,N_22049);
or U22669 (N_22669,N_22466,N_22340);
nor U22670 (N_22670,N_22253,N_22303);
and U22671 (N_22671,N_22209,N_22371);
or U22672 (N_22672,N_21900,N_22334);
nor U22673 (N_22673,N_21909,N_21921);
nor U22674 (N_22674,N_22321,N_22276);
or U22675 (N_22675,N_22153,N_22155);
nand U22676 (N_22676,N_22201,N_22487);
nor U22677 (N_22677,N_21990,N_21918);
nand U22678 (N_22678,N_22488,N_22154);
and U22679 (N_22679,N_22040,N_22485);
and U22680 (N_22680,N_21911,N_22419);
nand U22681 (N_22681,N_22213,N_22265);
nor U22682 (N_22682,N_22143,N_22053);
and U22683 (N_22683,N_22475,N_22026);
nand U22684 (N_22684,N_21995,N_22491);
and U22685 (N_22685,N_21910,N_21904);
nor U22686 (N_22686,N_22065,N_22159);
nand U22687 (N_22687,N_22164,N_21917);
and U22688 (N_22688,N_22423,N_22412);
nand U22689 (N_22689,N_22170,N_21969);
nor U22690 (N_22690,N_21962,N_22365);
nor U22691 (N_22691,N_22496,N_22119);
nor U22692 (N_22692,N_22134,N_22402);
and U22693 (N_22693,N_22437,N_22315);
nor U22694 (N_22694,N_22151,N_21989);
nand U22695 (N_22695,N_21945,N_22070);
or U22696 (N_22696,N_22425,N_22319);
nand U22697 (N_22697,N_22224,N_21997);
or U22698 (N_22698,N_22066,N_22441);
nand U22699 (N_22699,N_22000,N_22478);
xnor U22700 (N_22700,N_22418,N_22123);
or U22701 (N_22701,N_21901,N_22007);
and U22702 (N_22702,N_21913,N_22432);
nand U22703 (N_22703,N_22459,N_22372);
xnor U22704 (N_22704,N_22107,N_22443);
xor U22705 (N_22705,N_22471,N_22375);
or U22706 (N_22706,N_22222,N_21988);
nor U22707 (N_22707,N_22379,N_22048);
and U22708 (N_22708,N_22328,N_22018);
and U22709 (N_22709,N_22294,N_21949);
nor U22710 (N_22710,N_22362,N_22131);
nand U22711 (N_22711,N_22247,N_22196);
nor U22712 (N_22712,N_21984,N_22019);
and U22713 (N_22713,N_22325,N_22004);
nor U22714 (N_22714,N_21975,N_22045);
nand U22715 (N_22715,N_21974,N_22193);
and U22716 (N_22716,N_21998,N_22133);
and U22717 (N_22717,N_22330,N_21920);
xor U22718 (N_22718,N_22103,N_22271);
nand U22719 (N_22719,N_22318,N_22320);
and U22720 (N_22720,N_21977,N_22061);
or U22721 (N_22721,N_22071,N_22132);
and U22722 (N_22722,N_22301,N_22357);
and U22723 (N_22723,N_22231,N_22095);
xor U22724 (N_22724,N_22358,N_22428);
nand U22725 (N_22725,N_22197,N_22326);
nand U22726 (N_22726,N_22398,N_22262);
or U22727 (N_22727,N_22283,N_22100);
nor U22728 (N_22728,N_22453,N_21948);
and U22729 (N_22729,N_22228,N_22157);
nor U22730 (N_22730,N_22126,N_21915);
nor U22731 (N_22731,N_22230,N_22038);
and U22732 (N_22732,N_22346,N_22285);
nand U22733 (N_22733,N_22187,N_22244);
and U22734 (N_22734,N_22104,N_21886);
or U22735 (N_22735,N_22060,N_22081);
nand U22736 (N_22736,N_21938,N_22406);
xnor U22737 (N_22737,N_22206,N_22027);
or U22738 (N_22738,N_22376,N_22189);
or U22739 (N_22739,N_22181,N_22288);
nand U22740 (N_22740,N_21916,N_22047);
and U22741 (N_22741,N_22096,N_22094);
nand U22742 (N_22742,N_21878,N_22235);
xnor U22743 (N_22743,N_22327,N_21919);
and U22744 (N_22744,N_22140,N_22415);
nor U22745 (N_22745,N_21991,N_21898);
or U22746 (N_22746,N_22446,N_22256);
and U22747 (N_22747,N_22148,N_22407);
or U22748 (N_22748,N_21943,N_22417);
nand U22749 (N_22749,N_22205,N_22116);
and U22750 (N_22750,N_22015,N_22269);
xnor U22751 (N_22751,N_22260,N_22088);
nand U22752 (N_22752,N_22137,N_22074);
and U22753 (N_22753,N_22085,N_22044);
nand U22754 (N_22754,N_22429,N_22086);
nor U22755 (N_22755,N_21922,N_21884);
or U22756 (N_22756,N_21887,N_21939);
nand U22757 (N_22757,N_22267,N_22309);
nand U22758 (N_22758,N_22166,N_22216);
or U22759 (N_22759,N_22494,N_22236);
nand U22760 (N_22760,N_22249,N_21970);
nand U22761 (N_22761,N_22067,N_22127);
nand U22762 (N_22762,N_22125,N_22399);
and U22763 (N_22763,N_22008,N_22114);
nor U22764 (N_22764,N_22261,N_22422);
or U22765 (N_22765,N_22057,N_22403);
nor U22766 (N_22766,N_22090,N_22208);
and U22767 (N_22767,N_21946,N_21928);
xnor U22768 (N_22768,N_22076,N_21895);
nor U22769 (N_22769,N_22290,N_22447);
and U22770 (N_22770,N_22270,N_22324);
and U22771 (N_22771,N_21894,N_21959);
and U22772 (N_22772,N_21992,N_22024);
and U22773 (N_22773,N_21926,N_21968);
and U22774 (N_22774,N_21952,N_22414);
nand U22775 (N_22775,N_21893,N_22072);
or U22776 (N_22776,N_22333,N_21907);
or U22777 (N_22777,N_22176,N_22122);
xor U22778 (N_22778,N_22180,N_21964);
xor U22779 (N_22779,N_21925,N_22240);
nand U22780 (N_22780,N_22279,N_22084);
nand U22781 (N_22781,N_22397,N_22312);
nor U22782 (N_22782,N_22190,N_22341);
nor U22783 (N_22783,N_21905,N_22388);
xnor U22784 (N_22784,N_22033,N_22390);
or U22785 (N_22785,N_22391,N_22105);
nand U22786 (N_22786,N_21902,N_22093);
or U22787 (N_22787,N_22218,N_22400);
or U22788 (N_22788,N_22455,N_22313);
or U22789 (N_22789,N_22322,N_22167);
nor U22790 (N_22790,N_22192,N_21906);
and U22791 (N_22791,N_21947,N_21993);
xor U22792 (N_22792,N_22194,N_22449);
nor U22793 (N_22793,N_22113,N_22202);
or U22794 (N_22794,N_22420,N_22338);
and U22795 (N_22795,N_21983,N_22077);
and U22796 (N_22796,N_22347,N_21941);
nor U22797 (N_22797,N_22214,N_22130);
or U22798 (N_22798,N_22448,N_22025);
nor U22799 (N_22799,N_22041,N_22462);
and U22800 (N_22800,N_22237,N_22242);
nor U22801 (N_22801,N_22054,N_22484);
nor U22802 (N_22802,N_22436,N_21889);
nor U22803 (N_22803,N_22158,N_22102);
and U22804 (N_22804,N_22413,N_22035);
xnor U22805 (N_22805,N_22178,N_21882);
nor U22806 (N_22806,N_22383,N_22451);
and U22807 (N_22807,N_22101,N_22141);
or U22808 (N_22808,N_22426,N_21936);
nand U22809 (N_22809,N_22149,N_22307);
or U22810 (N_22810,N_21875,N_22263);
or U22811 (N_22811,N_22210,N_21885);
or U22812 (N_22812,N_22394,N_22346);
xnor U22813 (N_22813,N_22471,N_22443);
nand U22814 (N_22814,N_21960,N_22102);
and U22815 (N_22815,N_21997,N_22339);
and U22816 (N_22816,N_22029,N_22228);
or U22817 (N_22817,N_22145,N_22231);
and U22818 (N_22818,N_21894,N_22207);
nand U22819 (N_22819,N_22439,N_22396);
nor U22820 (N_22820,N_22281,N_22063);
and U22821 (N_22821,N_22052,N_21955);
nor U22822 (N_22822,N_22455,N_21942);
nand U22823 (N_22823,N_22466,N_22341);
xnor U22824 (N_22824,N_22389,N_22114);
and U22825 (N_22825,N_22341,N_22405);
nor U22826 (N_22826,N_22200,N_22182);
or U22827 (N_22827,N_22313,N_22220);
or U22828 (N_22828,N_22134,N_22302);
xnor U22829 (N_22829,N_22286,N_22074);
nand U22830 (N_22830,N_22386,N_22184);
nor U22831 (N_22831,N_22490,N_22390);
nor U22832 (N_22832,N_22236,N_22200);
or U22833 (N_22833,N_22454,N_22328);
xnor U22834 (N_22834,N_21912,N_22166);
or U22835 (N_22835,N_21942,N_22084);
nand U22836 (N_22836,N_22478,N_22429);
and U22837 (N_22837,N_21949,N_22090);
or U22838 (N_22838,N_22195,N_22194);
or U22839 (N_22839,N_22444,N_22111);
nand U22840 (N_22840,N_21981,N_22346);
nor U22841 (N_22841,N_22234,N_21929);
nor U22842 (N_22842,N_22132,N_22453);
nor U22843 (N_22843,N_22096,N_22492);
and U22844 (N_22844,N_22443,N_22141);
nand U22845 (N_22845,N_22440,N_22027);
and U22846 (N_22846,N_22436,N_21965);
xnor U22847 (N_22847,N_21961,N_22228);
nor U22848 (N_22848,N_22090,N_22078);
or U22849 (N_22849,N_22289,N_22400);
and U22850 (N_22850,N_22287,N_22369);
or U22851 (N_22851,N_22144,N_22447);
or U22852 (N_22852,N_22047,N_22329);
xor U22853 (N_22853,N_22147,N_22123);
and U22854 (N_22854,N_22401,N_22295);
and U22855 (N_22855,N_22474,N_22237);
and U22856 (N_22856,N_21888,N_22063);
nand U22857 (N_22857,N_22086,N_22258);
xnor U22858 (N_22858,N_22186,N_22033);
and U22859 (N_22859,N_21944,N_22281);
or U22860 (N_22860,N_21986,N_21997);
and U22861 (N_22861,N_22376,N_22084);
or U22862 (N_22862,N_21936,N_22287);
or U22863 (N_22863,N_21952,N_22407);
or U22864 (N_22864,N_22178,N_22001);
and U22865 (N_22865,N_22212,N_21912);
xor U22866 (N_22866,N_21941,N_22378);
nand U22867 (N_22867,N_22496,N_22000);
or U22868 (N_22868,N_22304,N_22251);
or U22869 (N_22869,N_22068,N_22246);
or U22870 (N_22870,N_22253,N_22002);
or U22871 (N_22871,N_22416,N_21880);
or U22872 (N_22872,N_22211,N_22357);
nand U22873 (N_22873,N_22400,N_22388);
nand U22874 (N_22874,N_22434,N_22485);
nand U22875 (N_22875,N_22013,N_22170);
nor U22876 (N_22876,N_21886,N_22127);
or U22877 (N_22877,N_22167,N_22490);
xor U22878 (N_22878,N_22488,N_22425);
nand U22879 (N_22879,N_22360,N_22463);
xnor U22880 (N_22880,N_21960,N_22454);
nand U22881 (N_22881,N_21888,N_22003);
nand U22882 (N_22882,N_22007,N_22117);
and U22883 (N_22883,N_22140,N_22449);
nand U22884 (N_22884,N_21915,N_22244);
nor U22885 (N_22885,N_22116,N_22135);
and U22886 (N_22886,N_22171,N_22193);
and U22887 (N_22887,N_22147,N_22405);
nand U22888 (N_22888,N_22021,N_22110);
xnor U22889 (N_22889,N_22042,N_22159);
and U22890 (N_22890,N_22356,N_22164);
and U22891 (N_22891,N_22130,N_22179);
or U22892 (N_22892,N_22407,N_22124);
nand U22893 (N_22893,N_22192,N_22276);
and U22894 (N_22894,N_22309,N_22299);
nor U22895 (N_22895,N_22330,N_22185);
nor U22896 (N_22896,N_22165,N_22301);
or U22897 (N_22897,N_22442,N_22304);
and U22898 (N_22898,N_21888,N_22386);
nor U22899 (N_22899,N_22027,N_22323);
nand U22900 (N_22900,N_22113,N_22354);
nand U22901 (N_22901,N_22416,N_22000);
or U22902 (N_22902,N_22331,N_22316);
nor U22903 (N_22903,N_22240,N_22140);
and U22904 (N_22904,N_22352,N_22063);
nor U22905 (N_22905,N_22284,N_22078);
nand U22906 (N_22906,N_22370,N_22411);
and U22907 (N_22907,N_21903,N_22003);
nor U22908 (N_22908,N_21878,N_22434);
nand U22909 (N_22909,N_22238,N_21986);
nand U22910 (N_22910,N_22140,N_21934);
or U22911 (N_22911,N_22468,N_22250);
nor U22912 (N_22912,N_22094,N_22495);
nand U22913 (N_22913,N_21896,N_22020);
or U22914 (N_22914,N_22102,N_22414);
nor U22915 (N_22915,N_22098,N_22118);
nand U22916 (N_22916,N_21893,N_22465);
nand U22917 (N_22917,N_22232,N_22139);
nor U22918 (N_22918,N_22083,N_22081);
xor U22919 (N_22919,N_22478,N_22008);
nor U22920 (N_22920,N_21979,N_22202);
and U22921 (N_22921,N_22007,N_22358);
or U22922 (N_22922,N_21889,N_21930);
nor U22923 (N_22923,N_21956,N_22151);
nand U22924 (N_22924,N_22129,N_22489);
nand U22925 (N_22925,N_22358,N_21889);
nand U22926 (N_22926,N_22331,N_22305);
and U22927 (N_22927,N_22167,N_22462);
or U22928 (N_22928,N_22283,N_22026);
and U22929 (N_22929,N_21892,N_21951);
and U22930 (N_22930,N_22179,N_21917);
nand U22931 (N_22931,N_22499,N_21988);
xor U22932 (N_22932,N_22072,N_22140);
nand U22933 (N_22933,N_22156,N_22219);
and U22934 (N_22934,N_22193,N_22315);
nor U22935 (N_22935,N_22463,N_22215);
nand U22936 (N_22936,N_22452,N_22119);
and U22937 (N_22937,N_22103,N_22163);
and U22938 (N_22938,N_22139,N_22065);
and U22939 (N_22939,N_22496,N_22403);
or U22940 (N_22940,N_22238,N_21965);
or U22941 (N_22941,N_22261,N_22367);
nor U22942 (N_22942,N_22121,N_22466);
nand U22943 (N_22943,N_22280,N_22040);
or U22944 (N_22944,N_22275,N_22171);
xnor U22945 (N_22945,N_22160,N_21908);
nand U22946 (N_22946,N_22091,N_22244);
nor U22947 (N_22947,N_22184,N_22346);
or U22948 (N_22948,N_22324,N_22069);
nor U22949 (N_22949,N_21890,N_22338);
or U22950 (N_22950,N_21941,N_21898);
nand U22951 (N_22951,N_22417,N_21947);
xnor U22952 (N_22952,N_22355,N_22172);
nor U22953 (N_22953,N_22054,N_21974);
xor U22954 (N_22954,N_22451,N_22124);
or U22955 (N_22955,N_22430,N_22200);
xor U22956 (N_22956,N_22137,N_22308);
nand U22957 (N_22957,N_21932,N_22177);
xnor U22958 (N_22958,N_21906,N_22138);
or U22959 (N_22959,N_22232,N_22043);
and U22960 (N_22960,N_22241,N_22097);
and U22961 (N_22961,N_22307,N_22346);
nand U22962 (N_22962,N_22468,N_22474);
or U22963 (N_22963,N_22331,N_22063);
and U22964 (N_22964,N_22055,N_22371);
and U22965 (N_22965,N_22156,N_21921);
or U22966 (N_22966,N_22493,N_22061);
and U22967 (N_22967,N_22399,N_22484);
nand U22968 (N_22968,N_22030,N_21876);
or U22969 (N_22969,N_21878,N_22234);
and U22970 (N_22970,N_22064,N_22314);
xor U22971 (N_22971,N_22293,N_21951);
and U22972 (N_22972,N_22284,N_22414);
nor U22973 (N_22973,N_22027,N_22380);
nor U22974 (N_22974,N_22327,N_22136);
xnor U22975 (N_22975,N_22193,N_22463);
and U22976 (N_22976,N_21944,N_21991);
and U22977 (N_22977,N_22065,N_22014);
or U22978 (N_22978,N_22278,N_21884);
nand U22979 (N_22979,N_22268,N_22344);
and U22980 (N_22980,N_22050,N_21969);
or U22981 (N_22981,N_22083,N_22309);
or U22982 (N_22982,N_22031,N_22362);
nand U22983 (N_22983,N_22389,N_21923);
or U22984 (N_22984,N_22485,N_22234);
nand U22985 (N_22985,N_22275,N_22366);
nand U22986 (N_22986,N_22233,N_21901);
nor U22987 (N_22987,N_22457,N_22485);
nand U22988 (N_22988,N_22260,N_22322);
or U22989 (N_22989,N_22106,N_22392);
or U22990 (N_22990,N_21952,N_22243);
nor U22991 (N_22991,N_21887,N_22116);
and U22992 (N_22992,N_22018,N_22453);
or U22993 (N_22993,N_22201,N_22316);
nand U22994 (N_22994,N_22273,N_22062);
xnor U22995 (N_22995,N_22383,N_22104);
nor U22996 (N_22996,N_22467,N_21964);
and U22997 (N_22997,N_22044,N_22211);
or U22998 (N_22998,N_22236,N_22483);
nor U22999 (N_22999,N_21938,N_22447);
nor U23000 (N_23000,N_22115,N_21877);
nor U23001 (N_23001,N_22375,N_21988);
or U23002 (N_23002,N_21886,N_22008);
nand U23003 (N_23003,N_22250,N_22022);
and U23004 (N_23004,N_22230,N_22064);
nand U23005 (N_23005,N_22297,N_22124);
nand U23006 (N_23006,N_22005,N_22046);
nor U23007 (N_23007,N_21997,N_21968);
or U23008 (N_23008,N_22463,N_22192);
or U23009 (N_23009,N_22388,N_22145);
xnor U23010 (N_23010,N_22317,N_22220);
nand U23011 (N_23011,N_22356,N_22134);
nor U23012 (N_23012,N_22218,N_22127);
or U23013 (N_23013,N_21973,N_22181);
or U23014 (N_23014,N_22344,N_22252);
nand U23015 (N_23015,N_22492,N_22475);
nor U23016 (N_23016,N_22488,N_22394);
nand U23017 (N_23017,N_22137,N_22202);
nor U23018 (N_23018,N_22112,N_22412);
nand U23019 (N_23019,N_22178,N_22402);
nand U23020 (N_23020,N_22230,N_21997);
xnor U23021 (N_23021,N_21913,N_22049);
nor U23022 (N_23022,N_22027,N_22247);
nor U23023 (N_23023,N_21986,N_22020);
nor U23024 (N_23024,N_22434,N_22477);
nor U23025 (N_23025,N_22142,N_22387);
nand U23026 (N_23026,N_22297,N_22319);
nand U23027 (N_23027,N_22263,N_22165);
nand U23028 (N_23028,N_22278,N_22104);
and U23029 (N_23029,N_21950,N_22306);
xor U23030 (N_23030,N_21923,N_21931);
nand U23031 (N_23031,N_22458,N_22215);
nand U23032 (N_23032,N_22226,N_22469);
nand U23033 (N_23033,N_22354,N_22088);
nor U23034 (N_23034,N_22316,N_22441);
nor U23035 (N_23035,N_21947,N_22249);
or U23036 (N_23036,N_22098,N_22442);
or U23037 (N_23037,N_22333,N_22473);
or U23038 (N_23038,N_22134,N_22174);
nand U23039 (N_23039,N_21973,N_22269);
and U23040 (N_23040,N_21920,N_22334);
and U23041 (N_23041,N_22350,N_21891);
or U23042 (N_23042,N_22357,N_21950);
nand U23043 (N_23043,N_22337,N_22415);
nor U23044 (N_23044,N_22342,N_21881);
and U23045 (N_23045,N_22184,N_22024);
or U23046 (N_23046,N_22011,N_22058);
or U23047 (N_23047,N_22452,N_22252);
nor U23048 (N_23048,N_22377,N_21984);
and U23049 (N_23049,N_22192,N_21990);
and U23050 (N_23050,N_22116,N_22109);
nor U23051 (N_23051,N_22461,N_22333);
xor U23052 (N_23052,N_21911,N_21948);
or U23053 (N_23053,N_22203,N_22342);
nor U23054 (N_23054,N_21948,N_22492);
nor U23055 (N_23055,N_22008,N_22136);
nand U23056 (N_23056,N_22342,N_22335);
and U23057 (N_23057,N_22431,N_22294);
nor U23058 (N_23058,N_22491,N_22268);
and U23059 (N_23059,N_22165,N_21969);
or U23060 (N_23060,N_22322,N_22030);
or U23061 (N_23061,N_22069,N_22494);
xor U23062 (N_23062,N_22372,N_22344);
nor U23063 (N_23063,N_22173,N_22000);
nor U23064 (N_23064,N_22347,N_22334);
or U23065 (N_23065,N_22459,N_22376);
xnor U23066 (N_23066,N_22103,N_22145);
and U23067 (N_23067,N_22277,N_22289);
nor U23068 (N_23068,N_21920,N_22475);
xnor U23069 (N_23069,N_22361,N_22477);
nor U23070 (N_23070,N_22325,N_22236);
nand U23071 (N_23071,N_21889,N_22252);
xnor U23072 (N_23072,N_22442,N_22047);
xor U23073 (N_23073,N_22428,N_22434);
xor U23074 (N_23074,N_22384,N_22310);
nor U23075 (N_23075,N_22030,N_22063);
xor U23076 (N_23076,N_22049,N_21985);
and U23077 (N_23077,N_22332,N_22355);
nor U23078 (N_23078,N_22456,N_22382);
nor U23079 (N_23079,N_22030,N_22083);
nand U23080 (N_23080,N_22106,N_21881);
nand U23081 (N_23081,N_22064,N_21888);
or U23082 (N_23082,N_22130,N_22222);
and U23083 (N_23083,N_22012,N_22133);
nor U23084 (N_23084,N_21886,N_22466);
xor U23085 (N_23085,N_22163,N_22487);
nand U23086 (N_23086,N_22259,N_21996);
nand U23087 (N_23087,N_22273,N_21879);
nand U23088 (N_23088,N_22171,N_22315);
nor U23089 (N_23089,N_22405,N_22175);
or U23090 (N_23090,N_21890,N_22375);
xor U23091 (N_23091,N_22009,N_22120);
xor U23092 (N_23092,N_22336,N_22364);
or U23093 (N_23093,N_22022,N_21891);
nor U23094 (N_23094,N_21926,N_22233);
nand U23095 (N_23095,N_21919,N_22299);
nor U23096 (N_23096,N_22004,N_21892);
or U23097 (N_23097,N_22019,N_22191);
nor U23098 (N_23098,N_22184,N_22342);
nand U23099 (N_23099,N_22401,N_22379);
xor U23100 (N_23100,N_22485,N_22277);
xnor U23101 (N_23101,N_21937,N_22287);
nor U23102 (N_23102,N_22000,N_22085);
and U23103 (N_23103,N_22491,N_22279);
nor U23104 (N_23104,N_22478,N_22230);
nor U23105 (N_23105,N_22332,N_22194);
nor U23106 (N_23106,N_22320,N_22397);
nand U23107 (N_23107,N_22376,N_22299);
nor U23108 (N_23108,N_22231,N_22281);
nor U23109 (N_23109,N_22100,N_22351);
nand U23110 (N_23110,N_21921,N_21979);
and U23111 (N_23111,N_22125,N_22438);
nand U23112 (N_23112,N_22294,N_22101);
nand U23113 (N_23113,N_22431,N_22115);
and U23114 (N_23114,N_22241,N_22329);
and U23115 (N_23115,N_22115,N_22216);
nand U23116 (N_23116,N_22308,N_22071);
nor U23117 (N_23117,N_22360,N_22019);
or U23118 (N_23118,N_22175,N_22057);
nor U23119 (N_23119,N_22161,N_22422);
nand U23120 (N_23120,N_22383,N_22480);
nor U23121 (N_23121,N_22400,N_22394);
and U23122 (N_23122,N_22017,N_22157);
or U23123 (N_23123,N_22383,N_22227);
or U23124 (N_23124,N_22491,N_22255);
or U23125 (N_23125,N_22837,N_22566);
or U23126 (N_23126,N_22900,N_22869);
or U23127 (N_23127,N_22724,N_22942);
xnor U23128 (N_23128,N_23010,N_23042);
or U23129 (N_23129,N_22635,N_22644);
xor U23130 (N_23130,N_22736,N_22611);
and U23131 (N_23131,N_22512,N_23069);
nor U23132 (N_23132,N_22692,N_23014);
and U23133 (N_23133,N_22698,N_22506);
and U23134 (N_23134,N_23076,N_22679);
nand U23135 (N_23135,N_22632,N_22733);
nor U23136 (N_23136,N_22553,N_22822);
or U23137 (N_23137,N_22951,N_22538);
or U23138 (N_23138,N_22815,N_22569);
nand U23139 (N_23139,N_22563,N_22818);
or U23140 (N_23140,N_23025,N_22661);
and U23141 (N_23141,N_22691,N_22988);
nand U23142 (N_23142,N_22609,N_22823);
or U23143 (N_23143,N_22825,N_22990);
and U23144 (N_23144,N_22802,N_22849);
and U23145 (N_23145,N_22788,N_22856);
nor U23146 (N_23146,N_22547,N_22540);
xor U23147 (N_23147,N_22713,N_22941);
xnor U23148 (N_23148,N_22916,N_22722);
and U23149 (N_23149,N_23079,N_22574);
xnor U23150 (N_23150,N_22675,N_23034);
nor U23151 (N_23151,N_22643,N_22863);
nand U23152 (N_23152,N_23098,N_23011);
or U23153 (N_23153,N_22639,N_22575);
nand U23154 (N_23154,N_22517,N_22545);
or U23155 (N_23155,N_22687,N_22748);
nand U23156 (N_23156,N_22721,N_22752);
nand U23157 (N_23157,N_22972,N_22804);
nor U23158 (N_23158,N_23001,N_22896);
nand U23159 (N_23159,N_22854,N_22688);
and U23160 (N_23160,N_22555,N_22511);
nor U23161 (N_23161,N_22989,N_22557);
nor U23162 (N_23162,N_22806,N_22562);
and U23163 (N_23163,N_22992,N_23081);
and U23164 (N_23164,N_23045,N_22646);
nor U23165 (N_23165,N_22925,N_22979);
or U23166 (N_23166,N_22875,N_22515);
nand U23167 (N_23167,N_23036,N_22514);
and U23168 (N_23168,N_22743,N_22626);
or U23169 (N_23169,N_23047,N_22791);
nor U23170 (N_23170,N_23080,N_23095);
and U23171 (N_23171,N_23029,N_22573);
or U23172 (N_23172,N_22812,N_22607);
and U23173 (N_23173,N_23055,N_23090);
and U23174 (N_23174,N_22739,N_22922);
or U23175 (N_23175,N_22530,N_22910);
xnor U23176 (N_23176,N_22581,N_22582);
nor U23177 (N_23177,N_23088,N_23005);
and U23178 (N_23178,N_22982,N_22872);
or U23179 (N_23179,N_22807,N_22765);
nor U23180 (N_23180,N_22954,N_22940);
nand U23181 (N_23181,N_22923,N_22543);
nand U23182 (N_23182,N_22795,N_23075);
and U23183 (N_23183,N_23065,N_22882);
nand U23184 (N_23184,N_22985,N_22601);
nor U23185 (N_23185,N_22732,N_22873);
and U23186 (N_23186,N_22755,N_22668);
nor U23187 (N_23187,N_22667,N_23041);
or U23188 (N_23188,N_22997,N_23031);
and U23189 (N_23189,N_22741,N_22546);
nor U23190 (N_23190,N_23062,N_22513);
or U23191 (N_23191,N_22917,N_22583);
nand U23192 (N_23192,N_23097,N_22636);
nor U23193 (N_23193,N_23108,N_23051);
nor U23194 (N_23194,N_22758,N_22783);
nand U23195 (N_23195,N_23017,N_22851);
nor U23196 (N_23196,N_23089,N_23121);
or U23197 (N_23197,N_22571,N_22831);
or U23198 (N_23198,N_22544,N_22949);
nand U23199 (N_23199,N_22664,N_22966);
and U23200 (N_23200,N_22728,N_22535);
nand U23201 (N_23201,N_22684,N_22857);
nor U23202 (N_23202,N_22836,N_22706);
or U23203 (N_23203,N_22630,N_22671);
nand U23204 (N_23204,N_22803,N_22805);
or U23205 (N_23205,N_23072,N_22669);
xor U23206 (N_23206,N_22879,N_23087);
nand U23207 (N_23207,N_22683,N_22508);
or U23208 (N_23208,N_22919,N_22766);
nor U23209 (N_23209,N_23120,N_23049);
or U23210 (N_23210,N_22572,N_22811);
and U23211 (N_23211,N_22880,N_23105);
or U23212 (N_23212,N_22763,N_22701);
xor U23213 (N_23213,N_22974,N_22981);
nand U23214 (N_23214,N_23033,N_23030);
nor U23215 (N_23215,N_23022,N_22786);
and U23216 (N_23216,N_22693,N_22780);
or U23217 (N_23217,N_23000,N_22702);
xnor U23218 (N_23218,N_22595,N_22767);
nand U23219 (N_23219,N_23052,N_23114);
xor U23220 (N_23220,N_23053,N_22907);
nand U23221 (N_23221,N_22887,N_22821);
and U23222 (N_23222,N_23091,N_22745);
nand U23223 (N_23223,N_23019,N_22850);
nand U23224 (N_23224,N_22648,N_22604);
nor U23225 (N_23225,N_23018,N_22817);
nor U23226 (N_23226,N_22605,N_22936);
or U23227 (N_23227,N_23106,N_23060);
xnor U23228 (N_23228,N_22772,N_23123);
nand U23229 (N_23229,N_23073,N_22841);
nor U23230 (N_23230,N_22777,N_22623);
nand U23231 (N_23231,N_22677,N_22962);
or U23232 (N_23232,N_22738,N_22799);
and U23233 (N_23233,N_22602,N_22507);
and U23234 (N_23234,N_23103,N_22603);
or U23235 (N_23235,N_22600,N_22718);
nand U23236 (N_23236,N_22933,N_22678);
nand U23237 (N_23237,N_22889,N_22897);
nand U23238 (N_23238,N_22835,N_22510);
nor U23239 (N_23239,N_22531,N_22820);
nand U23240 (N_23240,N_23124,N_22958);
or U23241 (N_23241,N_22627,N_22565);
nand U23242 (N_23242,N_22696,N_22534);
nand U23243 (N_23243,N_22610,N_22628);
nor U23244 (N_23244,N_22700,N_22971);
or U23245 (N_23245,N_22935,N_22924);
or U23246 (N_23246,N_23084,N_22580);
nand U23247 (N_23247,N_22541,N_22597);
or U23248 (N_23248,N_22893,N_22524);
nand U23249 (N_23249,N_23006,N_22877);
nor U23250 (N_23250,N_23077,N_22899);
or U23251 (N_23251,N_22537,N_23064);
or U23252 (N_23252,N_23093,N_23015);
and U23253 (N_23253,N_22797,N_22902);
nor U23254 (N_23254,N_22742,N_22699);
and U23255 (N_23255,N_22542,N_22930);
xnor U23256 (N_23256,N_22614,N_23050);
or U23257 (N_23257,N_22686,N_22615);
xnor U23258 (N_23258,N_22593,N_22960);
nand U23259 (N_23259,N_22551,N_22659);
nor U23260 (N_23260,N_22697,N_22734);
or U23261 (N_23261,N_23061,N_23119);
and U23262 (N_23262,N_22654,N_22918);
nor U23263 (N_23263,N_22640,N_22726);
xor U23264 (N_23264,N_23044,N_22584);
nor U23265 (N_23265,N_22596,N_23054);
or U23266 (N_23266,N_22682,N_22898);
nor U23267 (N_23267,N_22859,N_22874);
and U23268 (N_23268,N_22764,N_22525);
nor U23269 (N_23269,N_23099,N_23104);
nand U23270 (N_23270,N_23026,N_23122);
nor U23271 (N_23271,N_23043,N_22860);
and U23272 (N_23272,N_22550,N_22529);
nand U23273 (N_23273,N_22886,N_22617);
and U23274 (N_23274,N_22946,N_22800);
and U23275 (N_23275,N_22968,N_22681);
nor U23276 (N_23276,N_22503,N_22782);
and U23277 (N_23277,N_22599,N_23063);
or U23278 (N_23278,N_22528,N_22618);
nand U23279 (N_23279,N_22754,N_22865);
and U23280 (N_23280,N_22789,N_22901);
or U23281 (N_23281,N_22526,N_22913);
and U23282 (N_23282,N_22813,N_22578);
or U23283 (N_23283,N_22711,N_22650);
xnor U23284 (N_23284,N_22921,N_23048);
nor U23285 (N_23285,N_22554,N_22839);
nor U23286 (N_23286,N_22756,N_22939);
and U23287 (N_23287,N_23059,N_22883);
xnor U23288 (N_23288,N_22827,N_22908);
and U23289 (N_23289,N_22927,N_22703);
or U23290 (N_23290,N_22660,N_22655);
xor U23291 (N_23291,N_22533,N_23021);
or U23292 (N_23292,N_22751,N_22714);
nand U23293 (N_23293,N_22621,N_22613);
or U23294 (N_23294,N_22991,N_22967);
and U23295 (N_23295,N_22852,N_22505);
nor U23296 (N_23296,N_22504,N_22984);
nor U23297 (N_23297,N_22938,N_23007);
nand U23298 (N_23298,N_22964,N_22931);
nor U23299 (N_23299,N_22824,N_22846);
and U23300 (N_23300,N_22568,N_22536);
nor U23301 (N_23301,N_22976,N_22769);
nor U23302 (N_23302,N_23115,N_23038);
nor U23303 (N_23303,N_22816,N_23102);
and U23304 (N_23304,N_22830,N_22905);
or U23305 (N_23305,N_22522,N_22776);
or U23306 (N_23306,N_23012,N_23113);
and U23307 (N_23307,N_23068,N_22729);
nand U23308 (N_23308,N_22892,N_22556);
nand U23309 (N_23309,N_22548,N_22651);
nand U23310 (N_23310,N_22674,N_22740);
or U23311 (N_23311,N_22787,N_22987);
and U23312 (N_23312,N_22737,N_22768);
or U23313 (N_23313,N_22774,N_22832);
nor U23314 (N_23314,N_22624,N_22727);
and U23315 (N_23315,N_23037,N_22868);
or U23316 (N_23316,N_23056,N_22956);
xnor U23317 (N_23317,N_22619,N_23111);
nand U23318 (N_23318,N_22770,N_22871);
xnor U23319 (N_23319,N_23040,N_22500);
and U23320 (N_23320,N_22773,N_22878);
nor U23321 (N_23321,N_22999,N_22712);
nand U23322 (N_23322,N_23094,N_22761);
nor U23323 (N_23323,N_22746,N_22502);
or U23324 (N_23324,N_22666,N_22558);
nor U23325 (N_23325,N_23071,N_23066);
and U23326 (N_23326,N_22663,N_22749);
nor U23327 (N_23327,N_23027,N_23058);
nand U23328 (N_23328,N_22784,N_22523);
nor U23329 (N_23329,N_23085,N_22590);
nand U23330 (N_23330,N_22915,N_22779);
and U23331 (N_23331,N_22649,N_23035);
nor U23332 (N_23332,N_23092,N_22567);
xor U23333 (N_23333,N_22520,N_23046);
nand U23334 (N_23334,N_22785,N_22808);
or U23335 (N_23335,N_23003,N_23070);
nor U23336 (N_23336,N_23008,N_22828);
or U23337 (N_23337,N_22759,N_22670);
or U23338 (N_23338,N_22676,N_22909);
or U23339 (N_23339,N_22680,N_22929);
nand U23340 (N_23340,N_22570,N_22801);
or U23341 (N_23341,N_22589,N_23110);
or U23342 (N_23342,N_23118,N_22980);
nand U23343 (N_23343,N_22906,N_22973);
nand U23344 (N_23344,N_22716,N_22564);
nor U23345 (N_23345,N_22717,N_22744);
nor U23346 (N_23346,N_22620,N_22559);
nor U23347 (N_23347,N_22634,N_22945);
or U23348 (N_23348,N_22731,N_22842);
nor U23349 (N_23349,N_22920,N_22689);
and U23350 (N_23350,N_22519,N_22955);
nor U23351 (N_23351,N_22895,N_23002);
and U23352 (N_23352,N_22747,N_22709);
and U23353 (N_23353,N_23023,N_22993);
and U23354 (N_23354,N_22735,N_22793);
nand U23355 (N_23355,N_22598,N_22961);
xor U23356 (N_23356,N_22750,N_22986);
xnor U23357 (N_23357,N_22652,N_22876);
or U23358 (N_23358,N_22965,N_22778);
and U23359 (N_23359,N_22638,N_22969);
and U23360 (N_23360,N_23112,N_22994);
nor U23361 (N_23361,N_22707,N_22995);
nor U23362 (N_23362,N_22608,N_22685);
xnor U23363 (N_23363,N_22588,N_22890);
nor U23364 (N_23364,N_23057,N_22794);
or U23365 (N_23365,N_22975,N_22844);
nand U23366 (N_23366,N_22587,N_22633);
xnor U23367 (N_23367,N_22723,N_23013);
or U23368 (N_23368,N_22937,N_23078);
nand U23369 (N_23369,N_23067,N_23109);
or U23370 (N_23370,N_22532,N_22911);
nand U23371 (N_23371,N_23096,N_22864);
and U23372 (N_23372,N_23107,N_22586);
or U23373 (N_23373,N_22781,N_22710);
xnor U23374 (N_23374,N_23117,N_22527);
nor U23375 (N_23375,N_22725,N_22792);
nor U23376 (N_23376,N_22862,N_22577);
and U23377 (N_23377,N_22957,N_22891);
and U23378 (N_23378,N_22591,N_22539);
or U23379 (N_23379,N_22673,N_22653);
xnor U23380 (N_23380,N_22730,N_22845);
and U23381 (N_23381,N_22855,N_22848);
nand U23382 (N_23382,N_23100,N_22977);
nor U23383 (N_23383,N_22509,N_22983);
and U23384 (N_23384,N_22826,N_22561);
nor U23385 (N_23385,N_23083,N_22616);
nand U23386 (N_23386,N_22959,N_22625);
and U23387 (N_23387,N_23020,N_22885);
nor U23388 (N_23388,N_22771,N_22829);
or U23389 (N_23389,N_22810,N_22847);
or U23390 (N_23390,N_22704,N_22978);
and U23391 (N_23391,N_22858,N_22775);
nor U23392 (N_23392,N_22833,N_23116);
and U23393 (N_23393,N_23082,N_22762);
or U23394 (N_23394,N_22884,N_22943);
nand U23395 (N_23395,N_22903,N_22690);
nor U23396 (N_23396,N_22612,N_22861);
or U23397 (N_23397,N_22594,N_22658);
and U23398 (N_23398,N_22870,N_22708);
and U23399 (N_23399,N_22888,N_22576);
or U23400 (N_23400,N_22894,N_23039);
and U23401 (N_23401,N_22867,N_22970);
or U23402 (N_23402,N_22926,N_22952);
and U23403 (N_23403,N_22552,N_22996);
nor U23404 (N_23404,N_22622,N_23101);
or U23405 (N_23405,N_22705,N_22695);
nor U23406 (N_23406,N_23032,N_22672);
or U23407 (N_23407,N_22518,N_22760);
nor U23408 (N_23408,N_23009,N_22928);
and U23409 (N_23409,N_22656,N_22840);
or U23410 (N_23410,N_22715,N_22866);
nand U23411 (N_23411,N_23004,N_22665);
nand U23412 (N_23412,N_22834,N_22516);
xor U23413 (N_23413,N_22645,N_22814);
and U23414 (N_23414,N_22932,N_22819);
or U23415 (N_23415,N_22753,N_22881);
and U23416 (N_23416,N_22796,N_22998);
or U23417 (N_23417,N_22647,N_23028);
xnor U23418 (N_23418,N_22579,N_22719);
nand U23419 (N_23419,N_22904,N_22798);
or U23420 (N_23420,N_22934,N_22790);
or U23421 (N_23421,N_22501,N_22947);
nor U23422 (N_23422,N_22662,N_22585);
and U23423 (N_23423,N_23024,N_22838);
nand U23424 (N_23424,N_22720,N_22950);
nor U23425 (N_23425,N_22521,N_22944);
and U23426 (N_23426,N_22843,N_22757);
or U23427 (N_23427,N_22549,N_23016);
nand U23428 (N_23428,N_22657,N_23074);
or U23429 (N_23429,N_22853,N_22631);
or U23430 (N_23430,N_22606,N_22914);
or U23431 (N_23431,N_22809,N_22963);
and U23432 (N_23432,N_22642,N_23086);
xnor U23433 (N_23433,N_22912,N_22694);
or U23434 (N_23434,N_22953,N_22592);
nand U23435 (N_23435,N_22948,N_22637);
and U23436 (N_23436,N_22560,N_22641);
nor U23437 (N_23437,N_22629,N_22991);
or U23438 (N_23438,N_22599,N_22873);
and U23439 (N_23439,N_22771,N_22984);
nor U23440 (N_23440,N_22907,N_23052);
or U23441 (N_23441,N_23011,N_22872);
xor U23442 (N_23442,N_22918,N_22665);
nand U23443 (N_23443,N_22917,N_22889);
nor U23444 (N_23444,N_22767,N_22515);
and U23445 (N_23445,N_23068,N_22967);
nand U23446 (N_23446,N_22536,N_22906);
and U23447 (N_23447,N_22935,N_22610);
and U23448 (N_23448,N_23053,N_22866);
nor U23449 (N_23449,N_22778,N_22534);
xor U23450 (N_23450,N_22905,N_23029);
nand U23451 (N_23451,N_23023,N_22828);
and U23452 (N_23452,N_22543,N_22829);
nor U23453 (N_23453,N_22890,N_23085);
nand U23454 (N_23454,N_23118,N_23041);
and U23455 (N_23455,N_22674,N_22949);
and U23456 (N_23456,N_22701,N_22869);
or U23457 (N_23457,N_22578,N_22536);
or U23458 (N_23458,N_23121,N_23124);
nand U23459 (N_23459,N_22561,N_22527);
nor U23460 (N_23460,N_22735,N_22739);
nor U23461 (N_23461,N_22655,N_22628);
or U23462 (N_23462,N_22665,N_23060);
nor U23463 (N_23463,N_22579,N_22636);
or U23464 (N_23464,N_22604,N_22568);
nand U23465 (N_23465,N_22717,N_22772);
or U23466 (N_23466,N_22791,N_22685);
or U23467 (N_23467,N_22878,N_22741);
nor U23468 (N_23468,N_22717,N_22856);
nand U23469 (N_23469,N_22652,N_22566);
nor U23470 (N_23470,N_22609,N_23011);
nor U23471 (N_23471,N_22999,N_23023);
nor U23472 (N_23472,N_23009,N_23046);
nor U23473 (N_23473,N_22940,N_22997);
nor U23474 (N_23474,N_22599,N_22784);
or U23475 (N_23475,N_22505,N_22793);
and U23476 (N_23476,N_22854,N_22625);
and U23477 (N_23477,N_22656,N_22832);
nand U23478 (N_23478,N_22917,N_22726);
nand U23479 (N_23479,N_23028,N_22574);
xor U23480 (N_23480,N_22715,N_22707);
nor U23481 (N_23481,N_22863,N_23046);
nand U23482 (N_23482,N_22851,N_22795);
or U23483 (N_23483,N_22870,N_22720);
nand U23484 (N_23484,N_22770,N_22655);
nor U23485 (N_23485,N_23000,N_22668);
and U23486 (N_23486,N_22871,N_22637);
and U23487 (N_23487,N_23025,N_23042);
and U23488 (N_23488,N_23036,N_22727);
and U23489 (N_23489,N_22557,N_22869);
xor U23490 (N_23490,N_22855,N_23086);
and U23491 (N_23491,N_22519,N_22658);
nand U23492 (N_23492,N_23082,N_22781);
or U23493 (N_23493,N_22906,N_22961);
nor U23494 (N_23494,N_23057,N_22970);
nand U23495 (N_23495,N_22535,N_23000);
nor U23496 (N_23496,N_22623,N_22856);
nand U23497 (N_23497,N_22721,N_22736);
xor U23498 (N_23498,N_22944,N_22764);
nand U23499 (N_23499,N_23094,N_23069);
nor U23500 (N_23500,N_22649,N_22894);
or U23501 (N_23501,N_22974,N_22966);
or U23502 (N_23502,N_22556,N_22633);
nor U23503 (N_23503,N_22903,N_22715);
and U23504 (N_23504,N_22654,N_23067);
nor U23505 (N_23505,N_22967,N_23034);
and U23506 (N_23506,N_23068,N_22806);
nor U23507 (N_23507,N_22678,N_22904);
or U23508 (N_23508,N_22809,N_22626);
nand U23509 (N_23509,N_22626,N_23031);
or U23510 (N_23510,N_22960,N_22885);
and U23511 (N_23511,N_22596,N_22750);
nand U23512 (N_23512,N_22805,N_23043);
nor U23513 (N_23513,N_22676,N_22989);
nand U23514 (N_23514,N_22577,N_22913);
and U23515 (N_23515,N_23091,N_22614);
nand U23516 (N_23516,N_22927,N_23085);
nor U23517 (N_23517,N_22552,N_22955);
and U23518 (N_23518,N_23108,N_23122);
or U23519 (N_23519,N_22568,N_22552);
or U23520 (N_23520,N_23085,N_22724);
or U23521 (N_23521,N_22723,N_22721);
nand U23522 (N_23522,N_23083,N_22796);
and U23523 (N_23523,N_22803,N_22838);
nor U23524 (N_23524,N_22639,N_22908);
nand U23525 (N_23525,N_22849,N_22611);
or U23526 (N_23526,N_23016,N_22776);
and U23527 (N_23527,N_23008,N_22934);
nand U23528 (N_23528,N_22991,N_22714);
nand U23529 (N_23529,N_22830,N_22969);
and U23530 (N_23530,N_22629,N_22928);
nand U23531 (N_23531,N_23027,N_22961);
nand U23532 (N_23532,N_22958,N_22560);
or U23533 (N_23533,N_22885,N_22661);
and U23534 (N_23534,N_22553,N_22961);
xnor U23535 (N_23535,N_22877,N_22888);
and U23536 (N_23536,N_22825,N_22709);
or U23537 (N_23537,N_22854,N_22826);
xnor U23538 (N_23538,N_22723,N_23105);
nand U23539 (N_23539,N_22914,N_22958);
nand U23540 (N_23540,N_22740,N_22972);
nand U23541 (N_23541,N_22819,N_22750);
nand U23542 (N_23542,N_23122,N_22641);
or U23543 (N_23543,N_22917,N_22786);
or U23544 (N_23544,N_22665,N_22951);
or U23545 (N_23545,N_22707,N_22876);
nand U23546 (N_23546,N_22553,N_22903);
or U23547 (N_23547,N_22876,N_22601);
and U23548 (N_23548,N_22693,N_23117);
and U23549 (N_23549,N_22627,N_22553);
and U23550 (N_23550,N_23111,N_23068);
and U23551 (N_23551,N_22757,N_22828);
nand U23552 (N_23552,N_22583,N_22956);
and U23553 (N_23553,N_22652,N_22759);
and U23554 (N_23554,N_22960,N_22770);
or U23555 (N_23555,N_23047,N_22705);
nor U23556 (N_23556,N_22893,N_22520);
nand U23557 (N_23557,N_22539,N_22819);
nor U23558 (N_23558,N_22751,N_22985);
nor U23559 (N_23559,N_22808,N_22524);
and U23560 (N_23560,N_22594,N_22580);
and U23561 (N_23561,N_22582,N_22648);
nand U23562 (N_23562,N_23111,N_23043);
xor U23563 (N_23563,N_22685,N_22876);
nand U23564 (N_23564,N_22950,N_22728);
and U23565 (N_23565,N_22845,N_22743);
xnor U23566 (N_23566,N_22716,N_23013);
and U23567 (N_23567,N_23039,N_22882);
nor U23568 (N_23568,N_23083,N_22788);
nand U23569 (N_23569,N_22878,N_22718);
nor U23570 (N_23570,N_23118,N_22522);
xor U23571 (N_23571,N_23124,N_22839);
and U23572 (N_23572,N_22753,N_22879);
nor U23573 (N_23573,N_22807,N_22572);
and U23574 (N_23574,N_22674,N_22894);
and U23575 (N_23575,N_22711,N_22604);
nor U23576 (N_23576,N_22886,N_22633);
nor U23577 (N_23577,N_22769,N_22679);
or U23578 (N_23578,N_22853,N_22994);
or U23579 (N_23579,N_22517,N_22901);
or U23580 (N_23580,N_22842,N_22741);
xor U23581 (N_23581,N_22704,N_22683);
or U23582 (N_23582,N_22638,N_22818);
and U23583 (N_23583,N_22547,N_22831);
nand U23584 (N_23584,N_23018,N_22962);
xor U23585 (N_23585,N_22758,N_22677);
and U23586 (N_23586,N_22587,N_22509);
xor U23587 (N_23587,N_23044,N_22564);
nor U23588 (N_23588,N_22716,N_23033);
nor U23589 (N_23589,N_22746,N_22622);
and U23590 (N_23590,N_22600,N_22964);
nand U23591 (N_23591,N_22596,N_23050);
xnor U23592 (N_23592,N_23098,N_23052);
and U23593 (N_23593,N_22845,N_23023);
and U23594 (N_23594,N_23115,N_22982);
or U23595 (N_23595,N_22700,N_22588);
nor U23596 (N_23596,N_22625,N_22980);
nand U23597 (N_23597,N_22995,N_22782);
nand U23598 (N_23598,N_22571,N_22811);
nor U23599 (N_23599,N_22568,N_23031);
or U23600 (N_23600,N_22780,N_22898);
nor U23601 (N_23601,N_22761,N_23104);
or U23602 (N_23602,N_22561,N_23064);
or U23603 (N_23603,N_22931,N_23060);
and U23604 (N_23604,N_22872,N_22841);
nand U23605 (N_23605,N_22882,N_22979);
nand U23606 (N_23606,N_22867,N_22993);
or U23607 (N_23607,N_22866,N_22830);
nor U23608 (N_23608,N_22585,N_22540);
nor U23609 (N_23609,N_22598,N_22700);
and U23610 (N_23610,N_22538,N_22924);
nand U23611 (N_23611,N_22625,N_22966);
and U23612 (N_23612,N_23025,N_22843);
or U23613 (N_23613,N_23043,N_23100);
nand U23614 (N_23614,N_22915,N_22508);
nand U23615 (N_23615,N_22537,N_22637);
and U23616 (N_23616,N_22651,N_23113);
xnor U23617 (N_23617,N_23121,N_22937);
or U23618 (N_23618,N_22690,N_22813);
nor U23619 (N_23619,N_22692,N_22830);
and U23620 (N_23620,N_22607,N_23089);
and U23621 (N_23621,N_22939,N_22602);
nor U23622 (N_23622,N_22529,N_22800);
nor U23623 (N_23623,N_22907,N_22578);
nor U23624 (N_23624,N_23108,N_22910);
xor U23625 (N_23625,N_22819,N_22971);
nor U23626 (N_23626,N_22766,N_22696);
xnor U23627 (N_23627,N_23035,N_22706);
nor U23628 (N_23628,N_22779,N_22868);
nand U23629 (N_23629,N_22667,N_22876);
or U23630 (N_23630,N_22866,N_22843);
xor U23631 (N_23631,N_22555,N_23079);
or U23632 (N_23632,N_22991,N_22606);
or U23633 (N_23633,N_22859,N_22654);
xnor U23634 (N_23634,N_22500,N_23026);
or U23635 (N_23635,N_22726,N_23063);
nor U23636 (N_23636,N_22969,N_22873);
or U23637 (N_23637,N_22767,N_22824);
and U23638 (N_23638,N_22788,N_22693);
or U23639 (N_23639,N_22863,N_22754);
xnor U23640 (N_23640,N_22621,N_23067);
nor U23641 (N_23641,N_22503,N_22921);
or U23642 (N_23642,N_23063,N_22670);
nor U23643 (N_23643,N_22617,N_22993);
or U23644 (N_23644,N_22854,N_22700);
nor U23645 (N_23645,N_22532,N_22604);
nor U23646 (N_23646,N_22544,N_22788);
or U23647 (N_23647,N_22728,N_22730);
or U23648 (N_23648,N_22545,N_22743);
nand U23649 (N_23649,N_22598,N_22938);
nand U23650 (N_23650,N_22594,N_22993);
nand U23651 (N_23651,N_22997,N_22535);
or U23652 (N_23652,N_22938,N_23096);
nand U23653 (N_23653,N_22878,N_22775);
nor U23654 (N_23654,N_22910,N_22572);
nand U23655 (N_23655,N_23110,N_23039);
nand U23656 (N_23656,N_22540,N_22600);
nor U23657 (N_23657,N_23070,N_22892);
nand U23658 (N_23658,N_22668,N_22864);
or U23659 (N_23659,N_22961,N_22798);
nand U23660 (N_23660,N_22708,N_22927);
or U23661 (N_23661,N_23079,N_22599);
and U23662 (N_23662,N_23055,N_22745);
nor U23663 (N_23663,N_22962,N_22521);
or U23664 (N_23664,N_22978,N_22517);
nand U23665 (N_23665,N_22952,N_22524);
nor U23666 (N_23666,N_23116,N_22892);
nand U23667 (N_23667,N_23084,N_23018);
nand U23668 (N_23668,N_22847,N_22882);
nor U23669 (N_23669,N_22920,N_23015);
nand U23670 (N_23670,N_22664,N_22953);
nor U23671 (N_23671,N_22987,N_22727);
nor U23672 (N_23672,N_22709,N_23083);
nor U23673 (N_23673,N_23043,N_22923);
nor U23674 (N_23674,N_22723,N_23087);
xor U23675 (N_23675,N_22678,N_22666);
and U23676 (N_23676,N_22537,N_22559);
or U23677 (N_23677,N_22769,N_22719);
nor U23678 (N_23678,N_23011,N_22547);
nor U23679 (N_23679,N_22726,N_22741);
nor U23680 (N_23680,N_22956,N_22860);
nand U23681 (N_23681,N_22589,N_23111);
or U23682 (N_23682,N_22765,N_22946);
or U23683 (N_23683,N_22981,N_22941);
nor U23684 (N_23684,N_23120,N_22931);
or U23685 (N_23685,N_22921,N_23017);
nand U23686 (N_23686,N_22544,N_22611);
nand U23687 (N_23687,N_22668,N_22992);
and U23688 (N_23688,N_23104,N_23111);
nand U23689 (N_23689,N_22551,N_23010);
xor U23690 (N_23690,N_23097,N_23094);
nand U23691 (N_23691,N_22968,N_22791);
and U23692 (N_23692,N_22931,N_22555);
nand U23693 (N_23693,N_22718,N_22793);
nand U23694 (N_23694,N_22778,N_23095);
and U23695 (N_23695,N_22917,N_23017);
nand U23696 (N_23696,N_22741,N_22690);
nor U23697 (N_23697,N_22628,N_23095);
and U23698 (N_23698,N_22610,N_22787);
and U23699 (N_23699,N_22566,N_23114);
and U23700 (N_23700,N_22561,N_23120);
or U23701 (N_23701,N_22509,N_22589);
or U23702 (N_23702,N_22571,N_22970);
nand U23703 (N_23703,N_23065,N_22739);
xnor U23704 (N_23704,N_22867,N_22521);
and U23705 (N_23705,N_23086,N_23115);
nor U23706 (N_23706,N_23124,N_22829);
and U23707 (N_23707,N_22902,N_22748);
xnor U23708 (N_23708,N_23024,N_22586);
and U23709 (N_23709,N_23123,N_22670);
nand U23710 (N_23710,N_22625,N_22853);
or U23711 (N_23711,N_22551,N_22827);
nor U23712 (N_23712,N_23112,N_22598);
xor U23713 (N_23713,N_22677,N_22672);
nand U23714 (N_23714,N_22876,N_22551);
nand U23715 (N_23715,N_22788,N_22570);
xnor U23716 (N_23716,N_22965,N_22505);
nor U23717 (N_23717,N_22819,N_23108);
nand U23718 (N_23718,N_22883,N_22502);
or U23719 (N_23719,N_22839,N_22561);
nor U23720 (N_23720,N_22992,N_22522);
and U23721 (N_23721,N_22711,N_22810);
xnor U23722 (N_23722,N_23018,N_22707);
nand U23723 (N_23723,N_22516,N_23097);
nor U23724 (N_23724,N_22535,N_22766);
or U23725 (N_23725,N_22538,N_22688);
nor U23726 (N_23726,N_23032,N_23044);
or U23727 (N_23727,N_23119,N_22711);
nand U23728 (N_23728,N_23077,N_22729);
xor U23729 (N_23729,N_22814,N_22831);
or U23730 (N_23730,N_22625,N_22539);
nor U23731 (N_23731,N_22608,N_22963);
nand U23732 (N_23732,N_23028,N_23013);
or U23733 (N_23733,N_22889,N_22531);
nor U23734 (N_23734,N_23002,N_22757);
xor U23735 (N_23735,N_22579,N_22891);
nor U23736 (N_23736,N_22578,N_22711);
nand U23737 (N_23737,N_22910,N_22595);
nor U23738 (N_23738,N_22562,N_22568);
and U23739 (N_23739,N_22895,N_22833);
xnor U23740 (N_23740,N_22586,N_22736);
or U23741 (N_23741,N_22870,N_22927);
nor U23742 (N_23742,N_22611,N_23086);
nor U23743 (N_23743,N_22719,N_22833);
nand U23744 (N_23744,N_22553,N_22646);
nor U23745 (N_23745,N_22553,N_22639);
xnor U23746 (N_23746,N_22551,N_22522);
or U23747 (N_23747,N_23121,N_22878);
xor U23748 (N_23748,N_22914,N_22512);
nor U23749 (N_23749,N_22804,N_22673);
and U23750 (N_23750,N_23729,N_23389);
or U23751 (N_23751,N_23524,N_23257);
and U23752 (N_23752,N_23459,N_23648);
nor U23753 (N_23753,N_23720,N_23712);
and U23754 (N_23754,N_23695,N_23657);
nor U23755 (N_23755,N_23614,N_23673);
and U23756 (N_23756,N_23711,N_23302);
and U23757 (N_23757,N_23377,N_23368);
nand U23758 (N_23758,N_23486,N_23195);
nand U23759 (N_23759,N_23227,N_23410);
and U23760 (N_23760,N_23393,N_23228);
and U23761 (N_23761,N_23719,N_23483);
nor U23762 (N_23762,N_23422,N_23613);
and U23763 (N_23763,N_23445,N_23285);
xor U23764 (N_23764,N_23557,N_23206);
nor U23765 (N_23765,N_23588,N_23623);
and U23766 (N_23766,N_23490,N_23456);
nand U23767 (N_23767,N_23622,N_23237);
nand U23768 (N_23768,N_23531,N_23736);
or U23769 (N_23769,N_23662,N_23376);
xor U23770 (N_23770,N_23168,N_23266);
or U23771 (N_23771,N_23273,N_23163);
or U23772 (N_23772,N_23504,N_23357);
nor U23773 (N_23773,N_23731,N_23161);
xor U23774 (N_23774,N_23587,N_23723);
nand U23775 (N_23775,N_23295,N_23217);
and U23776 (N_23776,N_23272,N_23668);
or U23777 (N_23777,N_23496,N_23378);
and U23778 (N_23778,N_23555,N_23604);
nand U23779 (N_23779,N_23724,N_23380);
nor U23780 (N_23780,N_23575,N_23331);
xor U23781 (N_23781,N_23355,N_23324);
nand U23782 (N_23782,N_23564,N_23291);
and U23783 (N_23783,N_23430,N_23586);
nor U23784 (N_23784,N_23129,N_23451);
or U23785 (N_23785,N_23443,N_23289);
nor U23786 (N_23786,N_23427,N_23669);
nor U23787 (N_23787,N_23245,N_23157);
or U23788 (N_23788,N_23678,N_23691);
or U23789 (N_23789,N_23314,N_23322);
nand U23790 (N_23790,N_23585,N_23740);
nand U23791 (N_23791,N_23342,N_23628);
nand U23792 (N_23792,N_23126,N_23374);
or U23793 (N_23793,N_23419,N_23609);
and U23794 (N_23794,N_23714,N_23685);
xnor U23795 (N_23795,N_23280,N_23382);
or U23796 (N_23796,N_23498,N_23592);
or U23797 (N_23797,N_23379,N_23310);
xor U23798 (N_23798,N_23646,N_23385);
or U23799 (N_23799,N_23572,N_23461);
xnor U23800 (N_23800,N_23381,N_23529);
nor U23801 (N_23801,N_23611,N_23674);
and U23802 (N_23802,N_23655,N_23544);
nand U23803 (N_23803,N_23641,N_23661);
nand U23804 (N_23804,N_23260,N_23703);
or U23805 (N_23805,N_23455,N_23696);
and U23806 (N_23806,N_23239,N_23316);
and U23807 (N_23807,N_23642,N_23710);
nand U23808 (N_23808,N_23681,N_23463);
and U23809 (N_23809,N_23677,N_23166);
nor U23810 (N_23810,N_23347,N_23296);
and U23811 (N_23811,N_23580,N_23256);
xnor U23812 (N_23812,N_23560,N_23233);
nor U23813 (N_23813,N_23559,N_23432);
and U23814 (N_23814,N_23503,N_23436);
and U23815 (N_23815,N_23689,N_23699);
and U23816 (N_23816,N_23701,N_23267);
xor U23817 (N_23817,N_23337,N_23251);
nand U23818 (N_23818,N_23537,N_23748);
and U23819 (N_23819,N_23420,N_23246);
and U23820 (N_23820,N_23312,N_23694);
and U23821 (N_23821,N_23183,N_23299);
nand U23822 (N_23822,N_23713,N_23290);
nor U23823 (N_23823,N_23424,N_23511);
xor U23824 (N_23824,N_23154,N_23412);
nand U23825 (N_23825,N_23199,N_23640);
xor U23826 (N_23826,N_23541,N_23474);
nand U23827 (N_23827,N_23632,N_23200);
or U23828 (N_23828,N_23526,N_23261);
nor U23829 (N_23829,N_23244,N_23178);
xnor U23830 (N_23830,N_23247,N_23563);
nor U23831 (N_23831,N_23358,N_23679);
xnor U23832 (N_23832,N_23313,N_23321);
or U23833 (N_23833,N_23666,N_23465);
xor U23834 (N_23834,N_23718,N_23530);
nor U23835 (N_23835,N_23308,N_23513);
xor U23836 (N_23836,N_23220,N_23594);
nor U23837 (N_23837,N_23505,N_23743);
nor U23838 (N_23838,N_23225,N_23721);
nor U23839 (N_23839,N_23131,N_23392);
nand U23840 (N_23840,N_23464,N_23578);
and U23841 (N_23841,N_23545,N_23462);
nand U23842 (N_23842,N_23649,N_23730);
nor U23843 (N_23843,N_23734,N_23143);
or U23844 (N_23844,N_23230,N_23472);
or U23845 (N_23845,N_23287,N_23335);
and U23846 (N_23846,N_23401,N_23521);
nor U23847 (N_23847,N_23600,N_23151);
and U23848 (N_23848,N_23282,N_23134);
or U23849 (N_23849,N_23387,N_23664);
nor U23850 (N_23850,N_23305,N_23350);
nor U23851 (N_23851,N_23692,N_23619);
and U23852 (N_23852,N_23405,N_23468);
xnor U23853 (N_23853,N_23739,N_23400);
or U23854 (N_23854,N_23608,N_23454);
and U23855 (N_23855,N_23727,N_23492);
or U23856 (N_23856,N_23277,N_23449);
nor U23857 (N_23857,N_23232,N_23271);
nand U23858 (N_23858,N_23127,N_23680);
or U23859 (N_23859,N_23255,N_23738);
nand U23860 (N_23860,N_23212,N_23334);
xnor U23861 (N_23861,N_23589,N_23169);
nor U23862 (N_23862,N_23687,N_23698);
nor U23863 (N_23863,N_23582,N_23629);
and U23864 (N_23864,N_23144,N_23571);
nor U23865 (N_23865,N_23403,N_23415);
or U23866 (N_23866,N_23621,N_23136);
nor U23867 (N_23867,N_23643,N_23749);
nand U23868 (N_23868,N_23573,N_23138);
and U23869 (N_23869,N_23439,N_23336);
nand U23870 (N_23870,N_23333,N_23360);
nand U23871 (N_23871,N_23229,N_23323);
nor U23872 (N_23872,N_23515,N_23610);
nor U23873 (N_23873,N_23517,N_23522);
and U23874 (N_23874,N_23583,N_23485);
or U23875 (N_23875,N_23510,N_23605);
nand U23876 (N_23876,N_23325,N_23702);
xor U23877 (N_23877,N_23384,N_23561);
xor U23878 (N_23878,N_23431,N_23684);
nand U23879 (N_23879,N_23181,N_23663);
or U23880 (N_23880,N_23140,N_23269);
nand U23881 (N_23881,N_23265,N_23187);
nor U23882 (N_23882,N_23162,N_23735);
and U23883 (N_23883,N_23448,N_23453);
or U23884 (N_23884,N_23351,N_23519);
nor U23885 (N_23885,N_23469,N_23327);
or U23886 (N_23886,N_23128,N_23471);
and U23887 (N_23887,N_23215,N_23473);
and U23888 (N_23888,N_23328,N_23319);
nor U23889 (N_23889,N_23165,N_23624);
nor U23890 (N_23890,N_23137,N_23356);
and U23891 (N_23891,N_23362,N_23716);
and U23892 (N_23892,N_23341,N_23184);
or U23893 (N_23893,N_23437,N_23425);
or U23894 (N_23894,N_23235,N_23219);
xor U23895 (N_23895,N_23366,N_23398);
nand U23896 (N_23896,N_23388,N_23390);
and U23897 (N_23897,N_23447,N_23656);
and U23898 (N_23898,N_23307,N_23482);
or U23899 (N_23899,N_23155,N_23645);
nand U23900 (N_23900,N_23532,N_23476);
nand U23901 (N_23901,N_23139,N_23250);
or U23902 (N_23902,N_23226,N_23675);
and U23903 (N_23903,N_23213,N_23450);
nand U23904 (N_23904,N_23676,N_23682);
nor U23905 (N_23905,N_23202,N_23315);
or U23906 (N_23906,N_23527,N_23238);
nand U23907 (N_23907,N_23574,N_23533);
and U23908 (N_23908,N_23494,N_23566);
or U23909 (N_23909,N_23596,N_23556);
and U23910 (N_23910,N_23345,N_23276);
nor U23911 (N_23911,N_23705,N_23216);
or U23912 (N_23912,N_23528,N_23491);
nor U23913 (N_23913,N_23547,N_23242);
xor U23914 (N_23914,N_23402,N_23647);
and U23915 (N_23915,N_23683,N_23218);
and U23916 (N_23916,N_23552,N_23297);
or U23917 (N_23917,N_23413,N_23733);
and U23918 (N_23918,N_23177,N_23475);
or U23919 (N_23919,N_23577,N_23383);
nor U23920 (N_23920,N_23330,N_23516);
and U23921 (N_23921,N_23627,N_23214);
xnor U23922 (N_23922,N_23135,N_23576);
and U23923 (N_23923,N_23654,N_23700);
nor U23924 (N_23924,N_23174,N_23644);
and U23925 (N_23925,N_23301,N_23543);
nand U23926 (N_23926,N_23637,N_23525);
nor U23927 (N_23927,N_23708,N_23317);
or U23928 (N_23928,N_23147,N_23466);
and U23929 (N_23929,N_23286,N_23371);
and U23930 (N_23930,N_23599,N_23222);
nand U23931 (N_23931,N_23591,N_23597);
nor U23932 (N_23932,N_23236,N_23241);
and U23933 (N_23933,N_23444,N_23514);
nor U23934 (N_23934,N_23429,N_23565);
nor U23935 (N_23935,N_23534,N_23292);
nor U23936 (N_23936,N_23185,N_23340);
and U23937 (N_23937,N_23421,N_23745);
nor U23938 (N_23938,N_23570,N_23620);
nand U23939 (N_23939,N_23159,N_23553);
and U23940 (N_23940,N_23192,N_23262);
and U23941 (N_23941,N_23369,N_23259);
nor U23942 (N_23942,N_23634,N_23132);
or U23943 (N_23943,N_23567,N_23602);
and U23944 (N_23944,N_23332,N_23279);
xnor U23945 (N_23945,N_23542,N_23326);
nor U23946 (N_23946,N_23359,N_23338);
xor U23947 (N_23947,N_23508,N_23520);
and U23948 (N_23948,N_23441,N_23499);
xnor U23949 (N_23949,N_23497,N_23709);
xnor U23950 (N_23950,N_23460,N_23615);
and U23951 (N_23951,N_23142,N_23467);
nand U23952 (N_23952,N_23258,N_23551);
or U23953 (N_23953,N_23367,N_23593);
or U23954 (N_23954,N_23631,N_23300);
or U23955 (N_23955,N_23651,N_23414);
or U23956 (N_23956,N_23281,N_23211);
nor U23957 (N_23957,N_23728,N_23732);
and U23958 (N_23958,N_23125,N_23480);
or U23959 (N_23959,N_23607,N_23550);
nor U23960 (N_23960,N_23660,N_23523);
and U23961 (N_23961,N_23478,N_23617);
and U23962 (N_23962,N_23416,N_23391);
or U23963 (N_23963,N_23397,N_23606);
and U23964 (N_23964,N_23409,N_23506);
nor U23965 (N_23965,N_23659,N_23579);
and U23966 (N_23966,N_23386,N_23538);
nand U23967 (N_23967,N_23562,N_23288);
and U23968 (N_23968,N_23423,N_23428);
nor U23969 (N_23969,N_23275,N_23725);
or U23970 (N_23970,N_23540,N_23500);
and U23971 (N_23971,N_23318,N_23363);
and U23972 (N_23972,N_23194,N_23417);
nor U23973 (N_23973,N_23370,N_23433);
nor U23974 (N_23974,N_23470,N_23518);
nand U23975 (N_23975,N_23149,N_23343);
xnor U23976 (N_23976,N_23306,N_23512);
or U23977 (N_23977,N_23264,N_23672);
or U23978 (N_23978,N_23688,N_23175);
nand U23979 (N_23979,N_23130,N_23191);
and U23980 (N_23980,N_23435,N_23329);
nand U23981 (N_23981,N_23584,N_23548);
and U23982 (N_23982,N_23186,N_23141);
nand U23983 (N_23983,N_23304,N_23747);
and U23984 (N_23984,N_23243,N_23742);
and U23985 (N_23985,N_23536,N_23442);
or U23986 (N_23986,N_23148,N_23373);
nor U23987 (N_23987,N_23170,N_23179);
nand U23988 (N_23988,N_23457,N_23190);
xnor U23989 (N_23989,N_23481,N_23223);
and U23990 (N_23990,N_23653,N_23221);
nor U23991 (N_23991,N_23156,N_23693);
and U23992 (N_23992,N_23633,N_23590);
nand U23993 (N_23993,N_23352,N_23549);
nor U23994 (N_23994,N_23509,N_23320);
nor U23995 (N_23995,N_23197,N_23690);
and U23996 (N_23996,N_23180,N_23717);
and U23997 (N_23997,N_23133,N_23198);
and U23998 (N_23998,N_23344,N_23395);
nand U23999 (N_23999,N_23210,N_23535);
nor U24000 (N_24000,N_23746,N_23361);
nand U24001 (N_24001,N_23458,N_23204);
or U24002 (N_24002,N_23372,N_23167);
and U24003 (N_24003,N_23152,N_23346);
and U24004 (N_24004,N_23193,N_23704);
nand U24005 (N_24005,N_23440,N_23446);
or U24006 (N_24006,N_23375,N_23626);
and U24007 (N_24007,N_23353,N_23348);
or U24008 (N_24008,N_23635,N_23278);
nor U24009 (N_24009,N_23612,N_23270);
and U24010 (N_24010,N_23150,N_23404);
nand U24011 (N_24011,N_23487,N_23636);
nand U24012 (N_24012,N_23737,N_23434);
and U24013 (N_24013,N_23595,N_23546);
nand U24014 (N_24014,N_23493,N_23309);
nor U24015 (N_24015,N_23618,N_23396);
and U24016 (N_24016,N_23426,N_23207);
or U24017 (N_24017,N_23188,N_23686);
and U24018 (N_24018,N_23502,N_23252);
nor U24019 (N_24019,N_23697,N_23418);
nor U24020 (N_24020,N_23598,N_23158);
nor U24021 (N_24021,N_23298,N_23639);
xor U24022 (N_24022,N_23146,N_23254);
nor U24023 (N_24023,N_23630,N_23452);
nand U24024 (N_24024,N_23715,N_23408);
and U24025 (N_24025,N_23670,N_23164);
and U24026 (N_24026,N_23394,N_23501);
nand U24027 (N_24027,N_23650,N_23365);
or U24028 (N_24028,N_23196,N_23479);
nor U24029 (N_24029,N_23160,N_23311);
and U24030 (N_24030,N_23569,N_23249);
or U24031 (N_24031,N_23581,N_23744);
and U24032 (N_24032,N_23652,N_23407);
nand U24033 (N_24033,N_23707,N_23283);
nor U24034 (N_24034,N_23484,N_23234);
nand U24035 (N_24035,N_23671,N_23201);
nor U24036 (N_24036,N_23601,N_23706);
nor U24037 (N_24037,N_23488,N_23349);
xor U24038 (N_24038,N_23263,N_23658);
and U24039 (N_24039,N_23209,N_23477);
nand U24040 (N_24040,N_23625,N_23176);
and U24041 (N_24041,N_23554,N_23145);
nor U24042 (N_24042,N_23240,N_23171);
nor U24043 (N_24043,N_23294,N_23603);
nand U24044 (N_24044,N_23399,N_23205);
and U24045 (N_24045,N_23568,N_23354);
nand U24046 (N_24046,N_23303,N_23284);
or U24047 (N_24047,N_23665,N_23253);
or U24048 (N_24048,N_23722,N_23268);
and U24049 (N_24049,N_23224,N_23489);
or U24050 (N_24050,N_23189,N_23558);
and U24051 (N_24051,N_23173,N_23203);
nand U24052 (N_24052,N_23406,N_23364);
nand U24053 (N_24053,N_23438,N_23667);
nand U24054 (N_24054,N_23182,N_23495);
nor U24055 (N_24055,N_23616,N_23411);
or U24056 (N_24056,N_23726,N_23231);
and U24057 (N_24057,N_23638,N_23507);
or U24058 (N_24058,N_23248,N_23208);
nor U24059 (N_24059,N_23339,N_23293);
nand U24060 (N_24060,N_23153,N_23172);
and U24061 (N_24061,N_23539,N_23741);
and U24062 (N_24062,N_23274,N_23456);
and U24063 (N_24063,N_23561,N_23357);
or U24064 (N_24064,N_23518,N_23689);
or U24065 (N_24065,N_23456,N_23524);
nor U24066 (N_24066,N_23190,N_23156);
nand U24067 (N_24067,N_23162,N_23629);
xor U24068 (N_24068,N_23275,N_23247);
xor U24069 (N_24069,N_23147,N_23490);
and U24070 (N_24070,N_23454,N_23528);
and U24071 (N_24071,N_23677,N_23334);
nor U24072 (N_24072,N_23246,N_23162);
nand U24073 (N_24073,N_23594,N_23190);
and U24074 (N_24074,N_23372,N_23565);
or U24075 (N_24075,N_23175,N_23206);
nand U24076 (N_24076,N_23587,N_23589);
nor U24077 (N_24077,N_23263,N_23524);
or U24078 (N_24078,N_23644,N_23671);
nand U24079 (N_24079,N_23275,N_23720);
nor U24080 (N_24080,N_23515,N_23228);
and U24081 (N_24081,N_23686,N_23280);
and U24082 (N_24082,N_23265,N_23194);
nand U24083 (N_24083,N_23129,N_23308);
nor U24084 (N_24084,N_23352,N_23305);
and U24085 (N_24085,N_23551,N_23129);
and U24086 (N_24086,N_23220,N_23518);
or U24087 (N_24087,N_23617,N_23225);
and U24088 (N_24088,N_23387,N_23312);
or U24089 (N_24089,N_23725,N_23331);
nor U24090 (N_24090,N_23581,N_23502);
nand U24091 (N_24091,N_23600,N_23657);
or U24092 (N_24092,N_23267,N_23494);
nor U24093 (N_24093,N_23505,N_23617);
and U24094 (N_24094,N_23728,N_23742);
nor U24095 (N_24095,N_23683,N_23210);
and U24096 (N_24096,N_23548,N_23467);
nand U24097 (N_24097,N_23395,N_23744);
nor U24098 (N_24098,N_23447,N_23237);
nor U24099 (N_24099,N_23615,N_23239);
nand U24100 (N_24100,N_23133,N_23646);
nand U24101 (N_24101,N_23454,N_23242);
or U24102 (N_24102,N_23310,N_23502);
nor U24103 (N_24103,N_23401,N_23163);
or U24104 (N_24104,N_23613,N_23410);
or U24105 (N_24105,N_23353,N_23443);
nand U24106 (N_24106,N_23523,N_23177);
nor U24107 (N_24107,N_23430,N_23361);
nor U24108 (N_24108,N_23716,N_23379);
and U24109 (N_24109,N_23566,N_23561);
xnor U24110 (N_24110,N_23257,N_23658);
and U24111 (N_24111,N_23172,N_23588);
and U24112 (N_24112,N_23550,N_23725);
nor U24113 (N_24113,N_23604,N_23295);
and U24114 (N_24114,N_23700,N_23170);
nor U24115 (N_24115,N_23670,N_23649);
nor U24116 (N_24116,N_23180,N_23641);
or U24117 (N_24117,N_23240,N_23323);
and U24118 (N_24118,N_23368,N_23458);
or U24119 (N_24119,N_23255,N_23262);
or U24120 (N_24120,N_23719,N_23556);
nor U24121 (N_24121,N_23591,N_23350);
nor U24122 (N_24122,N_23732,N_23608);
and U24123 (N_24123,N_23232,N_23174);
nor U24124 (N_24124,N_23544,N_23165);
nand U24125 (N_24125,N_23511,N_23690);
or U24126 (N_24126,N_23640,N_23612);
xnor U24127 (N_24127,N_23729,N_23235);
nand U24128 (N_24128,N_23584,N_23254);
nor U24129 (N_24129,N_23333,N_23217);
and U24130 (N_24130,N_23741,N_23649);
or U24131 (N_24131,N_23513,N_23516);
or U24132 (N_24132,N_23371,N_23517);
or U24133 (N_24133,N_23365,N_23453);
and U24134 (N_24134,N_23549,N_23634);
nand U24135 (N_24135,N_23569,N_23314);
nand U24136 (N_24136,N_23176,N_23305);
nor U24137 (N_24137,N_23305,N_23653);
xor U24138 (N_24138,N_23265,N_23744);
nand U24139 (N_24139,N_23421,N_23272);
and U24140 (N_24140,N_23161,N_23133);
nor U24141 (N_24141,N_23299,N_23560);
or U24142 (N_24142,N_23514,N_23195);
nand U24143 (N_24143,N_23318,N_23565);
nand U24144 (N_24144,N_23730,N_23703);
or U24145 (N_24145,N_23371,N_23166);
nor U24146 (N_24146,N_23317,N_23419);
and U24147 (N_24147,N_23248,N_23434);
nor U24148 (N_24148,N_23506,N_23483);
and U24149 (N_24149,N_23308,N_23421);
nor U24150 (N_24150,N_23511,N_23221);
nand U24151 (N_24151,N_23129,N_23266);
and U24152 (N_24152,N_23366,N_23359);
xor U24153 (N_24153,N_23686,N_23602);
and U24154 (N_24154,N_23137,N_23479);
nand U24155 (N_24155,N_23240,N_23387);
nor U24156 (N_24156,N_23661,N_23459);
nor U24157 (N_24157,N_23561,N_23660);
and U24158 (N_24158,N_23151,N_23652);
xnor U24159 (N_24159,N_23649,N_23613);
or U24160 (N_24160,N_23386,N_23293);
nand U24161 (N_24161,N_23439,N_23303);
nor U24162 (N_24162,N_23187,N_23593);
or U24163 (N_24163,N_23528,N_23546);
and U24164 (N_24164,N_23140,N_23134);
nor U24165 (N_24165,N_23341,N_23405);
nor U24166 (N_24166,N_23673,N_23313);
and U24167 (N_24167,N_23473,N_23379);
and U24168 (N_24168,N_23157,N_23458);
nor U24169 (N_24169,N_23584,N_23323);
nand U24170 (N_24170,N_23587,N_23531);
nand U24171 (N_24171,N_23425,N_23248);
and U24172 (N_24172,N_23475,N_23381);
xor U24173 (N_24173,N_23722,N_23523);
nand U24174 (N_24174,N_23516,N_23710);
nand U24175 (N_24175,N_23269,N_23387);
xor U24176 (N_24176,N_23493,N_23566);
nor U24177 (N_24177,N_23206,N_23571);
and U24178 (N_24178,N_23141,N_23565);
nand U24179 (N_24179,N_23265,N_23702);
or U24180 (N_24180,N_23363,N_23428);
nand U24181 (N_24181,N_23351,N_23657);
xor U24182 (N_24182,N_23543,N_23722);
or U24183 (N_24183,N_23569,N_23252);
or U24184 (N_24184,N_23390,N_23664);
nand U24185 (N_24185,N_23206,N_23456);
nor U24186 (N_24186,N_23276,N_23620);
or U24187 (N_24187,N_23549,N_23719);
nand U24188 (N_24188,N_23144,N_23255);
and U24189 (N_24189,N_23586,N_23264);
nor U24190 (N_24190,N_23171,N_23612);
or U24191 (N_24191,N_23646,N_23310);
or U24192 (N_24192,N_23310,N_23153);
and U24193 (N_24193,N_23127,N_23183);
nand U24194 (N_24194,N_23682,N_23353);
and U24195 (N_24195,N_23158,N_23413);
and U24196 (N_24196,N_23540,N_23681);
nor U24197 (N_24197,N_23331,N_23528);
or U24198 (N_24198,N_23161,N_23294);
and U24199 (N_24199,N_23680,N_23156);
or U24200 (N_24200,N_23662,N_23599);
nand U24201 (N_24201,N_23373,N_23382);
nand U24202 (N_24202,N_23150,N_23705);
nand U24203 (N_24203,N_23445,N_23419);
and U24204 (N_24204,N_23665,N_23167);
nand U24205 (N_24205,N_23369,N_23220);
nand U24206 (N_24206,N_23418,N_23684);
and U24207 (N_24207,N_23591,N_23548);
nor U24208 (N_24208,N_23623,N_23332);
nor U24209 (N_24209,N_23367,N_23167);
and U24210 (N_24210,N_23431,N_23478);
and U24211 (N_24211,N_23637,N_23193);
nor U24212 (N_24212,N_23503,N_23376);
or U24213 (N_24213,N_23278,N_23249);
or U24214 (N_24214,N_23240,N_23559);
or U24215 (N_24215,N_23535,N_23616);
nor U24216 (N_24216,N_23592,N_23320);
or U24217 (N_24217,N_23748,N_23562);
or U24218 (N_24218,N_23570,N_23226);
xor U24219 (N_24219,N_23179,N_23428);
or U24220 (N_24220,N_23538,N_23140);
nor U24221 (N_24221,N_23390,N_23201);
nor U24222 (N_24222,N_23423,N_23550);
or U24223 (N_24223,N_23741,N_23406);
xor U24224 (N_24224,N_23504,N_23749);
and U24225 (N_24225,N_23364,N_23427);
nand U24226 (N_24226,N_23134,N_23559);
nor U24227 (N_24227,N_23744,N_23539);
or U24228 (N_24228,N_23377,N_23648);
and U24229 (N_24229,N_23476,N_23602);
nor U24230 (N_24230,N_23358,N_23530);
and U24231 (N_24231,N_23385,N_23205);
nor U24232 (N_24232,N_23593,N_23606);
nand U24233 (N_24233,N_23221,N_23194);
and U24234 (N_24234,N_23550,N_23298);
or U24235 (N_24235,N_23550,N_23575);
nand U24236 (N_24236,N_23361,N_23578);
nor U24237 (N_24237,N_23365,N_23294);
nor U24238 (N_24238,N_23648,N_23249);
nor U24239 (N_24239,N_23408,N_23540);
nor U24240 (N_24240,N_23632,N_23608);
nand U24241 (N_24241,N_23145,N_23174);
and U24242 (N_24242,N_23222,N_23491);
nand U24243 (N_24243,N_23602,N_23233);
nand U24244 (N_24244,N_23523,N_23371);
nand U24245 (N_24245,N_23411,N_23479);
nand U24246 (N_24246,N_23663,N_23471);
nand U24247 (N_24247,N_23606,N_23694);
or U24248 (N_24248,N_23684,N_23621);
nand U24249 (N_24249,N_23210,N_23353);
nand U24250 (N_24250,N_23638,N_23600);
xnor U24251 (N_24251,N_23282,N_23541);
nand U24252 (N_24252,N_23748,N_23380);
and U24253 (N_24253,N_23673,N_23253);
and U24254 (N_24254,N_23716,N_23449);
nor U24255 (N_24255,N_23131,N_23347);
nor U24256 (N_24256,N_23172,N_23711);
xor U24257 (N_24257,N_23598,N_23730);
nand U24258 (N_24258,N_23163,N_23350);
and U24259 (N_24259,N_23674,N_23431);
and U24260 (N_24260,N_23217,N_23239);
nor U24261 (N_24261,N_23713,N_23633);
and U24262 (N_24262,N_23582,N_23419);
nor U24263 (N_24263,N_23695,N_23547);
xnor U24264 (N_24264,N_23728,N_23364);
nor U24265 (N_24265,N_23632,N_23527);
and U24266 (N_24266,N_23150,N_23606);
nor U24267 (N_24267,N_23389,N_23280);
xnor U24268 (N_24268,N_23353,N_23221);
and U24269 (N_24269,N_23312,N_23637);
nor U24270 (N_24270,N_23268,N_23641);
or U24271 (N_24271,N_23420,N_23301);
nor U24272 (N_24272,N_23529,N_23339);
nand U24273 (N_24273,N_23527,N_23573);
or U24274 (N_24274,N_23656,N_23406);
xnor U24275 (N_24275,N_23162,N_23722);
or U24276 (N_24276,N_23353,N_23471);
and U24277 (N_24277,N_23592,N_23643);
nand U24278 (N_24278,N_23252,N_23144);
nand U24279 (N_24279,N_23283,N_23251);
nor U24280 (N_24280,N_23449,N_23296);
or U24281 (N_24281,N_23204,N_23270);
and U24282 (N_24282,N_23250,N_23535);
nor U24283 (N_24283,N_23602,N_23188);
or U24284 (N_24284,N_23495,N_23341);
nor U24285 (N_24285,N_23691,N_23590);
xor U24286 (N_24286,N_23150,N_23294);
nor U24287 (N_24287,N_23168,N_23584);
nand U24288 (N_24288,N_23471,N_23148);
or U24289 (N_24289,N_23437,N_23375);
nor U24290 (N_24290,N_23437,N_23663);
nand U24291 (N_24291,N_23253,N_23682);
nor U24292 (N_24292,N_23465,N_23249);
nand U24293 (N_24293,N_23634,N_23642);
nor U24294 (N_24294,N_23199,N_23739);
and U24295 (N_24295,N_23220,N_23648);
and U24296 (N_24296,N_23573,N_23336);
and U24297 (N_24297,N_23400,N_23157);
nand U24298 (N_24298,N_23465,N_23241);
nand U24299 (N_24299,N_23168,N_23421);
xor U24300 (N_24300,N_23211,N_23260);
nand U24301 (N_24301,N_23574,N_23629);
or U24302 (N_24302,N_23180,N_23358);
nor U24303 (N_24303,N_23261,N_23586);
or U24304 (N_24304,N_23271,N_23222);
nand U24305 (N_24305,N_23271,N_23423);
or U24306 (N_24306,N_23246,N_23497);
and U24307 (N_24307,N_23425,N_23368);
and U24308 (N_24308,N_23510,N_23202);
nor U24309 (N_24309,N_23454,N_23351);
or U24310 (N_24310,N_23307,N_23600);
or U24311 (N_24311,N_23429,N_23685);
xor U24312 (N_24312,N_23327,N_23638);
nor U24313 (N_24313,N_23337,N_23710);
nand U24314 (N_24314,N_23416,N_23173);
xor U24315 (N_24315,N_23469,N_23744);
nand U24316 (N_24316,N_23250,N_23166);
or U24317 (N_24317,N_23648,N_23611);
and U24318 (N_24318,N_23364,N_23318);
or U24319 (N_24319,N_23539,N_23428);
and U24320 (N_24320,N_23735,N_23542);
and U24321 (N_24321,N_23407,N_23217);
or U24322 (N_24322,N_23598,N_23720);
nor U24323 (N_24323,N_23703,N_23588);
and U24324 (N_24324,N_23198,N_23332);
nor U24325 (N_24325,N_23177,N_23300);
nand U24326 (N_24326,N_23720,N_23151);
nor U24327 (N_24327,N_23532,N_23267);
nand U24328 (N_24328,N_23493,N_23316);
nor U24329 (N_24329,N_23214,N_23152);
xor U24330 (N_24330,N_23211,N_23272);
nor U24331 (N_24331,N_23215,N_23644);
nand U24332 (N_24332,N_23603,N_23713);
nor U24333 (N_24333,N_23261,N_23695);
and U24334 (N_24334,N_23220,N_23646);
nand U24335 (N_24335,N_23391,N_23506);
nor U24336 (N_24336,N_23518,N_23332);
nor U24337 (N_24337,N_23374,N_23370);
nand U24338 (N_24338,N_23359,N_23469);
or U24339 (N_24339,N_23407,N_23651);
and U24340 (N_24340,N_23153,N_23688);
nand U24341 (N_24341,N_23623,N_23708);
and U24342 (N_24342,N_23607,N_23715);
nor U24343 (N_24343,N_23504,N_23257);
nor U24344 (N_24344,N_23346,N_23343);
nor U24345 (N_24345,N_23616,N_23297);
and U24346 (N_24346,N_23307,N_23614);
xnor U24347 (N_24347,N_23737,N_23222);
and U24348 (N_24348,N_23435,N_23730);
nor U24349 (N_24349,N_23551,N_23714);
or U24350 (N_24350,N_23161,N_23203);
xnor U24351 (N_24351,N_23194,N_23611);
and U24352 (N_24352,N_23287,N_23666);
nand U24353 (N_24353,N_23419,N_23457);
nor U24354 (N_24354,N_23240,N_23430);
and U24355 (N_24355,N_23185,N_23393);
nor U24356 (N_24356,N_23650,N_23215);
nor U24357 (N_24357,N_23345,N_23425);
and U24358 (N_24358,N_23351,N_23398);
and U24359 (N_24359,N_23650,N_23722);
nand U24360 (N_24360,N_23176,N_23323);
and U24361 (N_24361,N_23139,N_23541);
and U24362 (N_24362,N_23253,N_23177);
nor U24363 (N_24363,N_23412,N_23458);
or U24364 (N_24364,N_23678,N_23570);
nor U24365 (N_24365,N_23275,N_23548);
and U24366 (N_24366,N_23193,N_23272);
nand U24367 (N_24367,N_23600,N_23636);
nand U24368 (N_24368,N_23440,N_23490);
and U24369 (N_24369,N_23589,N_23447);
xor U24370 (N_24370,N_23208,N_23306);
nand U24371 (N_24371,N_23259,N_23686);
or U24372 (N_24372,N_23488,N_23260);
nand U24373 (N_24373,N_23223,N_23663);
nor U24374 (N_24374,N_23526,N_23638);
nor U24375 (N_24375,N_24140,N_24176);
nor U24376 (N_24376,N_24245,N_24304);
and U24377 (N_24377,N_23950,N_24111);
and U24378 (N_24378,N_23822,N_23760);
nor U24379 (N_24379,N_24058,N_24204);
xor U24380 (N_24380,N_24073,N_23866);
and U24381 (N_24381,N_24233,N_23959);
nor U24382 (N_24382,N_23989,N_24185);
nand U24383 (N_24383,N_24187,N_23787);
xor U24384 (N_24384,N_23773,N_23981);
and U24385 (N_24385,N_24170,N_23759);
and U24386 (N_24386,N_23842,N_24227);
nand U24387 (N_24387,N_23938,N_24045);
and U24388 (N_24388,N_24306,N_24283);
and U24389 (N_24389,N_24094,N_23847);
and U24390 (N_24390,N_23881,N_23836);
and U24391 (N_24391,N_23808,N_23967);
nor U24392 (N_24392,N_23924,N_24365);
and U24393 (N_24393,N_24166,N_24067);
nand U24394 (N_24394,N_23770,N_24355);
and U24395 (N_24395,N_24028,N_23761);
xor U24396 (N_24396,N_24345,N_24263);
xor U24397 (N_24397,N_23794,N_24279);
nor U24398 (N_24398,N_24211,N_24226);
and U24399 (N_24399,N_24196,N_24148);
nand U24400 (N_24400,N_24260,N_23915);
or U24401 (N_24401,N_24017,N_23806);
or U24402 (N_24402,N_24186,N_24206);
or U24403 (N_24403,N_24179,N_24139);
or U24404 (N_24404,N_24291,N_23828);
nand U24405 (N_24405,N_24331,N_24029);
and U24406 (N_24406,N_24228,N_23751);
nand U24407 (N_24407,N_24343,N_23974);
or U24408 (N_24408,N_23945,N_24302);
nand U24409 (N_24409,N_24298,N_23800);
xor U24410 (N_24410,N_24025,N_23810);
xnor U24411 (N_24411,N_24205,N_24201);
and U24412 (N_24412,N_24070,N_24059);
nor U24413 (N_24413,N_23921,N_24071);
nor U24414 (N_24414,N_24044,N_23965);
xor U24415 (N_24415,N_24224,N_24155);
nand U24416 (N_24416,N_24225,N_24002);
and U24417 (N_24417,N_24040,N_23801);
xor U24418 (N_24418,N_24316,N_23750);
nand U24419 (N_24419,N_24216,N_23803);
nand U24420 (N_24420,N_23902,N_24190);
or U24421 (N_24421,N_23823,N_23785);
nor U24422 (N_24422,N_24213,N_24270);
nand U24423 (N_24423,N_23900,N_23953);
and U24424 (N_24424,N_24237,N_24021);
or U24425 (N_24425,N_24266,N_23934);
nor U24426 (N_24426,N_24099,N_23976);
nor U24427 (N_24427,N_23825,N_23908);
or U24428 (N_24428,N_24314,N_24280);
or U24429 (N_24429,N_24235,N_24009);
nor U24430 (N_24430,N_24092,N_23771);
nand U24431 (N_24431,N_23817,N_24246);
or U24432 (N_24432,N_24181,N_24035);
and U24433 (N_24433,N_23916,N_24311);
nand U24434 (N_24434,N_24320,N_24004);
nor U24435 (N_24435,N_24130,N_23867);
and U24436 (N_24436,N_24103,N_23997);
nor U24437 (N_24437,N_24284,N_24313);
nor U24438 (N_24438,N_23789,N_24281);
or U24439 (N_24439,N_24164,N_24356);
nand U24440 (N_24440,N_23978,N_23892);
nand U24441 (N_24441,N_23756,N_23765);
nand U24442 (N_24442,N_23766,N_24084);
nor U24443 (N_24443,N_24309,N_24091);
nand U24444 (N_24444,N_24156,N_24317);
or U24445 (N_24445,N_23906,N_23821);
and U24446 (N_24446,N_24057,N_24119);
nor U24447 (N_24447,N_24022,N_24341);
nand U24448 (N_24448,N_23988,N_24020);
and U24449 (N_24449,N_24325,N_23877);
or U24450 (N_24450,N_24294,N_24238);
xor U24451 (N_24451,N_23849,N_24049);
nand U24452 (N_24452,N_24348,N_24026);
and U24453 (N_24453,N_24212,N_24367);
and U24454 (N_24454,N_24121,N_24330);
nand U24455 (N_24455,N_24300,N_24167);
and U24456 (N_24456,N_23772,N_23947);
xor U24457 (N_24457,N_24077,N_24189);
and U24458 (N_24458,N_24333,N_24267);
or U24459 (N_24459,N_24122,N_24096);
and U24460 (N_24460,N_23853,N_23949);
xor U24461 (N_24461,N_23896,N_24141);
nand U24462 (N_24462,N_24042,N_24310);
nor U24463 (N_24463,N_24328,N_24039);
xnor U24464 (N_24464,N_24287,N_24292);
nand U24465 (N_24465,N_24242,N_24015);
or U24466 (N_24466,N_23986,N_23863);
nand U24467 (N_24467,N_23954,N_24098);
nor U24468 (N_24468,N_24289,N_23793);
and U24469 (N_24469,N_24043,N_23777);
nor U24470 (N_24470,N_24162,N_24048);
nor U24471 (N_24471,N_24363,N_23873);
and U24472 (N_24472,N_24210,N_24274);
or U24473 (N_24473,N_23832,N_23929);
nand U24474 (N_24474,N_24172,N_24258);
and U24475 (N_24475,N_24334,N_24082);
nor U24476 (N_24476,N_24244,N_24090);
xnor U24477 (N_24477,N_23980,N_23797);
nor U24478 (N_24478,N_24193,N_23975);
nand U24479 (N_24479,N_24299,N_24230);
and U24480 (N_24480,N_24150,N_23861);
or U24481 (N_24481,N_23907,N_23802);
or U24482 (N_24482,N_23848,N_23805);
nor U24483 (N_24483,N_24038,N_24036);
and U24484 (N_24484,N_24138,N_23911);
nand U24485 (N_24485,N_23844,N_24135);
or U24486 (N_24486,N_24159,N_23790);
xor U24487 (N_24487,N_24322,N_23811);
nor U24488 (N_24488,N_24307,N_24072);
and U24489 (N_24489,N_24034,N_24183);
nor U24490 (N_24490,N_23833,N_24372);
nor U24491 (N_24491,N_24056,N_24006);
or U24492 (N_24492,N_24282,N_24231);
xnor U24493 (N_24493,N_24342,N_23996);
or U24494 (N_24494,N_23851,N_24197);
or U24495 (N_24495,N_24194,N_23786);
and U24496 (N_24496,N_24218,N_24066);
or U24497 (N_24497,N_24276,N_24312);
xnor U24498 (N_24498,N_24163,N_24340);
or U24499 (N_24499,N_23884,N_24188);
or U24500 (N_24500,N_23969,N_24338);
xnor U24501 (N_24501,N_23871,N_24359);
nand U24502 (N_24502,N_24327,N_24217);
nor U24503 (N_24503,N_23767,N_23769);
or U24504 (N_24504,N_23942,N_24142);
and U24505 (N_24505,N_24182,N_24200);
or U24506 (N_24506,N_24125,N_23925);
or U24507 (N_24507,N_23857,N_24132);
nor U24508 (N_24508,N_24123,N_24000);
nor U24509 (N_24509,N_24364,N_24089);
nand U24510 (N_24510,N_24250,N_24199);
nand U24511 (N_24511,N_24080,N_23961);
and U24512 (N_24512,N_23809,N_23798);
xnor U24513 (N_24513,N_23788,N_24368);
or U24514 (N_24514,N_24052,N_24168);
nand U24515 (N_24515,N_24151,N_24175);
and U24516 (N_24516,N_23876,N_23846);
or U24517 (N_24517,N_24074,N_23839);
or U24518 (N_24518,N_24027,N_24318);
and U24519 (N_24519,N_24290,N_23917);
nor U24520 (N_24520,N_23973,N_24223);
xnor U24521 (N_24521,N_24243,N_23984);
nor U24522 (N_24522,N_24319,N_24102);
xnor U24523 (N_24523,N_23928,N_24335);
nor U24524 (N_24524,N_24208,N_23992);
nand U24525 (N_24525,N_24014,N_23991);
nand U24526 (N_24526,N_24350,N_24303);
nor U24527 (N_24527,N_24301,N_23885);
or U24528 (N_24528,N_24326,N_24088);
nand U24529 (N_24529,N_24234,N_24174);
and U24530 (N_24530,N_23913,N_23904);
or U24531 (N_24531,N_24296,N_24055);
nand U24532 (N_24532,N_23918,N_23887);
or U24533 (N_24533,N_23827,N_23762);
xor U24534 (N_24534,N_23837,N_24161);
xor U24535 (N_24535,N_23998,N_24005);
nand U24536 (N_24536,N_24269,N_23854);
nand U24537 (N_24537,N_23764,N_24352);
nand U24538 (N_24538,N_23752,N_24347);
and U24539 (N_24539,N_24249,N_24154);
nor U24540 (N_24540,N_24128,N_24112);
or U24541 (N_24541,N_24337,N_24129);
xor U24542 (N_24542,N_24202,N_24146);
and U24543 (N_24543,N_23905,N_24143);
and U24544 (N_24544,N_24024,N_24262);
nor U24545 (N_24545,N_24371,N_23952);
nand U24546 (N_24546,N_24149,N_24297);
and U24547 (N_24547,N_23999,N_23994);
nor U24548 (N_24548,N_23880,N_23964);
and U24549 (N_24549,N_24346,N_24033);
or U24550 (N_24550,N_24054,N_23971);
nand U24551 (N_24551,N_24209,N_24195);
xor U24552 (N_24552,N_24252,N_23920);
or U24553 (N_24553,N_23946,N_23774);
and U24554 (N_24554,N_23966,N_23859);
nor U24555 (N_24555,N_23910,N_23956);
or U24556 (N_24556,N_23845,N_23977);
nand U24557 (N_24557,N_24256,N_23869);
nor U24558 (N_24558,N_24013,N_24308);
or U24559 (N_24559,N_24083,N_24214);
nand U24560 (N_24560,N_23931,N_23912);
and U24561 (N_24561,N_23815,N_24255);
or U24562 (N_24562,N_24241,N_24113);
nor U24563 (N_24563,N_23835,N_24007);
or U24564 (N_24564,N_23933,N_24011);
and U24565 (N_24565,N_24360,N_24062);
and U24566 (N_24566,N_23784,N_24321);
and U24567 (N_24567,N_24012,N_24171);
and U24568 (N_24568,N_24023,N_23865);
nor U24569 (N_24569,N_24215,N_24265);
xor U24570 (N_24570,N_23882,N_23855);
xor U24571 (N_24571,N_24061,N_23799);
and U24572 (N_24572,N_23757,N_23922);
or U24573 (N_24573,N_24133,N_24239);
nor U24574 (N_24574,N_24184,N_24259);
and U24575 (N_24575,N_24107,N_23963);
xnor U24576 (N_24576,N_23957,N_24085);
or U24577 (N_24577,N_24104,N_23955);
xor U24578 (N_24578,N_23990,N_24169);
nor U24579 (N_24579,N_23914,N_24374);
nor U24580 (N_24580,N_23982,N_24093);
and U24581 (N_24581,N_24158,N_23783);
nor U24582 (N_24582,N_24079,N_23893);
nor U24583 (N_24583,N_23778,N_24081);
and U24584 (N_24584,N_23795,N_24087);
nand U24585 (N_24585,N_24229,N_24323);
and U24586 (N_24586,N_24019,N_24064);
or U24587 (N_24587,N_23923,N_24068);
or U24588 (N_24588,N_24293,N_23886);
and U24589 (N_24589,N_23943,N_23872);
or U24590 (N_24590,N_24351,N_23824);
xnor U24591 (N_24591,N_24016,N_24145);
nor U24592 (N_24592,N_23754,N_24086);
nor U24593 (N_24593,N_24353,N_24105);
nor U24594 (N_24594,N_24286,N_24253);
and U24595 (N_24595,N_23895,N_24124);
nand U24596 (N_24596,N_24100,N_24277);
nor U24597 (N_24597,N_24192,N_23883);
nor U24598 (N_24598,N_24152,N_23983);
and U24599 (N_24599,N_23962,N_24203);
nand U24600 (N_24600,N_23753,N_23776);
nand U24601 (N_24601,N_23834,N_24221);
nor U24602 (N_24602,N_24339,N_23820);
nor U24603 (N_24603,N_24050,N_23940);
xor U24604 (N_24604,N_24329,N_24136);
nor U24605 (N_24605,N_24065,N_23979);
and U24606 (N_24606,N_23819,N_23935);
xor U24607 (N_24607,N_23782,N_23843);
nor U24608 (N_24608,N_24106,N_24248);
and U24609 (N_24609,N_24010,N_23941);
nor U24610 (N_24610,N_23894,N_23960);
or U24611 (N_24611,N_24373,N_24078);
and U24612 (N_24612,N_23791,N_24305);
xnor U24613 (N_24613,N_24268,N_23856);
nand U24614 (N_24614,N_24285,N_23829);
nand U24615 (N_24615,N_24332,N_23987);
or U24616 (N_24616,N_23891,N_24295);
nand U24617 (N_24617,N_24220,N_24247);
or U24618 (N_24618,N_24261,N_24236);
nand U24619 (N_24619,N_24003,N_24041);
nand U24620 (N_24620,N_24095,N_24037);
xnor U24621 (N_24621,N_23875,N_24366);
and U24622 (N_24622,N_24254,N_23796);
nor U24623 (N_24623,N_24354,N_23930);
xnor U24624 (N_24624,N_23879,N_24147);
nand U24625 (N_24625,N_24069,N_23972);
nor U24626 (N_24626,N_24097,N_24051);
or U24627 (N_24627,N_23852,N_24173);
nand U24628 (N_24628,N_23927,N_23890);
nor U24629 (N_24629,N_24063,N_23958);
and U24630 (N_24630,N_23758,N_24018);
xor U24631 (N_24631,N_23951,N_23899);
and U24632 (N_24632,N_23903,N_23818);
nand U24633 (N_24633,N_24032,N_23944);
or U24634 (N_24634,N_24358,N_24153);
and U24635 (N_24635,N_23985,N_23860);
nand U24636 (N_24636,N_23813,N_23840);
xor U24637 (N_24637,N_24137,N_23936);
xor U24638 (N_24638,N_24116,N_24120);
or U24639 (N_24639,N_23868,N_24198);
nand U24640 (N_24640,N_24349,N_24180);
nand U24641 (N_24641,N_23838,N_23864);
nand U24642 (N_24642,N_24075,N_24232);
nand U24643 (N_24643,N_24031,N_24060);
or U24644 (N_24644,N_23812,N_24369);
nand U24645 (N_24645,N_24001,N_24324);
nor U24646 (N_24646,N_23780,N_23932);
nand U24647 (N_24647,N_23897,N_24117);
or U24648 (N_24648,N_24165,N_24046);
and U24649 (N_24649,N_24178,N_24144);
and U24650 (N_24650,N_24177,N_24101);
nor U24651 (N_24651,N_24110,N_23826);
or U24652 (N_24652,N_23878,N_24127);
or U24653 (N_24653,N_24362,N_24222);
or U24654 (N_24654,N_24315,N_23755);
nor U24655 (N_24655,N_24361,N_24126);
and U24656 (N_24656,N_23858,N_24219);
xnor U24657 (N_24657,N_23763,N_24288);
nor U24658 (N_24658,N_23804,N_24264);
and U24659 (N_24659,N_24114,N_23816);
and U24660 (N_24660,N_23909,N_23995);
nand U24661 (N_24661,N_24109,N_24257);
and U24662 (N_24662,N_24240,N_24344);
nand U24663 (N_24663,N_23874,N_23768);
and U24664 (N_24664,N_23862,N_23939);
nor U24665 (N_24665,N_24275,N_24115);
xor U24666 (N_24666,N_23814,N_24336);
and U24667 (N_24667,N_23901,N_24273);
or U24668 (N_24668,N_24118,N_23919);
or U24669 (N_24669,N_23937,N_24278);
xor U24670 (N_24670,N_23926,N_23831);
and U24671 (N_24671,N_24008,N_24134);
or U24672 (N_24672,N_24370,N_23968);
or U24673 (N_24673,N_23775,N_24191);
or U24674 (N_24674,N_23970,N_23781);
nand U24675 (N_24675,N_24076,N_23792);
and U24676 (N_24676,N_24157,N_24160);
nand U24677 (N_24677,N_23830,N_23850);
nor U24678 (N_24678,N_23870,N_23889);
nor U24679 (N_24679,N_23948,N_23993);
nor U24680 (N_24680,N_23841,N_24357);
nor U24681 (N_24681,N_24030,N_23888);
and U24682 (N_24682,N_23807,N_24251);
or U24683 (N_24683,N_24272,N_23898);
nand U24684 (N_24684,N_23779,N_24047);
or U24685 (N_24685,N_24108,N_24131);
nor U24686 (N_24686,N_24207,N_24053);
nand U24687 (N_24687,N_24271,N_23852);
nor U24688 (N_24688,N_23990,N_23838);
and U24689 (N_24689,N_24112,N_23977);
or U24690 (N_24690,N_24233,N_24130);
nand U24691 (N_24691,N_24063,N_24259);
or U24692 (N_24692,N_23893,N_24278);
nand U24693 (N_24693,N_24113,N_24258);
and U24694 (N_24694,N_23967,N_24362);
nand U24695 (N_24695,N_23760,N_24057);
and U24696 (N_24696,N_24092,N_23998);
nand U24697 (N_24697,N_24017,N_24243);
and U24698 (N_24698,N_24248,N_24063);
or U24699 (N_24699,N_24282,N_24004);
nand U24700 (N_24700,N_24344,N_24260);
and U24701 (N_24701,N_24098,N_23920);
or U24702 (N_24702,N_23934,N_23913);
nor U24703 (N_24703,N_23847,N_24294);
or U24704 (N_24704,N_24032,N_23996);
nor U24705 (N_24705,N_23820,N_24360);
and U24706 (N_24706,N_23860,N_24239);
nor U24707 (N_24707,N_23886,N_24075);
nand U24708 (N_24708,N_24207,N_24221);
nand U24709 (N_24709,N_24311,N_23995);
or U24710 (N_24710,N_24310,N_23979);
nor U24711 (N_24711,N_24310,N_23977);
xor U24712 (N_24712,N_23830,N_24336);
nor U24713 (N_24713,N_24151,N_24122);
nor U24714 (N_24714,N_23785,N_24016);
and U24715 (N_24715,N_24122,N_24068);
xnor U24716 (N_24716,N_23783,N_24230);
and U24717 (N_24717,N_24349,N_24279);
xor U24718 (N_24718,N_24209,N_24361);
and U24719 (N_24719,N_24253,N_24365);
or U24720 (N_24720,N_24050,N_23788);
or U24721 (N_24721,N_24195,N_23844);
nand U24722 (N_24722,N_24248,N_23901);
and U24723 (N_24723,N_23837,N_23970);
nor U24724 (N_24724,N_24301,N_24337);
nor U24725 (N_24725,N_24160,N_24203);
or U24726 (N_24726,N_24234,N_24322);
nor U24727 (N_24727,N_24282,N_24016);
nor U24728 (N_24728,N_24045,N_24309);
and U24729 (N_24729,N_23876,N_23918);
nand U24730 (N_24730,N_23776,N_23997);
and U24731 (N_24731,N_24069,N_23815);
nand U24732 (N_24732,N_23855,N_23926);
or U24733 (N_24733,N_23957,N_23999);
and U24734 (N_24734,N_24017,N_24199);
or U24735 (N_24735,N_24112,N_24329);
nand U24736 (N_24736,N_23874,N_23986);
or U24737 (N_24737,N_24028,N_24336);
or U24738 (N_24738,N_24292,N_24223);
xnor U24739 (N_24739,N_23917,N_23861);
nand U24740 (N_24740,N_23832,N_23890);
or U24741 (N_24741,N_23952,N_24284);
nand U24742 (N_24742,N_24367,N_24022);
nand U24743 (N_24743,N_23959,N_24226);
and U24744 (N_24744,N_24294,N_23803);
nand U24745 (N_24745,N_23930,N_23968);
xnor U24746 (N_24746,N_24105,N_24296);
and U24747 (N_24747,N_23960,N_23846);
or U24748 (N_24748,N_24034,N_23971);
xnor U24749 (N_24749,N_23793,N_24259);
or U24750 (N_24750,N_24147,N_24094);
nor U24751 (N_24751,N_23908,N_24242);
or U24752 (N_24752,N_23928,N_24153);
nand U24753 (N_24753,N_24278,N_24131);
nor U24754 (N_24754,N_23995,N_24224);
or U24755 (N_24755,N_24026,N_24241);
and U24756 (N_24756,N_23825,N_23826);
xor U24757 (N_24757,N_24013,N_24139);
and U24758 (N_24758,N_24102,N_24217);
and U24759 (N_24759,N_24234,N_24286);
and U24760 (N_24760,N_24361,N_23752);
nand U24761 (N_24761,N_24046,N_23931);
nand U24762 (N_24762,N_23835,N_24212);
or U24763 (N_24763,N_23995,N_24278);
xor U24764 (N_24764,N_23885,N_23917);
or U24765 (N_24765,N_24036,N_24292);
nand U24766 (N_24766,N_23773,N_23977);
or U24767 (N_24767,N_23865,N_23944);
nand U24768 (N_24768,N_24244,N_23802);
or U24769 (N_24769,N_23876,N_24124);
nor U24770 (N_24770,N_23877,N_24033);
or U24771 (N_24771,N_24353,N_24230);
xnor U24772 (N_24772,N_23775,N_24281);
nand U24773 (N_24773,N_24001,N_24177);
xor U24774 (N_24774,N_23951,N_23815);
nand U24775 (N_24775,N_23951,N_23860);
nand U24776 (N_24776,N_24045,N_23964);
or U24777 (N_24777,N_23778,N_24199);
nand U24778 (N_24778,N_24106,N_23981);
or U24779 (N_24779,N_24287,N_24091);
nor U24780 (N_24780,N_23966,N_24006);
nor U24781 (N_24781,N_24235,N_24316);
or U24782 (N_24782,N_23879,N_24324);
nor U24783 (N_24783,N_24075,N_23966);
nand U24784 (N_24784,N_23921,N_24257);
and U24785 (N_24785,N_24154,N_24096);
nand U24786 (N_24786,N_24080,N_24291);
or U24787 (N_24787,N_24316,N_24347);
nand U24788 (N_24788,N_24080,N_23927);
nand U24789 (N_24789,N_24020,N_24010);
and U24790 (N_24790,N_23933,N_23857);
and U24791 (N_24791,N_24301,N_23968);
nand U24792 (N_24792,N_23998,N_24199);
nor U24793 (N_24793,N_24094,N_24313);
nor U24794 (N_24794,N_24274,N_24294);
nor U24795 (N_24795,N_24128,N_24037);
and U24796 (N_24796,N_24118,N_23964);
nand U24797 (N_24797,N_23837,N_23897);
nor U24798 (N_24798,N_23873,N_24216);
nor U24799 (N_24799,N_24075,N_23811);
nor U24800 (N_24800,N_23980,N_23875);
xor U24801 (N_24801,N_23814,N_24357);
and U24802 (N_24802,N_24032,N_24121);
or U24803 (N_24803,N_24355,N_24208);
nor U24804 (N_24804,N_23899,N_23919);
or U24805 (N_24805,N_24081,N_23798);
and U24806 (N_24806,N_24315,N_23814);
and U24807 (N_24807,N_24364,N_23951);
nor U24808 (N_24808,N_24177,N_24231);
or U24809 (N_24809,N_23926,N_23834);
xnor U24810 (N_24810,N_23959,N_24244);
nor U24811 (N_24811,N_24296,N_23781);
nor U24812 (N_24812,N_24288,N_24285);
and U24813 (N_24813,N_24157,N_23815);
and U24814 (N_24814,N_24259,N_23778);
or U24815 (N_24815,N_23797,N_24134);
and U24816 (N_24816,N_23780,N_23946);
and U24817 (N_24817,N_24252,N_23832);
or U24818 (N_24818,N_24332,N_23805);
nand U24819 (N_24819,N_23986,N_24220);
or U24820 (N_24820,N_23760,N_24338);
nor U24821 (N_24821,N_23946,N_24137);
or U24822 (N_24822,N_24330,N_24004);
xnor U24823 (N_24823,N_24337,N_23826);
and U24824 (N_24824,N_23974,N_24319);
nand U24825 (N_24825,N_23793,N_24303);
or U24826 (N_24826,N_24099,N_24171);
nor U24827 (N_24827,N_23984,N_24072);
nand U24828 (N_24828,N_24343,N_23764);
nand U24829 (N_24829,N_23917,N_23768);
nor U24830 (N_24830,N_23891,N_24122);
and U24831 (N_24831,N_23885,N_24116);
or U24832 (N_24832,N_24245,N_24268);
or U24833 (N_24833,N_24372,N_23794);
nor U24834 (N_24834,N_23981,N_23759);
nand U24835 (N_24835,N_24008,N_23971);
or U24836 (N_24836,N_23874,N_24310);
nand U24837 (N_24837,N_24114,N_23984);
nor U24838 (N_24838,N_24146,N_24256);
nor U24839 (N_24839,N_24313,N_23779);
or U24840 (N_24840,N_24051,N_24281);
nor U24841 (N_24841,N_24241,N_24183);
or U24842 (N_24842,N_24337,N_24239);
xnor U24843 (N_24843,N_23764,N_24359);
xnor U24844 (N_24844,N_23964,N_24008);
or U24845 (N_24845,N_24353,N_23785);
or U24846 (N_24846,N_24004,N_24254);
or U24847 (N_24847,N_24086,N_23851);
nor U24848 (N_24848,N_24027,N_24283);
nor U24849 (N_24849,N_24344,N_24229);
and U24850 (N_24850,N_24250,N_24081);
and U24851 (N_24851,N_24176,N_24193);
or U24852 (N_24852,N_24045,N_24084);
nor U24853 (N_24853,N_24006,N_23865);
nor U24854 (N_24854,N_24269,N_24178);
and U24855 (N_24855,N_24298,N_24145);
xor U24856 (N_24856,N_23892,N_24167);
xnor U24857 (N_24857,N_24116,N_24074);
and U24858 (N_24858,N_23777,N_24214);
nand U24859 (N_24859,N_24172,N_24311);
xnor U24860 (N_24860,N_24265,N_23951);
and U24861 (N_24861,N_24113,N_24244);
nor U24862 (N_24862,N_24289,N_23907);
nand U24863 (N_24863,N_24080,N_23997);
or U24864 (N_24864,N_23946,N_24261);
or U24865 (N_24865,N_24071,N_24297);
and U24866 (N_24866,N_24014,N_24263);
and U24867 (N_24867,N_23789,N_23907);
nor U24868 (N_24868,N_24365,N_24083);
and U24869 (N_24869,N_24165,N_24299);
or U24870 (N_24870,N_24309,N_24207);
and U24871 (N_24871,N_24332,N_24056);
or U24872 (N_24872,N_23909,N_23760);
or U24873 (N_24873,N_24085,N_24074);
or U24874 (N_24874,N_24321,N_23941);
nor U24875 (N_24875,N_24330,N_24293);
nor U24876 (N_24876,N_24032,N_24176);
and U24877 (N_24877,N_23959,N_24107);
and U24878 (N_24878,N_23826,N_23764);
or U24879 (N_24879,N_24011,N_24013);
nor U24880 (N_24880,N_24062,N_24008);
and U24881 (N_24881,N_23804,N_23929);
xnor U24882 (N_24882,N_23911,N_24215);
nor U24883 (N_24883,N_23914,N_24276);
nor U24884 (N_24884,N_23887,N_24313);
or U24885 (N_24885,N_24314,N_23777);
nand U24886 (N_24886,N_24040,N_24260);
or U24887 (N_24887,N_23800,N_24075);
or U24888 (N_24888,N_24254,N_23931);
nor U24889 (N_24889,N_24191,N_24105);
and U24890 (N_24890,N_24246,N_23850);
or U24891 (N_24891,N_23824,N_24247);
and U24892 (N_24892,N_24036,N_23828);
nor U24893 (N_24893,N_23816,N_24298);
xor U24894 (N_24894,N_23953,N_24054);
and U24895 (N_24895,N_23979,N_24326);
nand U24896 (N_24896,N_23988,N_23996);
and U24897 (N_24897,N_24269,N_24249);
xor U24898 (N_24898,N_24110,N_24273);
and U24899 (N_24899,N_23955,N_23918);
nand U24900 (N_24900,N_23868,N_23998);
or U24901 (N_24901,N_23977,N_24279);
nor U24902 (N_24902,N_23885,N_23976);
nor U24903 (N_24903,N_24256,N_23899);
nand U24904 (N_24904,N_24254,N_23911);
and U24905 (N_24905,N_23915,N_23990);
nor U24906 (N_24906,N_23822,N_24332);
nor U24907 (N_24907,N_24291,N_23850);
nand U24908 (N_24908,N_24357,N_23946);
or U24909 (N_24909,N_24170,N_23944);
nor U24910 (N_24910,N_24260,N_24113);
nor U24911 (N_24911,N_24099,N_23860);
or U24912 (N_24912,N_23911,N_24213);
or U24913 (N_24913,N_24307,N_24027);
nand U24914 (N_24914,N_24078,N_24013);
and U24915 (N_24915,N_24006,N_24244);
nand U24916 (N_24916,N_24034,N_24366);
nor U24917 (N_24917,N_24218,N_23774);
and U24918 (N_24918,N_23979,N_23954);
or U24919 (N_24919,N_24149,N_24052);
nor U24920 (N_24920,N_24140,N_23931);
or U24921 (N_24921,N_24112,N_23978);
or U24922 (N_24922,N_24064,N_23833);
xnor U24923 (N_24923,N_24362,N_24204);
and U24924 (N_24924,N_24196,N_24149);
xnor U24925 (N_24925,N_24373,N_23826);
or U24926 (N_24926,N_23767,N_24368);
nand U24927 (N_24927,N_24005,N_23783);
or U24928 (N_24928,N_24182,N_23982);
or U24929 (N_24929,N_24151,N_24283);
xnor U24930 (N_24930,N_24227,N_24065);
nand U24931 (N_24931,N_24151,N_23975);
or U24932 (N_24932,N_24149,N_23794);
xor U24933 (N_24933,N_24268,N_24210);
xor U24934 (N_24934,N_24236,N_24212);
and U24935 (N_24935,N_24221,N_24339);
and U24936 (N_24936,N_24037,N_23802);
or U24937 (N_24937,N_23983,N_24143);
or U24938 (N_24938,N_23824,N_23840);
nand U24939 (N_24939,N_24282,N_24095);
nor U24940 (N_24940,N_24015,N_24143);
nor U24941 (N_24941,N_24152,N_24330);
nor U24942 (N_24942,N_24184,N_24143);
nand U24943 (N_24943,N_23823,N_23764);
nand U24944 (N_24944,N_23784,N_23937);
or U24945 (N_24945,N_24007,N_24373);
nor U24946 (N_24946,N_24373,N_24228);
or U24947 (N_24947,N_24263,N_24255);
or U24948 (N_24948,N_24275,N_23795);
nor U24949 (N_24949,N_23826,N_24205);
nor U24950 (N_24950,N_23949,N_24274);
nor U24951 (N_24951,N_24051,N_23956);
and U24952 (N_24952,N_24022,N_24126);
or U24953 (N_24953,N_24288,N_24342);
or U24954 (N_24954,N_24219,N_23784);
xor U24955 (N_24955,N_24267,N_24215);
nor U24956 (N_24956,N_23791,N_23822);
xor U24957 (N_24957,N_23828,N_23919);
or U24958 (N_24958,N_23977,N_24189);
and U24959 (N_24959,N_24109,N_24113);
or U24960 (N_24960,N_23824,N_23902);
or U24961 (N_24961,N_24128,N_24215);
or U24962 (N_24962,N_23952,N_24304);
or U24963 (N_24963,N_23959,N_24369);
xor U24964 (N_24964,N_24373,N_23881);
nand U24965 (N_24965,N_23917,N_24351);
or U24966 (N_24966,N_23779,N_24073);
and U24967 (N_24967,N_24149,N_24112);
or U24968 (N_24968,N_24226,N_24282);
nor U24969 (N_24969,N_23932,N_24233);
and U24970 (N_24970,N_24237,N_24036);
or U24971 (N_24971,N_23811,N_23855);
xor U24972 (N_24972,N_24374,N_23920);
or U24973 (N_24973,N_24193,N_24306);
and U24974 (N_24974,N_24086,N_24045);
and U24975 (N_24975,N_24170,N_24155);
and U24976 (N_24976,N_24067,N_24185);
nor U24977 (N_24977,N_24348,N_24165);
nand U24978 (N_24978,N_23818,N_24263);
nor U24979 (N_24979,N_24168,N_23815);
nand U24980 (N_24980,N_24356,N_23836);
and U24981 (N_24981,N_23936,N_23788);
nor U24982 (N_24982,N_24272,N_23818);
nor U24983 (N_24983,N_24329,N_24012);
or U24984 (N_24984,N_23894,N_24042);
nand U24985 (N_24985,N_23868,N_24312);
or U24986 (N_24986,N_24137,N_24200);
nand U24987 (N_24987,N_24316,N_23821);
or U24988 (N_24988,N_24082,N_23974);
or U24989 (N_24989,N_24035,N_23936);
and U24990 (N_24990,N_24268,N_23922);
and U24991 (N_24991,N_23817,N_24036);
xnor U24992 (N_24992,N_23874,N_23765);
or U24993 (N_24993,N_23861,N_24041);
or U24994 (N_24994,N_23854,N_24044);
nand U24995 (N_24995,N_23836,N_23842);
and U24996 (N_24996,N_23796,N_24041);
nand U24997 (N_24997,N_24008,N_23889);
nand U24998 (N_24998,N_23853,N_24053);
nand U24999 (N_24999,N_24169,N_24031);
and UO_0 (O_0,N_24594,N_24826);
or UO_1 (O_1,N_24544,N_24546);
nand UO_2 (O_2,N_24605,N_24726);
nor UO_3 (O_3,N_24385,N_24378);
or UO_4 (O_4,N_24529,N_24450);
and UO_5 (O_5,N_24625,N_24487);
or UO_6 (O_6,N_24716,N_24603);
or UO_7 (O_7,N_24819,N_24630);
and UO_8 (O_8,N_24823,N_24380);
or UO_9 (O_9,N_24855,N_24542);
xor UO_10 (O_10,N_24668,N_24572);
nand UO_11 (O_11,N_24760,N_24938);
nor UO_12 (O_12,N_24587,N_24935);
and UO_13 (O_13,N_24772,N_24836);
xnor UO_14 (O_14,N_24618,N_24690);
xnor UO_15 (O_15,N_24900,N_24859);
and UO_16 (O_16,N_24545,N_24692);
nor UO_17 (O_17,N_24547,N_24914);
nand UO_18 (O_18,N_24850,N_24727);
nand UO_19 (O_19,N_24660,N_24803);
or UO_20 (O_20,N_24808,N_24469);
nor UO_21 (O_21,N_24585,N_24419);
or UO_22 (O_22,N_24426,N_24937);
nor UO_23 (O_23,N_24825,N_24944);
or UO_24 (O_24,N_24619,N_24551);
xnor UO_25 (O_25,N_24838,N_24467);
nor UO_26 (O_26,N_24767,N_24735);
nand UO_27 (O_27,N_24460,N_24746);
or UO_28 (O_28,N_24991,N_24595);
nand UO_29 (O_29,N_24701,N_24908);
nor UO_30 (O_30,N_24844,N_24533);
and UO_31 (O_31,N_24780,N_24503);
and UO_32 (O_32,N_24375,N_24440);
nor UO_33 (O_33,N_24854,N_24789);
nand UO_34 (O_34,N_24747,N_24834);
or UO_35 (O_35,N_24784,N_24428);
or UO_36 (O_36,N_24620,N_24764);
nor UO_37 (O_37,N_24430,N_24624);
xor UO_38 (O_38,N_24878,N_24442);
nor UO_39 (O_39,N_24591,N_24400);
nor UO_40 (O_40,N_24616,N_24664);
and UO_41 (O_41,N_24583,N_24961);
and UO_42 (O_42,N_24876,N_24970);
xor UO_43 (O_43,N_24897,N_24907);
or UO_44 (O_44,N_24699,N_24622);
and UO_45 (O_45,N_24665,N_24376);
or UO_46 (O_46,N_24471,N_24639);
nor UO_47 (O_47,N_24576,N_24980);
xor UO_48 (O_48,N_24738,N_24387);
nor UO_49 (O_49,N_24675,N_24636);
nor UO_50 (O_50,N_24882,N_24852);
or UO_51 (O_51,N_24996,N_24453);
or UO_52 (O_52,N_24475,N_24521);
xor UO_53 (O_53,N_24695,N_24895);
and UO_54 (O_54,N_24515,N_24885);
or UO_55 (O_55,N_24945,N_24432);
nand UO_56 (O_56,N_24557,N_24507);
and UO_57 (O_57,N_24439,N_24898);
and UO_58 (O_58,N_24959,N_24558);
nand UO_59 (O_59,N_24652,N_24863);
and UO_60 (O_60,N_24482,N_24593);
nand UO_61 (O_61,N_24653,N_24395);
or UO_62 (O_62,N_24802,N_24755);
nand UO_63 (O_63,N_24899,N_24661);
and UO_64 (O_64,N_24717,N_24614);
or UO_65 (O_65,N_24988,N_24797);
nand UO_66 (O_66,N_24833,N_24553);
nand UO_67 (O_67,N_24928,N_24912);
nand UO_68 (O_68,N_24768,N_24548);
nor UO_69 (O_69,N_24596,N_24924);
nor UO_70 (O_70,N_24990,N_24835);
and UO_71 (O_71,N_24511,N_24728);
nor UO_72 (O_72,N_24421,N_24401);
nand UO_73 (O_73,N_24436,N_24771);
or UO_74 (O_74,N_24444,N_24406);
or UO_75 (O_75,N_24659,N_24496);
nor UO_76 (O_76,N_24891,N_24472);
or UO_77 (O_77,N_24598,N_24848);
or UO_78 (O_78,N_24839,N_24677);
nand UO_79 (O_79,N_24589,N_24462);
xnor UO_80 (O_80,N_24381,N_24934);
xnor UO_81 (O_81,N_24402,N_24745);
nand UO_82 (O_82,N_24602,N_24555);
nand UO_83 (O_83,N_24447,N_24811);
nand UO_84 (O_84,N_24530,N_24657);
or UO_85 (O_85,N_24921,N_24386);
nor UO_86 (O_86,N_24520,N_24805);
and UO_87 (O_87,N_24643,N_24845);
nor UO_88 (O_88,N_24379,N_24902);
nand UO_89 (O_89,N_24497,N_24479);
and UO_90 (O_90,N_24989,N_24458);
nand UO_91 (O_91,N_24733,N_24568);
nor UO_92 (O_92,N_24837,N_24929);
nor UO_93 (O_93,N_24744,N_24398);
nor UO_94 (O_94,N_24654,N_24608);
nand UO_95 (O_95,N_24434,N_24474);
or UO_96 (O_96,N_24539,N_24886);
nand UO_97 (O_97,N_24470,N_24752);
nand UO_98 (O_98,N_24574,N_24392);
xor UO_99 (O_99,N_24600,N_24791);
nand UO_100 (O_100,N_24508,N_24906);
or UO_101 (O_101,N_24820,N_24864);
and UO_102 (O_102,N_24983,N_24810);
nor UO_103 (O_103,N_24667,N_24923);
or UO_104 (O_104,N_24627,N_24821);
xnor UO_105 (O_105,N_24623,N_24712);
nor UO_106 (O_106,N_24998,N_24851);
and UO_107 (O_107,N_24575,N_24681);
xor UO_108 (O_108,N_24679,N_24538);
nor UO_109 (O_109,N_24933,N_24713);
or UO_110 (O_110,N_24960,N_24455);
nor UO_111 (O_111,N_24765,N_24840);
or UO_112 (O_112,N_24707,N_24413);
nand UO_113 (O_113,N_24932,N_24941);
and UO_114 (O_114,N_24689,N_24957);
or UO_115 (O_115,N_24883,N_24815);
nor UO_116 (O_116,N_24422,N_24562);
nor UO_117 (O_117,N_24429,N_24448);
nand UO_118 (O_118,N_24865,N_24621);
nand UO_119 (O_119,N_24414,N_24971);
nor UO_120 (O_120,N_24409,N_24809);
nor UO_121 (O_121,N_24489,N_24952);
nor UO_122 (O_122,N_24749,N_24473);
nand UO_123 (O_123,N_24495,N_24441);
nand UO_124 (O_124,N_24869,N_24818);
or UO_125 (O_125,N_24706,N_24666);
nor UO_126 (O_126,N_24804,N_24569);
or UO_127 (O_127,N_24682,N_24676);
nand UO_128 (O_128,N_24955,N_24919);
nor UO_129 (O_129,N_24481,N_24947);
nand UO_130 (O_130,N_24564,N_24629);
nor UO_131 (O_131,N_24565,N_24377);
or UO_132 (O_132,N_24787,N_24829);
nor UO_133 (O_133,N_24531,N_24936);
xnor UO_134 (O_134,N_24581,N_24986);
nor UO_135 (O_135,N_24718,N_24425);
xnor UO_136 (O_136,N_24418,N_24396);
nand UO_137 (O_137,N_24563,N_24723);
nand UO_138 (O_138,N_24694,N_24650);
or UO_139 (O_139,N_24801,N_24451);
and UO_140 (O_140,N_24889,N_24856);
and UO_141 (O_141,N_24642,N_24662);
or UO_142 (O_142,N_24540,N_24720);
or UO_143 (O_143,N_24841,N_24527);
and UO_144 (O_144,N_24537,N_24601);
nand UO_145 (O_145,N_24758,N_24397);
and UO_146 (O_146,N_24948,N_24493);
or UO_147 (O_147,N_24740,N_24405);
nor UO_148 (O_148,N_24710,N_24794);
xor UO_149 (O_149,N_24751,N_24890);
and UO_150 (O_150,N_24590,N_24756);
or UO_151 (O_151,N_24696,N_24795);
nand UO_152 (O_152,N_24702,N_24862);
xnor UO_153 (O_153,N_24554,N_24573);
nand UO_154 (O_154,N_24817,N_24977);
nand UO_155 (O_155,N_24867,N_24644);
or UO_156 (O_156,N_24488,N_24832);
nand UO_157 (O_157,N_24582,N_24979);
nand UO_158 (O_158,N_24922,N_24670);
and UO_159 (O_159,N_24615,N_24995);
nor UO_160 (O_160,N_24592,N_24513);
nand UO_161 (O_161,N_24950,N_24648);
and UO_162 (O_162,N_24412,N_24438);
nor UO_163 (O_163,N_24927,N_24824);
nor UO_164 (O_164,N_24626,N_24431);
or UO_165 (O_165,N_24446,N_24478);
or UO_166 (O_166,N_24697,N_24466);
and UO_167 (O_167,N_24982,N_24394);
or UO_168 (O_168,N_24917,N_24655);
nor UO_169 (O_169,N_24516,N_24483);
and UO_170 (O_170,N_24584,N_24753);
nand UO_171 (O_171,N_24464,N_24500);
nand UO_172 (O_172,N_24484,N_24566);
xor UO_173 (O_173,N_24498,N_24816);
nor UO_174 (O_174,N_24671,N_24904);
nor UO_175 (O_175,N_24910,N_24762);
nand UO_176 (O_176,N_24777,N_24510);
nor UO_177 (O_177,N_24724,N_24393);
xnor UO_178 (O_178,N_24871,N_24857);
xor UO_179 (O_179,N_24509,N_24433);
or UO_180 (O_180,N_24388,N_24903);
nor UO_181 (O_181,N_24975,N_24452);
nand UO_182 (O_182,N_24609,N_24610);
and UO_183 (O_183,N_24637,N_24786);
nand UO_184 (O_184,N_24404,N_24981);
and UO_185 (O_185,N_24708,N_24522);
xor UO_186 (O_186,N_24965,N_24502);
nor UO_187 (O_187,N_24534,N_24514);
nand UO_188 (O_188,N_24651,N_24384);
or UO_189 (O_189,N_24663,N_24486);
nand UO_190 (O_190,N_24972,N_24407);
nand UO_191 (O_191,N_24750,N_24913);
nor UO_192 (O_192,N_24911,N_24640);
and UO_193 (O_193,N_24526,N_24577);
or UO_194 (O_194,N_24443,N_24847);
or UO_195 (O_195,N_24842,N_24783);
xor UO_196 (O_196,N_24992,N_24647);
or UO_197 (O_197,N_24870,N_24729);
nor UO_198 (O_198,N_24843,N_24491);
nor UO_199 (O_199,N_24631,N_24748);
xnor UO_200 (O_200,N_24814,N_24722);
and UO_201 (O_201,N_24549,N_24468);
or UO_202 (O_202,N_24456,N_24974);
and UO_203 (O_203,N_24628,N_24698);
and UO_204 (O_204,N_24711,N_24757);
or UO_205 (O_205,N_24427,N_24680);
nand UO_206 (O_206,N_24813,N_24459);
or UO_207 (O_207,N_24997,N_24683);
or UO_208 (O_208,N_24776,N_24967);
nor UO_209 (O_209,N_24408,N_24946);
or UO_210 (O_210,N_24705,N_24580);
nand UO_211 (O_211,N_24943,N_24861);
xor UO_212 (O_212,N_24480,N_24704);
or UO_213 (O_213,N_24918,N_24905);
nor UO_214 (O_214,N_24892,N_24492);
nand UO_215 (O_215,N_24822,N_24512);
and UO_216 (O_216,N_24968,N_24725);
xnor UO_217 (O_217,N_24930,N_24896);
nor UO_218 (O_218,N_24501,N_24881);
or UO_219 (O_219,N_24966,N_24523);
nor UO_220 (O_220,N_24411,N_24579);
nor UO_221 (O_221,N_24463,N_24763);
nand UO_222 (O_222,N_24963,N_24525);
and UO_223 (O_223,N_24672,N_24807);
nand UO_224 (O_224,N_24984,N_24812);
and UO_225 (O_225,N_24994,N_24504);
or UO_226 (O_226,N_24437,N_24449);
and UO_227 (O_227,N_24638,N_24737);
nand UO_228 (O_228,N_24956,N_24879);
and UO_229 (O_229,N_24828,N_24382);
nor UO_230 (O_230,N_24465,N_24939);
and UO_231 (O_231,N_24559,N_24949);
or UO_232 (O_232,N_24894,N_24773);
and UO_233 (O_233,N_24785,N_24417);
nor UO_234 (O_234,N_24798,N_24673);
and UO_235 (O_235,N_24688,N_24719);
nor UO_236 (O_236,N_24543,N_24477);
nand UO_237 (O_237,N_24714,N_24734);
nand UO_238 (O_238,N_24383,N_24742);
or UO_239 (O_239,N_24703,N_24953);
or UO_240 (O_240,N_24846,N_24390);
and UO_241 (O_241,N_24678,N_24779);
or UO_242 (O_242,N_24853,N_24646);
and UO_243 (O_243,N_24403,N_24769);
or UO_244 (O_244,N_24888,N_24641);
or UO_245 (O_245,N_24550,N_24873);
nor UO_246 (O_246,N_24860,N_24736);
or UO_247 (O_247,N_24391,N_24954);
xnor UO_248 (O_248,N_24759,N_24782);
and UO_249 (O_249,N_24790,N_24931);
nor UO_250 (O_250,N_24686,N_24920);
nand UO_251 (O_251,N_24399,N_24951);
nor UO_252 (O_252,N_24942,N_24887);
and UO_253 (O_253,N_24800,N_24506);
nand UO_254 (O_254,N_24490,N_24969);
nand UO_255 (O_255,N_24423,N_24872);
and UO_256 (O_256,N_24880,N_24674);
or UO_257 (O_257,N_24732,N_24962);
nor UO_258 (O_258,N_24754,N_24532);
xnor UO_259 (O_259,N_24987,N_24611);
or UO_260 (O_260,N_24877,N_24541);
nor UO_261 (O_261,N_24649,N_24617);
or UO_262 (O_262,N_24567,N_24536);
nor UO_263 (O_263,N_24519,N_24604);
or UO_264 (O_264,N_24976,N_24766);
or UO_265 (O_265,N_24739,N_24597);
or UO_266 (O_266,N_24978,N_24691);
nand UO_267 (O_267,N_24645,N_24517);
xor UO_268 (O_268,N_24830,N_24457);
nor UO_269 (O_269,N_24571,N_24461);
nor UO_270 (O_270,N_24633,N_24884);
nor UO_271 (O_271,N_24775,N_24424);
nand UO_272 (O_272,N_24792,N_24445);
nand UO_273 (O_273,N_24799,N_24858);
and UO_274 (O_274,N_24669,N_24999);
and UO_275 (O_275,N_24435,N_24925);
or UO_276 (O_276,N_24874,N_24410);
nand UO_277 (O_277,N_24687,N_24454);
nor UO_278 (O_278,N_24556,N_24709);
or UO_279 (O_279,N_24535,N_24586);
and UO_280 (O_280,N_24741,N_24893);
nand UO_281 (O_281,N_24875,N_24827);
nor UO_282 (O_282,N_24528,N_24743);
or UO_283 (O_283,N_24607,N_24774);
and UO_284 (O_284,N_24866,N_24389);
or UO_285 (O_285,N_24494,N_24721);
nor UO_286 (O_286,N_24909,N_24831);
and UO_287 (O_287,N_24700,N_24420);
or UO_288 (O_288,N_24916,N_24793);
or UO_289 (O_289,N_24485,N_24973);
nand UO_290 (O_290,N_24499,N_24761);
or UO_291 (O_291,N_24731,N_24505);
and UO_292 (O_292,N_24788,N_24901);
nand UO_293 (O_293,N_24415,N_24926);
xor UO_294 (O_294,N_24476,N_24606);
nor UO_295 (O_295,N_24570,N_24781);
or UO_296 (O_296,N_24552,N_24518);
xnor UO_297 (O_297,N_24578,N_24964);
and UO_298 (O_298,N_24658,N_24915);
and UO_299 (O_299,N_24560,N_24806);
nor UO_300 (O_300,N_24613,N_24561);
and UO_301 (O_301,N_24612,N_24524);
xnor UO_302 (O_302,N_24635,N_24685);
xor UO_303 (O_303,N_24634,N_24778);
and UO_304 (O_304,N_24868,N_24693);
nand UO_305 (O_305,N_24416,N_24684);
xnor UO_306 (O_306,N_24940,N_24993);
or UO_307 (O_307,N_24599,N_24715);
or UO_308 (O_308,N_24985,N_24632);
or UO_309 (O_309,N_24796,N_24958);
and UO_310 (O_310,N_24730,N_24656);
or UO_311 (O_311,N_24588,N_24770);
nand UO_312 (O_312,N_24849,N_24811);
xor UO_313 (O_313,N_24717,N_24735);
or UO_314 (O_314,N_24787,N_24534);
or UO_315 (O_315,N_24590,N_24661);
xor UO_316 (O_316,N_24552,N_24986);
and UO_317 (O_317,N_24970,N_24791);
and UO_318 (O_318,N_24610,N_24835);
nor UO_319 (O_319,N_24681,N_24407);
nand UO_320 (O_320,N_24442,N_24833);
nand UO_321 (O_321,N_24417,N_24606);
nor UO_322 (O_322,N_24481,N_24634);
nand UO_323 (O_323,N_24454,N_24789);
xor UO_324 (O_324,N_24565,N_24410);
or UO_325 (O_325,N_24549,N_24474);
nand UO_326 (O_326,N_24831,N_24627);
nor UO_327 (O_327,N_24878,N_24850);
and UO_328 (O_328,N_24487,N_24692);
nor UO_329 (O_329,N_24619,N_24990);
nand UO_330 (O_330,N_24780,N_24421);
and UO_331 (O_331,N_24861,N_24834);
and UO_332 (O_332,N_24772,N_24478);
and UO_333 (O_333,N_24701,N_24515);
nand UO_334 (O_334,N_24589,N_24851);
nand UO_335 (O_335,N_24508,N_24792);
or UO_336 (O_336,N_24635,N_24771);
or UO_337 (O_337,N_24717,N_24841);
xor UO_338 (O_338,N_24420,N_24797);
nand UO_339 (O_339,N_24880,N_24688);
nor UO_340 (O_340,N_24808,N_24770);
nor UO_341 (O_341,N_24782,N_24555);
or UO_342 (O_342,N_24517,N_24415);
nand UO_343 (O_343,N_24935,N_24956);
or UO_344 (O_344,N_24409,N_24787);
and UO_345 (O_345,N_24955,N_24515);
nor UO_346 (O_346,N_24448,N_24451);
or UO_347 (O_347,N_24660,N_24489);
nor UO_348 (O_348,N_24662,N_24634);
nand UO_349 (O_349,N_24443,N_24980);
xnor UO_350 (O_350,N_24472,N_24957);
nand UO_351 (O_351,N_24916,N_24470);
nor UO_352 (O_352,N_24376,N_24463);
or UO_353 (O_353,N_24960,N_24806);
nor UO_354 (O_354,N_24986,N_24573);
or UO_355 (O_355,N_24983,N_24505);
and UO_356 (O_356,N_24827,N_24823);
nor UO_357 (O_357,N_24713,N_24465);
and UO_358 (O_358,N_24998,N_24783);
nand UO_359 (O_359,N_24787,N_24385);
nor UO_360 (O_360,N_24755,N_24550);
nor UO_361 (O_361,N_24951,N_24609);
xnor UO_362 (O_362,N_24438,N_24967);
and UO_363 (O_363,N_24389,N_24391);
or UO_364 (O_364,N_24903,N_24722);
nor UO_365 (O_365,N_24387,N_24459);
nor UO_366 (O_366,N_24632,N_24694);
or UO_367 (O_367,N_24522,N_24783);
and UO_368 (O_368,N_24740,N_24739);
or UO_369 (O_369,N_24652,N_24942);
nand UO_370 (O_370,N_24870,N_24474);
nor UO_371 (O_371,N_24462,N_24763);
nor UO_372 (O_372,N_24965,N_24466);
or UO_373 (O_373,N_24493,N_24734);
nand UO_374 (O_374,N_24932,N_24487);
nand UO_375 (O_375,N_24940,N_24492);
or UO_376 (O_376,N_24947,N_24375);
or UO_377 (O_377,N_24509,N_24697);
nand UO_378 (O_378,N_24748,N_24715);
nor UO_379 (O_379,N_24996,N_24466);
or UO_380 (O_380,N_24773,N_24681);
or UO_381 (O_381,N_24477,N_24784);
nor UO_382 (O_382,N_24612,N_24903);
nor UO_383 (O_383,N_24638,N_24459);
and UO_384 (O_384,N_24886,N_24816);
nor UO_385 (O_385,N_24588,N_24701);
nor UO_386 (O_386,N_24741,N_24652);
or UO_387 (O_387,N_24587,N_24625);
and UO_388 (O_388,N_24615,N_24558);
xor UO_389 (O_389,N_24965,N_24921);
nand UO_390 (O_390,N_24483,N_24839);
and UO_391 (O_391,N_24410,N_24609);
nor UO_392 (O_392,N_24772,N_24585);
or UO_393 (O_393,N_24989,N_24457);
xnor UO_394 (O_394,N_24640,N_24755);
and UO_395 (O_395,N_24673,N_24890);
and UO_396 (O_396,N_24800,N_24650);
nor UO_397 (O_397,N_24386,N_24856);
or UO_398 (O_398,N_24407,N_24961);
nand UO_399 (O_399,N_24730,N_24587);
and UO_400 (O_400,N_24773,N_24445);
xnor UO_401 (O_401,N_24420,N_24403);
and UO_402 (O_402,N_24412,N_24479);
xnor UO_403 (O_403,N_24744,N_24864);
or UO_404 (O_404,N_24507,N_24901);
nor UO_405 (O_405,N_24751,N_24588);
and UO_406 (O_406,N_24793,N_24780);
or UO_407 (O_407,N_24731,N_24452);
and UO_408 (O_408,N_24821,N_24789);
nor UO_409 (O_409,N_24544,N_24384);
xnor UO_410 (O_410,N_24605,N_24704);
and UO_411 (O_411,N_24404,N_24776);
and UO_412 (O_412,N_24540,N_24425);
nand UO_413 (O_413,N_24610,N_24993);
nand UO_414 (O_414,N_24716,N_24895);
and UO_415 (O_415,N_24899,N_24598);
xnor UO_416 (O_416,N_24507,N_24849);
nor UO_417 (O_417,N_24500,N_24980);
or UO_418 (O_418,N_24430,N_24622);
or UO_419 (O_419,N_24923,N_24766);
or UO_420 (O_420,N_24901,N_24555);
and UO_421 (O_421,N_24896,N_24452);
and UO_422 (O_422,N_24620,N_24769);
and UO_423 (O_423,N_24442,N_24855);
and UO_424 (O_424,N_24922,N_24659);
xnor UO_425 (O_425,N_24526,N_24550);
and UO_426 (O_426,N_24982,N_24530);
and UO_427 (O_427,N_24525,N_24852);
or UO_428 (O_428,N_24590,N_24820);
xnor UO_429 (O_429,N_24907,N_24490);
nor UO_430 (O_430,N_24888,N_24886);
nand UO_431 (O_431,N_24385,N_24998);
or UO_432 (O_432,N_24573,N_24868);
or UO_433 (O_433,N_24729,N_24458);
nor UO_434 (O_434,N_24660,N_24593);
and UO_435 (O_435,N_24810,N_24542);
or UO_436 (O_436,N_24790,N_24724);
xor UO_437 (O_437,N_24958,N_24771);
xor UO_438 (O_438,N_24697,N_24607);
nand UO_439 (O_439,N_24632,N_24940);
nor UO_440 (O_440,N_24982,N_24743);
or UO_441 (O_441,N_24754,N_24622);
and UO_442 (O_442,N_24781,N_24730);
and UO_443 (O_443,N_24433,N_24518);
and UO_444 (O_444,N_24418,N_24700);
xnor UO_445 (O_445,N_24691,N_24966);
nor UO_446 (O_446,N_24617,N_24896);
or UO_447 (O_447,N_24905,N_24747);
nand UO_448 (O_448,N_24637,N_24749);
or UO_449 (O_449,N_24926,N_24574);
and UO_450 (O_450,N_24752,N_24972);
or UO_451 (O_451,N_24975,N_24807);
or UO_452 (O_452,N_24469,N_24425);
and UO_453 (O_453,N_24823,N_24639);
or UO_454 (O_454,N_24993,N_24726);
or UO_455 (O_455,N_24601,N_24832);
nor UO_456 (O_456,N_24618,N_24819);
and UO_457 (O_457,N_24877,N_24436);
and UO_458 (O_458,N_24593,N_24873);
nand UO_459 (O_459,N_24468,N_24560);
and UO_460 (O_460,N_24739,N_24789);
nor UO_461 (O_461,N_24472,N_24825);
and UO_462 (O_462,N_24962,N_24691);
and UO_463 (O_463,N_24400,N_24694);
and UO_464 (O_464,N_24526,N_24621);
nor UO_465 (O_465,N_24414,N_24766);
xor UO_466 (O_466,N_24685,N_24957);
xnor UO_467 (O_467,N_24928,N_24535);
or UO_468 (O_468,N_24825,N_24460);
nor UO_469 (O_469,N_24953,N_24738);
and UO_470 (O_470,N_24431,N_24575);
xnor UO_471 (O_471,N_24539,N_24560);
nand UO_472 (O_472,N_24954,N_24577);
and UO_473 (O_473,N_24856,N_24473);
nor UO_474 (O_474,N_24869,N_24458);
nand UO_475 (O_475,N_24748,N_24890);
xor UO_476 (O_476,N_24787,N_24813);
xnor UO_477 (O_477,N_24651,N_24923);
xor UO_478 (O_478,N_24610,N_24502);
nand UO_479 (O_479,N_24707,N_24863);
or UO_480 (O_480,N_24876,N_24520);
and UO_481 (O_481,N_24782,N_24937);
nand UO_482 (O_482,N_24446,N_24686);
or UO_483 (O_483,N_24656,N_24655);
nor UO_484 (O_484,N_24581,N_24895);
xnor UO_485 (O_485,N_24560,N_24900);
nand UO_486 (O_486,N_24813,N_24780);
or UO_487 (O_487,N_24801,N_24405);
or UO_488 (O_488,N_24511,N_24879);
nor UO_489 (O_489,N_24539,N_24758);
nor UO_490 (O_490,N_24629,N_24533);
xnor UO_491 (O_491,N_24761,N_24441);
nor UO_492 (O_492,N_24448,N_24839);
nor UO_493 (O_493,N_24887,N_24695);
nor UO_494 (O_494,N_24424,N_24839);
nand UO_495 (O_495,N_24998,N_24803);
nor UO_496 (O_496,N_24736,N_24994);
and UO_497 (O_497,N_24456,N_24936);
and UO_498 (O_498,N_24991,N_24907);
and UO_499 (O_499,N_24697,N_24615);
xor UO_500 (O_500,N_24397,N_24936);
or UO_501 (O_501,N_24587,N_24975);
nand UO_502 (O_502,N_24375,N_24583);
and UO_503 (O_503,N_24923,N_24845);
nor UO_504 (O_504,N_24677,N_24866);
nor UO_505 (O_505,N_24868,N_24678);
and UO_506 (O_506,N_24777,N_24547);
or UO_507 (O_507,N_24794,N_24590);
and UO_508 (O_508,N_24793,N_24646);
xor UO_509 (O_509,N_24907,N_24749);
or UO_510 (O_510,N_24824,N_24814);
and UO_511 (O_511,N_24453,N_24653);
or UO_512 (O_512,N_24450,N_24643);
and UO_513 (O_513,N_24789,N_24502);
and UO_514 (O_514,N_24920,N_24886);
nand UO_515 (O_515,N_24492,N_24657);
and UO_516 (O_516,N_24710,N_24407);
and UO_517 (O_517,N_24975,N_24700);
nand UO_518 (O_518,N_24775,N_24421);
or UO_519 (O_519,N_24526,N_24397);
and UO_520 (O_520,N_24501,N_24748);
and UO_521 (O_521,N_24590,N_24844);
or UO_522 (O_522,N_24495,N_24616);
and UO_523 (O_523,N_24491,N_24661);
or UO_524 (O_524,N_24994,N_24461);
nor UO_525 (O_525,N_24386,N_24431);
nor UO_526 (O_526,N_24553,N_24929);
nand UO_527 (O_527,N_24556,N_24921);
xor UO_528 (O_528,N_24798,N_24473);
nor UO_529 (O_529,N_24607,N_24513);
nor UO_530 (O_530,N_24787,N_24504);
or UO_531 (O_531,N_24552,N_24780);
nor UO_532 (O_532,N_24702,N_24695);
nand UO_533 (O_533,N_24759,N_24390);
xor UO_534 (O_534,N_24791,N_24709);
nor UO_535 (O_535,N_24404,N_24471);
nand UO_536 (O_536,N_24716,N_24844);
or UO_537 (O_537,N_24542,N_24817);
nor UO_538 (O_538,N_24964,N_24595);
xor UO_539 (O_539,N_24463,N_24629);
nor UO_540 (O_540,N_24955,N_24632);
nand UO_541 (O_541,N_24681,N_24876);
and UO_542 (O_542,N_24707,N_24881);
or UO_543 (O_543,N_24572,N_24895);
and UO_544 (O_544,N_24465,N_24753);
and UO_545 (O_545,N_24659,N_24961);
xor UO_546 (O_546,N_24834,N_24958);
nand UO_547 (O_547,N_24761,N_24984);
nor UO_548 (O_548,N_24796,N_24627);
and UO_549 (O_549,N_24674,N_24882);
and UO_550 (O_550,N_24602,N_24752);
xor UO_551 (O_551,N_24457,N_24950);
xnor UO_552 (O_552,N_24955,N_24936);
or UO_553 (O_553,N_24889,N_24694);
nor UO_554 (O_554,N_24434,N_24751);
nand UO_555 (O_555,N_24986,N_24937);
nand UO_556 (O_556,N_24781,N_24977);
and UO_557 (O_557,N_24501,N_24869);
nand UO_558 (O_558,N_24554,N_24967);
xor UO_559 (O_559,N_24884,N_24831);
nor UO_560 (O_560,N_24736,N_24608);
nand UO_561 (O_561,N_24676,N_24564);
nand UO_562 (O_562,N_24699,N_24405);
nand UO_563 (O_563,N_24486,N_24685);
xnor UO_564 (O_564,N_24795,N_24993);
or UO_565 (O_565,N_24599,N_24559);
xnor UO_566 (O_566,N_24978,N_24439);
and UO_567 (O_567,N_24471,N_24516);
nor UO_568 (O_568,N_24678,N_24866);
or UO_569 (O_569,N_24630,N_24861);
nor UO_570 (O_570,N_24956,N_24840);
or UO_571 (O_571,N_24795,N_24815);
nand UO_572 (O_572,N_24799,N_24931);
nor UO_573 (O_573,N_24859,N_24817);
nand UO_574 (O_574,N_24935,N_24779);
or UO_575 (O_575,N_24520,N_24551);
or UO_576 (O_576,N_24541,N_24673);
and UO_577 (O_577,N_24638,N_24891);
and UO_578 (O_578,N_24572,N_24426);
xnor UO_579 (O_579,N_24418,N_24544);
and UO_580 (O_580,N_24663,N_24441);
and UO_581 (O_581,N_24847,N_24417);
and UO_582 (O_582,N_24993,N_24621);
and UO_583 (O_583,N_24471,N_24863);
or UO_584 (O_584,N_24953,N_24705);
nand UO_585 (O_585,N_24893,N_24922);
nor UO_586 (O_586,N_24487,N_24849);
nor UO_587 (O_587,N_24415,N_24516);
nor UO_588 (O_588,N_24482,N_24379);
xnor UO_589 (O_589,N_24616,N_24813);
or UO_590 (O_590,N_24772,N_24638);
and UO_591 (O_591,N_24388,N_24624);
nand UO_592 (O_592,N_24938,N_24499);
or UO_593 (O_593,N_24844,N_24450);
or UO_594 (O_594,N_24842,N_24681);
or UO_595 (O_595,N_24734,N_24909);
nand UO_596 (O_596,N_24757,N_24894);
nor UO_597 (O_597,N_24575,N_24661);
or UO_598 (O_598,N_24491,N_24882);
nor UO_599 (O_599,N_24531,N_24956);
nand UO_600 (O_600,N_24655,N_24931);
or UO_601 (O_601,N_24977,N_24523);
nor UO_602 (O_602,N_24621,N_24630);
and UO_603 (O_603,N_24863,N_24937);
and UO_604 (O_604,N_24988,N_24598);
nor UO_605 (O_605,N_24537,N_24560);
nand UO_606 (O_606,N_24717,N_24454);
xor UO_607 (O_607,N_24415,N_24590);
xnor UO_608 (O_608,N_24528,N_24380);
nand UO_609 (O_609,N_24707,N_24883);
nand UO_610 (O_610,N_24911,N_24765);
and UO_611 (O_611,N_24830,N_24813);
nor UO_612 (O_612,N_24773,N_24697);
and UO_613 (O_613,N_24674,N_24937);
nand UO_614 (O_614,N_24993,N_24902);
or UO_615 (O_615,N_24544,N_24461);
nor UO_616 (O_616,N_24541,N_24664);
nor UO_617 (O_617,N_24894,N_24940);
nor UO_618 (O_618,N_24731,N_24937);
nor UO_619 (O_619,N_24992,N_24679);
and UO_620 (O_620,N_24584,N_24823);
or UO_621 (O_621,N_24613,N_24615);
nand UO_622 (O_622,N_24706,N_24461);
or UO_623 (O_623,N_24442,N_24941);
and UO_624 (O_624,N_24462,N_24732);
or UO_625 (O_625,N_24571,N_24566);
nand UO_626 (O_626,N_24550,N_24903);
nand UO_627 (O_627,N_24717,N_24727);
and UO_628 (O_628,N_24591,N_24479);
xnor UO_629 (O_629,N_24731,N_24674);
nor UO_630 (O_630,N_24958,N_24936);
nand UO_631 (O_631,N_24587,N_24458);
or UO_632 (O_632,N_24506,N_24608);
or UO_633 (O_633,N_24537,N_24491);
nor UO_634 (O_634,N_24527,N_24823);
nor UO_635 (O_635,N_24729,N_24500);
or UO_636 (O_636,N_24852,N_24644);
or UO_637 (O_637,N_24581,N_24561);
nor UO_638 (O_638,N_24430,N_24883);
or UO_639 (O_639,N_24627,N_24833);
nand UO_640 (O_640,N_24598,N_24673);
and UO_641 (O_641,N_24690,N_24752);
xor UO_642 (O_642,N_24623,N_24754);
nor UO_643 (O_643,N_24461,N_24845);
nand UO_644 (O_644,N_24796,N_24464);
nand UO_645 (O_645,N_24674,N_24382);
nor UO_646 (O_646,N_24593,N_24764);
nor UO_647 (O_647,N_24751,N_24836);
nand UO_648 (O_648,N_24883,N_24985);
and UO_649 (O_649,N_24612,N_24901);
or UO_650 (O_650,N_24914,N_24933);
nor UO_651 (O_651,N_24752,N_24821);
nor UO_652 (O_652,N_24418,N_24545);
nand UO_653 (O_653,N_24875,N_24921);
and UO_654 (O_654,N_24607,N_24400);
and UO_655 (O_655,N_24972,N_24436);
and UO_656 (O_656,N_24653,N_24485);
and UO_657 (O_657,N_24438,N_24680);
or UO_658 (O_658,N_24386,N_24944);
and UO_659 (O_659,N_24440,N_24873);
and UO_660 (O_660,N_24955,N_24469);
nand UO_661 (O_661,N_24829,N_24383);
or UO_662 (O_662,N_24854,N_24819);
or UO_663 (O_663,N_24990,N_24636);
nand UO_664 (O_664,N_24894,N_24472);
and UO_665 (O_665,N_24756,N_24682);
nand UO_666 (O_666,N_24403,N_24933);
and UO_667 (O_667,N_24533,N_24794);
nor UO_668 (O_668,N_24761,N_24846);
or UO_669 (O_669,N_24771,N_24686);
or UO_670 (O_670,N_24999,N_24922);
nand UO_671 (O_671,N_24684,N_24432);
nand UO_672 (O_672,N_24633,N_24469);
nor UO_673 (O_673,N_24897,N_24899);
nor UO_674 (O_674,N_24505,N_24890);
nand UO_675 (O_675,N_24567,N_24771);
or UO_676 (O_676,N_24411,N_24564);
and UO_677 (O_677,N_24867,N_24913);
nand UO_678 (O_678,N_24435,N_24715);
nand UO_679 (O_679,N_24866,N_24798);
nor UO_680 (O_680,N_24831,N_24490);
and UO_681 (O_681,N_24904,N_24500);
nand UO_682 (O_682,N_24848,N_24483);
nor UO_683 (O_683,N_24622,N_24878);
or UO_684 (O_684,N_24645,N_24971);
xor UO_685 (O_685,N_24849,N_24489);
and UO_686 (O_686,N_24702,N_24479);
or UO_687 (O_687,N_24390,N_24421);
nor UO_688 (O_688,N_24758,N_24656);
nand UO_689 (O_689,N_24862,N_24905);
or UO_690 (O_690,N_24814,N_24429);
xnor UO_691 (O_691,N_24770,N_24709);
nor UO_692 (O_692,N_24750,N_24446);
nand UO_693 (O_693,N_24663,N_24532);
xnor UO_694 (O_694,N_24619,N_24988);
or UO_695 (O_695,N_24755,N_24903);
or UO_696 (O_696,N_24693,N_24461);
xor UO_697 (O_697,N_24906,N_24498);
nor UO_698 (O_698,N_24994,N_24934);
and UO_699 (O_699,N_24761,N_24392);
or UO_700 (O_700,N_24377,N_24802);
nor UO_701 (O_701,N_24764,N_24683);
and UO_702 (O_702,N_24872,N_24655);
nor UO_703 (O_703,N_24748,N_24786);
or UO_704 (O_704,N_24799,N_24757);
or UO_705 (O_705,N_24697,N_24711);
or UO_706 (O_706,N_24746,N_24995);
and UO_707 (O_707,N_24520,N_24735);
or UO_708 (O_708,N_24482,N_24908);
or UO_709 (O_709,N_24991,N_24958);
and UO_710 (O_710,N_24489,N_24456);
nand UO_711 (O_711,N_24889,N_24483);
or UO_712 (O_712,N_24405,N_24942);
and UO_713 (O_713,N_24647,N_24710);
nor UO_714 (O_714,N_24555,N_24409);
nor UO_715 (O_715,N_24621,N_24613);
nand UO_716 (O_716,N_24415,N_24567);
nand UO_717 (O_717,N_24956,N_24411);
or UO_718 (O_718,N_24847,N_24524);
nor UO_719 (O_719,N_24798,N_24493);
xor UO_720 (O_720,N_24902,N_24412);
and UO_721 (O_721,N_24661,N_24972);
nand UO_722 (O_722,N_24529,N_24803);
or UO_723 (O_723,N_24635,N_24600);
and UO_724 (O_724,N_24593,N_24394);
nor UO_725 (O_725,N_24500,N_24822);
nor UO_726 (O_726,N_24820,N_24599);
nand UO_727 (O_727,N_24430,N_24872);
and UO_728 (O_728,N_24985,N_24686);
or UO_729 (O_729,N_24631,N_24522);
or UO_730 (O_730,N_24482,N_24527);
nand UO_731 (O_731,N_24938,N_24561);
nor UO_732 (O_732,N_24834,N_24787);
and UO_733 (O_733,N_24892,N_24963);
xnor UO_734 (O_734,N_24866,N_24894);
nor UO_735 (O_735,N_24744,N_24492);
nor UO_736 (O_736,N_24676,N_24821);
nand UO_737 (O_737,N_24812,N_24761);
nand UO_738 (O_738,N_24607,N_24838);
nor UO_739 (O_739,N_24768,N_24923);
or UO_740 (O_740,N_24606,N_24874);
nand UO_741 (O_741,N_24448,N_24924);
nor UO_742 (O_742,N_24567,N_24408);
or UO_743 (O_743,N_24643,N_24430);
and UO_744 (O_744,N_24702,N_24377);
nand UO_745 (O_745,N_24383,N_24839);
or UO_746 (O_746,N_24940,N_24630);
and UO_747 (O_747,N_24557,N_24596);
nand UO_748 (O_748,N_24578,N_24438);
and UO_749 (O_749,N_24959,N_24937);
and UO_750 (O_750,N_24702,N_24527);
and UO_751 (O_751,N_24946,N_24839);
and UO_752 (O_752,N_24887,N_24390);
xor UO_753 (O_753,N_24565,N_24944);
and UO_754 (O_754,N_24747,N_24592);
xnor UO_755 (O_755,N_24876,N_24822);
or UO_756 (O_756,N_24838,N_24970);
and UO_757 (O_757,N_24865,N_24625);
or UO_758 (O_758,N_24554,N_24785);
nor UO_759 (O_759,N_24869,N_24533);
and UO_760 (O_760,N_24875,N_24445);
or UO_761 (O_761,N_24757,N_24505);
nand UO_762 (O_762,N_24408,N_24951);
or UO_763 (O_763,N_24991,N_24500);
nor UO_764 (O_764,N_24415,N_24387);
nand UO_765 (O_765,N_24399,N_24956);
nor UO_766 (O_766,N_24378,N_24625);
and UO_767 (O_767,N_24449,N_24803);
and UO_768 (O_768,N_24853,N_24896);
nor UO_769 (O_769,N_24691,N_24772);
and UO_770 (O_770,N_24757,N_24584);
or UO_771 (O_771,N_24585,N_24489);
or UO_772 (O_772,N_24968,N_24489);
or UO_773 (O_773,N_24684,N_24536);
nand UO_774 (O_774,N_24414,N_24686);
nor UO_775 (O_775,N_24859,N_24603);
or UO_776 (O_776,N_24549,N_24473);
and UO_777 (O_777,N_24455,N_24836);
xor UO_778 (O_778,N_24535,N_24805);
nand UO_779 (O_779,N_24527,N_24778);
or UO_780 (O_780,N_24966,N_24825);
nand UO_781 (O_781,N_24510,N_24636);
or UO_782 (O_782,N_24624,N_24701);
xor UO_783 (O_783,N_24720,N_24780);
nor UO_784 (O_784,N_24900,N_24948);
xnor UO_785 (O_785,N_24775,N_24976);
nand UO_786 (O_786,N_24644,N_24583);
and UO_787 (O_787,N_24830,N_24605);
nand UO_788 (O_788,N_24419,N_24498);
and UO_789 (O_789,N_24908,N_24623);
nor UO_790 (O_790,N_24421,N_24656);
or UO_791 (O_791,N_24442,N_24702);
nand UO_792 (O_792,N_24593,N_24877);
nand UO_793 (O_793,N_24841,N_24496);
xnor UO_794 (O_794,N_24588,N_24439);
xnor UO_795 (O_795,N_24702,N_24545);
and UO_796 (O_796,N_24688,N_24752);
nand UO_797 (O_797,N_24419,N_24425);
or UO_798 (O_798,N_24641,N_24398);
nor UO_799 (O_799,N_24415,N_24544);
or UO_800 (O_800,N_24863,N_24600);
nand UO_801 (O_801,N_24562,N_24500);
nand UO_802 (O_802,N_24480,N_24529);
nor UO_803 (O_803,N_24695,N_24984);
nand UO_804 (O_804,N_24594,N_24632);
xor UO_805 (O_805,N_24932,N_24540);
and UO_806 (O_806,N_24508,N_24928);
nand UO_807 (O_807,N_24912,N_24728);
or UO_808 (O_808,N_24666,N_24523);
nor UO_809 (O_809,N_24621,N_24681);
and UO_810 (O_810,N_24593,N_24540);
and UO_811 (O_811,N_24443,N_24901);
or UO_812 (O_812,N_24680,N_24421);
or UO_813 (O_813,N_24858,N_24648);
nand UO_814 (O_814,N_24450,N_24995);
or UO_815 (O_815,N_24764,N_24981);
and UO_816 (O_816,N_24409,N_24720);
nor UO_817 (O_817,N_24956,N_24850);
xnor UO_818 (O_818,N_24648,N_24736);
and UO_819 (O_819,N_24969,N_24863);
or UO_820 (O_820,N_24701,N_24559);
and UO_821 (O_821,N_24485,N_24763);
and UO_822 (O_822,N_24919,N_24878);
nor UO_823 (O_823,N_24591,N_24747);
and UO_824 (O_824,N_24640,N_24482);
and UO_825 (O_825,N_24779,N_24668);
nor UO_826 (O_826,N_24775,N_24815);
nand UO_827 (O_827,N_24385,N_24647);
nand UO_828 (O_828,N_24966,N_24620);
nand UO_829 (O_829,N_24600,N_24575);
nor UO_830 (O_830,N_24707,N_24738);
and UO_831 (O_831,N_24446,N_24719);
nor UO_832 (O_832,N_24494,N_24945);
nand UO_833 (O_833,N_24672,N_24574);
nand UO_834 (O_834,N_24708,N_24733);
nor UO_835 (O_835,N_24653,N_24926);
nor UO_836 (O_836,N_24767,N_24709);
and UO_837 (O_837,N_24705,N_24991);
nor UO_838 (O_838,N_24705,N_24489);
nand UO_839 (O_839,N_24549,N_24850);
or UO_840 (O_840,N_24650,N_24685);
xnor UO_841 (O_841,N_24389,N_24715);
and UO_842 (O_842,N_24937,N_24574);
nand UO_843 (O_843,N_24716,N_24775);
and UO_844 (O_844,N_24989,N_24463);
nor UO_845 (O_845,N_24734,N_24421);
nor UO_846 (O_846,N_24603,N_24814);
and UO_847 (O_847,N_24739,N_24844);
nor UO_848 (O_848,N_24506,N_24440);
xor UO_849 (O_849,N_24891,N_24959);
nand UO_850 (O_850,N_24506,N_24830);
nor UO_851 (O_851,N_24998,N_24405);
nand UO_852 (O_852,N_24552,N_24640);
or UO_853 (O_853,N_24751,N_24942);
xnor UO_854 (O_854,N_24509,N_24525);
or UO_855 (O_855,N_24919,N_24913);
xnor UO_856 (O_856,N_24871,N_24533);
or UO_857 (O_857,N_24466,N_24842);
and UO_858 (O_858,N_24684,N_24749);
and UO_859 (O_859,N_24630,N_24735);
nor UO_860 (O_860,N_24708,N_24521);
and UO_861 (O_861,N_24482,N_24838);
nor UO_862 (O_862,N_24953,N_24485);
or UO_863 (O_863,N_24974,N_24626);
or UO_864 (O_864,N_24755,N_24586);
and UO_865 (O_865,N_24807,N_24605);
nand UO_866 (O_866,N_24852,N_24998);
nand UO_867 (O_867,N_24737,N_24924);
and UO_868 (O_868,N_24921,N_24575);
or UO_869 (O_869,N_24717,N_24516);
xor UO_870 (O_870,N_24863,N_24686);
or UO_871 (O_871,N_24432,N_24629);
and UO_872 (O_872,N_24750,N_24858);
nand UO_873 (O_873,N_24848,N_24999);
nor UO_874 (O_874,N_24621,N_24652);
or UO_875 (O_875,N_24806,N_24583);
or UO_876 (O_876,N_24557,N_24770);
and UO_877 (O_877,N_24579,N_24627);
and UO_878 (O_878,N_24820,N_24801);
or UO_879 (O_879,N_24921,N_24636);
or UO_880 (O_880,N_24964,N_24543);
nand UO_881 (O_881,N_24972,N_24440);
nor UO_882 (O_882,N_24818,N_24747);
nor UO_883 (O_883,N_24979,N_24414);
nor UO_884 (O_884,N_24841,N_24524);
or UO_885 (O_885,N_24460,N_24975);
nand UO_886 (O_886,N_24874,N_24941);
nand UO_887 (O_887,N_24655,N_24383);
nor UO_888 (O_888,N_24499,N_24757);
or UO_889 (O_889,N_24782,N_24431);
nand UO_890 (O_890,N_24661,N_24925);
nor UO_891 (O_891,N_24526,N_24975);
or UO_892 (O_892,N_24968,N_24389);
nand UO_893 (O_893,N_24488,N_24671);
nand UO_894 (O_894,N_24507,N_24702);
or UO_895 (O_895,N_24884,N_24897);
nor UO_896 (O_896,N_24476,N_24646);
nand UO_897 (O_897,N_24433,N_24413);
nand UO_898 (O_898,N_24589,N_24464);
and UO_899 (O_899,N_24625,N_24935);
and UO_900 (O_900,N_24543,N_24431);
or UO_901 (O_901,N_24501,N_24802);
nand UO_902 (O_902,N_24731,N_24717);
or UO_903 (O_903,N_24508,N_24894);
and UO_904 (O_904,N_24554,N_24583);
or UO_905 (O_905,N_24720,N_24577);
nand UO_906 (O_906,N_24839,N_24693);
and UO_907 (O_907,N_24453,N_24561);
and UO_908 (O_908,N_24751,N_24435);
xnor UO_909 (O_909,N_24476,N_24832);
or UO_910 (O_910,N_24657,N_24804);
and UO_911 (O_911,N_24819,N_24992);
nand UO_912 (O_912,N_24466,N_24987);
or UO_913 (O_913,N_24985,N_24402);
nor UO_914 (O_914,N_24562,N_24938);
nand UO_915 (O_915,N_24622,N_24417);
or UO_916 (O_916,N_24472,N_24744);
nand UO_917 (O_917,N_24916,N_24447);
xnor UO_918 (O_918,N_24714,N_24600);
xnor UO_919 (O_919,N_24638,N_24779);
nand UO_920 (O_920,N_24736,N_24732);
or UO_921 (O_921,N_24743,N_24686);
nand UO_922 (O_922,N_24909,N_24620);
and UO_923 (O_923,N_24549,N_24714);
nand UO_924 (O_924,N_24688,N_24390);
nor UO_925 (O_925,N_24385,N_24669);
xnor UO_926 (O_926,N_24780,N_24452);
nand UO_927 (O_927,N_24547,N_24645);
and UO_928 (O_928,N_24745,N_24823);
or UO_929 (O_929,N_24996,N_24429);
nand UO_930 (O_930,N_24812,N_24689);
or UO_931 (O_931,N_24606,N_24668);
or UO_932 (O_932,N_24389,N_24470);
nand UO_933 (O_933,N_24756,N_24527);
nor UO_934 (O_934,N_24510,N_24678);
xnor UO_935 (O_935,N_24464,N_24748);
and UO_936 (O_936,N_24852,N_24824);
or UO_937 (O_937,N_24639,N_24801);
xnor UO_938 (O_938,N_24870,N_24397);
nand UO_939 (O_939,N_24687,N_24460);
and UO_940 (O_940,N_24789,N_24725);
nand UO_941 (O_941,N_24729,N_24538);
nor UO_942 (O_942,N_24477,N_24963);
or UO_943 (O_943,N_24747,N_24502);
or UO_944 (O_944,N_24539,N_24620);
or UO_945 (O_945,N_24628,N_24852);
and UO_946 (O_946,N_24894,N_24892);
nand UO_947 (O_947,N_24814,N_24834);
nor UO_948 (O_948,N_24757,N_24628);
xnor UO_949 (O_949,N_24745,N_24507);
or UO_950 (O_950,N_24978,N_24729);
and UO_951 (O_951,N_24499,N_24535);
nor UO_952 (O_952,N_24801,N_24586);
xnor UO_953 (O_953,N_24688,N_24796);
and UO_954 (O_954,N_24848,N_24868);
and UO_955 (O_955,N_24767,N_24640);
nand UO_956 (O_956,N_24504,N_24967);
nor UO_957 (O_957,N_24900,N_24985);
or UO_958 (O_958,N_24638,N_24960);
or UO_959 (O_959,N_24720,N_24595);
xnor UO_960 (O_960,N_24707,N_24698);
nor UO_961 (O_961,N_24540,N_24661);
nand UO_962 (O_962,N_24671,N_24840);
nand UO_963 (O_963,N_24951,N_24655);
nor UO_964 (O_964,N_24893,N_24803);
nor UO_965 (O_965,N_24611,N_24653);
or UO_966 (O_966,N_24677,N_24492);
nor UO_967 (O_967,N_24595,N_24881);
nor UO_968 (O_968,N_24408,N_24579);
nand UO_969 (O_969,N_24603,N_24671);
xnor UO_970 (O_970,N_24838,N_24728);
nand UO_971 (O_971,N_24990,N_24939);
nor UO_972 (O_972,N_24616,N_24933);
nand UO_973 (O_973,N_24432,N_24635);
nor UO_974 (O_974,N_24940,N_24392);
or UO_975 (O_975,N_24499,N_24940);
or UO_976 (O_976,N_24383,N_24929);
nor UO_977 (O_977,N_24753,N_24448);
xnor UO_978 (O_978,N_24543,N_24614);
xnor UO_979 (O_979,N_24440,N_24520);
nor UO_980 (O_980,N_24729,N_24713);
and UO_981 (O_981,N_24443,N_24806);
and UO_982 (O_982,N_24676,N_24749);
and UO_983 (O_983,N_24453,N_24526);
nor UO_984 (O_984,N_24566,N_24874);
nand UO_985 (O_985,N_24630,N_24949);
and UO_986 (O_986,N_24679,N_24877);
xnor UO_987 (O_987,N_24696,N_24476);
nand UO_988 (O_988,N_24707,N_24882);
nand UO_989 (O_989,N_24697,N_24666);
and UO_990 (O_990,N_24436,N_24860);
nor UO_991 (O_991,N_24915,N_24793);
nor UO_992 (O_992,N_24711,N_24759);
nor UO_993 (O_993,N_24695,N_24389);
nor UO_994 (O_994,N_24765,N_24578);
nand UO_995 (O_995,N_24911,N_24653);
nand UO_996 (O_996,N_24413,N_24633);
and UO_997 (O_997,N_24888,N_24722);
and UO_998 (O_998,N_24544,N_24924);
and UO_999 (O_999,N_24758,N_24440);
xnor UO_1000 (O_1000,N_24393,N_24448);
nor UO_1001 (O_1001,N_24486,N_24802);
and UO_1002 (O_1002,N_24421,N_24952);
nor UO_1003 (O_1003,N_24467,N_24960);
nor UO_1004 (O_1004,N_24868,N_24438);
or UO_1005 (O_1005,N_24700,N_24811);
and UO_1006 (O_1006,N_24705,N_24801);
nand UO_1007 (O_1007,N_24515,N_24994);
nor UO_1008 (O_1008,N_24717,N_24547);
and UO_1009 (O_1009,N_24743,N_24477);
or UO_1010 (O_1010,N_24548,N_24587);
or UO_1011 (O_1011,N_24736,N_24655);
nand UO_1012 (O_1012,N_24913,N_24628);
and UO_1013 (O_1013,N_24905,N_24454);
or UO_1014 (O_1014,N_24750,N_24407);
xor UO_1015 (O_1015,N_24983,N_24603);
nor UO_1016 (O_1016,N_24560,N_24884);
nor UO_1017 (O_1017,N_24498,N_24504);
and UO_1018 (O_1018,N_24583,N_24688);
or UO_1019 (O_1019,N_24475,N_24410);
or UO_1020 (O_1020,N_24687,N_24774);
xor UO_1021 (O_1021,N_24827,N_24990);
and UO_1022 (O_1022,N_24510,N_24771);
nor UO_1023 (O_1023,N_24957,N_24593);
or UO_1024 (O_1024,N_24995,N_24457);
or UO_1025 (O_1025,N_24966,N_24969);
or UO_1026 (O_1026,N_24433,N_24447);
nand UO_1027 (O_1027,N_24464,N_24786);
nand UO_1028 (O_1028,N_24691,N_24449);
or UO_1029 (O_1029,N_24980,N_24493);
nor UO_1030 (O_1030,N_24389,N_24851);
or UO_1031 (O_1031,N_24583,N_24512);
xor UO_1032 (O_1032,N_24528,N_24739);
nor UO_1033 (O_1033,N_24648,N_24485);
or UO_1034 (O_1034,N_24377,N_24616);
nand UO_1035 (O_1035,N_24757,N_24726);
nor UO_1036 (O_1036,N_24426,N_24525);
and UO_1037 (O_1037,N_24857,N_24868);
or UO_1038 (O_1038,N_24735,N_24750);
and UO_1039 (O_1039,N_24375,N_24673);
nand UO_1040 (O_1040,N_24475,N_24872);
and UO_1041 (O_1041,N_24660,N_24789);
or UO_1042 (O_1042,N_24678,N_24726);
and UO_1043 (O_1043,N_24911,N_24886);
or UO_1044 (O_1044,N_24508,N_24775);
and UO_1045 (O_1045,N_24466,N_24514);
or UO_1046 (O_1046,N_24914,N_24620);
xnor UO_1047 (O_1047,N_24950,N_24730);
xor UO_1048 (O_1048,N_24665,N_24860);
nand UO_1049 (O_1049,N_24918,N_24696);
nor UO_1050 (O_1050,N_24830,N_24613);
or UO_1051 (O_1051,N_24611,N_24603);
nor UO_1052 (O_1052,N_24655,N_24530);
and UO_1053 (O_1053,N_24927,N_24562);
or UO_1054 (O_1054,N_24475,N_24479);
nor UO_1055 (O_1055,N_24590,N_24433);
and UO_1056 (O_1056,N_24377,N_24984);
nand UO_1057 (O_1057,N_24569,N_24913);
nand UO_1058 (O_1058,N_24745,N_24987);
and UO_1059 (O_1059,N_24853,N_24834);
and UO_1060 (O_1060,N_24913,N_24754);
nand UO_1061 (O_1061,N_24830,N_24984);
nor UO_1062 (O_1062,N_24755,N_24398);
and UO_1063 (O_1063,N_24641,N_24662);
nor UO_1064 (O_1064,N_24445,N_24631);
and UO_1065 (O_1065,N_24730,N_24596);
nand UO_1066 (O_1066,N_24588,N_24970);
and UO_1067 (O_1067,N_24572,N_24780);
or UO_1068 (O_1068,N_24915,N_24872);
nor UO_1069 (O_1069,N_24954,N_24666);
and UO_1070 (O_1070,N_24617,N_24691);
and UO_1071 (O_1071,N_24467,N_24638);
xor UO_1072 (O_1072,N_24663,N_24562);
nor UO_1073 (O_1073,N_24384,N_24786);
or UO_1074 (O_1074,N_24508,N_24447);
and UO_1075 (O_1075,N_24377,N_24533);
or UO_1076 (O_1076,N_24793,N_24702);
xnor UO_1077 (O_1077,N_24991,N_24744);
xnor UO_1078 (O_1078,N_24945,N_24382);
and UO_1079 (O_1079,N_24735,N_24578);
and UO_1080 (O_1080,N_24474,N_24941);
nor UO_1081 (O_1081,N_24618,N_24524);
or UO_1082 (O_1082,N_24927,N_24541);
or UO_1083 (O_1083,N_24623,N_24896);
or UO_1084 (O_1084,N_24924,N_24709);
nor UO_1085 (O_1085,N_24871,N_24999);
and UO_1086 (O_1086,N_24868,N_24592);
nand UO_1087 (O_1087,N_24447,N_24840);
nand UO_1088 (O_1088,N_24771,N_24422);
nor UO_1089 (O_1089,N_24423,N_24984);
and UO_1090 (O_1090,N_24611,N_24827);
nand UO_1091 (O_1091,N_24517,N_24428);
and UO_1092 (O_1092,N_24588,N_24915);
and UO_1093 (O_1093,N_24829,N_24437);
and UO_1094 (O_1094,N_24656,N_24603);
and UO_1095 (O_1095,N_24964,N_24456);
and UO_1096 (O_1096,N_24811,N_24843);
or UO_1097 (O_1097,N_24478,N_24971);
nor UO_1098 (O_1098,N_24940,N_24642);
and UO_1099 (O_1099,N_24979,N_24823);
or UO_1100 (O_1100,N_24728,N_24698);
nor UO_1101 (O_1101,N_24889,N_24816);
or UO_1102 (O_1102,N_24839,N_24532);
xnor UO_1103 (O_1103,N_24459,N_24707);
nor UO_1104 (O_1104,N_24901,N_24761);
or UO_1105 (O_1105,N_24390,N_24885);
nand UO_1106 (O_1106,N_24962,N_24398);
nand UO_1107 (O_1107,N_24771,N_24613);
nand UO_1108 (O_1108,N_24454,N_24418);
nor UO_1109 (O_1109,N_24648,N_24953);
or UO_1110 (O_1110,N_24794,N_24976);
or UO_1111 (O_1111,N_24917,N_24784);
and UO_1112 (O_1112,N_24585,N_24519);
and UO_1113 (O_1113,N_24687,N_24759);
xor UO_1114 (O_1114,N_24613,N_24793);
nand UO_1115 (O_1115,N_24490,N_24580);
and UO_1116 (O_1116,N_24415,N_24727);
or UO_1117 (O_1117,N_24677,N_24631);
nand UO_1118 (O_1118,N_24915,N_24653);
nor UO_1119 (O_1119,N_24847,N_24743);
nor UO_1120 (O_1120,N_24630,N_24878);
and UO_1121 (O_1121,N_24539,N_24841);
and UO_1122 (O_1122,N_24998,N_24801);
and UO_1123 (O_1123,N_24759,N_24535);
nand UO_1124 (O_1124,N_24522,N_24756);
or UO_1125 (O_1125,N_24862,N_24420);
nor UO_1126 (O_1126,N_24692,N_24567);
nand UO_1127 (O_1127,N_24895,N_24489);
and UO_1128 (O_1128,N_24768,N_24493);
nand UO_1129 (O_1129,N_24432,N_24854);
nand UO_1130 (O_1130,N_24800,N_24543);
nand UO_1131 (O_1131,N_24743,N_24438);
xor UO_1132 (O_1132,N_24707,N_24514);
xnor UO_1133 (O_1133,N_24762,N_24907);
xor UO_1134 (O_1134,N_24905,N_24726);
and UO_1135 (O_1135,N_24643,N_24957);
xor UO_1136 (O_1136,N_24529,N_24783);
nor UO_1137 (O_1137,N_24397,N_24634);
or UO_1138 (O_1138,N_24450,N_24644);
nand UO_1139 (O_1139,N_24401,N_24917);
and UO_1140 (O_1140,N_24376,N_24757);
nand UO_1141 (O_1141,N_24605,N_24715);
xor UO_1142 (O_1142,N_24949,N_24521);
or UO_1143 (O_1143,N_24936,N_24590);
or UO_1144 (O_1144,N_24983,N_24784);
and UO_1145 (O_1145,N_24611,N_24786);
or UO_1146 (O_1146,N_24946,N_24818);
nor UO_1147 (O_1147,N_24725,N_24567);
and UO_1148 (O_1148,N_24999,N_24602);
nor UO_1149 (O_1149,N_24791,N_24483);
nand UO_1150 (O_1150,N_24850,N_24838);
or UO_1151 (O_1151,N_24673,N_24574);
nor UO_1152 (O_1152,N_24856,N_24583);
or UO_1153 (O_1153,N_24971,N_24454);
nand UO_1154 (O_1154,N_24896,N_24391);
nand UO_1155 (O_1155,N_24494,N_24683);
or UO_1156 (O_1156,N_24690,N_24701);
and UO_1157 (O_1157,N_24459,N_24908);
nor UO_1158 (O_1158,N_24990,N_24459);
or UO_1159 (O_1159,N_24661,N_24597);
nor UO_1160 (O_1160,N_24398,N_24466);
nor UO_1161 (O_1161,N_24580,N_24675);
nor UO_1162 (O_1162,N_24492,N_24485);
and UO_1163 (O_1163,N_24589,N_24451);
nand UO_1164 (O_1164,N_24614,N_24545);
nand UO_1165 (O_1165,N_24672,N_24757);
or UO_1166 (O_1166,N_24854,N_24549);
and UO_1167 (O_1167,N_24750,N_24543);
nor UO_1168 (O_1168,N_24857,N_24536);
xor UO_1169 (O_1169,N_24865,N_24719);
nand UO_1170 (O_1170,N_24903,N_24972);
xnor UO_1171 (O_1171,N_24647,N_24749);
or UO_1172 (O_1172,N_24463,N_24803);
and UO_1173 (O_1173,N_24471,N_24711);
nand UO_1174 (O_1174,N_24699,N_24887);
nand UO_1175 (O_1175,N_24628,N_24734);
xor UO_1176 (O_1176,N_24859,N_24957);
nor UO_1177 (O_1177,N_24796,N_24995);
nand UO_1178 (O_1178,N_24895,N_24918);
or UO_1179 (O_1179,N_24551,N_24784);
nand UO_1180 (O_1180,N_24401,N_24457);
or UO_1181 (O_1181,N_24406,N_24928);
or UO_1182 (O_1182,N_24958,N_24585);
nor UO_1183 (O_1183,N_24510,N_24855);
nor UO_1184 (O_1184,N_24747,N_24772);
nor UO_1185 (O_1185,N_24661,N_24377);
nor UO_1186 (O_1186,N_24790,N_24822);
nand UO_1187 (O_1187,N_24738,N_24580);
or UO_1188 (O_1188,N_24574,N_24634);
nor UO_1189 (O_1189,N_24670,N_24738);
nor UO_1190 (O_1190,N_24379,N_24540);
nand UO_1191 (O_1191,N_24794,N_24739);
or UO_1192 (O_1192,N_24886,N_24464);
nor UO_1193 (O_1193,N_24492,N_24407);
and UO_1194 (O_1194,N_24470,N_24603);
or UO_1195 (O_1195,N_24842,N_24503);
nor UO_1196 (O_1196,N_24691,N_24812);
or UO_1197 (O_1197,N_24681,N_24956);
nor UO_1198 (O_1198,N_24879,N_24695);
and UO_1199 (O_1199,N_24633,N_24881);
or UO_1200 (O_1200,N_24575,N_24876);
nand UO_1201 (O_1201,N_24463,N_24398);
and UO_1202 (O_1202,N_24728,N_24410);
nand UO_1203 (O_1203,N_24750,N_24665);
and UO_1204 (O_1204,N_24376,N_24537);
or UO_1205 (O_1205,N_24448,N_24737);
xnor UO_1206 (O_1206,N_24479,N_24391);
nand UO_1207 (O_1207,N_24646,N_24722);
xor UO_1208 (O_1208,N_24709,N_24549);
nor UO_1209 (O_1209,N_24821,N_24509);
or UO_1210 (O_1210,N_24549,N_24697);
and UO_1211 (O_1211,N_24979,N_24873);
or UO_1212 (O_1212,N_24394,N_24420);
and UO_1213 (O_1213,N_24434,N_24507);
or UO_1214 (O_1214,N_24473,N_24792);
xor UO_1215 (O_1215,N_24965,N_24824);
nor UO_1216 (O_1216,N_24583,N_24627);
or UO_1217 (O_1217,N_24445,N_24837);
nor UO_1218 (O_1218,N_24929,N_24653);
nor UO_1219 (O_1219,N_24711,N_24886);
or UO_1220 (O_1220,N_24510,N_24685);
or UO_1221 (O_1221,N_24678,N_24662);
nand UO_1222 (O_1222,N_24776,N_24606);
nor UO_1223 (O_1223,N_24656,N_24586);
and UO_1224 (O_1224,N_24583,N_24706);
nand UO_1225 (O_1225,N_24983,N_24984);
nor UO_1226 (O_1226,N_24534,N_24864);
or UO_1227 (O_1227,N_24973,N_24876);
or UO_1228 (O_1228,N_24894,N_24840);
or UO_1229 (O_1229,N_24829,N_24379);
nor UO_1230 (O_1230,N_24883,N_24448);
and UO_1231 (O_1231,N_24619,N_24649);
and UO_1232 (O_1232,N_24812,N_24722);
nand UO_1233 (O_1233,N_24861,N_24854);
nand UO_1234 (O_1234,N_24829,N_24780);
and UO_1235 (O_1235,N_24479,N_24866);
nand UO_1236 (O_1236,N_24388,N_24552);
nor UO_1237 (O_1237,N_24494,N_24786);
xnor UO_1238 (O_1238,N_24654,N_24590);
or UO_1239 (O_1239,N_24503,N_24805);
or UO_1240 (O_1240,N_24594,N_24379);
and UO_1241 (O_1241,N_24447,N_24613);
and UO_1242 (O_1242,N_24829,N_24648);
nand UO_1243 (O_1243,N_24884,N_24481);
and UO_1244 (O_1244,N_24507,N_24669);
or UO_1245 (O_1245,N_24638,N_24615);
and UO_1246 (O_1246,N_24455,N_24513);
xnor UO_1247 (O_1247,N_24648,N_24940);
nor UO_1248 (O_1248,N_24479,N_24894);
and UO_1249 (O_1249,N_24938,N_24871);
or UO_1250 (O_1250,N_24503,N_24902);
and UO_1251 (O_1251,N_24381,N_24937);
nand UO_1252 (O_1252,N_24792,N_24571);
or UO_1253 (O_1253,N_24823,N_24536);
and UO_1254 (O_1254,N_24983,N_24379);
xnor UO_1255 (O_1255,N_24980,N_24575);
xor UO_1256 (O_1256,N_24920,N_24538);
or UO_1257 (O_1257,N_24467,N_24499);
nand UO_1258 (O_1258,N_24651,N_24548);
or UO_1259 (O_1259,N_24469,N_24774);
or UO_1260 (O_1260,N_24445,N_24583);
or UO_1261 (O_1261,N_24782,N_24515);
and UO_1262 (O_1262,N_24490,N_24600);
and UO_1263 (O_1263,N_24742,N_24952);
or UO_1264 (O_1264,N_24735,N_24452);
xnor UO_1265 (O_1265,N_24727,N_24500);
nand UO_1266 (O_1266,N_24407,N_24926);
and UO_1267 (O_1267,N_24565,N_24504);
nand UO_1268 (O_1268,N_24516,N_24820);
and UO_1269 (O_1269,N_24608,N_24423);
xnor UO_1270 (O_1270,N_24830,N_24831);
nor UO_1271 (O_1271,N_24873,N_24921);
or UO_1272 (O_1272,N_24406,N_24614);
nor UO_1273 (O_1273,N_24816,N_24983);
nand UO_1274 (O_1274,N_24712,N_24797);
or UO_1275 (O_1275,N_24964,N_24818);
nor UO_1276 (O_1276,N_24510,N_24507);
nand UO_1277 (O_1277,N_24508,N_24925);
nor UO_1278 (O_1278,N_24469,N_24758);
and UO_1279 (O_1279,N_24491,N_24649);
or UO_1280 (O_1280,N_24624,N_24610);
or UO_1281 (O_1281,N_24668,N_24713);
nor UO_1282 (O_1282,N_24725,N_24702);
nand UO_1283 (O_1283,N_24880,N_24994);
xnor UO_1284 (O_1284,N_24656,N_24957);
nand UO_1285 (O_1285,N_24645,N_24595);
nand UO_1286 (O_1286,N_24637,N_24705);
nor UO_1287 (O_1287,N_24627,N_24487);
nand UO_1288 (O_1288,N_24777,N_24536);
or UO_1289 (O_1289,N_24924,N_24990);
and UO_1290 (O_1290,N_24987,N_24746);
nand UO_1291 (O_1291,N_24495,N_24748);
and UO_1292 (O_1292,N_24887,N_24865);
nor UO_1293 (O_1293,N_24642,N_24639);
nor UO_1294 (O_1294,N_24564,N_24622);
and UO_1295 (O_1295,N_24981,N_24678);
and UO_1296 (O_1296,N_24895,N_24488);
nor UO_1297 (O_1297,N_24375,N_24462);
nor UO_1298 (O_1298,N_24568,N_24938);
nand UO_1299 (O_1299,N_24956,N_24553);
or UO_1300 (O_1300,N_24994,N_24906);
or UO_1301 (O_1301,N_24747,N_24949);
xnor UO_1302 (O_1302,N_24779,N_24547);
nor UO_1303 (O_1303,N_24946,N_24598);
nand UO_1304 (O_1304,N_24868,N_24502);
xnor UO_1305 (O_1305,N_24900,N_24896);
nand UO_1306 (O_1306,N_24436,N_24869);
and UO_1307 (O_1307,N_24586,N_24762);
nand UO_1308 (O_1308,N_24669,N_24632);
nor UO_1309 (O_1309,N_24894,N_24891);
nor UO_1310 (O_1310,N_24786,N_24949);
nor UO_1311 (O_1311,N_24490,N_24724);
and UO_1312 (O_1312,N_24532,N_24818);
nand UO_1313 (O_1313,N_24885,N_24420);
nand UO_1314 (O_1314,N_24815,N_24570);
or UO_1315 (O_1315,N_24883,N_24619);
nor UO_1316 (O_1316,N_24802,N_24820);
or UO_1317 (O_1317,N_24477,N_24646);
or UO_1318 (O_1318,N_24949,N_24934);
and UO_1319 (O_1319,N_24709,N_24928);
or UO_1320 (O_1320,N_24389,N_24724);
xnor UO_1321 (O_1321,N_24473,N_24709);
nand UO_1322 (O_1322,N_24780,N_24551);
or UO_1323 (O_1323,N_24890,N_24417);
nand UO_1324 (O_1324,N_24795,N_24749);
or UO_1325 (O_1325,N_24744,N_24532);
nor UO_1326 (O_1326,N_24926,N_24933);
nand UO_1327 (O_1327,N_24768,N_24533);
and UO_1328 (O_1328,N_24840,N_24795);
nor UO_1329 (O_1329,N_24589,N_24507);
nor UO_1330 (O_1330,N_24509,N_24436);
or UO_1331 (O_1331,N_24666,N_24948);
nand UO_1332 (O_1332,N_24730,N_24597);
nand UO_1333 (O_1333,N_24993,N_24814);
nor UO_1334 (O_1334,N_24687,N_24864);
or UO_1335 (O_1335,N_24777,N_24750);
xor UO_1336 (O_1336,N_24848,N_24923);
or UO_1337 (O_1337,N_24954,N_24454);
nand UO_1338 (O_1338,N_24451,N_24706);
and UO_1339 (O_1339,N_24465,N_24997);
or UO_1340 (O_1340,N_24983,N_24769);
nor UO_1341 (O_1341,N_24581,N_24647);
nand UO_1342 (O_1342,N_24847,N_24734);
and UO_1343 (O_1343,N_24825,N_24890);
or UO_1344 (O_1344,N_24549,N_24494);
nand UO_1345 (O_1345,N_24786,N_24824);
nor UO_1346 (O_1346,N_24839,N_24563);
nor UO_1347 (O_1347,N_24791,N_24889);
nand UO_1348 (O_1348,N_24813,N_24751);
nor UO_1349 (O_1349,N_24797,N_24976);
nor UO_1350 (O_1350,N_24794,N_24982);
nor UO_1351 (O_1351,N_24951,N_24702);
and UO_1352 (O_1352,N_24563,N_24825);
and UO_1353 (O_1353,N_24812,N_24501);
nand UO_1354 (O_1354,N_24754,N_24869);
nand UO_1355 (O_1355,N_24801,N_24702);
nand UO_1356 (O_1356,N_24543,N_24479);
and UO_1357 (O_1357,N_24868,N_24801);
and UO_1358 (O_1358,N_24897,N_24467);
or UO_1359 (O_1359,N_24767,N_24759);
nor UO_1360 (O_1360,N_24448,N_24507);
nand UO_1361 (O_1361,N_24622,N_24935);
or UO_1362 (O_1362,N_24445,N_24816);
nor UO_1363 (O_1363,N_24401,N_24800);
nor UO_1364 (O_1364,N_24813,N_24661);
nor UO_1365 (O_1365,N_24896,N_24402);
and UO_1366 (O_1366,N_24753,N_24967);
nand UO_1367 (O_1367,N_24660,N_24902);
nand UO_1368 (O_1368,N_24907,N_24559);
nor UO_1369 (O_1369,N_24463,N_24977);
xor UO_1370 (O_1370,N_24565,N_24626);
nand UO_1371 (O_1371,N_24725,N_24560);
nand UO_1372 (O_1372,N_24694,N_24594);
or UO_1373 (O_1373,N_24460,N_24675);
xor UO_1374 (O_1374,N_24818,N_24376);
and UO_1375 (O_1375,N_24870,N_24824);
and UO_1376 (O_1376,N_24696,N_24887);
or UO_1377 (O_1377,N_24916,N_24875);
and UO_1378 (O_1378,N_24751,N_24656);
xor UO_1379 (O_1379,N_24941,N_24620);
or UO_1380 (O_1380,N_24696,N_24742);
and UO_1381 (O_1381,N_24925,N_24974);
nand UO_1382 (O_1382,N_24829,N_24955);
and UO_1383 (O_1383,N_24585,N_24509);
or UO_1384 (O_1384,N_24929,N_24915);
and UO_1385 (O_1385,N_24574,N_24817);
or UO_1386 (O_1386,N_24765,N_24540);
or UO_1387 (O_1387,N_24691,N_24527);
nor UO_1388 (O_1388,N_24558,N_24539);
xor UO_1389 (O_1389,N_24840,N_24646);
nor UO_1390 (O_1390,N_24903,N_24898);
xnor UO_1391 (O_1391,N_24597,N_24485);
and UO_1392 (O_1392,N_24787,N_24728);
and UO_1393 (O_1393,N_24937,N_24871);
and UO_1394 (O_1394,N_24449,N_24739);
or UO_1395 (O_1395,N_24526,N_24863);
nor UO_1396 (O_1396,N_24847,N_24514);
and UO_1397 (O_1397,N_24478,N_24578);
nor UO_1398 (O_1398,N_24769,N_24840);
or UO_1399 (O_1399,N_24947,N_24743);
nand UO_1400 (O_1400,N_24585,N_24609);
and UO_1401 (O_1401,N_24558,N_24747);
nand UO_1402 (O_1402,N_24896,N_24829);
or UO_1403 (O_1403,N_24381,N_24840);
nor UO_1404 (O_1404,N_24962,N_24819);
and UO_1405 (O_1405,N_24523,N_24548);
nor UO_1406 (O_1406,N_24889,N_24824);
and UO_1407 (O_1407,N_24627,N_24744);
nand UO_1408 (O_1408,N_24534,N_24556);
nor UO_1409 (O_1409,N_24822,N_24808);
nand UO_1410 (O_1410,N_24594,N_24486);
nor UO_1411 (O_1411,N_24899,N_24815);
nand UO_1412 (O_1412,N_24898,N_24459);
and UO_1413 (O_1413,N_24427,N_24764);
and UO_1414 (O_1414,N_24991,N_24383);
or UO_1415 (O_1415,N_24949,N_24390);
nor UO_1416 (O_1416,N_24498,N_24788);
and UO_1417 (O_1417,N_24705,N_24769);
nor UO_1418 (O_1418,N_24806,N_24601);
or UO_1419 (O_1419,N_24773,N_24521);
nor UO_1420 (O_1420,N_24920,N_24829);
or UO_1421 (O_1421,N_24903,N_24699);
nand UO_1422 (O_1422,N_24804,N_24698);
or UO_1423 (O_1423,N_24400,N_24406);
and UO_1424 (O_1424,N_24715,N_24600);
or UO_1425 (O_1425,N_24859,N_24869);
nand UO_1426 (O_1426,N_24705,N_24663);
nor UO_1427 (O_1427,N_24911,N_24907);
nand UO_1428 (O_1428,N_24415,N_24890);
and UO_1429 (O_1429,N_24753,N_24539);
and UO_1430 (O_1430,N_24519,N_24427);
and UO_1431 (O_1431,N_24446,N_24597);
nor UO_1432 (O_1432,N_24675,N_24814);
nor UO_1433 (O_1433,N_24942,N_24764);
and UO_1434 (O_1434,N_24615,N_24495);
and UO_1435 (O_1435,N_24409,N_24631);
nor UO_1436 (O_1436,N_24976,N_24920);
and UO_1437 (O_1437,N_24952,N_24696);
xor UO_1438 (O_1438,N_24405,N_24923);
nand UO_1439 (O_1439,N_24411,N_24990);
nor UO_1440 (O_1440,N_24798,N_24918);
nor UO_1441 (O_1441,N_24668,N_24741);
nand UO_1442 (O_1442,N_24383,N_24482);
nand UO_1443 (O_1443,N_24619,N_24982);
nand UO_1444 (O_1444,N_24848,N_24479);
nor UO_1445 (O_1445,N_24404,N_24671);
xor UO_1446 (O_1446,N_24417,N_24466);
nor UO_1447 (O_1447,N_24441,N_24508);
nand UO_1448 (O_1448,N_24846,N_24474);
or UO_1449 (O_1449,N_24621,N_24917);
xnor UO_1450 (O_1450,N_24641,N_24975);
nand UO_1451 (O_1451,N_24545,N_24775);
and UO_1452 (O_1452,N_24606,N_24515);
nand UO_1453 (O_1453,N_24378,N_24918);
nand UO_1454 (O_1454,N_24881,N_24828);
nand UO_1455 (O_1455,N_24761,N_24756);
and UO_1456 (O_1456,N_24412,N_24581);
or UO_1457 (O_1457,N_24647,N_24784);
and UO_1458 (O_1458,N_24885,N_24449);
nand UO_1459 (O_1459,N_24544,N_24815);
or UO_1460 (O_1460,N_24781,N_24738);
and UO_1461 (O_1461,N_24422,N_24577);
or UO_1462 (O_1462,N_24698,N_24775);
nor UO_1463 (O_1463,N_24787,N_24596);
nor UO_1464 (O_1464,N_24457,N_24952);
and UO_1465 (O_1465,N_24604,N_24487);
or UO_1466 (O_1466,N_24983,N_24609);
xor UO_1467 (O_1467,N_24910,N_24921);
or UO_1468 (O_1468,N_24918,N_24780);
nor UO_1469 (O_1469,N_24402,N_24393);
or UO_1470 (O_1470,N_24720,N_24534);
nand UO_1471 (O_1471,N_24798,N_24896);
and UO_1472 (O_1472,N_24727,N_24977);
or UO_1473 (O_1473,N_24624,N_24721);
and UO_1474 (O_1474,N_24629,N_24763);
or UO_1475 (O_1475,N_24754,N_24789);
and UO_1476 (O_1476,N_24913,N_24581);
or UO_1477 (O_1477,N_24630,N_24505);
xnor UO_1478 (O_1478,N_24533,N_24544);
xor UO_1479 (O_1479,N_24999,N_24886);
nand UO_1480 (O_1480,N_24770,N_24649);
nor UO_1481 (O_1481,N_24932,N_24555);
or UO_1482 (O_1482,N_24880,N_24721);
and UO_1483 (O_1483,N_24628,N_24873);
or UO_1484 (O_1484,N_24742,N_24947);
and UO_1485 (O_1485,N_24932,N_24773);
or UO_1486 (O_1486,N_24954,N_24759);
nor UO_1487 (O_1487,N_24576,N_24810);
and UO_1488 (O_1488,N_24991,N_24743);
nor UO_1489 (O_1489,N_24995,N_24941);
or UO_1490 (O_1490,N_24866,N_24694);
xor UO_1491 (O_1491,N_24410,N_24734);
nor UO_1492 (O_1492,N_24826,N_24539);
nor UO_1493 (O_1493,N_24736,N_24414);
nand UO_1494 (O_1494,N_24765,N_24453);
and UO_1495 (O_1495,N_24479,N_24567);
nand UO_1496 (O_1496,N_24726,N_24743);
or UO_1497 (O_1497,N_24738,N_24865);
nand UO_1498 (O_1498,N_24786,N_24863);
or UO_1499 (O_1499,N_24790,N_24843);
xor UO_1500 (O_1500,N_24849,N_24576);
nand UO_1501 (O_1501,N_24605,N_24877);
or UO_1502 (O_1502,N_24762,N_24621);
nand UO_1503 (O_1503,N_24802,N_24590);
nand UO_1504 (O_1504,N_24872,N_24546);
nor UO_1505 (O_1505,N_24994,N_24403);
nor UO_1506 (O_1506,N_24389,N_24940);
xor UO_1507 (O_1507,N_24909,N_24538);
or UO_1508 (O_1508,N_24620,N_24631);
and UO_1509 (O_1509,N_24893,N_24866);
nand UO_1510 (O_1510,N_24934,N_24783);
or UO_1511 (O_1511,N_24523,N_24913);
nor UO_1512 (O_1512,N_24905,N_24475);
or UO_1513 (O_1513,N_24805,N_24640);
nand UO_1514 (O_1514,N_24851,N_24675);
nand UO_1515 (O_1515,N_24548,N_24871);
or UO_1516 (O_1516,N_24952,N_24585);
nand UO_1517 (O_1517,N_24459,N_24609);
or UO_1518 (O_1518,N_24667,N_24801);
nand UO_1519 (O_1519,N_24678,N_24918);
nand UO_1520 (O_1520,N_24817,N_24981);
nor UO_1521 (O_1521,N_24562,N_24983);
and UO_1522 (O_1522,N_24919,N_24439);
nor UO_1523 (O_1523,N_24752,N_24920);
nand UO_1524 (O_1524,N_24812,N_24921);
nor UO_1525 (O_1525,N_24689,N_24757);
xnor UO_1526 (O_1526,N_24787,N_24721);
xnor UO_1527 (O_1527,N_24716,N_24504);
nor UO_1528 (O_1528,N_24488,N_24918);
nand UO_1529 (O_1529,N_24995,N_24627);
and UO_1530 (O_1530,N_24500,N_24555);
or UO_1531 (O_1531,N_24812,N_24380);
nor UO_1532 (O_1532,N_24668,N_24631);
and UO_1533 (O_1533,N_24450,N_24435);
or UO_1534 (O_1534,N_24467,N_24828);
nand UO_1535 (O_1535,N_24775,N_24462);
and UO_1536 (O_1536,N_24848,N_24668);
nor UO_1537 (O_1537,N_24974,N_24971);
xnor UO_1538 (O_1538,N_24918,N_24598);
and UO_1539 (O_1539,N_24934,N_24965);
or UO_1540 (O_1540,N_24892,N_24886);
and UO_1541 (O_1541,N_24999,N_24663);
xnor UO_1542 (O_1542,N_24434,N_24820);
and UO_1543 (O_1543,N_24589,N_24880);
and UO_1544 (O_1544,N_24977,N_24740);
nor UO_1545 (O_1545,N_24589,N_24932);
nor UO_1546 (O_1546,N_24813,N_24392);
nand UO_1547 (O_1547,N_24857,N_24596);
nand UO_1548 (O_1548,N_24745,N_24486);
or UO_1549 (O_1549,N_24502,N_24500);
nand UO_1550 (O_1550,N_24415,N_24568);
and UO_1551 (O_1551,N_24723,N_24585);
xnor UO_1552 (O_1552,N_24758,N_24507);
or UO_1553 (O_1553,N_24408,N_24788);
nor UO_1554 (O_1554,N_24958,N_24541);
nand UO_1555 (O_1555,N_24728,N_24784);
nor UO_1556 (O_1556,N_24831,N_24778);
and UO_1557 (O_1557,N_24483,N_24492);
or UO_1558 (O_1558,N_24648,N_24589);
or UO_1559 (O_1559,N_24608,N_24714);
xnor UO_1560 (O_1560,N_24572,N_24431);
xnor UO_1561 (O_1561,N_24483,N_24530);
nor UO_1562 (O_1562,N_24778,N_24430);
and UO_1563 (O_1563,N_24615,N_24598);
and UO_1564 (O_1564,N_24551,N_24566);
or UO_1565 (O_1565,N_24937,N_24405);
nor UO_1566 (O_1566,N_24947,N_24629);
and UO_1567 (O_1567,N_24645,N_24447);
and UO_1568 (O_1568,N_24880,N_24460);
and UO_1569 (O_1569,N_24695,N_24489);
and UO_1570 (O_1570,N_24784,N_24547);
nor UO_1571 (O_1571,N_24956,N_24523);
or UO_1572 (O_1572,N_24686,N_24542);
or UO_1573 (O_1573,N_24721,N_24385);
nor UO_1574 (O_1574,N_24900,N_24908);
xor UO_1575 (O_1575,N_24959,N_24916);
or UO_1576 (O_1576,N_24937,N_24925);
nand UO_1577 (O_1577,N_24432,N_24543);
nand UO_1578 (O_1578,N_24778,N_24772);
nor UO_1579 (O_1579,N_24489,N_24910);
xor UO_1580 (O_1580,N_24720,N_24829);
nand UO_1581 (O_1581,N_24375,N_24853);
nand UO_1582 (O_1582,N_24416,N_24833);
or UO_1583 (O_1583,N_24424,N_24600);
nand UO_1584 (O_1584,N_24456,N_24843);
and UO_1585 (O_1585,N_24388,N_24934);
or UO_1586 (O_1586,N_24673,N_24904);
or UO_1587 (O_1587,N_24774,N_24525);
nor UO_1588 (O_1588,N_24472,N_24967);
and UO_1589 (O_1589,N_24402,N_24850);
nor UO_1590 (O_1590,N_24874,N_24869);
nor UO_1591 (O_1591,N_24805,N_24971);
nor UO_1592 (O_1592,N_24635,N_24551);
nor UO_1593 (O_1593,N_24481,N_24702);
and UO_1594 (O_1594,N_24722,N_24616);
and UO_1595 (O_1595,N_24844,N_24389);
and UO_1596 (O_1596,N_24977,N_24670);
or UO_1597 (O_1597,N_24748,N_24597);
nor UO_1598 (O_1598,N_24383,N_24982);
or UO_1599 (O_1599,N_24972,N_24461);
nor UO_1600 (O_1600,N_24931,N_24468);
nor UO_1601 (O_1601,N_24881,N_24546);
nand UO_1602 (O_1602,N_24711,N_24503);
nand UO_1603 (O_1603,N_24983,N_24487);
and UO_1604 (O_1604,N_24928,N_24470);
or UO_1605 (O_1605,N_24750,N_24456);
or UO_1606 (O_1606,N_24943,N_24832);
nand UO_1607 (O_1607,N_24463,N_24522);
nand UO_1608 (O_1608,N_24720,N_24742);
and UO_1609 (O_1609,N_24379,N_24945);
nand UO_1610 (O_1610,N_24449,N_24905);
nor UO_1611 (O_1611,N_24859,N_24823);
nor UO_1612 (O_1612,N_24906,N_24553);
and UO_1613 (O_1613,N_24381,N_24695);
or UO_1614 (O_1614,N_24654,N_24938);
and UO_1615 (O_1615,N_24746,N_24964);
nand UO_1616 (O_1616,N_24687,N_24629);
or UO_1617 (O_1617,N_24427,N_24750);
nand UO_1618 (O_1618,N_24485,N_24904);
nand UO_1619 (O_1619,N_24522,N_24666);
nor UO_1620 (O_1620,N_24435,N_24538);
xnor UO_1621 (O_1621,N_24695,N_24858);
and UO_1622 (O_1622,N_24898,N_24772);
and UO_1623 (O_1623,N_24574,N_24468);
and UO_1624 (O_1624,N_24868,N_24666);
and UO_1625 (O_1625,N_24673,N_24522);
and UO_1626 (O_1626,N_24923,N_24619);
and UO_1627 (O_1627,N_24861,N_24694);
or UO_1628 (O_1628,N_24681,N_24553);
nor UO_1629 (O_1629,N_24834,N_24716);
nand UO_1630 (O_1630,N_24620,N_24827);
or UO_1631 (O_1631,N_24730,N_24460);
and UO_1632 (O_1632,N_24926,N_24711);
and UO_1633 (O_1633,N_24679,N_24453);
nor UO_1634 (O_1634,N_24674,N_24843);
and UO_1635 (O_1635,N_24705,N_24485);
xnor UO_1636 (O_1636,N_24832,N_24418);
or UO_1637 (O_1637,N_24399,N_24972);
nand UO_1638 (O_1638,N_24569,N_24576);
nor UO_1639 (O_1639,N_24982,N_24556);
xor UO_1640 (O_1640,N_24743,N_24996);
and UO_1641 (O_1641,N_24705,N_24858);
xnor UO_1642 (O_1642,N_24939,N_24470);
and UO_1643 (O_1643,N_24828,N_24562);
or UO_1644 (O_1644,N_24696,N_24805);
nor UO_1645 (O_1645,N_24633,N_24523);
nor UO_1646 (O_1646,N_24739,N_24950);
nor UO_1647 (O_1647,N_24912,N_24931);
xnor UO_1648 (O_1648,N_24438,N_24917);
nand UO_1649 (O_1649,N_24419,N_24492);
or UO_1650 (O_1650,N_24979,N_24405);
or UO_1651 (O_1651,N_24765,N_24775);
and UO_1652 (O_1652,N_24627,N_24376);
or UO_1653 (O_1653,N_24405,N_24452);
xor UO_1654 (O_1654,N_24883,N_24938);
and UO_1655 (O_1655,N_24958,N_24559);
nand UO_1656 (O_1656,N_24732,N_24394);
and UO_1657 (O_1657,N_24786,N_24945);
or UO_1658 (O_1658,N_24874,N_24649);
nor UO_1659 (O_1659,N_24949,N_24537);
and UO_1660 (O_1660,N_24819,N_24864);
and UO_1661 (O_1661,N_24884,N_24804);
xnor UO_1662 (O_1662,N_24767,N_24880);
nor UO_1663 (O_1663,N_24822,N_24571);
nor UO_1664 (O_1664,N_24912,N_24510);
nor UO_1665 (O_1665,N_24399,N_24712);
xnor UO_1666 (O_1666,N_24751,N_24862);
nor UO_1667 (O_1667,N_24925,N_24444);
xor UO_1668 (O_1668,N_24402,N_24848);
nand UO_1669 (O_1669,N_24910,N_24863);
nand UO_1670 (O_1670,N_24860,N_24859);
or UO_1671 (O_1671,N_24423,N_24782);
nor UO_1672 (O_1672,N_24955,N_24405);
nor UO_1673 (O_1673,N_24823,N_24837);
or UO_1674 (O_1674,N_24934,N_24986);
nand UO_1675 (O_1675,N_24936,N_24833);
nor UO_1676 (O_1676,N_24507,N_24697);
or UO_1677 (O_1677,N_24375,N_24944);
or UO_1678 (O_1678,N_24893,N_24728);
nor UO_1679 (O_1679,N_24534,N_24958);
nand UO_1680 (O_1680,N_24529,N_24955);
nor UO_1681 (O_1681,N_24443,N_24852);
nor UO_1682 (O_1682,N_24466,N_24676);
or UO_1683 (O_1683,N_24409,N_24960);
nand UO_1684 (O_1684,N_24995,N_24836);
nor UO_1685 (O_1685,N_24867,N_24788);
or UO_1686 (O_1686,N_24423,N_24977);
nor UO_1687 (O_1687,N_24833,N_24669);
xnor UO_1688 (O_1688,N_24402,N_24384);
or UO_1689 (O_1689,N_24719,N_24447);
xor UO_1690 (O_1690,N_24896,N_24729);
and UO_1691 (O_1691,N_24856,N_24687);
nand UO_1692 (O_1692,N_24525,N_24447);
or UO_1693 (O_1693,N_24678,N_24596);
nand UO_1694 (O_1694,N_24734,N_24768);
nor UO_1695 (O_1695,N_24632,N_24670);
nand UO_1696 (O_1696,N_24413,N_24771);
xnor UO_1697 (O_1697,N_24866,N_24640);
nand UO_1698 (O_1698,N_24446,N_24518);
nand UO_1699 (O_1699,N_24408,N_24965);
nand UO_1700 (O_1700,N_24399,N_24442);
nand UO_1701 (O_1701,N_24699,N_24712);
or UO_1702 (O_1702,N_24919,N_24853);
or UO_1703 (O_1703,N_24493,N_24738);
nand UO_1704 (O_1704,N_24565,N_24433);
and UO_1705 (O_1705,N_24943,N_24512);
nand UO_1706 (O_1706,N_24490,N_24770);
nand UO_1707 (O_1707,N_24857,N_24821);
and UO_1708 (O_1708,N_24552,N_24727);
nand UO_1709 (O_1709,N_24462,N_24882);
nand UO_1710 (O_1710,N_24601,N_24385);
or UO_1711 (O_1711,N_24916,N_24921);
and UO_1712 (O_1712,N_24890,N_24612);
nor UO_1713 (O_1713,N_24741,N_24475);
or UO_1714 (O_1714,N_24691,N_24800);
and UO_1715 (O_1715,N_24623,N_24649);
nand UO_1716 (O_1716,N_24999,N_24381);
and UO_1717 (O_1717,N_24991,N_24968);
nand UO_1718 (O_1718,N_24637,N_24415);
and UO_1719 (O_1719,N_24773,N_24949);
xnor UO_1720 (O_1720,N_24608,N_24775);
or UO_1721 (O_1721,N_24912,N_24869);
or UO_1722 (O_1722,N_24431,N_24664);
xnor UO_1723 (O_1723,N_24994,N_24580);
nor UO_1724 (O_1724,N_24818,N_24679);
or UO_1725 (O_1725,N_24756,N_24420);
and UO_1726 (O_1726,N_24938,N_24904);
nor UO_1727 (O_1727,N_24792,N_24865);
nor UO_1728 (O_1728,N_24973,N_24732);
nor UO_1729 (O_1729,N_24904,N_24797);
nor UO_1730 (O_1730,N_24719,N_24559);
or UO_1731 (O_1731,N_24523,N_24431);
nand UO_1732 (O_1732,N_24479,N_24961);
or UO_1733 (O_1733,N_24878,N_24520);
and UO_1734 (O_1734,N_24394,N_24540);
xnor UO_1735 (O_1735,N_24526,N_24855);
nand UO_1736 (O_1736,N_24907,N_24744);
nand UO_1737 (O_1737,N_24861,N_24520);
nand UO_1738 (O_1738,N_24677,N_24464);
nor UO_1739 (O_1739,N_24989,N_24799);
nor UO_1740 (O_1740,N_24853,N_24706);
nand UO_1741 (O_1741,N_24533,N_24856);
nor UO_1742 (O_1742,N_24967,N_24837);
nor UO_1743 (O_1743,N_24729,N_24871);
nor UO_1744 (O_1744,N_24549,N_24752);
or UO_1745 (O_1745,N_24762,N_24536);
and UO_1746 (O_1746,N_24902,N_24908);
nand UO_1747 (O_1747,N_24468,N_24876);
nor UO_1748 (O_1748,N_24531,N_24835);
and UO_1749 (O_1749,N_24702,N_24614);
or UO_1750 (O_1750,N_24495,N_24772);
nand UO_1751 (O_1751,N_24673,N_24678);
nor UO_1752 (O_1752,N_24849,N_24861);
nor UO_1753 (O_1753,N_24708,N_24763);
nand UO_1754 (O_1754,N_24752,N_24578);
or UO_1755 (O_1755,N_24577,N_24811);
or UO_1756 (O_1756,N_24657,N_24400);
nor UO_1757 (O_1757,N_24790,N_24781);
or UO_1758 (O_1758,N_24608,N_24569);
xnor UO_1759 (O_1759,N_24630,N_24832);
nor UO_1760 (O_1760,N_24889,N_24408);
or UO_1761 (O_1761,N_24920,N_24834);
nor UO_1762 (O_1762,N_24468,N_24607);
and UO_1763 (O_1763,N_24484,N_24983);
or UO_1764 (O_1764,N_24528,N_24713);
nand UO_1765 (O_1765,N_24455,N_24905);
and UO_1766 (O_1766,N_24979,N_24860);
or UO_1767 (O_1767,N_24580,N_24839);
xor UO_1768 (O_1768,N_24959,N_24541);
and UO_1769 (O_1769,N_24998,N_24547);
nor UO_1770 (O_1770,N_24782,N_24448);
nor UO_1771 (O_1771,N_24464,N_24927);
nor UO_1772 (O_1772,N_24901,N_24924);
and UO_1773 (O_1773,N_24473,N_24783);
nor UO_1774 (O_1774,N_24733,N_24643);
nor UO_1775 (O_1775,N_24849,N_24442);
and UO_1776 (O_1776,N_24924,N_24618);
or UO_1777 (O_1777,N_24461,N_24454);
or UO_1778 (O_1778,N_24610,N_24732);
or UO_1779 (O_1779,N_24759,N_24417);
nor UO_1780 (O_1780,N_24559,N_24724);
nor UO_1781 (O_1781,N_24710,N_24723);
and UO_1782 (O_1782,N_24620,N_24745);
nand UO_1783 (O_1783,N_24720,N_24941);
or UO_1784 (O_1784,N_24786,N_24550);
xnor UO_1785 (O_1785,N_24741,N_24890);
and UO_1786 (O_1786,N_24903,N_24800);
or UO_1787 (O_1787,N_24816,N_24814);
nand UO_1788 (O_1788,N_24819,N_24507);
nand UO_1789 (O_1789,N_24744,N_24473);
and UO_1790 (O_1790,N_24590,N_24842);
and UO_1791 (O_1791,N_24917,N_24648);
nand UO_1792 (O_1792,N_24805,N_24463);
nor UO_1793 (O_1793,N_24626,N_24951);
xnor UO_1794 (O_1794,N_24445,N_24487);
or UO_1795 (O_1795,N_24720,N_24745);
nand UO_1796 (O_1796,N_24427,N_24592);
and UO_1797 (O_1797,N_24642,N_24984);
nor UO_1798 (O_1798,N_24983,N_24656);
and UO_1799 (O_1799,N_24425,N_24461);
or UO_1800 (O_1800,N_24693,N_24740);
and UO_1801 (O_1801,N_24629,N_24443);
or UO_1802 (O_1802,N_24731,N_24700);
nor UO_1803 (O_1803,N_24712,N_24616);
or UO_1804 (O_1804,N_24745,N_24965);
or UO_1805 (O_1805,N_24751,N_24479);
or UO_1806 (O_1806,N_24756,N_24449);
or UO_1807 (O_1807,N_24791,N_24899);
nand UO_1808 (O_1808,N_24832,N_24525);
nor UO_1809 (O_1809,N_24954,N_24430);
nor UO_1810 (O_1810,N_24533,N_24581);
nor UO_1811 (O_1811,N_24452,N_24442);
nand UO_1812 (O_1812,N_24645,N_24912);
nor UO_1813 (O_1813,N_24759,N_24896);
nor UO_1814 (O_1814,N_24761,N_24782);
and UO_1815 (O_1815,N_24633,N_24498);
nand UO_1816 (O_1816,N_24819,N_24711);
nand UO_1817 (O_1817,N_24455,N_24572);
or UO_1818 (O_1818,N_24854,N_24444);
nand UO_1819 (O_1819,N_24406,N_24428);
and UO_1820 (O_1820,N_24481,N_24989);
nor UO_1821 (O_1821,N_24791,N_24395);
nand UO_1822 (O_1822,N_24392,N_24746);
and UO_1823 (O_1823,N_24747,N_24638);
or UO_1824 (O_1824,N_24505,N_24625);
or UO_1825 (O_1825,N_24397,N_24676);
nand UO_1826 (O_1826,N_24745,N_24592);
nand UO_1827 (O_1827,N_24524,N_24684);
or UO_1828 (O_1828,N_24799,N_24857);
nand UO_1829 (O_1829,N_24688,N_24966);
and UO_1830 (O_1830,N_24618,N_24610);
and UO_1831 (O_1831,N_24679,N_24534);
or UO_1832 (O_1832,N_24613,N_24419);
or UO_1833 (O_1833,N_24672,N_24742);
xor UO_1834 (O_1834,N_24742,N_24429);
or UO_1835 (O_1835,N_24444,N_24537);
nor UO_1836 (O_1836,N_24565,N_24723);
nor UO_1837 (O_1837,N_24758,N_24543);
and UO_1838 (O_1838,N_24418,N_24717);
or UO_1839 (O_1839,N_24456,N_24473);
and UO_1840 (O_1840,N_24858,N_24537);
nand UO_1841 (O_1841,N_24491,N_24691);
and UO_1842 (O_1842,N_24561,N_24446);
nand UO_1843 (O_1843,N_24704,N_24912);
and UO_1844 (O_1844,N_24723,N_24495);
or UO_1845 (O_1845,N_24477,N_24486);
nor UO_1846 (O_1846,N_24776,N_24977);
nand UO_1847 (O_1847,N_24384,N_24732);
nor UO_1848 (O_1848,N_24733,N_24908);
and UO_1849 (O_1849,N_24451,N_24856);
nor UO_1850 (O_1850,N_24435,N_24750);
or UO_1851 (O_1851,N_24678,N_24498);
or UO_1852 (O_1852,N_24596,N_24697);
nor UO_1853 (O_1853,N_24548,N_24563);
or UO_1854 (O_1854,N_24799,N_24995);
nand UO_1855 (O_1855,N_24505,N_24607);
nand UO_1856 (O_1856,N_24916,N_24745);
and UO_1857 (O_1857,N_24869,N_24480);
xnor UO_1858 (O_1858,N_24421,N_24549);
or UO_1859 (O_1859,N_24812,N_24552);
xor UO_1860 (O_1860,N_24477,N_24790);
nor UO_1861 (O_1861,N_24489,N_24928);
or UO_1862 (O_1862,N_24693,N_24745);
nor UO_1863 (O_1863,N_24878,N_24837);
nand UO_1864 (O_1864,N_24591,N_24529);
nand UO_1865 (O_1865,N_24697,N_24584);
nor UO_1866 (O_1866,N_24548,N_24627);
nand UO_1867 (O_1867,N_24585,N_24750);
or UO_1868 (O_1868,N_24920,N_24557);
nor UO_1869 (O_1869,N_24743,N_24582);
nor UO_1870 (O_1870,N_24624,N_24806);
nand UO_1871 (O_1871,N_24750,N_24518);
and UO_1872 (O_1872,N_24703,N_24776);
nor UO_1873 (O_1873,N_24635,N_24721);
nand UO_1874 (O_1874,N_24526,N_24937);
or UO_1875 (O_1875,N_24422,N_24887);
and UO_1876 (O_1876,N_24593,N_24423);
nand UO_1877 (O_1877,N_24453,N_24813);
and UO_1878 (O_1878,N_24751,N_24981);
or UO_1879 (O_1879,N_24795,N_24962);
nand UO_1880 (O_1880,N_24824,N_24812);
nor UO_1881 (O_1881,N_24990,N_24957);
nand UO_1882 (O_1882,N_24392,N_24674);
nand UO_1883 (O_1883,N_24671,N_24796);
and UO_1884 (O_1884,N_24552,N_24980);
nor UO_1885 (O_1885,N_24591,N_24945);
or UO_1886 (O_1886,N_24402,N_24527);
and UO_1887 (O_1887,N_24676,N_24806);
or UO_1888 (O_1888,N_24420,N_24452);
nor UO_1889 (O_1889,N_24410,N_24756);
and UO_1890 (O_1890,N_24586,N_24462);
or UO_1891 (O_1891,N_24638,N_24688);
xnor UO_1892 (O_1892,N_24967,N_24756);
or UO_1893 (O_1893,N_24509,N_24748);
nand UO_1894 (O_1894,N_24701,N_24899);
nand UO_1895 (O_1895,N_24685,N_24547);
or UO_1896 (O_1896,N_24995,N_24553);
and UO_1897 (O_1897,N_24498,N_24620);
or UO_1898 (O_1898,N_24771,N_24566);
or UO_1899 (O_1899,N_24481,N_24433);
nand UO_1900 (O_1900,N_24513,N_24832);
xor UO_1901 (O_1901,N_24385,N_24598);
nand UO_1902 (O_1902,N_24844,N_24914);
nand UO_1903 (O_1903,N_24459,N_24560);
nand UO_1904 (O_1904,N_24973,N_24616);
nor UO_1905 (O_1905,N_24890,N_24452);
or UO_1906 (O_1906,N_24771,N_24391);
nor UO_1907 (O_1907,N_24775,N_24827);
nand UO_1908 (O_1908,N_24707,N_24594);
xnor UO_1909 (O_1909,N_24990,N_24814);
or UO_1910 (O_1910,N_24654,N_24963);
xor UO_1911 (O_1911,N_24512,N_24699);
nor UO_1912 (O_1912,N_24597,N_24876);
nor UO_1913 (O_1913,N_24672,N_24496);
xor UO_1914 (O_1914,N_24794,N_24760);
and UO_1915 (O_1915,N_24926,N_24685);
or UO_1916 (O_1916,N_24933,N_24580);
nor UO_1917 (O_1917,N_24883,N_24772);
or UO_1918 (O_1918,N_24557,N_24491);
nand UO_1919 (O_1919,N_24888,N_24745);
or UO_1920 (O_1920,N_24388,N_24503);
and UO_1921 (O_1921,N_24722,N_24914);
nand UO_1922 (O_1922,N_24913,N_24787);
nand UO_1923 (O_1923,N_24637,N_24612);
and UO_1924 (O_1924,N_24458,N_24598);
or UO_1925 (O_1925,N_24861,N_24447);
and UO_1926 (O_1926,N_24911,N_24970);
nand UO_1927 (O_1927,N_24424,N_24685);
nand UO_1928 (O_1928,N_24620,N_24744);
nor UO_1929 (O_1929,N_24497,N_24828);
nor UO_1930 (O_1930,N_24480,N_24970);
xor UO_1931 (O_1931,N_24706,N_24935);
nand UO_1932 (O_1932,N_24682,N_24597);
nor UO_1933 (O_1933,N_24478,N_24605);
nor UO_1934 (O_1934,N_24566,N_24692);
or UO_1935 (O_1935,N_24564,N_24669);
nor UO_1936 (O_1936,N_24787,N_24844);
nand UO_1937 (O_1937,N_24889,N_24687);
or UO_1938 (O_1938,N_24386,N_24501);
nor UO_1939 (O_1939,N_24793,N_24493);
nand UO_1940 (O_1940,N_24663,N_24831);
and UO_1941 (O_1941,N_24995,N_24501);
or UO_1942 (O_1942,N_24911,N_24731);
nand UO_1943 (O_1943,N_24959,N_24408);
and UO_1944 (O_1944,N_24567,N_24660);
and UO_1945 (O_1945,N_24530,N_24939);
xnor UO_1946 (O_1946,N_24662,N_24504);
or UO_1947 (O_1947,N_24433,N_24442);
nand UO_1948 (O_1948,N_24685,N_24932);
or UO_1949 (O_1949,N_24570,N_24493);
nand UO_1950 (O_1950,N_24823,N_24664);
nor UO_1951 (O_1951,N_24697,N_24629);
nor UO_1952 (O_1952,N_24511,N_24849);
nor UO_1953 (O_1953,N_24475,N_24726);
or UO_1954 (O_1954,N_24582,N_24860);
nor UO_1955 (O_1955,N_24788,N_24774);
nor UO_1956 (O_1956,N_24756,N_24376);
nand UO_1957 (O_1957,N_24517,N_24740);
nand UO_1958 (O_1958,N_24748,N_24376);
or UO_1959 (O_1959,N_24916,N_24435);
and UO_1960 (O_1960,N_24682,N_24890);
nor UO_1961 (O_1961,N_24923,N_24482);
nand UO_1962 (O_1962,N_24446,N_24436);
nor UO_1963 (O_1963,N_24419,N_24701);
nand UO_1964 (O_1964,N_24487,N_24634);
and UO_1965 (O_1965,N_24542,N_24588);
nor UO_1966 (O_1966,N_24659,N_24848);
nor UO_1967 (O_1967,N_24831,N_24839);
xnor UO_1968 (O_1968,N_24639,N_24542);
or UO_1969 (O_1969,N_24888,N_24881);
nand UO_1970 (O_1970,N_24643,N_24857);
xor UO_1971 (O_1971,N_24743,N_24645);
nand UO_1972 (O_1972,N_24632,N_24761);
nor UO_1973 (O_1973,N_24566,N_24593);
nand UO_1974 (O_1974,N_24500,N_24921);
nand UO_1975 (O_1975,N_24388,N_24718);
nand UO_1976 (O_1976,N_24661,N_24782);
or UO_1977 (O_1977,N_24388,N_24804);
nor UO_1978 (O_1978,N_24802,N_24471);
nor UO_1979 (O_1979,N_24768,N_24595);
and UO_1980 (O_1980,N_24906,N_24814);
nor UO_1981 (O_1981,N_24592,N_24771);
nor UO_1982 (O_1982,N_24771,N_24503);
nor UO_1983 (O_1983,N_24863,N_24714);
and UO_1984 (O_1984,N_24434,N_24813);
or UO_1985 (O_1985,N_24785,N_24730);
or UO_1986 (O_1986,N_24963,N_24933);
and UO_1987 (O_1987,N_24951,N_24936);
and UO_1988 (O_1988,N_24703,N_24824);
nand UO_1989 (O_1989,N_24719,N_24561);
or UO_1990 (O_1990,N_24814,N_24379);
nand UO_1991 (O_1991,N_24476,N_24662);
or UO_1992 (O_1992,N_24876,N_24752);
and UO_1993 (O_1993,N_24700,N_24375);
nor UO_1994 (O_1994,N_24621,N_24730);
xor UO_1995 (O_1995,N_24408,N_24575);
or UO_1996 (O_1996,N_24740,N_24380);
and UO_1997 (O_1997,N_24697,N_24734);
xor UO_1998 (O_1998,N_24836,N_24511);
nand UO_1999 (O_1999,N_24536,N_24679);
and UO_2000 (O_2000,N_24494,N_24814);
xnor UO_2001 (O_2001,N_24449,N_24823);
and UO_2002 (O_2002,N_24526,N_24465);
or UO_2003 (O_2003,N_24834,N_24593);
nor UO_2004 (O_2004,N_24769,N_24665);
nand UO_2005 (O_2005,N_24686,N_24546);
or UO_2006 (O_2006,N_24645,N_24911);
nor UO_2007 (O_2007,N_24827,N_24935);
and UO_2008 (O_2008,N_24503,N_24748);
nand UO_2009 (O_2009,N_24970,N_24828);
or UO_2010 (O_2010,N_24464,N_24552);
and UO_2011 (O_2011,N_24389,N_24813);
nor UO_2012 (O_2012,N_24756,N_24432);
nand UO_2013 (O_2013,N_24409,N_24519);
nand UO_2014 (O_2014,N_24375,N_24825);
nand UO_2015 (O_2015,N_24824,N_24466);
or UO_2016 (O_2016,N_24408,N_24762);
or UO_2017 (O_2017,N_24733,N_24982);
and UO_2018 (O_2018,N_24621,N_24386);
nand UO_2019 (O_2019,N_24570,N_24390);
or UO_2020 (O_2020,N_24608,N_24695);
and UO_2021 (O_2021,N_24615,N_24876);
nand UO_2022 (O_2022,N_24505,N_24842);
xnor UO_2023 (O_2023,N_24398,N_24383);
and UO_2024 (O_2024,N_24768,N_24551);
or UO_2025 (O_2025,N_24964,N_24990);
nand UO_2026 (O_2026,N_24613,N_24937);
nand UO_2027 (O_2027,N_24674,N_24690);
nand UO_2028 (O_2028,N_24469,N_24679);
nand UO_2029 (O_2029,N_24878,N_24949);
or UO_2030 (O_2030,N_24394,N_24930);
or UO_2031 (O_2031,N_24590,N_24812);
nor UO_2032 (O_2032,N_24888,N_24954);
or UO_2033 (O_2033,N_24628,N_24872);
nand UO_2034 (O_2034,N_24611,N_24913);
or UO_2035 (O_2035,N_24717,N_24885);
and UO_2036 (O_2036,N_24894,N_24743);
xnor UO_2037 (O_2037,N_24571,N_24827);
and UO_2038 (O_2038,N_24861,N_24518);
nor UO_2039 (O_2039,N_24613,N_24818);
and UO_2040 (O_2040,N_24703,N_24920);
or UO_2041 (O_2041,N_24394,N_24869);
nor UO_2042 (O_2042,N_24455,N_24618);
or UO_2043 (O_2043,N_24537,N_24515);
and UO_2044 (O_2044,N_24724,N_24802);
xnor UO_2045 (O_2045,N_24650,N_24983);
xor UO_2046 (O_2046,N_24777,N_24665);
nor UO_2047 (O_2047,N_24515,N_24656);
nor UO_2048 (O_2048,N_24915,N_24741);
nand UO_2049 (O_2049,N_24678,N_24916);
nor UO_2050 (O_2050,N_24943,N_24908);
nor UO_2051 (O_2051,N_24945,N_24706);
nand UO_2052 (O_2052,N_24854,N_24572);
and UO_2053 (O_2053,N_24810,N_24567);
nor UO_2054 (O_2054,N_24809,N_24995);
nor UO_2055 (O_2055,N_24651,N_24701);
or UO_2056 (O_2056,N_24988,N_24760);
xnor UO_2057 (O_2057,N_24908,N_24657);
nand UO_2058 (O_2058,N_24982,N_24977);
nor UO_2059 (O_2059,N_24893,N_24426);
or UO_2060 (O_2060,N_24435,N_24436);
xnor UO_2061 (O_2061,N_24909,N_24467);
and UO_2062 (O_2062,N_24875,N_24692);
or UO_2063 (O_2063,N_24631,N_24653);
and UO_2064 (O_2064,N_24428,N_24611);
or UO_2065 (O_2065,N_24566,N_24590);
and UO_2066 (O_2066,N_24615,N_24796);
nor UO_2067 (O_2067,N_24948,N_24651);
xnor UO_2068 (O_2068,N_24621,N_24446);
and UO_2069 (O_2069,N_24536,N_24426);
nand UO_2070 (O_2070,N_24709,N_24619);
nor UO_2071 (O_2071,N_24866,N_24700);
or UO_2072 (O_2072,N_24721,N_24440);
nand UO_2073 (O_2073,N_24710,N_24966);
or UO_2074 (O_2074,N_24969,N_24664);
or UO_2075 (O_2075,N_24696,N_24889);
nor UO_2076 (O_2076,N_24733,N_24845);
nand UO_2077 (O_2077,N_24723,N_24376);
nor UO_2078 (O_2078,N_24766,N_24459);
nor UO_2079 (O_2079,N_24580,N_24750);
and UO_2080 (O_2080,N_24648,N_24692);
nor UO_2081 (O_2081,N_24380,N_24855);
nor UO_2082 (O_2082,N_24501,N_24628);
nor UO_2083 (O_2083,N_24804,N_24986);
or UO_2084 (O_2084,N_24991,N_24908);
nand UO_2085 (O_2085,N_24877,N_24872);
and UO_2086 (O_2086,N_24868,N_24981);
or UO_2087 (O_2087,N_24394,N_24959);
or UO_2088 (O_2088,N_24590,N_24747);
xnor UO_2089 (O_2089,N_24535,N_24394);
nand UO_2090 (O_2090,N_24993,N_24765);
or UO_2091 (O_2091,N_24568,N_24975);
or UO_2092 (O_2092,N_24959,N_24855);
or UO_2093 (O_2093,N_24781,N_24959);
and UO_2094 (O_2094,N_24737,N_24415);
or UO_2095 (O_2095,N_24577,N_24726);
or UO_2096 (O_2096,N_24803,N_24798);
or UO_2097 (O_2097,N_24893,N_24465);
and UO_2098 (O_2098,N_24653,N_24437);
nand UO_2099 (O_2099,N_24499,N_24716);
and UO_2100 (O_2100,N_24827,N_24477);
nor UO_2101 (O_2101,N_24864,N_24831);
nand UO_2102 (O_2102,N_24712,N_24488);
nand UO_2103 (O_2103,N_24555,N_24865);
and UO_2104 (O_2104,N_24731,N_24585);
xnor UO_2105 (O_2105,N_24492,N_24733);
xnor UO_2106 (O_2106,N_24692,N_24979);
or UO_2107 (O_2107,N_24630,N_24738);
and UO_2108 (O_2108,N_24872,N_24418);
or UO_2109 (O_2109,N_24676,N_24395);
nor UO_2110 (O_2110,N_24806,N_24841);
nand UO_2111 (O_2111,N_24573,N_24452);
and UO_2112 (O_2112,N_24689,N_24525);
or UO_2113 (O_2113,N_24673,N_24617);
nand UO_2114 (O_2114,N_24710,N_24417);
nand UO_2115 (O_2115,N_24786,N_24585);
xnor UO_2116 (O_2116,N_24534,N_24381);
nand UO_2117 (O_2117,N_24965,N_24513);
and UO_2118 (O_2118,N_24719,N_24708);
and UO_2119 (O_2119,N_24883,N_24389);
nor UO_2120 (O_2120,N_24378,N_24588);
nand UO_2121 (O_2121,N_24867,N_24658);
nor UO_2122 (O_2122,N_24728,N_24779);
or UO_2123 (O_2123,N_24944,N_24575);
nor UO_2124 (O_2124,N_24957,N_24574);
nor UO_2125 (O_2125,N_24948,N_24640);
or UO_2126 (O_2126,N_24732,N_24826);
or UO_2127 (O_2127,N_24899,N_24574);
nor UO_2128 (O_2128,N_24579,N_24805);
nor UO_2129 (O_2129,N_24877,N_24635);
nor UO_2130 (O_2130,N_24761,N_24463);
or UO_2131 (O_2131,N_24698,N_24756);
xor UO_2132 (O_2132,N_24852,N_24844);
or UO_2133 (O_2133,N_24466,N_24596);
nand UO_2134 (O_2134,N_24455,N_24629);
nor UO_2135 (O_2135,N_24387,N_24790);
and UO_2136 (O_2136,N_24974,N_24850);
and UO_2137 (O_2137,N_24467,N_24409);
or UO_2138 (O_2138,N_24577,N_24915);
and UO_2139 (O_2139,N_24826,N_24741);
and UO_2140 (O_2140,N_24894,N_24921);
or UO_2141 (O_2141,N_24651,N_24596);
or UO_2142 (O_2142,N_24497,N_24543);
or UO_2143 (O_2143,N_24988,N_24726);
and UO_2144 (O_2144,N_24922,N_24810);
or UO_2145 (O_2145,N_24380,N_24581);
and UO_2146 (O_2146,N_24428,N_24460);
and UO_2147 (O_2147,N_24608,N_24637);
nor UO_2148 (O_2148,N_24580,N_24668);
nand UO_2149 (O_2149,N_24886,N_24453);
nor UO_2150 (O_2150,N_24840,N_24628);
nor UO_2151 (O_2151,N_24441,N_24583);
nand UO_2152 (O_2152,N_24833,N_24551);
or UO_2153 (O_2153,N_24804,N_24623);
nor UO_2154 (O_2154,N_24880,N_24776);
xnor UO_2155 (O_2155,N_24703,N_24933);
xnor UO_2156 (O_2156,N_24450,N_24947);
or UO_2157 (O_2157,N_24744,N_24401);
and UO_2158 (O_2158,N_24515,N_24712);
nand UO_2159 (O_2159,N_24703,N_24409);
nand UO_2160 (O_2160,N_24751,N_24833);
and UO_2161 (O_2161,N_24748,N_24780);
or UO_2162 (O_2162,N_24586,N_24514);
nand UO_2163 (O_2163,N_24502,N_24728);
xnor UO_2164 (O_2164,N_24826,N_24401);
and UO_2165 (O_2165,N_24748,N_24407);
or UO_2166 (O_2166,N_24845,N_24538);
xor UO_2167 (O_2167,N_24743,N_24895);
nand UO_2168 (O_2168,N_24796,N_24718);
and UO_2169 (O_2169,N_24939,N_24754);
nand UO_2170 (O_2170,N_24897,N_24828);
and UO_2171 (O_2171,N_24456,N_24975);
xnor UO_2172 (O_2172,N_24719,N_24690);
nand UO_2173 (O_2173,N_24549,N_24591);
nor UO_2174 (O_2174,N_24463,N_24728);
nand UO_2175 (O_2175,N_24944,N_24658);
or UO_2176 (O_2176,N_24916,N_24540);
or UO_2177 (O_2177,N_24938,N_24380);
xnor UO_2178 (O_2178,N_24375,N_24829);
xnor UO_2179 (O_2179,N_24536,N_24713);
nand UO_2180 (O_2180,N_24834,N_24678);
and UO_2181 (O_2181,N_24487,N_24951);
and UO_2182 (O_2182,N_24477,N_24623);
and UO_2183 (O_2183,N_24944,N_24878);
nor UO_2184 (O_2184,N_24722,N_24791);
nand UO_2185 (O_2185,N_24578,N_24542);
or UO_2186 (O_2186,N_24533,N_24552);
or UO_2187 (O_2187,N_24754,N_24817);
nand UO_2188 (O_2188,N_24984,N_24609);
xnor UO_2189 (O_2189,N_24491,N_24728);
xor UO_2190 (O_2190,N_24823,N_24483);
nand UO_2191 (O_2191,N_24618,N_24404);
nor UO_2192 (O_2192,N_24553,N_24745);
or UO_2193 (O_2193,N_24758,N_24426);
or UO_2194 (O_2194,N_24851,N_24884);
nand UO_2195 (O_2195,N_24942,N_24540);
or UO_2196 (O_2196,N_24998,N_24759);
nor UO_2197 (O_2197,N_24950,N_24653);
nand UO_2198 (O_2198,N_24835,N_24695);
nor UO_2199 (O_2199,N_24977,N_24750);
nor UO_2200 (O_2200,N_24659,N_24933);
nand UO_2201 (O_2201,N_24920,N_24603);
nor UO_2202 (O_2202,N_24907,N_24608);
nor UO_2203 (O_2203,N_24718,N_24747);
nand UO_2204 (O_2204,N_24422,N_24462);
nand UO_2205 (O_2205,N_24526,N_24805);
or UO_2206 (O_2206,N_24619,N_24504);
nand UO_2207 (O_2207,N_24500,N_24623);
nand UO_2208 (O_2208,N_24792,N_24554);
nor UO_2209 (O_2209,N_24933,N_24704);
nor UO_2210 (O_2210,N_24416,N_24582);
xor UO_2211 (O_2211,N_24800,N_24795);
or UO_2212 (O_2212,N_24799,N_24758);
nand UO_2213 (O_2213,N_24615,N_24731);
xor UO_2214 (O_2214,N_24509,N_24984);
or UO_2215 (O_2215,N_24725,N_24653);
or UO_2216 (O_2216,N_24424,N_24430);
nand UO_2217 (O_2217,N_24613,N_24869);
or UO_2218 (O_2218,N_24809,N_24731);
and UO_2219 (O_2219,N_24774,N_24817);
nor UO_2220 (O_2220,N_24874,N_24604);
xor UO_2221 (O_2221,N_24608,N_24437);
nor UO_2222 (O_2222,N_24582,N_24879);
xor UO_2223 (O_2223,N_24631,N_24834);
and UO_2224 (O_2224,N_24864,N_24402);
and UO_2225 (O_2225,N_24819,N_24455);
nor UO_2226 (O_2226,N_24494,N_24895);
and UO_2227 (O_2227,N_24734,N_24822);
nor UO_2228 (O_2228,N_24727,N_24649);
nand UO_2229 (O_2229,N_24883,N_24689);
and UO_2230 (O_2230,N_24802,N_24980);
nand UO_2231 (O_2231,N_24915,N_24554);
and UO_2232 (O_2232,N_24639,N_24687);
or UO_2233 (O_2233,N_24598,N_24562);
xnor UO_2234 (O_2234,N_24957,N_24589);
nand UO_2235 (O_2235,N_24512,N_24762);
or UO_2236 (O_2236,N_24994,N_24940);
and UO_2237 (O_2237,N_24685,N_24900);
or UO_2238 (O_2238,N_24655,N_24664);
nand UO_2239 (O_2239,N_24727,N_24900);
or UO_2240 (O_2240,N_24997,N_24604);
or UO_2241 (O_2241,N_24539,N_24941);
nand UO_2242 (O_2242,N_24887,N_24702);
and UO_2243 (O_2243,N_24429,N_24660);
nor UO_2244 (O_2244,N_24991,N_24376);
nand UO_2245 (O_2245,N_24812,N_24495);
xor UO_2246 (O_2246,N_24912,N_24913);
nand UO_2247 (O_2247,N_24724,N_24771);
and UO_2248 (O_2248,N_24950,N_24771);
and UO_2249 (O_2249,N_24584,N_24577);
and UO_2250 (O_2250,N_24914,N_24545);
nand UO_2251 (O_2251,N_24481,N_24590);
nand UO_2252 (O_2252,N_24764,N_24818);
and UO_2253 (O_2253,N_24480,N_24757);
and UO_2254 (O_2254,N_24920,N_24497);
xor UO_2255 (O_2255,N_24499,N_24849);
nand UO_2256 (O_2256,N_24516,N_24557);
nand UO_2257 (O_2257,N_24886,N_24956);
or UO_2258 (O_2258,N_24875,N_24441);
or UO_2259 (O_2259,N_24530,N_24725);
or UO_2260 (O_2260,N_24588,N_24676);
and UO_2261 (O_2261,N_24910,N_24833);
nor UO_2262 (O_2262,N_24397,N_24470);
xnor UO_2263 (O_2263,N_24832,N_24409);
or UO_2264 (O_2264,N_24624,N_24962);
xnor UO_2265 (O_2265,N_24523,N_24573);
and UO_2266 (O_2266,N_24805,N_24891);
nand UO_2267 (O_2267,N_24421,N_24875);
xnor UO_2268 (O_2268,N_24906,N_24793);
xor UO_2269 (O_2269,N_24562,N_24532);
or UO_2270 (O_2270,N_24606,N_24580);
or UO_2271 (O_2271,N_24693,N_24379);
or UO_2272 (O_2272,N_24389,N_24642);
nand UO_2273 (O_2273,N_24830,N_24961);
nand UO_2274 (O_2274,N_24376,N_24404);
nor UO_2275 (O_2275,N_24562,N_24525);
nor UO_2276 (O_2276,N_24951,N_24803);
or UO_2277 (O_2277,N_24655,N_24421);
nor UO_2278 (O_2278,N_24563,N_24575);
xnor UO_2279 (O_2279,N_24412,N_24414);
xor UO_2280 (O_2280,N_24533,N_24594);
nor UO_2281 (O_2281,N_24548,N_24398);
nor UO_2282 (O_2282,N_24897,N_24618);
or UO_2283 (O_2283,N_24637,N_24950);
or UO_2284 (O_2284,N_24931,N_24748);
xnor UO_2285 (O_2285,N_24510,N_24585);
nor UO_2286 (O_2286,N_24376,N_24925);
nor UO_2287 (O_2287,N_24802,N_24670);
and UO_2288 (O_2288,N_24924,N_24998);
and UO_2289 (O_2289,N_24613,N_24421);
nor UO_2290 (O_2290,N_24885,N_24608);
nand UO_2291 (O_2291,N_24953,N_24590);
nor UO_2292 (O_2292,N_24787,N_24908);
nor UO_2293 (O_2293,N_24744,N_24437);
nand UO_2294 (O_2294,N_24702,N_24891);
or UO_2295 (O_2295,N_24938,N_24762);
and UO_2296 (O_2296,N_24829,N_24942);
xor UO_2297 (O_2297,N_24934,N_24724);
nand UO_2298 (O_2298,N_24939,N_24562);
nor UO_2299 (O_2299,N_24396,N_24672);
and UO_2300 (O_2300,N_24517,N_24817);
nand UO_2301 (O_2301,N_24716,N_24699);
or UO_2302 (O_2302,N_24896,N_24607);
xnor UO_2303 (O_2303,N_24659,N_24939);
nand UO_2304 (O_2304,N_24493,N_24453);
nor UO_2305 (O_2305,N_24566,N_24612);
nand UO_2306 (O_2306,N_24482,N_24817);
xnor UO_2307 (O_2307,N_24537,N_24390);
nand UO_2308 (O_2308,N_24430,N_24947);
nor UO_2309 (O_2309,N_24648,N_24376);
nand UO_2310 (O_2310,N_24444,N_24576);
nor UO_2311 (O_2311,N_24515,N_24518);
or UO_2312 (O_2312,N_24638,N_24631);
and UO_2313 (O_2313,N_24895,N_24965);
nor UO_2314 (O_2314,N_24811,N_24935);
nand UO_2315 (O_2315,N_24638,N_24998);
or UO_2316 (O_2316,N_24569,N_24807);
or UO_2317 (O_2317,N_24531,N_24383);
nand UO_2318 (O_2318,N_24855,N_24987);
nor UO_2319 (O_2319,N_24489,N_24538);
nand UO_2320 (O_2320,N_24815,N_24933);
nand UO_2321 (O_2321,N_24862,N_24638);
nor UO_2322 (O_2322,N_24789,N_24811);
xnor UO_2323 (O_2323,N_24486,N_24910);
nor UO_2324 (O_2324,N_24486,N_24614);
nor UO_2325 (O_2325,N_24656,N_24594);
nand UO_2326 (O_2326,N_24557,N_24412);
or UO_2327 (O_2327,N_24546,N_24466);
nor UO_2328 (O_2328,N_24472,N_24625);
nor UO_2329 (O_2329,N_24424,N_24614);
nor UO_2330 (O_2330,N_24419,N_24441);
nor UO_2331 (O_2331,N_24385,N_24523);
xnor UO_2332 (O_2332,N_24386,N_24908);
or UO_2333 (O_2333,N_24645,N_24498);
or UO_2334 (O_2334,N_24759,N_24524);
nor UO_2335 (O_2335,N_24837,N_24714);
and UO_2336 (O_2336,N_24438,N_24754);
nor UO_2337 (O_2337,N_24386,N_24871);
nand UO_2338 (O_2338,N_24808,N_24922);
and UO_2339 (O_2339,N_24971,N_24612);
nand UO_2340 (O_2340,N_24573,N_24740);
xnor UO_2341 (O_2341,N_24655,N_24678);
nor UO_2342 (O_2342,N_24605,N_24534);
and UO_2343 (O_2343,N_24816,N_24810);
nor UO_2344 (O_2344,N_24992,N_24781);
nor UO_2345 (O_2345,N_24940,N_24577);
and UO_2346 (O_2346,N_24676,N_24511);
nand UO_2347 (O_2347,N_24729,N_24876);
and UO_2348 (O_2348,N_24791,N_24624);
and UO_2349 (O_2349,N_24579,N_24913);
xnor UO_2350 (O_2350,N_24887,N_24692);
nand UO_2351 (O_2351,N_24640,N_24661);
xnor UO_2352 (O_2352,N_24527,N_24500);
nand UO_2353 (O_2353,N_24718,N_24389);
nor UO_2354 (O_2354,N_24880,N_24917);
and UO_2355 (O_2355,N_24601,N_24988);
nand UO_2356 (O_2356,N_24662,N_24658);
nand UO_2357 (O_2357,N_24881,N_24603);
and UO_2358 (O_2358,N_24700,N_24900);
and UO_2359 (O_2359,N_24984,N_24909);
nor UO_2360 (O_2360,N_24455,N_24461);
or UO_2361 (O_2361,N_24686,N_24872);
and UO_2362 (O_2362,N_24996,N_24599);
and UO_2363 (O_2363,N_24919,N_24976);
nor UO_2364 (O_2364,N_24575,N_24910);
or UO_2365 (O_2365,N_24831,N_24690);
and UO_2366 (O_2366,N_24969,N_24376);
nor UO_2367 (O_2367,N_24616,N_24684);
nand UO_2368 (O_2368,N_24596,N_24728);
nor UO_2369 (O_2369,N_24584,N_24777);
and UO_2370 (O_2370,N_24860,N_24748);
and UO_2371 (O_2371,N_24622,N_24597);
or UO_2372 (O_2372,N_24884,N_24665);
and UO_2373 (O_2373,N_24877,N_24667);
and UO_2374 (O_2374,N_24472,N_24460);
nor UO_2375 (O_2375,N_24398,N_24658);
and UO_2376 (O_2376,N_24520,N_24919);
nand UO_2377 (O_2377,N_24667,N_24698);
nor UO_2378 (O_2378,N_24781,N_24682);
nand UO_2379 (O_2379,N_24655,N_24689);
and UO_2380 (O_2380,N_24648,N_24547);
and UO_2381 (O_2381,N_24782,N_24897);
nor UO_2382 (O_2382,N_24578,N_24780);
nand UO_2383 (O_2383,N_24908,N_24550);
or UO_2384 (O_2384,N_24868,N_24439);
nor UO_2385 (O_2385,N_24612,N_24609);
nand UO_2386 (O_2386,N_24829,N_24934);
nor UO_2387 (O_2387,N_24510,N_24982);
nand UO_2388 (O_2388,N_24973,N_24871);
xnor UO_2389 (O_2389,N_24768,N_24909);
and UO_2390 (O_2390,N_24762,N_24378);
and UO_2391 (O_2391,N_24431,N_24564);
nand UO_2392 (O_2392,N_24464,N_24949);
xnor UO_2393 (O_2393,N_24856,N_24837);
nand UO_2394 (O_2394,N_24975,N_24876);
nand UO_2395 (O_2395,N_24870,N_24546);
or UO_2396 (O_2396,N_24726,N_24812);
nor UO_2397 (O_2397,N_24788,N_24389);
nor UO_2398 (O_2398,N_24854,N_24400);
nand UO_2399 (O_2399,N_24944,N_24449);
and UO_2400 (O_2400,N_24524,N_24621);
or UO_2401 (O_2401,N_24633,N_24955);
nor UO_2402 (O_2402,N_24637,N_24738);
nor UO_2403 (O_2403,N_24789,N_24453);
nor UO_2404 (O_2404,N_24811,N_24852);
nor UO_2405 (O_2405,N_24687,N_24706);
or UO_2406 (O_2406,N_24918,N_24849);
or UO_2407 (O_2407,N_24522,N_24663);
nor UO_2408 (O_2408,N_24472,N_24569);
or UO_2409 (O_2409,N_24481,N_24752);
nor UO_2410 (O_2410,N_24537,N_24604);
xor UO_2411 (O_2411,N_24391,N_24746);
nor UO_2412 (O_2412,N_24954,N_24858);
nor UO_2413 (O_2413,N_24703,N_24473);
nor UO_2414 (O_2414,N_24967,N_24761);
or UO_2415 (O_2415,N_24575,N_24888);
and UO_2416 (O_2416,N_24902,N_24778);
xnor UO_2417 (O_2417,N_24493,N_24776);
or UO_2418 (O_2418,N_24445,N_24566);
and UO_2419 (O_2419,N_24801,N_24970);
or UO_2420 (O_2420,N_24605,N_24563);
nor UO_2421 (O_2421,N_24512,N_24554);
xor UO_2422 (O_2422,N_24952,N_24630);
nor UO_2423 (O_2423,N_24971,N_24547);
and UO_2424 (O_2424,N_24484,N_24666);
nor UO_2425 (O_2425,N_24965,N_24522);
or UO_2426 (O_2426,N_24525,N_24813);
nor UO_2427 (O_2427,N_24588,N_24728);
xnor UO_2428 (O_2428,N_24701,N_24691);
and UO_2429 (O_2429,N_24924,N_24419);
and UO_2430 (O_2430,N_24784,N_24794);
or UO_2431 (O_2431,N_24818,N_24711);
nor UO_2432 (O_2432,N_24669,N_24812);
nor UO_2433 (O_2433,N_24856,N_24893);
nand UO_2434 (O_2434,N_24747,N_24819);
nor UO_2435 (O_2435,N_24429,N_24532);
nand UO_2436 (O_2436,N_24419,N_24685);
and UO_2437 (O_2437,N_24437,N_24673);
nor UO_2438 (O_2438,N_24992,N_24682);
nor UO_2439 (O_2439,N_24760,N_24580);
nand UO_2440 (O_2440,N_24698,N_24557);
and UO_2441 (O_2441,N_24396,N_24945);
or UO_2442 (O_2442,N_24438,N_24567);
nor UO_2443 (O_2443,N_24788,N_24805);
nor UO_2444 (O_2444,N_24435,N_24774);
xor UO_2445 (O_2445,N_24633,N_24497);
or UO_2446 (O_2446,N_24798,N_24955);
xnor UO_2447 (O_2447,N_24932,N_24755);
xnor UO_2448 (O_2448,N_24993,N_24863);
nor UO_2449 (O_2449,N_24931,N_24934);
or UO_2450 (O_2450,N_24491,N_24951);
nand UO_2451 (O_2451,N_24852,N_24682);
nand UO_2452 (O_2452,N_24760,N_24544);
or UO_2453 (O_2453,N_24420,N_24753);
xor UO_2454 (O_2454,N_24612,N_24850);
nor UO_2455 (O_2455,N_24389,N_24531);
nor UO_2456 (O_2456,N_24776,N_24497);
nand UO_2457 (O_2457,N_24545,N_24892);
nor UO_2458 (O_2458,N_24994,N_24707);
xnor UO_2459 (O_2459,N_24512,N_24779);
xnor UO_2460 (O_2460,N_24402,N_24654);
nand UO_2461 (O_2461,N_24741,N_24576);
or UO_2462 (O_2462,N_24689,N_24760);
xor UO_2463 (O_2463,N_24939,N_24743);
or UO_2464 (O_2464,N_24710,N_24879);
or UO_2465 (O_2465,N_24754,N_24781);
and UO_2466 (O_2466,N_24653,N_24773);
nor UO_2467 (O_2467,N_24748,N_24785);
nor UO_2468 (O_2468,N_24678,N_24438);
or UO_2469 (O_2469,N_24875,N_24851);
and UO_2470 (O_2470,N_24781,N_24860);
nor UO_2471 (O_2471,N_24863,N_24925);
or UO_2472 (O_2472,N_24550,N_24442);
xor UO_2473 (O_2473,N_24990,N_24698);
xnor UO_2474 (O_2474,N_24544,N_24944);
nand UO_2475 (O_2475,N_24661,N_24638);
nand UO_2476 (O_2476,N_24896,N_24708);
nand UO_2477 (O_2477,N_24925,N_24920);
and UO_2478 (O_2478,N_24765,N_24479);
or UO_2479 (O_2479,N_24654,N_24472);
and UO_2480 (O_2480,N_24833,N_24424);
nand UO_2481 (O_2481,N_24615,N_24648);
or UO_2482 (O_2482,N_24758,N_24753);
nor UO_2483 (O_2483,N_24710,N_24430);
nor UO_2484 (O_2484,N_24755,N_24480);
nand UO_2485 (O_2485,N_24684,N_24482);
nand UO_2486 (O_2486,N_24505,N_24900);
xor UO_2487 (O_2487,N_24940,N_24916);
or UO_2488 (O_2488,N_24535,N_24645);
or UO_2489 (O_2489,N_24928,N_24604);
nor UO_2490 (O_2490,N_24462,N_24799);
or UO_2491 (O_2491,N_24945,N_24717);
nand UO_2492 (O_2492,N_24608,N_24459);
or UO_2493 (O_2493,N_24958,N_24875);
or UO_2494 (O_2494,N_24769,N_24818);
and UO_2495 (O_2495,N_24884,N_24465);
nand UO_2496 (O_2496,N_24985,N_24904);
and UO_2497 (O_2497,N_24397,N_24417);
nor UO_2498 (O_2498,N_24406,N_24566);
nor UO_2499 (O_2499,N_24955,N_24648);
nor UO_2500 (O_2500,N_24966,N_24697);
and UO_2501 (O_2501,N_24950,N_24984);
or UO_2502 (O_2502,N_24630,N_24902);
nor UO_2503 (O_2503,N_24444,N_24974);
or UO_2504 (O_2504,N_24624,N_24450);
nand UO_2505 (O_2505,N_24661,N_24727);
nor UO_2506 (O_2506,N_24475,N_24938);
nand UO_2507 (O_2507,N_24858,N_24576);
nand UO_2508 (O_2508,N_24701,N_24629);
or UO_2509 (O_2509,N_24541,N_24485);
xnor UO_2510 (O_2510,N_24860,N_24838);
nor UO_2511 (O_2511,N_24908,N_24888);
and UO_2512 (O_2512,N_24411,N_24855);
or UO_2513 (O_2513,N_24431,N_24960);
or UO_2514 (O_2514,N_24836,N_24798);
or UO_2515 (O_2515,N_24995,N_24473);
xnor UO_2516 (O_2516,N_24591,N_24446);
nor UO_2517 (O_2517,N_24865,N_24450);
and UO_2518 (O_2518,N_24655,N_24722);
and UO_2519 (O_2519,N_24488,N_24591);
nand UO_2520 (O_2520,N_24777,N_24465);
or UO_2521 (O_2521,N_24504,N_24533);
or UO_2522 (O_2522,N_24609,N_24397);
nand UO_2523 (O_2523,N_24659,N_24965);
nor UO_2524 (O_2524,N_24998,N_24390);
or UO_2525 (O_2525,N_24402,N_24949);
xnor UO_2526 (O_2526,N_24547,N_24951);
or UO_2527 (O_2527,N_24379,N_24551);
and UO_2528 (O_2528,N_24999,N_24970);
and UO_2529 (O_2529,N_24545,N_24756);
nand UO_2530 (O_2530,N_24713,N_24691);
or UO_2531 (O_2531,N_24619,N_24612);
and UO_2532 (O_2532,N_24766,N_24914);
nand UO_2533 (O_2533,N_24410,N_24792);
and UO_2534 (O_2534,N_24531,N_24698);
and UO_2535 (O_2535,N_24668,N_24440);
nor UO_2536 (O_2536,N_24990,N_24485);
or UO_2537 (O_2537,N_24538,N_24612);
and UO_2538 (O_2538,N_24637,N_24670);
nor UO_2539 (O_2539,N_24722,N_24740);
nor UO_2540 (O_2540,N_24540,N_24611);
or UO_2541 (O_2541,N_24376,N_24432);
nor UO_2542 (O_2542,N_24900,N_24579);
and UO_2543 (O_2543,N_24458,N_24863);
and UO_2544 (O_2544,N_24430,N_24878);
xor UO_2545 (O_2545,N_24959,N_24435);
and UO_2546 (O_2546,N_24470,N_24840);
xnor UO_2547 (O_2547,N_24925,N_24922);
nor UO_2548 (O_2548,N_24519,N_24801);
and UO_2549 (O_2549,N_24488,N_24659);
or UO_2550 (O_2550,N_24927,N_24605);
and UO_2551 (O_2551,N_24675,N_24824);
nand UO_2552 (O_2552,N_24853,N_24418);
nand UO_2553 (O_2553,N_24881,N_24502);
and UO_2554 (O_2554,N_24821,N_24661);
nand UO_2555 (O_2555,N_24577,N_24703);
and UO_2556 (O_2556,N_24723,N_24994);
or UO_2557 (O_2557,N_24488,N_24654);
nor UO_2558 (O_2558,N_24617,N_24743);
nor UO_2559 (O_2559,N_24396,N_24539);
or UO_2560 (O_2560,N_24462,N_24902);
nand UO_2561 (O_2561,N_24926,N_24756);
nand UO_2562 (O_2562,N_24892,N_24526);
xnor UO_2563 (O_2563,N_24829,N_24927);
and UO_2564 (O_2564,N_24544,N_24626);
and UO_2565 (O_2565,N_24980,N_24446);
nand UO_2566 (O_2566,N_24800,N_24410);
nand UO_2567 (O_2567,N_24608,N_24933);
nor UO_2568 (O_2568,N_24822,N_24991);
nand UO_2569 (O_2569,N_24600,N_24534);
xnor UO_2570 (O_2570,N_24633,N_24570);
xor UO_2571 (O_2571,N_24748,N_24704);
and UO_2572 (O_2572,N_24757,N_24997);
nand UO_2573 (O_2573,N_24914,N_24634);
nor UO_2574 (O_2574,N_24584,N_24935);
and UO_2575 (O_2575,N_24485,N_24397);
or UO_2576 (O_2576,N_24763,N_24608);
or UO_2577 (O_2577,N_24855,N_24611);
and UO_2578 (O_2578,N_24847,N_24389);
and UO_2579 (O_2579,N_24920,N_24677);
xnor UO_2580 (O_2580,N_24505,N_24477);
or UO_2581 (O_2581,N_24574,N_24632);
or UO_2582 (O_2582,N_24900,N_24719);
nor UO_2583 (O_2583,N_24818,N_24426);
or UO_2584 (O_2584,N_24670,N_24908);
or UO_2585 (O_2585,N_24559,N_24868);
nand UO_2586 (O_2586,N_24635,N_24970);
nand UO_2587 (O_2587,N_24431,N_24687);
and UO_2588 (O_2588,N_24640,N_24434);
nor UO_2589 (O_2589,N_24475,N_24744);
nor UO_2590 (O_2590,N_24396,N_24886);
nand UO_2591 (O_2591,N_24924,N_24554);
nand UO_2592 (O_2592,N_24850,N_24416);
nor UO_2593 (O_2593,N_24511,N_24543);
and UO_2594 (O_2594,N_24853,N_24536);
xor UO_2595 (O_2595,N_24790,N_24716);
nand UO_2596 (O_2596,N_24811,N_24424);
nor UO_2597 (O_2597,N_24849,N_24859);
and UO_2598 (O_2598,N_24836,N_24606);
nand UO_2599 (O_2599,N_24393,N_24435);
xor UO_2600 (O_2600,N_24931,N_24603);
or UO_2601 (O_2601,N_24834,N_24456);
xor UO_2602 (O_2602,N_24530,N_24985);
nand UO_2603 (O_2603,N_24961,N_24647);
nand UO_2604 (O_2604,N_24780,N_24768);
xnor UO_2605 (O_2605,N_24547,N_24435);
nand UO_2606 (O_2606,N_24660,N_24609);
nand UO_2607 (O_2607,N_24609,N_24826);
or UO_2608 (O_2608,N_24797,N_24941);
and UO_2609 (O_2609,N_24607,N_24397);
and UO_2610 (O_2610,N_24814,N_24715);
or UO_2611 (O_2611,N_24682,N_24451);
xor UO_2612 (O_2612,N_24830,N_24580);
nor UO_2613 (O_2613,N_24908,N_24650);
nand UO_2614 (O_2614,N_24619,N_24524);
nor UO_2615 (O_2615,N_24800,N_24960);
and UO_2616 (O_2616,N_24830,N_24681);
or UO_2617 (O_2617,N_24630,N_24530);
and UO_2618 (O_2618,N_24466,N_24695);
or UO_2619 (O_2619,N_24559,N_24615);
and UO_2620 (O_2620,N_24768,N_24386);
or UO_2621 (O_2621,N_24931,N_24986);
and UO_2622 (O_2622,N_24540,N_24641);
and UO_2623 (O_2623,N_24386,N_24444);
nand UO_2624 (O_2624,N_24693,N_24543);
nand UO_2625 (O_2625,N_24864,N_24830);
xnor UO_2626 (O_2626,N_24395,N_24885);
nor UO_2627 (O_2627,N_24597,N_24483);
and UO_2628 (O_2628,N_24545,N_24509);
or UO_2629 (O_2629,N_24949,N_24433);
and UO_2630 (O_2630,N_24503,N_24653);
and UO_2631 (O_2631,N_24992,N_24669);
and UO_2632 (O_2632,N_24547,N_24786);
xnor UO_2633 (O_2633,N_24614,N_24922);
xor UO_2634 (O_2634,N_24387,N_24997);
xor UO_2635 (O_2635,N_24820,N_24651);
nand UO_2636 (O_2636,N_24524,N_24929);
or UO_2637 (O_2637,N_24471,N_24920);
xor UO_2638 (O_2638,N_24554,N_24827);
or UO_2639 (O_2639,N_24668,N_24697);
nand UO_2640 (O_2640,N_24430,N_24386);
and UO_2641 (O_2641,N_24591,N_24844);
nand UO_2642 (O_2642,N_24747,N_24960);
nand UO_2643 (O_2643,N_24733,N_24650);
nor UO_2644 (O_2644,N_24630,N_24826);
nor UO_2645 (O_2645,N_24682,N_24579);
xor UO_2646 (O_2646,N_24777,N_24874);
or UO_2647 (O_2647,N_24932,N_24568);
and UO_2648 (O_2648,N_24707,N_24780);
or UO_2649 (O_2649,N_24574,N_24812);
nor UO_2650 (O_2650,N_24960,N_24738);
nor UO_2651 (O_2651,N_24528,N_24712);
nand UO_2652 (O_2652,N_24689,N_24458);
nand UO_2653 (O_2653,N_24748,N_24856);
nand UO_2654 (O_2654,N_24425,N_24479);
or UO_2655 (O_2655,N_24872,N_24979);
nor UO_2656 (O_2656,N_24849,N_24649);
or UO_2657 (O_2657,N_24471,N_24497);
nor UO_2658 (O_2658,N_24852,N_24643);
xnor UO_2659 (O_2659,N_24378,N_24463);
or UO_2660 (O_2660,N_24944,N_24907);
nand UO_2661 (O_2661,N_24580,N_24993);
and UO_2662 (O_2662,N_24722,N_24660);
and UO_2663 (O_2663,N_24435,N_24982);
and UO_2664 (O_2664,N_24610,N_24935);
nand UO_2665 (O_2665,N_24506,N_24747);
and UO_2666 (O_2666,N_24967,N_24759);
nand UO_2667 (O_2667,N_24826,N_24452);
nand UO_2668 (O_2668,N_24570,N_24976);
nor UO_2669 (O_2669,N_24668,N_24651);
xnor UO_2670 (O_2670,N_24418,N_24533);
and UO_2671 (O_2671,N_24842,N_24432);
nand UO_2672 (O_2672,N_24419,N_24794);
nor UO_2673 (O_2673,N_24852,N_24483);
and UO_2674 (O_2674,N_24962,N_24458);
nand UO_2675 (O_2675,N_24806,N_24769);
and UO_2676 (O_2676,N_24729,N_24588);
nand UO_2677 (O_2677,N_24410,N_24908);
or UO_2678 (O_2678,N_24615,N_24857);
and UO_2679 (O_2679,N_24950,N_24954);
or UO_2680 (O_2680,N_24634,N_24982);
or UO_2681 (O_2681,N_24747,N_24900);
and UO_2682 (O_2682,N_24997,N_24461);
nor UO_2683 (O_2683,N_24667,N_24962);
nor UO_2684 (O_2684,N_24426,N_24745);
or UO_2685 (O_2685,N_24598,N_24952);
or UO_2686 (O_2686,N_24698,N_24443);
and UO_2687 (O_2687,N_24518,N_24476);
or UO_2688 (O_2688,N_24853,N_24442);
xor UO_2689 (O_2689,N_24614,N_24866);
or UO_2690 (O_2690,N_24610,N_24964);
nor UO_2691 (O_2691,N_24842,N_24383);
and UO_2692 (O_2692,N_24989,N_24822);
or UO_2693 (O_2693,N_24959,N_24813);
nand UO_2694 (O_2694,N_24696,N_24939);
or UO_2695 (O_2695,N_24737,N_24967);
xnor UO_2696 (O_2696,N_24918,N_24511);
nor UO_2697 (O_2697,N_24486,N_24414);
nor UO_2698 (O_2698,N_24698,N_24456);
nand UO_2699 (O_2699,N_24765,N_24791);
and UO_2700 (O_2700,N_24755,N_24879);
xor UO_2701 (O_2701,N_24521,N_24605);
and UO_2702 (O_2702,N_24713,N_24615);
nand UO_2703 (O_2703,N_24966,N_24551);
nand UO_2704 (O_2704,N_24468,N_24612);
and UO_2705 (O_2705,N_24675,N_24710);
nor UO_2706 (O_2706,N_24869,N_24632);
nand UO_2707 (O_2707,N_24423,N_24435);
nor UO_2708 (O_2708,N_24443,N_24929);
or UO_2709 (O_2709,N_24764,N_24794);
or UO_2710 (O_2710,N_24863,N_24966);
and UO_2711 (O_2711,N_24612,N_24990);
nand UO_2712 (O_2712,N_24938,N_24923);
nor UO_2713 (O_2713,N_24720,N_24876);
nor UO_2714 (O_2714,N_24838,N_24693);
and UO_2715 (O_2715,N_24513,N_24857);
and UO_2716 (O_2716,N_24531,N_24867);
nand UO_2717 (O_2717,N_24521,N_24539);
nand UO_2718 (O_2718,N_24388,N_24803);
and UO_2719 (O_2719,N_24980,N_24755);
nor UO_2720 (O_2720,N_24694,N_24702);
nand UO_2721 (O_2721,N_24913,N_24897);
xor UO_2722 (O_2722,N_24908,N_24591);
xor UO_2723 (O_2723,N_24488,N_24619);
xnor UO_2724 (O_2724,N_24571,N_24459);
nor UO_2725 (O_2725,N_24650,N_24464);
nor UO_2726 (O_2726,N_24625,N_24403);
nor UO_2727 (O_2727,N_24646,N_24687);
nand UO_2728 (O_2728,N_24841,N_24434);
nor UO_2729 (O_2729,N_24909,N_24392);
nand UO_2730 (O_2730,N_24810,N_24935);
xor UO_2731 (O_2731,N_24826,N_24807);
nand UO_2732 (O_2732,N_24641,N_24408);
and UO_2733 (O_2733,N_24609,N_24729);
nand UO_2734 (O_2734,N_24846,N_24681);
or UO_2735 (O_2735,N_24677,N_24919);
nand UO_2736 (O_2736,N_24719,N_24399);
or UO_2737 (O_2737,N_24405,N_24970);
nor UO_2738 (O_2738,N_24606,N_24823);
nand UO_2739 (O_2739,N_24844,N_24428);
or UO_2740 (O_2740,N_24729,N_24611);
and UO_2741 (O_2741,N_24903,N_24572);
nor UO_2742 (O_2742,N_24859,N_24468);
xnor UO_2743 (O_2743,N_24832,N_24634);
and UO_2744 (O_2744,N_24776,N_24930);
nor UO_2745 (O_2745,N_24622,N_24854);
nand UO_2746 (O_2746,N_24934,N_24831);
nand UO_2747 (O_2747,N_24441,N_24732);
xor UO_2748 (O_2748,N_24704,N_24706);
nand UO_2749 (O_2749,N_24571,N_24561);
nor UO_2750 (O_2750,N_24800,N_24704);
or UO_2751 (O_2751,N_24379,N_24926);
or UO_2752 (O_2752,N_24819,N_24756);
or UO_2753 (O_2753,N_24389,N_24648);
nor UO_2754 (O_2754,N_24545,N_24921);
and UO_2755 (O_2755,N_24643,N_24485);
nand UO_2756 (O_2756,N_24898,N_24839);
nand UO_2757 (O_2757,N_24447,N_24686);
nand UO_2758 (O_2758,N_24398,N_24689);
nor UO_2759 (O_2759,N_24943,N_24793);
nand UO_2760 (O_2760,N_24520,N_24951);
or UO_2761 (O_2761,N_24979,N_24615);
xnor UO_2762 (O_2762,N_24445,N_24529);
nand UO_2763 (O_2763,N_24761,N_24930);
and UO_2764 (O_2764,N_24473,N_24779);
nor UO_2765 (O_2765,N_24646,N_24753);
and UO_2766 (O_2766,N_24882,N_24460);
or UO_2767 (O_2767,N_24604,N_24711);
nand UO_2768 (O_2768,N_24668,N_24919);
nor UO_2769 (O_2769,N_24402,N_24657);
or UO_2770 (O_2770,N_24974,N_24376);
or UO_2771 (O_2771,N_24667,N_24820);
nand UO_2772 (O_2772,N_24763,N_24436);
nor UO_2773 (O_2773,N_24662,N_24869);
nand UO_2774 (O_2774,N_24946,N_24787);
nor UO_2775 (O_2775,N_24813,N_24419);
xor UO_2776 (O_2776,N_24850,N_24427);
nor UO_2777 (O_2777,N_24589,N_24420);
nor UO_2778 (O_2778,N_24597,N_24674);
nand UO_2779 (O_2779,N_24390,N_24958);
nand UO_2780 (O_2780,N_24934,N_24450);
nor UO_2781 (O_2781,N_24722,N_24522);
nor UO_2782 (O_2782,N_24759,N_24913);
and UO_2783 (O_2783,N_24682,N_24464);
nand UO_2784 (O_2784,N_24633,N_24378);
nor UO_2785 (O_2785,N_24716,N_24946);
or UO_2786 (O_2786,N_24420,N_24387);
nor UO_2787 (O_2787,N_24932,N_24698);
nor UO_2788 (O_2788,N_24861,N_24594);
nor UO_2789 (O_2789,N_24800,N_24757);
nand UO_2790 (O_2790,N_24740,N_24980);
or UO_2791 (O_2791,N_24973,N_24714);
xor UO_2792 (O_2792,N_24469,N_24698);
nand UO_2793 (O_2793,N_24955,N_24689);
and UO_2794 (O_2794,N_24882,N_24381);
nor UO_2795 (O_2795,N_24691,N_24782);
xnor UO_2796 (O_2796,N_24878,N_24710);
or UO_2797 (O_2797,N_24748,N_24391);
nand UO_2798 (O_2798,N_24484,N_24558);
xnor UO_2799 (O_2799,N_24390,N_24845);
xnor UO_2800 (O_2800,N_24848,N_24935);
nand UO_2801 (O_2801,N_24504,N_24599);
or UO_2802 (O_2802,N_24987,N_24801);
nand UO_2803 (O_2803,N_24771,N_24548);
nor UO_2804 (O_2804,N_24538,N_24688);
or UO_2805 (O_2805,N_24989,N_24742);
and UO_2806 (O_2806,N_24561,N_24404);
nand UO_2807 (O_2807,N_24726,N_24638);
nor UO_2808 (O_2808,N_24757,N_24648);
and UO_2809 (O_2809,N_24559,N_24860);
xor UO_2810 (O_2810,N_24983,N_24504);
and UO_2811 (O_2811,N_24999,N_24438);
nand UO_2812 (O_2812,N_24441,N_24769);
or UO_2813 (O_2813,N_24824,N_24566);
nor UO_2814 (O_2814,N_24695,N_24762);
or UO_2815 (O_2815,N_24645,N_24985);
nand UO_2816 (O_2816,N_24898,N_24511);
and UO_2817 (O_2817,N_24599,N_24653);
nor UO_2818 (O_2818,N_24454,N_24906);
and UO_2819 (O_2819,N_24632,N_24599);
or UO_2820 (O_2820,N_24669,N_24806);
nor UO_2821 (O_2821,N_24666,N_24888);
nor UO_2822 (O_2822,N_24622,N_24550);
nor UO_2823 (O_2823,N_24675,N_24408);
or UO_2824 (O_2824,N_24561,N_24506);
nor UO_2825 (O_2825,N_24647,N_24996);
nor UO_2826 (O_2826,N_24752,N_24659);
and UO_2827 (O_2827,N_24898,N_24826);
or UO_2828 (O_2828,N_24728,N_24889);
nor UO_2829 (O_2829,N_24966,N_24730);
or UO_2830 (O_2830,N_24974,N_24898);
and UO_2831 (O_2831,N_24676,N_24833);
nand UO_2832 (O_2832,N_24471,N_24971);
and UO_2833 (O_2833,N_24671,N_24446);
xnor UO_2834 (O_2834,N_24386,N_24966);
nand UO_2835 (O_2835,N_24383,N_24718);
xor UO_2836 (O_2836,N_24458,N_24658);
or UO_2837 (O_2837,N_24850,N_24934);
and UO_2838 (O_2838,N_24998,N_24680);
nor UO_2839 (O_2839,N_24617,N_24778);
nor UO_2840 (O_2840,N_24531,N_24579);
nor UO_2841 (O_2841,N_24386,N_24512);
nand UO_2842 (O_2842,N_24592,N_24581);
nand UO_2843 (O_2843,N_24591,N_24781);
nand UO_2844 (O_2844,N_24835,N_24496);
nor UO_2845 (O_2845,N_24796,N_24788);
nand UO_2846 (O_2846,N_24533,N_24805);
nor UO_2847 (O_2847,N_24561,N_24414);
or UO_2848 (O_2848,N_24635,N_24647);
nand UO_2849 (O_2849,N_24436,N_24904);
nand UO_2850 (O_2850,N_24620,N_24859);
and UO_2851 (O_2851,N_24479,N_24919);
or UO_2852 (O_2852,N_24783,N_24941);
nand UO_2853 (O_2853,N_24437,N_24455);
or UO_2854 (O_2854,N_24721,N_24931);
nor UO_2855 (O_2855,N_24547,N_24746);
nand UO_2856 (O_2856,N_24959,N_24961);
nand UO_2857 (O_2857,N_24933,N_24826);
or UO_2858 (O_2858,N_24977,N_24464);
nor UO_2859 (O_2859,N_24957,N_24531);
nand UO_2860 (O_2860,N_24992,N_24796);
xor UO_2861 (O_2861,N_24688,N_24422);
or UO_2862 (O_2862,N_24577,N_24806);
and UO_2863 (O_2863,N_24775,N_24431);
and UO_2864 (O_2864,N_24394,N_24737);
or UO_2865 (O_2865,N_24819,N_24951);
xor UO_2866 (O_2866,N_24838,N_24495);
nor UO_2867 (O_2867,N_24935,N_24611);
nor UO_2868 (O_2868,N_24907,N_24999);
nand UO_2869 (O_2869,N_24871,N_24398);
or UO_2870 (O_2870,N_24686,N_24656);
nand UO_2871 (O_2871,N_24507,N_24426);
nand UO_2872 (O_2872,N_24451,N_24398);
nand UO_2873 (O_2873,N_24744,N_24537);
or UO_2874 (O_2874,N_24984,N_24580);
or UO_2875 (O_2875,N_24857,N_24843);
nand UO_2876 (O_2876,N_24947,N_24532);
nand UO_2877 (O_2877,N_24411,N_24936);
or UO_2878 (O_2878,N_24730,N_24990);
and UO_2879 (O_2879,N_24377,N_24896);
or UO_2880 (O_2880,N_24604,N_24619);
or UO_2881 (O_2881,N_24869,N_24766);
nand UO_2882 (O_2882,N_24768,N_24453);
xnor UO_2883 (O_2883,N_24634,N_24522);
or UO_2884 (O_2884,N_24830,N_24850);
nor UO_2885 (O_2885,N_24987,N_24936);
nor UO_2886 (O_2886,N_24514,N_24872);
and UO_2887 (O_2887,N_24709,N_24960);
nor UO_2888 (O_2888,N_24695,N_24920);
and UO_2889 (O_2889,N_24513,N_24998);
nor UO_2890 (O_2890,N_24444,N_24706);
or UO_2891 (O_2891,N_24596,N_24956);
xor UO_2892 (O_2892,N_24562,N_24528);
nand UO_2893 (O_2893,N_24428,N_24996);
xnor UO_2894 (O_2894,N_24493,N_24854);
and UO_2895 (O_2895,N_24735,N_24942);
nor UO_2896 (O_2896,N_24925,N_24426);
and UO_2897 (O_2897,N_24602,N_24725);
nand UO_2898 (O_2898,N_24600,N_24646);
or UO_2899 (O_2899,N_24737,N_24412);
and UO_2900 (O_2900,N_24781,N_24592);
or UO_2901 (O_2901,N_24637,N_24702);
nand UO_2902 (O_2902,N_24867,N_24978);
nor UO_2903 (O_2903,N_24873,N_24763);
or UO_2904 (O_2904,N_24964,N_24381);
or UO_2905 (O_2905,N_24944,N_24700);
and UO_2906 (O_2906,N_24622,N_24617);
xor UO_2907 (O_2907,N_24806,N_24700);
or UO_2908 (O_2908,N_24401,N_24989);
xor UO_2909 (O_2909,N_24586,N_24886);
xnor UO_2910 (O_2910,N_24592,N_24792);
nor UO_2911 (O_2911,N_24970,N_24437);
nor UO_2912 (O_2912,N_24506,N_24639);
or UO_2913 (O_2913,N_24690,N_24953);
nand UO_2914 (O_2914,N_24743,N_24379);
nor UO_2915 (O_2915,N_24496,N_24494);
and UO_2916 (O_2916,N_24544,N_24704);
nor UO_2917 (O_2917,N_24996,N_24446);
nand UO_2918 (O_2918,N_24603,N_24456);
and UO_2919 (O_2919,N_24791,N_24879);
nor UO_2920 (O_2920,N_24875,N_24584);
or UO_2921 (O_2921,N_24450,N_24986);
or UO_2922 (O_2922,N_24743,N_24713);
nand UO_2923 (O_2923,N_24999,N_24722);
and UO_2924 (O_2924,N_24695,N_24670);
nand UO_2925 (O_2925,N_24673,N_24447);
and UO_2926 (O_2926,N_24799,N_24898);
and UO_2927 (O_2927,N_24539,N_24912);
xor UO_2928 (O_2928,N_24433,N_24999);
or UO_2929 (O_2929,N_24930,N_24893);
nand UO_2930 (O_2930,N_24744,N_24405);
nor UO_2931 (O_2931,N_24961,N_24993);
nand UO_2932 (O_2932,N_24414,N_24763);
nor UO_2933 (O_2933,N_24720,N_24504);
and UO_2934 (O_2934,N_24496,N_24896);
nor UO_2935 (O_2935,N_24429,N_24893);
or UO_2936 (O_2936,N_24457,N_24602);
nor UO_2937 (O_2937,N_24811,N_24649);
or UO_2938 (O_2938,N_24660,N_24531);
xor UO_2939 (O_2939,N_24894,N_24581);
and UO_2940 (O_2940,N_24513,N_24745);
or UO_2941 (O_2941,N_24797,N_24597);
nor UO_2942 (O_2942,N_24434,N_24997);
nand UO_2943 (O_2943,N_24734,N_24625);
xor UO_2944 (O_2944,N_24404,N_24476);
nor UO_2945 (O_2945,N_24545,N_24860);
nor UO_2946 (O_2946,N_24733,N_24477);
or UO_2947 (O_2947,N_24717,N_24618);
or UO_2948 (O_2948,N_24866,N_24583);
nand UO_2949 (O_2949,N_24905,N_24407);
nand UO_2950 (O_2950,N_24885,N_24433);
nand UO_2951 (O_2951,N_24711,N_24529);
nand UO_2952 (O_2952,N_24962,N_24895);
or UO_2953 (O_2953,N_24735,N_24439);
and UO_2954 (O_2954,N_24646,N_24839);
or UO_2955 (O_2955,N_24542,N_24854);
nor UO_2956 (O_2956,N_24395,N_24652);
and UO_2957 (O_2957,N_24576,N_24931);
nand UO_2958 (O_2958,N_24539,N_24496);
or UO_2959 (O_2959,N_24992,N_24832);
xnor UO_2960 (O_2960,N_24437,N_24746);
and UO_2961 (O_2961,N_24530,N_24772);
or UO_2962 (O_2962,N_24888,N_24956);
nand UO_2963 (O_2963,N_24825,N_24907);
and UO_2964 (O_2964,N_24883,N_24889);
and UO_2965 (O_2965,N_24782,N_24793);
or UO_2966 (O_2966,N_24799,N_24733);
nand UO_2967 (O_2967,N_24551,N_24894);
nand UO_2968 (O_2968,N_24484,N_24431);
nand UO_2969 (O_2969,N_24558,N_24672);
or UO_2970 (O_2970,N_24708,N_24382);
or UO_2971 (O_2971,N_24703,N_24791);
nand UO_2972 (O_2972,N_24888,N_24890);
xor UO_2973 (O_2973,N_24555,N_24519);
and UO_2974 (O_2974,N_24480,N_24672);
nor UO_2975 (O_2975,N_24530,N_24773);
nor UO_2976 (O_2976,N_24759,N_24842);
nor UO_2977 (O_2977,N_24396,N_24811);
nor UO_2978 (O_2978,N_24975,N_24577);
and UO_2979 (O_2979,N_24398,N_24508);
nand UO_2980 (O_2980,N_24637,N_24640);
or UO_2981 (O_2981,N_24998,N_24474);
and UO_2982 (O_2982,N_24502,N_24739);
nor UO_2983 (O_2983,N_24808,N_24900);
nand UO_2984 (O_2984,N_24936,N_24490);
and UO_2985 (O_2985,N_24544,N_24425);
nor UO_2986 (O_2986,N_24560,N_24816);
or UO_2987 (O_2987,N_24397,N_24459);
xnor UO_2988 (O_2988,N_24616,N_24671);
and UO_2989 (O_2989,N_24995,N_24758);
or UO_2990 (O_2990,N_24902,N_24579);
nor UO_2991 (O_2991,N_24644,N_24556);
nand UO_2992 (O_2992,N_24704,N_24962);
and UO_2993 (O_2993,N_24409,N_24427);
nand UO_2994 (O_2994,N_24998,N_24664);
and UO_2995 (O_2995,N_24377,N_24926);
xnor UO_2996 (O_2996,N_24551,N_24642);
nand UO_2997 (O_2997,N_24945,N_24773);
xor UO_2998 (O_2998,N_24770,N_24375);
and UO_2999 (O_2999,N_24440,N_24508);
endmodule