module basic_500_3000_500_60_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_458,In_26);
xnor U1 (N_1,In_360,In_162);
or U2 (N_2,In_386,In_347);
and U3 (N_3,In_95,In_21);
nand U4 (N_4,In_8,In_80);
nor U5 (N_5,In_158,In_471);
nor U6 (N_6,In_277,In_290);
nor U7 (N_7,In_307,In_313);
nand U8 (N_8,In_185,In_165);
nand U9 (N_9,In_73,In_300);
xnor U10 (N_10,In_330,In_480);
xor U11 (N_11,In_303,In_134);
nand U12 (N_12,In_312,In_132);
nand U13 (N_13,In_87,In_44);
nand U14 (N_14,In_208,In_319);
and U15 (N_15,In_262,In_177);
and U16 (N_16,In_12,In_126);
and U17 (N_17,In_127,In_7);
and U18 (N_18,In_389,In_308);
and U19 (N_19,In_199,In_148);
nand U20 (N_20,In_397,In_157);
or U21 (N_21,In_202,In_184);
or U22 (N_22,In_230,In_244);
nor U23 (N_23,In_20,In_10);
nand U24 (N_24,In_451,In_54);
or U25 (N_25,In_197,In_286);
nor U26 (N_26,In_440,In_228);
or U27 (N_27,In_392,In_407);
nor U28 (N_28,In_255,In_142);
nor U29 (N_29,In_324,In_427);
nor U30 (N_30,In_305,In_346);
or U31 (N_31,In_498,In_221);
xor U32 (N_32,In_273,In_193);
nor U33 (N_33,In_376,In_144);
nand U34 (N_34,In_90,In_245);
and U35 (N_35,In_470,In_116);
nor U36 (N_36,In_370,In_355);
or U37 (N_37,In_261,In_188);
nand U38 (N_38,In_117,In_326);
nand U39 (N_39,In_112,In_192);
and U40 (N_40,In_30,In_24);
and U41 (N_41,In_212,In_461);
nand U42 (N_42,In_409,In_491);
nor U43 (N_43,In_110,In_70);
nor U44 (N_44,In_260,In_433);
nor U45 (N_45,In_168,In_11);
and U46 (N_46,In_292,In_466);
nand U47 (N_47,In_129,In_190);
or U48 (N_48,In_425,In_482);
nand U49 (N_49,In_42,In_375);
nand U50 (N_50,In_310,In_85);
nand U51 (N_51,In_53,In_83);
nor U52 (N_52,N_35,In_379);
nor U53 (N_53,In_264,In_374);
and U54 (N_54,N_9,In_69);
nor U55 (N_55,In_422,In_51);
or U56 (N_56,In_338,In_384);
or U57 (N_57,N_14,In_31);
or U58 (N_58,In_497,In_79);
nor U59 (N_59,In_98,In_373);
or U60 (N_60,In_265,In_74);
and U61 (N_61,In_280,In_123);
or U62 (N_62,In_194,In_443);
nor U63 (N_63,N_34,In_234);
nor U64 (N_64,N_28,In_13);
nor U65 (N_65,In_487,In_316);
and U66 (N_66,In_344,In_203);
nand U67 (N_67,N_21,In_249);
nor U68 (N_68,In_325,In_86);
nor U69 (N_69,In_39,N_18);
xor U70 (N_70,N_40,In_89);
nor U71 (N_71,In_459,N_5);
nand U72 (N_72,In_105,In_329);
nor U73 (N_73,In_122,In_315);
nand U74 (N_74,In_258,In_195);
and U75 (N_75,In_267,In_309);
nor U76 (N_76,N_17,In_170);
nand U77 (N_77,In_299,In_27);
nand U78 (N_78,In_334,In_133);
nor U79 (N_79,In_223,In_76);
nor U80 (N_80,In_320,In_270);
and U81 (N_81,In_108,N_4);
nand U82 (N_82,In_363,In_456);
nor U83 (N_83,In_17,In_484);
and U84 (N_84,In_57,In_455);
nor U85 (N_85,In_169,In_444);
and U86 (N_86,In_231,In_254);
or U87 (N_87,In_109,In_413);
or U88 (N_88,In_287,In_166);
nor U89 (N_89,In_240,In_357);
or U90 (N_90,In_404,In_36);
and U91 (N_91,In_350,In_367);
or U92 (N_92,In_473,In_336);
and U93 (N_93,In_414,In_47);
or U94 (N_94,In_29,In_428);
or U95 (N_95,In_256,In_340);
and U96 (N_96,In_388,In_318);
and U97 (N_97,In_15,In_136);
or U98 (N_98,In_359,In_121);
nor U99 (N_99,In_38,In_181);
or U100 (N_100,In_101,N_37);
or U101 (N_101,In_5,In_479);
nor U102 (N_102,In_63,In_489);
nand U103 (N_103,N_76,In_285);
nor U104 (N_104,N_44,In_145);
or U105 (N_105,In_191,N_93);
nor U106 (N_106,In_3,In_151);
and U107 (N_107,In_353,In_486);
and U108 (N_108,In_218,In_75);
and U109 (N_109,In_405,In_421);
or U110 (N_110,In_115,In_284);
or U111 (N_111,N_45,N_47);
or U112 (N_112,N_7,In_365);
and U113 (N_113,N_78,In_84);
nor U114 (N_114,In_411,N_68);
nor U115 (N_115,In_442,N_43);
and U116 (N_116,In_345,N_26);
nand U117 (N_117,In_328,In_217);
and U118 (N_118,N_69,In_61);
nor U119 (N_119,In_435,N_94);
nor U120 (N_120,In_141,N_99);
and U121 (N_121,In_288,In_395);
and U122 (N_122,N_90,In_278);
or U123 (N_123,In_232,N_12);
or U124 (N_124,In_14,In_393);
or U125 (N_125,In_100,N_96);
and U126 (N_126,In_463,In_56);
nand U127 (N_127,In_135,In_175);
or U128 (N_128,In_156,N_65);
nor U129 (N_129,N_97,In_275);
nand U130 (N_130,In_483,In_174);
nand U131 (N_131,N_77,N_29);
nor U132 (N_132,In_352,In_253);
nor U133 (N_133,In_94,In_402);
nand U134 (N_134,In_387,N_62);
nand U135 (N_135,In_130,N_20);
nand U136 (N_136,N_30,In_55);
nand U137 (N_137,In_178,In_446);
or U138 (N_138,In_301,In_335);
nor U139 (N_139,In_283,In_92);
and U140 (N_140,In_362,In_454);
or U141 (N_141,N_64,In_317);
nor U142 (N_142,In_206,In_0);
or U143 (N_143,In_189,In_16);
or U144 (N_144,In_306,In_460);
nor U145 (N_145,In_160,In_227);
nand U146 (N_146,In_182,N_72);
or U147 (N_147,N_2,In_28);
or U148 (N_148,In_293,In_64);
nor U149 (N_149,In_147,In_67);
or U150 (N_150,In_257,N_67);
nand U151 (N_151,In_294,In_274);
and U152 (N_152,In_97,In_396);
nor U153 (N_153,In_468,N_49);
or U154 (N_154,In_476,In_48);
nand U155 (N_155,In_424,In_415);
or U156 (N_156,In_241,In_226);
or U157 (N_157,In_248,In_243);
or U158 (N_158,In_222,In_91);
or U159 (N_159,N_129,In_321);
nor U160 (N_160,In_469,In_279);
nand U161 (N_161,In_143,N_125);
nor U162 (N_162,In_366,In_173);
nand U163 (N_163,In_172,N_108);
nand U164 (N_164,N_82,N_84);
nor U165 (N_165,In_445,In_50);
nor U166 (N_166,N_23,N_104);
and U167 (N_167,N_114,N_105);
nor U168 (N_168,N_101,In_485);
nand U169 (N_169,In_412,In_235);
nor U170 (N_170,N_33,In_45);
nor U171 (N_171,N_106,N_137);
nand U172 (N_172,In_137,In_96);
nand U173 (N_173,In_211,N_39);
nand U174 (N_174,In_364,In_35);
or U175 (N_175,N_127,N_10);
and U176 (N_176,In_146,In_210);
or U177 (N_177,In_449,N_38);
nor U178 (N_178,In_431,In_474);
nor U179 (N_179,In_272,In_58);
nor U180 (N_180,In_448,In_420);
nand U181 (N_181,N_140,In_499);
and U182 (N_182,In_349,In_399);
nand U183 (N_183,In_66,In_103);
nand U184 (N_184,In_383,N_128);
nand U185 (N_185,N_91,In_416);
nor U186 (N_186,In_381,In_113);
and U187 (N_187,In_1,In_207);
nand U188 (N_188,N_115,N_144);
and U189 (N_189,In_247,N_66);
nor U190 (N_190,N_41,In_266);
nand U191 (N_191,N_79,N_42);
and U192 (N_192,N_102,In_417);
and U193 (N_193,In_400,In_436);
nor U194 (N_194,N_46,N_61);
nand U195 (N_195,In_200,N_56);
nor U196 (N_196,In_60,In_333);
nor U197 (N_197,In_4,In_472);
or U198 (N_198,In_419,N_19);
nand U199 (N_199,N_113,N_80);
nand U200 (N_200,N_176,N_89);
nor U201 (N_201,In_439,In_401);
and U202 (N_202,N_193,In_37);
nand U203 (N_203,In_22,N_22);
nand U204 (N_204,N_117,In_385);
xnor U205 (N_205,N_135,In_155);
nand U206 (N_206,In_19,In_239);
nor U207 (N_207,In_390,N_27);
or U208 (N_208,In_297,N_51);
and U209 (N_209,N_191,In_441);
or U210 (N_210,In_40,In_496);
nor U211 (N_211,N_124,In_298);
or U212 (N_212,N_195,In_216);
nor U213 (N_213,In_426,N_153);
nand U214 (N_214,N_50,In_371);
and U215 (N_215,N_54,In_140);
nand U216 (N_216,In_125,In_356);
nand U217 (N_217,In_119,N_166);
nand U218 (N_218,In_337,N_58);
nor U219 (N_219,In_33,N_98);
and U220 (N_220,N_189,In_490);
and U221 (N_221,N_192,In_167);
and U222 (N_222,N_143,In_201);
nand U223 (N_223,In_323,N_118);
or U224 (N_224,N_151,In_152);
and U225 (N_225,In_198,In_281);
or U226 (N_226,N_103,In_6);
or U227 (N_227,N_107,In_204);
and U228 (N_228,N_146,In_139);
or U229 (N_229,In_327,In_423);
nand U230 (N_230,In_229,N_85);
nand U231 (N_231,In_467,N_187);
nor U232 (N_232,In_251,In_492);
and U233 (N_233,N_184,N_198);
nand U234 (N_234,N_134,In_88);
nor U235 (N_235,N_48,N_75);
or U236 (N_236,In_9,In_351);
nand U237 (N_237,In_495,N_116);
or U238 (N_238,N_110,In_59);
nor U239 (N_239,In_233,In_271);
nand U240 (N_240,In_23,In_219);
or U241 (N_241,In_450,N_152);
nand U242 (N_242,In_224,N_169);
nor U243 (N_243,N_92,In_361);
nor U244 (N_244,In_209,N_149);
nor U245 (N_245,In_118,In_296);
or U246 (N_246,In_434,N_13);
or U247 (N_247,N_70,In_183);
and U248 (N_248,N_31,N_138);
nand U249 (N_249,In_382,In_378);
xor U250 (N_250,N_236,In_339);
nand U251 (N_251,N_174,N_177);
or U252 (N_252,In_32,In_149);
and U253 (N_253,In_398,In_481);
nor U254 (N_254,N_234,N_130);
nor U255 (N_255,In_418,N_55);
nor U256 (N_256,In_380,N_60);
nor U257 (N_257,N_6,N_157);
and U258 (N_258,In_322,In_161);
nand U259 (N_259,N_119,In_447);
or U260 (N_260,In_282,N_222);
and U261 (N_261,N_207,In_403);
and U262 (N_262,In_269,In_494);
nand U263 (N_263,N_243,N_247);
nor U264 (N_264,In_49,N_246);
or U265 (N_265,In_372,In_289);
or U266 (N_266,N_231,In_408);
nand U267 (N_267,N_217,N_112);
nor U268 (N_268,N_142,N_156);
nand U269 (N_269,In_138,In_46);
or U270 (N_270,In_332,N_73);
nor U271 (N_271,In_164,In_153);
nand U272 (N_272,In_314,N_148);
nand U273 (N_273,In_180,N_214);
and U274 (N_274,In_196,N_219);
nand U275 (N_275,N_167,In_72);
and U276 (N_276,N_178,In_107);
or U277 (N_277,In_462,N_242);
and U278 (N_278,N_163,N_81);
and U279 (N_279,N_52,N_186);
and U280 (N_280,N_175,N_206);
or U281 (N_281,N_100,N_185);
nand U282 (N_282,In_41,In_268);
and U283 (N_283,N_160,In_406);
and U284 (N_284,In_331,N_223);
and U285 (N_285,N_216,In_263);
nor U286 (N_286,N_190,N_181);
nor U287 (N_287,In_341,N_201);
and U288 (N_288,In_71,In_52);
and U289 (N_289,In_179,In_2);
and U290 (N_290,In_394,In_354);
nand U291 (N_291,N_154,In_150);
or U292 (N_292,In_213,N_16);
and U293 (N_293,N_173,N_233);
or U294 (N_294,In_452,In_236);
nor U295 (N_295,N_87,N_126);
nand U296 (N_296,In_304,N_3);
and U297 (N_297,In_163,N_210);
and U298 (N_298,N_229,N_199);
nand U299 (N_299,In_77,N_196);
or U300 (N_300,N_204,In_82);
nor U301 (N_301,N_285,N_268);
nor U302 (N_302,N_272,N_287);
nor U303 (N_303,N_256,N_269);
nor U304 (N_304,N_59,In_391);
or U305 (N_305,N_57,In_342);
nand U306 (N_306,N_182,In_465);
or U307 (N_307,In_93,In_215);
and U308 (N_308,N_71,N_265);
and U309 (N_309,N_288,N_227);
nand U310 (N_310,In_477,In_464);
nor U311 (N_311,In_493,N_297);
nor U312 (N_312,N_238,In_104);
or U313 (N_313,N_259,In_348);
nand U314 (N_314,N_120,N_1);
nand U315 (N_315,In_475,N_278);
nor U316 (N_316,In_43,In_429);
nor U317 (N_317,In_377,In_457);
nand U318 (N_318,N_179,N_248);
and U319 (N_319,N_271,N_266);
and U320 (N_320,N_228,N_250);
nor U321 (N_321,N_183,N_224);
and U322 (N_322,In_186,In_488);
and U323 (N_323,N_239,In_252);
and U324 (N_324,N_133,N_215);
nor U325 (N_325,N_245,In_311);
nand U326 (N_326,In_176,In_124);
and U327 (N_327,In_302,In_68);
and U328 (N_328,N_53,N_136);
or U329 (N_329,N_208,N_158);
or U330 (N_330,N_289,N_277);
nor U331 (N_331,In_242,N_244);
or U332 (N_332,N_171,N_273);
and U333 (N_333,N_209,N_164);
nand U334 (N_334,N_282,N_170);
nor U335 (N_335,In_159,N_132);
and U336 (N_336,N_63,In_453);
or U337 (N_337,N_202,N_279);
and U338 (N_338,N_257,N_200);
and U339 (N_339,In_369,N_292);
nand U340 (N_340,N_295,N_218);
or U341 (N_341,N_188,N_203);
or U342 (N_342,N_291,In_430);
nor U343 (N_343,In_250,N_25);
nor U344 (N_344,N_220,N_74);
nor U345 (N_345,N_274,In_478);
nor U346 (N_346,N_141,In_214);
nor U347 (N_347,N_212,N_275);
nor U348 (N_348,N_286,N_36);
or U349 (N_349,In_78,In_25);
or U350 (N_350,N_168,N_83);
and U351 (N_351,N_334,N_290);
nand U352 (N_352,In_187,In_410);
nor U353 (N_353,N_333,In_65);
nor U354 (N_354,N_131,N_213);
and U355 (N_355,In_437,N_255);
or U356 (N_356,N_0,N_8);
and U357 (N_357,N_342,N_237);
or U358 (N_358,In_259,N_330);
nor U359 (N_359,N_122,In_81);
nand U360 (N_360,In_128,N_260);
nand U361 (N_361,In_295,In_237);
or U362 (N_362,N_348,N_258);
nand U363 (N_363,N_264,N_336);
or U364 (N_364,N_263,N_32);
or U365 (N_365,N_24,In_171);
or U366 (N_366,N_109,N_298);
or U367 (N_367,N_254,N_232);
nor U368 (N_368,N_139,N_284);
and U369 (N_369,N_155,N_121);
and U370 (N_370,N_347,In_62);
and U371 (N_371,N_338,N_270);
nand U372 (N_372,N_162,N_280);
nand U373 (N_373,N_318,N_314);
and U374 (N_374,N_345,N_253);
nor U375 (N_375,In_368,In_131);
or U376 (N_376,In_220,N_283);
or U377 (N_377,In_120,N_15);
nand U378 (N_378,In_18,In_225);
and U379 (N_379,In_102,N_306);
nor U380 (N_380,N_111,N_249);
nand U381 (N_381,N_340,N_300);
and U382 (N_382,In_34,N_88);
and U383 (N_383,In_246,N_305);
or U384 (N_384,N_328,N_332);
nand U385 (N_385,N_145,In_291);
or U386 (N_386,N_321,N_299);
and U387 (N_387,N_276,In_276);
and U388 (N_388,N_261,N_325);
and U389 (N_389,N_303,N_240);
and U390 (N_390,N_317,N_315);
nand U391 (N_391,In_438,N_225);
and U392 (N_392,In_432,N_327);
nand U393 (N_393,N_180,N_316);
xor U394 (N_394,N_346,N_307);
or U395 (N_395,In_99,N_251);
and U396 (N_396,N_329,N_343);
or U397 (N_397,N_165,In_106);
or U398 (N_398,N_322,N_211);
nor U399 (N_399,In_111,In_238);
nor U400 (N_400,N_360,N_150);
or U401 (N_401,N_364,N_319);
and U402 (N_402,N_381,N_302);
and U403 (N_403,In_154,N_147);
nand U404 (N_404,N_367,N_312);
and U405 (N_405,N_382,N_358);
nor U406 (N_406,N_378,N_351);
nor U407 (N_407,N_361,N_313);
xnor U408 (N_408,N_262,N_326);
nand U409 (N_409,N_172,N_301);
nand U410 (N_410,In_358,N_365);
nand U411 (N_411,N_161,N_324);
nor U412 (N_412,N_241,N_359);
nand U413 (N_413,N_379,N_383);
nor U414 (N_414,N_389,N_323);
and U415 (N_415,N_252,N_384);
or U416 (N_416,N_357,N_337);
nor U417 (N_417,N_353,N_397);
xor U418 (N_418,N_398,N_374);
nor U419 (N_419,N_375,N_386);
and U420 (N_420,N_394,N_311);
or U421 (N_421,N_372,In_114);
and U422 (N_422,N_335,N_86);
nor U423 (N_423,N_373,N_293);
nand U424 (N_424,N_320,N_205);
nand U425 (N_425,N_390,N_296);
nor U426 (N_426,N_370,N_194);
nand U427 (N_427,N_356,N_304);
nand U428 (N_428,N_352,N_380);
nand U429 (N_429,N_354,N_230);
or U430 (N_430,N_371,N_350);
nand U431 (N_431,N_362,N_235);
or U432 (N_432,N_226,N_309);
nor U433 (N_433,N_355,N_368);
and U434 (N_434,N_267,N_308);
or U435 (N_435,N_281,N_391);
and U436 (N_436,N_396,N_392);
or U437 (N_437,N_123,N_341);
nand U438 (N_438,N_393,N_221);
nand U439 (N_439,N_331,N_366);
nor U440 (N_440,N_387,N_369);
or U441 (N_441,N_376,N_310);
or U442 (N_442,N_339,N_388);
and U443 (N_443,N_349,In_205);
nand U444 (N_444,N_399,N_363);
nor U445 (N_445,N_294,N_344);
nor U446 (N_446,N_377,N_385);
nand U447 (N_447,N_395,N_159);
nor U448 (N_448,In_343,N_95);
or U449 (N_449,N_11,N_197);
and U450 (N_450,N_432,N_441);
and U451 (N_451,N_434,N_435);
and U452 (N_452,N_440,N_426);
or U453 (N_453,N_407,N_428);
nor U454 (N_454,N_401,N_439);
or U455 (N_455,N_446,N_420);
nand U456 (N_456,N_424,N_412);
xnor U457 (N_457,N_418,N_409);
or U458 (N_458,N_429,N_442);
nor U459 (N_459,N_425,N_447);
and U460 (N_460,N_405,N_437);
or U461 (N_461,N_433,N_438);
nor U462 (N_462,N_419,N_400);
nor U463 (N_463,N_427,N_404);
and U464 (N_464,N_422,N_411);
and U465 (N_465,N_414,N_410);
nor U466 (N_466,N_445,N_423);
nor U467 (N_467,N_421,N_415);
nor U468 (N_468,N_449,N_443);
or U469 (N_469,N_413,N_430);
nor U470 (N_470,N_444,N_448);
nand U471 (N_471,N_403,N_402);
nand U472 (N_472,N_436,N_417);
nand U473 (N_473,N_431,N_416);
nor U474 (N_474,N_406,N_408);
nor U475 (N_475,N_445,N_405);
and U476 (N_476,N_429,N_436);
nand U477 (N_477,N_447,N_413);
nand U478 (N_478,N_406,N_413);
nand U479 (N_479,N_435,N_412);
and U480 (N_480,N_410,N_428);
and U481 (N_481,N_433,N_440);
nand U482 (N_482,N_440,N_413);
nor U483 (N_483,N_411,N_433);
nor U484 (N_484,N_417,N_400);
nor U485 (N_485,N_414,N_402);
nand U486 (N_486,N_422,N_433);
nor U487 (N_487,N_411,N_403);
nor U488 (N_488,N_411,N_427);
nand U489 (N_489,N_423,N_439);
xnor U490 (N_490,N_426,N_418);
and U491 (N_491,N_430,N_448);
nand U492 (N_492,N_441,N_411);
or U493 (N_493,N_421,N_425);
or U494 (N_494,N_415,N_434);
and U495 (N_495,N_441,N_436);
nand U496 (N_496,N_403,N_414);
and U497 (N_497,N_410,N_438);
nor U498 (N_498,N_439,N_424);
and U499 (N_499,N_445,N_404);
or U500 (N_500,N_495,N_474);
nor U501 (N_501,N_460,N_491);
nor U502 (N_502,N_497,N_467);
nand U503 (N_503,N_478,N_485);
nand U504 (N_504,N_464,N_489);
or U505 (N_505,N_452,N_471);
nor U506 (N_506,N_492,N_483);
nor U507 (N_507,N_469,N_458);
nand U508 (N_508,N_488,N_476);
or U509 (N_509,N_462,N_494);
nand U510 (N_510,N_466,N_461);
and U511 (N_511,N_481,N_496);
and U512 (N_512,N_455,N_472);
nor U513 (N_513,N_457,N_468);
nand U514 (N_514,N_487,N_477);
and U515 (N_515,N_475,N_459);
and U516 (N_516,N_493,N_484);
nand U517 (N_517,N_486,N_463);
nor U518 (N_518,N_453,N_473);
and U519 (N_519,N_480,N_499);
nor U520 (N_520,N_482,N_451);
or U521 (N_521,N_454,N_490);
nor U522 (N_522,N_456,N_498);
or U523 (N_523,N_450,N_470);
nand U524 (N_524,N_465,N_479);
or U525 (N_525,N_482,N_471);
or U526 (N_526,N_483,N_478);
nor U527 (N_527,N_483,N_475);
and U528 (N_528,N_459,N_471);
and U529 (N_529,N_469,N_456);
nand U530 (N_530,N_483,N_463);
nand U531 (N_531,N_480,N_467);
nor U532 (N_532,N_482,N_477);
and U533 (N_533,N_461,N_476);
nand U534 (N_534,N_451,N_480);
nand U535 (N_535,N_479,N_466);
or U536 (N_536,N_455,N_497);
and U537 (N_537,N_480,N_486);
nand U538 (N_538,N_464,N_475);
nand U539 (N_539,N_451,N_471);
nor U540 (N_540,N_483,N_465);
nor U541 (N_541,N_470,N_455);
and U542 (N_542,N_451,N_464);
and U543 (N_543,N_451,N_473);
or U544 (N_544,N_460,N_454);
or U545 (N_545,N_493,N_467);
nor U546 (N_546,N_456,N_475);
nor U547 (N_547,N_453,N_498);
and U548 (N_548,N_468,N_472);
xnor U549 (N_549,N_494,N_459);
and U550 (N_550,N_517,N_533);
and U551 (N_551,N_521,N_506);
nand U552 (N_552,N_515,N_546);
or U553 (N_553,N_519,N_532);
and U554 (N_554,N_505,N_500);
and U555 (N_555,N_535,N_508);
or U556 (N_556,N_507,N_511);
nor U557 (N_557,N_524,N_513);
nor U558 (N_558,N_502,N_510);
nor U559 (N_559,N_509,N_534);
and U560 (N_560,N_549,N_503);
nand U561 (N_561,N_547,N_541);
and U562 (N_562,N_525,N_516);
and U563 (N_563,N_501,N_529);
and U564 (N_564,N_545,N_514);
and U565 (N_565,N_542,N_543);
or U566 (N_566,N_536,N_548);
nand U567 (N_567,N_504,N_537);
or U568 (N_568,N_540,N_512);
nand U569 (N_569,N_522,N_518);
or U570 (N_570,N_530,N_527);
and U571 (N_571,N_526,N_539);
or U572 (N_572,N_544,N_528);
and U573 (N_573,N_520,N_538);
or U574 (N_574,N_531,N_523);
nand U575 (N_575,N_517,N_531);
nor U576 (N_576,N_517,N_534);
or U577 (N_577,N_530,N_533);
and U578 (N_578,N_501,N_513);
and U579 (N_579,N_533,N_519);
nor U580 (N_580,N_526,N_529);
or U581 (N_581,N_520,N_535);
nand U582 (N_582,N_515,N_529);
and U583 (N_583,N_505,N_507);
nor U584 (N_584,N_548,N_510);
nor U585 (N_585,N_505,N_549);
nand U586 (N_586,N_539,N_530);
nand U587 (N_587,N_509,N_543);
nor U588 (N_588,N_543,N_510);
or U589 (N_589,N_511,N_531);
or U590 (N_590,N_542,N_540);
nand U591 (N_591,N_522,N_502);
nor U592 (N_592,N_501,N_537);
and U593 (N_593,N_543,N_532);
and U594 (N_594,N_511,N_528);
nand U595 (N_595,N_531,N_509);
nor U596 (N_596,N_533,N_507);
and U597 (N_597,N_545,N_532);
and U598 (N_598,N_529,N_503);
nor U599 (N_599,N_524,N_528);
or U600 (N_600,N_599,N_580);
nand U601 (N_601,N_587,N_551);
and U602 (N_602,N_550,N_553);
nand U603 (N_603,N_564,N_576);
or U604 (N_604,N_595,N_578);
nor U605 (N_605,N_566,N_562);
nor U606 (N_606,N_589,N_555);
nor U607 (N_607,N_563,N_556);
and U608 (N_608,N_571,N_596);
or U609 (N_609,N_577,N_581);
nand U610 (N_610,N_557,N_574);
nand U611 (N_611,N_558,N_590);
nand U612 (N_612,N_584,N_559);
and U613 (N_613,N_560,N_565);
and U614 (N_614,N_570,N_575);
nor U615 (N_615,N_552,N_567);
nor U616 (N_616,N_592,N_573);
and U617 (N_617,N_585,N_588);
nor U618 (N_618,N_597,N_561);
nor U619 (N_619,N_569,N_591);
and U620 (N_620,N_572,N_583);
and U621 (N_621,N_582,N_586);
nand U622 (N_622,N_594,N_568);
nor U623 (N_623,N_598,N_579);
nor U624 (N_624,N_593,N_554);
or U625 (N_625,N_562,N_582);
and U626 (N_626,N_586,N_571);
or U627 (N_627,N_553,N_585);
nand U628 (N_628,N_585,N_557);
nand U629 (N_629,N_584,N_585);
nand U630 (N_630,N_574,N_555);
or U631 (N_631,N_599,N_562);
nand U632 (N_632,N_557,N_593);
or U633 (N_633,N_555,N_551);
or U634 (N_634,N_569,N_587);
nand U635 (N_635,N_563,N_565);
and U636 (N_636,N_599,N_582);
nand U637 (N_637,N_559,N_571);
or U638 (N_638,N_569,N_590);
nand U639 (N_639,N_599,N_586);
or U640 (N_640,N_569,N_570);
or U641 (N_641,N_587,N_560);
or U642 (N_642,N_588,N_589);
and U643 (N_643,N_580,N_573);
nor U644 (N_644,N_554,N_584);
or U645 (N_645,N_597,N_562);
or U646 (N_646,N_583,N_577);
nand U647 (N_647,N_550,N_556);
nor U648 (N_648,N_580,N_576);
and U649 (N_649,N_565,N_564);
or U650 (N_650,N_603,N_620);
or U651 (N_651,N_605,N_616);
nand U652 (N_652,N_612,N_643);
or U653 (N_653,N_633,N_614);
and U654 (N_654,N_649,N_629);
nand U655 (N_655,N_645,N_624);
or U656 (N_656,N_648,N_622);
and U657 (N_657,N_606,N_636);
xnor U658 (N_658,N_619,N_610);
or U659 (N_659,N_627,N_641);
and U660 (N_660,N_604,N_644);
nand U661 (N_661,N_637,N_625);
nor U662 (N_662,N_600,N_607);
and U663 (N_663,N_617,N_613);
or U664 (N_664,N_601,N_602);
nand U665 (N_665,N_623,N_608);
nand U666 (N_666,N_628,N_634);
nand U667 (N_667,N_626,N_630);
nand U668 (N_668,N_638,N_631);
or U669 (N_669,N_640,N_647);
nand U670 (N_670,N_609,N_611);
or U671 (N_671,N_618,N_632);
or U672 (N_672,N_615,N_635);
nor U673 (N_673,N_639,N_646);
nor U674 (N_674,N_642,N_621);
and U675 (N_675,N_612,N_623);
and U676 (N_676,N_612,N_618);
and U677 (N_677,N_601,N_619);
or U678 (N_678,N_600,N_606);
and U679 (N_679,N_602,N_635);
nand U680 (N_680,N_642,N_628);
or U681 (N_681,N_620,N_619);
nand U682 (N_682,N_607,N_648);
or U683 (N_683,N_639,N_637);
or U684 (N_684,N_625,N_642);
nand U685 (N_685,N_635,N_631);
or U686 (N_686,N_600,N_640);
and U687 (N_687,N_606,N_623);
and U688 (N_688,N_607,N_620);
nor U689 (N_689,N_612,N_642);
and U690 (N_690,N_602,N_600);
nor U691 (N_691,N_630,N_646);
nand U692 (N_692,N_624,N_613);
or U693 (N_693,N_600,N_611);
or U694 (N_694,N_629,N_639);
and U695 (N_695,N_626,N_601);
nand U696 (N_696,N_609,N_621);
or U697 (N_697,N_639,N_619);
nand U698 (N_698,N_617,N_625);
nor U699 (N_699,N_603,N_600);
and U700 (N_700,N_687,N_683);
nor U701 (N_701,N_662,N_664);
and U702 (N_702,N_696,N_654);
and U703 (N_703,N_666,N_675);
nor U704 (N_704,N_693,N_698);
nand U705 (N_705,N_690,N_672);
nand U706 (N_706,N_658,N_682);
nor U707 (N_707,N_691,N_677);
nor U708 (N_708,N_657,N_681);
and U709 (N_709,N_694,N_653);
or U710 (N_710,N_652,N_689);
or U711 (N_711,N_680,N_655);
nor U712 (N_712,N_676,N_660);
nor U713 (N_713,N_692,N_668);
nor U714 (N_714,N_665,N_685);
nor U715 (N_715,N_667,N_684);
or U716 (N_716,N_699,N_688);
and U717 (N_717,N_673,N_674);
or U718 (N_718,N_656,N_679);
and U719 (N_719,N_669,N_686);
or U720 (N_720,N_678,N_659);
and U721 (N_721,N_695,N_650);
nand U722 (N_722,N_697,N_661);
nand U723 (N_723,N_670,N_651);
nand U724 (N_724,N_663,N_671);
nor U725 (N_725,N_676,N_687);
and U726 (N_726,N_684,N_658);
nor U727 (N_727,N_656,N_677);
nor U728 (N_728,N_652,N_662);
nand U729 (N_729,N_655,N_682);
nor U730 (N_730,N_668,N_699);
nor U731 (N_731,N_671,N_690);
nor U732 (N_732,N_669,N_696);
and U733 (N_733,N_676,N_668);
and U734 (N_734,N_657,N_650);
nand U735 (N_735,N_697,N_660);
and U736 (N_736,N_687,N_662);
xnor U737 (N_737,N_676,N_664);
nor U738 (N_738,N_657,N_661);
nor U739 (N_739,N_655,N_651);
or U740 (N_740,N_681,N_662);
nor U741 (N_741,N_695,N_653);
nor U742 (N_742,N_679,N_682);
nand U743 (N_743,N_671,N_684);
or U744 (N_744,N_677,N_650);
nor U745 (N_745,N_699,N_684);
nor U746 (N_746,N_661,N_699);
and U747 (N_747,N_696,N_665);
and U748 (N_748,N_669,N_662);
and U749 (N_749,N_697,N_652);
nor U750 (N_750,N_727,N_735);
and U751 (N_751,N_707,N_721);
nor U752 (N_752,N_720,N_738);
and U753 (N_753,N_713,N_749);
and U754 (N_754,N_747,N_709);
nor U755 (N_755,N_723,N_743);
and U756 (N_756,N_728,N_725);
nor U757 (N_757,N_736,N_729);
or U758 (N_758,N_704,N_710);
nand U759 (N_759,N_703,N_712);
nand U760 (N_760,N_711,N_731);
nor U761 (N_761,N_717,N_746);
nand U762 (N_762,N_700,N_748);
nand U763 (N_763,N_734,N_708);
nand U764 (N_764,N_724,N_737);
and U765 (N_765,N_745,N_744);
nor U766 (N_766,N_715,N_741);
nand U767 (N_767,N_714,N_733);
nor U768 (N_768,N_719,N_740);
nand U769 (N_769,N_726,N_742);
nand U770 (N_770,N_702,N_730);
or U771 (N_771,N_722,N_706);
or U772 (N_772,N_701,N_732);
nor U773 (N_773,N_739,N_705);
and U774 (N_774,N_716,N_718);
nand U775 (N_775,N_736,N_731);
nand U776 (N_776,N_726,N_722);
nand U777 (N_777,N_734,N_709);
nand U778 (N_778,N_730,N_725);
or U779 (N_779,N_706,N_725);
nand U780 (N_780,N_722,N_705);
xnor U781 (N_781,N_746,N_708);
and U782 (N_782,N_722,N_700);
nand U783 (N_783,N_706,N_720);
or U784 (N_784,N_723,N_724);
or U785 (N_785,N_716,N_730);
nor U786 (N_786,N_711,N_712);
nor U787 (N_787,N_741,N_702);
or U788 (N_788,N_704,N_723);
nand U789 (N_789,N_712,N_733);
nor U790 (N_790,N_709,N_724);
or U791 (N_791,N_740,N_721);
nand U792 (N_792,N_730,N_746);
nor U793 (N_793,N_749,N_709);
or U794 (N_794,N_728,N_700);
nor U795 (N_795,N_722,N_720);
nor U796 (N_796,N_707,N_748);
or U797 (N_797,N_729,N_725);
nand U798 (N_798,N_745,N_728);
and U799 (N_799,N_723,N_728);
or U800 (N_800,N_776,N_790);
nor U801 (N_801,N_782,N_794);
and U802 (N_802,N_766,N_750);
nand U803 (N_803,N_770,N_771);
and U804 (N_804,N_787,N_792);
nor U805 (N_805,N_784,N_767);
or U806 (N_806,N_777,N_786);
nand U807 (N_807,N_780,N_772);
nor U808 (N_808,N_797,N_754);
or U809 (N_809,N_795,N_781);
and U810 (N_810,N_761,N_765);
nand U811 (N_811,N_791,N_778);
nor U812 (N_812,N_759,N_788);
and U813 (N_813,N_760,N_758);
nor U814 (N_814,N_773,N_764);
and U815 (N_815,N_752,N_796);
nand U816 (N_816,N_755,N_789);
nand U817 (N_817,N_775,N_753);
and U818 (N_818,N_769,N_799);
or U819 (N_819,N_762,N_774);
and U820 (N_820,N_793,N_783);
or U821 (N_821,N_779,N_768);
nand U822 (N_822,N_763,N_756);
or U823 (N_823,N_751,N_798);
nand U824 (N_824,N_785,N_757);
nor U825 (N_825,N_753,N_762);
nor U826 (N_826,N_797,N_771);
nand U827 (N_827,N_758,N_799);
and U828 (N_828,N_754,N_783);
nand U829 (N_829,N_774,N_778);
nand U830 (N_830,N_753,N_766);
nand U831 (N_831,N_772,N_773);
or U832 (N_832,N_776,N_763);
and U833 (N_833,N_763,N_785);
and U834 (N_834,N_799,N_787);
nand U835 (N_835,N_796,N_761);
and U836 (N_836,N_791,N_784);
nand U837 (N_837,N_795,N_770);
and U838 (N_838,N_768,N_750);
or U839 (N_839,N_788,N_751);
nand U840 (N_840,N_751,N_795);
or U841 (N_841,N_760,N_757);
xnor U842 (N_842,N_762,N_758);
nor U843 (N_843,N_796,N_762);
or U844 (N_844,N_791,N_796);
and U845 (N_845,N_775,N_792);
nand U846 (N_846,N_774,N_766);
nor U847 (N_847,N_784,N_761);
nand U848 (N_848,N_758,N_751);
nor U849 (N_849,N_750,N_781);
and U850 (N_850,N_831,N_844);
nand U851 (N_851,N_819,N_836);
or U852 (N_852,N_805,N_817);
nor U853 (N_853,N_839,N_843);
or U854 (N_854,N_834,N_824);
nor U855 (N_855,N_823,N_806);
nor U856 (N_856,N_818,N_814);
nor U857 (N_857,N_807,N_840);
or U858 (N_858,N_815,N_822);
or U859 (N_859,N_804,N_813);
or U860 (N_860,N_842,N_845);
or U861 (N_861,N_809,N_800);
nor U862 (N_862,N_826,N_846);
nor U863 (N_863,N_802,N_847);
or U864 (N_864,N_835,N_837);
nor U865 (N_865,N_848,N_830);
nand U866 (N_866,N_811,N_816);
nor U867 (N_867,N_832,N_833);
nand U868 (N_868,N_828,N_808);
and U869 (N_869,N_810,N_820);
xnor U870 (N_870,N_821,N_801);
or U871 (N_871,N_829,N_827);
nand U872 (N_872,N_849,N_812);
nand U873 (N_873,N_838,N_803);
nor U874 (N_874,N_841,N_825);
or U875 (N_875,N_837,N_840);
nand U876 (N_876,N_809,N_831);
or U877 (N_877,N_826,N_842);
nor U878 (N_878,N_804,N_848);
or U879 (N_879,N_829,N_834);
and U880 (N_880,N_833,N_830);
xor U881 (N_881,N_849,N_847);
nor U882 (N_882,N_849,N_848);
and U883 (N_883,N_801,N_827);
and U884 (N_884,N_834,N_839);
nor U885 (N_885,N_800,N_838);
and U886 (N_886,N_804,N_823);
nand U887 (N_887,N_820,N_847);
or U888 (N_888,N_838,N_849);
nand U889 (N_889,N_838,N_836);
nor U890 (N_890,N_801,N_822);
nor U891 (N_891,N_802,N_829);
and U892 (N_892,N_846,N_812);
nand U893 (N_893,N_815,N_836);
nor U894 (N_894,N_842,N_835);
and U895 (N_895,N_811,N_809);
and U896 (N_896,N_835,N_847);
nor U897 (N_897,N_830,N_842);
or U898 (N_898,N_830,N_846);
and U899 (N_899,N_815,N_821);
or U900 (N_900,N_874,N_891);
nand U901 (N_901,N_882,N_895);
nor U902 (N_902,N_881,N_878);
nor U903 (N_903,N_887,N_897);
and U904 (N_904,N_875,N_853);
and U905 (N_905,N_873,N_855);
nor U906 (N_906,N_883,N_852);
or U907 (N_907,N_892,N_864);
and U908 (N_908,N_859,N_850);
and U909 (N_909,N_898,N_876);
nand U910 (N_910,N_857,N_863);
nand U911 (N_911,N_869,N_860);
nand U912 (N_912,N_899,N_856);
or U913 (N_913,N_861,N_862);
or U914 (N_914,N_870,N_880);
or U915 (N_915,N_867,N_885);
nor U916 (N_916,N_865,N_866);
nand U917 (N_917,N_851,N_894);
and U918 (N_918,N_896,N_872);
nand U919 (N_919,N_868,N_888);
nor U920 (N_920,N_889,N_871);
nand U921 (N_921,N_890,N_886);
nor U922 (N_922,N_858,N_884);
or U923 (N_923,N_854,N_893);
nand U924 (N_924,N_877,N_879);
or U925 (N_925,N_891,N_863);
and U926 (N_926,N_875,N_859);
nor U927 (N_927,N_879,N_850);
or U928 (N_928,N_893,N_895);
nand U929 (N_929,N_865,N_855);
or U930 (N_930,N_867,N_895);
and U931 (N_931,N_874,N_871);
and U932 (N_932,N_854,N_875);
or U933 (N_933,N_852,N_873);
and U934 (N_934,N_876,N_897);
or U935 (N_935,N_871,N_895);
or U936 (N_936,N_859,N_881);
or U937 (N_937,N_869,N_896);
or U938 (N_938,N_852,N_867);
nor U939 (N_939,N_879,N_851);
nor U940 (N_940,N_868,N_869);
or U941 (N_941,N_890,N_858);
or U942 (N_942,N_877,N_872);
nand U943 (N_943,N_887,N_892);
or U944 (N_944,N_874,N_862);
nand U945 (N_945,N_852,N_896);
nand U946 (N_946,N_852,N_892);
or U947 (N_947,N_878,N_874);
nand U948 (N_948,N_867,N_853);
and U949 (N_949,N_889,N_883);
or U950 (N_950,N_933,N_949);
nor U951 (N_951,N_911,N_919);
and U952 (N_952,N_923,N_906);
nand U953 (N_953,N_913,N_935);
nand U954 (N_954,N_900,N_939);
and U955 (N_955,N_918,N_917);
nor U956 (N_956,N_926,N_934);
nor U957 (N_957,N_942,N_924);
and U958 (N_958,N_901,N_938);
nor U959 (N_959,N_940,N_927);
and U960 (N_960,N_920,N_931);
or U961 (N_961,N_945,N_930);
nand U962 (N_962,N_928,N_947);
or U963 (N_963,N_908,N_943);
or U964 (N_964,N_925,N_915);
nor U965 (N_965,N_936,N_903);
nand U966 (N_966,N_929,N_948);
and U967 (N_967,N_909,N_941);
nor U968 (N_968,N_946,N_944);
or U969 (N_969,N_921,N_902);
nor U970 (N_970,N_932,N_907);
nor U971 (N_971,N_910,N_922);
nor U972 (N_972,N_904,N_905);
and U973 (N_973,N_912,N_916);
and U974 (N_974,N_937,N_914);
nand U975 (N_975,N_913,N_920);
or U976 (N_976,N_949,N_906);
and U977 (N_977,N_949,N_942);
or U978 (N_978,N_948,N_920);
nor U979 (N_979,N_934,N_920);
nand U980 (N_980,N_916,N_943);
or U981 (N_981,N_935,N_921);
or U982 (N_982,N_935,N_939);
nor U983 (N_983,N_918,N_902);
nor U984 (N_984,N_929,N_902);
and U985 (N_985,N_922,N_921);
nor U986 (N_986,N_926,N_929);
and U987 (N_987,N_945,N_926);
and U988 (N_988,N_917,N_913);
or U989 (N_989,N_916,N_922);
or U990 (N_990,N_904,N_925);
nor U991 (N_991,N_900,N_932);
or U992 (N_992,N_940,N_902);
or U993 (N_993,N_921,N_943);
and U994 (N_994,N_936,N_944);
and U995 (N_995,N_947,N_942);
xor U996 (N_996,N_933,N_920);
nand U997 (N_997,N_941,N_939);
and U998 (N_998,N_906,N_942);
nand U999 (N_999,N_915,N_907);
nor U1000 (N_1000,N_986,N_969);
and U1001 (N_1001,N_982,N_991);
or U1002 (N_1002,N_984,N_999);
and U1003 (N_1003,N_973,N_975);
and U1004 (N_1004,N_997,N_994);
and U1005 (N_1005,N_970,N_988);
nor U1006 (N_1006,N_958,N_962);
nor U1007 (N_1007,N_952,N_977);
nand U1008 (N_1008,N_985,N_992);
or U1009 (N_1009,N_989,N_961);
nand U1010 (N_1010,N_996,N_954);
or U1011 (N_1011,N_957,N_983);
nand U1012 (N_1012,N_968,N_980);
or U1013 (N_1013,N_953,N_998);
nor U1014 (N_1014,N_978,N_987);
nor U1015 (N_1015,N_981,N_964);
and U1016 (N_1016,N_956,N_979);
nor U1017 (N_1017,N_993,N_965);
nand U1018 (N_1018,N_951,N_990);
or U1019 (N_1019,N_966,N_976);
or U1020 (N_1020,N_950,N_967);
or U1021 (N_1021,N_955,N_963);
nand U1022 (N_1022,N_972,N_959);
xor U1023 (N_1023,N_960,N_974);
and U1024 (N_1024,N_995,N_971);
or U1025 (N_1025,N_981,N_973);
nor U1026 (N_1026,N_967,N_988);
nand U1027 (N_1027,N_981,N_994);
nor U1028 (N_1028,N_977,N_956);
nor U1029 (N_1029,N_996,N_976);
nor U1030 (N_1030,N_971,N_988);
or U1031 (N_1031,N_971,N_985);
or U1032 (N_1032,N_958,N_999);
nor U1033 (N_1033,N_995,N_950);
nand U1034 (N_1034,N_975,N_953);
nor U1035 (N_1035,N_993,N_992);
and U1036 (N_1036,N_973,N_961);
or U1037 (N_1037,N_977,N_962);
nor U1038 (N_1038,N_969,N_951);
nand U1039 (N_1039,N_959,N_968);
or U1040 (N_1040,N_965,N_969);
nor U1041 (N_1041,N_956,N_962);
nor U1042 (N_1042,N_976,N_995);
and U1043 (N_1043,N_967,N_971);
and U1044 (N_1044,N_953,N_958);
nor U1045 (N_1045,N_992,N_996);
nand U1046 (N_1046,N_975,N_996);
nor U1047 (N_1047,N_970,N_968);
nand U1048 (N_1048,N_986,N_966);
or U1049 (N_1049,N_966,N_953);
nor U1050 (N_1050,N_1043,N_1003);
nor U1051 (N_1051,N_1029,N_1039);
nor U1052 (N_1052,N_1044,N_1027);
nor U1053 (N_1053,N_1015,N_1005);
or U1054 (N_1054,N_1013,N_1016);
nor U1055 (N_1055,N_1000,N_1012);
nor U1056 (N_1056,N_1035,N_1010);
or U1057 (N_1057,N_1049,N_1046);
and U1058 (N_1058,N_1030,N_1001);
or U1059 (N_1059,N_1002,N_1042);
nand U1060 (N_1060,N_1018,N_1028);
nor U1061 (N_1061,N_1019,N_1040);
nand U1062 (N_1062,N_1034,N_1045);
nor U1063 (N_1063,N_1036,N_1032);
nand U1064 (N_1064,N_1022,N_1007);
nor U1065 (N_1065,N_1041,N_1008);
or U1066 (N_1066,N_1009,N_1017);
nand U1067 (N_1067,N_1047,N_1033);
nand U1068 (N_1068,N_1024,N_1038);
or U1069 (N_1069,N_1023,N_1031);
nand U1070 (N_1070,N_1004,N_1014);
nand U1071 (N_1071,N_1026,N_1011);
or U1072 (N_1072,N_1021,N_1025);
nand U1073 (N_1073,N_1006,N_1048);
or U1074 (N_1074,N_1037,N_1020);
nand U1075 (N_1075,N_1040,N_1044);
nand U1076 (N_1076,N_1031,N_1043);
nand U1077 (N_1077,N_1003,N_1037);
or U1078 (N_1078,N_1042,N_1012);
or U1079 (N_1079,N_1044,N_1037);
and U1080 (N_1080,N_1032,N_1044);
nand U1081 (N_1081,N_1040,N_1027);
or U1082 (N_1082,N_1006,N_1013);
nor U1083 (N_1083,N_1037,N_1045);
nand U1084 (N_1084,N_1021,N_1038);
or U1085 (N_1085,N_1004,N_1033);
nor U1086 (N_1086,N_1012,N_1003);
and U1087 (N_1087,N_1041,N_1028);
nand U1088 (N_1088,N_1029,N_1043);
nand U1089 (N_1089,N_1026,N_1016);
nor U1090 (N_1090,N_1045,N_1040);
nand U1091 (N_1091,N_1039,N_1044);
nor U1092 (N_1092,N_1007,N_1005);
or U1093 (N_1093,N_1049,N_1013);
nand U1094 (N_1094,N_1027,N_1024);
nor U1095 (N_1095,N_1005,N_1026);
or U1096 (N_1096,N_1034,N_1027);
nand U1097 (N_1097,N_1048,N_1001);
and U1098 (N_1098,N_1038,N_1040);
nor U1099 (N_1099,N_1024,N_1042);
nor U1100 (N_1100,N_1072,N_1083);
nor U1101 (N_1101,N_1076,N_1050);
nor U1102 (N_1102,N_1075,N_1089);
and U1103 (N_1103,N_1070,N_1090);
or U1104 (N_1104,N_1097,N_1055);
nor U1105 (N_1105,N_1063,N_1085);
and U1106 (N_1106,N_1093,N_1078);
or U1107 (N_1107,N_1074,N_1054);
and U1108 (N_1108,N_1079,N_1053);
nor U1109 (N_1109,N_1086,N_1052);
or U1110 (N_1110,N_1088,N_1073);
or U1111 (N_1111,N_1060,N_1061);
nor U1112 (N_1112,N_1080,N_1051);
nand U1113 (N_1113,N_1099,N_1098);
or U1114 (N_1114,N_1096,N_1059);
nor U1115 (N_1115,N_1091,N_1077);
and U1116 (N_1116,N_1062,N_1084);
nand U1117 (N_1117,N_1057,N_1095);
or U1118 (N_1118,N_1081,N_1087);
nor U1119 (N_1119,N_1067,N_1066);
and U1120 (N_1120,N_1069,N_1082);
and U1121 (N_1121,N_1071,N_1064);
and U1122 (N_1122,N_1092,N_1065);
nor U1123 (N_1123,N_1094,N_1068);
nor U1124 (N_1124,N_1058,N_1056);
or U1125 (N_1125,N_1050,N_1061);
nor U1126 (N_1126,N_1054,N_1051);
and U1127 (N_1127,N_1057,N_1085);
nand U1128 (N_1128,N_1068,N_1063);
or U1129 (N_1129,N_1052,N_1065);
or U1130 (N_1130,N_1084,N_1081);
or U1131 (N_1131,N_1051,N_1097);
nand U1132 (N_1132,N_1078,N_1058);
nand U1133 (N_1133,N_1061,N_1082);
nor U1134 (N_1134,N_1099,N_1067);
or U1135 (N_1135,N_1082,N_1054);
nor U1136 (N_1136,N_1056,N_1084);
nor U1137 (N_1137,N_1070,N_1063);
nor U1138 (N_1138,N_1093,N_1056);
nand U1139 (N_1139,N_1069,N_1080);
and U1140 (N_1140,N_1066,N_1077);
nor U1141 (N_1141,N_1067,N_1053);
and U1142 (N_1142,N_1054,N_1069);
nand U1143 (N_1143,N_1056,N_1053);
or U1144 (N_1144,N_1050,N_1082);
or U1145 (N_1145,N_1087,N_1080);
nor U1146 (N_1146,N_1064,N_1062);
nand U1147 (N_1147,N_1099,N_1062);
nand U1148 (N_1148,N_1070,N_1058);
and U1149 (N_1149,N_1062,N_1069);
xor U1150 (N_1150,N_1138,N_1144);
nor U1151 (N_1151,N_1116,N_1105);
nand U1152 (N_1152,N_1142,N_1113);
and U1153 (N_1153,N_1140,N_1109);
and U1154 (N_1154,N_1107,N_1118);
or U1155 (N_1155,N_1112,N_1122);
nand U1156 (N_1156,N_1126,N_1119);
nand U1157 (N_1157,N_1124,N_1146);
and U1158 (N_1158,N_1114,N_1100);
and U1159 (N_1159,N_1121,N_1132);
or U1160 (N_1160,N_1106,N_1128);
or U1161 (N_1161,N_1133,N_1103);
or U1162 (N_1162,N_1101,N_1111);
and U1163 (N_1163,N_1125,N_1117);
and U1164 (N_1164,N_1145,N_1147);
and U1165 (N_1165,N_1129,N_1127);
nor U1166 (N_1166,N_1148,N_1130);
and U1167 (N_1167,N_1149,N_1139);
or U1168 (N_1168,N_1110,N_1136);
nor U1169 (N_1169,N_1108,N_1120);
nand U1170 (N_1170,N_1141,N_1134);
or U1171 (N_1171,N_1135,N_1123);
nand U1172 (N_1172,N_1115,N_1102);
and U1173 (N_1173,N_1131,N_1143);
nor U1174 (N_1174,N_1104,N_1137);
and U1175 (N_1175,N_1104,N_1119);
nand U1176 (N_1176,N_1120,N_1119);
nor U1177 (N_1177,N_1105,N_1124);
nor U1178 (N_1178,N_1104,N_1114);
nand U1179 (N_1179,N_1147,N_1109);
and U1180 (N_1180,N_1138,N_1110);
and U1181 (N_1181,N_1120,N_1126);
or U1182 (N_1182,N_1105,N_1122);
nor U1183 (N_1183,N_1137,N_1126);
nand U1184 (N_1184,N_1107,N_1110);
nor U1185 (N_1185,N_1101,N_1142);
and U1186 (N_1186,N_1126,N_1142);
nand U1187 (N_1187,N_1142,N_1139);
nand U1188 (N_1188,N_1141,N_1133);
or U1189 (N_1189,N_1127,N_1131);
nor U1190 (N_1190,N_1110,N_1125);
nor U1191 (N_1191,N_1137,N_1105);
and U1192 (N_1192,N_1132,N_1138);
nand U1193 (N_1193,N_1114,N_1122);
nor U1194 (N_1194,N_1126,N_1102);
nand U1195 (N_1195,N_1113,N_1103);
nor U1196 (N_1196,N_1132,N_1124);
nor U1197 (N_1197,N_1144,N_1149);
nor U1198 (N_1198,N_1121,N_1104);
nand U1199 (N_1199,N_1141,N_1139);
nand U1200 (N_1200,N_1193,N_1164);
xnor U1201 (N_1201,N_1172,N_1195);
or U1202 (N_1202,N_1162,N_1167);
nor U1203 (N_1203,N_1191,N_1197);
nor U1204 (N_1204,N_1198,N_1157);
nand U1205 (N_1205,N_1165,N_1163);
and U1206 (N_1206,N_1196,N_1152);
and U1207 (N_1207,N_1199,N_1153);
and U1208 (N_1208,N_1175,N_1180);
and U1209 (N_1209,N_1187,N_1166);
and U1210 (N_1210,N_1189,N_1183);
and U1211 (N_1211,N_1176,N_1159);
or U1212 (N_1212,N_1190,N_1171);
or U1213 (N_1213,N_1192,N_1185);
or U1214 (N_1214,N_1174,N_1184);
nor U1215 (N_1215,N_1150,N_1177);
nand U1216 (N_1216,N_1169,N_1160);
or U1217 (N_1217,N_1173,N_1194);
or U1218 (N_1218,N_1181,N_1151);
and U1219 (N_1219,N_1182,N_1170);
or U1220 (N_1220,N_1188,N_1168);
nand U1221 (N_1221,N_1186,N_1155);
or U1222 (N_1222,N_1156,N_1154);
or U1223 (N_1223,N_1158,N_1179);
nor U1224 (N_1224,N_1161,N_1178);
and U1225 (N_1225,N_1198,N_1171);
and U1226 (N_1226,N_1169,N_1170);
nand U1227 (N_1227,N_1175,N_1183);
nor U1228 (N_1228,N_1181,N_1188);
nor U1229 (N_1229,N_1196,N_1172);
or U1230 (N_1230,N_1199,N_1181);
and U1231 (N_1231,N_1157,N_1161);
or U1232 (N_1232,N_1161,N_1164);
and U1233 (N_1233,N_1190,N_1196);
nand U1234 (N_1234,N_1162,N_1175);
nand U1235 (N_1235,N_1193,N_1163);
or U1236 (N_1236,N_1158,N_1160);
nor U1237 (N_1237,N_1160,N_1165);
and U1238 (N_1238,N_1193,N_1199);
or U1239 (N_1239,N_1198,N_1151);
nor U1240 (N_1240,N_1160,N_1167);
nor U1241 (N_1241,N_1188,N_1176);
nand U1242 (N_1242,N_1197,N_1158);
nor U1243 (N_1243,N_1151,N_1164);
nand U1244 (N_1244,N_1198,N_1170);
nand U1245 (N_1245,N_1162,N_1155);
and U1246 (N_1246,N_1173,N_1176);
nand U1247 (N_1247,N_1160,N_1177);
nand U1248 (N_1248,N_1180,N_1158);
and U1249 (N_1249,N_1156,N_1188);
or U1250 (N_1250,N_1243,N_1219);
nor U1251 (N_1251,N_1235,N_1214);
nand U1252 (N_1252,N_1241,N_1222);
and U1253 (N_1253,N_1221,N_1249);
nor U1254 (N_1254,N_1203,N_1218);
nand U1255 (N_1255,N_1242,N_1204);
nor U1256 (N_1256,N_1244,N_1237);
nor U1257 (N_1257,N_1232,N_1202);
nand U1258 (N_1258,N_1211,N_1225);
nand U1259 (N_1259,N_1248,N_1239);
nand U1260 (N_1260,N_1247,N_1209);
nor U1261 (N_1261,N_1224,N_1230);
nand U1262 (N_1262,N_1246,N_1217);
nor U1263 (N_1263,N_1220,N_1238);
nand U1264 (N_1264,N_1231,N_1207);
and U1265 (N_1265,N_1229,N_1205);
nor U1266 (N_1266,N_1236,N_1200);
and U1267 (N_1267,N_1210,N_1227);
nor U1268 (N_1268,N_1213,N_1245);
nand U1269 (N_1269,N_1201,N_1212);
and U1270 (N_1270,N_1216,N_1234);
nand U1271 (N_1271,N_1240,N_1206);
or U1272 (N_1272,N_1228,N_1215);
nand U1273 (N_1273,N_1208,N_1233);
nand U1274 (N_1274,N_1226,N_1223);
and U1275 (N_1275,N_1213,N_1235);
and U1276 (N_1276,N_1234,N_1246);
xnor U1277 (N_1277,N_1224,N_1206);
nand U1278 (N_1278,N_1214,N_1234);
or U1279 (N_1279,N_1215,N_1218);
or U1280 (N_1280,N_1207,N_1224);
or U1281 (N_1281,N_1230,N_1210);
nor U1282 (N_1282,N_1203,N_1215);
nand U1283 (N_1283,N_1235,N_1201);
nor U1284 (N_1284,N_1232,N_1210);
and U1285 (N_1285,N_1247,N_1206);
nor U1286 (N_1286,N_1230,N_1225);
or U1287 (N_1287,N_1227,N_1200);
and U1288 (N_1288,N_1216,N_1235);
nor U1289 (N_1289,N_1209,N_1208);
nor U1290 (N_1290,N_1232,N_1216);
nor U1291 (N_1291,N_1234,N_1219);
and U1292 (N_1292,N_1220,N_1201);
and U1293 (N_1293,N_1234,N_1244);
and U1294 (N_1294,N_1238,N_1213);
nor U1295 (N_1295,N_1238,N_1249);
and U1296 (N_1296,N_1219,N_1242);
and U1297 (N_1297,N_1224,N_1220);
nand U1298 (N_1298,N_1209,N_1231);
nand U1299 (N_1299,N_1202,N_1241);
nand U1300 (N_1300,N_1295,N_1251);
nor U1301 (N_1301,N_1273,N_1276);
nand U1302 (N_1302,N_1287,N_1284);
and U1303 (N_1303,N_1282,N_1271);
nand U1304 (N_1304,N_1254,N_1292);
and U1305 (N_1305,N_1285,N_1268);
and U1306 (N_1306,N_1263,N_1293);
or U1307 (N_1307,N_1281,N_1262);
and U1308 (N_1308,N_1264,N_1267);
nor U1309 (N_1309,N_1256,N_1260);
or U1310 (N_1310,N_1257,N_1294);
xor U1311 (N_1311,N_1277,N_1283);
nor U1312 (N_1312,N_1290,N_1299);
nor U1313 (N_1313,N_1253,N_1291);
or U1314 (N_1314,N_1298,N_1269);
and U1315 (N_1315,N_1289,N_1296);
nand U1316 (N_1316,N_1270,N_1266);
nand U1317 (N_1317,N_1252,N_1288);
and U1318 (N_1318,N_1280,N_1265);
and U1319 (N_1319,N_1275,N_1261);
nor U1320 (N_1320,N_1274,N_1259);
nor U1321 (N_1321,N_1297,N_1279);
and U1322 (N_1322,N_1272,N_1255);
nor U1323 (N_1323,N_1258,N_1286);
nor U1324 (N_1324,N_1250,N_1278);
and U1325 (N_1325,N_1263,N_1257);
or U1326 (N_1326,N_1295,N_1294);
nor U1327 (N_1327,N_1277,N_1260);
nor U1328 (N_1328,N_1298,N_1254);
nor U1329 (N_1329,N_1271,N_1268);
and U1330 (N_1330,N_1279,N_1272);
and U1331 (N_1331,N_1273,N_1254);
nand U1332 (N_1332,N_1256,N_1268);
or U1333 (N_1333,N_1295,N_1289);
and U1334 (N_1334,N_1250,N_1258);
nor U1335 (N_1335,N_1265,N_1284);
or U1336 (N_1336,N_1274,N_1270);
nand U1337 (N_1337,N_1298,N_1270);
or U1338 (N_1338,N_1289,N_1256);
and U1339 (N_1339,N_1282,N_1260);
and U1340 (N_1340,N_1284,N_1294);
or U1341 (N_1341,N_1273,N_1270);
and U1342 (N_1342,N_1268,N_1293);
or U1343 (N_1343,N_1252,N_1283);
nand U1344 (N_1344,N_1293,N_1281);
nand U1345 (N_1345,N_1267,N_1263);
nor U1346 (N_1346,N_1263,N_1266);
and U1347 (N_1347,N_1273,N_1278);
or U1348 (N_1348,N_1296,N_1287);
and U1349 (N_1349,N_1292,N_1271);
nor U1350 (N_1350,N_1343,N_1324);
nor U1351 (N_1351,N_1300,N_1331);
nor U1352 (N_1352,N_1339,N_1344);
or U1353 (N_1353,N_1334,N_1308);
nand U1354 (N_1354,N_1314,N_1341);
and U1355 (N_1355,N_1302,N_1313);
nand U1356 (N_1356,N_1316,N_1342);
nor U1357 (N_1357,N_1303,N_1337);
and U1358 (N_1358,N_1330,N_1322);
or U1359 (N_1359,N_1328,N_1307);
and U1360 (N_1360,N_1335,N_1317);
nor U1361 (N_1361,N_1325,N_1327);
nor U1362 (N_1362,N_1301,N_1318);
or U1363 (N_1363,N_1315,N_1348);
nor U1364 (N_1364,N_1323,N_1312);
or U1365 (N_1365,N_1346,N_1345);
or U1366 (N_1366,N_1311,N_1309);
and U1367 (N_1367,N_1326,N_1338);
and U1368 (N_1368,N_1336,N_1347);
nor U1369 (N_1369,N_1340,N_1306);
or U1370 (N_1370,N_1320,N_1319);
and U1371 (N_1371,N_1333,N_1329);
nand U1372 (N_1372,N_1349,N_1310);
and U1373 (N_1373,N_1305,N_1321);
and U1374 (N_1374,N_1304,N_1332);
nand U1375 (N_1375,N_1312,N_1340);
nand U1376 (N_1376,N_1339,N_1308);
and U1377 (N_1377,N_1335,N_1342);
nand U1378 (N_1378,N_1340,N_1303);
nand U1379 (N_1379,N_1345,N_1336);
nand U1380 (N_1380,N_1308,N_1349);
nand U1381 (N_1381,N_1315,N_1330);
xor U1382 (N_1382,N_1311,N_1340);
and U1383 (N_1383,N_1333,N_1307);
or U1384 (N_1384,N_1340,N_1309);
nand U1385 (N_1385,N_1345,N_1303);
or U1386 (N_1386,N_1334,N_1312);
nor U1387 (N_1387,N_1335,N_1314);
or U1388 (N_1388,N_1331,N_1326);
nand U1389 (N_1389,N_1302,N_1330);
nor U1390 (N_1390,N_1301,N_1347);
nor U1391 (N_1391,N_1332,N_1320);
and U1392 (N_1392,N_1331,N_1304);
nor U1393 (N_1393,N_1337,N_1329);
or U1394 (N_1394,N_1331,N_1346);
nor U1395 (N_1395,N_1328,N_1341);
or U1396 (N_1396,N_1302,N_1323);
nand U1397 (N_1397,N_1339,N_1310);
or U1398 (N_1398,N_1319,N_1339);
and U1399 (N_1399,N_1323,N_1314);
or U1400 (N_1400,N_1388,N_1376);
nor U1401 (N_1401,N_1386,N_1372);
nand U1402 (N_1402,N_1351,N_1393);
nand U1403 (N_1403,N_1390,N_1382);
nor U1404 (N_1404,N_1368,N_1354);
or U1405 (N_1405,N_1358,N_1365);
or U1406 (N_1406,N_1352,N_1392);
nand U1407 (N_1407,N_1385,N_1384);
nor U1408 (N_1408,N_1387,N_1366);
nor U1409 (N_1409,N_1378,N_1380);
nor U1410 (N_1410,N_1364,N_1396);
nand U1411 (N_1411,N_1359,N_1398);
nand U1412 (N_1412,N_1383,N_1375);
and U1413 (N_1413,N_1371,N_1379);
nand U1414 (N_1414,N_1374,N_1367);
nand U1415 (N_1415,N_1361,N_1350);
nor U1416 (N_1416,N_1399,N_1391);
nor U1417 (N_1417,N_1397,N_1394);
nand U1418 (N_1418,N_1353,N_1356);
nand U1419 (N_1419,N_1355,N_1373);
nand U1420 (N_1420,N_1395,N_1377);
or U1421 (N_1421,N_1389,N_1360);
nor U1422 (N_1422,N_1370,N_1362);
or U1423 (N_1423,N_1357,N_1381);
nor U1424 (N_1424,N_1363,N_1369);
and U1425 (N_1425,N_1392,N_1372);
xnor U1426 (N_1426,N_1382,N_1379);
nor U1427 (N_1427,N_1378,N_1377);
nand U1428 (N_1428,N_1360,N_1397);
nor U1429 (N_1429,N_1358,N_1388);
and U1430 (N_1430,N_1376,N_1354);
nand U1431 (N_1431,N_1385,N_1399);
or U1432 (N_1432,N_1365,N_1398);
and U1433 (N_1433,N_1390,N_1351);
or U1434 (N_1434,N_1369,N_1370);
and U1435 (N_1435,N_1371,N_1385);
nand U1436 (N_1436,N_1354,N_1353);
nor U1437 (N_1437,N_1395,N_1352);
or U1438 (N_1438,N_1399,N_1392);
and U1439 (N_1439,N_1399,N_1364);
nor U1440 (N_1440,N_1358,N_1354);
and U1441 (N_1441,N_1350,N_1373);
and U1442 (N_1442,N_1382,N_1362);
and U1443 (N_1443,N_1360,N_1357);
nand U1444 (N_1444,N_1368,N_1393);
or U1445 (N_1445,N_1390,N_1393);
or U1446 (N_1446,N_1391,N_1359);
or U1447 (N_1447,N_1385,N_1375);
nor U1448 (N_1448,N_1363,N_1389);
or U1449 (N_1449,N_1362,N_1357);
nor U1450 (N_1450,N_1422,N_1440);
or U1451 (N_1451,N_1447,N_1418);
and U1452 (N_1452,N_1401,N_1429);
nand U1453 (N_1453,N_1416,N_1432);
nor U1454 (N_1454,N_1424,N_1435);
nand U1455 (N_1455,N_1439,N_1430);
nor U1456 (N_1456,N_1417,N_1449);
nor U1457 (N_1457,N_1414,N_1404);
nor U1458 (N_1458,N_1442,N_1433);
nor U1459 (N_1459,N_1431,N_1410);
and U1460 (N_1460,N_1437,N_1415);
and U1461 (N_1461,N_1423,N_1443);
nor U1462 (N_1462,N_1405,N_1408);
nand U1463 (N_1463,N_1438,N_1409);
xnor U1464 (N_1464,N_1434,N_1427);
nand U1465 (N_1465,N_1436,N_1448);
nor U1466 (N_1466,N_1446,N_1419);
nand U1467 (N_1467,N_1403,N_1420);
and U1468 (N_1468,N_1407,N_1406);
or U1469 (N_1469,N_1445,N_1428);
and U1470 (N_1470,N_1441,N_1402);
nor U1471 (N_1471,N_1425,N_1421);
nand U1472 (N_1472,N_1400,N_1412);
or U1473 (N_1473,N_1413,N_1411);
nand U1474 (N_1474,N_1444,N_1426);
nor U1475 (N_1475,N_1446,N_1437);
nor U1476 (N_1476,N_1408,N_1407);
nor U1477 (N_1477,N_1426,N_1446);
or U1478 (N_1478,N_1422,N_1431);
or U1479 (N_1479,N_1416,N_1441);
nor U1480 (N_1480,N_1439,N_1410);
nand U1481 (N_1481,N_1437,N_1435);
nand U1482 (N_1482,N_1442,N_1409);
or U1483 (N_1483,N_1430,N_1431);
or U1484 (N_1484,N_1419,N_1428);
nor U1485 (N_1485,N_1443,N_1416);
and U1486 (N_1486,N_1406,N_1410);
or U1487 (N_1487,N_1403,N_1439);
nand U1488 (N_1488,N_1438,N_1414);
nor U1489 (N_1489,N_1441,N_1433);
or U1490 (N_1490,N_1419,N_1416);
nand U1491 (N_1491,N_1405,N_1432);
or U1492 (N_1492,N_1405,N_1426);
nand U1493 (N_1493,N_1412,N_1417);
or U1494 (N_1494,N_1409,N_1437);
nor U1495 (N_1495,N_1434,N_1403);
nor U1496 (N_1496,N_1414,N_1443);
nor U1497 (N_1497,N_1423,N_1404);
and U1498 (N_1498,N_1435,N_1434);
or U1499 (N_1499,N_1421,N_1422);
and U1500 (N_1500,N_1483,N_1496);
or U1501 (N_1501,N_1455,N_1450);
or U1502 (N_1502,N_1468,N_1475);
nand U1503 (N_1503,N_1453,N_1479);
and U1504 (N_1504,N_1460,N_1457);
nand U1505 (N_1505,N_1489,N_1497);
or U1506 (N_1506,N_1480,N_1485);
and U1507 (N_1507,N_1462,N_1484);
or U1508 (N_1508,N_1463,N_1456);
nand U1509 (N_1509,N_1474,N_1490);
and U1510 (N_1510,N_1470,N_1459);
nor U1511 (N_1511,N_1488,N_1465);
nand U1512 (N_1512,N_1478,N_1466);
nor U1513 (N_1513,N_1494,N_1476);
nor U1514 (N_1514,N_1491,N_1486);
nor U1515 (N_1515,N_1495,N_1493);
nand U1516 (N_1516,N_1477,N_1498);
nand U1517 (N_1517,N_1472,N_1482);
or U1518 (N_1518,N_1499,N_1467);
and U1519 (N_1519,N_1487,N_1452);
xor U1520 (N_1520,N_1492,N_1461);
and U1521 (N_1521,N_1451,N_1469);
and U1522 (N_1522,N_1454,N_1473);
and U1523 (N_1523,N_1481,N_1471);
or U1524 (N_1524,N_1458,N_1464);
nand U1525 (N_1525,N_1480,N_1498);
and U1526 (N_1526,N_1462,N_1471);
or U1527 (N_1527,N_1490,N_1465);
nand U1528 (N_1528,N_1454,N_1459);
nand U1529 (N_1529,N_1468,N_1450);
and U1530 (N_1530,N_1491,N_1454);
and U1531 (N_1531,N_1473,N_1450);
or U1532 (N_1532,N_1491,N_1465);
nor U1533 (N_1533,N_1495,N_1455);
and U1534 (N_1534,N_1494,N_1485);
nor U1535 (N_1535,N_1458,N_1467);
and U1536 (N_1536,N_1451,N_1485);
or U1537 (N_1537,N_1478,N_1485);
and U1538 (N_1538,N_1469,N_1489);
nand U1539 (N_1539,N_1474,N_1457);
nor U1540 (N_1540,N_1497,N_1493);
and U1541 (N_1541,N_1470,N_1469);
and U1542 (N_1542,N_1465,N_1476);
and U1543 (N_1543,N_1487,N_1482);
or U1544 (N_1544,N_1466,N_1455);
and U1545 (N_1545,N_1495,N_1491);
nand U1546 (N_1546,N_1453,N_1452);
or U1547 (N_1547,N_1480,N_1496);
or U1548 (N_1548,N_1459,N_1481);
or U1549 (N_1549,N_1489,N_1499);
nor U1550 (N_1550,N_1519,N_1545);
nor U1551 (N_1551,N_1511,N_1520);
and U1552 (N_1552,N_1508,N_1506);
nor U1553 (N_1553,N_1532,N_1528);
or U1554 (N_1554,N_1549,N_1515);
nand U1555 (N_1555,N_1529,N_1524);
nand U1556 (N_1556,N_1546,N_1518);
nor U1557 (N_1557,N_1504,N_1512);
or U1558 (N_1558,N_1503,N_1509);
or U1559 (N_1559,N_1548,N_1522);
and U1560 (N_1560,N_1516,N_1542);
and U1561 (N_1561,N_1526,N_1537);
or U1562 (N_1562,N_1523,N_1538);
and U1563 (N_1563,N_1525,N_1534);
or U1564 (N_1564,N_1527,N_1501);
nand U1565 (N_1565,N_1535,N_1513);
or U1566 (N_1566,N_1505,N_1541);
nor U1567 (N_1567,N_1514,N_1521);
or U1568 (N_1568,N_1530,N_1543);
and U1569 (N_1569,N_1507,N_1533);
nand U1570 (N_1570,N_1531,N_1500);
and U1571 (N_1571,N_1544,N_1539);
and U1572 (N_1572,N_1536,N_1510);
and U1573 (N_1573,N_1547,N_1502);
nand U1574 (N_1574,N_1517,N_1540);
and U1575 (N_1575,N_1504,N_1548);
and U1576 (N_1576,N_1519,N_1544);
nand U1577 (N_1577,N_1516,N_1512);
nor U1578 (N_1578,N_1549,N_1547);
and U1579 (N_1579,N_1530,N_1522);
or U1580 (N_1580,N_1538,N_1512);
nand U1581 (N_1581,N_1513,N_1532);
or U1582 (N_1582,N_1501,N_1508);
nor U1583 (N_1583,N_1538,N_1511);
and U1584 (N_1584,N_1500,N_1512);
or U1585 (N_1585,N_1504,N_1508);
nor U1586 (N_1586,N_1515,N_1507);
and U1587 (N_1587,N_1532,N_1543);
nor U1588 (N_1588,N_1523,N_1507);
or U1589 (N_1589,N_1546,N_1506);
nor U1590 (N_1590,N_1542,N_1548);
or U1591 (N_1591,N_1521,N_1548);
or U1592 (N_1592,N_1528,N_1529);
nor U1593 (N_1593,N_1506,N_1539);
nand U1594 (N_1594,N_1504,N_1537);
and U1595 (N_1595,N_1533,N_1527);
nor U1596 (N_1596,N_1521,N_1512);
or U1597 (N_1597,N_1516,N_1523);
nor U1598 (N_1598,N_1535,N_1538);
nor U1599 (N_1599,N_1543,N_1502);
or U1600 (N_1600,N_1574,N_1558);
or U1601 (N_1601,N_1592,N_1555);
nor U1602 (N_1602,N_1564,N_1568);
or U1603 (N_1603,N_1561,N_1552);
or U1604 (N_1604,N_1593,N_1562);
and U1605 (N_1605,N_1553,N_1569);
nor U1606 (N_1606,N_1578,N_1567);
nor U1607 (N_1607,N_1559,N_1584);
and U1608 (N_1608,N_1582,N_1576);
xnor U1609 (N_1609,N_1557,N_1589);
nand U1610 (N_1610,N_1590,N_1566);
nand U1611 (N_1611,N_1595,N_1563);
nand U1612 (N_1612,N_1583,N_1575);
or U1613 (N_1613,N_1598,N_1565);
and U1614 (N_1614,N_1580,N_1570);
or U1615 (N_1615,N_1586,N_1551);
and U1616 (N_1616,N_1588,N_1573);
nand U1617 (N_1617,N_1560,N_1571);
nor U1618 (N_1618,N_1577,N_1579);
nor U1619 (N_1619,N_1556,N_1597);
or U1620 (N_1620,N_1591,N_1572);
nand U1621 (N_1621,N_1587,N_1596);
and U1622 (N_1622,N_1550,N_1599);
or U1623 (N_1623,N_1594,N_1585);
and U1624 (N_1624,N_1581,N_1554);
nor U1625 (N_1625,N_1571,N_1588);
or U1626 (N_1626,N_1566,N_1551);
nand U1627 (N_1627,N_1575,N_1555);
and U1628 (N_1628,N_1597,N_1576);
and U1629 (N_1629,N_1573,N_1597);
or U1630 (N_1630,N_1584,N_1597);
or U1631 (N_1631,N_1570,N_1558);
and U1632 (N_1632,N_1575,N_1574);
nand U1633 (N_1633,N_1594,N_1591);
and U1634 (N_1634,N_1564,N_1566);
nor U1635 (N_1635,N_1558,N_1552);
nor U1636 (N_1636,N_1550,N_1568);
nor U1637 (N_1637,N_1569,N_1576);
and U1638 (N_1638,N_1593,N_1563);
nor U1639 (N_1639,N_1555,N_1586);
nor U1640 (N_1640,N_1569,N_1554);
nand U1641 (N_1641,N_1569,N_1592);
or U1642 (N_1642,N_1563,N_1561);
or U1643 (N_1643,N_1574,N_1551);
nor U1644 (N_1644,N_1563,N_1594);
nor U1645 (N_1645,N_1581,N_1556);
and U1646 (N_1646,N_1596,N_1559);
nor U1647 (N_1647,N_1599,N_1558);
nand U1648 (N_1648,N_1554,N_1560);
or U1649 (N_1649,N_1589,N_1593);
nand U1650 (N_1650,N_1621,N_1644);
or U1651 (N_1651,N_1616,N_1626);
and U1652 (N_1652,N_1643,N_1604);
or U1653 (N_1653,N_1649,N_1625);
nor U1654 (N_1654,N_1601,N_1628);
nand U1655 (N_1655,N_1634,N_1612);
nor U1656 (N_1656,N_1605,N_1638);
nor U1657 (N_1657,N_1631,N_1617);
nand U1658 (N_1658,N_1608,N_1613);
nand U1659 (N_1659,N_1624,N_1619);
or U1660 (N_1660,N_1633,N_1606);
nor U1661 (N_1661,N_1636,N_1620);
and U1662 (N_1662,N_1647,N_1609);
and U1663 (N_1663,N_1641,N_1629);
or U1664 (N_1664,N_1611,N_1614);
or U1665 (N_1665,N_1610,N_1603);
or U1666 (N_1666,N_1645,N_1642);
and U1667 (N_1667,N_1618,N_1632);
nor U1668 (N_1668,N_1637,N_1640);
nand U1669 (N_1669,N_1622,N_1623);
and U1670 (N_1670,N_1607,N_1600);
nand U1671 (N_1671,N_1648,N_1639);
or U1672 (N_1672,N_1627,N_1630);
nor U1673 (N_1673,N_1646,N_1615);
and U1674 (N_1674,N_1635,N_1602);
nor U1675 (N_1675,N_1602,N_1608);
or U1676 (N_1676,N_1648,N_1615);
and U1677 (N_1677,N_1614,N_1642);
nand U1678 (N_1678,N_1617,N_1636);
nand U1679 (N_1679,N_1613,N_1614);
or U1680 (N_1680,N_1623,N_1613);
and U1681 (N_1681,N_1606,N_1641);
nor U1682 (N_1682,N_1621,N_1600);
nor U1683 (N_1683,N_1601,N_1632);
nand U1684 (N_1684,N_1643,N_1633);
or U1685 (N_1685,N_1622,N_1641);
or U1686 (N_1686,N_1613,N_1627);
and U1687 (N_1687,N_1634,N_1606);
nand U1688 (N_1688,N_1646,N_1603);
or U1689 (N_1689,N_1645,N_1603);
nand U1690 (N_1690,N_1624,N_1640);
nand U1691 (N_1691,N_1610,N_1609);
or U1692 (N_1692,N_1643,N_1628);
and U1693 (N_1693,N_1608,N_1633);
or U1694 (N_1694,N_1621,N_1636);
nand U1695 (N_1695,N_1639,N_1617);
and U1696 (N_1696,N_1624,N_1607);
nand U1697 (N_1697,N_1629,N_1606);
nor U1698 (N_1698,N_1644,N_1613);
or U1699 (N_1699,N_1608,N_1618);
or U1700 (N_1700,N_1650,N_1671);
or U1701 (N_1701,N_1688,N_1662);
nor U1702 (N_1702,N_1687,N_1680);
nand U1703 (N_1703,N_1677,N_1695);
nor U1704 (N_1704,N_1673,N_1692);
nand U1705 (N_1705,N_1653,N_1661);
and U1706 (N_1706,N_1682,N_1693);
or U1707 (N_1707,N_1676,N_1660);
nand U1708 (N_1708,N_1669,N_1665);
nor U1709 (N_1709,N_1690,N_1694);
or U1710 (N_1710,N_1672,N_1684);
nor U1711 (N_1711,N_1670,N_1658);
nand U1712 (N_1712,N_1667,N_1675);
nor U1713 (N_1713,N_1654,N_1664);
nor U1714 (N_1714,N_1699,N_1652);
or U1715 (N_1715,N_1651,N_1666);
or U1716 (N_1716,N_1698,N_1663);
and U1717 (N_1717,N_1685,N_1686);
and U1718 (N_1718,N_1655,N_1659);
and U1719 (N_1719,N_1696,N_1697);
nand U1720 (N_1720,N_1681,N_1657);
nor U1721 (N_1721,N_1656,N_1674);
nor U1722 (N_1722,N_1683,N_1679);
nand U1723 (N_1723,N_1668,N_1678);
xnor U1724 (N_1724,N_1689,N_1691);
nand U1725 (N_1725,N_1698,N_1678);
and U1726 (N_1726,N_1683,N_1670);
and U1727 (N_1727,N_1685,N_1653);
nor U1728 (N_1728,N_1699,N_1684);
and U1729 (N_1729,N_1692,N_1658);
or U1730 (N_1730,N_1684,N_1667);
and U1731 (N_1731,N_1660,N_1670);
and U1732 (N_1732,N_1674,N_1653);
or U1733 (N_1733,N_1666,N_1660);
or U1734 (N_1734,N_1681,N_1666);
and U1735 (N_1735,N_1656,N_1697);
and U1736 (N_1736,N_1698,N_1691);
nor U1737 (N_1737,N_1650,N_1658);
nand U1738 (N_1738,N_1691,N_1659);
and U1739 (N_1739,N_1670,N_1679);
nor U1740 (N_1740,N_1653,N_1681);
nor U1741 (N_1741,N_1684,N_1681);
nor U1742 (N_1742,N_1667,N_1687);
or U1743 (N_1743,N_1699,N_1675);
or U1744 (N_1744,N_1672,N_1661);
and U1745 (N_1745,N_1688,N_1654);
and U1746 (N_1746,N_1685,N_1662);
xnor U1747 (N_1747,N_1698,N_1688);
or U1748 (N_1748,N_1650,N_1674);
nand U1749 (N_1749,N_1686,N_1689);
or U1750 (N_1750,N_1743,N_1737);
and U1751 (N_1751,N_1733,N_1701);
nor U1752 (N_1752,N_1727,N_1717);
and U1753 (N_1753,N_1726,N_1719);
and U1754 (N_1754,N_1716,N_1747);
and U1755 (N_1755,N_1721,N_1725);
or U1756 (N_1756,N_1744,N_1713);
nor U1757 (N_1757,N_1706,N_1748);
or U1758 (N_1758,N_1711,N_1742);
nand U1759 (N_1759,N_1745,N_1720);
nor U1760 (N_1760,N_1715,N_1749);
or U1761 (N_1761,N_1735,N_1731);
nand U1762 (N_1762,N_1730,N_1712);
nand U1763 (N_1763,N_1718,N_1710);
nand U1764 (N_1764,N_1702,N_1707);
and U1765 (N_1765,N_1714,N_1736);
or U1766 (N_1766,N_1724,N_1728);
nor U1767 (N_1767,N_1703,N_1708);
nor U1768 (N_1768,N_1729,N_1746);
nor U1769 (N_1769,N_1709,N_1700);
nor U1770 (N_1770,N_1722,N_1739);
and U1771 (N_1771,N_1738,N_1723);
or U1772 (N_1772,N_1732,N_1740);
or U1773 (N_1773,N_1741,N_1734);
nand U1774 (N_1774,N_1704,N_1705);
nand U1775 (N_1775,N_1721,N_1729);
nor U1776 (N_1776,N_1748,N_1740);
or U1777 (N_1777,N_1732,N_1708);
nor U1778 (N_1778,N_1727,N_1723);
xor U1779 (N_1779,N_1732,N_1711);
or U1780 (N_1780,N_1739,N_1745);
nor U1781 (N_1781,N_1731,N_1745);
and U1782 (N_1782,N_1716,N_1748);
and U1783 (N_1783,N_1744,N_1708);
and U1784 (N_1784,N_1706,N_1716);
nor U1785 (N_1785,N_1705,N_1735);
nor U1786 (N_1786,N_1744,N_1709);
nand U1787 (N_1787,N_1705,N_1731);
nand U1788 (N_1788,N_1708,N_1746);
and U1789 (N_1789,N_1720,N_1709);
nand U1790 (N_1790,N_1730,N_1706);
and U1791 (N_1791,N_1726,N_1717);
or U1792 (N_1792,N_1748,N_1739);
nor U1793 (N_1793,N_1705,N_1737);
nand U1794 (N_1794,N_1702,N_1739);
and U1795 (N_1795,N_1730,N_1738);
nand U1796 (N_1796,N_1744,N_1723);
nand U1797 (N_1797,N_1730,N_1726);
nand U1798 (N_1798,N_1732,N_1744);
nand U1799 (N_1799,N_1747,N_1711);
and U1800 (N_1800,N_1755,N_1775);
nor U1801 (N_1801,N_1783,N_1779);
and U1802 (N_1802,N_1794,N_1763);
and U1803 (N_1803,N_1776,N_1757);
nor U1804 (N_1804,N_1796,N_1784);
nand U1805 (N_1805,N_1765,N_1770);
and U1806 (N_1806,N_1781,N_1786);
nand U1807 (N_1807,N_1785,N_1759);
nor U1808 (N_1808,N_1778,N_1790);
nor U1809 (N_1809,N_1792,N_1780);
and U1810 (N_1810,N_1750,N_1764);
nor U1811 (N_1811,N_1753,N_1751);
nand U1812 (N_1812,N_1752,N_1799);
or U1813 (N_1813,N_1771,N_1767);
nor U1814 (N_1814,N_1774,N_1787);
nor U1815 (N_1815,N_1766,N_1797);
nor U1816 (N_1816,N_1760,N_1782);
nor U1817 (N_1817,N_1793,N_1788);
nor U1818 (N_1818,N_1762,N_1769);
and U1819 (N_1819,N_1772,N_1761);
nor U1820 (N_1820,N_1756,N_1777);
and U1821 (N_1821,N_1768,N_1754);
and U1822 (N_1822,N_1789,N_1795);
or U1823 (N_1823,N_1798,N_1758);
nor U1824 (N_1824,N_1773,N_1791);
nor U1825 (N_1825,N_1758,N_1770);
nand U1826 (N_1826,N_1781,N_1768);
nand U1827 (N_1827,N_1780,N_1760);
nand U1828 (N_1828,N_1769,N_1795);
and U1829 (N_1829,N_1772,N_1796);
and U1830 (N_1830,N_1777,N_1772);
or U1831 (N_1831,N_1772,N_1771);
and U1832 (N_1832,N_1796,N_1783);
or U1833 (N_1833,N_1778,N_1792);
nand U1834 (N_1834,N_1784,N_1754);
or U1835 (N_1835,N_1764,N_1780);
nand U1836 (N_1836,N_1752,N_1768);
nand U1837 (N_1837,N_1793,N_1782);
or U1838 (N_1838,N_1786,N_1787);
and U1839 (N_1839,N_1758,N_1752);
nor U1840 (N_1840,N_1762,N_1760);
nor U1841 (N_1841,N_1761,N_1787);
nor U1842 (N_1842,N_1756,N_1788);
and U1843 (N_1843,N_1764,N_1785);
nand U1844 (N_1844,N_1774,N_1752);
and U1845 (N_1845,N_1759,N_1762);
nor U1846 (N_1846,N_1762,N_1755);
or U1847 (N_1847,N_1753,N_1772);
and U1848 (N_1848,N_1795,N_1773);
nor U1849 (N_1849,N_1767,N_1783);
nor U1850 (N_1850,N_1808,N_1839);
nor U1851 (N_1851,N_1847,N_1819);
nand U1852 (N_1852,N_1811,N_1832);
and U1853 (N_1853,N_1807,N_1800);
or U1854 (N_1854,N_1843,N_1828);
or U1855 (N_1855,N_1815,N_1810);
nor U1856 (N_1856,N_1806,N_1809);
nor U1857 (N_1857,N_1846,N_1816);
nand U1858 (N_1858,N_1830,N_1801);
or U1859 (N_1859,N_1803,N_1829);
nor U1860 (N_1860,N_1841,N_1833);
nor U1861 (N_1861,N_1838,N_1823);
or U1862 (N_1862,N_1831,N_1804);
nor U1863 (N_1863,N_1812,N_1814);
or U1864 (N_1864,N_1840,N_1844);
and U1865 (N_1865,N_1834,N_1824);
nand U1866 (N_1866,N_1826,N_1805);
nor U1867 (N_1867,N_1820,N_1825);
nand U1868 (N_1868,N_1835,N_1849);
or U1869 (N_1869,N_1822,N_1836);
or U1870 (N_1870,N_1818,N_1802);
or U1871 (N_1871,N_1817,N_1848);
nand U1872 (N_1872,N_1842,N_1813);
nand U1873 (N_1873,N_1845,N_1837);
or U1874 (N_1874,N_1827,N_1821);
and U1875 (N_1875,N_1826,N_1801);
or U1876 (N_1876,N_1817,N_1823);
nand U1877 (N_1877,N_1830,N_1843);
nand U1878 (N_1878,N_1819,N_1830);
nand U1879 (N_1879,N_1837,N_1846);
or U1880 (N_1880,N_1823,N_1803);
and U1881 (N_1881,N_1821,N_1833);
and U1882 (N_1882,N_1802,N_1834);
nand U1883 (N_1883,N_1813,N_1841);
or U1884 (N_1884,N_1822,N_1813);
or U1885 (N_1885,N_1818,N_1833);
nor U1886 (N_1886,N_1841,N_1808);
nor U1887 (N_1887,N_1810,N_1831);
nand U1888 (N_1888,N_1844,N_1841);
and U1889 (N_1889,N_1824,N_1806);
and U1890 (N_1890,N_1845,N_1836);
or U1891 (N_1891,N_1823,N_1802);
and U1892 (N_1892,N_1811,N_1834);
or U1893 (N_1893,N_1806,N_1823);
nor U1894 (N_1894,N_1826,N_1806);
xor U1895 (N_1895,N_1833,N_1801);
nand U1896 (N_1896,N_1808,N_1849);
and U1897 (N_1897,N_1816,N_1827);
or U1898 (N_1898,N_1810,N_1841);
nand U1899 (N_1899,N_1840,N_1836);
and U1900 (N_1900,N_1885,N_1887);
nand U1901 (N_1901,N_1857,N_1896);
nand U1902 (N_1902,N_1897,N_1880);
and U1903 (N_1903,N_1858,N_1851);
and U1904 (N_1904,N_1876,N_1863);
nand U1905 (N_1905,N_1862,N_1854);
or U1906 (N_1906,N_1893,N_1861);
and U1907 (N_1907,N_1875,N_1869);
or U1908 (N_1908,N_1855,N_1879);
or U1909 (N_1909,N_1882,N_1874);
and U1910 (N_1910,N_1873,N_1889);
and U1911 (N_1911,N_1868,N_1894);
nor U1912 (N_1912,N_1860,N_1891);
nor U1913 (N_1913,N_1850,N_1865);
and U1914 (N_1914,N_1856,N_1852);
or U1915 (N_1915,N_1872,N_1864);
and U1916 (N_1916,N_1877,N_1892);
nand U1917 (N_1917,N_1871,N_1881);
nand U1918 (N_1918,N_1898,N_1859);
nor U1919 (N_1919,N_1886,N_1853);
nand U1920 (N_1920,N_1895,N_1888);
nand U1921 (N_1921,N_1870,N_1866);
or U1922 (N_1922,N_1890,N_1899);
nor U1923 (N_1923,N_1867,N_1878);
and U1924 (N_1924,N_1884,N_1883);
and U1925 (N_1925,N_1893,N_1890);
nor U1926 (N_1926,N_1893,N_1867);
or U1927 (N_1927,N_1857,N_1855);
and U1928 (N_1928,N_1871,N_1859);
and U1929 (N_1929,N_1888,N_1893);
and U1930 (N_1930,N_1895,N_1855);
nor U1931 (N_1931,N_1880,N_1857);
and U1932 (N_1932,N_1874,N_1857);
nand U1933 (N_1933,N_1857,N_1883);
or U1934 (N_1934,N_1867,N_1876);
nor U1935 (N_1935,N_1880,N_1875);
and U1936 (N_1936,N_1896,N_1895);
or U1937 (N_1937,N_1887,N_1872);
nor U1938 (N_1938,N_1862,N_1864);
and U1939 (N_1939,N_1891,N_1863);
or U1940 (N_1940,N_1859,N_1875);
nor U1941 (N_1941,N_1884,N_1866);
nand U1942 (N_1942,N_1876,N_1882);
nor U1943 (N_1943,N_1860,N_1883);
or U1944 (N_1944,N_1888,N_1856);
or U1945 (N_1945,N_1867,N_1879);
or U1946 (N_1946,N_1877,N_1899);
or U1947 (N_1947,N_1878,N_1875);
and U1948 (N_1948,N_1864,N_1893);
nand U1949 (N_1949,N_1871,N_1867);
or U1950 (N_1950,N_1913,N_1930);
and U1951 (N_1951,N_1904,N_1941);
and U1952 (N_1952,N_1938,N_1918);
nand U1953 (N_1953,N_1916,N_1946);
or U1954 (N_1954,N_1909,N_1933);
nor U1955 (N_1955,N_1902,N_1925);
or U1956 (N_1956,N_1935,N_1943);
nor U1957 (N_1957,N_1937,N_1940);
and U1958 (N_1958,N_1906,N_1949);
xnor U1959 (N_1959,N_1936,N_1920);
or U1960 (N_1960,N_1942,N_1929);
nand U1961 (N_1961,N_1934,N_1928);
or U1962 (N_1962,N_1901,N_1915);
and U1963 (N_1963,N_1944,N_1932);
nor U1964 (N_1964,N_1945,N_1931);
nor U1965 (N_1965,N_1917,N_1927);
nand U1966 (N_1966,N_1922,N_1912);
nor U1967 (N_1967,N_1926,N_1905);
nand U1968 (N_1968,N_1924,N_1903);
nand U1969 (N_1969,N_1910,N_1947);
nor U1970 (N_1970,N_1914,N_1939);
and U1971 (N_1971,N_1919,N_1923);
and U1972 (N_1972,N_1900,N_1948);
nand U1973 (N_1973,N_1908,N_1911);
nor U1974 (N_1974,N_1921,N_1907);
nor U1975 (N_1975,N_1948,N_1918);
and U1976 (N_1976,N_1948,N_1922);
nor U1977 (N_1977,N_1917,N_1926);
or U1978 (N_1978,N_1947,N_1927);
nand U1979 (N_1979,N_1908,N_1921);
and U1980 (N_1980,N_1916,N_1939);
and U1981 (N_1981,N_1943,N_1921);
or U1982 (N_1982,N_1918,N_1932);
and U1983 (N_1983,N_1918,N_1904);
and U1984 (N_1984,N_1924,N_1901);
nor U1985 (N_1985,N_1940,N_1910);
or U1986 (N_1986,N_1932,N_1936);
or U1987 (N_1987,N_1902,N_1936);
or U1988 (N_1988,N_1900,N_1922);
nor U1989 (N_1989,N_1938,N_1949);
and U1990 (N_1990,N_1942,N_1916);
nor U1991 (N_1991,N_1925,N_1908);
nor U1992 (N_1992,N_1937,N_1920);
or U1993 (N_1993,N_1933,N_1924);
nand U1994 (N_1994,N_1902,N_1912);
nand U1995 (N_1995,N_1938,N_1924);
nor U1996 (N_1996,N_1923,N_1916);
and U1997 (N_1997,N_1935,N_1913);
or U1998 (N_1998,N_1903,N_1926);
nand U1999 (N_1999,N_1940,N_1941);
and U2000 (N_2000,N_1988,N_1974);
or U2001 (N_2001,N_1957,N_1990);
and U2002 (N_2002,N_1994,N_1968);
nand U2003 (N_2003,N_1984,N_1965);
nor U2004 (N_2004,N_1995,N_1973);
and U2005 (N_2005,N_1999,N_1989);
and U2006 (N_2006,N_1971,N_1952);
and U2007 (N_2007,N_1963,N_1983);
nand U2008 (N_2008,N_1956,N_1985);
and U2009 (N_2009,N_1964,N_1958);
nor U2010 (N_2010,N_1996,N_1993);
nand U2011 (N_2011,N_1976,N_1992);
or U2012 (N_2012,N_1981,N_1991);
nor U2013 (N_2013,N_1959,N_1953);
nand U2014 (N_2014,N_1950,N_1998);
nand U2015 (N_2015,N_1951,N_1972);
or U2016 (N_2016,N_1982,N_1977);
and U2017 (N_2017,N_1967,N_1960);
nor U2018 (N_2018,N_1955,N_1969);
nor U2019 (N_2019,N_1970,N_1962);
or U2020 (N_2020,N_1966,N_1954);
and U2021 (N_2021,N_1961,N_1980);
nand U2022 (N_2022,N_1986,N_1975);
nand U2023 (N_2023,N_1979,N_1997);
nand U2024 (N_2024,N_1987,N_1978);
and U2025 (N_2025,N_1980,N_1999);
nand U2026 (N_2026,N_1962,N_1957);
nand U2027 (N_2027,N_1995,N_1987);
nand U2028 (N_2028,N_1981,N_1950);
nand U2029 (N_2029,N_1997,N_1999);
and U2030 (N_2030,N_1999,N_1973);
and U2031 (N_2031,N_1976,N_1964);
nand U2032 (N_2032,N_1969,N_1982);
or U2033 (N_2033,N_1958,N_1973);
and U2034 (N_2034,N_1951,N_1950);
nand U2035 (N_2035,N_1974,N_1975);
nand U2036 (N_2036,N_1999,N_1993);
nand U2037 (N_2037,N_1989,N_1998);
nand U2038 (N_2038,N_1987,N_1956);
or U2039 (N_2039,N_1964,N_1991);
xnor U2040 (N_2040,N_1952,N_1967);
nand U2041 (N_2041,N_1969,N_1964);
nand U2042 (N_2042,N_1970,N_1974);
or U2043 (N_2043,N_1973,N_1970);
nand U2044 (N_2044,N_1976,N_1953);
and U2045 (N_2045,N_1978,N_1992);
and U2046 (N_2046,N_1950,N_1992);
or U2047 (N_2047,N_1988,N_1953);
or U2048 (N_2048,N_1989,N_1983);
or U2049 (N_2049,N_1997,N_1974);
and U2050 (N_2050,N_2035,N_2001);
or U2051 (N_2051,N_2008,N_2024);
or U2052 (N_2052,N_2046,N_2002);
nand U2053 (N_2053,N_2038,N_2020);
or U2054 (N_2054,N_2000,N_2018);
or U2055 (N_2055,N_2003,N_2015);
nor U2056 (N_2056,N_2027,N_2016);
nor U2057 (N_2057,N_2011,N_2012);
nor U2058 (N_2058,N_2021,N_2025);
nand U2059 (N_2059,N_2007,N_2048);
nand U2060 (N_2060,N_2045,N_2023);
and U2061 (N_2061,N_2017,N_2005);
or U2062 (N_2062,N_2049,N_2019);
and U2063 (N_2063,N_2040,N_2004);
and U2064 (N_2064,N_2031,N_2041);
nor U2065 (N_2065,N_2034,N_2044);
nand U2066 (N_2066,N_2036,N_2043);
or U2067 (N_2067,N_2014,N_2028);
or U2068 (N_2068,N_2029,N_2042);
nand U2069 (N_2069,N_2047,N_2006);
or U2070 (N_2070,N_2037,N_2026);
nand U2071 (N_2071,N_2022,N_2039);
or U2072 (N_2072,N_2032,N_2013);
nor U2073 (N_2073,N_2033,N_2030);
nor U2074 (N_2074,N_2010,N_2009);
and U2075 (N_2075,N_2046,N_2048);
and U2076 (N_2076,N_2049,N_2011);
and U2077 (N_2077,N_2019,N_2037);
and U2078 (N_2078,N_2025,N_2019);
nand U2079 (N_2079,N_2016,N_2000);
and U2080 (N_2080,N_2010,N_2019);
or U2081 (N_2081,N_2047,N_2041);
nand U2082 (N_2082,N_2028,N_2038);
or U2083 (N_2083,N_2017,N_2041);
nand U2084 (N_2084,N_2005,N_2024);
nand U2085 (N_2085,N_2042,N_2024);
or U2086 (N_2086,N_2024,N_2049);
or U2087 (N_2087,N_2011,N_2044);
nand U2088 (N_2088,N_2046,N_2024);
nand U2089 (N_2089,N_2041,N_2023);
and U2090 (N_2090,N_2012,N_2025);
or U2091 (N_2091,N_2040,N_2048);
and U2092 (N_2092,N_2012,N_2010);
nor U2093 (N_2093,N_2044,N_2013);
or U2094 (N_2094,N_2004,N_2038);
or U2095 (N_2095,N_2035,N_2011);
nor U2096 (N_2096,N_2046,N_2043);
nand U2097 (N_2097,N_2018,N_2044);
nand U2098 (N_2098,N_2047,N_2015);
nand U2099 (N_2099,N_2002,N_2031);
and U2100 (N_2100,N_2070,N_2054);
or U2101 (N_2101,N_2084,N_2058);
and U2102 (N_2102,N_2069,N_2074);
and U2103 (N_2103,N_2066,N_2089);
and U2104 (N_2104,N_2068,N_2056);
and U2105 (N_2105,N_2060,N_2078);
or U2106 (N_2106,N_2077,N_2085);
nand U2107 (N_2107,N_2064,N_2065);
nor U2108 (N_2108,N_2053,N_2055);
or U2109 (N_2109,N_2098,N_2087);
or U2110 (N_2110,N_2081,N_2073);
nand U2111 (N_2111,N_2057,N_2050);
or U2112 (N_2112,N_2061,N_2094);
nor U2113 (N_2113,N_2063,N_2080);
nand U2114 (N_2114,N_2082,N_2091);
nand U2115 (N_2115,N_2079,N_2099);
nand U2116 (N_2116,N_2076,N_2086);
and U2117 (N_2117,N_2075,N_2096);
and U2118 (N_2118,N_2052,N_2093);
nand U2119 (N_2119,N_2097,N_2059);
nor U2120 (N_2120,N_2090,N_2072);
nor U2121 (N_2121,N_2071,N_2051);
nand U2122 (N_2122,N_2062,N_2095);
or U2123 (N_2123,N_2088,N_2083);
nand U2124 (N_2124,N_2092,N_2067);
and U2125 (N_2125,N_2093,N_2084);
and U2126 (N_2126,N_2059,N_2052);
nor U2127 (N_2127,N_2068,N_2081);
and U2128 (N_2128,N_2084,N_2098);
or U2129 (N_2129,N_2065,N_2098);
or U2130 (N_2130,N_2075,N_2086);
nand U2131 (N_2131,N_2053,N_2076);
nor U2132 (N_2132,N_2074,N_2064);
nor U2133 (N_2133,N_2092,N_2059);
nand U2134 (N_2134,N_2096,N_2094);
and U2135 (N_2135,N_2095,N_2063);
nor U2136 (N_2136,N_2062,N_2089);
or U2137 (N_2137,N_2096,N_2061);
or U2138 (N_2138,N_2066,N_2080);
nor U2139 (N_2139,N_2091,N_2076);
nor U2140 (N_2140,N_2094,N_2054);
and U2141 (N_2141,N_2076,N_2069);
nand U2142 (N_2142,N_2065,N_2071);
nand U2143 (N_2143,N_2063,N_2064);
nand U2144 (N_2144,N_2091,N_2085);
or U2145 (N_2145,N_2051,N_2075);
nor U2146 (N_2146,N_2062,N_2096);
xor U2147 (N_2147,N_2077,N_2094);
or U2148 (N_2148,N_2064,N_2092);
nand U2149 (N_2149,N_2069,N_2081);
nor U2150 (N_2150,N_2143,N_2111);
and U2151 (N_2151,N_2123,N_2126);
and U2152 (N_2152,N_2105,N_2107);
or U2153 (N_2153,N_2148,N_2128);
and U2154 (N_2154,N_2139,N_2135);
nand U2155 (N_2155,N_2141,N_2118);
and U2156 (N_2156,N_2127,N_2129);
and U2157 (N_2157,N_2110,N_2136);
and U2158 (N_2158,N_2149,N_2144);
and U2159 (N_2159,N_2109,N_2103);
or U2160 (N_2160,N_2124,N_2112);
or U2161 (N_2161,N_2117,N_2115);
nand U2162 (N_2162,N_2147,N_2113);
and U2163 (N_2163,N_2108,N_2130);
nor U2164 (N_2164,N_2132,N_2104);
xnor U2165 (N_2165,N_2119,N_2102);
and U2166 (N_2166,N_2114,N_2131);
nor U2167 (N_2167,N_2140,N_2145);
and U2168 (N_2168,N_2120,N_2101);
or U2169 (N_2169,N_2134,N_2125);
nor U2170 (N_2170,N_2146,N_2138);
and U2171 (N_2171,N_2133,N_2137);
nand U2172 (N_2172,N_2122,N_2116);
or U2173 (N_2173,N_2106,N_2121);
nand U2174 (N_2174,N_2100,N_2142);
or U2175 (N_2175,N_2109,N_2122);
nand U2176 (N_2176,N_2139,N_2122);
nor U2177 (N_2177,N_2117,N_2149);
and U2178 (N_2178,N_2124,N_2148);
and U2179 (N_2179,N_2142,N_2117);
nor U2180 (N_2180,N_2130,N_2145);
or U2181 (N_2181,N_2149,N_2131);
or U2182 (N_2182,N_2105,N_2129);
or U2183 (N_2183,N_2125,N_2145);
and U2184 (N_2184,N_2110,N_2126);
nand U2185 (N_2185,N_2142,N_2140);
and U2186 (N_2186,N_2129,N_2101);
or U2187 (N_2187,N_2135,N_2131);
and U2188 (N_2188,N_2141,N_2117);
nor U2189 (N_2189,N_2102,N_2146);
and U2190 (N_2190,N_2103,N_2104);
and U2191 (N_2191,N_2123,N_2101);
nor U2192 (N_2192,N_2133,N_2111);
nand U2193 (N_2193,N_2138,N_2117);
nor U2194 (N_2194,N_2106,N_2138);
or U2195 (N_2195,N_2102,N_2148);
nand U2196 (N_2196,N_2124,N_2129);
nor U2197 (N_2197,N_2103,N_2108);
nand U2198 (N_2198,N_2131,N_2118);
nor U2199 (N_2199,N_2140,N_2147);
or U2200 (N_2200,N_2160,N_2158);
nand U2201 (N_2201,N_2168,N_2189);
nor U2202 (N_2202,N_2178,N_2151);
or U2203 (N_2203,N_2184,N_2153);
nand U2204 (N_2204,N_2166,N_2174);
or U2205 (N_2205,N_2181,N_2171);
nand U2206 (N_2206,N_2162,N_2164);
or U2207 (N_2207,N_2163,N_2196);
and U2208 (N_2208,N_2154,N_2155);
nor U2209 (N_2209,N_2175,N_2179);
or U2210 (N_2210,N_2180,N_2194);
nand U2211 (N_2211,N_2172,N_2177);
nand U2212 (N_2212,N_2191,N_2195);
nand U2213 (N_2213,N_2185,N_2165);
or U2214 (N_2214,N_2167,N_2159);
nor U2215 (N_2215,N_2192,N_2197);
xor U2216 (N_2216,N_2152,N_2193);
and U2217 (N_2217,N_2157,N_2170);
and U2218 (N_2218,N_2176,N_2161);
or U2219 (N_2219,N_2150,N_2156);
and U2220 (N_2220,N_2169,N_2190);
nor U2221 (N_2221,N_2199,N_2186);
and U2222 (N_2222,N_2183,N_2182);
nand U2223 (N_2223,N_2173,N_2187);
nor U2224 (N_2224,N_2188,N_2198);
nor U2225 (N_2225,N_2169,N_2162);
nand U2226 (N_2226,N_2195,N_2153);
nor U2227 (N_2227,N_2154,N_2160);
nor U2228 (N_2228,N_2190,N_2182);
xor U2229 (N_2229,N_2199,N_2160);
and U2230 (N_2230,N_2176,N_2196);
or U2231 (N_2231,N_2175,N_2153);
nand U2232 (N_2232,N_2162,N_2156);
nand U2233 (N_2233,N_2154,N_2167);
and U2234 (N_2234,N_2192,N_2158);
nor U2235 (N_2235,N_2185,N_2163);
nand U2236 (N_2236,N_2188,N_2173);
and U2237 (N_2237,N_2197,N_2154);
nor U2238 (N_2238,N_2199,N_2171);
or U2239 (N_2239,N_2181,N_2157);
or U2240 (N_2240,N_2193,N_2162);
nor U2241 (N_2241,N_2177,N_2153);
or U2242 (N_2242,N_2196,N_2191);
or U2243 (N_2243,N_2192,N_2173);
or U2244 (N_2244,N_2173,N_2170);
and U2245 (N_2245,N_2174,N_2157);
or U2246 (N_2246,N_2164,N_2185);
nand U2247 (N_2247,N_2175,N_2190);
and U2248 (N_2248,N_2163,N_2191);
and U2249 (N_2249,N_2186,N_2156);
or U2250 (N_2250,N_2215,N_2201);
nand U2251 (N_2251,N_2204,N_2203);
and U2252 (N_2252,N_2214,N_2235);
and U2253 (N_2253,N_2209,N_2249);
and U2254 (N_2254,N_2213,N_2211);
or U2255 (N_2255,N_2246,N_2200);
nand U2256 (N_2256,N_2230,N_2242);
or U2257 (N_2257,N_2218,N_2207);
nand U2258 (N_2258,N_2228,N_2244);
nor U2259 (N_2259,N_2241,N_2216);
nand U2260 (N_2260,N_2221,N_2234);
nor U2261 (N_2261,N_2202,N_2219);
and U2262 (N_2262,N_2243,N_2208);
or U2263 (N_2263,N_2238,N_2210);
nand U2264 (N_2264,N_2247,N_2245);
nand U2265 (N_2265,N_2236,N_2205);
nand U2266 (N_2266,N_2217,N_2248);
nand U2267 (N_2267,N_2232,N_2231);
and U2268 (N_2268,N_2237,N_2233);
nand U2269 (N_2269,N_2226,N_2240);
and U2270 (N_2270,N_2225,N_2212);
and U2271 (N_2271,N_2227,N_2220);
and U2272 (N_2272,N_2206,N_2223);
and U2273 (N_2273,N_2229,N_2239);
nor U2274 (N_2274,N_2224,N_2222);
nor U2275 (N_2275,N_2238,N_2230);
or U2276 (N_2276,N_2204,N_2237);
nor U2277 (N_2277,N_2230,N_2237);
and U2278 (N_2278,N_2214,N_2200);
nor U2279 (N_2279,N_2217,N_2239);
nand U2280 (N_2280,N_2206,N_2242);
nor U2281 (N_2281,N_2205,N_2227);
and U2282 (N_2282,N_2224,N_2225);
and U2283 (N_2283,N_2241,N_2245);
and U2284 (N_2284,N_2207,N_2200);
nand U2285 (N_2285,N_2217,N_2219);
nor U2286 (N_2286,N_2204,N_2219);
and U2287 (N_2287,N_2237,N_2205);
nor U2288 (N_2288,N_2243,N_2239);
nand U2289 (N_2289,N_2228,N_2243);
and U2290 (N_2290,N_2247,N_2217);
and U2291 (N_2291,N_2244,N_2219);
and U2292 (N_2292,N_2233,N_2216);
nand U2293 (N_2293,N_2230,N_2241);
or U2294 (N_2294,N_2209,N_2232);
or U2295 (N_2295,N_2233,N_2207);
nor U2296 (N_2296,N_2209,N_2202);
or U2297 (N_2297,N_2202,N_2236);
and U2298 (N_2298,N_2220,N_2248);
nor U2299 (N_2299,N_2218,N_2235);
or U2300 (N_2300,N_2254,N_2263);
and U2301 (N_2301,N_2285,N_2280);
nand U2302 (N_2302,N_2253,N_2292);
and U2303 (N_2303,N_2268,N_2261);
and U2304 (N_2304,N_2250,N_2297);
nand U2305 (N_2305,N_2274,N_2286);
and U2306 (N_2306,N_2288,N_2272);
and U2307 (N_2307,N_2270,N_2267);
or U2308 (N_2308,N_2279,N_2275);
and U2309 (N_2309,N_2282,N_2269);
and U2310 (N_2310,N_2283,N_2266);
and U2311 (N_2311,N_2278,N_2257);
or U2312 (N_2312,N_2294,N_2251);
nand U2313 (N_2313,N_2256,N_2273);
nand U2314 (N_2314,N_2295,N_2252);
nor U2315 (N_2315,N_2293,N_2258);
or U2316 (N_2316,N_2277,N_2299);
nand U2317 (N_2317,N_2259,N_2281);
nand U2318 (N_2318,N_2276,N_2289);
nor U2319 (N_2319,N_2284,N_2271);
nor U2320 (N_2320,N_2262,N_2264);
and U2321 (N_2321,N_2290,N_2298);
nor U2322 (N_2322,N_2255,N_2260);
nor U2323 (N_2323,N_2291,N_2287);
or U2324 (N_2324,N_2296,N_2265);
or U2325 (N_2325,N_2250,N_2296);
or U2326 (N_2326,N_2283,N_2269);
nor U2327 (N_2327,N_2278,N_2291);
and U2328 (N_2328,N_2276,N_2272);
and U2329 (N_2329,N_2263,N_2272);
nor U2330 (N_2330,N_2251,N_2286);
nor U2331 (N_2331,N_2280,N_2279);
nand U2332 (N_2332,N_2261,N_2293);
nor U2333 (N_2333,N_2259,N_2252);
or U2334 (N_2334,N_2265,N_2256);
or U2335 (N_2335,N_2258,N_2272);
nor U2336 (N_2336,N_2298,N_2297);
nor U2337 (N_2337,N_2285,N_2289);
nand U2338 (N_2338,N_2264,N_2263);
nand U2339 (N_2339,N_2297,N_2267);
or U2340 (N_2340,N_2290,N_2282);
and U2341 (N_2341,N_2289,N_2274);
nor U2342 (N_2342,N_2277,N_2266);
or U2343 (N_2343,N_2257,N_2256);
and U2344 (N_2344,N_2275,N_2251);
nor U2345 (N_2345,N_2283,N_2290);
nand U2346 (N_2346,N_2295,N_2281);
nand U2347 (N_2347,N_2259,N_2254);
or U2348 (N_2348,N_2264,N_2265);
nand U2349 (N_2349,N_2283,N_2254);
or U2350 (N_2350,N_2324,N_2313);
and U2351 (N_2351,N_2334,N_2333);
or U2352 (N_2352,N_2349,N_2309);
nand U2353 (N_2353,N_2319,N_2345);
nor U2354 (N_2354,N_2312,N_2320);
and U2355 (N_2355,N_2329,N_2306);
nor U2356 (N_2356,N_2339,N_2344);
or U2357 (N_2357,N_2315,N_2310);
nor U2358 (N_2358,N_2340,N_2300);
and U2359 (N_2359,N_2314,N_2326);
or U2360 (N_2360,N_2335,N_2307);
nand U2361 (N_2361,N_2323,N_2327);
nand U2362 (N_2362,N_2311,N_2348);
and U2363 (N_2363,N_2332,N_2301);
nand U2364 (N_2364,N_2343,N_2328);
nand U2365 (N_2365,N_2330,N_2325);
nor U2366 (N_2366,N_2318,N_2346);
nand U2367 (N_2367,N_2302,N_2336);
and U2368 (N_2368,N_2338,N_2305);
xor U2369 (N_2369,N_2337,N_2316);
or U2370 (N_2370,N_2308,N_2304);
nand U2371 (N_2371,N_2317,N_2347);
nor U2372 (N_2372,N_2342,N_2303);
nor U2373 (N_2373,N_2321,N_2331);
or U2374 (N_2374,N_2322,N_2341);
nand U2375 (N_2375,N_2300,N_2322);
nor U2376 (N_2376,N_2311,N_2304);
and U2377 (N_2377,N_2301,N_2327);
or U2378 (N_2378,N_2302,N_2340);
or U2379 (N_2379,N_2300,N_2326);
or U2380 (N_2380,N_2312,N_2306);
xnor U2381 (N_2381,N_2303,N_2341);
nand U2382 (N_2382,N_2344,N_2323);
or U2383 (N_2383,N_2320,N_2349);
and U2384 (N_2384,N_2302,N_2324);
nand U2385 (N_2385,N_2348,N_2342);
and U2386 (N_2386,N_2343,N_2345);
or U2387 (N_2387,N_2323,N_2318);
or U2388 (N_2388,N_2333,N_2345);
nand U2389 (N_2389,N_2301,N_2317);
nor U2390 (N_2390,N_2313,N_2311);
nor U2391 (N_2391,N_2317,N_2310);
or U2392 (N_2392,N_2346,N_2310);
nor U2393 (N_2393,N_2310,N_2333);
or U2394 (N_2394,N_2300,N_2303);
nor U2395 (N_2395,N_2304,N_2337);
nor U2396 (N_2396,N_2327,N_2310);
nor U2397 (N_2397,N_2347,N_2322);
or U2398 (N_2398,N_2308,N_2303);
or U2399 (N_2399,N_2306,N_2304);
and U2400 (N_2400,N_2397,N_2386);
nor U2401 (N_2401,N_2363,N_2383);
nand U2402 (N_2402,N_2393,N_2350);
and U2403 (N_2403,N_2370,N_2352);
and U2404 (N_2404,N_2360,N_2398);
nand U2405 (N_2405,N_2373,N_2381);
nor U2406 (N_2406,N_2368,N_2353);
nor U2407 (N_2407,N_2359,N_2389);
nor U2408 (N_2408,N_2376,N_2388);
or U2409 (N_2409,N_2387,N_2364);
and U2410 (N_2410,N_2378,N_2361);
nand U2411 (N_2411,N_2380,N_2369);
or U2412 (N_2412,N_2384,N_2356);
nand U2413 (N_2413,N_2372,N_2358);
and U2414 (N_2414,N_2351,N_2366);
nor U2415 (N_2415,N_2396,N_2395);
or U2416 (N_2416,N_2371,N_2390);
and U2417 (N_2417,N_2375,N_2377);
and U2418 (N_2418,N_2365,N_2382);
nand U2419 (N_2419,N_2367,N_2391);
nor U2420 (N_2420,N_2362,N_2392);
nand U2421 (N_2421,N_2394,N_2355);
or U2422 (N_2422,N_2374,N_2354);
and U2423 (N_2423,N_2399,N_2379);
nor U2424 (N_2424,N_2385,N_2357);
nor U2425 (N_2425,N_2393,N_2365);
and U2426 (N_2426,N_2382,N_2386);
nor U2427 (N_2427,N_2356,N_2376);
nand U2428 (N_2428,N_2360,N_2361);
nor U2429 (N_2429,N_2388,N_2391);
and U2430 (N_2430,N_2376,N_2397);
nor U2431 (N_2431,N_2395,N_2376);
or U2432 (N_2432,N_2396,N_2376);
nand U2433 (N_2433,N_2387,N_2351);
or U2434 (N_2434,N_2380,N_2364);
or U2435 (N_2435,N_2373,N_2356);
nand U2436 (N_2436,N_2382,N_2388);
or U2437 (N_2437,N_2351,N_2395);
nand U2438 (N_2438,N_2389,N_2367);
nand U2439 (N_2439,N_2381,N_2360);
or U2440 (N_2440,N_2351,N_2375);
nand U2441 (N_2441,N_2384,N_2362);
and U2442 (N_2442,N_2386,N_2391);
nor U2443 (N_2443,N_2364,N_2352);
nor U2444 (N_2444,N_2367,N_2396);
nand U2445 (N_2445,N_2362,N_2363);
xnor U2446 (N_2446,N_2385,N_2392);
or U2447 (N_2447,N_2358,N_2378);
or U2448 (N_2448,N_2375,N_2368);
or U2449 (N_2449,N_2393,N_2396);
nand U2450 (N_2450,N_2420,N_2418);
nand U2451 (N_2451,N_2433,N_2426);
and U2452 (N_2452,N_2417,N_2423);
nand U2453 (N_2453,N_2443,N_2405);
or U2454 (N_2454,N_2432,N_2442);
or U2455 (N_2455,N_2445,N_2416);
nor U2456 (N_2456,N_2434,N_2437);
or U2457 (N_2457,N_2422,N_2447);
and U2458 (N_2458,N_2401,N_2425);
and U2459 (N_2459,N_2419,N_2412);
nand U2460 (N_2460,N_2438,N_2427);
nor U2461 (N_2461,N_2435,N_2403);
or U2462 (N_2462,N_2440,N_2436);
or U2463 (N_2463,N_2406,N_2441);
nor U2464 (N_2464,N_2431,N_2448);
nand U2465 (N_2465,N_2404,N_2414);
nand U2466 (N_2466,N_2421,N_2410);
nand U2467 (N_2467,N_2402,N_2424);
and U2468 (N_2468,N_2444,N_2408);
or U2469 (N_2469,N_2439,N_2429);
nor U2470 (N_2470,N_2415,N_2409);
nor U2471 (N_2471,N_2449,N_2411);
or U2472 (N_2472,N_2413,N_2446);
and U2473 (N_2473,N_2407,N_2428);
nor U2474 (N_2474,N_2400,N_2430);
nor U2475 (N_2475,N_2422,N_2409);
nand U2476 (N_2476,N_2409,N_2421);
nand U2477 (N_2477,N_2411,N_2436);
nor U2478 (N_2478,N_2406,N_2436);
nor U2479 (N_2479,N_2404,N_2447);
nand U2480 (N_2480,N_2429,N_2412);
or U2481 (N_2481,N_2427,N_2437);
nor U2482 (N_2482,N_2446,N_2431);
nand U2483 (N_2483,N_2425,N_2402);
and U2484 (N_2484,N_2446,N_2443);
nand U2485 (N_2485,N_2448,N_2425);
and U2486 (N_2486,N_2417,N_2400);
nand U2487 (N_2487,N_2419,N_2432);
and U2488 (N_2488,N_2433,N_2412);
nand U2489 (N_2489,N_2446,N_2435);
or U2490 (N_2490,N_2441,N_2410);
nor U2491 (N_2491,N_2406,N_2448);
nand U2492 (N_2492,N_2437,N_2404);
or U2493 (N_2493,N_2438,N_2424);
nor U2494 (N_2494,N_2441,N_2408);
or U2495 (N_2495,N_2414,N_2446);
nor U2496 (N_2496,N_2400,N_2448);
nand U2497 (N_2497,N_2430,N_2433);
nand U2498 (N_2498,N_2431,N_2407);
nor U2499 (N_2499,N_2430,N_2428);
or U2500 (N_2500,N_2471,N_2461);
and U2501 (N_2501,N_2490,N_2474);
nor U2502 (N_2502,N_2462,N_2467);
nor U2503 (N_2503,N_2466,N_2451);
nand U2504 (N_2504,N_2483,N_2494);
nand U2505 (N_2505,N_2450,N_2489);
nand U2506 (N_2506,N_2458,N_2495);
nand U2507 (N_2507,N_2493,N_2455);
nand U2508 (N_2508,N_2478,N_2499);
nand U2509 (N_2509,N_2481,N_2469);
nand U2510 (N_2510,N_2473,N_2477);
nor U2511 (N_2511,N_2487,N_2480);
or U2512 (N_2512,N_2460,N_2465);
nor U2513 (N_2513,N_2453,N_2476);
nand U2514 (N_2514,N_2472,N_2464);
or U2515 (N_2515,N_2456,N_2457);
and U2516 (N_2516,N_2491,N_2486);
nor U2517 (N_2517,N_2482,N_2479);
nor U2518 (N_2518,N_2485,N_2475);
nor U2519 (N_2519,N_2498,N_2497);
or U2520 (N_2520,N_2459,N_2496);
and U2521 (N_2521,N_2492,N_2484);
nand U2522 (N_2522,N_2463,N_2454);
nor U2523 (N_2523,N_2488,N_2470);
nor U2524 (N_2524,N_2452,N_2468);
nor U2525 (N_2525,N_2464,N_2491);
or U2526 (N_2526,N_2462,N_2490);
nand U2527 (N_2527,N_2476,N_2488);
nor U2528 (N_2528,N_2468,N_2499);
nand U2529 (N_2529,N_2487,N_2469);
nand U2530 (N_2530,N_2459,N_2457);
nand U2531 (N_2531,N_2482,N_2475);
or U2532 (N_2532,N_2458,N_2480);
nand U2533 (N_2533,N_2480,N_2460);
or U2534 (N_2534,N_2454,N_2466);
or U2535 (N_2535,N_2466,N_2474);
nand U2536 (N_2536,N_2487,N_2475);
nand U2537 (N_2537,N_2487,N_2494);
nand U2538 (N_2538,N_2483,N_2457);
nand U2539 (N_2539,N_2469,N_2484);
and U2540 (N_2540,N_2465,N_2494);
or U2541 (N_2541,N_2487,N_2456);
and U2542 (N_2542,N_2461,N_2475);
nor U2543 (N_2543,N_2459,N_2474);
nor U2544 (N_2544,N_2484,N_2472);
nand U2545 (N_2545,N_2467,N_2481);
nor U2546 (N_2546,N_2471,N_2484);
and U2547 (N_2547,N_2479,N_2476);
and U2548 (N_2548,N_2470,N_2464);
nor U2549 (N_2549,N_2493,N_2462);
and U2550 (N_2550,N_2539,N_2534);
and U2551 (N_2551,N_2519,N_2528);
nor U2552 (N_2552,N_2517,N_2535);
or U2553 (N_2553,N_2537,N_2522);
and U2554 (N_2554,N_2548,N_2505);
nor U2555 (N_2555,N_2507,N_2541);
nor U2556 (N_2556,N_2510,N_2543);
or U2557 (N_2557,N_2503,N_2545);
or U2558 (N_2558,N_2504,N_2506);
nand U2559 (N_2559,N_2538,N_2516);
nor U2560 (N_2560,N_2531,N_2527);
or U2561 (N_2561,N_2509,N_2512);
or U2562 (N_2562,N_2530,N_2544);
nand U2563 (N_2563,N_2549,N_2540);
nor U2564 (N_2564,N_2523,N_2511);
and U2565 (N_2565,N_2546,N_2525);
or U2566 (N_2566,N_2514,N_2524);
nand U2567 (N_2567,N_2533,N_2515);
nand U2568 (N_2568,N_2500,N_2526);
and U2569 (N_2569,N_2547,N_2520);
nand U2570 (N_2570,N_2521,N_2513);
or U2571 (N_2571,N_2508,N_2529);
and U2572 (N_2572,N_2501,N_2542);
and U2573 (N_2573,N_2536,N_2502);
and U2574 (N_2574,N_2518,N_2532);
or U2575 (N_2575,N_2542,N_2520);
nand U2576 (N_2576,N_2548,N_2513);
or U2577 (N_2577,N_2501,N_2521);
nor U2578 (N_2578,N_2514,N_2547);
nand U2579 (N_2579,N_2532,N_2524);
nor U2580 (N_2580,N_2526,N_2540);
nor U2581 (N_2581,N_2509,N_2530);
or U2582 (N_2582,N_2509,N_2536);
xnor U2583 (N_2583,N_2519,N_2524);
or U2584 (N_2584,N_2527,N_2522);
or U2585 (N_2585,N_2538,N_2525);
or U2586 (N_2586,N_2505,N_2538);
nor U2587 (N_2587,N_2546,N_2517);
nor U2588 (N_2588,N_2507,N_2530);
and U2589 (N_2589,N_2500,N_2521);
and U2590 (N_2590,N_2501,N_2537);
nand U2591 (N_2591,N_2547,N_2516);
nor U2592 (N_2592,N_2501,N_2515);
and U2593 (N_2593,N_2510,N_2525);
nor U2594 (N_2594,N_2534,N_2544);
and U2595 (N_2595,N_2513,N_2530);
or U2596 (N_2596,N_2547,N_2507);
nor U2597 (N_2597,N_2522,N_2525);
or U2598 (N_2598,N_2511,N_2539);
nor U2599 (N_2599,N_2501,N_2544);
or U2600 (N_2600,N_2564,N_2587);
nand U2601 (N_2601,N_2562,N_2570);
nand U2602 (N_2602,N_2559,N_2550);
nor U2603 (N_2603,N_2573,N_2583);
and U2604 (N_2604,N_2597,N_2554);
nand U2605 (N_2605,N_2574,N_2569);
or U2606 (N_2606,N_2568,N_2582);
nand U2607 (N_2607,N_2593,N_2590);
or U2608 (N_2608,N_2552,N_2556);
nor U2609 (N_2609,N_2555,N_2579);
nor U2610 (N_2610,N_2561,N_2566);
nand U2611 (N_2611,N_2586,N_2591);
nand U2612 (N_2612,N_2594,N_2598);
or U2613 (N_2613,N_2577,N_2580);
nor U2614 (N_2614,N_2565,N_2567);
nand U2615 (N_2615,N_2575,N_2551);
and U2616 (N_2616,N_2588,N_2557);
and U2617 (N_2617,N_2560,N_2571);
nor U2618 (N_2618,N_2558,N_2581);
nor U2619 (N_2619,N_2596,N_2584);
and U2620 (N_2620,N_2595,N_2563);
and U2621 (N_2621,N_2585,N_2599);
nor U2622 (N_2622,N_2589,N_2592);
nor U2623 (N_2623,N_2578,N_2553);
nand U2624 (N_2624,N_2572,N_2576);
and U2625 (N_2625,N_2562,N_2573);
or U2626 (N_2626,N_2593,N_2586);
nor U2627 (N_2627,N_2597,N_2587);
nand U2628 (N_2628,N_2550,N_2579);
and U2629 (N_2629,N_2552,N_2573);
and U2630 (N_2630,N_2587,N_2585);
xor U2631 (N_2631,N_2578,N_2554);
nand U2632 (N_2632,N_2575,N_2558);
nand U2633 (N_2633,N_2550,N_2589);
nor U2634 (N_2634,N_2583,N_2564);
and U2635 (N_2635,N_2599,N_2551);
and U2636 (N_2636,N_2558,N_2572);
and U2637 (N_2637,N_2592,N_2586);
or U2638 (N_2638,N_2574,N_2592);
and U2639 (N_2639,N_2598,N_2558);
nor U2640 (N_2640,N_2559,N_2563);
nand U2641 (N_2641,N_2574,N_2557);
and U2642 (N_2642,N_2569,N_2597);
nand U2643 (N_2643,N_2573,N_2560);
and U2644 (N_2644,N_2597,N_2578);
or U2645 (N_2645,N_2553,N_2580);
and U2646 (N_2646,N_2552,N_2584);
or U2647 (N_2647,N_2579,N_2568);
and U2648 (N_2648,N_2566,N_2574);
nand U2649 (N_2649,N_2599,N_2584);
nor U2650 (N_2650,N_2638,N_2642);
nand U2651 (N_2651,N_2645,N_2635);
and U2652 (N_2652,N_2632,N_2605);
or U2653 (N_2653,N_2643,N_2630);
or U2654 (N_2654,N_2627,N_2615);
and U2655 (N_2655,N_2636,N_2607);
nand U2656 (N_2656,N_2614,N_2646);
and U2657 (N_2657,N_2612,N_2648);
or U2658 (N_2658,N_2621,N_2610);
or U2659 (N_2659,N_2641,N_2608);
or U2660 (N_2660,N_2629,N_2604);
xnor U2661 (N_2661,N_2640,N_2606);
xnor U2662 (N_2662,N_2622,N_2613);
nand U2663 (N_2663,N_2618,N_2619);
and U2664 (N_2664,N_2620,N_2602);
or U2665 (N_2665,N_2625,N_2616);
or U2666 (N_2666,N_2634,N_2628);
or U2667 (N_2667,N_2626,N_2639);
and U2668 (N_2668,N_2647,N_2600);
or U2669 (N_2669,N_2603,N_2617);
nor U2670 (N_2670,N_2611,N_2601);
nor U2671 (N_2671,N_2644,N_2623);
and U2672 (N_2672,N_2649,N_2624);
and U2673 (N_2673,N_2633,N_2631);
or U2674 (N_2674,N_2609,N_2637);
nand U2675 (N_2675,N_2634,N_2618);
and U2676 (N_2676,N_2609,N_2645);
or U2677 (N_2677,N_2649,N_2617);
nand U2678 (N_2678,N_2625,N_2605);
or U2679 (N_2679,N_2632,N_2612);
and U2680 (N_2680,N_2610,N_2619);
or U2681 (N_2681,N_2630,N_2607);
and U2682 (N_2682,N_2637,N_2622);
and U2683 (N_2683,N_2623,N_2632);
and U2684 (N_2684,N_2634,N_2644);
or U2685 (N_2685,N_2621,N_2602);
nor U2686 (N_2686,N_2640,N_2649);
or U2687 (N_2687,N_2642,N_2605);
nor U2688 (N_2688,N_2615,N_2604);
or U2689 (N_2689,N_2625,N_2610);
nand U2690 (N_2690,N_2604,N_2617);
or U2691 (N_2691,N_2645,N_2637);
nor U2692 (N_2692,N_2647,N_2611);
and U2693 (N_2693,N_2606,N_2634);
and U2694 (N_2694,N_2644,N_2609);
and U2695 (N_2695,N_2602,N_2648);
nand U2696 (N_2696,N_2622,N_2600);
nand U2697 (N_2697,N_2631,N_2605);
or U2698 (N_2698,N_2608,N_2632);
or U2699 (N_2699,N_2606,N_2622);
nor U2700 (N_2700,N_2683,N_2696);
nor U2701 (N_2701,N_2681,N_2654);
and U2702 (N_2702,N_2659,N_2650);
or U2703 (N_2703,N_2652,N_2674);
nor U2704 (N_2704,N_2651,N_2658);
nor U2705 (N_2705,N_2697,N_2662);
and U2706 (N_2706,N_2676,N_2689);
and U2707 (N_2707,N_2671,N_2686);
nand U2708 (N_2708,N_2694,N_2663);
nor U2709 (N_2709,N_2660,N_2679);
or U2710 (N_2710,N_2669,N_2672);
or U2711 (N_2711,N_2675,N_2664);
nor U2712 (N_2712,N_2668,N_2657);
nand U2713 (N_2713,N_2685,N_2666);
nand U2714 (N_2714,N_2680,N_2661);
nand U2715 (N_2715,N_2690,N_2691);
and U2716 (N_2716,N_2665,N_2673);
nor U2717 (N_2717,N_2695,N_2655);
or U2718 (N_2718,N_2699,N_2678);
nand U2719 (N_2719,N_2677,N_2692);
nor U2720 (N_2720,N_2698,N_2656);
or U2721 (N_2721,N_2687,N_2653);
and U2722 (N_2722,N_2684,N_2693);
nor U2723 (N_2723,N_2682,N_2667);
or U2724 (N_2724,N_2688,N_2670);
and U2725 (N_2725,N_2688,N_2657);
and U2726 (N_2726,N_2654,N_2661);
or U2727 (N_2727,N_2653,N_2650);
nand U2728 (N_2728,N_2696,N_2698);
nand U2729 (N_2729,N_2693,N_2678);
nand U2730 (N_2730,N_2650,N_2654);
nand U2731 (N_2731,N_2689,N_2696);
nor U2732 (N_2732,N_2666,N_2688);
nand U2733 (N_2733,N_2665,N_2666);
nand U2734 (N_2734,N_2683,N_2667);
nor U2735 (N_2735,N_2693,N_2652);
nand U2736 (N_2736,N_2680,N_2665);
nand U2737 (N_2737,N_2690,N_2656);
or U2738 (N_2738,N_2657,N_2694);
or U2739 (N_2739,N_2678,N_2658);
nor U2740 (N_2740,N_2666,N_2672);
or U2741 (N_2741,N_2662,N_2687);
nor U2742 (N_2742,N_2694,N_2688);
and U2743 (N_2743,N_2662,N_2651);
and U2744 (N_2744,N_2692,N_2662);
nor U2745 (N_2745,N_2667,N_2657);
nor U2746 (N_2746,N_2685,N_2658);
or U2747 (N_2747,N_2655,N_2664);
nand U2748 (N_2748,N_2696,N_2682);
or U2749 (N_2749,N_2665,N_2679);
nand U2750 (N_2750,N_2715,N_2737);
and U2751 (N_2751,N_2748,N_2703);
nor U2752 (N_2752,N_2702,N_2736);
nand U2753 (N_2753,N_2742,N_2723);
and U2754 (N_2754,N_2701,N_2714);
and U2755 (N_2755,N_2711,N_2722);
nand U2756 (N_2756,N_2731,N_2747);
nand U2757 (N_2757,N_2745,N_2708);
nor U2758 (N_2758,N_2712,N_2726);
or U2759 (N_2759,N_2704,N_2705);
nand U2760 (N_2760,N_2744,N_2743);
nand U2761 (N_2761,N_2734,N_2738);
nor U2762 (N_2762,N_2732,N_2709);
or U2763 (N_2763,N_2719,N_2724);
nand U2764 (N_2764,N_2720,N_2733);
nor U2765 (N_2765,N_2730,N_2739);
and U2766 (N_2766,N_2707,N_2718);
and U2767 (N_2767,N_2717,N_2740);
and U2768 (N_2768,N_2749,N_2716);
and U2769 (N_2769,N_2713,N_2729);
nor U2770 (N_2770,N_2710,N_2700);
nand U2771 (N_2771,N_2721,N_2746);
nor U2772 (N_2772,N_2741,N_2728);
nand U2773 (N_2773,N_2725,N_2735);
nor U2774 (N_2774,N_2727,N_2706);
nand U2775 (N_2775,N_2724,N_2707);
nand U2776 (N_2776,N_2746,N_2749);
and U2777 (N_2777,N_2718,N_2729);
nand U2778 (N_2778,N_2723,N_2743);
or U2779 (N_2779,N_2749,N_2726);
or U2780 (N_2780,N_2706,N_2709);
or U2781 (N_2781,N_2735,N_2729);
or U2782 (N_2782,N_2719,N_2720);
nand U2783 (N_2783,N_2707,N_2717);
nand U2784 (N_2784,N_2742,N_2713);
and U2785 (N_2785,N_2714,N_2741);
or U2786 (N_2786,N_2723,N_2722);
and U2787 (N_2787,N_2729,N_2746);
or U2788 (N_2788,N_2710,N_2740);
nand U2789 (N_2789,N_2727,N_2709);
nor U2790 (N_2790,N_2719,N_2732);
nor U2791 (N_2791,N_2711,N_2730);
and U2792 (N_2792,N_2724,N_2728);
and U2793 (N_2793,N_2719,N_2703);
and U2794 (N_2794,N_2745,N_2730);
nand U2795 (N_2795,N_2715,N_2703);
or U2796 (N_2796,N_2704,N_2741);
and U2797 (N_2797,N_2732,N_2705);
xor U2798 (N_2798,N_2748,N_2733);
or U2799 (N_2799,N_2745,N_2713);
nor U2800 (N_2800,N_2765,N_2775);
or U2801 (N_2801,N_2753,N_2778);
nor U2802 (N_2802,N_2793,N_2750);
nor U2803 (N_2803,N_2762,N_2758);
or U2804 (N_2804,N_2751,N_2792);
nor U2805 (N_2805,N_2754,N_2788);
nor U2806 (N_2806,N_2773,N_2755);
and U2807 (N_2807,N_2784,N_2756);
nand U2808 (N_2808,N_2790,N_2795);
nand U2809 (N_2809,N_2767,N_2771);
nand U2810 (N_2810,N_2772,N_2799);
nor U2811 (N_2811,N_2763,N_2764);
and U2812 (N_2812,N_2796,N_2768);
nand U2813 (N_2813,N_2789,N_2798);
xnor U2814 (N_2814,N_2761,N_2794);
or U2815 (N_2815,N_2786,N_2791);
or U2816 (N_2816,N_2785,N_2759);
and U2817 (N_2817,N_2760,N_2769);
or U2818 (N_2818,N_2797,N_2757);
nor U2819 (N_2819,N_2783,N_2770);
nand U2820 (N_2820,N_2787,N_2779);
or U2821 (N_2821,N_2766,N_2782);
nand U2822 (N_2822,N_2776,N_2752);
and U2823 (N_2823,N_2781,N_2780);
nand U2824 (N_2824,N_2777,N_2774);
nand U2825 (N_2825,N_2773,N_2761);
or U2826 (N_2826,N_2775,N_2769);
nor U2827 (N_2827,N_2759,N_2789);
nor U2828 (N_2828,N_2798,N_2786);
nand U2829 (N_2829,N_2795,N_2784);
nor U2830 (N_2830,N_2793,N_2783);
or U2831 (N_2831,N_2786,N_2764);
nor U2832 (N_2832,N_2788,N_2786);
xor U2833 (N_2833,N_2773,N_2794);
nor U2834 (N_2834,N_2769,N_2761);
nor U2835 (N_2835,N_2768,N_2775);
and U2836 (N_2836,N_2785,N_2763);
and U2837 (N_2837,N_2758,N_2761);
nand U2838 (N_2838,N_2783,N_2751);
and U2839 (N_2839,N_2770,N_2754);
or U2840 (N_2840,N_2790,N_2783);
or U2841 (N_2841,N_2771,N_2797);
nand U2842 (N_2842,N_2769,N_2767);
or U2843 (N_2843,N_2782,N_2756);
nand U2844 (N_2844,N_2793,N_2760);
and U2845 (N_2845,N_2752,N_2754);
or U2846 (N_2846,N_2765,N_2797);
and U2847 (N_2847,N_2780,N_2778);
nand U2848 (N_2848,N_2777,N_2780);
and U2849 (N_2849,N_2761,N_2795);
or U2850 (N_2850,N_2820,N_2809);
nand U2851 (N_2851,N_2827,N_2837);
nand U2852 (N_2852,N_2818,N_2832);
or U2853 (N_2853,N_2834,N_2831);
or U2854 (N_2854,N_2848,N_2825);
or U2855 (N_2855,N_2802,N_2846);
or U2856 (N_2856,N_2836,N_2824);
nor U2857 (N_2857,N_2828,N_2823);
and U2858 (N_2858,N_2807,N_2819);
nor U2859 (N_2859,N_2810,N_2840);
or U2860 (N_2860,N_2813,N_2839);
nand U2861 (N_2861,N_2815,N_2849);
and U2862 (N_2862,N_2814,N_2806);
or U2863 (N_2863,N_2841,N_2811);
or U2864 (N_2864,N_2808,N_2842);
nand U2865 (N_2865,N_2826,N_2821);
nor U2866 (N_2866,N_2812,N_2845);
nor U2867 (N_2867,N_2803,N_2844);
nand U2868 (N_2868,N_2833,N_2843);
or U2869 (N_2869,N_2804,N_2816);
nand U2870 (N_2870,N_2835,N_2801);
nor U2871 (N_2871,N_2830,N_2817);
or U2872 (N_2872,N_2847,N_2800);
nor U2873 (N_2873,N_2822,N_2805);
nor U2874 (N_2874,N_2838,N_2829);
nand U2875 (N_2875,N_2835,N_2839);
nor U2876 (N_2876,N_2841,N_2822);
and U2877 (N_2877,N_2819,N_2847);
or U2878 (N_2878,N_2846,N_2845);
or U2879 (N_2879,N_2807,N_2802);
nor U2880 (N_2880,N_2813,N_2818);
or U2881 (N_2881,N_2807,N_2836);
nor U2882 (N_2882,N_2824,N_2804);
or U2883 (N_2883,N_2843,N_2845);
and U2884 (N_2884,N_2843,N_2830);
and U2885 (N_2885,N_2828,N_2824);
nor U2886 (N_2886,N_2804,N_2823);
nor U2887 (N_2887,N_2808,N_2800);
or U2888 (N_2888,N_2803,N_2824);
and U2889 (N_2889,N_2841,N_2824);
nor U2890 (N_2890,N_2822,N_2825);
and U2891 (N_2891,N_2821,N_2839);
and U2892 (N_2892,N_2834,N_2835);
nor U2893 (N_2893,N_2834,N_2840);
or U2894 (N_2894,N_2839,N_2843);
nor U2895 (N_2895,N_2800,N_2813);
nand U2896 (N_2896,N_2830,N_2842);
and U2897 (N_2897,N_2830,N_2811);
nand U2898 (N_2898,N_2832,N_2800);
nand U2899 (N_2899,N_2842,N_2845);
nor U2900 (N_2900,N_2855,N_2888);
or U2901 (N_2901,N_2885,N_2881);
and U2902 (N_2902,N_2869,N_2879);
nand U2903 (N_2903,N_2884,N_2857);
nor U2904 (N_2904,N_2866,N_2858);
nand U2905 (N_2905,N_2882,N_2865);
and U2906 (N_2906,N_2868,N_2867);
nor U2907 (N_2907,N_2859,N_2862);
nand U2908 (N_2908,N_2891,N_2861);
nor U2909 (N_2909,N_2897,N_2886);
nand U2910 (N_2910,N_2893,N_2876);
and U2911 (N_2911,N_2895,N_2898);
nor U2912 (N_2912,N_2883,N_2872);
and U2913 (N_2913,N_2871,N_2877);
and U2914 (N_2914,N_2889,N_2887);
and U2915 (N_2915,N_2875,N_2890);
nand U2916 (N_2916,N_2850,N_2852);
nand U2917 (N_2917,N_2894,N_2896);
and U2918 (N_2918,N_2892,N_2851);
and U2919 (N_2919,N_2853,N_2863);
or U2920 (N_2920,N_2874,N_2880);
nor U2921 (N_2921,N_2860,N_2864);
nand U2922 (N_2922,N_2899,N_2854);
nor U2923 (N_2923,N_2856,N_2878);
or U2924 (N_2924,N_2873,N_2870);
and U2925 (N_2925,N_2896,N_2886);
and U2926 (N_2926,N_2875,N_2894);
or U2927 (N_2927,N_2881,N_2899);
nor U2928 (N_2928,N_2891,N_2870);
or U2929 (N_2929,N_2852,N_2883);
and U2930 (N_2930,N_2891,N_2857);
nor U2931 (N_2931,N_2894,N_2857);
nor U2932 (N_2932,N_2860,N_2896);
xor U2933 (N_2933,N_2878,N_2864);
and U2934 (N_2934,N_2857,N_2887);
nand U2935 (N_2935,N_2870,N_2868);
nand U2936 (N_2936,N_2898,N_2853);
nor U2937 (N_2937,N_2861,N_2865);
and U2938 (N_2938,N_2895,N_2873);
or U2939 (N_2939,N_2869,N_2851);
and U2940 (N_2940,N_2862,N_2884);
nand U2941 (N_2941,N_2882,N_2879);
nand U2942 (N_2942,N_2866,N_2886);
and U2943 (N_2943,N_2883,N_2891);
nand U2944 (N_2944,N_2885,N_2863);
or U2945 (N_2945,N_2861,N_2850);
and U2946 (N_2946,N_2882,N_2866);
nor U2947 (N_2947,N_2855,N_2898);
or U2948 (N_2948,N_2889,N_2895);
and U2949 (N_2949,N_2868,N_2858);
and U2950 (N_2950,N_2926,N_2929);
nand U2951 (N_2951,N_2945,N_2909);
or U2952 (N_2952,N_2937,N_2932);
nand U2953 (N_2953,N_2928,N_2936);
nand U2954 (N_2954,N_2908,N_2944);
nand U2955 (N_2955,N_2911,N_2931);
and U2956 (N_2956,N_2921,N_2941);
and U2957 (N_2957,N_2902,N_2940);
and U2958 (N_2958,N_2930,N_2903);
nand U2959 (N_2959,N_2916,N_2927);
nand U2960 (N_2960,N_2923,N_2946);
and U2961 (N_2961,N_2913,N_2947);
nor U2962 (N_2962,N_2900,N_2942);
nor U2963 (N_2963,N_2910,N_2914);
and U2964 (N_2964,N_2948,N_2906);
xor U2965 (N_2965,N_2934,N_2915);
and U2966 (N_2966,N_2920,N_2904);
nor U2967 (N_2967,N_2939,N_2907);
or U2968 (N_2968,N_2943,N_2917);
nor U2969 (N_2969,N_2919,N_2938);
nor U2970 (N_2970,N_2935,N_2905);
nand U2971 (N_2971,N_2918,N_2933);
nand U2972 (N_2972,N_2949,N_2922);
nand U2973 (N_2973,N_2901,N_2912);
and U2974 (N_2974,N_2924,N_2925);
or U2975 (N_2975,N_2932,N_2947);
or U2976 (N_2976,N_2904,N_2935);
and U2977 (N_2977,N_2927,N_2924);
and U2978 (N_2978,N_2923,N_2909);
nor U2979 (N_2979,N_2907,N_2935);
nor U2980 (N_2980,N_2946,N_2926);
and U2981 (N_2981,N_2938,N_2903);
nand U2982 (N_2982,N_2935,N_2942);
and U2983 (N_2983,N_2923,N_2913);
and U2984 (N_2984,N_2933,N_2925);
and U2985 (N_2985,N_2949,N_2909);
or U2986 (N_2986,N_2927,N_2931);
or U2987 (N_2987,N_2936,N_2945);
or U2988 (N_2988,N_2916,N_2920);
nand U2989 (N_2989,N_2942,N_2933);
nand U2990 (N_2990,N_2904,N_2909);
nor U2991 (N_2991,N_2920,N_2927);
and U2992 (N_2992,N_2910,N_2946);
or U2993 (N_2993,N_2908,N_2928);
nor U2994 (N_2994,N_2915,N_2939);
or U2995 (N_2995,N_2948,N_2946);
or U2996 (N_2996,N_2905,N_2921);
nand U2997 (N_2997,N_2920,N_2900);
or U2998 (N_2998,N_2910,N_2902);
or U2999 (N_2999,N_2938,N_2937);
nor UO_0 (O_0,N_2997,N_2969);
xnor UO_1 (O_1,N_2967,N_2961);
nand UO_2 (O_2,N_2962,N_2979);
nand UO_3 (O_3,N_2974,N_2985);
and UO_4 (O_4,N_2986,N_2995);
or UO_5 (O_5,N_2993,N_2972);
nand UO_6 (O_6,N_2980,N_2977);
or UO_7 (O_7,N_2953,N_2968);
nand UO_8 (O_8,N_2958,N_2978);
or UO_9 (O_9,N_2982,N_2951);
nand UO_10 (O_10,N_2963,N_2989);
or UO_11 (O_11,N_2991,N_2966);
nand UO_12 (O_12,N_2954,N_2970);
or UO_13 (O_13,N_2976,N_2956);
and UO_14 (O_14,N_2999,N_2950);
and UO_15 (O_15,N_2983,N_2987);
or UO_16 (O_16,N_2960,N_2988);
nor UO_17 (O_17,N_2996,N_2984);
nand UO_18 (O_18,N_2964,N_2998);
or UO_19 (O_19,N_2955,N_2965);
and UO_20 (O_20,N_2952,N_2975);
or UO_21 (O_21,N_2990,N_2992);
nor UO_22 (O_22,N_2957,N_2973);
nor UO_23 (O_23,N_2994,N_2981);
or UO_24 (O_24,N_2959,N_2971);
nand UO_25 (O_25,N_2990,N_2964);
nor UO_26 (O_26,N_2991,N_2970);
or UO_27 (O_27,N_2978,N_2973);
nor UO_28 (O_28,N_2970,N_2986);
and UO_29 (O_29,N_2968,N_2996);
nand UO_30 (O_30,N_2954,N_2955);
nor UO_31 (O_31,N_2983,N_2971);
nor UO_32 (O_32,N_2978,N_2959);
nor UO_33 (O_33,N_2965,N_2953);
xor UO_34 (O_34,N_2959,N_2955);
or UO_35 (O_35,N_2966,N_2951);
and UO_36 (O_36,N_2961,N_2966);
nor UO_37 (O_37,N_2987,N_2961);
and UO_38 (O_38,N_2986,N_2983);
and UO_39 (O_39,N_2965,N_2990);
and UO_40 (O_40,N_2998,N_2990);
nor UO_41 (O_41,N_2990,N_2997);
and UO_42 (O_42,N_2979,N_2980);
nand UO_43 (O_43,N_2976,N_2951);
and UO_44 (O_44,N_2968,N_2950);
nand UO_45 (O_45,N_2954,N_2973);
and UO_46 (O_46,N_2980,N_2968);
and UO_47 (O_47,N_2988,N_2954);
or UO_48 (O_48,N_2957,N_2971);
nor UO_49 (O_49,N_2987,N_2970);
nor UO_50 (O_50,N_2989,N_2965);
nand UO_51 (O_51,N_2991,N_2956);
and UO_52 (O_52,N_2992,N_2989);
nor UO_53 (O_53,N_2966,N_2978);
and UO_54 (O_54,N_2992,N_2985);
nand UO_55 (O_55,N_2999,N_2986);
nand UO_56 (O_56,N_2966,N_2971);
nor UO_57 (O_57,N_2990,N_2959);
and UO_58 (O_58,N_2996,N_2951);
and UO_59 (O_59,N_2959,N_2965);
and UO_60 (O_60,N_2955,N_2996);
nand UO_61 (O_61,N_2954,N_2958);
nor UO_62 (O_62,N_2977,N_2981);
or UO_63 (O_63,N_2998,N_2979);
or UO_64 (O_64,N_2989,N_2952);
nor UO_65 (O_65,N_2955,N_2971);
and UO_66 (O_66,N_2992,N_2961);
and UO_67 (O_67,N_2979,N_2973);
nor UO_68 (O_68,N_2963,N_2999);
nand UO_69 (O_69,N_2998,N_2950);
and UO_70 (O_70,N_2976,N_2971);
and UO_71 (O_71,N_2966,N_2992);
or UO_72 (O_72,N_2961,N_2984);
or UO_73 (O_73,N_2967,N_2960);
or UO_74 (O_74,N_2991,N_2951);
and UO_75 (O_75,N_2995,N_2979);
or UO_76 (O_76,N_2951,N_2998);
nor UO_77 (O_77,N_2982,N_2969);
nand UO_78 (O_78,N_2979,N_2989);
and UO_79 (O_79,N_2952,N_2999);
nor UO_80 (O_80,N_2970,N_2985);
or UO_81 (O_81,N_2980,N_2997);
and UO_82 (O_82,N_2988,N_2967);
or UO_83 (O_83,N_2994,N_2972);
and UO_84 (O_84,N_2952,N_2974);
nand UO_85 (O_85,N_2979,N_2984);
nor UO_86 (O_86,N_2987,N_2960);
nor UO_87 (O_87,N_2975,N_2980);
nand UO_88 (O_88,N_2975,N_2961);
nor UO_89 (O_89,N_2975,N_2967);
or UO_90 (O_90,N_2976,N_2968);
nand UO_91 (O_91,N_2972,N_2970);
and UO_92 (O_92,N_2955,N_2995);
and UO_93 (O_93,N_2976,N_2959);
nand UO_94 (O_94,N_2995,N_2982);
xnor UO_95 (O_95,N_2950,N_2978);
or UO_96 (O_96,N_2977,N_2992);
nand UO_97 (O_97,N_2990,N_2972);
nand UO_98 (O_98,N_2958,N_2956);
nor UO_99 (O_99,N_2968,N_2985);
or UO_100 (O_100,N_2955,N_2997);
and UO_101 (O_101,N_2977,N_2965);
or UO_102 (O_102,N_2962,N_2977);
nand UO_103 (O_103,N_2984,N_2976);
nor UO_104 (O_104,N_2988,N_2989);
and UO_105 (O_105,N_2975,N_2958);
or UO_106 (O_106,N_2982,N_2998);
and UO_107 (O_107,N_2980,N_2963);
or UO_108 (O_108,N_2981,N_2992);
nand UO_109 (O_109,N_2999,N_2962);
or UO_110 (O_110,N_2972,N_2995);
nor UO_111 (O_111,N_2967,N_2957);
nand UO_112 (O_112,N_2980,N_2950);
nand UO_113 (O_113,N_2953,N_2962);
and UO_114 (O_114,N_2962,N_2987);
or UO_115 (O_115,N_2973,N_2960);
or UO_116 (O_116,N_2975,N_2983);
and UO_117 (O_117,N_2990,N_2994);
or UO_118 (O_118,N_2994,N_2966);
and UO_119 (O_119,N_2997,N_2992);
xnor UO_120 (O_120,N_2976,N_2966);
and UO_121 (O_121,N_2983,N_2988);
nor UO_122 (O_122,N_2959,N_2994);
or UO_123 (O_123,N_2965,N_2993);
nand UO_124 (O_124,N_2952,N_2954);
nor UO_125 (O_125,N_2952,N_2984);
and UO_126 (O_126,N_2996,N_2983);
or UO_127 (O_127,N_2998,N_2974);
nand UO_128 (O_128,N_2983,N_2990);
and UO_129 (O_129,N_2994,N_2969);
nand UO_130 (O_130,N_2950,N_2985);
nand UO_131 (O_131,N_2963,N_2990);
nand UO_132 (O_132,N_2985,N_2956);
nand UO_133 (O_133,N_2974,N_2957);
nor UO_134 (O_134,N_2968,N_2973);
and UO_135 (O_135,N_2979,N_2994);
nand UO_136 (O_136,N_2956,N_2996);
or UO_137 (O_137,N_2973,N_2961);
or UO_138 (O_138,N_2987,N_2984);
and UO_139 (O_139,N_2991,N_2976);
nor UO_140 (O_140,N_2954,N_2980);
nand UO_141 (O_141,N_2996,N_2970);
and UO_142 (O_142,N_2999,N_2984);
nor UO_143 (O_143,N_2968,N_2952);
or UO_144 (O_144,N_2996,N_2950);
and UO_145 (O_145,N_2950,N_2964);
nand UO_146 (O_146,N_2963,N_2975);
or UO_147 (O_147,N_2966,N_2962);
nand UO_148 (O_148,N_2996,N_2963);
nand UO_149 (O_149,N_2986,N_2990);
or UO_150 (O_150,N_2990,N_2987);
nand UO_151 (O_151,N_2970,N_2968);
nor UO_152 (O_152,N_2983,N_2960);
nor UO_153 (O_153,N_2982,N_2972);
nor UO_154 (O_154,N_2964,N_2962);
nand UO_155 (O_155,N_2995,N_2967);
nand UO_156 (O_156,N_2962,N_2994);
nor UO_157 (O_157,N_2975,N_2973);
or UO_158 (O_158,N_2973,N_2989);
nand UO_159 (O_159,N_2971,N_2996);
nor UO_160 (O_160,N_2987,N_2989);
and UO_161 (O_161,N_2956,N_2980);
nor UO_162 (O_162,N_2991,N_2977);
nor UO_163 (O_163,N_2981,N_2980);
and UO_164 (O_164,N_2996,N_2992);
or UO_165 (O_165,N_2950,N_2981);
nand UO_166 (O_166,N_2963,N_2974);
or UO_167 (O_167,N_2997,N_2954);
nor UO_168 (O_168,N_2959,N_2960);
nand UO_169 (O_169,N_2958,N_2955);
or UO_170 (O_170,N_2965,N_2981);
and UO_171 (O_171,N_2984,N_2988);
xor UO_172 (O_172,N_2971,N_2973);
xnor UO_173 (O_173,N_2952,N_2998);
and UO_174 (O_174,N_2962,N_2991);
and UO_175 (O_175,N_2957,N_2953);
or UO_176 (O_176,N_2954,N_2971);
and UO_177 (O_177,N_2951,N_2993);
and UO_178 (O_178,N_2997,N_2999);
and UO_179 (O_179,N_2999,N_2972);
nand UO_180 (O_180,N_2978,N_2964);
and UO_181 (O_181,N_2993,N_2989);
or UO_182 (O_182,N_2962,N_2997);
nor UO_183 (O_183,N_2973,N_2969);
xnor UO_184 (O_184,N_2976,N_2952);
or UO_185 (O_185,N_2959,N_2984);
and UO_186 (O_186,N_2982,N_2996);
or UO_187 (O_187,N_2995,N_2960);
nand UO_188 (O_188,N_2978,N_2990);
and UO_189 (O_189,N_2958,N_2957);
nand UO_190 (O_190,N_2972,N_2992);
nor UO_191 (O_191,N_2975,N_2981);
nand UO_192 (O_192,N_2952,N_2996);
nand UO_193 (O_193,N_2960,N_2972);
or UO_194 (O_194,N_2987,N_2951);
nor UO_195 (O_195,N_2992,N_2952);
nand UO_196 (O_196,N_2981,N_2988);
and UO_197 (O_197,N_2971,N_2978);
and UO_198 (O_198,N_2999,N_2983);
nand UO_199 (O_199,N_2986,N_2953);
or UO_200 (O_200,N_2962,N_2957);
and UO_201 (O_201,N_2952,N_2967);
nor UO_202 (O_202,N_2973,N_2955);
nand UO_203 (O_203,N_2968,N_2951);
nand UO_204 (O_204,N_2962,N_2973);
nor UO_205 (O_205,N_2950,N_2972);
nor UO_206 (O_206,N_2991,N_2969);
and UO_207 (O_207,N_2969,N_2958);
or UO_208 (O_208,N_2960,N_2950);
or UO_209 (O_209,N_2965,N_2969);
or UO_210 (O_210,N_2985,N_2963);
and UO_211 (O_211,N_2993,N_2966);
and UO_212 (O_212,N_2994,N_2982);
and UO_213 (O_213,N_2972,N_2962);
nand UO_214 (O_214,N_2990,N_2962);
nand UO_215 (O_215,N_2993,N_2997);
or UO_216 (O_216,N_2989,N_2953);
and UO_217 (O_217,N_2958,N_2967);
and UO_218 (O_218,N_2985,N_2966);
nor UO_219 (O_219,N_2980,N_2986);
and UO_220 (O_220,N_2978,N_2998);
and UO_221 (O_221,N_2986,N_2984);
nand UO_222 (O_222,N_2951,N_2983);
or UO_223 (O_223,N_2996,N_2981);
and UO_224 (O_224,N_2963,N_2987);
and UO_225 (O_225,N_2971,N_2970);
or UO_226 (O_226,N_2990,N_2954);
and UO_227 (O_227,N_2992,N_2987);
nand UO_228 (O_228,N_2981,N_2987);
nand UO_229 (O_229,N_2978,N_2962);
nor UO_230 (O_230,N_2954,N_2972);
nor UO_231 (O_231,N_2962,N_2970);
and UO_232 (O_232,N_2954,N_2950);
nand UO_233 (O_233,N_2974,N_2996);
nand UO_234 (O_234,N_2988,N_2968);
or UO_235 (O_235,N_2990,N_2974);
and UO_236 (O_236,N_2991,N_2953);
nand UO_237 (O_237,N_2974,N_2989);
nand UO_238 (O_238,N_2984,N_2962);
and UO_239 (O_239,N_2967,N_2971);
and UO_240 (O_240,N_2983,N_2989);
nor UO_241 (O_241,N_2968,N_2960);
or UO_242 (O_242,N_2987,N_2977);
nor UO_243 (O_243,N_2983,N_2963);
nor UO_244 (O_244,N_2975,N_2993);
nand UO_245 (O_245,N_2960,N_2991);
nand UO_246 (O_246,N_2971,N_2960);
and UO_247 (O_247,N_2993,N_2953);
nand UO_248 (O_248,N_2960,N_2957);
nor UO_249 (O_249,N_2963,N_2981);
nand UO_250 (O_250,N_2963,N_2977);
nand UO_251 (O_251,N_2961,N_2983);
and UO_252 (O_252,N_2970,N_2959);
nand UO_253 (O_253,N_2970,N_2997);
or UO_254 (O_254,N_2984,N_2950);
and UO_255 (O_255,N_2963,N_2961);
nand UO_256 (O_256,N_2969,N_2962);
nor UO_257 (O_257,N_2973,N_2997);
and UO_258 (O_258,N_2992,N_2998);
or UO_259 (O_259,N_2993,N_2963);
nand UO_260 (O_260,N_2975,N_2953);
nand UO_261 (O_261,N_2955,N_2953);
and UO_262 (O_262,N_2952,N_2980);
nor UO_263 (O_263,N_2976,N_2978);
or UO_264 (O_264,N_2986,N_2958);
or UO_265 (O_265,N_2967,N_2981);
or UO_266 (O_266,N_2975,N_2964);
nand UO_267 (O_267,N_2998,N_2981);
and UO_268 (O_268,N_2988,N_2966);
nand UO_269 (O_269,N_2995,N_2981);
and UO_270 (O_270,N_2967,N_2992);
nor UO_271 (O_271,N_2987,N_2964);
and UO_272 (O_272,N_2950,N_2955);
or UO_273 (O_273,N_2999,N_2995);
nand UO_274 (O_274,N_2970,N_2993);
nor UO_275 (O_275,N_2994,N_2967);
nor UO_276 (O_276,N_2971,N_2952);
nor UO_277 (O_277,N_2981,N_2972);
nand UO_278 (O_278,N_2974,N_2987);
nand UO_279 (O_279,N_2951,N_2995);
nor UO_280 (O_280,N_2953,N_2960);
and UO_281 (O_281,N_2976,N_2975);
or UO_282 (O_282,N_2984,N_2990);
nor UO_283 (O_283,N_2960,N_2992);
nand UO_284 (O_284,N_2950,N_2991);
nor UO_285 (O_285,N_2978,N_2968);
and UO_286 (O_286,N_2968,N_2956);
nand UO_287 (O_287,N_2984,N_2991);
nand UO_288 (O_288,N_2985,N_2972);
nand UO_289 (O_289,N_2970,N_2978);
nand UO_290 (O_290,N_2999,N_2970);
xnor UO_291 (O_291,N_2950,N_2990);
and UO_292 (O_292,N_2967,N_2982);
and UO_293 (O_293,N_2988,N_2990);
nor UO_294 (O_294,N_2976,N_2998);
or UO_295 (O_295,N_2972,N_2968);
nand UO_296 (O_296,N_2964,N_2953);
nand UO_297 (O_297,N_2981,N_2956);
nand UO_298 (O_298,N_2962,N_2958);
or UO_299 (O_299,N_2990,N_2960);
nor UO_300 (O_300,N_2978,N_2999);
or UO_301 (O_301,N_2969,N_2956);
nand UO_302 (O_302,N_2955,N_2977);
nand UO_303 (O_303,N_2952,N_2997);
or UO_304 (O_304,N_2969,N_2984);
nand UO_305 (O_305,N_2959,N_2988);
or UO_306 (O_306,N_2967,N_2999);
or UO_307 (O_307,N_2992,N_2976);
nand UO_308 (O_308,N_2998,N_2968);
nand UO_309 (O_309,N_2982,N_2987);
nand UO_310 (O_310,N_2979,N_2988);
or UO_311 (O_311,N_2955,N_2988);
and UO_312 (O_312,N_2953,N_2958);
nand UO_313 (O_313,N_2965,N_2956);
and UO_314 (O_314,N_2969,N_2998);
and UO_315 (O_315,N_2974,N_2992);
nand UO_316 (O_316,N_2994,N_2971);
and UO_317 (O_317,N_2967,N_2979);
or UO_318 (O_318,N_2958,N_2992);
nand UO_319 (O_319,N_2958,N_2996);
and UO_320 (O_320,N_2952,N_2962);
nand UO_321 (O_321,N_2991,N_2994);
and UO_322 (O_322,N_2975,N_2986);
nand UO_323 (O_323,N_2958,N_2990);
and UO_324 (O_324,N_2954,N_2957);
nand UO_325 (O_325,N_2994,N_2985);
or UO_326 (O_326,N_2994,N_2997);
nor UO_327 (O_327,N_2987,N_2972);
or UO_328 (O_328,N_2983,N_2997);
and UO_329 (O_329,N_2973,N_2983);
or UO_330 (O_330,N_2985,N_2952);
or UO_331 (O_331,N_2973,N_2966);
and UO_332 (O_332,N_2953,N_2976);
nor UO_333 (O_333,N_2993,N_2952);
nor UO_334 (O_334,N_2960,N_2974);
xnor UO_335 (O_335,N_2952,N_2970);
nand UO_336 (O_336,N_2956,N_2997);
and UO_337 (O_337,N_2989,N_2961);
or UO_338 (O_338,N_2968,N_2992);
nand UO_339 (O_339,N_2951,N_2980);
nor UO_340 (O_340,N_2985,N_2953);
xnor UO_341 (O_341,N_2981,N_2990);
or UO_342 (O_342,N_2998,N_2966);
nor UO_343 (O_343,N_2953,N_2987);
nor UO_344 (O_344,N_2987,N_2976);
and UO_345 (O_345,N_2975,N_2978);
nand UO_346 (O_346,N_2983,N_2959);
xnor UO_347 (O_347,N_2961,N_2972);
or UO_348 (O_348,N_2971,N_2974);
and UO_349 (O_349,N_2981,N_2991);
nor UO_350 (O_350,N_2996,N_2957);
or UO_351 (O_351,N_2993,N_2986);
or UO_352 (O_352,N_2961,N_2994);
nand UO_353 (O_353,N_2957,N_2990);
or UO_354 (O_354,N_2972,N_2965);
nand UO_355 (O_355,N_2959,N_2998);
and UO_356 (O_356,N_2975,N_2951);
nor UO_357 (O_357,N_2981,N_2979);
nand UO_358 (O_358,N_2963,N_2998);
nand UO_359 (O_359,N_2951,N_2964);
and UO_360 (O_360,N_2979,N_2951);
or UO_361 (O_361,N_2950,N_2952);
or UO_362 (O_362,N_2955,N_2990);
nand UO_363 (O_363,N_2951,N_2974);
and UO_364 (O_364,N_2988,N_2963);
nor UO_365 (O_365,N_2965,N_2967);
nand UO_366 (O_366,N_2956,N_2990);
or UO_367 (O_367,N_2994,N_2964);
or UO_368 (O_368,N_2968,N_2983);
nand UO_369 (O_369,N_2969,N_2979);
and UO_370 (O_370,N_2970,N_2979);
and UO_371 (O_371,N_2954,N_2956);
or UO_372 (O_372,N_2965,N_2973);
or UO_373 (O_373,N_2959,N_2985);
nand UO_374 (O_374,N_2956,N_2989);
or UO_375 (O_375,N_2959,N_2973);
nor UO_376 (O_376,N_2998,N_2967);
or UO_377 (O_377,N_2957,N_2956);
and UO_378 (O_378,N_2952,N_2972);
or UO_379 (O_379,N_2991,N_2986);
and UO_380 (O_380,N_2960,N_2951);
nand UO_381 (O_381,N_2973,N_2956);
and UO_382 (O_382,N_2965,N_2975);
or UO_383 (O_383,N_2959,N_2958);
or UO_384 (O_384,N_2982,N_2965);
and UO_385 (O_385,N_2997,N_2988);
nor UO_386 (O_386,N_2976,N_2993);
nor UO_387 (O_387,N_2998,N_2987);
nor UO_388 (O_388,N_2979,N_2965);
and UO_389 (O_389,N_2979,N_2999);
nand UO_390 (O_390,N_2958,N_2963);
and UO_391 (O_391,N_2951,N_2950);
or UO_392 (O_392,N_2985,N_2980);
and UO_393 (O_393,N_2990,N_2979);
or UO_394 (O_394,N_2969,N_2999);
nor UO_395 (O_395,N_2960,N_2996);
nor UO_396 (O_396,N_2970,N_2963);
and UO_397 (O_397,N_2972,N_2975);
or UO_398 (O_398,N_2971,N_2991);
nor UO_399 (O_399,N_2971,N_2982);
nand UO_400 (O_400,N_2981,N_2973);
or UO_401 (O_401,N_2991,N_2968);
and UO_402 (O_402,N_2957,N_2981);
nor UO_403 (O_403,N_2996,N_2990);
xor UO_404 (O_404,N_2952,N_2978);
nand UO_405 (O_405,N_2987,N_2980);
or UO_406 (O_406,N_2977,N_2973);
and UO_407 (O_407,N_2980,N_2998);
nor UO_408 (O_408,N_2998,N_2971);
nand UO_409 (O_409,N_2970,N_2977);
or UO_410 (O_410,N_2954,N_2995);
nor UO_411 (O_411,N_2971,N_2953);
nor UO_412 (O_412,N_2992,N_2984);
nor UO_413 (O_413,N_2976,N_2999);
and UO_414 (O_414,N_2991,N_2989);
nor UO_415 (O_415,N_2985,N_2965);
nand UO_416 (O_416,N_2964,N_2979);
nand UO_417 (O_417,N_2981,N_2958);
nor UO_418 (O_418,N_2968,N_2984);
nand UO_419 (O_419,N_2964,N_2952);
or UO_420 (O_420,N_2968,N_2957);
or UO_421 (O_421,N_2961,N_2997);
nand UO_422 (O_422,N_2952,N_2969);
nor UO_423 (O_423,N_2987,N_2968);
nand UO_424 (O_424,N_2960,N_2964);
or UO_425 (O_425,N_2964,N_2971);
and UO_426 (O_426,N_2996,N_2954);
and UO_427 (O_427,N_2988,N_2972);
and UO_428 (O_428,N_2958,N_2964);
and UO_429 (O_429,N_2991,N_2963);
nor UO_430 (O_430,N_2950,N_2963);
nor UO_431 (O_431,N_2979,N_2961);
or UO_432 (O_432,N_2950,N_2973);
and UO_433 (O_433,N_2957,N_2984);
or UO_434 (O_434,N_2978,N_2982);
and UO_435 (O_435,N_2992,N_2956);
nand UO_436 (O_436,N_2980,N_2999);
and UO_437 (O_437,N_2968,N_2966);
and UO_438 (O_438,N_2959,N_2952);
nand UO_439 (O_439,N_2985,N_2975);
or UO_440 (O_440,N_2984,N_2989);
and UO_441 (O_441,N_2995,N_2994);
nand UO_442 (O_442,N_2961,N_2969);
or UO_443 (O_443,N_2956,N_2978);
nor UO_444 (O_444,N_2960,N_2997);
and UO_445 (O_445,N_2979,N_2997);
and UO_446 (O_446,N_2969,N_2975);
and UO_447 (O_447,N_2987,N_2955);
nor UO_448 (O_448,N_2985,N_2961);
or UO_449 (O_449,N_2991,N_2965);
or UO_450 (O_450,N_2965,N_2983);
nor UO_451 (O_451,N_2997,N_2959);
nor UO_452 (O_452,N_2980,N_2955);
nor UO_453 (O_453,N_2955,N_2981);
or UO_454 (O_454,N_2976,N_2997);
nand UO_455 (O_455,N_2995,N_2985);
or UO_456 (O_456,N_2958,N_2952);
and UO_457 (O_457,N_2965,N_2962);
or UO_458 (O_458,N_2959,N_2987);
or UO_459 (O_459,N_2950,N_2988);
nand UO_460 (O_460,N_2982,N_2983);
or UO_461 (O_461,N_2979,N_2950);
nand UO_462 (O_462,N_2999,N_2974);
nand UO_463 (O_463,N_2990,N_2980);
or UO_464 (O_464,N_2970,N_2965);
or UO_465 (O_465,N_2953,N_2997);
nor UO_466 (O_466,N_2988,N_2965);
nand UO_467 (O_467,N_2985,N_2977);
or UO_468 (O_468,N_2992,N_2954);
and UO_469 (O_469,N_2953,N_2979);
nand UO_470 (O_470,N_2957,N_2983);
nor UO_471 (O_471,N_2995,N_2963);
nor UO_472 (O_472,N_2951,N_2973);
and UO_473 (O_473,N_2962,N_2967);
and UO_474 (O_474,N_2963,N_2992);
nand UO_475 (O_475,N_2951,N_2953);
or UO_476 (O_476,N_2957,N_2950);
and UO_477 (O_477,N_2964,N_2977);
and UO_478 (O_478,N_2996,N_2959);
nand UO_479 (O_479,N_2957,N_2952);
or UO_480 (O_480,N_2961,N_2999);
nand UO_481 (O_481,N_2992,N_2980);
and UO_482 (O_482,N_2967,N_2984);
nand UO_483 (O_483,N_2969,N_2985);
nor UO_484 (O_484,N_2951,N_2999);
nor UO_485 (O_485,N_2976,N_2973);
and UO_486 (O_486,N_2960,N_2986);
and UO_487 (O_487,N_2977,N_2975);
or UO_488 (O_488,N_2984,N_2994);
or UO_489 (O_489,N_2987,N_2969);
and UO_490 (O_490,N_2977,N_2972);
and UO_491 (O_491,N_2997,N_2996);
nor UO_492 (O_492,N_2994,N_2989);
and UO_493 (O_493,N_2968,N_2982);
nand UO_494 (O_494,N_2951,N_2986);
nand UO_495 (O_495,N_2989,N_2975);
nand UO_496 (O_496,N_2951,N_2972);
nor UO_497 (O_497,N_2961,N_2968);
or UO_498 (O_498,N_2968,N_2962);
and UO_499 (O_499,N_2998,N_2994);
endmodule