module basic_750_5000_1000_25_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_293,In_576);
nand U1 (N_1,In_149,In_172);
nand U2 (N_2,In_747,In_409);
or U3 (N_3,In_197,In_243);
nor U4 (N_4,In_353,In_166);
nand U5 (N_5,In_402,In_464);
nor U6 (N_6,In_686,In_392);
or U7 (N_7,In_313,In_399);
nor U8 (N_8,In_514,In_400);
or U9 (N_9,In_126,In_196);
nand U10 (N_10,In_365,In_634);
and U11 (N_11,In_257,In_109);
nand U12 (N_12,In_667,In_596);
or U13 (N_13,In_411,In_419);
nand U14 (N_14,In_98,In_462);
and U15 (N_15,In_52,In_709);
nand U16 (N_16,In_61,In_454);
and U17 (N_17,In_473,In_532);
or U18 (N_18,In_2,In_696);
nor U19 (N_19,In_22,In_442);
and U20 (N_20,In_631,In_675);
or U21 (N_21,In_116,In_272);
or U22 (N_22,In_12,In_106);
nand U23 (N_23,In_512,In_190);
nor U24 (N_24,In_413,In_683);
or U25 (N_25,In_453,In_37);
nand U26 (N_26,In_628,In_32);
or U27 (N_27,In_223,In_232);
or U28 (N_28,In_387,In_296);
nor U29 (N_29,In_488,In_630);
and U30 (N_30,In_171,In_489);
nand U31 (N_31,In_26,In_498);
or U32 (N_32,In_134,In_440);
nand U33 (N_33,In_485,In_513);
nand U34 (N_34,In_508,In_10);
or U35 (N_35,In_352,In_209);
and U36 (N_36,In_550,In_502);
or U37 (N_37,In_282,In_523);
or U38 (N_38,In_7,In_671);
nor U39 (N_39,In_67,In_518);
nand U40 (N_40,In_715,In_378);
nor U41 (N_41,In_96,In_557);
nor U42 (N_42,In_469,In_122);
nor U43 (N_43,In_21,In_640);
nor U44 (N_44,In_139,In_565);
or U45 (N_45,In_541,In_48);
nor U46 (N_46,In_605,In_194);
or U47 (N_47,In_94,In_140);
nor U48 (N_48,In_129,In_414);
or U49 (N_49,In_570,In_704);
or U50 (N_50,In_688,In_620);
nand U51 (N_51,In_504,In_625);
and U52 (N_52,In_522,In_292);
nor U53 (N_53,In_707,In_8);
or U54 (N_54,In_213,In_653);
nand U55 (N_55,In_535,In_721);
and U56 (N_56,In_598,In_319);
or U57 (N_57,In_566,In_638);
nand U58 (N_58,In_58,In_0);
nor U59 (N_59,In_136,In_569);
and U60 (N_60,In_374,In_192);
nand U61 (N_61,In_644,In_115);
or U62 (N_62,In_57,In_538);
or U63 (N_63,In_274,In_158);
and U64 (N_64,In_597,In_314);
nand U65 (N_65,In_446,In_287);
nand U66 (N_66,In_626,In_348);
nand U67 (N_67,In_471,In_410);
nand U68 (N_68,In_280,In_269);
or U69 (N_69,In_177,In_678);
nor U70 (N_70,In_623,In_449);
nand U71 (N_71,In_66,In_334);
nand U72 (N_72,In_231,In_295);
or U73 (N_73,In_593,In_679);
or U74 (N_74,In_289,In_74);
nand U75 (N_75,In_216,In_635);
nor U76 (N_76,In_609,In_492);
nand U77 (N_77,In_191,In_568);
or U78 (N_78,In_36,In_380);
nor U79 (N_79,In_564,In_19);
and U80 (N_80,In_450,In_478);
and U81 (N_81,In_256,In_180);
nand U82 (N_82,In_349,In_415);
nor U83 (N_83,In_211,In_515);
or U84 (N_84,In_212,In_544);
or U85 (N_85,In_418,In_375);
xnor U86 (N_86,In_543,In_680);
nand U87 (N_87,In_80,In_712);
and U88 (N_88,In_340,In_746);
nand U89 (N_89,In_438,In_560);
and U90 (N_90,In_252,In_218);
and U91 (N_91,In_86,In_408);
nand U92 (N_92,In_719,In_416);
or U93 (N_93,In_713,In_341);
nand U94 (N_94,In_435,In_526);
or U95 (N_95,In_308,In_527);
and U96 (N_96,In_281,In_143);
or U97 (N_97,In_101,In_107);
or U98 (N_98,In_728,In_24);
nand U99 (N_99,In_244,In_494);
nor U100 (N_100,In_509,In_729);
and U101 (N_101,In_606,In_15);
nand U102 (N_102,In_674,In_738);
or U103 (N_103,In_481,In_639);
or U104 (N_104,In_29,In_84);
nor U105 (N_105,In_725,In_703);
or U106 (N_106,In_175,In_91);
nand U107 (N_107,In_451,In_322);
nor U108 (N_108,In_317,In_458);
and U109 (N_109,In_503,In_394);
nand U110 (N_110,In_384,In_441);
nor U111 (N_111,In_720,In_553);
nor U112 (N_112,In_137,In_506);
and U113 (N_113,In_382,In_370);
nor U114 (N_114,In_432,In_173);
nor U115 (N_115,In_693,In_682);
nand U116 (N_116,In_50,In_654);
and U117 (N_117,In_684,In_371);
nand U118 (N_118,In_663,In_737);
and U119 (N_119,In_25,In_176);
or U120 (N_120,In_562,In_239);
nor U121 (N_121,In_62,In_277);
and U122 (N_122,In_398,In_582);
or U123 (N_123,In_297,In_381);
or U124 (N_124,In_586,In_304);
or U125 (N_125,In_161,In_412);
nand U126 (N_126,In_230,In_210);
or U127 (N_127,In_363,In_16);
and U128 (N_128,In_629,In_55);
nor U129 (N_129,In_339,In_660);
nand U130 (N_130,In_439,In_561);
or U131 (N_131,In_595,In_3);
and U132 (N_132,In_480,In_141);
nand U133 (N_133,In_487,In_445);
nor U134 (N_134,In_236,In_283);
nand U135 (N_135,In_463,In_676);
or U136 (N_136,In_123,In_324);
and U137 (N_137,In_148,In_189);
nor U138 (N_138,In_266,In_315);
or U139 (N_139,In_132,In_602);
nand U140 (N_140,In_685,In_612);
or U141 (N_141,In_310,In_69);
or U142 (N_142,In_345,In_208);
nand U143 (N_143,In_6,In_227);
and U144 (N_144,In_429,In_649);
and U145 (N_145,In_475,In_336);
and U146 (N_146,In_40,In_695);
nor U147 (N_147,In_133,In_495);
or U148 (N_148,In_54,In_567);
and U149 (N_149,In_240,In_291);
nor U150 (N_150,In_155,In_53);
nand U151 (N_151,In_253,In_591);
nand U152 (N_152,In_534,In_611);
nor U153 (N_153,In_184,In_531);
and U154 (N_154,In_455,In_174);
or U155 (N_155,In_689,In_170);
nor U156 (N_156,In_732,In_650);
nand U157 (N_157,In_519,In_536);
and U158 (N_158,In_619,In_181);
nand U159 (N_159,In_298,In_431);
nor U160 (N_160,In_337,In_546);
and U161 (N_161,In_267,In_264);
or U162 (N_162,In_233,In_585);
and U163 (N_163,In_262,In_332);
nor U164 (N_164,In_436,In_539);
or U165 (N_165,In_670,In_367);
and U166 (N_166,In_470,In_162);
or U167 (N_167,In_320,In_112);
nand U168 (N_168,In_270,In_601);
nor U169 (N_169,In_219,In_658);
nor U170 (N_170,In_717,In_698);
nand U171 (N_171,In_205,In_376);
and U172 (N_172,In_554,In_364);
nor U173 (N_173,In_276,In_457);
nand U174 (N_174,In_27,In_119);
or U175 (N_175,In_130,In_311);
nor U176 (N_176,In_379,In_726);
or U177 (N_177,In_648,In_97);
nand U178 (N_178,In_479,In_486);
nor U179 (N_179,In_517,In_357);
and U180 (N_180,In_372,In_484);
and U181 (N_181,In_105,In_723);
nor U182 (N_182,In_202,In_497);
nand U183 (N_183,In_113,In_290);
and U184 (N_184,In_520,In_589);
nand U185 (N_185,In_714,In_579);
nand U186 (N_186,In_43,In_263);
and U187 (N_187,In_271,In_299);
nor U188 (N_188,In_393,In_499);
or U189 (N_189,In_745,In_248);
or U190 (N_190,In_433,In_187);
nor U191 (N_191,In_425,In_476);
or U192 (N_192,In_82,In_168);
and U193 (N_193,In_128,In_448);
or U194 (N_194,In_354,In_668);
and U195 (N_195,In_228,In_20);
nand U196 (N_196,In_103,In_120);
and U197 (N_197,In_700,In_42);
or U198 (N_198,In_571,In_138);
and U199 (N_199,In_511,In_1);
and U200 (N_200,N_196,In_551);
and U201 (N_201,In_603,N_160);
and U202 (N_202,In_691,In_330);
nor U203 (N_203,In_160,In_510);
and U204 (N_204,N_199,In_305);
nor U205 (N_205,N_176,N_42);
xor U206 (N_206,In_246,In_92);
nand U207 (N_207,In_373,N_156);
and U208 (N_208,In_427,N_192);
and U209 (N_209,N_44,N_103);
nor U210 (N_210,In_739,In_18);
and U211 (N_211,In_328,In_124);
or U212 (N_212,In_724,N_20);
and U213 (N_213,In_258,N_70);
xor U214 (N_214,In_377,N_92);
nor U215 (N_215,N_56,In_241);
nor U216 (N_216,In_51,In_102);
and U217 (N_217,In_45,N_146);
and U218 (N_218,In_238,In_659);
and U219 (N_219,In_617,In_677);
nor U220 (N_220,In_718,In_744);
or U221 (N_221,In_577,In_616);
and U222 (N_222,N_165,In_355);
or U223 (N_223,N_126,In_154);
nor U224 (N_224,In_87,N_65);
nand U225 (N_225,In_749,In_386);
nand U226 (N_226,N_178,N_124);
nand U227 (N_227,N_141,In_95);
or U228 (N_228,N_57,In_636);
and U229 (N_229,N_169,N_120);
or U230 (N_230,In_11,N_136);
nand U231 (N_231,In_548,In_261);
nor U232 (N_232,N_6,In_188);
or U233 (N_233,N_43,In_607);
nand U234 (N_234,In_613,In_383);
nor U235 (N_235,In_641,N_151);
or U236 (N_236,In_642,In_655);
nand U237 (N_237,N_24,In_615);
nor U238 (N_238,N_171,N_123);
or U239 (N_239,N_61,In_474);
and U240 (N_240,N_22,In_4);
nor U241 (N_241,In_59,In_88);
and U242 (N_242,N_99,N_168);
and U243 (N_243,In_279,In_77);
nand U244 (N_244,In_286,In_574);
and U245 (N_245,In_83,In_563);
nor U246 (N_246,In_63,N_180);
nor U247 (N_247,In_652,N_79);
nand U248 (N_248,In_23,N_100);
and U249 (N_249,In_403,N_164);
or U250 (N_250,In_633,N_167);
and U251 (N_251,In_41,In_198);
or U252 (N_252,N_132,In_316);
nand U253 (N_253,In_145,N_114);
nand U254 (N_254,N_26,In_199);
or U255 (N_255,N_197,N_163);
nor U256 (N_256,N_1,In_70);
or U257 (N_257,In_588,In_621);
or U258 (N_258,N_187,In_666);
or U259 (N_259,In_235,In_608);
nand U260 (N_260,In_742,N_135);
nand U261 (N_261,In_524,In_28);
nand U262 (N_262,In_207,In_420);
nand U263 (N_263,In_366,In_285);
or U264 (N_264,In_60,N_2);
and U265 (N_265,In_467,N_38);
or U266 (N_266,In_251,N_31);
and U267 (N_267,In_100,In_333);
nor U268 (N_268,In_301,In_278);
or U269 (N_269,In_443,N_148);
nor U270 (N_270,In_220,In_396);
nand U271 (N_271,In_627,N_127);
or U272 (N_272,In_584,N_119);
or U273 (N_273,In_482,N_69);
and U274 (N_274,N_53,N_64);
and U275 (N_275,In_590,In_34);
or U276 (N_276,N_32,In_552);
and U277 (N_277,In_423,N_181);
or U278 (N_278,N_109,In_156);
nand U279 (N_279,N_45,In_163);
nand U280 (N_280,In_672,In_89);
nand U281 (N_281,N_162,In_662);
and U282 (N_282,In_637,In_39);
nand U283 (N_283,In_369,In_104);
nand U284 (N_284,In_558,In_645);
nand U285 (N_285,N_66,N_55);
or U286 (N_286,N_3,N_86);
and U287 (N_287,In_385,In_159);
nand U288 (N_288,In_131,In_669);
nor U289 (N_289,N_125,In_705);
or U290 (N_290,N_183,In_193);
nand U291 (N_291,In_710,N_128);
nand U292 (N_292,In_323,In_401);
or U293 (N_293,In_73,In_533);
or U294 (N_294,N_71,N_52);
or U295 (N_295,In_362,In_144);
or U296 (N_296,In_730,In_748);
nand U297 (N_297,In_165,N_186);
nand U298 (N_298,N_130,N_84);
nor U299 (N_299,In_643,In_444);
nand U300 (N_300,In_150,N_191);
nor U301 (N_301,In_245,N_46);
or U302 (N_302,In_731,In_356);
nor U303 (N_303,N_108,N_21);
or U304 (N_304,N_139,In_581);
and U305 (N_305,In_306,In_434);
and U306 (N_306,N_90,In_72);
nand U307 (N_307,N_4,N_85);
nor U308 (N_308,N_15,In_578);
or U309 (N_309,In_632,In_618);
nor U310 (N_310,N_102,In_583);
and U311 (N_311,In_335,In_234);
and U312 (N_312,In_716,In_247);
and U313 (N_313,In_575,In_14);
or U314 (N_314,N_110,N_145);
or U315 (N_315,N_76,In_651);
nand U316 (N_316,N_8,N_134);
and U317 (N_317,N_188,In_456);
and U318 (N_318,N_159,In_195);
nand U319 (N_319,In_447,In_201);
nor U320 (N_320,In_351,N_101);
and U321 (N_321,In_147,N_144);
and U322 (N_322,N_88,In_17);
nor U323 (N_323,In_13,In_587);
nand U324 (N_324,In_549,N_11);
nand U325 (N_325,In_275,N_9);
and U326 (N_326,In_214,N_154);
and U327 (N_327,In_203,N_10);
and U328 (N_328,In_390,N_33);
and U329 (N_329,In_344,In_342);
and U330 (N_330,In_624,N_170);
nor U331 (N_331,N_51,In_38);
nor U332 (N_332,In_326,In_422);
or U333 (N_333,In_559,In_225);
nor U334 (N_334,In_388,N_62);
and U335 (N_335,In_664,In_312);
nor U336 (N_336,In_490,N_67);
nor U337 (N_337,In_483,In_259);
nand U338 (N_338,N_25,In_226);
or U339 (N_339,In_260,N_174);
nand U340 (N_340,N_182,N_49);
nand U341 (N_341,In_360,In_516);
and U342 (N_342,In_33,In_708);
nor U343 (N_343,In_350,N_118);
or U344 (N_344,N_94,N_34);
and U345 (N_345,N_12,In_78);
and U346 (N_346,In_646,N_89);
or U347 (N_347,In_507,In_540);
nor U348 (N_348,In_665,N_16);
or U349 (N_349,In_76,N_98);
nand U350 (N_350,In_318,In_182);
nor U351 (N_351,N_58,In_85);
nor U352 (N_352,In_31,N_13);
nor U353 (N_353,In_229,In_417);
or U354 (N_354,In_254,In_421);
nand U355 (N_355,In_65,In_547);
nor U356 (N_356,In_204,N_39);
or U357 (N_357,N_111,In_224);
nor U358 (N_358,In_465,N_184);
or U359 (N_359,N_72,In_206);
and U360 (N_360,N_28,In_610);
or U361 (N_361,N_19,In_200);
nand U362 (N_362,In_740,In_706);
nor U363 (N_363,In_542,N_81);
and U364 (N_364,In_284,N_5);
nor U365 (N_365,In_68,In_30);
nor U366 (N_366,In_321,In_300);
nand U367 (N_367,N_105,In_529);
nor U368 (N_368,In_500,N_194);
and U369 (N_369,N_37,In_167);
nand U370 (N_370,In_501,N_175);
and U371 (N_371,N_35,In_169);
nor U372 (N_372,N_14,N_190);
and U373 (N_373,In_64,N_117);
and U374 (N_374,In_426,In_268);
and U375 (N_375,In_397,N_121);
or U376 (N_376,In_699,In_329);
and U377 (N_377,N_193,In_657);
or U378 (N_378,In_505,N_122);
and U379 (N_379,In_90,N_95);
or U380 (N_380,In_164,In_125);
and U381 (N_381,In_250,In_604);
nand U382 (N_382,N_140,In_521);
nor U383 (N_383,N_68,In_359);
and U384 (N_384,In_594,N_198);
or U385 (N_385,In_302,N_47);
nand U386 (N_386,In_249,N_173);
nand U387 (N_387,In_118,In_142);
and U388 (N_388,In_325,N_96);
nand U389 (N_389,In_309,N_112);
nor U390 (N_390,In_44,In_430);
and U391 (N_391,N_131,N_115);
or U392 (N_392,In_157,In_466);
nor U393 (N_393,N_138,N_87);
and U394 (N_394,N_97,In_528);
or U395 (N_395,N_93,In_153);
nand U396 (N_396,In_47,N_143);
or U397 (N_397,In_110,N_116);
nand U398 (N_398,N_91,In_237);
nand U399 (N_399,N_189,N_29);
and U400 (N_400,N_258,N_23);
or U401 (N_401,N_236,In_687);
nand U402 (N_402,In_461,N_338);
or U403 (N_403,N_331,N_353);
nor U404 (N_404,N_241,N_217);
and U405 (N_405,N_266,In_599);
nor U406 (N_406,N_200,N_356);
nand U407 (N_407,In_46,N_289);
and U408 (N_408,In_580,N_265);
nand U409 (N_409,N_395,In_733);
nor U410 (N_410,N_208,N_272);
and U411 (N_411,In_491,N_161);
nand U412 (N_412,In_735,In_673);
and U413 (N_413,In_572,In_727);
and U414 (N_414,N_80,In_75);
nor U415 (N_415,N_17,N_351);
and U416 (N_416,N_303,N_291);
nor U417 (N_417,N_295,N_36);
or U418 (N_418,N_239,N_367);
and U419 (N_419,In_690,N_300);
or U420 (N_420,N_365,N_7);
and U421 (N_421,In_346,N_388);
nor U422 (N_422,In_459,N_259);
and U423 (N_423,In_114,N_73);
nand U424 (N_424,N_363,N_249);
nor U425 (N_425,N_344,N_333);
and U426 (N_426,In_151,In_146);
nor U427 (N_427,In_99,N_220);
nand U428 (N_428,In_391,In_294);
nand U429 (N_429,N_314,N_390);
or U430 (N_430,N_210,N_381);
or U431 (N_431,In_681,N_166);
and U432 (N_432,N_346,In_656);
nand U433 (N_433,In_743,In_273);
and U434 (N_434,N_288,N_347);
and U435 (N_435,N_375,N_30);
or U436 (N_436,N_271,N_306);
and U437 (N_437,In_472,N_230);
or U438 (N_438,In_395,N_292);
nor U439 (N_439,N_231,N_153);
nor U440 (N_440,N_370,N_238);
nand U441 (N_441,In_347,N_325);
nand U442 (N_442,In_81,N_77);
and U443 (N_443,N_229,N_224);
nand U444 (N_444,N_219,N_234);
and U445 (N_445,N_252,N_104);
or U446 (N_446,N_225,N_316);
nand U447 (N_447,N_255,N_279);
nand U448 (N_448,N_386,N_348);
nand U449 (N_449,In_614,In_405);
nor U450 (N_450,N_275,N_273);
nor U451 (N_451,In_452,N_343);
or U452 (N_452,N_318,N_205);
nand U453 (N_453,In_741,N_142);
nand U454 (N_454,In_530,N_0);
or U455 (N_455,In_179,In_56);
nor U456 (N_456,In_121,N_328);
or U457 (N_457,N_250,N_382);
and U458 (N_458,N_216,N_380);
nor U459 (N_459,N_358,N_397);
nand U460 (N_460,In_178,In_437);
and U461 (N_461,In_331,N_357);
and U462 (N_462,N_277,N_221);
or U463 (N_463,N_297,In_186);
or U464 (N_464,N_232,N_309);
or U465 (N_465,In_555,N_281);
nand U466 (N_466,N_133,In_5);
nand U467 (N_467,In_711,N_322);
or U468 (N_468,N_147,In_222);
nor U469 (N_469,In_468,N_399);
or U470 (N_470,N_74,In_525);
nand U471 (N_471,N_327,N_362);
or U472 (N_472,N_63,N_263);
nand U473 (N_473,N_237,N_366);
nor U474 (N_474,N_260,In_79);
and U475 (N_475,N_329,N_195);
or U476 (N_476,N_280,N_284);
nand U477 (N_477,N_50,N_227);
nand U478 (N_478,N_377,N_319);
or U479 (N_479,In_361,N_340);
nand U480 (N_480,N_257,N_78);
nand U481 (N_481,N_209,N_206);
and U482 (N_482,N_312,N_387);
nor U483 (N_483,In_692,N_394);
or U484 (N_484,N_359,N_372);
nor U485 (N_485,N_323,In_592);
or U486 (N_486,N_83,N_203);
xor U487 (N_487,N_293,N_149);
and U488 (N_488,In_183,N_317);
nor U489 (N_489,In_493,In_343);
nand U490 (N_490,N_245,N_296);
nor U491 (N_491,In_288,N_313);
nand U492 (N_492,N_256,In_477);
or U493 (N_493,N_212,N_341);
or U494 (N_494,In_389,N_321);
or U495 (N_495,In_127,N_228);
or U496 (N_496,N_267,N_305);
or U497 (N_497,N_244,N_251);
and U498 (N_498,N_207,N_48);
or U499 (N_499,In_600,N_215);
or U500 (N_500,N_82,N_150);
and U501 (N_501,N_285,In_702);
nand U502 (N_502,N_307,N_389);
nand U503 (N_503,N_376,N_233);
and U504 (N_504,N_276,N_27);
or U505 (N_505,N_301,N_214);
nand U506 (N_506,In_307,In_255);
nor U507 (N_507,In_428,In_694);
nor U508 (N_508,In_573,N_177);
nor U509 (N_509,In_71,N_18);
nor U510 (N_510,N_222,In_358);
or U511 (N_511,N_352,In_93);
or U512 (N_512,N_286,N_339);
nand U513 (N_513,N_211,N_315);
or U514 (N_514,In_215,In_338);
nor U515 (N_515,N_213,N_294);
and U516 (N_516,In_722,In_556);
nor U517 (N_517,In_35,In_406);
nand U518 (N_518,N_385,N_242);
nor U519 (N_519,N_157,N_360);
and U520 (N_520,N_373,In_327);
and U521 (N_521,N_113,In_185);
nand U522 (N_522,N_158,N_330);
or U523 (N_523,N_247,N_226);
or U524 (N_524,N_383,N_240);
nor U525 (N_525,N_218,N_172);
nor U526 (N_526,In_424,N_392);
xor U527 (N_527,N_155,N_396);
or U528 (N_528,N_282,In_111);
or U529 (N_529,N_299,In_622);
nor U530 (N_530,In_49,In_303);
and U531 (N_531,In_701,In_496);
or U532 (N_532,N_398,N_246);
nor U533 (N_533,In_242,In_404);
nor U534 (N_534,N_254,N_202);
and U535 (N_535,N_334,In_697);
or U536 (N_536,In_368,N_379);
nand U537 (N_537,N_369,N_253);
and U538 (N_538,N_345,N_106);
nor U539 (N_539,N_54,In_135);
nand U540 (N_540,N_261,N_204);
and U541 (N_541,N_290,N_264);
and U542 (N_542,N_201,N_75);
nand U543 (N_543,In_661,N_223);
nor U544 (N_544,N_324,N_368);
nor U545 (N_545,N_311,N_278);
nand U546 (N_546,N_350,N_378);
nand U547 (N_547,N_320,N_355);
xor U548 (N_548,N_374,N_248);
xnor U549 (N_549,N_371,N_137);
and U550 (N_550,In_221,In_545);
and U551 (N_551,N_304,N_335);
nor U552 (N_552,N_262,In_108);
or U553 (N_553,N_274,N_129);
nor U554 (N_554,N_243,In_460);
nor U555 (N_555,N_310,In_537);
nand U556 (N_556,N_336,N_269);
and U557 (N_557,In_9,In_152);
nand U558 (N_558,N_302,N_349);
nor U559 (N_559,N_326,N_268);
nor U560 (N_560,In_736,N_287);
nand U561 (N_561,N_332,In_217);
and U562 (N_562,N_361,N_235);
or U563 (N_563,N_354,N_107);
and U564 (N_564,N_283,N_40);
or U565 (N_565,N_60,N_364);
nand U566 (N_566,In_117,N_41);
nand U567 (N_567,N_152,N_384);
nor U568 (N_568,In_407,N_337);
and U569 (N_569,N_391,N_59);
nand U570 (N_570,N_185,N_342);
or U571 (N_571,In_265,In_647);
nand U572 (N_572,N_179,N_298);
nand U573 (N_573,N_393,N_308);
nand U574 (N_574,In_734,N_270);
nand U575 (N_575,In_222,N_254);
nor U576 (N_576,In_111,N_373);
nand U577 (N_577,N_360,In_217);
nand U578 (N_578,N_350,In_294);
and U579 (N_579,N_205,In_288);
nor U580 (N_580,In_661,In_255);
and U581 (N_581,N_224,In_331);
or U582 (N_582,In_572,N_246);
and U583 (N_583,In_361,N_63);
nor U584 (N_584,In_221,N_278);
or U585 (N_585,N_268,In_35);
nand U586 (N_586,N_155,In_734);
or U587 (N_587,N_281,N_217);
xnor U588 (N_588,N_350,N_253);
nand U589 (N_589,N_73,N_306);
nor U590 (N_590,N_294,In_49);
nor U591 (N_591,In_545,N_275);
nor U592 (N_592,N_367,In_530);
and U593 (N_593,In_661,N_201);
nor U594 (N_594,In_461,N_249);
nor U595 (N_595,In_687,N_368);
and U596 (N_596,In_406,N_277);
nand U597 (N_597,N_323,N_266);
nand U598 (N_598,In_733,N_333);
or U599 (N_599,N_209,In_121);
nor U600 (N_600,N_554,N_441);
nor U601 (N_601,N_433,N_431);
nand U602 (N_602,N_513,N_591);
and U603 (N_603,N_411,N_409);
or U604 (N_604,N_527,N_518);
nor U605 (N_605,N_510,N_501);
nor U606 (N_606,N_559,N_484);
nand U607 (N_607,N_438,N_564);
nand U608 (N_608,N_516,N_524);
and U609 (N_609,N_592,N_486);
xor U610 (N_610,N_556,N_493);
nor U611 (N_611,N_577,N_598);
nor U612 (N_612,N_440,N_508);
nor U613 (N_613,N_422,N_545);
nand U614 (N_614,N_580,N_490);
nor U615 (N_615,N_473,N_407);
or U616 (N_616,N_520,N_595);
and U617 (N_617,N_412,N_487);
or U618 (N_618,N_504,N_555);
or U619 (N_619,N_457,N_472);
nor U620 (N_620,N_413,N_435);
nor U621 (N_621,N_528,N_464);
or U622 (N_622,N_587,N_567);
nand U623 (N_623,N_400,N_405);
or U624 (N_624,N_455,N_525);
or U625 (N_625,N_542,N_461);
or U626 (N_626,N_563,N_427);
or U627 (N_627,N_477,N_537);
or U628 (N_628,N_458,N_467);
nand U629 (N_629,N_459,N_443);
nand U630 (N_630,N_583,N_492);
xor U631 (N_631,N_565,N_446);
and U632 (N_632,N_454,N_415);
nand U633 (N_633,N_538,N_535);
nor U634 (N_634,N_489,N_581);
nand U635 (N_635,N_485,N_588);
nand U636 (N_636,N_590,N_529);
nand U637 (N_637,N_522,N_406);
or U638 (N_638,N_566,N_579);
nand U639 (N_639,N_517,N_449);
or U640 (N_640,N_582,N_552);
or U641 (N_641,N_547,N_476);
and U642 (N_642,N_557,N_442);
nand U643 (N_643,N_465,N_423);
and U644 (N_644,N_597,N_499);
nand U645 (N_645,N_507,N_491);
nand U646 (N_646,N_421,N_483);
or U647 (N_647,N_434,N_462);
nor U648 (N_648,N_539,N_551);
nor U649 (N_649,N_479,N_426);
and U650 (N_650,N_550,N_512);
and U651 (N_651,N_502,N_404);
and U652 (N_652,N_451,N_488);
nor U653 (N_653,N_466,N_578);
or U654 (N_654,N_474,N_469);
and U655 (N_655,N_543,N_568);
or U656 (N_656,N_573,N_445);
nor U657 (N_657,N_500,N_589);
nor U658 (N_658,N_439,N_478);
or U659 (N_659,N_436,N_561);
and U660 (N_660,N_414,N_560);
or U661 (N_661,N_428,N_541);
nor U662 (N_662,N_585,N_594);
or U663 (N_663,N_599,N_570);
nand U664 (N_664,N_584,N_403);
and U665 (N_665,N_497,N_509);
and U666 (N_666,N_546,N_470);
or U667 (N_667,N_417,N_514);
nand U668 (N_668,N_515,N_429);
nand U669 (N_669,N_544,N_530);
xor U670 (N_670,N_430,N_549);
and U671 (N_671,N_495,N_437);
and U672 (N_672,N_519,N_408);
nand U673 (N_673,N_416,N_419);
nand U674 (N_674,N_534,N_410);
and U675 (N_675,N_432,N_463);
or U676 (N_676,N_468,N_540);
nor U677 (N_677,N_576,N_575);
xor U678 (N_678,N_553,N_526);
and U679 (N_679,N_456,N_548);
or U680 (N_680,N_569,N_521);
or U681 (N_681,N_460,N_523);
and U682 (N_682,N_532,N_471);
and U683 (N_683,N_506,N_571);
nor U684 (N_684,N_572,N_533);
or U685 (N_685,N_503,N_482);
nand U686 (N_686,N_574,N_494);
nor U687 (N_687,N_452,N_531);
and U688 (N_688,N_498,N_401);
nor U689 (N_689,N_450,N_424);
nor U690 (N_690,N_593,N_586);
or U691 (N_691,N_596,N_505);
and U692 (N_692,N_481,N_420);
or U693 (N_693,N_511,N_562);
nand U694 (N_694,N_480,N_558);
nand U695 (N_695,N_496,N_425);
and U696 (N_696,N_453,N_447);
nor U697 (N_697,N_448,N_402);
nand U698 (N_698,N_536,N_475);
nor U699 (N_699,N_444,N_418);
or U700 (N_700,N_481,N_594);
or U701 (N_701,N_586,N_549);
or U702 (N_702,N_557,N_479);
nor U703 (N_703,N_450,N_556);
or U704 (N_704,N_476,N_481);
and U705 (N_705,N_591,N_500);
or U706 (N_706,N_579,N_421);
or U707 (N_707,N_406,N_458);
nand U708 (N_708,N_400,N_595);
or U709 (N_709,N_482,N_439);
nor U710 (N_710,N_466,N_409);
and U711 (N_711,N_427,N_599);
or U712 (N_712,N_583,N_498);
or U713 (N_713,N_442,N_576);
nor U714 (N_714,N_491,N_511);
nand U715 (N_715,N_475,N_467);
or U716 (N_716,N_507,N_485);
nor U717 (N_717,N_584,N_474);
and U718 (N_718,N_514,N_475);
nand U719 (N_719,N_420,N_552);
nor U720 (N_720,N_454,N_469);
xnor U721 (N_721,N_418,N_469);
nand U722 (N_722,N_586,N_542);
nor U723 (N_723,N_507,N_419);
and U724 (N_724,N_417,N_511);
nand U725 (N_725,N_587,N_458);
nand U726 (N_726,N_577,N_555);
or U727 (N_727,N_437,N_430);
nor U728 (N_728,N_497,N_575);
and U729 (N_729,N_437,N_527);
nor U730 (N_730,N_546,N_457);
nor U731 (N_731,N_505,N_462);
nor U732 (N_732,N_472,N_576);
nand U733 (N_733,N_538,N_465);
or U734 (N_734,N_533,N_445);
nand U735 (N_735,N_447,N_436);
or U736 (N_736,N_589,N_414);
and U737 (N_737,N_426,N_541);
and U738 (N_738,N_444,N_599);
or U739 (N_739,N_443,N_435);
nand U740 (N_740,N_489,N_509);
or U741 (N_741,N_550,N_468);
nand U742 (N_742,N_431,N_468);
or U743 (N_743,N_517,N_505);
and U744 (N_744,N_550,N_504);
or U745 (N_745,N_557,N_481);
or U746 (N_746,N_488,N_440);
nor U747 (N_747,N_434,N_470);
xnor U748 (N_748,N_403,N_480);
and U749 (N_749,N_402,N_511);
nand U750 (N_750,N_401,N_532);
or U751 (N_751,N_583,N_448);
nor U752 (N_752,N_453,N_518);
nor U753 (N_753,N_480,N_459);
nor U754 (N_754,N_579,N_451);
and U755 (N_755,N_513,N_413);
and U756 (N_756,N_444,N_438);
nand U757 (N_757,N_478,N_524);
nand U758 (N_758,N_533,N_511);
nand U759 (N_759,N_521,N_460);
nor U760 (N_760,N_492,N_587);
or U761 (N_761,N_589,N_568);
nand U762 (N_762,N_569,N_588);
and U763 (N_763,N_553,N_573);
and U764 (N_764,N_594,N_577);
nand U765 (N_765,N_491,N_520);
nor U766 (N_766,N_501,N_447);
or U767 (N_767,N_425,N_551);
or U768 (N_768,N_593,N_520);
or U769 (N_769,N_544,N_586);
or U770 (N_770,N_562,N_464);
or U771 (N_771,N_533,N_579);
or U772 (N_772,N_514,N_423);
and U773 (N_773,N_599,N_438);
xnor U774 (N_774,N_587,N_558);
nor U775 (N_775,N_406,N_444);
and U776 (N_776,N_414,N_463);
and U777 (N_777,N_541,N_587);
nor U778 (N_778,N_569,N_564);
or U779 (N_779,N_576,N_514);
or U780 (N_780,N_587,N_559);
or U781 (N_781,N_483,N_428);
or U782 (N_782,N_455,N_574);
or U783 (N_783,N_484,N_473);
and U784 (N_784,N_420,N_542);
nor U785 (N_785,N_414,N_500);
or U786 (N_786,N_559,N_477);
or U787 (N_787,N_480,N_567);
and U788 (N_788,N_419,N_483);
nor U789 (N_789,N_413,N_599);
nand U790 (N_790,N_493,N_548);
nor U791 (N_791,N_571,N_464);
nor U792 (N_792,N_569,N_553);
and U793 (N_793,N_504,N_557);
nand U794 (N_794,N_414,N_453);
and U795 (N_795,N_402,N_473);
and U796 (N_796,N_407,N_500);
nand U797 (N_797,N_491,N_518);
nor U798 (N_798,N_530,N_519);
and U799 (N_799,N_567,N_494);
nand U800 (N_800,N_792,N_795);
nor U801 (N_801,N_748,N_708);
nor U802 (N_802,N_674,N_619);
nor U803 (N_803,N_760,N_740);
nor U804 (N_804,N_762,N_625);
or U805 (N_805,N_682,N_673);
nand U806 (N_806,N_735,N_722);
and U807 (N_807,N_796,N_645);
nor U808 (N_808,N_692,N_771);
or U809 (N_809,N_607,N_642);
or U810 (N_810,N_749,N_777);
xor U811 (N_811,N_773,N_661);
nor U812 (N_812,N_641,N_744);
or U813 (N_813,N_751,N_711);
nand U814 (N_814,N_780,N_624);
nand U815 (N_815,N_772,N_649);
nand U816 (N_816,N_681,N_732);
or U817 (N_817,N_791,N_782);
and U818 (N_818,N_669,N_626);
or U819 (N_819,N_657,N_739);
xnor U820 (N_820,N_761,N_654);
nand U821 (N_821,N_627,N_710);
nand U822 (N_822,N_726,N_724);
and U823 (N_823,N_629,N_653);
and U824 (N_824,N_754,N_636);
nand U825 (N_825,N_755,N_676);
or U826 (N_826,N_769,N_737);
or U827 (N_827,N_746,N_701);
nand U828 (N_828,N_656,N_672);
nor U829 (N_829,N_721,N_664);
or U830 (N_830,N_678,N_714);
nand U831 (N_831,N_610,N_717);
nand U832 (N_832,N_774,N_671);
or U833 (N_833,N_750,N_702);
nand U834 (N_834,N_757,N_712);
nor U835 (N_835,N_727,N_639);
nor U836 (N_836,N_734,N_693);
nor U837 (N_837,N_675,N_763);
or U838 (N_838,N_686,N_652);
nand U839 (N_839,N_747,N_781);
or U840 (N_840,N_759,N_666);
or U841 (N_841,N_600,N_770);
nor U842 (N_842,N_731,N_696);
nor U843 (N_843,N_650,N_784);
or U844 (N_844,N_709,N_703);
nor U845 (N_845,N_799,N_758);
nand U846 (N_846,N_677,N_638);
nand U847 (N_847,N_786,N_643);
nand U848 (N_848,N_658,N_651);
or U849 (N_849,N_706,N_659);
or U850 (N_850,N_715,N_690);
nor U851 (N_851,N_668,N_623);
and U852 (N_852,N_628,N_768);
or U853 (N_853,N_662,N_718);
and U854 (N_854,N_753,N_707);
or U855 (N_855,N_633,N_640);
or U856 (N_856,N_660,N_679);
nor U857 (N_857,N_743,N_602);
and U858 (N_858,N_601,N_797);
nor U859 (N_859,N_729,N_745);
nand U860 (N_860,N_765,N_631);
and U861 (N_861,N_635,N_752);
and U862 (N_862,N_788,N_608);
nand U863 (N_863,N_719,N_697);
nor U864 (N_864,N_728,N_670);
or U865 (N_865,N_720,N_616);
or U866 (N_866,N_646,N_783);
or U867 (N_867,N_667,N_775);
or U868 (N_868,N_716,N_700);
nand U869 (N_869,N_611,N_680);
nand U870 (N_870,N_766,N_794);
or U871 (N_871,N_609,N_764);
and U872 (N_872,N_689,N_699);
or U873 (N_873,N_685,N_742);
or U874 (N_874,N_606,N_778);
or U875 (N_875,N_798,N_756);
and U876 (N_876,N_691,N_790);
and U877 (N_877,N_713,N_603);
or U878 (N_878,N_644,N_698);
nand U879 (N_879,N_621,N_665);
nand U880 (N_880,N_684,N_632);
nor U881 (N_881,N_655,N_695);
or U882 (N_882,N_620,N_787);
or U883 (N_883,N_618,N_683);
and U884 (N_884,N_694,N_704);
and U885 (N_885,N_617,N_604);
nor U886 (N_886,N_688,N_725);
or U887 (N_887,N_647,N_730);
or U888 (N_888,N_613,N_738);
or U889 (N_889,N_779,N_605);
nand U890 (N_890,N_741,N_630);
nor U891 (N_891,N_615,N_767);
or U892 (N_892,N_789,N_614);
and U893 (N_893,N_733,N_663);
nor U894 (N_894,N_723,N_705);
and U895 (N_895,N_736,N_622);
and U896 (N_896,N_776,N_637);
and U897 (N_897,N_612,N_785);
or U898 (N_898,N_687,N_648);
or U899 (N_899,N_634,N_793);
nor U900 (N_900,N_734,N_624);
and U901 (N_901,N_687,N_617);
nor U902 (N_902,N_606,N_763);
or U903 (N_903,N_787,N_714);
and U904 (N_904,N_631,N_711);
nor U905 (N_905,N_619,N_600);
or U906 (N_906,N_795,N_651);
and U907 (N_907,N_619,N_690);
nand U908 (N_908,N_728,N_796);
nor U909 (N_909,N_640,N_737);
nor U910 (N_910,N_604,N_709);
and U911 (N_911,N_670,N_716);
xnor U912 (N_912,N_600,N_650);
xor U913 (N_913,N_660,N_721);
or U914 (N_914,N_741,N_680);
and U915 (N_915,N_695,N_798);
and U916 (N_916,N_722,N_669);
and U917 (N_917,N_710,N_693);
or U918 (N_918,N_657,N_737);
and U919 (N_919,N_678,N_771);
nand U920 (N_920,N_636,N_611);
or U921 (N_921,N_719,N_732);
and U922 (N_922,N_727,N_611);
nand U923 (N_923,N_637,N_737);
nor U924 (N_924,N_605,N_623);
nand U925 (N_925,N_689,N_775);
nor U926 (N_926,N_627,N_624);
nand U927 (N_927,N_787,N_660);
nand U928 (N_928,N_759,N_615);
nor U929 (N_929,N_621,N_743);
nor U930 (N_930,N_788,N_657);
or U931 (N_931,N_710,N_765);
nor U932 (N_932,N_750,N_647);
or U933 (N_933,N_788,N_747);
or U934 (N_934,N_754,N_701);
or U935 (N_935,N_601,N_760);
nand U936 (N_936,N_646,N_715);
and U937 (N_937,N_624,N_735);
and U938 (N_938,N_731,N_724);
or U939 (N_939,N_645,N_765);
or U940 (N_940,N_712,N_731);
nor U941 (N_941,N_700,N_791);
or U942 (N_942,N_655,N_768);
and U943 (N_943,N_724,N_671);
or U944 (N_944,N_677,N_770);
xor U945 (N_945,N_637,N_665);
nor U946 (N_946,N_656,N_616);
or U947 (N_947,N_769,N_766);
nand U948 (N_948,N_777,N_657);
nand U949 (N_949,N_656,N_668);
nand U950 (N_950,N_602,N_618);
or U951 (N_951,N_665,N_604);
and U952 (N_952,N_731,N_638);
and U953 (N_953,N_798,N_626);
or U954 (N_954,N_648,N_622);
nand U955 (N_955,N_705,N_714);
nand U956 (N_956,N_735,N_754);
nor U957 (N_957,N_793,N_621);
nor U958 (N_958,N_787,N_618);
nand U959 (N_959,N_748,N_627);
or U960 (N_960,N_746,N_665);
and U961 (N_961,N_778,N_675);
and U962 (N_962,N_662,N_613);
or U963 (N_963,N_657,N_640);
and U964 (N_964,N_702,N_700);
and U965 (N_965,N_730,N_684);
nor U966 (N_966,N_677,N_602);
and U967 (N_967,N_786,N_695);
nor U968 (N_968,N_712,N_621);
nor U969 (N_969,N_629,N_678);
nor U970 (N_970,N_655,N_769);
and U971 (N_971,N_671,N_691);
and U972 (N_972,N_665,N_755);
and U973 (N_973,N_788,N_755);
nand U974 (N_974,N_717,N_754);
nor U975 (N_975,N_606,N_733);
and U976 (N_976,N_731,N_607);
or U977 (N_977,N_747,N_720);
xor U978 (N_978,N_674,N_728);
or U979 (N_979,N_647,N_723);
or U980 (N_980,N_615,N_763);
and U981 (N_981,N_652,N_659);
or U982 (N_982,N_748,N_736);
and U983 (N_983,N_752,N_711);
or U984 (N_984,N_760,N_789);
and U985 (N_985,N_638,N_764);
or U986 (N_986,N_752,N_636);
nand U987 (N_987,N_659,N_644);
nand U988 (N_988,N_638,N_664);
or U989 (N_989,N_797,N_666);
nand U990 (N_990,N_634,N_695);
and U991 (N_991,N_679,N_739);
nand U992 (N_992,N_757,N_603);
and U993 (N_993,N_683,N_795);
nand U994 (N_994,N_616,N_690);
or U995 (N_995,N_690,N_699);
and U996 (N_996,N_712,N_781);
or U997 (N_997,N_725,N_704);
nor U998 (N_998,N_686,N_775);
and U999 (N_999,N_785,N_666);
or U1000 (N_1000,N_951,N_984);
or U1001 (N_1001,N_834,N_953);
or U1002 (N_1002,N_904,N_988);
nand U1003 (N_1003,N_913,N_852);
nor U1004 (N_1004,N_908,N_932);
nor U1005 (N_1005,N_896,N_828);
and U1006 (N_1006,N_931,N_808);
nand U1007 (N_1007,N_959,N_999);
nand U1008 (N_1008,N_895,N_872);
nor U1009 (N_1009,N_880,N_843);
or U1010 (N_1010,N_874,N_830);
nor U1011 (N_1011,N_985,N_964);
or U1012 (N_1012,N_983,N_922);
nor U1013 (N_1013,N_822,N_975);
and U1014 (N_1014,N_831,N_813);
xor U1015 (N_1015,N_883,N_957);
nand U1016 (N_1016,N_936,N_812);
or U1017 (N_1017,N_920,N_942);
nand U1018 (N_1018,N_898,N_899);
nand U1019 (N_1019,N_995,N_979);
and U1020 (N_1020,N_844,N_960);
and U1021 (N_1021,N_864,N_832);
nor U1022 (N_1022,N_819,N_954);
nor U1023 (N_1023,N_937,N_980);
and U1024 (N_1024,N_890,N_863);
or U1025 (N_1025,N_862,N_800);
and U1026 (N_1026,N_962,N_933);
or U1027 (N_1027,N_835,N_892);
nor U1028 (N_1028,N_914,N_909);
nand U1029 (N_1029,N_935,N_943);
or U1030 (N_1030,N_807,N_925);
nor U1031 (N_1031,N_861,N_845);
and U1032 (N_1032,N_981,N_838);
or U1033 (N_1033,N_894,N_986);
nor U1034 (N_1034,N_804,N_850);
nor U1035 (N_1035,N_948,N_860);
and U1036 (N_1036,N_972,N_934);
nor U1037 (N_1037,N_967,N_833);
or U1038 (N_1038,N_857,N_961);
nand U1039 (N_1039,N_939,N_958);
or U1040 (N_1040,N_823,N_940);
nor U1041 (N_1041,N_809,N_841);
and U1042 (N_1042,N_884,N_888);
nand U1043 (N_1043,N_846,N_801);
or U1044 (N_1044,N_911,N_901);
nor U1045 (N_1045,N_916,N_849);
and U1046 (N_1046,N_919,N_867);
nand U1047 (N_1047,N_817,N_978);
or U1048 (N_1048,N_971,N_856);
and U1049 (N_1049,N_987,N_869);
and U1050 (N_1050,N_886,N_938);
or U1051 (N_1051,N_929,N_915);
nand U1052 (N_1052,N_930,N_875);
nor U1053 (N_1053,N_806,N_923);
or U1054 (N_1054,N_821,N_847);
or U1055 (N_1055,N_866,N_881);
or U1056 (N_1056,N_897,N_965);
or U1057 (N_1057,N_976,N_868);
nand U1058 (N_1058,N_945,N_855);
nor U1059 (N_1059,N_858,N_865);
nand U1060 (N_1060,N_926,N_891);
nor U1061 (N_1061,N_816,N_982);
nand U1062 (N_1062,N_815,N_949);
and U1063 (N_1063,N_992,N_842);
nor U1064 (N_1064,N_946,N_907);
and U1065 (N_1065,N_944,N_903);
nor U1066 (N_1066,N_956,N_826);
or U1067 (N_1067,N_973,N_970);
nor U1068 (N_1068,N_996,N_839);
or U1069 (N_1069,N_820,N_851);
and U1070 (N_1070,N_829,N_968);
nor U1071 (N_1071,N_917,N_977);
or U1072 (N_1072,N_989,N_877);
or U1073 (N_1073,N_836,N_811);
nor U1074 (N_1074,N_814,N_950);
or U1075 (N_1075,N_837,N_889);
nor U1076 (N_1076,N_924,N_941);
or U1077 (N_1077,N_993,N_893);
and U1078 (N_1078,N_991,N_998);
and U1079 (N_1079,N_974,N_928);
or U1080 (N_1080,N_871,N_947);
or U1081 (N_1081,N_969,N_882);
nand U1082 (N_1082,N_966,N_879);
nor U1083 (N_1083,N_885,N_905);
nor U1084 (N_1084,N_902,N_918);
and U1085 (N_1085,N_848,N_818);
nor U1086 (N_1086,N_853,N_873);
nand U1087 (N_1087,N_825,N_955);
or U1088 (N_1088,N_810,N_910);
and U1089 (N_1089,N_878,N_827);
or U1090 (N_1090,N_870,N_990);
nand U1091 (N_1091,N_824,N_921);
and U1092 (N_1092,N_840,N_876);
nor U1093 (N_1093,N_802,N_859);
nor U1094 (N_1094,N_906,N_912);
and U1095 (N_1095,N_952,N_805);
or U1096 (N_1096,N_803,N_854);
nand U1097 (N_1097,N_994,N_927);
or U1098 (N_1098,N_900,N_887);
nand U1099 (N_1099,N_963,N_997);
or U1100 (N_1100,N_887,N_919);
and U1101 (N_1101,N_908,N_895);
nand U1102 (N_1102,N_816,N_895);
nand U1103 (N_1103,N_861,N_848);
and U1104 (N_1104,N_938,N_902);
nor U1105 (N_1105,N_897,N_933);
and U1106 (N_1106,N_969,N_989);
nor U1107 (N_1107,N_895,N_959);
nand U1108 (N_1108,N_921,N_904);
nor U1109 (N_1109,N_917,N_981);
and U1110 (N_1110,N_845,N_972);
nand U1111 (N_1111,N_931,N_971);
or U1112 (N_1112,N_888,N_881);
nor U1113 (N_1113,N_895,N_975);
nand U1114 (N_1114,N_950,N_830);
and U1115 (N_1115,N_937,N_901);
nor U1116 (N_1116,N_986,N_828);
nand U1117 (N_1117,N_996,N_863);
nor U1118 (N_1118,N_910,N_914);
and U1119 (N_1119,N_820,N_819);
or U1120 (N_1120,N_826,N_960);
nor U1121 (N_1121,N_983,N_880);
and U1122 (N_1122,N_975,N_883);
or U1123 (N_1123,N_923,N_976);
nor U1124 (N_1124,N_881,N_944);
or U1125 (N_1125,N_879,N_860);
nand U1126 (N_1126,N_976,N_901);
and U1127 (N_1127,N_836,N_871);
nand U1128 (N_1128,N_860,N_813);
and U1129 (N_1129,N_802,N_842);
nand U1130 (N_1130,N_975,N_965);
and U1131 (N_1131,N_815,N_916);
and U1132 (N_1132,N_869,N_848);
or U1133 (N_1133,N_986,N_941);
and U1134 (N_1134,N_874,N_864);
and U1135 (N_1135,N_892,N_963);
or U1136 (N_1136,N_913,N_919);
nor U1137 (N_1137,N_913,N_876);
nor U1138 (N_1138,N_810,N_953);
nand U1139 (N_1139,N_894,N_991);
or U1140 (N_1140,N_937,N_803);
or U1141 (N_1141,N_939,N_957);
nor U1142 (N_1142,N_877,N_929);
nand U1143 (N_1143,N_859,N_900);
and U1144 (N_1144,N_949,N_960);
or U1145 (N_1145,N_822,N_982);
or U1146 (N_1146,N_895,N_859);
and U1147 (N_1147,N_988,N_977);
nor U1148 (N_1148,N_894,N_863);
nand U1149 (N_1149,N_810,N_854);
nor U1150 (N_1150,N_840,N_856);
or U1151 (N_1151,N_913,N_980);
nand U1152 (N_1152,N_935,N_854);
or U1153 (N_1153,N_823,N_972);
nor U1154 (N_1154,N_987,N_842);
and U1155 (N_1155,N_819,N_854);
and U1156 (N_1156,N_977,N_916);
and U1157 (N_1157,N_884,N_933);
nand U1158 (N_1158,N_910,N_949);
or U1159 (N_1159,N_881,N_883);
and U1160 (N_1160,N_993,N_880);
and U1161 (N_1161,N_952,N_809);
or U1162 (N_1162,N_822,N_945);
nand U1163 (N_1163,N_845,N_822);
and U1164 (N_1164,N_835,N_904);
or U1165 (N_1165,N_900,N_829);
and U1166 (N_1166,N_949,N_946);
and U1167 (N_1167,N_932,N_838);
nor U1168 (N_1168,N_816,N_979);
nor U1169 (N_1169,N_927,N_941);
or U1170 (N_1170,N_817,N_806);
nor U1171 (N_1171,N_807,N_826);
nand U1172 (N_1172,N_948,N_839);
and U1173 (N_1173,N_893,N_948);
or U1174 (N_1174,N_990,N_940);
or U1175 (N_1175,N_900,N_932);
or U1176 (N_1176,N_975,N_837);
or U1177 (N_1177,N_888,N_814);
or U1178 (N_1178,N_975,N_972);
nand U1179 (N_1179,N_812,N_815);
nand U1180 (N_1180,N_866,N_956);
or U1181 (N_1181,N_935,N_804);
nor U1182 (N_1182,N_860,N_833);
or U1183 (N_1183,N_921,N_967);
nor U1184 (N_1184,N_962,N_959);
nand U1185 (N_1185,N_892,N_916);
nor U1186 (N_1186,N_825,N_930);
nand U1187 (N_1187,N_882,N_898);
nor U1188 (N_1188,N_828,N_885);
or U1189 (N_1189,N_904,N_978);
or U1190 (N_1190,N_813,N_893);
or U1191 (N_1191,N_875,N_888);
nand U1192 (N_1192,N_817,N_937);
nand U1193 (N_1193,N_847,N_975);
or U1194 (N_1194,N_879,N_994);
nor U1195 (N_1195,N_911,N_910);
nor U1196 (N_1196,N_827,N_942);
and U1197 (N_1197,N_913,N_976);
and U1198 (N_1198,N_951,N_829);
nand U1199 (N_1199,N_875,N_898);
or U1200 (N_1200,N_1109,N_1148);
nand U1201 (N_1201,N_1147,N_1068);
nor U1202 (N_1202,N_1052,N_1045);
or U1203 (N_1203,N_1025,N_1119);
or U1204 (N_1204,N_1050,N_1092);
nand U1205 (N_1205,N_1062,N_1072);
nand U1206 (N_1206,N_1125,N_1124);
nand U1207 (N_1207,N_1195,N_1059);
nand U1208 (N_1208,N_1011,N_1107);
nor U1209 (N_1209,N_1091,N_1078);
nor U1210 (N_1210,N_1117,N_1085);
and U1211 (N_1211,N_1076,N_1069);
or U1212 (N_1212,N_1039,N_1056);
or U1213 (N_1213,N_1080,N_1028);
and U1214 (N_1214,N_1009,N_1186);
or U1215 (N_1215,N_1182,N_1035);
nor U1216 (N_1216,N_1007,N_1176);
and U1217 (N_1217,N_1089,N_1114);
nand U1218 (N_1218,N_1067,N_1196);
nor U1219 (N_1219,N_1074,N_1161);
or U1220 (N_1220,N_1152,N_1171);
nor U1221 (N_1221,N_1105,N_1136);
nand U1222 (N_1222,N_1033,N_1197);
and U1223 (N_1223,N_1058,N_1173);
and U1224 (N_1224,N_1086,N_1168);
nor U1225 (N_1225,N_1004,N_1179);
or U1226 (N_1226,N_1047,N_1008);
and U1227 (N_1227,N_1120,N_1097);
and U1228 (N_1228,N_1127,N_1166);
nand U1229 (N_1229,N_1108,N_1019);
nor U1230 (N_1230,N_1165,N_1135);
and U1231 (N_1231,N_1010,N_1103);
nand U1232 (N_1232,N_1126,N_1040);
or U1233 (N_1233,N_1192,N_1174);
or U1234 (N_1234,N_1156,N_1121);
or U1235 (N_1235,N_1157,N_1150);
nand U1236 (N_1236,N_1030,N_1053);
nor U1237 (N_1237,N_1049,N_1015);
or U1238 (N_1238,N_1187,N_1163);
or U1239 (N_1239,N_1073,N_1083);
nand U1240 (N_1240,N_1042,N_1075);
nand U1241 (N_1241,N_1041,N_1101);
nand U1242 (N_1242,N_1034,N_1063);
or U1243 (N_1243,N_1038,N_1118);
nor U1244 (N_1244,N_1128,N_1199);
and U1245 (N_1245,N_1137,N_1031);
nand U1246 (N_1246,N_1082,N_1023);
or U1247 (N_1247,N_1016,N_1132);
nor U1248 (N_1248,N_1003,N_1081);
or U1249 (N_1249,N_1141,N_1088);
nor U1250 (N_1250,N_1175,N_1142);
nor U1251 (N_1251,N_1046,N_1145);
nand U1252 (N_1252,N_1032,N_1021);
nand U1253 (N_1253,N_1112,N_1066);
or U1254 (N_1254,N_1094,N_1198);
and U1255 (N_1255,N_1190,N_1194);
or U1256 (N_1256,N_1172,N_1129);
nand U1257 (N_1257,N_1185,N_1012);
or U1258 (N_1258,N_1160,N_1155);
and U1259 (N_1259,N_1110,N_1054);
and U1260 (N_1260,N_1122,N_1167);
or U1261 (N_1261,N_1143,N_1188);
and U1262 (N_1262,N_1006,N_1139);
nand U1263 (N_1263,N_1146,N_1154);
nand U1264 (N_1264,N_1099,N_1095);
and U1265 (N_1265,N_1077,N_1149);
nor U1266 (N_1266,N_1071,N_1113);
nor U1267 (N_1267,N_1180,N_1193);
nor U1268 (N_1268,N_1014,N_1106);
and U1269 (N_1269,N_1177,N_1115);
nand U1270 (N_1270,N_1064,N_1090);
xnor U1271 (N_1271,N_1140,N_1051);
nand U1272 (N_1272,N_1153,N_1151);
nor U1273 (N_1273,N_1133,N_1098);
or U1274 (N_1274,N_1065,N_1018);
and U1275 (N_1275,N_1104,N_1060);
and U1276 (N_1276,N_1183,N_1070);
nor U1277 (N_1277,N_1102,N_1024);
and U1278 (N_1278,N_1189,N_1043);
or U1279 (N_1279,N_1178,N_1134);
nor U1280 (N_1280,N_1164,N_1191);
nor U1281 (N_1281,N_1144,N_1169);
nor U1282 (N_1282,N_1017,N_1159);
nor U1283 (N_1283,N_1184,N_1044);
xnor U1284 (N_1284,N_1027,N_1048);
or U1285 (N_1285,N_1061,N_1037);
nor U1286 (N_1286,N_1093,N_1100);
or U1287 (N_1287,N_1162,N_1079);
nor U1288 (N_1288,N_1000,N_1036);
nor U1289 (N_1289,N_1029,N_1020);
nor U1290 (N_1290,N_1096,N_1001);
nor U1291 (N_1291,N_1022,N_1130);
nor U1292 (N_1292,N_1158,N_1057);
xor U1293 (N_1293,N_1002,N_1111);
and U1294 (N_1294,N_1026,N_1013);
nor U1295 (N_1295,N_1138,N_1170);
nor U1296 (N_1296,N_1181,N_1084);
nand U1297 (N_1297,N_1116,N_1123);
nand U1298 (N_1298,N_1131,N_1055);
nand U1299 (N_1299,N_1005,N_1087);
nor U1300 (N_1300,N_1092,N_1072);
nand U1301 (N_1301,N_1199,N_1183);
and U1302 (N_1302,N_1145,N_1181);
and U1303 (N_1303,N_1014,N_1078);
or U1304 (N_1304,N_1073,N_1020);
or U1305 (N_1305,N_1108,N_1045);
or U1306 (N_1306,N_1050,N_1012);
or U1307 (N_1307,N_1035,N_1101);
and U1308 (N_1308,N_1100,N_1033);
and U1309 (N_1309,N_1060,N_1078);
or U1310 (N_1310,N_1064,N_1143);
and U1311 (N_1311,N_1056,N_1188);
nand U1312 (N_1312,N_1186,N_1185);
or U1313 (N_1313,N_1092,N_1035);
nand U1314 (N_1314,N_1112,N_1120);
nand U1315 (N_1315,N_1050,N_1138);
or U1316 (N_1316,N_1016,N_1041);
nor U1317 (N_1317,N_1026,N_1006);
nand U1318 (N_1318,N_1048,N_1003);
nor U1319 (N_1319,N_1191,N_1110);
and U1320 (N_1320,N_1033,N_1166);
nand U1321 (N_1321,N_1083,N_1165);
nor U1322 (N_1322,N_1067,N_1074);
nor U1323 (N_1323,N_1026,N_1161);
or U1324 (N_1324,N_1180,N_1058);
xor U1325 (N_1325,N_1116,N_1120);
nand U1326 (N_1326,N_1073,N_1131);
or U1327 (N_1327,N_1024,N_1188);
nor U1328 (N_1328,N_1046,N_1070);
nand U1329 (N_1329,N_1035,N_1132);
or U1330 (N_1330,N_1196,N_1115);
and U1331 (N_1331,N_1177,N_1057);
or U1332 (N_1332,N_1017,N_1119);
nor U1333 (N_1333,N_1090,N_1078);
or U1334 (N_1334,N_1114,N_1017);
and U1335 (N_1335,N_1062,N_1046);
nor U1336 (N_1336,N_1001,N_1080);
nand U1337 (N_1337,N_1029,N_1014);
nor U1338 (N_1338,N_1105,N_1114);
nor U1339 (N_1339,N_1060,N_1107);
or U1340 (N_1340,N_1130,N_1120);
nand U1341 (N_1341,N_1193,N_1045);
nor U1342 (N_1342,N_1149,N_1012);
and U1343 (N_1343,N_1119,N_1171);
and U1344 (N_1344,N_1134,N_1072);
nand U1345 (N_1345,N_1031,N_1013);
and U1346 (N_1346,N_1080,N_1189);
and U1347 (N_1347,N_1120,N_1188);
or U1348 (N_1348,N_1047,N_1146);
and U1349 (N_1349,N_1004,N_1100);
and U1350 (N_1350,N_1173,N_1190);
nor U1351 (N_1351,N_1115,N_1188);
or U1352 (N_1352,N_1140,N_1162);
and U1353 (N_1353,N_1132,N_1099);
nor U1354 (N_1354,N_1173,N_1035);
or U1355 (N_1355,N_1072,N_1067);
nor U1356 (N_1356,N_1069,N_1071);
and U1357 (N_1357,N_1178,N_1127);
nand U1358 (N_1358,N_1110,N_1160);
and U1359 (N_1359,N_1008,N_1033);
and U1360 (N_1360,N_1093,N_1179);
nand U1361 (N_1361,N_1176,N_1092);
and U1362 (N_1362,N_1084,N_1045);
nor U1363 (N_1363,N_1031,N_1166);
nor U1364 (N_1364,N_1020,N_1143);
and U1365 (N_1365,N_1064,N_1194);
and U1366 (N_1366,N_1142,N_1114);
nor U1367 (N_1367,N_1183,N_1095);
nand U1368 (N_1368,N_1025,N_1137);
or U1369 (N_1369,N_1182,N_1193);
nand U1370 (N_1370,N_1129,N_1169);
nor U1371 (N_1371,N_1101,N_1069);
or U1372 (N_1372,N_1184,N_1006);
xnor U1373 (N_1373,N_1022,N_1153);
nand U1374 (N_1374,N_1013,N_1051);
or U1375 (N_1375,N_1060,N_1054);
or U1376 (N_1376,N_1159,N_1038);
or U1377 (N_1377,N_1045,N_1146);
nand U1378 (N_1378,N_1070,N_1186);
nand U1379 (N_1379,N_1079,N_1093);
or U1380 (N_1380,N_1163,N_1010);
nor U1381 (N_1381,N_1076,N_1039);
nor U1382 (N_1382,N_1095,N_1100);
nor U1383 (N_1383,N_1151,N_1184);
nand U1384 (N_1384,N_1195,N_1199);
and U1385 (N_1385,N_1110,N_1192);
nor U1386 (N_1386,N_1082,N_1128);
nand U1387 (N_1387,N_1178,N_1007);
nor U1388 (N_1388,N_1095,N_1014);
or U1389 (N_1389,N_1120,N_1152);
nor U1390 (N_1390,N_1162,N_1043);
nor U1391 (N_1391,N_1007,N_1107);
nor U1392 (N_1392,N_1069,N_1051);
or U1393 (N_1393,N_1158,N_1046);
and U1394 (N_1394,N_1111,N_1055);
or U1395 (N_1395,N_1181,N_1073);
nand U1396 (N_1396,N_1080,N_1126);
or U1397 (N_1397,N_1167,N_1113);
nand U1398 (N_1398,N_1166,N_1172);
nand U1399 (N_1399,N_1066,N_1056);
nor U1400 (N_1400,N_1339,N_1225);
and U1401 (N_1401,N_1290,N_1231);
and U1402 (N_1402,N_1357,N_1346);
or U1403 (N_1403,N_1350,N_1232);
nand U1404 (N_1404,N_1252,N_1372);
nand U1405 (N_1405,N_1257,N_1288);
and U1406 (N_1406,N_1247,N_1293);
or U1407 (N_1407,N_1296,N_1300);
nor U1408 (N_1408,N_1388,N_1279);
nor U1409 (N_1409,N_1351,N_1284);
nor U1410 (N_1410,N_1345,N_1343);
and U1411 (N_1411,N_1266,N_1303);
or U1412 (N_1412,N_1223,N_1393);
or U1413 (N_1413,N_1299,N_1370);
nor U1414 (N_1414,N_1208,N_1368);
and U1415 (N_1415,N_1387,N_1255);
and U1416 (N_1416,N_1272,N_1265);
and U1417 (N_1417,N_1276,N_1254);
nor U1418 (N_1418,N_1383,N_1287);
nor U1419 (N_1419,N_1360,N_1399);
and U1420 (N_1420,N_1201,N_1329);
or U1421 (N_1421,N_1253,N_1369);
or U1422 (N_1422,N_1327,N_1356);
or U1423 (N_1423,N_1309,N_1242);
nand U1424 (N_1424,N_1269,N_1262);
and U1425 (N_1425,N_1301,N_1233);
and U1426 (N_1426,N_1245,N_1306);
and U1427 (N_1427,N_1317,N_1352);
nand U1428 (N_1428,N_1209,N_1365);
nand U1429 (N_1429,N_1324,N_1263);
or U1430 (N_1430,N_1358,N_1398);
nand U1431 (N_1431,N_1313,N_1271);
and U1432 (N_1432,N_1335,N_1326);
nor U1433 (N_1433,N_1280,N_1302);
and U1434 (N_1434,N_1328,N_1246);
nand U1435 (N_1435,N_1294,N_1385);
or U1436 (N_1436,N_1334,N_1361);
nor U1437 (N_1437,N_1212,N_1367);
or U1438 (N_1438,N_1362,N_1314);
and U1439 (N_1439,N_1282,N_1218);
nor U1440 (N_1440,N_1392,N_1376);
nor U1441 (N_1441,N_1251,N_1318);
nand U1442 (N_1442,N_1250,N_1204);
nor U1443 (N_1443,N_1386,N_1321);
nor U1444 (N_1444,N_1226,N_1205);
or U1445 (N_1445,N_1230,N_1366);
and U1446 (N_1446,N_1375,N_1289);
nand U1447 (N_1447,N_1203,N_1396);
nand U1448 (N_1448,N_1258,N_1364);
or U1449 (N_1449,N_1323,N_1273);
nor U1450 (N_1450,N_1286,N_1354);
and U1451 (N_1451,N_1240,N_1241);
and U1452 (N_1452,N_1312,N_1373);
nor U1453 (N_1453,N_1347,N_1261);
nor U1454 (N_1454,N_1344,N_1381);
nand U1455 (N_1455,N_1297,N_1374);
nand U1456 (N_1456,N_1342,N_1363);
and U1457 (N_1457,N_1292,N_1237);
nor U1458 (N_1458,N_1319,N_1234);
or U1459 (N_1459,N_1395,N_1210);
nand U1460 (N_1460,N_1268,N_1308);
nand U1461 (N_1461,N_1349,N_1267);
or U1462 (N_1462,N_1213,N_1338);
or U1463 (N_1463,N_1331,N_1207);
nand U1464 (N_1464,N_1382,N_1310);
and U1465 (N_1465,N_1325,N_1238);
nand U1466 (N_1466,N_1371,N_1236);
and U1467 (N_1467,N_1315,N_1394);
nor U1468 (N_1468,N_1391,N_1216);
or U1469 (N_1469,N_1380,N_1304);
nand U1470 (N_1470,N_1384,N_1320);
or U1471 (N_1471,N_1222,N_1311);
and U1472 (N_1472,N_1316,N_1219);
or U1473 (N_1473,N_1211,N_1259);
nand U1474 (N_1474,N_1291,N_1277);
or U1475 (N_1475,N_1348,N_1217);
and U1476 (N_1476,N_1378,N_1305);
nor U1477 (N_1477,N_1341,N_1377);
nor U1478 (N_1478,N_1248,N_1220);
xor U1479 (N_1479,N_1336,N_1285);
and U1480 (N_1480,N_1227,N_1275);
or U1481 (N_1481,N_1397,N_1379);
or U1482 (N_1482,N_1260,N_1243);
nand U1483 (N_1483,N_1389,N_1224);
nor U1484 (N_1484,N_1206,N_1249);
nor U1485 (N_1485,N_1353,N_1264);
nor U1486 (N_1486,N_1283,N_1215);
or U1487 (N_1487,N_1244,N_1281);
and U1488 (N_1488,N_1359,N_1228);
and U1489 (N_1489,N_1333,N_1200);
nor U1490 (N_1490,N_1330,N_1322);
nor U1491 (N_1491,N_1298,N_1202);
and U1492 (N_1492,N_1214,N_1337);
nand U1493 (N_1493,N_1355,N_1278);
or U1494 (N_1494,N_1390,N_1256);
and U1495 (N_1495,N_1295,N_1307);
or U1496 (N_1496,N_1270,N_1340);
or U1497 (N_1497,N_1332,N_1274);
nand U1498 (N_1498,N_1235,N_1239);
or U1499 (N_1499,N_1221,N_1229);
nor U1500 (N_1500,N_1260,N_1272);
nor U1501 (N_1501,N_1325,N_1279);
and U1502 (N_1502,N_1247,N_1254);
or U1503 (N_1503,N_1270,N_1230);
nand U1504 (N_1504,N_1254,N_1242);
xor U1505 (N_1505,N_1362,N_1356);
or U1506 (N_1506,N_1329,N_1234);
nor U1507 (N_1507,N_1249,N_1272);
and U1508 (N_1508,N_1334,N_1339);
nand U1509 (N_1509,N_1246,N_1218);
and U1510 (N_1510,N_1318,N_1277);
or U1511 (N_1511,N_1332,N_1292);
nor U1512 (N_1512,N_1217,N_1323);
nor U1513 (N_1513,N_1270,N_1399);
nor U1514 (N_1514,N_1243,N_1212);
and U1515 (N_1515,N_1220,N_1339);
nor U1516 (N_1516,N_1338,N_1273);
nand U1517 (N_1517,N_1390,N_1215);
nand U1518 (N_1518,N_1241,N_1271);
or U1519 (N_1519,N_1353,N_1206);
nand U1520 (N_1520,N_1319,N_1312);
or U1521 (N_1521,N_1394,N_1225);
and U1522 (N_1522,N_1380,N_1226);
nor U1523 (N_1523,N_1263,N_1212);
nor U1524 (N_1524,N_1262,N_1294);
nand U1525 (N_1525,N_1299,N_1293);
and U1526 (N_1526,N_1354,N_1281);
nand U1527 (N_1527,N_1222,N_1271);
nor U1528 (N_1528,N_1368,N_1275);
or U1529 (N_1529,N_1267,N_1276);
or U1530 (N_1530,N_1297,N_1342);
or U1531 (N_1531,N_1377,N_1217);
and U1532 (N_1532,N_1273,N_1203);
and U1533 (N_1533,N_1283,N_1204);
or U1534 (N_1534,N_1222,N_1338);
or U1535 (N_1535,N_1317,N_1341);
and U1536 (N_1536,N_1357,N_1275);
and U1537 (N_1537,N_1238,N_1291);
xor U1538 (N_1538,N_1252,N_1319);
or U1539 (N_1539,N_1376,N_1292);
or U1540 (N_1540,N_1239,N_1384);
or U1541 (N_1541,N_1299,N_1290);
nor U1542 (N_1542,N_1389,N_1353);
nand U1543 (N_1543,N_1379,N_1374);
nor U1544 (N_1544,N_1240,N_1242);
or U1545 (N_1545,N_1209,N_1307);
nand U1546 (N_1546,N_1308,N_1284);
nor U1547 (N_1547,N_1291,N_1339);
nor U1548 (N_1548,N_1314,N_1382);
or U1549 (N_1549,N_1318,N_1363);
nand U1550 (N_1550,N_1354,N_1370);
or U1551 (N_1551,N_1244,N_1369);
or U1552 (N_1552,N_1315,N_1377);
or U1553 (N_1553,N_1245,N_1246);
nand U1554 (N_1554,N_1258,N_1297);
or U1555 (N_1555,N_1205,N_1248);
nor U1556 (N_1556,N_1345,N_1283);
nand U1557 (N_1557,N_1216,N_1355);
and U1558 (N_1558,N_1346,N_1265);
or U1559 (N_1559,N_1224,N_1319);
nor U1560 (N_1560,N_1220,N_1381);
nand U1561 (N_1561,N_1287,N_1288);
nand U1562 (N_1562,N_1312,N_1395);
nand U1563 (N_1563,N_1322,N_1367);
nand U1564 (N_1564,N_1334,N_1390);
nor U1565 (N_1565,N_1236,N_1361);
nor U1566 (N_1566,N_1349,N_1299);
or U1567 (N_1567,N_1231,N_1205);
nand U1568 (N_1568,N_1374,N_1326);
or U1569 (N_1569,N_1279,N_1234);
nand U1570 (N_1570,N_1257,N_1379);
or U1571 (N_1571,N_1280,N_1274);
and U1572 (N_1572,N_1360,N_1321);
or U1573 (N_1573,N_1299,N_1223);
nand U1574 (N_1574,N_1312,N_1368);
nor U1575 (N_1575,N_1238,N_1288);
and U1576 (N_1576,N_1273,N_1354);
or U1577 (N_1577,N_1364,N_1293);
and U1578 (N_1578,N_1221,N_1206);
nand U1579 (N_1579,N_1360,N_1258);
nor U1580 (N_1580,N_1257,N_1226);
or U1581 (N_1581,N_1344,N_1391);
or U1582 (N_1582,N_1258,N_1230);
nand U1583 (N_1583,N_1266,N_1251);
and U1584 (N_1584,N_1312,N_1248);
nor U1585 (N_1585,N_1279,N_1217);
and U1586 (N_1586,N_1336,N_1315);
nand U1587 (N_1587,N_1381,N_1385);
nand U1588 (N_1588,N_1339,N_1357);
nand U1589 (N_1589,N_1258,N_1283);
nor U1590 (N_1590,N_1292,N_1374);
and U1591 (N_1591,N_1349,N_1245);
nor U1592 (N_1592,N_1226,N_1290);
nand U1593 (N_1593,N_1395,N_1225);
nand U1594 (N_1594,N_1215,N_1332);
nand U1595 (N_1595,N_1229,N_1254);
nand U1596 (N_1596,N_1308,N_1300);
nand U1597 (N_1597,N_1278,N_1328);
or U1598 (N_1598,N_1270,N_1302);
nor U1599 (N_1599,N_1232,N_1332);
nand U1600 (N_1600,N_1475,N_1564);
or U1601 (N_1601,N_1425,N_1516);
or U1602 (N_1602,N_1487,N_1498);
or U1603 (N_1603,N_1580,N_1560);
nand U1604 (N_1604,N_1426,N_1477);
nand U1605 (N_1605,N_1531,N_1540);
xnor U1606 (N_1606,N_1527,N_1595);
nand U1607 (N_1607,N_1405,N_1568);
or U1608 (N_1608,N_1440,N_1403);
and U1609 (N_1609,N_1465,N_1413);
nor U1610 (N_1610,N_1453,N_1534);
and U1611 (N_1611,N_1448,N_1515);
nor U1612 (N_1612,N_1429,N_1472);
nand U1613 (N_1613,N_1565,N_1419);
or U1614 (N_1614,N_1482,N_1467);
nor U1615 (N_1615,N_1486,N_1592);
and U1616 (N_1616,N_1507,N_1442);
or U1617 (N_1617,N_1599,N_1444);
and U1618 (N_1618,N_1538,N_1416);
and U1619 (N_1619,N_1420,N_1566);
or U1620 (N_1620,N_1578,N_1559);
or U1621 (N_1621,N_1509,N_1473);
nor U1622 (N_1622,N_1431,N_1589);
and U1623 (N_1623,N_1481,N_1490);
nor U1624 (N_1624,N_1411,N_1503);
nor U1625 (N_1625,N_1410,N_1581);
and U1626 (N_1626,N_1526,N_1464);
and U1627 (N_1627,N_1584,N_1548);
nor U1628 (N_1628,N_1458,N_1533);
or U1629 (N_1629,N_1468,N_1511);
nor U1630 (N_1630,N_1479,N_1459);
and U1631 (N_1631,N_1450,N_1446);
nor U1632 (N_1632,N_1434,N_1549);
nand U1633 (N_1633,N_1567,N_1579);
or U1634 (N_1634,N_1590,N_1497);
or U1635 (N_1635,N_1552,N_1517);
or U1636 (N_1636,N_1430,N_1588);
nor U1637 (N_1637,N_1528,N_1547);
and U1638 (N_1638,N_1572,N_1409);
nor U1639 (N_1639,N_1417,N_1408);
nand U1640 (N_1640,N_1596,N_1400);
and U1641 (N_1641,N_1502,N_1499);
and U1642 (N_1642,N_1447,N_1428);
or U1643 (N_1643,N_1582,N_1491);
nand U1644 (N_1644,N_1525,N_1587);
nor U1645 (N_1645,N_1529,N_1523);
nand U1646 (N_1646,N_1461,N_1501);
or U1647 (N_1647,N_1493,N_1539);
and U1648 (N_1648,N_1519,N_1577);
and U1649 (N_1649,N_1575,N_1557);
or U1650 (N_1650,N_1573,N_1508);
xnor U1651 (N_1651,N_1551,N_1506);
nand U1652 (N_1652,N_1488,N_1483);
nand U1653 (N_1653,N_1570,N_1471);
or U1654 (N_1654,N_1569,N_1406);
and U1655 (N_1655,N_1550,N_1495);
and U1656 (N_1656,N_1574,N_1441);
or U1657 (N_1657,N_1522,N_1598);
nor U1658 (N_1658,N_1422,N_1455);
nor U1659 (N_1659,N_1474,N_1423);
and U1660 (N_1660,N_1583,N_1591);
nor U1661 (N_1661,N_1556,N_1470);
nor U1662 (N_1662,N_1546,N_1407);
or U1663 (N_1663,N_1433,N_1460);
nand U1664 (N_1664,N_1521,N_1484);
nor U1665 (N_1665,N_1542,N_1415);
and U1666 (N_1666,N_1586,N_1432);
or U1667 (N_1667,N_1489,N_1597);
and U1668 (N_1668,N_1510,N_1402);
and U1669 (N_1669,N_1424,N_1585);
and U1670 (N_1670,N_1480,N_1494);
or U1671 (N_1671,N_1541,N_1537);
nand U1672 (N_1672,N_1454,N_1437);
or U1673 (N_1673,N_1593,N_1562);
or U1674 (N_1674,N_1443,N_1449);
nand U1675 (N_1675,N_1553,N_1427);
and U1676 (N_1676,N_1496,N_1576);
or U1677 (N_1677,N_1401,N_1438);
nor U1678 (N_1678,N_1543,N_1451);
nand U1679 (N_1679,N_1514,N_1535);
or U1680 (N_1680,N_1445,N_1421);
nor U1681 (N_1681,N_1476,N_1457);
nor U1682 (N_1682,N_1513,N_1561);
and U1683 (N_1683,N_1594,N_1463);
nand U1684 (N_1684,N_1545,N_1558);
or U1685 (N_1685,N_1555,N_1518);
nand U1686 (N_1686,N_1456,N_1436);
and U1687 (N_1687,N_1466,N_1512);
and U1688 (N_1688,N_1469,N_1418);
nand U1689 (N_1689,N_1544,N_1485);
and U1690 (N_1690,N_1504,N_1462);
and U1691 (N_1691,N_1404,N_1530);
or U1692 (N_1692,N_1520,N_1554);
nand U1693 (N_1693,N_1492,N_1524);
and U1694 (N_1694,N_1452,N_1414);
or U1695 (N_1695,N_1478,N_1563);
nor U1696 (N_1696,N_1435,N_1571);
nand U1697 (N_1697,N_1536,N_1500);
or U1698 (N_1698,N_1532,N_1439);
or U1699 (N_1699,N_1505,N_1412);
nand U1700 (N_1700,N_1577,N_1576);
or U1701 (N_1701,N_1515,N_1568);
nor U1702 (N_1702,N_1505,N_1482);
and U1703 (N_1703,N_1561,N_1466);
or U1704 (N_1704,N_1584,N_1405);
or U1705 (N_1705,N_1555,N_1560);
nor U1706 (N_1706,N_1411,N_1489);
nor U1707 (N_1707,N_1513,N_1568);
and U1708 (N_1708,N_1567,N_1590);
nand U1709 (N_1709,N_1577,N_1424);
nor U1710 (N_1710,N_1438,N_1508);
nor U1711 (N_1711,N_1482,N_1496);
nand U1712 (N_1712,N_1539,N_1583);
and U1713 (N_1713,N_1485,N_1419);
or U1714 (N_1714,N_1555,N_1474);
nand U1715 (N_1715,N_1590,N_1471);
and U1716 (N_1716,N_1515,N_1502);
nand U1717 (N_1717,N_1475,N_1599);
and U1718 (N_1718,N_1463,N_1434);
nor U1719 (N_1719,N_1569,N_1405);
and U1720 (N_1720,N_1437,N_1408);
or U1721 (N_1721,N_1458,N_1576);
and U1722 (N_1722,N_1414,N_1561);
and U1723 (N_1723,N_1407,N_1459);
and U1724 (N_1724,N_1596,N_1408);
nand U1725 (N_1725,N_1589,N_1521);
nand U1726 (N_1726,N_1582,N_1488);
nand U1727 (N_1727,N_1447,N_1544);
nor U1728 (N_1728,N_1451,N_1422);
nor U1729 (N_1729,N_1565,N_1414);
or U1730 (N_1730,N_1474,N_1447);
nor U1731 (N_1731,N_1494,N_1508);
and U1732 (N_1732,N_1583,N_1404);
and U1733 (N_1733,N_1483,N_1441);
and U1734 (N_1734,N_1429,N_1425);
nand U1735 (N_1735,N_1405,N_1597);
nand U1736 (N_1736,N_1513,N_1424);
and U1737 (N_1737,N_1524,N_1473);
and U1738 (N_1738,N_1558,N_1400);
nor U1739 (N_1739,N_1505,N_1478);
or U1740 (N_1740,N_1536,N_1534);
nand U1741 (N_1741,N_1504,N_1465);
and U1742 (N_1742,N_1571,N_1554);
and U1743 (N_1743,N_1580,N_1415);
or U1744 (N_1744,N_1401,N_1472);
and U1745 (N_1745,N_1421,N_1548);
nor U1746 (N_1746,N_1431,N_1447);
nor U1747 (N_1747,N_1471,N_1544);
and U1748 (N_1748,N_1402,N_1427);
nor U1749 (N_1749,N_1599,N_1443);
nand U1750 (N_1750,N_1467,N_1479);
nor U1751 (N_1751,N_1543,N_1578);
and U1752 (N_1752,N_1466,N_1463);
or U1753 (N_1753,N_1525,N_1572);
and U1754 (N_1754,N_1574,N_1567);
or U1755 (N_1755,N_1489,N_1417);
and U1756 (N_1756,N_1461,N_1443);
nand U1757 (N_1757,N_1453,N_1556);
and U1758 (N_1758,N_1414,N_1482);
nand U1759 (N_1759,N_1516,N_1496);
and U1760 (N_1760,N_1584,N_1469);
or U1761 (N_1761,N_1535,N_1536);
nand U1762 (N_1762,N_1416,N_1567);
or U1763 (N_1763,N_1403,N_1528);
or U1764 (N_1764,N_1470,N_1516);
and U1765 (N_1765,N_1467,N_1534);
and U1766 (N_1766,N_1490,N_1542);
or U1767 (N_1767,N_1586,N_1520);
and U1768 (N_1768,N_1445,N_1593);
or U1769 (N_1769,N_1446,N_1431);
and U1770 (N_1770,N_1540,N_1435);
nor U1771 (N_1771,N_1433,N_1411);
and U1772 (N_1772,N_1502,N_1510);
nand U1773 (N_1773,N_1448,N_1575);
nor U1774 (N_1774,N_1509,N_1522);
nand U1775 (N_1775,N_1436,N_1475);
or U1776 (N_1776,N_1594,N_1497);
nand U1777 (N_1777,N_1585,N_1599);
and U1778 (N_1778,N_1470,N_1404);
and U1779 (N_1779,N_1587,N_1570);
nor U1780 (N_1780,N_1455,N_1467);
or U1781 (N_1781,N_1403,N_1511);
nor U1782 (N_1782,N_1479,N_1424);
nor U1783 (N_1783,N_1496,N_1530);
or U1784 (N_1784,N_1588,N_1472);
and U1785 (N_1785,N_1477,N_1497);
or U1786 (N_1786,N_1566,N_1486);
and U1787 (N_1787,N_1418,N_1485);
nor U1788 (N_1788,N_1539,N_1451);
or U1789 (N_1789,N_1453,N_1582);
or U1790 (N_1790,N_1438,N_1557);
nor U1791 (N_1791,N_1531,N_1433);
nor U1792 (N_1792,N_1416,N_1529);
and U1793 (N_1793,N_1438,N_1534);
nand U1794 (N_1794,N_1534,N_1515);
nor U1795 (N_1795,N_1430,N_1577);
or U1796 (N_1796,N_1408,N_1409);
nor U1797 (N_1797,N_1569,N_1513);
nor U1798 (N_1798,N_1567,N_1422);
and U1799 (N_1799,N_1589,N_1523);
nand U1800 (N_1800,N_1604,N_1665);
or U1801 (N_1801,N_1749,N_1625);
and U1802 (N_1802,N_1636,N_1775);
or U1803 (N_1803,N_1700,N_1778);
or U1804 (N_1804,N_1677,N_1783);
xor U1805 (N_1805,N_1777,N_1764);
nor U1806 (N_1806,N_1765,N_1756);
and U1807 (N_1807,N_1717,N_1794);
nand U1808 (N_1808,N_1671,N_1757);
nor U1809 (N_1809,N_1759,N_1795);
nor U1810 (N_1810,N_1767,N_1686);
and U1811 (N_1811,N_1768,N_1748);
nand U1812 (N_1812,N_1718,N_1793);
nand U1813 (N_1813,N_1676,N_1620);
or U1814 (N_1814,N_1791,N_1739);
and U1815 (N_1815,N_1745,N_1702);
or U1816 (N_1816,N_1674,N_1743);
and U1817 (N_1817,N_1752,N_1753);
and U1818 (N_1818,N_1719,N_1699);
and U1819 (N_1819,N_1725,N_1648);
and U1820 (N_1820,N_1728,N_1784);
nor U1821 (N_1821,N_1798,N_1645);
and U1822 (N_1822,N_1796,N_1736);
nand U1823 (N_1823,N_1754,N_1704);
nor U1824 (N_1824,N_1723,N_1616);
and U1825 (N_1825,N_1644,N_1642);
and U1826 (N_1826,N_1619,N_1720);
and U1827 (N_1827,N_1773,N_1659);
nor U1828 (N_1828,N_1682,N_1713);
nand U1829 (N_1829,N_1782,N_1760);
and U1830 (N_1830,N_1761,N_1626);
and U1831 (N_1831,N_1670,N_1668);
and U1832 (N_1832,N_1660,N_1694);
or U1833 (N_1833,N_1672,N_1643);
or U1834 (N_1834,N_1751,N_1797);
and U1835 (N_1835,N_1612,N_1630);
nor U1836 (N_1836,N_1740,N_1780);
nor U1837 (N_1837,N_1657,N_1661);
nand U1838 (N_1838,N_1774,N_1770);
or U1839 (N_1839,N_1664,N_1662);
and U1840 (N_1840,N_1787,N_1709);
nor U1841 (N_1841,N_1680,N_1678);
and U1842 (N_1842,N_1701,N_1785);
and U1843 (N_1843,N_1714,N_1640);
nand U1844 (N_1844,N_1744,N_1687);
nand U1845 (N_1845,N_1675,N_1649);
nand U1846 (N_1846,N_1646,N_1666);
or U1847 (N_1847,N_1790,N_1639);
nand U1848 (N_1848,N_1673,N_1710);
nor U1849 (N_1849,N_1603,N_1741);
xnor U1850 (N_1850,N_1635,N_1746);
or U1851 (N_1851,N_1727,N_1608);
and U1852 (N_1852,N_1632,N_1618);
or U1853 (N_1853,N_1755,N_1658);
nor U1854 (N_1854,N_1669,N_1772);
nand U1855 (N_1855,N_1683,N_1623);
nand U1856 (N_1856,N_1734,N_1656);
nand U1857 (N_1857,N_1697,N_1724);
nor U1858 (N_1858,N_1690,N_1654);
and U1859 (N_1859,N_1695,N_1721);
nor U1860 (N_1860,N_1788,N_1651);
and U1861 (N_1861,N_1605,N_1733);
or U1862 (N_1862,N_1722,N_1663);
nand U1863 (N_1863,N_1617,N_1705);
and U1864 (N_1864,N_1730,N_1628);
nand U1865 (N_1865,N_1613,N_1779);
nor U1866 (N_1866,N_1602,N_1688);
and U1867 (N_1867,N_1691,N_1771);
nor U1868 (N_1868,N_1667,N_1711);
nand U1869 (N_1869,N_1615,N_1627);
nor U1870 (N_1870,N_1600,N_1735);
and U1871 (N_1871,N_1781,N_1776);
nand U1872 (N_1872,N_1799,N_1685);
or U1873 (N_1873,N_1689,N_1698);
xor U1874 (N_1874,N_1738,N_1763);
nand U1875 (N_1875,N_1637,N_1732);
or U1876 (N_1876,N_1696,N_1681);
or U1877 (N_1877,N_1715,N_1786);
nor U1878 (N_1878,N_1716,N_1633);
and U1879 (N_1879,N_1631,N_1647);
or U1880 (N_1880,N_1693,N_1789);
and U1881 (N_1881,N_1758,N_1726);
and U1882 (N_1882,N_1750,N_1729);
and U1883 (N_1883,N_1708,N_1731);
nand U1884 (N_1884,N_1679,N_1655);
and U1885 (N_1885,N_1706,N_1742);
and U1886 (N_1886,N_1792,N_1762);
nand U1887 (N_1887,N_1607,N_1638);
nand U1888 (N_1888,N_1606,N_1652);
and U1889 (N_1889,N_1611,N_1629);
nor U1890 (N_1890,N_1737,N_1622);
nand U1891 (N_1891,N_1692,N_1641);
or U1892 (N_1892,N_1609,N_1601);
nor U1893 (N_1893,N_1634,N_1684);
nand U1894 (N_1894,N_1769,N_1610);
nand U1895 (N_1895,N_1624,N_1707);
and U1896 (N_1896,N_1766,N_1703);
or U1897 (N_1897,N_1614,N_1650);
nor U1898 (N_1898,N_1712,N_1653);
and U1899 (N_1899,N_1747,N_1621);
and U1900 (N_1900,N_1716,N_1744);
or U1901 (N_1901,N_1640,N_1638);
and U1902 (N_1902,N_1794,N_1750);
nand U1903 (N_1903,N_1625,N_1650);
nor U1904 (N_1904,N_1795,N_1683);
nor U1905 (N_1905,N_1678,N_1617);
nor U1906 (N_1906,N_1658,N_1779);
and U1907 (N_1907,N_1659,N_1763);
nand U1908 (N_1908,N_1770,N_1781);
or U1909 (N_1909,N_1719,N_1779);
and U1910 (N_1910,N_1746,N_1725);
or U1911 (N_1911,N_1654,N_1612);
nor U1912 (N_1912,N_1774,N_1639);
nor U1913 (N_1913,N_1615,N_1749);
nand U1914 (N_1914,N_1761,N_1601);
nand U1915 (N_1915,N_1717,N_1687);
or U1916 (N_1916,N_1706,N_1755);
or U1917 (N_1917,N_1679,N_1779);
nor U1918 (N_1918,N_1786,N_1681);
and U1919 (N_1919,N_1658,N_1771);
and U1920 (N_1920,N_1630,N_1758);
and U1921 (N_1921,N_1712,N_1635);
nor U1922 (N_1922,N_1686,N_1710);
nand U1923 (N_1923,N_1635,N_1781);
and U1924 (N_1924,N_1774,N_1757);
or U1925 (N_1925,N_1769,N_1721);
nor U1926 (N_1926,N_1766,N_1601);
or U1927 (N_1927,N_1716,N_1657);
and U1928 (N_1928,N_1737,N_1643);
or U1929 (N_1929,N_1752,N_1743);
nand U1930 (N_1930,N_1696,N_1612);
or U1931 (N_1931,N_1669,N_1675);
nand U1932 (N_1932,N_1754,N_1765);
nor U1933 (N_1933,N_1640,N_1719);
nand U1934 (N_1934,N_1737,N_1785);
nor U1935 (N_1935,N_1667,N_1626);
or U1936 (N_1936,N_1607,N_1678);
nor U1937 (N_1937,N_1723,N_1774);
and U1938 (N_1938,N_1759,N_1619);
and U1939 (N_1939,N_1692,N_1635);
nand U1940 (N_1940,N_1753,N_1744);
nand U1941 (N_1941,N_1697,N_1653);
nor U1942 (N_1942,N_1639,N_1716);
or U1943 (N_1943,N_1601,N_1697);
xnor U1944 (N_1944,N_1653,N_1799);
nor U1945 (N_1945,N_1697,N_1620);
nor U1946 (N_1946,N_1760,N_1770);
nand U1947 (N_1947,N_1630,N_1723);
and U1948 (N_1948,N_1678,N_1695);
nor U1949 (N_1949,N_1669,N_1750);
or U1950 (N_1950,N_1667,N_1699);
or U1951 (N_1951,N_1673,N_1755);
nand U1952 (N_1952,N_1713,N_1712);
and U1953 (N_1953,N_1620,N_1763);
nand U1954 (N_1954,N_1602,N_1623);
nor U1955 (N_1955,N_1754,N_1697);
nand U1956 (N_1956,N_1617,N_1777);
or U1957 (N_1957,N_1756,N_1723);
or U1958 (N_1958,N_1798,N_1735);
or U1959 (N_1959,N_1768,N_1644);
and U1960 (N_1960,N_1767,N_1723);
or U1961 (N_1961,N_1731,N_1637);
nand U1962 (N_1962,N_1741,N_1792);
nor U1963 (N_1963,N_1661,N_1700);
nor U1964 (N_1964,N_1648,N_1667);
nor U1965 (N_1965,N_1614,N_1688);
or U1966 (N_1966,N_1716,N_1651);
nor U1967 (N_1967,N_1767,N_1666);
and U1968 (N_1968,N_1783,N_1799);
and U1969 (N_1969,N_1766,N_1626);
and U1970 (N_1970,N_1689,N_1785);
nor U1971 (N_1971,N_1601,N_1774);
or U1972 (N_1972,N_1756,N_1615);
and U1973 (N_1973,N_1677,N_1736);
nor U1974 (N_1974,N_1769,N_1637);
nor U1975 (N_1975,N_1669,N_1737);
or U1976 (N_1976,N_1662,N_1718);
or U1977 (N_1977,N_1729,N_1761);
nor U1978 (N_1978,N_1640,N_1626);
nor U1979 (N_1979,N_1630,N_1742);
and U1980 (N_1980,N_1711,N_1781);
nand U1981 (N_1981,N_1736,N_1623);
or U1982 (N_1982,N_1782,N_1614);
xor U1983 (N_1983,N_1688,N_1646);
nor U1984 (N_1984,N_1682,N_1670);
nor U1985 (N_1985,N_1691,N_1720);
and U1986 (N_1986,N_1771,N_1659);
and U1987 (N_1987,N_1694,N_1759);
nor U1988 (N_1988,N_1605,N_1752);
nand U1989 (N_1989,N_1623,N_1601);
nand U1990 (N_1990,N_1701,N_1783);
nand U1991 (N_1991,N_1725,N_1629);
and U1992 (N_1992,N_1724,N_1688);
nor U1993 (N_1993,N_1745,N_1750);
or U1994 (N_1994,N_1656,N_1761);
or U1995 (N_1995,N_1650,N_1686);
nor U1996 (N_1996,N_1675,N_1672);
or U1997 (N_1997,N_1616,N_1749);
nand U1998 (N_1998,N_1765,N_1646);
and U1999 (N_1999,N_1631,N_1677);
or U2000 (N_2000,N_1961,N_1938);
nand U2001 (N_2001,N_1811,N_1944);
or U2002 (N_2002,N_1925,N_1991);
or U2003 (N_2003,N_1955,N_1846);
nor U2004 (N_2004,N_1948,N_1974);
nor U2005 (N_2005,N_1899,N_1920);
nand U2006 (N_2006,N_1894,N_1966);
nor U2007 (N_2007,N_1877,N_1989);
nand U2008 (N_2008,N_1883,N_1875);
nand U2009 (N_2009,N_1819,N_1953);
or U2010 (N_2010,N_1994,N_1968);
nor U2011 (N_2011,N_1995,N_1900);
nor U2012 (N_2012,N_1977,N_1837);
nand U2013 (N_2013,N_1835,N_1911);
nand U2014 (N_2014,N_1874,N_1910);
nor U2015 (N_2015,N_1892,N_1993);
nand U2016 (N_2016,N_1949,N_1915);
and U2017 (N_2017,N_1902,N_1861);
and U2018 (N_2018,N_1978,N_1801);
nor U2019 (N_2019,N_1880,N_1836);
and U2020 (N_2020,N_1878,N_1828);
and U2021 (N_2021,N_1946,N_1913);
or U2022 (N_2022,N_1919,N_1873);
nand U2023 (N_2023,N_1807,N_1976);
nor U2024 (N_2024,N_1996,N_1983);
or U2025 (N_2025,N_1926,N_1981);
and U2026 (N_2026,N_1992,N_1936);
nor U2027 (N_2027,N_1849,N_1942);
nor U2028 (N_2028,N_1998,N_1973);
or U2029 (N_2029,N_1943,N_1839);
nor U2030 (N_2030,N_1945,N_1986);
nor U2031 (N_2031,N_1906,N_1962);
nand U2032 (N_2032,N_1890,N_1820);
nor U2033 (N_2033,N_1806,N_1823);
or U2034 (N_2034,N_1845,N_1941);
nor U2035 (N_2035,N_1927,N_1904);
nand U2036 (N_2036,N_1821,N_1912);
and U2037 (N_2037,N_1853,N_1847);
nor U2038 (N_2038,N_1803,N_1922);
or U2039 (N_2039,N_1959,N_1870);
and U2040 (N_2040,N_1869,N_1963);
nand U2041 (N_2041,N_1908,N_1997);
nand U2042 (N_2042,N_1832,N_1848);
nor U2043 (N_2043,N_1813,N_1972);
nor U2044 (N_2044,N_1805,N_1933);
nor U2045 (N_2045,N_1868,N_1950);
nor U2046 (N_2046,N_1979,N_1816);
and U2047 (N_2047,N_1897,N_1957);
or U2048 (N_2048,N_1982,N_1905);
or U2049 (N_2049,N_1939,N_1815);
nand U2050 (N_2050,N_1842,N_1951);
nand U2051 (N_2051,N_1872,N_1889);
xor U2052 (N_2052,N_1952,N_1929);
nor U2053 (N_2053,N_1924,N_1809);
nand U2054 (N_2054,N_1931,N_1812);
or U2055 (N_2055,N_1808,N_1887);
nand U2056 (N_2056,N_1826,N_1802);
or U2057 (N_2057,N_1830,N_1888);
nor U2058 (N_2058,N_1818,N_1916);
or U2059 (N_2059,N_1930,N_1884);
nor U2060 (N_2060,N_1918,N_1817);
or U2061 (N_2061,N_1990,N_1935);
and U2062 (N_2062,N_1917,N_1831);
nand U2063 (N_2063,N_1850,N_1804);
nor U2064 (N_2064,N_1999,N_1855);
nor U2065 (N_2065,N_1980,N_1984);
or U2066 (N_2066,N_1891,N_1840);
and U2067 (N_2067,N_1886,N_1825);
nor U2068 (N_2068,N_1829,N_1858);
nand U2069 (N_2069,N_1844,N_1985);
nor U2070 (N_2070,N_1987,N_1863);
or U2071 (N_2071,N_1859,N_1885);
nor U2072 (N_2072,N_1876,N_1909);
or U2073 (N_2073,N_1907,N_1882);
or U2074 (N_2074,N_1958,N_1865);
and U2075 (N_2075,N_1854,N_1970);
or U2076 (N_2076,N_1862,N_1810);
or U2077 (N_2077,N_1857,N_1967);
or U2078 (N_2078,N_1901,N_1834);
nor U2079 (N_2079,N_1903,N_1937);
and U2080 (N_2080,N_1833,N_1964);
and U2081 (N_2081,N_1954,N_1871);
nand U2082 (N_2082,N_1843,N_1928);
and U2083 (N_2083,N_1965,N_1860);
or U2084 (N_2084,N_1866,N_1914);
nor U2085 (N_2085,N_1881,N_1841);
or U2086 (N_2086,N_1940,N_1934);
nor U2087 (N_2087,N_1947,N_1814);
nand U2088 (N_2088,N_1969,N_1956);
and U2089 (N_2089,N_1822,N_1895);
or U2090 (N_2090,N_1856,N_1988);
or U2091 (N_2091,N_1898,N_1921);
and U2092 (N_2092,N_1893,N_1879);
nor U2093 (N_2093,N_1923,N_1827);
nand U2094 (N_2094,N_1867,N_1800);
nor U2095 (N_2095,N_1838,N_1896);
and U2096 (N_2096,N_1851,N_1971);
nor U2097 (N_2097,N_1824,N_1852);
or U2098 (N_2098,N_1932,N_1975);
or U2099 (N_2099,N_1864,N_1960);
or U2100 (N_2100,N_1924,N_1850);
or U2101 (N_2101,N_1997,N_1823);
nor U2102 (N_2102,N_1833,N_1992);
and U2103 (N_2103,N_1894,N_1982);
or U2104 (N_2104,N_1854,N_1932);
nand U2105 (N_2105,N_1966,N_1861);
nand U2106 (N_2106,N_1892,N_1879);
or U2107 (N_2107,N_1906,N_1831);
nand U2108 (N_2108,N_1868,N_1871);
nand U2109 (N_2109,N_1820,N_1972);
nand U2110 (N_2110,N_1809,N_1939);
and U2111 (N_2111,N_1958,N_1856);
nand U2112 (N_2112,N_1869,N_1968);
nand U2113 (N_2113,N_1938,N_1864);
or U2114 (N_2114,N_1904,N_1815);
or U2115 (N_2115,N_1887,N_1836);
nand U2116 (N_2116,N_1922,N_1898);
and U2117 (N_2117,N_1986,N_1836);
nand U2118 (N_2118,N_1975,N_1812);
nand U2119 (N_2119,N_1874,N_1827);
nor U2120 (N_2120,N_1938,N_1944);
nand U2121 (N_2121,N_1913,N_1947);
or U2122 (N_2122,N_1883,N_1839);
and U2123 (N_2123,N_1885,N_1984);
nand U2124 (N_2124,N_1848,N_1812);
nand U2125 (N_2125,N_1849,N_1839);
and U2126 (N_2126,N_1826,N_1843);
nand U2127 (N_2127,N_1968,N_1950);
or U2128 (N_2128,N_1902,N_1801);
and U2129 (N_2129,N_1801,N_1821);
nand U2130 (N_2130,N_1990,N_1861);
and U2131 (N_2131,N_1883,N_1807);
and U2132 (N_2132,N_1920,N_1985);
or U2133 (N_2133,N_1872,N_1824);
nor U2134 (N_2134,N_1805,N_1866);
nor U2135 (N_2135,N_1967,N_1914);
and U2136 (N_2136,N_1842,N_1901);
and U2137 (N_2137,N_1899,N_1834);
nor U2138 (N_2138,N_1897,N_1841);
or U2139 (N_2139,N_1976,N_1949);
nor U2140 (N_2140,N_1935,N_1807);
or U2141 (N_2141,N_1961,N_1951);
nand U2142 (N_2142,N_1874,N_1905);
nor U2143 (N_2143,N_1994,N_1960);
nor U2144 (N_2144,N_1870,N_1869);
nor U2145 (N_2145,N_1848,N_1857);
or U2146 (N_2146,N_1849,N_1937);
or U2147 (N_2147,N_1822,N_1818);
nand U2148 (N_2148,N_1802,N_1892);
and U2149 (N_2149,N_1811,N_1963);
nor U2150 (N_2150,N_1887,N_1958);
and U2151 (N_2151,N_1863,N_1973);
and U2152 (N_2152,N_1840,N_1981);
or U2153 (N_2153,N_1877,N_1802);
or U2154 (N_2154,N_1988,N_1847);
or U2155 (N_2155,N_1992,N_1975);
and U2156 (N_2156,N_1832,N_1808);
nor U2157 (N_2157,N_1974,N_1924);
and U2158 (N_2158,N_1993,N_1979);
or U2159 (N_2159,N_1807,N_1881);
nor U2160 (N_2160,N_1912,N_1818);
nand U2161 (N_2161,N_1994,N_1837);
or U2162 (N_2162,N_1904,N_1828);
nor U2163 (N_2163,N_1904,N_1873);
nand U2164 (N_2164,N_1834,N_1977);
nor U2165 (N_2165,N_1866,N_1840);
or U2166 (N_2166,N_1972,N_1816);
or U2167 (N_2167,N_1810,N_1815);
nor U2168 (N_2168,N_1807,N_1821);
nand U2169 (N_2169,N_1871,N_1996);
nor U2170 (N_2170,N_1916,N_1848);
and U2171 (N_2171,N_1995,N_1923);
nor U2172 (N_2172,N_1847,N_1871);
and U2173 (N_2173,N_1994,N_1985);
and U2174 (N_2174,N_1893,N_1894);
or U2175 (N_2175,N_1950,N_1955);
and U2176 (N_2176,N_1907,N_1967);
or U2177 (N_2177,N_1989,N_1963);
or U2178 (N_2178,N_1993,N_1835);
or U2179 (N_2179,N_1800,N_1910);
nor U2180 (N_2180,N_1840,N_1974);
nand U2181 (N_2181,N_1887,N_1949);
nor U2182 (N_2182,N_1939,N_1941);
nor U2183 (N_2183,N_1845,N_1989);
nor U2184 (N_2184,N_1968,N_1959);
nor U2185 (N_2185,N_1992,N_1942);
nand U2186 (N_2186,N_1938,N_1879);
or U2187 (N_2187,N_1972,N_1898);
nand U2188 (N_2188,N_1802,N_1932);
and U2189 (N_2189,N_1803,N_1914);
and U2190 (N_2190,N_1919,N_1962);
nand U2191 (N_2191,N_1810,N_1928);
or U2192 (N_2192,N_1880,N_1851);
or U2193 (N_2193,N_1850,N_1874);
nor U2194 (N_2194,N_1817,N_1806);
nand U2195 (N_2195,N_1842,N_1930);
and U2196 (N_2196,N_1881,N_1910);
nand U2197 (N_2197,N_1855,N_1810);
or U2198 (N_2198,N_1903,N_1985);
nand U2199 (N_2199,N_1957,N_1890);
and U2200 (N_2200,N_2008,N_2121);
nor U2201 (N_2201,N_2048,N_2004);
or U2202 (N_2202,N_2029,N_2170);
and U2203 (N_2203,N_2034,N_2118);
and U2204 (N_2204,N_2134,N_2058);
or U2205 (N_2205,N_2169,N_2087);
and U2206 (N_2206,N_2174,N_2076);
nand U2207 (N_2207,N_2083,N_2041);
and U2208 (N_2208,N_2192,N_2081);
nand U2209 (N_2209,N_2013,N_2086);
nor U2210 (N_2210,N_2062,N_2094);
xnor U2211 (N_2211,N_2042,N_2059);
or U2212 (N_2212,N_2054,N_2128);
nor U2213 (N_2213,N_2175,N_2142);
and U2214 (N_2214,N_2148,N_2088);
nand U2215 (N_2215,N_2178,N_2098);
or U2216 (N_2216,N_2166,N_2049);
nand U2217 (N_2217,N_2194,N_2114);
or U2218 (N_2218,N_2130,N_2187);
nand U2219 (N_2219,N_2043,N_2075);
and U2220 (N_2220,N_2039,N_2153);
nor U2221 (N_2221,N_2012,N_2154);
and U2222 (N_2222,N_2085,N_2031);
and U2223 (N_2223,N_2106,N_2109);
or U2224 (N_2224,N_2111,N_2033);
nor U2225 (N_2225,N_2028,N_2161);
nor U2226 (N_2226,N_2127,N_2159);
nor U2227 (N_2227,N_2019,N_2052);
and U2228 (N_2228,N_2030,N_2020);
nor U2229 (N_2229,N_2093,N_2167);
nand U2230 (N_2230,N_2023,N_2000);
nor U2231 (N_2231,N_2001,N_2018);
nor U2232 (N_2232,N_2158,N_2070);
nand U2233 (N_2233,N_2104,N_2003);
nand U2234 (N_2234,N_2191,N_2097);
nor U2235 (N_2235,N_2186,N_2196);
and U2236 (N_2236,N_2080,N_2151);
and U2237 (N_2237,N_2156,N_2010);
nand U2238 (N_2238,N_2091,N_2171);
nor U2239 (N_2239,N_2055,N_2068);
nor U2240 (N_2240,N_2040,N_2162);
xnor U2241 (N_2241,N_2135,N_2032);
or U2242 (N_2242,N_2071,N_2197);
nand U2243 (N_2243,N_2176,N_2037);
nor U2244 (N_2244,N_2146,N_2073);
and U2245 (N_2245,N_2172,N_2129);
and U2246 (N_2246,N_2108,N_2017);
nor U2247 (N_2247,N_2045,N_2066);
and U2248 (N_2248,N_2155,N_2082);
xnor U2249 (N_2249,N_2079,N_2163);
and U2250 (N_2250,N_2044,N_2089);
nand U2251 (N_2251,N_2160,N_2025);
or U2252 (N_2252,N_2057,N_2005);
nor U2253 (N_2253,N_2053,N_2189);
and U2254 (N_2254,N_2064,N_2188);
or U2255 (N_2255,N_2072,N_2113);
nand U2256 (N_2256,N_2078,N_2116);
nor U2257 (N_2257,N_2050,N_2047);
and U2258 (N_2258,N_2164,N_2105);
or U2259 (N_2259,N_2077,N_2133);
or U2260 (N_2260,N_2193,N_2063);
and U2261 (N_2261,N_2143,N_2179);
or U2262 (N_2262,N_2185,N_2056);
and U2263 (N_2263,N_2046,N_2141);
or U2264 (N_2264,N_2136,N_2024);
nand U2265 (N_2265,N_2096,N_2006);
nor U2266 (N_2266,N_2198,N_2107);
and U2267 (N_2267,N_2181,N_2157);
or U2268 (N_2268,N_2011,N_2124);
nand U2269 (N_2269,N_2182,N_2180);
nand U2270 (N_2270,N_2061,N_2123);
nand U2271 (N_2271,N_2195,N_2150);
or U2272 (N_2272,N_2126,N_2007);
or U2273 (N_2273,N_2103,N_2112);
and U2274 (N_2274,N_2021,N_2149);
nor U2275 (N_2275,N_2190,N_2092);
nor U2276 (N_2276,N_2110,N_2095);
or U2277 (N_2277,N_2102,N_2038);
or U2278 (N_2278,N_2117,N_2016);
or U2279 (N_2279,N_2132,N_2100);
and U2280 (N_2280,N_2184,N_2035);
nor U2281 (N_2281,N_2036,N_2060);
or U2282 (N_2282,N_2137,N_2065);
and U2283 (N_2283,N_2165,N_2122);
nor U2284 (N_2284,N_2119,N_2027);
and U2285 (N_2285,N_2139,N_2144);
and U2286 (N_2286,N_2140,N_2168);
nor U2287 (N_2287,N_2051,N_2084);
or U2288 (N_2288,N_2002,N_2090);
nand U2289 (N_2289,N_2120,N_2069);
and U2290 (N_2290,N_2026,N_2014);
or U2291 (N_2291,N_2199,N_2101);
nor U2292 (N_2292,N_2173,N_2138);
nand U2293 (N_2293,N_2147,N_2183);
nor U2294 (N_2294,N_2099,N_2015);
nor U2295 (N_2295,N_2125,N_2074);
or U2296 (N_2296,N_2009,N_2145);
and U2297 (N_2297,N_2022,N_2131);
or U2298 (N_2298,N_2152,N_2115);
and U2299 (N_2299,N_2177,N_2067);
and U2300 (N_2300,N_2140,N_2003);
nand U2301 (N_2301,N_2122,N_2116);
nor U2302 (N_2302,N_2086,N_2137);
nand U2303 (N_2303,N_2172,N_2188);
nor U2304 (N_2304,N_2068,N_2009);
nor U2305 (N_2305,N_2161,N_2085);
or U2306 (N_2306,N_2010,N_2024);
and U2307 (N_2307,N_2039,N_2047);
or U2308 (N_2308,N_2149,N_2120);
and U2309 (N_2309,N_2107,N_2125);
or U2310 (N_2310,N_2025,N_2114);
nand U2311 (N_2311,N_2145,N_2153);
nor U2312 (N_2312,N_2142,N_2161);
or U2313 (N_2313,N_2150,N_2154);
xor U2314 (N_2314,N_2137,N_2145);
and U2315 (N_2315,N_2005,N_2023);
and U2316 (N_2316,N_2168,N_2128);
or U2317 (N_2317,N_2151,N_2005);
and U2318 (N_2318,N_2032,N_2014);
and U2319 (N_2319,N_2040,N_2074);
and U2320 (N_2320,N_2009,N_2143);
nor U2321 (N_2321,N_2006,N_2122);
or U2322 (N_2322,N_2183,N_2177);
nand U2323 (N_2323,N_2140,N_2090);
nand U2324 (N_2324,N_2020,N_2194);
and U2325 (N_2325,N_2152,N_2098);
or U2326 (N_2326,N_2067,N_2099);
nor U2327 (N_2327,N_2099,N_2196);
nand U2328 (N_2328,N_2140,N_2137);
nor U2329 (N_2329,N_2064,N_2186);
and U2330 (N_2330,N_2156,N_2139);
nor U2331 (N_2331,N_2155,N_2143);
nor U2332 (N_2332,N_2071,N_2103);
and U2333 (N_2333,N_2112,N_2125);
nand U2334 (N_2334,N_2046,N_2087);
and U2335 (N_2335,N_2157,N_2035);
nand U2336 (N_2336,N_2106,N_2067);
nor U2337 (N_2337,N_2127,N_2111);
nand U2338 (N_2338,N_2091,N_2135);
nor U2339 (N_2339,N_2192,N_2163);
nand U2340 (N_2340,N_2131,N_2166);
nand U2341 (N_2341,N_2006,N_2054);
nor U2342 (N_2342,N_2061,N_2038);
and U2343 (N_2343,N_2027,N_2047);
or U2344 (N_2344,N_2087,N_2090);
nand U2345 (N_2345,N_2134,N_2194);
nor U2346 (N_2346,N_2049,N_2185);
nand U2347 (N_2347,N_2154,N_2134);
xnor U2348 (N_2348,N_2169,N_2105);
and U2349 (N_2349,N_2145,N_2120);
nor U2350 (N_2350,N_2150,N_2076);
or U2351 (N_2351,N_2168,N_2121);
nor U2352 (N_2352,N_2027,N_2111);
or U2353 (N_2353,N_2162,N_2025);
nand U2354 (N_2354,N_2035,N_2188);
nor U2355 (N_2355,N_2011,N_2163);
and U2356 (N_2356,N_2171,N_2097);
and U2357 (N_2357,N_2002,N_2067);
nand U2358 (N_2358,N_2085,N_2026);
nand U2359 (N_2359,N_2031,N_2101);
nor U2360 (N_2360,N_2018,N_2134);
and U2361 (N_2361,N_2118,N_2064);
or U2362 (N_2362,N_2135,N_2158);
and U2363 (N_2363,N_2158,N_2055);
nor U2364 (N_2364,N_2060,N_2147);
or U2365 (N_2365,N_2133,N_2024);
nand U2366 (N_2366,N_2199,N_2138);
nor U2367 (N_2367,N_2049,N_2148);
nand U2368 (N_2368,N_2102,N_2183);
or U2369 (N_2369,N_2009,N_2129);
or U2370 (N_2370,N_2077,N_2152);
xor U2371 (N_2371,N_2016,N_2094);
nor U2372 (N_2372,N_2113,N_2108);
and U2373 (N_2373,N_2113,N_2048);
or U2374 (N_2374,N_2083,N_2089);
and U2375 (N_2375,N_2198,N_2127);
nor U2376 (N_2376,N_2082,N_2197);
nor U2377 (N_2377,N_2031,N_2018);
nor U2378 (N_2378,N_2120,N_2076);
nand U2379 (N_2379,N_2027,N_2038);
and U2380 (N_2380,N_2168,N_2027);
nor U2381 (N_2381,N_2154,N_2077);
nand U2382 (N_2382,N_2020,N_2072);
nand U2383 (N_2383,N_2039,N_2052);
and U2384 (N_2384,N_2092,N_2106);
or U2385 (N_2385,N_2046,N_2026);
nor U2386 (N_2386,N_2015,N_2051);
nor U2387 (N_2387,N_2019,N_2107);
and U2388 (N_2388,N_2165,N_2053);
or U2389 (N_2389,N_2062,N_2193);
or U2390 (N_2390,N_2088,N_2187);
nor U2391 (N_2391,N_2024,N_2106);
or U2392 (N_2392,N_2007,N_2102);
nand U2393 (N_2393,N_2035,N_2121);
and U2394 (N_2394,N_2135,N_2094);
nand U2395 (N_2395,N_2158,N_2176);
or U2396 (N_2396,N_2118,N_2199);
or U2397 (N_2397,N_2192,N_2176);
xor U2398 (N_2398,N_2082,N_2050);
nand U2399 (N_2399,N_2157,N_2150);
or U2400 (N_2400,N_2386,N_2243);
nor U2401 (N_2401,N_2389,N_2373);
nor U2402 (N_2402,N_2315,N_2325);
or U2403 (N_2403,N_2328,N_2394);
nor U2404 (N_2404,N_2376,N_2237);
and U2405 (N_2405,N_2399,N_2344);
nor U2406 (N_2406,N_2253,N_2366);
or U2407 (N_2407,N_2278,N_2252);
and U2408 (N_2408,N_2365,N_2321);
and U2409 (N_2409,N_2244,N_2273);
and U2410 (N_2410,N_2268,N_2370);
nor U2411 (N_2411,N_2327,N_2326);
and U2412 (N_2412,N_2342,N_2357);
nand U2413 (N_2413,N_2387,N_2230);
and U2414 (N_2414,N_2350,N_2360);
or U2415 (N_2415,N_2287,N_2383);
or U2416 (N_2416,N_2332,N_2235);
nor U2417 (N_2417,N_2208,N_2228);
nor U2418 (N_2418,N_2364,N_2358);
nand U2419 (N_2419,N_2353,N_2356);
nand U2420 (N_2420,N_2222,N_2262);
or U2421 (N_2421,N_2207,N_2374);
and U2422 (N_2422,N_2294,N_2368);
nor U2423 (N_2423,N_2363,N_2379);
and U2424 (N_2424,N_2331,N_2265);
nor U2425 (N_2425,N_2362,N_2256);
nor U2426 (N_2426,N_2267,N_2302);
nand U2427 (N_2427,N_2220,N_2203);
or U2428 (N_2428,N_2313,N_2248);
nor U2429 (N_2429,N_2232,N_2254);
nor U2430 (N_2430,N_2334,N_2255);
or U2431 (N_2431,N_2247,N_2223);
or U2432 (N_2432,N_2311,N_2337);
or U2433 (N_2433,N_2291,N_2380);
or U2434 (N_2434,N_2233,N_2209);
or U2435 (N_2435,N_2216,N_2289);
or U2436 (N_2436,N_2296,N_2293);
nand U2437 (N_2437,N_2210,N_2234);
or U2438 (N_2438,N_2226,N_2347);
nand U2439 (N_2439,N_2245,N_2258);
or U2440 (N_2440,N_2242,N_2206);
nand U2441 (N_2441,N_2336,N_2390);
nor U2442 (N_2442,N_2283,N_2264);
nand U2443 (N_2443,N_2260,N_2246);
or U2444 (N_2444,N_2297,N_2241);
and U2445 (N_2445,N_2303,N_2304);
or U2446 (N_2446,N_2263,N_2318);
or U2447 (N_2447,N_2249,N_2316);
nor U2448 (N_2448,N_2295,N_2300);
or U2449 (N_2449,N_2384,N_2280);
nand U2450 (N_2450,N_2284,N_2352);
nand U2451 (N_2451,N_2346,N_2224);
nor U2452 (N_2452,N_2301,N_2231);
nor U2453 (N_2453,N_2261,N_2201);
nand U2454 (N_2454,N_2305,N_2345);
and U2455 (N_2455,N_2323,N_2277);
nand U2456 (N_2456,N_2269,N_2214);
nor U2457 (N_2457,N_2377,N_2212);
nor U2458 (N_2458,N_2349,N_2298);
nand U2459 (N_2459,N_2333,N_2211);
and U2460 (N_2460,N_2217,N_2392);
nor U2461 (N_2461,N_2398,N_2229);
nand U2462 (N_2462,N_2382,N_2202);
or U2463 (N_2463,N_2381,N_2391);
nor U2464 (N_2464,N_2314,N_2215);
nor U2465 (N_2465,N_2385,N_2348);
nor U2466 (N_2466,N_2341,N_2355);
or U2467 (N_2467,N_2361,N_2282);
and U2468 (N_2468,N_2250,N_2259);
and U2469 (N_2469,N_2388,N_2272);
or U2470 (N_2470,N_2274,N_2286);
and U2471 (N_2471,N_2317,N_2306);
nor U2472 (N_2472,N_2351,N_2319);
nor U2473 (N_2473,N_2307,N_2240);
and U2474 (N_2474,N_2219,N_2367);
nand U2475 (N_2475,N_2204,N_2335);
and U2476 (N_2476,N_2285,N_2270);
nand U2477 (N_2477,N_2218,N_2227);
and U2478 (N_2478,N_2396,N_2359);
nand U2479 (N_2479,N_2338,N_2292);
or U2480 (N_2480,N_2310,N_2257);
nor U2481 (N_2481,N_2375,N_2266);
nor U2482 (N_2482,N_2279,N_2309);
nor U2483 (N_2483,N_2308,N_2329);
or U2484 (N_2484,N_2200,N_2213);
or U2485 (N_2485,N_2397,N_2339);
or U2486 (N_2486,N_2312,N_2320);
nand U2487 (N_2487,N_2221,N_2330);
nor U2488 (N_2488,N_2340,N_2236);
nand U2489 (N_2489,N_2225,N_2395);
nor U2490 (N_2490,N_2281,N_2275);
and U2491 (N_2491,N_2271,N_2371);
or U2492 (N_2492,N_2393,N_2238);
nor U2493 (N_2493,N_2378,N_2369);
and U2494 (N_2494,N_2205,N_2239);
or U2495 (N_2495,N_2251,N_2324);
nand U2496 (N_2496,N_2290,N_2322);
and U2497 (N_2497,N_2343,N_2299);
nand U2498 (N_2498,N_2372,N_2354);
nor U2499 (N_2499,N_2288,N_2276);
nand U2500 (N_2500,N_2362,N_2244);
and U2501 (N_2501,N_2331,N_2358);
or U2502 (N_2502,N_2215,N_2245);
nor U2503 (N_2503,N_2346,N_2320);
and U2504 (N_2504,N_2328,N_2291);
and U2505 (N_2505,N_2260,N_2296);
nand U2506 (N_2506,N_2267,N_2340);
nor U2507 (N_2507,N_2242,N_2268);
and U2508 (N_2508,N_2396,N_2231);
nor U2509 (N_2509,N_2287,N_2257);
nand U2510 (N_2510,N_2366,N_2375);
or U2511 (N_2511,N_2397,N_2228);
nand U2512 (N_2512,N_2221,N_2273);
nand U2513 (N_2513,N_2246,N_2296);
and U2514 (N_2514,N_2258,N_2309);
and U2515 (N_2515,N_2210,N_2285);
nand U2516 (N_2516,N_2270,N_2325);
nor U2517 (N_2517,N_2347,N_2295);
and U2518 (N_2518,N_2384,N_2241);
nand U2519 (N_2519,N_2335,N_2322);
nand U2520 (N_2520,N_2274,N_2346);
and U2521 (N_2521,N_2284,N_2347);
and U2522 (N_2522,N_2245,N_2213);
and U2523 (N_2523,N_2374,N_2399);
and U2524 (N_2524,N_2232,N_2319);
nor U2525 (N_2525,N_2356,N_2272);
and U2526 (N_2526,N_2377,N_2287);
nor U2527 (N_2527,N_2204,N_2228);
and U2528 (N_2528,N_2368,N_2397);
nand U2529 (N_2529,N_2362,N_2341);
or U2530 (N_2530,N_2321,N_2371);
nor U2531 (N_2531,N_2216,N_2382);
and U2532 (N_2532,N_2375,N_2223);
or U2533 (N_2533,N_2361,N_2201);
nand U2534 (N_2534,N_2374,N_2328);
and U2535 (N_2535,N_2231,N_2398);
or U2536 (N_2536,N_2309,N_2374);
nand U2537 (N_2537,N_2368,N_2325);
or U2538 (N_2538,N_2360,N_2256);
or U2539 (N_2539,N_2341,N_2382);
nand U2540 (N_2540,N_2257,N_2372);
nand U2541 (N_2541,N_2204,N_2213);
and U2542 (N_2542,N_2254,N_2237);
nor U2543 (N_2543,N_2296,N_2396);
nor U2544 (N_2544,N_2377,N_2206);
nand U2545 (N_2545,N_2244,N_2221);
nand U2546 (N_2546,N_2321,N_2235);
nand U2547 (N_2547,N_2249,N_2355);
nand U2548 (N_2548,N_2269,N_2284);
or U2549 (N_2549,N_2305,N_2340);
nand U2550 (N_2550,N_2228,N_2384);
nor U2551 (N_2551,N_2369,N_2355);
nand U2552 (N_2552,N_2363,N_2307);
nor U2553 (N_2553,N_2388,N_2282);
or U2554 (N_2554,N_2399,N_2391);
or U2555 (N_2555,N_2301,N_2262);
and U2556 (N_2556,N_2341,N_2309);
or U2557 (N_2557,N_2269,N_2226);
nor U2558 (N_2558,N_2390,N_2367);
and U2559 (N_2559,N_2274,N_2213);
and U2560 (N_2560,N_2324,N_2385);
nand U2561 (N_2561,N_2244,N_2262);
nand U2562 (N_2562,N_2318,N_2275);
and U2563 (N_2563,N_2259,N_2238);
nand U2564 (N_2564,N_2381,N_2294);
nand U2565 (N_2565,N_2293,N_2392);
or U2566 (N_2566,N_2221,N_2337);
nor U2567 (N_2567,N_2277,N_2342);
nor U2568 (N_2568,N_2381,N_2338);
nor U2569 (N_2569,N_2242,N_2272);
and U2570 (N_2570,N_2214,N_2239);
and U2571 (N_2571,N_2202,N_2257);
or U2572 (N_2572,N_2215,N_2360);
nand U2573 (N_2573,N_2283,N_2261);
nor U2574 (N_2574,N_2257,N_2382);
nor U2575 (N_2575,N_2350,N_2318);
nand U2576 (N_2576,N_2277,N_2305);
nand U2577 (N_2577,N_2390,N_2234);
or U2578 (N_2578,N_2372,N_2310);
nand U2579 (N_2579,N_2262,N_2390);
or U2580 (N_2580,N_2271,N_2269);
nand U2581 (N_2581,N_2385,N_2386);
or U2582 (N_2582,N_2261,N_2235);
nand U2583 (N_2583,N_2364,N_2276);
nor U2584 (N_2584,N_2379,N_2227);
nor U2585 (N_2585,N_2212,N_2313);
nand U2586 (N_2586,N_2344,N_2207);
or U2587 (N_2587,N_2224,N_2242);
or U2588 (N_2588,N_2297,N_2340);
and U2589 (N_2589,N_2213,N_2365);
or U2590 (N_2590,N_2262,N_2376);
nor U2591 (N_2591,N_2351,N_2361);
nand U2592 (N_2592,N_2270,N_2209);
nor U2593 (N_2593,N_2262,N_2392);
or U2594 (N_2594,N_2377,N_2360);
nor U2595 (N_2595,N_2265,N_2364);
and U2596 (N_2596,N_2271,N_2241);
nor U2597 (N_2597,N_2345,N_2399);
or U2598 (N_2598,N_2281,N_2223);
or U2599 (N_2599,N_2325,N_2227);
and U2600 (N_2600,N_2409,N_2427);
and U2601 (N_2601,N_2507,N_2578);
nor U2602 (N_2602,N_2486,N_2589);
nand U2603 (N_2603,N_2525,N_2544);
or U2604 (N_2604,N_2562,N_2433);
nand U2605 (N_2605,N_2460,N_2450);
or U2606 (N_2606,N_2476,N_2453);
or U2607 (N_2607,N_2466,N_2521);
nor U2608 (N_2608,N_2502,N_2595);
and U2609 (N_2609,N_2551,N_2526);
nand U2610 (N_2610,N_2567,N_2559);
and U2611 (N_2611,N_2423,N_2556);
nand U2612 (N_2612,N_2419,N_2594);
nand U2613 (N_2613,N_2519,N_2527);
nor U2614 (N_2614,N_2553,N_2477);
nor U2615 (N_2615,N_2541,N_2547);
nor U2616 (N_2616,N_2542,N_2407);
or U2617 (N_2617,N_2443,N_2574);
nor U2618 (N_2618,N_2517,N_2588);
or U2619 (N_2619,N_2463,N_2456);
nand U2620 (N_2620,N_2508,N_2487);
nand U2621 (N_2621,N_2441,N_2585);
nor U2622 (N_2622,N_2451,N_2492);
or U2623 (N_2623,N_2418,N_2566);
or U2624 (N_2624,N_2429,N_2509);
xor U2625 (N_2625,N_2415,N_2572);
or U2626 (N_2626,N_2532,N_2428);
nand U2627 (N_2627,N_2454,N_2472);
nor U2628 (N_2628,N_2539,N_2555);
nor U2629 (N_2629,N_2400,N_2599);
or U2630 (N_2630,N_2565,N_2446);
nor U2631 (N_2631,N_2505,N_2596);
nand U2632 (N_2632,N_2564,N_2404);
nand U2633 (N_2633,N_2401,N_2490);
and U2634 (N_2634,N_2590,N_2455);
or U2635 (N_2635,N_2437,N_2436);
or U2636 (N_2636,N_2405,N_2501);
nand U2637 (N_2637,N_2425,N_2563);
or U2638 (N_2638,N_2471,N_2503);
or U2639 (N_2639,N_2438,N_2481);
and U2640 (N_2640,N_2430,N_2432);
nand U2641 (N_2641,N_2518,N_2560);
nor U2642 (N_2642,N_2411,N_2579);
nor U2643 (N_2643,N_2554,N_2537);
nor U2644 (N_2644,N_2403,N_2488);
nor U2645 (N_2645,N_2420,N_2422);
and U2646 (N_2646,N_2511,N_2546);
or U2647 (N_2647,N_2474,N_2557);
and U2648 (N_2648,N_2410,N_2449);
and U2649 (N_2649,N_2484,N_2458);
and U2650 (N_2650,N_2402,N_2470);
nand U2651 (N_2651,N_2483,N_2597);
or U2652 (N_2652,N_2442,N_2576);
nand U2653 (N_2653,N_2457,N_2431);
nand U2654 (N_2654,N_2582,N_2558);
nand U2655 (N_2655,N_2584,N_2489);
nor U2656 (N_2656,N_2513,N_2533);
nor U2657 (N_2657,N_2491,N_2467);
nand U2658 (N_2658,N_2468,N_2552);
nand U2659 (N_2659,N_2408,N_2529);
nand U2660 (N_2660,N_2591,N_2448);
nand U2661 (N_2661,N_2440,N_2497);
nand U2662 (N_2662,N_2478,N_2495);
nand U2663 (N_2663,N_2499,N_2516);
nor U2664 (N_2664,N_2549,N_2462);
and U2665 (N_2665,N_2514,N_2452);
and U2666 (N_2666,N_2461,N_2583);
nor U2667 (N_2667,N_2538,N_2577);
nand U2668 (N_2668,N_2473,N_2498);
nor U2669 (N_2669,N_2580,N_2475);
and U2670 (N_2670,N_2439,N_2573);
or U2671 (N_2671,N_2550,N_2587);
and U2672 (N_2672,N_2531,N_2523);
nand U2673 (N_2673,N_2413,N_2575);
xnor U2674 (N_2674,N_2569,N_2540);
or U2675 (N_2675,N_2434,N_2480);
or U2676 (N_2676,N_2479,N_2485);
nor U2677 (N_2677,N_2414,N_2530);
nor U2678 (N_2678,N_2464,N_2548);
nand U2679 (N_2679,N_2543,N_2571);
and U2680 (N_2680,N_2592,N_2482);
and U2681 (N_2681,N_2524,N_2417);
and U2682 (N_2682,N_2506,N_2581);
nand U2683 (N_2683,N_2512,N_2522);
and U2684 (N_2684,N_2510,N_2416);
nand U2685 (N_2685,N_2412,N_2515);
and U2686 (N_2686,N_2586,N_2561);
or U2687 (N_2687,N_2421,N_2447);
nand U2688 (N_2688,N_2435,N_2465);
nand U2689 (N_2689,N_2496,N_2444);
and U2690 (N_2690,N_2534,N_2445);
nor U2691 (N_2691,N_2528,N_2424);
nand U2692 (N_2692,N_2494,N_2570);
or U2693 (N_2693,N_2568,N_2406);
nor U2694 (N_2694,N_2598,N_2520);
nand U2695 (N_2695,N_2593,N_2459);
and U2696 (N_2696,N_2500,N_2469);
nor U2697 (N_2697,N_2504,N_2536);
and U2698 (N_2698,N_2535,N_2545);
and U2699 (N_2699,N_2493,N_2426);
nand U2700 (N_2700,N_2415,N_2524);
or U2701 (N_2701,N_2514,N_2447);
or U2702 (N_2702,N_2567,N_2435);
nor U2703 (N_2703,N_2407,N_2479);
nor U2704 (N_2704,N_2432,N_2477);
and U2705 (N_2705,N_2588,N_2427);
nor U2706 (N_2706,N_2448,N_2484);
nor U2707 (N_2707,N_2456,N_2484);
or U2708 (N_2708,N_2468,N_2526);
and U2709 (N_2709,N_2458,N_2488);
and U2710 (N_2710,N_2430,N_2494);
and U2711 (N_2711,N_2549,N_2437);
or U2712 (N_2712,N_2508,N_2512);
nor U2713 (N_2713,N_2500,N_2513);
nor U2714 (N_2714,N_2522,N_2468);
xor U2715 (N_2715,N_2524,N_2430);
nand U2716 (N_2716,N_2503,N_2588);
nor U2717 (N_2717,N_2450,N_2566);
and U2718 (N_2718,N_2414,N_2430);
or U2719 (N_2719,N_2493,N_2519);
nand U2720 (N_2720,N_2598,N_2571);
or U2721 (N_2721,N_2587,N_2467);
and U2722 (N_2722,N_2529,N_2465);
and U2723 (N_2723,N_2454,N_2437);
nand U2724 (N_2724,N_2405,N_2516);
nand U2725 (N_2725,N_2518,N_2495);
nor U2726 (N_2726,N_2446,N_2454);
and U2727 (N_2727,N_2538,N_2506);
or U2728 (N_2728,N_2483,N_2555);
or U2729 (N_2729,N_2460,N_2574);
nor U2730 (N_2730,N_2546,N_2505);
or U2731 (N_2731,N_2535,N_2537);
nor U2732 (N_2732,N_2510,N_2559);
or U2733 (N_2733,N_2581,N_2570);
nor U2734 (N_2734,N_2410,N_2555);
or U2735 (N_2735,N_2446,N_2502);
and U2736 (N_2736,N_2496,N_2520);
nand U2737 (N_2737,N_2593,N_2403);
or U2738 (N_2738,N_2427,N_2570);
nand U2739 (N_2739,N_2490,N_2537);
nor U2740 (N_2740,N_2594,N_2463);
nor U2741 (N_2741,N_2417,N_2521);
nand U2742 (N_2742,N_2573,N_2462);
nor U2743 (N_2743,N_2400,N_2593);
nor U2744 (N_2744,N_2422,N_2589);
or U2745 (N_2745,N_2414,N_2445);
nor U2746 (N_2746,N_2510,N_2533);
and U2747 (N_2747,N_2492,N_2493);
or U2748 (N_2748,N_2520,N_2587);
or U2749 (N_2749,N_2589,N_2449);
or U2750 (N_2750,N_2462,N_2413);
and U2751 (N_2751,N_2569,N_2442);
or U2752 (N_2752,N_2579,N_2566);
and U2753 (N_2753,N_2580,N_2508);
nor U2754 (N_2754,N_2482,N_2491);
or U2755 (N_2755,N_2478,N_2526);
nand U2756 (N_2756,N_2524,N_2556);
nand U2757 (N_2757,N_2513,N_2422);
nand U2758 (N_2758,N_2400,N_2404);
nor U2759 (N_2759,N_2490,N_2460);
and U2760 (N_2760,N_2426,N_2412);
nand U2761 (N_2761,N_2489,N_2491);
nor U2762 (N_2762,N_2593,N_2463);
and U2763 (N_2763,N_2560,N_2572);
or U2764 (N_2764,N_2471,N_2464);
nand U2765 (N_2765,N_2503,N_2574);
and U2766 (N_2766,N_2573,N_2581);
nor U2767 (N_2767,N_2414,N_2541);
nor U2768 (N_2768,N_2406,N_2430);
nor U2769 (N_2769,N_2465,N_2491);
or U2770 (N_2770,N_2570,N_2447);
nor U2771 (N_2771,N_2464,N_2538);
and U2772 (N_2772,N_2430,N_2523);
and U2773 (N_2773,N_2515,N_2546);
or U2774 (N_2774,N_2530,N_2537);
nand U2775 (N_2775,N_2461,N_2462);
and U2776 (N_2776,N_2587,N_2499);
nor U2777 (N_2777,N_2583,N_2527);
nor U2778 (N_2778,N_2481,N_2471);
nor U2779 (N_2779,N_2433,N_2524);
nand U2780 (N_2780,N_2582,N_2426);
nor U2781 (N_2781,N_2404,N_2471);
or U2782 (N_2782,N_2499,N_2569);
or U2783 (N_2783,N_2418,N_2595);
nand U2784 (N_2784,N_2556,N_2501);
nand U2785 (N_2785,N_2580,N_2575);
nand U2786 (N_2786,N_2445,N_2588);
nand U2787 (N_2787,N_2449,N_2564);
nor U2788 (N_2788,N_2405,N_2572);
nand U2789 (N_2789,N_2571,N_2584);
nand U2790 (N_2790,N_2475,N_2479);
nand U2791 (N_2791,N_2485,N_2546);
and U2792 (N_2792,N_2539,N_2503);
nor U2793 (N_2793,N_2506,N_2570);
and U2794 (N_2794,N_2461,N_2568);
and U2795 (N_2795,N_2434,N_2435);
or U2796 (N_2796,N_2462,N_2513);
and U2797 (N_2797,N_2525,N_2409);
nand U2798 (N_2798,N_2478,N_2505);
nor U2799 (N_2799,N_2436,N_2530);
nand U2800 (N_2800,N_2780,N_2689);
nor U2801 (N_2801,N_2736,N_2798);
nor U2802 (N_2802,N_2762,N_2748);
and U2803 (N_2803,N_2675,N_2737);
nand U2804 (N_2804,N_2754,N_2769);
or U2805 (N_2805,N_2683,N_2687);
or U2806 (N_2806,N_2646,N_2793);
nand U2807 (N_2807,N_2701,N_2786);
xnor U2808 (N_2808,N_2613,N_2690);
nor U2809 (N_2809,N_2697,N_2691);
nor U2810 (N_2810,N_2696,N_2787);
or U2811 (N_2811,N_2742,N_2650);
nand U2812 (N_2812,N_2700,N_2681);
nand U2813 (N_2813,N_2710,N_2686);
nand U2814 (N_2814,N_2728,N_2743);
nor U2815 (N_2815,N_2712,N_2719);
nor U2816 (N_2816,N_2771,N_2717);
or U2817 (N_2817,N_2789,N_2795);
xnor U2818 (N_2818,N_2661,N_2722);
and U2819 (N_2819,N_2709,N_2669);
nor U2820 (N_2820,N_2617,N_2635);
xor U2821 (N_2821,N_2667,N_2643);
nor U2822 (N_2822,N_2615,N_2633);
and U2823 (N_2823,N_2725,N_2660);
nand U2824 (N_2824,N_2738,N_2665);
nand U2825 (N_2825,N_2799,N_2677);
nand U2826 (N_2826,N_2674,N_2778);
nor U2827 (N_2827,N_2735,N_2772);
nor U2828 (N_2828,N_2761,N_2783);
nand U2829 (N_2829,N_2682,N_2776);
and U2830 (N_2830,N_2666,N_2781);
nor U2831 (N_2831,N_2610,N_2631);
or U2832 (N_2832,N_2708,N_2653);
nand U2833 (N_2833,N_2622,N_2758);
and U2834 (N_2834,N_2618,N_2760);
and U2835 (N_2835,N_2628,N_2785);
nor U2836 (N_2836,N_2768,N_2611);
nand U2837 (N_2837,N_2766,N_2605);
or U2838 (N_2838,N_2692,N_2641);
or U2839 (N_2839,N_2625,N_2705);
and U2840 (N_2840,N_2729,N_2680);
and U2841 (N_2841,N_2648,N_2656);
nand U2842 (N_2842,N_2797,N_2654);
nand U2843 (N_2843,N_2619,N_2688);
or U2844 (N_2844,N_2627,N_2779);
or U2845 (N_2845,N_2637,N_2733);
nand U2846 (N_2846,N_2752,N_2732);
nor U2847 (N_2847,N_2621,N_2607);
and U2848 (N_2848,N_2698,N_2788);
or U2849 (N_2849,N_2706,N_2600);
and U2850 (N_2850,N_2759,N_2639);
nand U2851 (N_2851,N_2757,N_2658);
nand U2852 (N_2852,N_2749,N_2745);
nand U2853 (N_2853,N_2636,N_2773);
xnor U2854 (N_2854,N_2649,N_2770);
nand U2855 (N_2855,N_2676,N_2671);
and U2856 (N_2856,N_2782,N_2703);
or U2857 (N_2857,N_2644,N_2734);
and U2858 (N_2858,N_2704,N_2731);
or U2859 (N_2859,N_2624,N_2747);
xor U2860 (N_2860,N_2629,N_2796);
and U2861 (N_2861,N_2684,N_2604);
xor U2862 (N_2862,N_2694,N_2645);
and U2863 (N_2863,N_2640,N_2721);
and U2864 (N_2864,N_2744,N_2713);
nand U2865 (N_2865,N_2647,N_2652);
nand U2866 (N_2866,N_2784,N_2727);
and U2867 (N_2867,N_2601,N_2606);
nor U2868 (N_2868,N_2711,N_2791);
nand U2869 (N_2869,N_2634,N_2741);
nor U2870 (N_2870,N_2774,N_2756);
and U2871 (N_2871,N_2672,N_2679);
nor U2872 (N_2872,N_2699,N_2726);
nand U2873 (N_2873,N_2724,N_2664);
or U2874 (N_2874,N_2638,N_2657);
nor U2875 (N_2875,N_2775,N_2602);
and U2876 (N_2876,N_2651,N_2632);
nand U2877 (N_2877,N_2609,N_2707);
nand U2878 (N_2878,N_2763,N_2670);
nor U2879 (N_2879,N_2751,N_2723);
nor U2880 (N_2880,N_2767,N_2720);
nand U2881 (N_2881,N_2765,N_2659);
and U2882 (N_2882,N_2668,N_2673);
or U2883 (N_2883,N_2718,N_2612);
nor U2884 (N_2884,N_2655,N_2603);
xor U2885 (N_2885,N_2630,N_2739);
nor U2886 (N_2886,N_2608,N_2702);
and U2887 (N_2887,N_2662,N_2685);
nand U2888 (N_2888,N_2777,N_2663);
or U2889 (N_2889,N_2623,N_2730);
nor U2890 (N_2890,N_2693,N_2750);
and U2891 (N_2891,N_2620,N_2614);
nor U2892 (N_2892,N_2716,N_2715);
nand U2893 (N_2893,N_2764,N_2746);
nand U2894 (N_2894,N_2794,N_2626);
nand U2895 (N_2895,N_2755,N_2616);
and U2896 (N_2896,N_2790,N_2714);
and U2897 (N_2897,N_2695,N_2642);
or U2898 (N_2898,N_2740,N_2753);
or U2899 (N_2899,N_2792,N_2678);
nand U2900 (N_2900,N_2752,N_2776);
and U2901 (N_2901,N_2757,N_2784);
nor U2902 (N_2902,N_2794,N_2779);
or U2903 (N_2903,N_2718,N_2712);
and U2904 (N_2904,N_2766,N_2651);
and U2905 (N_2905,N_2736,N_2717);
and U2906 (N_2906,N_2790,N_2692);
nand U2907 (N_2907,N_2615,N_2607);
or U2908 (N_2908,N_2639,N_2717);
and U2909 (N_2909,N_2681,N_2771);
nor U2910 (N_2910,N_2648,N_2719);
nor U2911 (N_2911,N_2661,N_2606);
nand U2912 (N_2912,N_2742,N_2693);
nand U2913 (N_2913,N_2749,N_2750);
nor U2914 (N_2914,N_2764,N_2750);
or U2915 (N_2915,N_2793,N_2605);
and U2916 (N_2916,N_2614,N_2694);
nor U2917 (N_2917,N_2660,N_2665);
or U2918 (N_2918,N_2658,N_2707);
and U2919 (N_2919,N_2721,N_2752);
and U2920 (N_2920,N_2664,N_2645);
nand U2921 (N_2921,N_2620,N_2618);
nand U2922 (N_2922,N_2692,N_2680);
or U2923 (N_2923,N_2682,N_2782);
and U2924 (N_2924,N_2624,N_2735);
and U2925 (N_2925,N_2654,N_2627);
or U2926 (N_2926,N_2735,N_2664);
nand U2927 (N_2927,N_2635,N_2607);
and U2928 (N_2928,N_2647,N_2672);
nand U2929 (N_2929,N_2612,N_2683);
and U2930 (N_2930,N_2675,N_2609);
and U2931 (N_2931,N_2665,N_2638);
nor U2932 (N_2932,N_2638,N_2790);
and U2933 (N_2933,N_2728,N_2670);
nor U2934 (N_2934,N_2771,N_2752);
nand U2935 (N_2935,N_2706,N_2774);
nand U2936 (N_2936,N_2758,N_2653);
nand U2937 (N_2937,N_2606,N_2684);
nor U2938 (N_2938,N_2762,N_2731);
and U2939 (N_2939,N_2671,N_2799);
nand U2940 (N_2940,N_2706,N_2673);
or U2941 (N_2941,N_2766,N_2664);
nor U2942 (N_2942,N_2738,N_2787);
and U2943 (N_2943,N_2739,N_2760);
nor U2944 (N_2944,N_2605,N_2790);
nor U2945 (N_2945,N_2649,N_2749);
nand U2946 (N_2946,N_2606,N_2741);
or U2947 (N_2947,N_2667,N_2678);
and U2948 (N_2948,N_2779,N_2665);
nand U2949 (N_2949,N_2604,N_2733);
and U2950 (N_2950,N_2706,N_2768);
nor U2951 (N_2951,N_2777,N_2784);
nor U2952 (N_2952,N_2703,N_2768);
nor U2953 (N_2953,N_2660,N_2632);
nor U2954 (N_2954,N_2773,N_2618);
nor U2955 (N_2955,N_2662,N_2783);
nor U2956 (N_2956,N_2650,N_2752);
or U2957 (N_2957,N_2754,N_2744);
and U2958 (N_2958,N_2712,N_2672);
nor U2959 (N_2959,N_2614,N_2726);
nor U2960 (N_2960,N_2749,N_2714);
nor U2961 (N_2961,N_2778,N_2774);
nor U2962 (N_2962,N_2624,N_2692);
and U2963 (N_2963,N_2674,N_2790);
or U2964 (N_2964,N_2749,N_2755);
nand U2965 (N_2965,N_2639,N_2789);
nand U2966 (N_2966,N_2697,N_2657);
nor U2967 (N_2967,N_2724,N_2620);
nor U2968 (N_2968,N_2627,N_2783);
and U2969 (N_2969,N_2716,N_2625);
and U2970 (N_2970,N_2628,N_2617);
xnor U2971 (N_2971,N_2701,N_2680);
or U2972 (N_2972,N_2602,N_2621);
nand U2973 (N_2973,N_2785,N_2735);
nand U2974 (N_2974,N_2703,N_2739);
nor U2975 (N_2975,N_2771,N_2639);
and U2976 (N_2976,N_2780,N_2713);
or U2977 (N_2977,N_2639,N_2779);
nand U2978 (N_2978,N_2778,N_2682);
and U2979 (N_2979,N_2617,N_2637);
nor U2980 (N_2980,N_2667,N_2645);
nor U2981 (N_2981,N_2603,N_2764);
and U2982 (N_2982,N_2697,N_2655);
nor U2983 (N_2983,N_2621,N_2649);
nand U2984 (N_2984,N_2723,N_2759);
or U2985 (N_2985,N_2701,N_2704);
nand U2986 (N_2986,N_2617,N_2650);
and U2987 (N_2987,N_2618,N_2634);
nand U2988 (N_2988,N_2618,N_2762);
nor U2989 (N_2989,N_2763,N_2633);
nor U2990 (N_2990,N_2719,N_2692);
nor U2991 (N_2991,N_2713,N_2760);
and U2992 (N_2992,N_2669,N_2692);
nor U2993 (N_2993,N_2793,N_2777);
nand U2994 (N_2994,N_2747,N_2779);
or U2995 (N_2995,N_2715,N_2747);
and U2996 (N_2996,N_2641,N_2773);
and U2997 (N_2997,N_2725,N_2698);
nand U2998 (N_2998,N_2730,N_2725);
nor U2999 (N_2999,N_2745,N_2703);
nor U3000 (N_3000,N_2909,N_2953);
nand U3001 (N_3001,N_2878,N_2907);
nor U3002 (N_3002,N_2916,N_2877);
and U3003 (N_3003,N_2930,N_2847);
or U3004 (N_3004,N_2820,N_2856);
nand U3005 (N_3005,N_2974,N_2897);
nor U3006 (N_3006,N_2873,N_2830);
nor U3007 (N_3007,N_2908,N_2813);
and U3008 (N_3008,N_2898,N_2901);
or U3009 (N_3009,N_2894,N_2848);
nand U3010 (N_3010,N_2927,N_2812);
and U3011 (N_3011,N_2838,N_2976);
nor U3012 (N_3012,N_2867,N_2837);
and U3013 (N_3013,N_2925,N_2824);
and U3014 (N_3014,N_2851,N_2924);
nor U3015 (N_3015,N_2825,N_2922);
or U3016 (N_3016,N_2859,N_2979);
or U3017 (N_3017,N_2884,N_2862);
and U3018 (N_3018,N_2842,N_2886);
or U3019 (N_3019,N_2810,N_2822);
nor U3020 (N_3020,N_2855,N_2872);
or U3021 (N_3021,N_2891,N_2947);
nor U3022 (N_3022,N_2803,N_2941);
and U3023 (N_3023,N_2817,N_2943);
nor U3024 (N_3024,N_2915,N_2971);
and U3025 (N_3025,N_2942,N_2883);
and U3026 (N_3026,N_2945,N_2966);
and U3027 (N_3027,N_2964,N_2931);
nor U3028 (N_3028,N_2829,N_2879);
nor U3029 (N_3029,N_2954,N_2984);
nor U3030 (N_3030,N_2962,N_2814);
nor U3031 (N_3031,N_2918,N_2904);
nand U3032 (N_3032,N_2973,N_2977);
nand U3033 (N_3033,N_2928,N_2832);
or U3034 (N_3034,N_2895,N_2853);
xnor U3035 (N_3035,N_2934,N_2999);
nor U3036 (N_3036,N_2880,N_2885);
and U3037 (N_3037,N_2998,N_2882);
nand U3038 (N_3038,N_2949,N_2913);
nand U3039 (N_3039,N_2874,N_2957);
nand U3040 (N_3040,N_2911,N_2818);
or U3041 (N_3041,N_2811,N_2960);
xnor U3042 (N_3042,N_2933,N_2804);
and U3043 (N_3043,N_2869,N_2961);
or U3044 (N_3044,N_2846,N_2835);
nand U3045 (N_3045,N_2956,N_2932);
nor U3046 (N_3046,N_2887,N_2863);
nand U3047 (N_3047,N_2819,N_2840);
nand U3048 (N_3048,N_2967,N_2997);
or U3049 (N_3049,N_2965,N_2975);
and U3050 (N_3050,N_2850,N_2866);
nand U3051 (N_3051,N_2809,N_2988);
nor U3052 (N_3052,N_2923,N_2944);
nand U3053 (N_3053,N_2919,N_2900);
nand U3054 (N_3054,N_2910,N_2861);
or U3055 (N_3055,N_2969,N_2937);
nand U3056 (N_3056,N_2994,N_2963);
and U3057 (N_3057,N_2821,N_2936);
nand U3058 (N_3058,N_2806,N_2992);
and U3059 (N_3059,N_2905,N_2860);
nand U3060 (N_3060,N_2876,N_2805);
and U3061 (N_3061,N_2870,N_2959);
nand U3062 (N_3062,N_2980,N_2987);
nand U3063 (N_3063,N_2844,N_2968);
nor U3064 (N_3064,N_2868,N_2871);
or U3065 (N_3065,N_2986,N_2836);
and U3066 (N_3066,N_2807,N_2935);
nor U3067 (N_3067,N_2982,N_2865);
and U3068 (N_3068,N_2828,N_2938);
or U3069 (N_3069,N_2906,N_2801);
or U3070 (N_3070,N_2823,N_2995);
nand U3071 (N_3071,N_2940,N_2948);
xor U3072 (N_3072,N_2991,N_2889);
nor U3073 (N_3073,N_2826,N_2890);
or U3074 (N_3074,N_2972,N_2858);
or U3075 (N_3075,N_2926,N_2802);
or U3076 (N_3076,N_2834,N_2833);
nor U3077 (N_3077,N_2946,N_2996);
nand U3078 (N_3078,N_2983,N_2951);
nor U3079 (N_3079,N_2857,N_2950);
nor U3080 (N_3080,N_2815,N_2981);
nor U3081 (N_3081,N_2808,N_2917);
and U3082 (N_3082,N_2849,N_2978);
and U3083 (N_3083,N_2990,N_2893);
nor U3084 (N_3084,N_2902,N_2843);
nand U3085 (N_3085,N_2921,N_2841);
or U3086 (N_3086,N_2955,N_2816);
and U3087 (N_3087,N_2875,N_2939);
nand U3088 (N_3088,N_2800,N_2831);
and U3089 (N_3089,N_2881,N_2929);
nand U3090 (N_3090,N_2845,N_2864);
nor U3091 (N_3091,N_2903,N_2989);
nor U3092 (N_3092,N_2899,N_2952);
nor U3093 (N_3093,N_2970,N_2914);
nand U3094 (N_3094,N_2985,N_2912);
nor U3095 (N_3095,N_2920,N_2839);
nand U3096 (N_3096,N_2958,N_2852);
nand U3097 (N_3097,N_2993,N_2892);
nand U3098 (N_3098,N_2896,N_2827);
and U3099 (N_3099,N_2888,N_2854);
and U3100 (N_3100,N_2904,N_2917);
or U3101 (N_3101,N_2840,N_2967);
nor U3102 (N_3102,N_2986,N_2939);
or U3103 (N_3103,N_2897,N_2844);
or U3104 (N_3104,N_2881,N_2800);
nand U3105 (N_3105,N_2839,N_2885);
and U3106 (N_3106,N_2923,N_2981);
nand U3107 (N_3107,N_2932,N_2863);
and U3108 (N_3108,N_2944,N_2927);
nor U3109 (N_3109,N_2929,N_2990);
and U3110 (N_3110,N_2902,N_2989);
and U3111 (N_3111,N_2824,N_2839);
nor U3112 (N_3112,N_2961,N_2863);
or U3113 (N_3113,N_2984,N_2902);
and U3114 (N_3114,N_2808,N_2885);
nor U3115 (N_3115,N_2881,N_2903);
nand U3116 (N_3116,N_2986,N_2997);
nand U3117 (N_3117,N_2945,N_2886);
nor U3118 (N_3118,N_2860,N_2904);
nor U3119 (N_3119,N_2867,N_2848);
nor U3120 (N_3120,N_2921,N_2826);
or U3121 (N_3121,N_2862,N_2836);
nand U3122 (N_3122,N_2805,N_2938);
nor U3123 (N_3123,N_2859,N_2821);
or U3124 (N_3124,N_2898,N_2819);
nor U3125 (N_3125,N_2923,N_2913);
nor U3126 (N_3126,N_2920,N_2967);
or U3127 (N_3127,N_2865,N_2886);
or U3128 (N_3128,N_2865,N_2903);
nand U3129 (N_3129,N_2987,N_2866);
nand U3130 (N_3130,N_2995,N_2916);
or U3131 (N_3131,N_2990,N_2856);
and U3132 (N_3132,N_2898,N_2877);
or U3133 (N_3133,N_2865,N_2849);
and U3134 (N_3134,N_2937,N_2839);
or U3135 (N_3135,N_2811,N_2954);
and U3136 (N_3136,N_2965,N_2894);
or U3137 (N_3137,N_2932,N_2896);
or U3138 (N_3138,N_2844,N_2832);
nor U3139 (N_3139,N_2837,N_2885);
nand U3140 (N_3140,N_2917,N_2909);
or U3141 (N_3141,N_2833,N_2947);
nand U3142 (N_3142,N_2848,N_2811);
nor U3143 (N_3143,N_2842,N_2903);
nand U3144 (N_3144,N_2886,N_2805);
nand U3145 (N_3145,N_2828,N_2950);
nand U3146 (N_3146,N_2987,N_2967);
nand U3147 (N_3147,N_2962,N_2847);
nand U3148 (N_3148,N_2947,N_2945);
and U3149 (N_3149,N_2978,N_2945);
and U3150 (N_3150,N_2878,N_2839);
nor U3151 (N_3151,N_2901,N_2938);
or U3152 (N_3152,N_2976,N_2882);
or U3153 (N_3153,N_2914,N_2953);
nor U3154 (N_3154,N_2932,N_2817);
nand U3155 (N_3155,N_2829,N_2944);
nor U3156 (N_3156,N_2981,N_2944);
nor U3157 (N_3157,N_2929,N_2840);
nand U3158 (N_3158,N_2892,N_2983);
and U3159 (N_3159,N_2880,N_2854);
nor U3160 (N_3160,N_2820,N_2977);
or U3161 (N_3161,N_2897,N_2850);
and U3162 (N_3162,N_2844,N_2957);
nor U3163 (N_3163,N_2885,N_2817);
or U3164 (N_3164,N_2964,N_2892);
nor U3165 (N_3165,N_2947,N_2905);
and U3166 (N_3166,N_2933,N_2949);
nand U3167 (N_3167,N_2916,N_2961);
nand U3168 (N_3168,N_2985,N_2844);
or U3169 (N_3169,N_2874,N_2839);
or U3170 (N_3170,N_2992,N_2801);
or U3171 (N_3171,N_2917,N_2885);
xor U3172 (N_3172,N_2919,N_2819);
nor U3173 (N_3173,N_2929,N_2863);
or U3174 (N_3174,N_2928,N_2886);
and U3175 (N_3175,N_2911,N_2917);
nand U3176 (N_3176,N_2853,N_2837);
nand U3177 (N_3177,N_2809,N_2906);
nand U3178 (N_3178,N_2990,N_2821);
nor U3179 (N_3179,N_2886,N_2858);
or U3180 (N_3180,N_2820,N_2840);
or U3181 (N_3181,N_2967,N_2966);
nor U3182 (N_3182,N_2854,N_2924);
nor U3183 (N_3183,N_2842,N_2925);
nor U3184 (N_3184,N_2819,N_2802);
nor U3185 (N_3185,N_2963,N_2908);
nand U3186 (N_3186,N_2904,N_2896);
and U3187 (N_3187,N_2916,N_2817);
nor U3188 (N_3188,N_2880,N_2847);
and U3189 (N_3189,N_2874,N_2878);
or U3190 (N_3190,N_2866,N_2950);
or U3191 (N_3191,N_2869,N_2893);
nor U3192 (N_3192,N_2990,N_2855);
nor U3193 (N_3193,N_2952,N_2878);
nand U3194 (N_3194,N_2974,N_2869);
and U3195 (N_3195,N_2911,N_2899);
nand U3196 (N_3196,N_2884,N_2879);
or U3197 (N_3197,N_2958,N_2813);
nand U3198 (N_3198,N_2831,N_2989);
nand U3199 (N_3199,N_2887,N_2977);
nor U3200 (N_3200,N_3044,N_3058);
nand U3201 (N_3201,N_3163,N_3195);
nand U3202 (N_3202,N_3008,N_3009);
or U3203 (N_3203,N_3057,N_3090);
nor U3204 (N_3204,N_3066,N_3134);
and U3205 (N_3205,N_3020,N_3122);
nor U3206 (N_3206,N_3086,N_3186);
nand U3207 (N_3207,N_3055,N_3101);
nor U3208 (N_3208,N_3080,N_3091);
nor U3209 (N_3209,N_3072,N_3171);
and U3210 (N_3210,N_3099,N_3102);
or U3211 (N_3211,N_3187,N_3159);
and U3212 (N_3212,N_3000,N_3136);
nor U3213 (N_3213,N_3184,N_3193);
nand U3214 (N_3214,N_3125,N_3160);
and U3215 (N_3215,N_3164,N_3036);
or U3216 (N_3216,N_3010,N_3165);
and U3217 (N_3217,N_3022,N_3005);
nand U3218 (N_3218,N_3061,N_3052);
nor U3219 (N_3219,N_3069,N_3140);
and U3220 (N_3220,N_3083,N_3162);
nor U3221 (N_3221,N_3161,N_3188);
or U3222 (N_3222,N_3096,N_3149);
nor U3223 (N_3223,N_3157,N_3176);
and U3224 (N_3224,N_3037,N_3143);
or U3225 (N_3225,N_3146,N_3130);
nand U3226 (N_3226,N_3013,N_3041);
nor U3227 (N_3227,N_3097,N_3035);
nand U3228 (N_3228,N_3132,N_3135);
and U3229 (N_3229,N_3119,N_3084);
nand U3230 (N_3230,N_3133,N_3172);
nand U3231 (N_3231,N_3145,N_3088);
or U3232 (N_3232,N_3060,N_3137);
and U3233 (N_3233,N_3003,N_3199);
or U3234 (N_3234,N_3026,N_3039);
and U3235 (N_3235,N_3148,N_3100);
or U3236 (N_3236,N_3175,N_3150);
nand U3237 (N_3237,N_3004,N_3177);
or U3238 (N_3238,N_3007,N_3185);
or U3239 (N_3239,N_3023,N_3049);
or U3240 (N_3240,N_3179,N_3191);
or U3241 (N_3241,N_3151,N_3012);
and U3242 (N_3242,N_3015,N_3028);
and U3243 (N_3243,N_3105,N_3112);
nor U3244 (N_3244,N_3152,N_3183);
nand U3245 (N_3245,N_3181,N_3095);
or U3246 (N_3246,N_3138,N_3129);
nand U3247 (N_3247,N_3045,N_3131);
and U3248 (N_3248,N_3128,N_3018);
nand U3249 (N_3249,N_3021,N_3114);
nor U3250 (N_3250,N_3124,N_3142);
or U3251 (N_3251,N_3156,N_3081);
nand U3252 (N_3252,N_3115,N_3040);
nand U3253 (N_3253,N_3074,N_3032);
nand U3254 (N_3254,N_3190,N_3197);
nand U3255 (N_3255,N_3110,N_3111);
or U3256 (N_3256,N_3158,N_3048);
nor U3257 (N_3257,N_3141,N_3107);
nand U3258 (N_3258,N_3198,N_3071);
nor U3259 (N_3259,N_3079,N_3103);
nand U3260 (N_3260,N_3062,N_3155);
and U3261 (N_3261,N_3168,N_3070);
or U3262 (N_3262,N_3068,N_3121);
nor U3263 (N_3263,N_3089,N_3067);
and U3264 (N_3264,N_3034,N_3180);
nand U3265 (N_3265,N_3082,N_3116);
and U3266 (N_3266,N_3031,N_3194);
nor U3267 (N_3267,N_3078,N_3027);
nand U3268 (N_3268,N_3033,N_3051);
and U3269 (N_3269,N_3038,N_3094);
and U3270 (N_3270,N_3092,N_3050);
and U3271 (N_3271,N_3056,N_3126);
nand U3272 (N_3272,N_3006,N_3014);
nor U3273 (N_3273,N_3030,N_3108);
nor U3274 (N_3274,N_3117,N_3167);
nor U3275 (N_3275,N_3196,N_3192);
or U3276 (N_3276,N_3063,N_3064);
nor U3277 (N_3277,N_3170,N_3144);
nand U3278 (N_3278,N_3073,N_3123);
or U3279 (N_3279,N_3169,N_3024);
and U3280 (N_3280,N_3029,N_3025);
and U3281 (N_3281,N_3182,N_3077);
and U3282 (N_3282,N_3053,N_3139);
or U3283 (N_3283,N_3109,N_3153);
nor U3284 (N_3284,N_3104,N_3001);
nor U3285 (N_3285,N_3046,N_3065);
nor U3286 (N_3286,N_3113,N_3166);
nand U3287 (N_3287,N_3178,N_3173);
nand U3288 (N_3288,N_3016,N_3002);
nor U3289 (N_3289,N_3047,N_3017);
nor U3290 (N_3290,N_3147,N_3059);
nor U3291 (N_3291,N_3019,N_3127);
nor U3292 (N_3292,N_3118,N_3043);
nand U3293 (N_3293,N_3106,N_3042);
nor U3294 (N_3294,N_3098,N_3075);
and U3295 (N_3295,N_3174,N_3120);
nor U3296 (N_3296,N_3054,N_3087);
nand U3297 (N_3297,N_3011,N_3076);
nor U3298 (N_3298,N_3189,N_3085);
and U3299 (N_3299,N_3093,N_3154);
nand U3300 (N_3300,N_3084,N_3183);
xnor U3301 (N_3301,N_3055,N_3179);
nor U3302 (N_3302,N_3194,N_3039);
nand U3303 (N_3303,N_3103,N_3197);
or U3304 (N_3304,N_3000,N_3045);
nor U3305 (N_3305,N_3194,N_3095);
or U3306 (N_3306,N_3020,N_3042);
nand U3307 (N_3307,N_3151,N_3138);
nand U3308 (N_3308,N_3017,N_3139);
nand U3309 (N_3309,N_3151,N_3053);
nand U3310 (N_3310,N_3056,N_3023);
nand U3311 (N_3311,N_3101,N_3020);
and U3312 (N_3312,N_3041,N_3196);
and U3313 (N_3313,N_3165,N_3000);
or U3314 (N_3314,N_3069,N_3146);
or U3315 (N_3315,N_3143,N_3086);
or U3316 (N_3316,N_3043,N_3004);
nand U3317 (N_3317,N_3124,N_3025);
and U3318 (N_3318,N_3085,N_3123);
or U3319 (N_3319,N_3023,N_3041);
nor U3320 (N_3320,N_3166,N_3065);
nand U3321 (N_3321,N_3134,N_3099);
nand U3322 (N_3322,N_3121,N_3091);
nand U3323 (N_3323,N_3019,N_3187);
nand U3324 (N_3324,N_3133,N_3136);
nor U3325 (N_3325,N_3010,N_3125);
nand U3326 (N_3326,N_3064,N_3170);
nor U3327 (N_3327,N_3041,N_3069);
nor U3328 (N_3328,N_3192,N_3124);
and U3329 (N_3329,N_3060,N_3046);
nor U3330 (N_3330,N_3038,N_3066);
or U3331 (N_3331,N_3068,N_3024);
nand U3332 (N_3332,N_3137,N_3102);
nor U3333 (N_3333,N_3129,N_3005);
nand U3334 (N_3334,N_3174,N_3171);
nand U3335 (N_3335,N_3109,N_3148);
and U3336 (N_3336,N_3008,N_3115);
nand U3337 (N_3337,N_3072,N_3018);
nor U3338 (N_3338,N_3033,N_3007);
and U3339 (N_3339,N_3056,N_3122);
nand U3340 (N_3340,N_3019,N_3156);
and U3341 (N_3341,N_3014,N_3005);
or U3342 (N_3342,N_3145,N_3097);
and U3343 (N_3343,N_3057,N_3128);
nor U3344 (N_3344,N_3058,N_3189);
or U3345 (N_3345,N_3061,N_3101);
or U3346 (N_3346,N_3176,N_3169);
nor U3347 (N_3347,N_3003,N_3070);
and U3348 (N_3348,N_3149,N_3074);
nand U3349 (N_3349,N_3152,N_3178);
or U3350 (N_3350,N_3108,N_3191);
or U3351 (N_3351,N_3061,N_3133);
nor U3352 (N_3352,N_3039,N_3128);
nor U3353 (N_3353,N_3196,N_3063);
or U3354 (N_3354,N_3133,N_3075);
or U3355 (N_3355,N_3153,N_3013);
or U3356 (N_3356,N_3034,N_3194);
nor U3357 (N_3357,N_3047,N_3149);
nand U3358 (N_3358,N_3033,N_3028);
nand U3359 (N_3359,N_3097,N_3095);
or U3360 (N_3360,N_3069,N_3097);
or U3361 (N_3361,N_3074,N_3027);
or U3362 (N_3362,N_3169,N_3183);
nand U3363 (N_3363,N_3181,N_3156);
nand U3364 (N_3364,N_3083,N_3060);
nand U3365 (N_3365,N_3145,N_3030);
nor U3366 (N_3366,N_3186,N_3124);
or U3367 (N_3367,N_3105,N_3123);
nor U3368 (N_3368,N_3106,N_3029);
nor U3369 (N_3369,N_3087,N_3069);
and U3370 (N_3370,N_3034,N_3068);
nand U3371 (N_3371,N_3113,N_3169);
nand U3372 (N_3372,N_3071,N_3113);
nand U3373 (N_3373,N_3019,N_3133);
or U3374 (N_3374,N_3175,N_3031);
nor U3375 (N_3375,N_3041,N_3015);
nand U3376 (N_3376,N_3064,N_3103);
nor U3377 (N_3377,N_3077,N_3140);
and U3378 (N_3378,N_3193,N_3108);
or U3379 (N_3379,N_3081,N_3154);
or U3380 (N_3380,N_3183,N_3140);
and U3381 (N_3381,N_3198,N_3182);
and U3382 (N_3382,N_3163,N_3076);
or U3383 (N_3383,N_3099,N_3159);
or U3384 (N_3384,N_3087,N_3198);
nor U3385 (N_3385,N_3031,N_3034);
and U3386 (N_3386,N_3168,N_3113);
nor U3387 (N_3387,N_3192,N_3037);
nand U3388 (N_3388,N_3093,N_3158);
and U3389 (N_3389,N_3179,N_3116);
nand U3390 (N_3390,N_3165,N_3142);
nand U3391 (N_3391,N_3094,N_3029);
nand U3392 (N_3392,N_3123,N_3026);
and U3393 (N_3393,N_3118,N_3142);
and U3394 (N_3394,N_3178,N_3107);
nor U3395 (N_3395,N_3112,N_3157);
nor U3396 (N_3396,N_3084,N_3133);
nor U3397 (N_3397,N_3075,N_3183);
nor U3398 (N_3398,N_3123,N_3126);
nor U3399 (N_3399,N_3178,N_3071);
or U3400 (N_3400,N_3290,N_3244);
nand U3401 (N_3401,N_3383,N_3210);
nor U3402 (N_3402,N_3232,N_3295);
nor U3403 (N_3403,N_3289,N_3321);
nand U3404 (N_3404,N_3281,N_3360);
nor U3405 (N_3405,N_3307,N_3315);
or U3406 (N_3406,N_3283,N_3390);
nor U3407 (N_3407,N_3313,N_3312);
or U3408 (N_3408,N_3309,N_3242);
nor U3409 (N_3409,N_3240,N_3393);
nor U3410 (N_3410,N_3279,N_3341);
and U3411 (N_3411,N_3363,N_3247);
or U3412 (N_3412,N_3357,N_3369);
nor U3413 (N_3413,N_3370,N_3226);
and U3414 (N_3414,N_3231,N_3397);
nand U3415 (N_3415,N_3392,N_3284);
nor U3416 (N_3416,N_3345,N_3213);
nor U3417 (N_3417,N_3338,N_3396);
or U3418 (N_3418,N_3320,N_3288);
and U3419 (N_3419,N_3361,N_3253);
nor U3420 (N_3420,N_3222,N_3300);
or U3421 (N_3421,N_3229,N_3344);
or U3422 (N_3422,N_3218,N_3330);
nor U3423 (N_3423,N_3276,N_3319);
and U3424 (N_3424,N_3327,N_3260);
nand U3425 (N_3425,N_3381,N_3372);
or U3426 (N_3426,N_3323,N_3375);
or U3427 (N_3427,N_3332,N_3227);
and U3428 (N_3428,N_3267,N_3326);
nor U3429 (N_3429,N_3265,N_3202);
nand U3430 (N_3430,N_3365,N_3395);
nand U3431 (N_3431,N_3234,N_3301);
nor U3432 (N_3432,N_3349,N_3249);
and U3433 (N_3433,N_3324,N_3264);
and U3434 (N_3434,N_3259,N_3251);
nand U3435 (N_3435,N_3306,N_3386);
nand U3436 (N_3436,N_3316,N_3200);
and U3437 (N_3437,N_3248,N_3358);
and U3438 (N_3438,N_3245,N_3205);
nor U3439 (N_3439,N_3353,N_3355);
nand U3440 (N_3440,N_3388,N_3209);
nor U3441 (N_3441,N_3230,N_3286);
nor U3442 (N_3442,N_3238,N_3262);
or U3443 (N_3443,N_3376,N_3221);
or U3444 (N_3444,N_3246,N_3346);
nand U3445 (N_3445,N_3356,N_3257);
or U3446 (N_3446,N_3261,N_3255);
or U3447 (N_3447,N_3371,N_3206);
and U3448 (N_3448,N_3329,N_3366);
and U3449 (N_3449,N_3252,N_3325);
and U3450 (N_3450,N_3351,N_3278);
and U3451 (N_3451,N_3239,N_3219);
or U3452 (N_3452,N_3215,N_3380);
or U3453 (N_3453,N_3367,N_3354);
nand U3454 (N_3454,N_3272,N_3394);
or U3455 (N_3455,N_3243,N_3382);
and U3456 (N_3456,N_3333,N_3352);
nor U3457 (N_3457,N_3378,N_3308);
and U3458 (N_3458,N_3311,N_3362);
nand U3459 (N_3459,N_3317,N_3336);
or U3460 (N_3460,N_3391,N_3223);
nor U3461 (N_3461,N_3368,N_3297);
nor U3462 (N_3462,N_3379,N_3292);
nor U3463 (N_3463,N_3377,N_3233);
and U3464 (N_3464,N_3337,N_3373);
nor U3465 (N_3465,N_3214,N_3269);
and U3466 (N_3466,N_3225,N_3224);
and U3467 (N_3467,N_3280,N_3294);
nor U3468 (N_3468,N_3347,N_3266);
or U3469 (N_3469,N_3364,N_3303);
nand U3470 (N_3470,N_3298,N_3340);
nand U3471 (N_3471,N_3216,N_3212);
nor U3472 (N_3472,N_3254,N_3302);
or U3473 (N_3473,N_3314,N_3350);
and U3474 (N_3474,N_3207,N_3228);
and U3475 (N_3475,N_3237,N_3334);
or U3476 (N_3476,N_3387,N_3305);
or U3477 (N_3477,N_3322,N_3287);
nor U3478 (N_3478,N_3299,N_3291);
nor U3479 (N_3479,N_3256,N_3250);
nand U3480 (N_3480,N_3385,N_3270);
nand U3481 (N_3481,N_3201,N_3359);
and U3482 (N_3482,N_3268,N_3236);
and U3483 (N_3483,N_3217,N_3273);
and U3484 (N_3484,N_3235,N_3282);
and U3485 (N_3485,N_3374,N_3389);
nand U3486 (N_3486,N_3296,N_3211);
nor U3487 (N_3487,N_3220,N_3293);
nor U3488 (N_3488,N_3274,N_3241);
and U3489 (N_3489,N_3339,N_3277);
xnor U3490 (N_3490,N_3343,N_3271);
nand U3491 (N_3491,N_3304,N_3342);
or U3492 (N_3492,N_3203,N_3328);
or U3493 (N_3493,N_3318,N_3258);
or U3494 (N_3494,N_3335,N_3399);
and U3495 (N_3495,N_3398,N_3204);
nand U3496 (N_3496,N_3263,N_3310);
and U3497 (N_3497,N_3331,N_3348);
and U3498 (N_3498,N_3384,N_3285);
nor U3499 (N_3499,N_3275,N_3208);
or U3500 (N_3500,N_3200,N_3216);
and U3501 (N_3501,N_3379,N_3357);
and U3502 (N_3502,N_3264,N_3369);
nand U3503 (N_3503,N_3319,N_3354);
nor U3504 (N_3504,N_3359,N_3378);
and U3505 (N_3505,N_3309,N_3201);
nor U3506 (N_3506,N_3285,N_3317);
nand U3507 (N_3507,N_3308,N_3271);
nand U3508 (N_3508,N_3320,N_3337);
and U3509 (N_3509,N_3248,N_3329);
nand U3510 (N_3510,N_3341,N_3348);
nor U3511 (N_3511,N_3295,N_3334);
and U3512 (N_3512,N_3278,N_3293);
and U3513 (N_3513,N_3207,N_3209);
nand U3514 (N_3514,N_3398,N_3225);
and U3515 (N_3515,N_3392,N_3389);
nand U3516 (N_3516,N_3228,N_3351);
nand U3517 (N_3517,N_3395,N_3356);
nor U3518 (N_3518,N_3395,N_3344);
nor U3519 (N_3519,N_3322,N_3378);
and U3520 (N_3520,N_3242,N_3255);
or U3521 (N_3521,N_3377,N_3372);
or U3522 (N_3522,N_3230,N_3214);
nor U3523 (N_3523,N_3327,N_3285);
nor U3524 (N_3524,N_3362,N_3236);
and U3525 (N_3525,N_3214,N_3260);
or U3526 (N_3526,N_3254,N_3207);
and U3527 (N_3527,N_3312,N_3367);
and U3528 (N_3528,N_3369,N_3337);
nand U3529 (N_3529,N_3348,N_3384);
nand U3530 (N_3530,N_3394,N_3371);
xnor U3531 (N_3531,N_3383,N_3220);
and U3532 (N_3532,N_3264,N_3329);
and U3533 (N_3533,N_3212,N_3299);
nand U3534 (N_3534,N_3286,N_3345);
nor U3535 (N_3535,N_3362,N_3336);
or U3536 (N_3536,N_3380,N_3396);
nand U3537 (N_3537,N_3209,N_3369);
nor U3538 (N_3538,N_3228,N_3214);
nand U3539 (N_3539,N_3326,N_3281);
nor U3540 (N_3540,N_3316,N_3263);
or U3541 (N_3541,N_3333,N_3224);
or U3542 (N_3542,N_3321,N_3346);
nand U3543 (N_3543,N_3378,N_3202);
nor U3544 (N_3544,N_3336,N_3208);
or U3545 (N_3545,N_3260,N_3352);
and U3546 (N_3546,N_3303,N_3311);
nand U3547 (N_3547,N_3209,N_3260);
nand U3548 (N_3548,N_3225,N_3329);
nor U3549 (N_3549,N_3300,N_3372);
and U3550 (N_3550,N_3332,N_3270);
nand U3551 (N_3551,N_3250,N_3317);
and U3552 (N_3552,N_3320,N_3278);
nand U3553 (N_3553,N_3297,N_3385);
or U3554 (N_3554,N_3303,N_3366);
and U3555 (N_3555,N_3293,N_3269);
nand U3556 (N_3556,N_3363,N_3326);
nor U3557 (N_3557,N_3233,N_3288);
xor U3558 (N_3558,N_3298,N_3369);
and U3559 (N_3559,N_3206,N_3281);
nor U3560 (N_3560,N_3246,N_3315);
and U3561 (N_3561,N_3298,N_3237);
nor U3562 (N_3562,N_3385,N_3283);
nand U3563 (N_3563,N_3353,N_3206);
or U3564 (N_3564,N_3348,N_3346);
and U3565 (N_3565,N_3261,N_3323);
nand U3566 (N_3566,N_3315,N_3317);
nor U3567 (N_3567,N_3263,N_3393);
nand U3568 (N_3568,N_3308,N_3241);
xor U3569 (N_3569,N_3328,N_3362);
xnor U3570 (N_3570,N_3367,N_3207);
or U3571 (N_3571,N_3367,N_3336);
nand U3572 (N_3572,N_3377,N_3283);
and U3573 (N_3573,N_3378,N_3262);
nand U3574 (N_3574,N_3373,N_3293);
and U3575 (N_3575,N_3218,N_3221);
nand U3576 (N_3576,N_3322,N_3369);
nand U3577 (N_3577,N_3214,N_3273);
nand U3578 (N_3578,N_3237,N_3266);
nand U3579 (N_3579,N_3209,N_3341);
or U3580 (N_3580,N_3343,N_3388);
nor U3581 (N_3581,N_3350,N_3373);
and U3582 (N_3582,N_3238,N_3201);
nor U3583 (N_3583,N_3317,N_3223);
or U3584 (N_3584,N_3398,N_3251);
or U3585 (N_3585,N_3304,N_3200);
or U3586 (N_3586,N_3314,N_3381);
nand U3587 (N_3587,N_3282,N_3304);
or U3588 (N_3588,N_3277,N_3354);
nand U3589 (N_3589,N_3235,N_3365);
or U3590 (N_3590,N_3206,N_3266);
nand U3591 (N_3591,N_3290,N_3370);
or U3592 (N_3592,N_3385,N_3242);
nand U3593 (N_3593,N_3210,N_3203);
nor U3594 (N_3594,N_3269,N_3371);
and U3595 (N_3595,N_3393,N_3377);
and U3596 (N_3596,N_3394,N_3310);
or U3597 (N_3597,N_3357,N_3310);
or U3598 (N_3598,N_3349,N_3257);
nand U3599 (N_3599,N_3259,N_3370);
nand U3600 (N_3600,N_3487,N_3545);
or U3601 (N_3601,N_3510,N_3596);
and U3602 (N_3602,N_3404,N_3467);
nand U3603 (N_3603,N_3482,N_3594);
or U3604 (N_3604,N_3416,N_3598);
nor U3605 (N_3605,N_3518,N_3400);
nand U3606 (N_3606,N_3529,N_3507);
nand U3607 (N_3607,N_3523,N_3429);
nand U3608 (N_3608,N_3484,N_3458);
nand U3609 (N_3609,N_3468,N_3474);
nor U3610 (N_3610,N_3494,N_3436);
nand U3611 (N_3611,N_3502,N_3514);
and U3612 (N_3612,N_3534,N_3528);
or U3613 (N_3613,N_3562,N_3493);
or U3614 (N_3614,N_3541,N_3411);
and U3615 (N_3615,N_3491,N_3505);
nand U3616 (N_3616,N_3587,N_3441);
and U3617 (N_3617,N_3439,N_3437);
and U3618 (N_3618,N_3585,N_3572);
nand U3619 (N_3619,N_3595,N_3536);
or U3620 (N_3620,N_3576,N_3427);
and U3621 (N_3621,N_3535,N_3470);
or U3622 (N_3622,N_3466,N_3559);
nand U3623 (N_3623,N_3471,N_3461);
and U3624 (N_3624,N_3420,N_3425);
nor U3625 (N_3625,N_3492,N_3503);
and U3626 (N_3626,N_3408,N_3443);
nor U3627 (N_3627,N_3430,N_3453);
or U3628 (N_3628,N_3463,N_3549);
and U3629 (N_3629,N_3574,N_3433);
and U3630 (N_3630,N_3477,N_3563);
or U3631 (N_3631,N_3588,N_3511);
or U3632 (N_3632,N_3557,N_3578);
nor U3633 (N_3633,N_3583,N_3584);
nand U3634 (N_3634,N_3449,N_3516);
nor U3635 (N_3635,N_3517,N_3451);
or U3636 (N_3636,N_3465,N_3531);
or U3637 (N_3637,N_3550,N_3409);
nor U3638 (N_3638,N_3490,N_3472);
nor U3639 (N_3639,N_3519,N_3406);
nor U3640 (N_3640,N_3582,N_3459);
nand U3641 (N_3641,N_3464,N_3570);
or U3642 (N_3642,N_3543,N_3560);
nor U3643 (N_3643,N_3489,N_3552);
and U3644 (N_3644,N_3575,N_3448);
nand U3645 (N_3645,N_3533,N_3548);
nor U3646 (N_3646,N_3546,N_3593);
nor U3647 (N_3647,N_3539,N_3540);
or U3648 (N_3648,N_3415,N_3520);
nand U3649 (N_3649,N_3592,N_3499);
nor U3650 (N_3650,N_3456,N_3551);
or U3651 (N_3651,N_3410,N_3506);
nor U3652 (N_3652,N_3526,N_3555);
and U3653 (N_3653,N_3403,N_3530);
or U3654 (N_3654,N_3424,N_3554);
nor U3655 (N_3655,N_3579,N_3571);
nand U3656 (N_3656,N_3475,N_3504);
or U3657 (N_3657,N_3591,N_3401);
xnor U3658 (N_3658,N_3573,N_3479);
nor U3659 (N_3659,N_3417,N_3407);
nand U3660 (N_3660,N_3564,N_3515);
nand U3661 (N_3661,N_3547,N_3447);
and U3662 (N_3662,N_3444,N_3485);
nand U3663 (N_3663,N_3561,N_3438);
or U3664 (N_3664,N_3455,N_3590);
nand U3665 (N_3665,N_3422,N_3597);
nor U3666 (N_3666,N_3426,N_3446);
and U3667 (N_3667,N_3412,N_3542);
or U3668 (N_3668,N_3580,N_3501);
or U3669 (N_3669,N_3440,N_3421);
or U3670 (N_3670,N_3532,N_3513);
nor U3671 (N_3671,N_3432,N_3498);
nand U3672 (N_3672,N_3556,N_3431);
and U3673 (N_3673,N_3577,N_3473);
nor U3674 (N_3674,N_3405,N_3457);
nand U3675 (N_3675,N_3599,N_3460);
xnor U3676 (N_3676,N_3525,N_3483);
nor U3677 (N_3677,N_3462,N_3414);
or U3678 (N_3678,N_3586,N_3445);
nand U3679 (N_3679,N_3434,N_3589);
and U3680 (N_3680,N_3537,N_3428);
and U3681 (N_3681,N_3419,N_3480);
nand U3682 (N_3682,N_3538,N_3486);
and U3683 (N_3683,N_3478,N_3413);
or U3684 (N_3684,N_3509,N_3527);
nor U3685 (N_3685,N_3558,N_3423);
or U3686 (N_3686,N_3469,N_3508);
and U3687 (N_3687,N_3418,N_3450);
and U3688 (N_3688,N_3442,N_3402);
and U3689 (N_3689,N_3497,N_3569);
nor U3690 (N_3690,N_3581,N_3496);
or U3691 (N_3691,N_3512,N_3553);
nor U3692 (N_3692,N_3476,N_3565);
nor U3693 (N_3693,N_3522,N_3495);
and U3694 (N_3694,N_3567,N_3481);
and U3695 (N_3695,N_3452,N_3454);
and U3696 (N_3696,N_3500,N_3566);
nand U3697 (N_3697,N_3521,N_3544);
or U3698 (N_3698,N_3568,N_3524);
nor U3699 (N_3699,N_3435,N_3488);
or U3700 (N_3700,N_3558,N_3428);
or U3701 (N_3701,N_3463,N_3456);
or U3702 (N_3702,N_3531,N_3500);
or U3703 (N_3703,N_3463,N_3478);
nor U3704 (N_3704,N_3581,N_3535);
nor U3705 (N_3705,N_3591,N_3441);
nor U3706 (N_3706,N_3482,N_3564);
xnor U3707 (N_3707,N_3420,N_3441);
and U3708 (N_3708,N_3418,N_3507);
or U3709 (N_3709,N_3421,N_3543);
nand U3710 (N_3710,N_3452,N_3526);
nor U3711 (N_3711,N_3468,N_3571);
or U3712 (N_3712,N_3473,N_3429);
xnor U3713 (N_3713,N_3433,N_3428);
and U3714 (N_3714,N_3486,N_3441);
nor U3715 (N_3715,N_3534,N_3524);
nand U3716 (N_3716,N_3464,N_3581);
or U3717 (N_3717,N_3531,N_3576);
nor U3718 (N_3718,N_3493,N_3468);
nand U3719 (N_3719,N_3468,N_3401);
nand U3720 (N_3720,N_3402,N_3436);
nand U3721 (N_3721,N_3487,N_3573);
nor U3722 (N_3722,N_3548,N_3504);
nor U3723 (N_3723,N_3547,N_3526);
nand U3724 (N_3724,N_3467,N_3424);
or U3725 (N_3725,N_3487,N_3501);
nor U3726 (N_3726,N_3449,N_3481);
or U3727 (N_3727,N_3538,N_3593);
and U3728 (N_3728,N_3446,N_3453);
nor U3729 (N_3729,N_3418,N_3516);
nand U3730 (N_3730,N_3514,N_3557);
nand U3731 (N_3731,N_3501,N_3521);
or U3732 (N_3732,N_3590,N_3475);
nand U3733 (N_3733,N_3579,N_3480);
and U3734 (N_3734,N_3487,N_3590);
or U3735 (N_3735,N_3410,N_3542);
and U3736 (N_3736,N_3481,N_3548);
and U3737 (N_3737,N_3521,N_3480);
and U3738 (N_3738,N_3522,N_3481);
xor U3739 (N_3739,N_3467,N_3497);
or U3740 (N_3740,N_3504,N_3505);
nand U3741 (N_3741,N_3425,N_3435);
and U3742 (N_3742,N_3453,N_3500);
and U3743 (N_3743,N_3579,N_3482);
or U3744 (N_3744,N_3498,N_3478);
nand U3745 (N_3745,N_3543,N_3569);
or U3746 (N_3746,N_3426,N_3435);
or U3747 (N_3747,N_3532,N_3470);
or U3748 (N_3748,N_3545,N_3538);
and U3749 (N_3749,N_3552,N_3569);
or U3750 (N_3750,N_3540,N_3439);
or U3751 (N_3751,N_3489,N_3424);
and U3752 (N_3752,N_3424,N_3529);
nor U3753 (N_3753,N_3452,N_3546);
nand U3754 (N_3754,N_3535,N_3421);
and U3755 (N_3755,N_3557,N_3458);
nand U3756 (N_3756,N_3463,N_3568);
nand U3757 (N_3757,N_3457,N_3487);
nand U3758 (N_3758,N_3440,N_3431);
nand U3759 (N_3759,N_3568,N_3474);
nor U3760 (N_3760,N_3555,N_3590);
xor U3761 (N_3761,N_3572,N_3423);
nand U3762 (N_3762,N_3426,N_3535);
or U3763 (N_3763,N_3556,N_3543);
nor U3764 (N_3764,N_3520,N_3593);
and U3765 (N_3765,N_3410,N_3413);
nand U3766 (N_3766,N_3439,N_3421);
nand U3767 (N_3767,N_3576,N_3597);
nor U3768 (N_3768,N_3458,N_3540);
or U3769 (N_3769,N_3411,N_3452);
and U3770 (N_3770,N_3509,N_3405);
or U3771 (N_3771,N_3574,N_3521);
or U3772 (N_3772,N_3435,N_3438);
nor U3773 (N_3773,N_3477,N_3571);
and U3774 (N_3774,N_3528,N_3412);
and U3775 (N_3775,N_3510,N_3546);
nand U3776 (N_3776,N_3438,N_3566);
or U3777 (N_3777,N_3518,N_3495);
nor U3778 (N_3778,N_3573,N_3502);
nor U3779 (N_3779,N_3409,N_3406);
or U3780 (N_3780,N_3586,N_3599);
nand U3781 (N_3781,N_3542,N_3547);
or U3782 (N_3782,N_3523,N_3587);
nand U3783 (N_3783,N_3521,N_3539);
nor U3784 (N_3784,N_3438,N_3449);
or U3785 (N_3785,N_3443,N_3564);
nor U3786 (N_3786,N_3506,N_3488);
or U3787 (N_3787,N_3419,N_3534);
or U3788 (N_3788,N_3437,N_3457);
and U3789 (N_3789,N_3546,N_3431);
or U3790 (N_3790,N_3453,N_3452);
or U3791 (N_3791,N_3495,N_3418);
or U3792 (N_3792,N_3508,N_3495);
nand U3793 (N_3793,N_3413,N_3488);
nor U3794 (N_3794,N_3581,N_3467);
nor U3795 (N_3795,N_3572,N_3530);
or U3796 (N_3796,N_3420,N_3541);
or U3797 (N_3797,N_3499,N_3426);
nand U3798 (N_3798,N_3555,N_3583);
nand U3799 (N_3799,N_3512,N_3487);
nor U3800 (N_3800,N_3693,N_3683);
nor U3801 (N_3801,N_3631,N_3662);
and U3802 (N_3802,N_3624,N_3610);
nor U3803 (N_3803,N_3730,N_3675);
and U3804 (N_3804,N_3770,N_3689);
or U3805 (N_3805,N_3714,N_3760);
nor U3806 (N_3806,N_3703,N_3724);
or U3807 (N_3807,N_3615,N_3665);
nor U3808 (N_3808,N_3772,N_3782);
and U3809 (N_3809,N_3745,N_3698);
or U3810 (N_3810,N_3647,N_3655);
nor U3811 (N_3811,N_3712,N_3781);
nand U3812 (N_3812,N_3713,N_3758);
nand U3813 (N_3813,N_3743,N_3605);
nor U3814 (N_3814,N_3754,N_3696);
or U3815 (N_3815,N_3741,N_3704);
nor U3816 (N_3816,N_3701,N_3729);
and U3817 (N_3817,N_3785,N_3670);
nand U3818 (N_3818,N_3656,N_3674);
or U3819 (N_3819,N_3722,N_3721);
or U3820 (N_3820,N_3669,N_3793);
and U3821 (N_3821,N_3613,N_3723);
nor U3822 (N_3822,N_3755,N_3709);
nand U3823 (N_3823,N_3769,N_3620);
nor U3824 (N_3824,N_3606,N_3695);
nor U3825 (N_3825,N_3671,N_3614);
or U3826 (N_3826,N_3708,N_3632);
nand U3827 (N_3827,N_3638,N_3688);
and U3828 (N_3828,N_3641,N_3750);
nor U3829 (N_3829,N_3654,N_3679);
nand U3830 (N_3830,N_3667,N_3691);
nand U3831 (N_3831,N_3734,N_3700);
nor U3832 (N_3832,N_3771,N_3681);
nand U3833 (N_3833,N_3759,N_3652);
or U3834 (N_3834,N_3780,N_3775);
or U3835 (N_3835,N_3702,N_3682);
nor U3836 (N_3836,N_3715,N_3797);
and U3837 (N_3837,N_3753,N_3676);
nand U3838 (N_3838,N_3608,N_3643);
and U3839 (N_3839,N_3799,N_3744);
nor U3840 (N_3840,N_3789,N_3672);
nand U3841 (N_3841,N_3707,N_3650);
and U3842 (N_3842,N_3727,N_3751);
nor U3843 (N_3843,N_3765,N_3763);
nand U3844 (N_3844,N_3663,N_3680);
nand U3845 (N_3845,N_3623,N_3711);
or U3846 (N_3846,N_3653,N_3659);
or U3847 (N_3847,N_3749,N_3795);
and U3848 (N_3848,N_3735,N_3746);
nor U3849 (N_3849,N_3686,N_3739);
nor U3850 (N_3850,N_3604,N_3778);
nor U3851 (N_3851,N_3645,N_3777);
or U3852 (N_3852,N_3738,N_3784);
or U3853 (N_3853,N_3621,N_3609);
or U3854 (N_3854,N_3619,N_3661);
and U3855 (N_3855,N_3639,N_3791);
and U3856 (N_3856,N_3612,N_3697);
and U3857 (N_3857,N_3685,N_3786);
nand U3858 (N_3858,N_3756,N_3783);
nand U3859 (N_3859,N_3600,N_3673);
xnor U3860 (N_3860,N_3699,N_3617);
and U3861 (N_3861,N_3690,N_3634);
or U3862 (N_3862,N_3790,N_3625);
or U3863 (N_3863,N_3719,N_3628);
nand U3864 (N_3864,N_3694,N_3635);
or U3865 (N_3865,N_3607,N_3706);
nand U3866 (N_3866,N_3657,N_3716);
nor U3867 (N_3867,N_3792,N_3717);
nand U3868 (N_3868,N_3630,N_3774);
nor U3869 (N_3869,N_3629,N_3787);
nand U3870 (N_3870,N_3768,N_3677);
nor U3871 (N_3871,N_3640,N_3798);
nand U3872 (N_3872,N_3603,N_3788);
and U3873 (N_3873,N_3796,N_3733);
nand U3874 (N_3874,N_3651,N_3710);
nand U3875 (N_3875,N_3705,N_3740);
and U3876 (N_3876,N_3794,N_3761);
and U3877 (N_3877,N_3601,N_3725);
nor U3878 (N_3878,N_3776,N_3736);
and U3879 (N_3879,N_3762,N_3748);
and U3880 (N_3880,N_3637,N_3649);
or U3881 (N_3881,N_3622,N_3752);
and U3882 (N_3882,N_3644,N_3636);
nand U3883 (N_3883,N_3773,N_3618);
nand U3884 (N_3884,N_3767,N_3678);
or U3885 (N_3885,N_3692,N_3660);
and U3886 (N_3886,N_3602,N_3648);
or U3887 (N_3887,N_3642,N_3728);
nor U3888 (N_3888,N_3684,N_3764);
nand U3889 (N_3889,N_3626,N_3668);
or U3890 (N_3890,N_3732,N_3766);
nand U3891 (N_3891,N_3718,N_3779);
or U3892 (N_3892,N_3757,N_3687);
nor U3893 (N_3893,N_3633,N_3747);
xnor U3894 (N_3894,N_3611,N_3737);
or U3895 (N_3895,N_3664,N_3731);
or U3896 (N_3896,N_3742,N_3646);
nand U3897 (N_3897,N_3658,N_3726);
nand U3898 (N_3898,N_3616,N_3666);
nand U3899 (N_3899,N_3627,N_3720);
nand U3900 (N_3900,N_3737,N_3617);
and U3901 (N_3901,N_3713,N_3681);
nor U3902 (N_3902,N_3626,N_3621);
nand U3903 (N_3903,N_3777,N_3745);
and U3904 (N_3904,N_3666,N_3619);
nor U3905 (N_3905,N_3737,N_3604);
nand U3906 (N_3906,N_3637,N_3704);
nand U3907 (N_3907,N_3605,N_3711);
or U3908 (N_3908,N_3620,N_3688);
nor U3909 (N_3909,N_3698,N_3784);
or U3910 (N_3910,N_3633,N_3600);
nor U3911 (N_3911,N_3660,N_3750);
nor U3912 (N_3912,N_3745,N_3755);
or U3913 (N_3913,N_3733,N_3640);
and U3914 (N_3914,N_3761,N_3688);
nor U3915 (N_3915,N_3650,N_3671);
and U3916 (N_3916,N_3693,N_3725);
and U3917 (N_3917,N_3754,N_3665);
or U3918 (N_3918,N_3632,N_3698);
and U3919 (N_3919,N_3647,N_3646);
and U3920 (N_3920,N_3681,N_3754);
nand U3921 (N_3921,N_3745,N_3799);
or U3922 (N_3922,N_3702,N_3625);
or U3923 (N_3923,N_3770,N_3683);
nand U3924 (N_3924,N_3786,N_3728);
nand U3925 (N_3925,N_3744,N_3663);
nand U3926 (N_3926,N_3768,N_3684);
nor U3927 (N_3927,N_3627,N_3747);
or U3928 (N_3928,N_3769,N_3632);
and U3929 (N_3929,N_3671,N_3669);
or U3930 (N_3930,N_3655,N_3728);
nand U3931 (N_3931,N_3670,N_3780);
and U3932 (N_3932,N_3625,N_3676);
nor U3933 (N_3933,N_3750,N_3707);
nor U3934 (N_3934,N_3768,N_3717);
and U3935 (N_3935,N_3657,N_3799);
and U3936 (N_3936,N_3616,N_3748);
or U3937 (N_3937,N_3650,N_3681);
and U3938 (N_3938,N_3711,N_3727);
nand U3939 (N_3939,N_3701,N_3645);
nor U3940 (N_3940,N_3637,N_3746);
and U3941 (N_3941,N_3644,N_3696);
or U3942 (N_3942,N_3701,N_3723);
nor U3943 (N_3943,N_3721,N_3600);
nand U3944 (N_3944,N_3730,N_3775);
nand U3945 (N_3945,N_3795,N_3665);
and U3946 (N_3946,N_3745,N_3649);
or U3947 (N_3947,N_3690,N_3644);
nand U3948 (N_3948,N_3785,N_3772);
nor U3949 (N_3949,N_3784,N_3638);
nor U3950 (N_3950,N_3792,N_3632);
or U3951 (N_3951,N_3656,N_3743);
or U3952 (N_3952,N_3607,N_3745);
and U3953 (N_3953,N_3754,N_3634);
nand U3954 (N_3954,N_3761,N_3749);
nor U3955 (N_3955,N_3758,N_3648);
nor U3956 (N_3956,N_3635,N_3752);
nand U3957 (N_3957,N_3746,N_3744);
nor U3958 (N_3958,N_3760,N_3786);
nand U3959 (N_3959,N_3631,N_3609);
nand U3960 (N_3960,N_3728,N_3777);
nand U3961 (N_3961,N_3672,N_3761);
and U3962 (N_3962,N_3696,N_3726);
nor U3963 (N_3963,N_3618,N_3617);
or U3964 (N_3964,N_3631,N_3693);
or U3965 (N_3965,N_3659,N_3615);
nand U3966 (N_3966,N_3692,N_3629);
nor U3967 (N_3967,N_3664,N_3682);
nand U3968 (N_3968,N_3680,N_3622);
nand U3969 (N_3969,N_3706,N_3686);
and U3970 (N_3970,N_3607,N_3771);
nand U3971 (N_3971,N_3676,N_3666);
and U3972 (N_3972,N_3660,N_3728);
and U3973 (N_3973,N_3622,N_3797);
and U3974 (N_3974,N_3796,N_3636);
or U3975 (N_3975,N_3677,N_3641);
nand U3976 (N_3976,N_3717,N_3709);
nand U3977 (N_3977,N_3720,N_3761);
nand U3978 (N_3978,N_3646,N_3613);
or U3979 (N_3979,N_3775,N_3751);
nand U3980 (N_3980,N_3673,N_3784);
or U3981 (N_3981,N_3777,N_3604);
nand U3982 (N_3982,N_3603,N_3797);
and U3983 (N_3983,N_3652,N_3623);
nor U3984 (N_3984,N_3628,N_3737);
or U3985 (N_3985,N_3728,N_3755);
nor U3986 (N_3986,N_3753,N_3600);
nor U3987 (N_3987,N_3772,N_3685);
and U3988 (N_3988,N_3703,N_3714);
and U3989 (N_3989,N_3658,N_3643);
nand U3990 (N_3990,N_3681,N_3699);
or U3991 (N_3991,N_3602,N_3702);
nor U3992 (N_3992,N_3726,N_3723);
and U3993 (N_3993,N_3741,N_3793);
nand U3994 (N_3994,N_3759,N_3783);
or U3995 (N_3995,N_3639,N_3696);
or U3996 (N_3996,N_3735,N_3662);
nor U3997 (N_3997,N_3760,N_3737);
or U3998 (N_3998,N_3624,N_3679);
nand U3999 (N_3999,N_3615,N_3755);
and U4000 (N_4000,N_3965,N_3976);
and U4001 (N_4001,N_3810,N_3925);
nor U4002 (N_4002,N_3885,N_3975);
nand U4003 (N_4003,N_3846,N_3871);
or U4004 (N_4004,N_3926,N_3806);
and U4005 (N_4005,N_3948,N_3977);
or U4006 (N_4006,N_3942,N_3919);
nor U4007 (N_4007,N_3999,N_3936);
or U4008 (N_4008,N_3863,N_3868);
nor U4009 (N_4009,N_3876,N_3913);
nor U4010 (N_4010,N_3865,N_3823);
and U4011 (N_4011,N_3809,N_3923);
or U4012 (N_4012,N_3990,N_3860);
and U4013 (N_4013,N_3934,N_3896);
and U4014 (N_4014,N_3981,N_3829);
and U4015 (N_4015,N_3931,N_3830);
or U4016 (N_4016,N_3803,N_3912);
or U4017 (N_4017,N_3992,N_3964);
nor U4018 (N_4018,N_3812,N_3894);
nand U4019 (N_4019,N_3997,N_3956);
and U4020 (N_4020,N_3859,N_3927);
nand U4021 (N_4021,N_3850,N_3849);
or U4022 (N_4022,N_3881,N_3983);
nor U4023 (N_4023,N_3935,N_3838);
and U4024 (N_4024,N_3945,N_3840);
or U4025 (N_4025,N_3958,N_3819);
xor U4026 (N_4026,N_3902,N_3946);
nor U4027 (N_4027,N_3968,N_3973);
nor U4028 (N_4028,N_3834,N_3938);
and U4029 (N_4029,N_3899,N_3933);
nand U4030 (N_4030,N_3993,N_3982);
and U4031 (N_4031,N_3879,N_3842);
and U4032 (N_4032,N_3832,N_3855);
and U4033 (N_4033,N_3893,N_3886);
nand U4034 (N_4034,N_3955,N_3906);
or U4035 (N_4035,N_3874,N_3970);
or U4036 (N_4036,N_3873,N_3937);
nor U4037 (N_4037,N_3811,N_3959);
nand U4038 (N_4038,N_3820,N_3870);
and U4039 (N_4039,N_3862,N_3943);
and U4040 (N_4040,N_3867,N_3817);
nand U4041 (N_4041,N_3816,N_3883);
or U4042 (N_4042,N_3951,N_3911);
nor U4043 (N_4043,N_3984,N_3839);
nor U4044 (N_4044,N_3844,N_3978);
or U4045 (N_4045,N_3875,N_3947);
nor U4046 (N_4046,N_3954,N_3872);
or U4047 (N_4047,N_3905,N_3808);
nor U4048 (N_4048,N_3805,N_3914);
nor U4049 (N_4049,N_3944,N_3857);
or U4050 (N_4050,N_3833,N_3949);
nand U4051 (N_4051,N_3891,N_3920);
nor U4052 (N_4052,N_3827,N_3826);
nand U4053 (N_4053,N_3845,N_3898);
or U4054 (N_4054,N_3831,N_3979);
and U4055 (N_4055,N_3847,N_3996);
nand U4056 (N_4056,N_3835,N_3961);
nor U4057 (N_4057,N_3966,N_3910);
nor U4058 (N_4058,N_3929,N_3957);
nor U4059 (N_4059,N_3841,N_3916);
nor U4060 (N_4060,N_3971,N_3907);
and U4061 (N_4061,N_3995,N_3864);
and U4062 (N_4062,N_3908,N_3904);
nand U4063 (N_4063,N_3807,N_3989);
nand U4064 (N_4064,N_3918,N_3960);
nand U4065 (N_4065,N_3852,N_3941);
nand U4066 (N_4066,N_3939,N_3821);
or U4067 (N_4067,N_3962,N_3887);
or U4068 (N_4068,N_3998,N_3822);
nand U4069 (N_4069,N_3878,N_3980);
and U4070 (N_4070,N_3917,N_3856);
nand U4071 (N_4071,N_3988,N_3837);
nand U4072 (N_4072,N_3861,N_3928);
nor U4073 (N_4073,N_3915,N_3900);
nor U4074 (N_4074,N_3877,N_3854);
and U4075 (N_4075,N_3986,N_3880);
nor U4076 (N_4076,N_3932,N_3818);
and U4077 (N_4077,N_3866,N_3825);
or U4078 (N_4078,N_3967,N_3952);
nand U4079 (N_4079,N_3801,N_3969);
nor U4080 (N_4080,N_3824,N_3953);
and U4081 (N_4081,N_3882,N_3987);
or U4082 (N_4082,N_3853,N_3909);
or U4083 (N_4083,N_3994,N_3889);
and U4084 (N_4084,N_3815,N_3922);
nand U4085 (N_4085,N_3991,N_3804);
nor U4086 (N_4086,N_3890,N_3985);
and U4087 (N_4087,N_3930,N_3950);
nor U4088 (N_4088,N_3924,N_3921);
and U4089 (N_4089,N_3802,N_3843);
and U4090 (N_4090,N_3800,N_3851);
nor U4091 (N_4091,N_3828,N_3901);
or U4092 (N_4092,N_3888,N_3814);
nand U4093 (N_4093,N_3897,N_3940);
or U4094 (N_4094,N_3869,N_3903);
or U4095 (N_4095,N_3813,N_3848);
and U4096 (N_4096,N_3858,N_3836);
or U4097 (N_4097,N_3892,N_3974);
and U4098 (N_4098,N_3884,N_3895);
nor U4099 (N_4099,N_3963,N_3972);
nor U4100 (N_4100,N_3853,N_3898);
nor U4101 (N_4101,N_3855,N_3968);
and U4102 (N_4102,N_3814,N_3869);
or U4103 (N_4103,N_3928,N_3887);
xnor U4104 (N_4104,N_3824,N_3850);
or U4105 (N_4105,N_3937,N_3993);
and U4106 (N_4106,N_3921,N_3803);
and U4107 (N_4107,N_3853,N_3907);
and U4108 (N_4108,N_3953,N_3858);
nand U4109 (N_4109,N_3883,N_3971);
nand U4110 (N_4110,N_3825,N_3801);
or U4111 (N_4111,N_3917,N_3833);
or U4112 (N_4112,N_3827,N_3911);
and U4113 (N_4113,N_3857,N_3949);
nand U4114 (N_4114,N_3973,N_3872);
nand U4115 (N_4115,N_3836,N_3888);
nor U4116 (N_4116,N_3940,N_3961);
nand U4117 (N_4117,N_3817,N_3806);
and U4118 (N_4118,N_3852,N_3928);
or U4119 (N_4119,N_3921,N_3995);
and U4120 (N_4120,N_3970,N_3950);
nand U4121 (N_4121,N_3993,N_3954);
and U4122 (N_4122,N_3914,N_3843);
and U4123 (N_4123,N_3805,N_3899);
and U4124 (N_4124,N_3967,N_3981);
nand U4125 (N_4125,N_3875,N_3852);
nand U4126 (N_4126,N_3870,N_3896);
nor U4127 (N_4127,N_3964,N_3837);
nor U4128 (N_4128,N_3819,N_3957);
or U4129 (N_4129,N_3852,N_3817);
nand U4130 (N_4130,N_3877,N_3907);
nor U4131 (N_4131,N_3822,N_3886);
nor U4132 (N_4132,N_3849,N_3816);
and U4133 (N_4133,N_3859,N_3969);
nand U4134 (N_4134,N_3903,N_3807);
nand U4135 (N_4135,N_3996,N_3804);
and U4136 (N_4136,N_3990,N_3985);
nor U4137 (N_4137,N_3921,N_3936);
and U4138 (N_4138,N_3971,N_3972);
and U4139 (N_4139,N_3896,N_3811);
nand U4140 (N_4140,N_3962,N_3827);
and U4141 (N_4141,N_3928,N_3998);
and U4142 (N_4142,N_3856,N_3973);
nor U4143 (N_4143,N_3934,N_3823);
or U4144 (N_4144,N_3983,N_3982);
and U4145 (N_4145,N_3957,N_3831);
nor U4146 (N_4146,N_3893,N_3828);
xor U4147 (N_4147,N_3976,N_3868);
nand U4148 (N_4148,N_3843,N_3883);
and U4149 (N_4149,N_3976,N_3834);
and U4150 (N_4150,N_3929,N_3926);
and U4151 (N_4151,N_3885,N_3932);
and U4152 (N_4152,N_3812,N_3915);
nor U4153 (N_4153,N_3888,N_3952);
nand U4154 (N_4154,N_3827,N_3867);
or U4155 (N_4155,N_3863,N_3846);
nor U4156 (N_4156,N_3975,N_3966);
nor U4157 (N_4157,N_3801,N_3840);
and U4158 (N_4158,N_3868,N_3950);
or U4159 (N_4159,N_3812,N_3861);
and U4160 (N_4160,N_3881,N_3853);
nor U4161 (N_4161,N_3855,N_3931);
nand U4162 (N_4162,N_3890,N_3996);
or U4163 (N_4163,N_3899,N_3908);
nor U4164 (N_4164,N_3939,N_3835);
nor U4165 (N_4165,N_3873,N_3868);
and U4166 (N_4166,N_3982,N_3864);
or U4167 (N_4167,N_3804,N_3941);
or U4168 (N_4168,N_3885,N_3833);
nand U4169 (N_4169,N_3978,N_3955);
or U4170 (N_4170,N_3857,N_3853);
or U4171 (N_4171,N_3892,N_3871);
nand U4172 (N_4172,N_3960,N_3895);
and U4173 (N_4173,N_3929,N_3913);
nand U4174 (N_4174,N_3857,N_3958);
nand U4175 (N_4175,N_3879,N_3961);
or U4176 (N_4176,N_3962,N_3803);
and U4177 (N_4177,N_3959,N_3997);
and U4178 (N_4178,N_3842,N_3838);
nand U4179 (N_4179,N_3914,N_3817);
nor U4180 (N_4180,N_3856,N_3869);
or U4181 (N_4181,N_3804,N_3832);
or U4182 (N_4182,N_3867,N_3957);
nand U4183 (N_4183,N_3943,N_3947);
or U4184 (N_4184,N_3951,N_3804);
and U4185 (N_4185,N_3919,N_3866);
nand U4186 (N_4186,N_3850,N_3865);
or U4187 (N_4187,N_3980,N_3972);
nor U4188 (N_4188,N_3838,N_3971);
nor U4189 (N_4189,N_3992,N_3966);
or U4190 (N_4190,N_3820,N_3837);
or U4191 (N_4191,N_3977,N_3993);
nand U4192 (N_4192,N_3961,N_3978);
and U4193 (N_4193,N_3958,N_3815);
and U4194 (N_4194,N_3832,N_3939);
and U4195 (N_4195,N_3967,N_3927);
or U4196 (N_4196,N_3827,N_3860);
nor U4197 (N_4197,N_3896,N_3807);
nor U4198 (N_4198,N_3973,N_3904);
or U4199 (N_4199,N_3811,N_3802);
nor U4200 (N_4200,N_4089,N_4192);
nand U4201 (N_4201,N_4057,N_4082);
and U4202 (N_4202,N_4079,N_4153);
nor U4203 (N_4203,N_4035,N_4066);
nor U4204 (N_4204,N_4074,N_4036);
nor U4205 (N_4205,N_4008,N_4083);
and U4206 (N_4206,N_4026,N_4034);
nand U4207 (N_4207,N_4168,N_4080);
nor U4208 (N_4208,N_4131,N_4069);
or U4209 (N_4209,N_4110,N_4124);
nand U4210 (N_4210,N_4064,N_4091);
nand U4211 (N_4211,N_4076,N_4187);
nor U4212 (N_4212,N_4135,N_4019);
nor U4213 (N_4213,N_4121,N_4154);
or U4214 (N_4214,N_4052,N_4127);
and U4215 (N_4215,N_4163,N_4198);
nand U4216 (N_4216,N_4123,N_4112);
or U4217 (N_4217,N_4063,N_4177);
nand U4218 (N_4218,N_4119,N_4143);
nand U4219 (N_4219,N_4013,N_4175);
nand U4220 (N_4220,N_4050,N_4094);
or U4221 (N_4221,N_4138,N_4140);
nand U4222 (N_4222,N_4146,N_4166);
nor U4223 (N_4223,N_4020,N_4027);
nand U4224 (N_4224,N_4186,N_4105);
or U4225 (N_4225,N_4157,N_4049);
nand U4226 (N_4226,N_4075,N_4183);
or U4227 (N_4227,N_4058,N_4073);
nor U4228 (N_4228,N_4015,N_4045);
nor U4229 (N_4229,N_4071,N_4059);
or U4230 (N_4230,N_4164,N_4011);
nor U4231 (N_4231,N_4196,N_4185);
nand U4232 (N_4232,N_4150,N_4047);
and U4233 (N_4233,N_4025,N_4044);
and U4234 (N_4234,N_4030,N_4098);
nand U4235 (N_4235,N_4068,N_4055);
nor U4236 (N_4236,N_4014,N_4161);
nor U4237 (N_4237,N_4042,N_4165);
nor U4238 (N_4238,N_4199,N_4130);
nand U4239 (N_4239,N_4088,N_4065);
nor U4240 (N_4240,N_4085,N_4142);
and U4241 (N_4241,N_4111,N_4133);
or U4242 (N_4242,N_4005,N_4113);
nand U4243 (N_4243,N_4132,N_4171);
and U4244 (N_4244,N_4170,N_4017);
nand U4245 (N_4245,N_4197,N_4141);
or U4246 (N_4246,N_4158,N_4033);
and U4247 (N_4247,N_4002,N_4179);
nand U4248 (N_4248,N_4039,N_4077);
nor U4249 (N_4249,N_4120,N_4016);
nand U4250 (N_4250,N_4115,N_4101);
or U4251 (N_4251,N_4003,N_4012);
xor U4252 (N_4252,N_4149,N_4128);
or U4253 (N_4253,N_4028,N_4095);
nor U4254 (N_4254,N_4181,N_4117);
and U4255 (N_4255,N_4087,N_4021);
and U4256 (N_4256,N_4126,N_4061);
or U4257 (N_4257,N_4037,N_4041);
or U4258 (N_4258,N_4040,N_4046);
nand U4259 (N_4259,N_4053,N_4152);
nor U4260 (N_4260,N_4067,N_4189);
nand U4261 (N_4261,N_4102,N_4107);
or U4262 (N_4262,N_4096,N_4148);
nor U4263 (N_4263,N_4029,N_4032);
nor U4264 (N_4264,N_4188,N_4092);
and U4265 (N_4265,N_4001,N_4000);
nor U4266 (N_4266,N_4156,N_4118);
xnor U4267 (N_4267,N_4099,N_4169);
nand U4268 (N_4268,N_4100,N_4056);
nand U4269 (N_4269,N_4178,N_4051);
and U4270 (N_4270,N_4078,N_4172);
and U4271 (N_4271,N_4116,N_4086);
and U4272 (N_4272,N_4160,N_4173);
and U4273 (N_4273,N_4144,N_4125);
nor U4274 (N_4274,N_4176,N_4097);
nand U4275 (N_4275,N_4009,N_4093);
or U4276 (N_4276,N_4109,N_4007);
and U4277 (N_4277,N_4004,N_4180);
nor U4278 (N_4278,N_4054,N_4024);
nor U4279 (N_4279,N_4023,N_4191);
and U4280 (N_4280,N_4129,N_4108);
nor U4281 (N_4281,N_4048,N_4043);
and U4282 (N_4282,N_4010,N_4159);
and U4283 (N_4283,N_4134,N_4145);
or U4284 (N_4284,N_4006,N_4194);
and U4285 (N_4285,N_4137,N_4062);
or U4286 (N_4286,N_4084,N_4155);
nand U4287 (N_4287,N_4122,N_4114);
or U4288 (N_4288,N_4162,N_4167);
nor U4289 (N_4289,N_4060,N_4018);
nand U4290 (N_4290,N_4136,N_4031);
nand U4291 (N_4291,N_4193,N_4104);
nor U4292 (N_4292,N_4184,N_4174);
nor U4293 (N_4293,N_4182,N_4038);
nand U4294 (N_4294,N_4139,N_4090);
nand U4295 (N_4295,N_4106,N_4190);
nand U4296 (N_4296,N_4070,N_4195);
nand U4297 (N_4297,N_4072,N_4103);
or U4298 (N_4298,N_4147,N_4022);
nor U4299 (N_4299,N_4151,N_4081);
and U4300 (N_4300,N_4183,N_4140);
nor U4301 (N_4301,N_4175,N_4082);
nand U4302 (N_4302,N_4182,N_4059);
or U4303 (N_4303,N_4104,N_4145);
nor U4304 (N_4304,N_4074,N_4018);
and U4305 (N_4305,N_4119,N_4052);
xnor U4306 (N_4306,N_4084,N_4175);
nand U4307 (N_4307,N_4145,N_4043);
nand U4308 (N_4308,N_4105,N_4060);
and U4309 (N_4309,N_4050,N_4182);
or U4310 (N_4310,N_4158,N_4197);
and U4311 (N_4311,N_4174,N_4149);
nand U4312 (N_4312,N_4159,N_4185);
and U4313 (N_4313,N_4082,N_4086);
and U4314 (N_4314,N_4095,N_4086);
nor U4315 (N_4315,N_4151,N_4114);
or U4316 (N_4316,N_4027,N_4141);
nor U4317 (N_4317,N_4158,N_4123);
or U4318 (N_4318,N_4091,N_4169);
nor U4319 (N_4319,N_4124,N_4169);
or U4320 (N_4320,N_4122,N_4062);
nor U4321 (N_4321,N_4101,N_4016);
nor U4322 (N_4322,N_4169,N_4017);
nor U4323 (N_4323,N_4131,N_4091);
nor U4324 (N_4324,N_4143,N_4078);
or U4325 (N_4325,N_4191,N_4018);
nand U4326 (N_4326,N_4125,N_4171);
or U4327 (N_4327,N_4028,N_4104);
or U4328 (N_4328,N_4166,N_4188);
nor U4329 (N_4329,N_4093,N_4072);
and U4330 (N_4330,N_4178,N_4040);
and U4331 (N_4331,N_4193,N_4165);
and U4332 (N_4332,N_4176,N_4066);
nand U4333 (N_4333,N_4079,N_4053);
xor U4334 (N_4334,N_4087,N_4133);
nor U4335 (N_4335,N_4128,N_4054);
nand U4336 (N_4336,N_4074,N_4139);
nand U4337 (N_4337,N_4127,N_4149);
nand U4338 (N_4338,N_4046,N_4057);
or U4339 (N_4339,N_4062,N_4176);
nor U4340 (N_4340,N_4109,N_4036);
or U4341 (N_4341,N_4147,N_4028);
or U4342 (N_4342,N_4102,N_4060);
nand U4343 (N_4343,N_4118,N_4086);
nand U4344 (N_4344,N_4122,N_4146);
nand U4345 (N_4345,N_4066,N_4118);
nor U4346 (N_4346,N_4040,N_4013);
or U4347 (N_4347,N_4010,N_4027);
and U4348 (N_4348,N_4195,N_4096);
nand U4349 (N_4349,N_4099,N_4067);
or U4350 (N_4350,N_4009,N_4163);
nand U4351 (N_4351,N_4030,N_4089);
nor U4352 (N_4352,N_4145,N_4127);
and U4353 (N_4353,N_4066,N_4061);
or U4354 (N_4354,N_4152,N_4062);
nand U4355 (N_4355,N_4021,N_4148);
nand U4356 (N_4356,N_4171,N_4192);
nand U4357 (N_4357,N_4141,N_4043);
and U4358 (N_4358,N_4032,N_4114);
or U4359 (N_4359,N_4155,N_4030);
or U4360 (N_4360,N_4116,N_4172);
nor U4361 (N_4361,N_4159,N_4167);
nor U4362 (N_4362,N_4077,N_4170);
nand U4363 (N_4363,N_4107,N_4027);
nand U4364 (N_4364,N_4134,N_4162);
nor U4365 (N_4365,N_4187,N_4128);
nand U4366 (N_4366,N_4141,N_4163);
nor U4367 (N_4367,N_4076,N_4089);
and U4368 (N_4368,N_4165,N_4161);
nand U4369 (N_4369,N_4175,N_4008);
and U4370 (N_4370,N_4153,N_4029);
and U4371 (N_4371,N_4014,N_4194);
nor U4372 (N_4372,N_4138,N_4084);
or U4373 (N_4373,N_4120,N_4034);
nor U4374 (N_4374,N_4144,N_4087);
and U4375 (N_4375,N_4066,N_4014);
and U4376 (N_4376,N_4185,N_4184);
or U4377 (N_4377,N_4106,N_4062);
or U4378 (N_4378,N_4147,N_4174);
nor U4379 (N_4379,N_4058,N_4047);
or U4380 (N_4380,N_4153,N_4057);
and U4381 (N_4381,N_4003,N_4139);
and U4382 (N_4382,N_4184,N_4025);
and U4383 (N_4383,N_4160,N_4067);
and U4384 (N_4384,N_4187,N_4000);
or U4385 (N_4385,N_4068,N_4072);
or U4386 (N_4386,N_4184,N_4077);
or U4387 (N_4387,N_4116,N_4087);
or U4388 (N_4388,N_4131,N_4146);
and U4389 (N_4389,N_4072,N_4075);
or U4390 (N_4390,N_4120,N_4023);
or U4391 (N_4391,N_4092,N_4186);
and U4392 (N_4392,N_4095,N_4058);
nand U4393 (N_4393,N_4006,N_4004);
or U4394 (N_4394,N_4131,N_4087);
and U4395 (N_4395,N_4063,N_4021);
or U4396 (N_4396,N_4038,N_4120);
nor U4397 (N_4397,N_4072,N_4170);
nor U4398 (N_4398,N_4122,N_4110);
nor U4399 (N_4399,N_4128,N_4106);
nand U4400 (N_4400,N_4292,N_4348);
nand U4401 (N_4401,N_4347,N_4342);
and U4402 (N_4402,N_4244,N_4273);
nor U4403 (N_4403,N_4246,N_4313);
nor U4404 (N_4404,N_4207,N_4304);
and U4405 (N_4405,N_4306,N_4212);
and U4406 (N_4406,N_4365,N_4202);
and U4407 (N_4407,N_4320,N_4235);
nor U4408 (N_4408,N_4318,N_4255);
nand U4409 (N_4409,N_4307,N_4383);
nand U4410 (N_4410,N_4262,N_4370);
nor U4411 (N_4411,N_4269,N_4302);
nor U4412 (N_4412,N_4206,N_4381);
and U4413 (N_4413,N_4366,N_4253);
nor U4414 (N_4414,N_4200,N_4279);
or U4415 (N_4415,N_4205,N_4360);
and U4416 (N_4416,N_4277,N_4225);
or U4417 (N_4417,N_4276,N_4204);
nand U4418 (N_4418,N_4329,N_4355);
and U4419 (N_4419,N_4346,N_4295);
or U4420 (N_4420,N_4374,N_4397);
nand U4421 (N_4421,N_4311,N_4266);
nor U4422 (N_4422,N_4331,N_4268);
nor U4423 (N_4423,N_4267,N_4376);
and U4424 (N_4424,N_4245,N_4251);
nor U4425 (N_4425,N_4362,N_4315);
and U4426 (N_4426,N_4394,N_4248);
nand U4427 (N_4427,N_4389,N_4211);
nor U4428 (N_4428,N_4340,N_4236);
and U4429 (N_4429,N_4231,N_4361);
nor U4430 (N_4430,N_4343,N_4285);
nor U4431 (N_4431,N_4289,N_4378);
nor U4432 (N_4432,N_4221,N_4291);
and U4433 (N_4433,N_4264,N_4241);
or U4434 (N_4434,N_4377,N_4368);
nand U4435 (N_4435,N_4338,N_4300);
nand U4436 (N_4436,N_4336,N_4201);
nor U4437 (N_4437,N_4363,N_4259);
and U4438 (N_4438,N_4213,N_4252);
or U4439 (N_4439,N_4278,N_4274);
nor U4440 (N_4440,N_4327,N_4228);
nand U4441 (N_4441,N_4293,N_4230);
nor U4442 (N_4442,N_4356,N_4287);
xnor U4443 (N_4443,N_4358,N_4271);
and U4444 (N_4444,N_4232,N_4238);
and U4445 (N_4445,N_4284,N_4280);
nand U4446 (N_4446,N_4334,N_4385);
nand U4447 (N_4447,N_4237,N_4314);
or U4448 (N_4448,N_4239,N_4249);
or U4449 (N_4449,N_4233,N_4282);
or U4450 (N_4450,N_4303,N_4390);
xnor U4451 (N_4451,N_4222,N_4240);
and U4452 (N_4452,N_4395,N_4301);
nor U4453 (N_4453,N_4387,N_4257);
or U4454 (N_4454,N_4234,N_4350);
nor U4455 (N_4455,N_4396,N_4321);
nor U4456 (N_4456,N_4261,N_4333);
nor U4457 (N_4457,N_4297,N_4369);
or U4458 (N_4458,N_4217,N_4218);
nor U4459 (N_4459,N_4220,N_4345);
or U4460 (N_4460,N_4226,N_4353);
nor U4461 (N_4461,N_4290,N_4392);
nand U4462 (N_4462,N_4312,N_4281);
or U4463 (N_4463,N_4243,N_4299);
nor U4464 (N_4464,N_4349,N_4323);
nand U4465 (N_4465,N_4382,N_4393);
nor U4466 (N_4466,N_4351,N_4324);
and U4467 (N_4467,N_4247,N_4317);
and U4468 (N_4468,N_4364,N_4332);
or U4469 (N_4469,N_4399,N_4316);
nor U4470 (N_4470,N_4254,N_4341);
and U4471 (N_4471,N_4319,N_4337);
nor U4472 (N_4472,N_4250,N_4258);
nand U4473 (N_4473,N_4270,N_4242);
nor U4474 (N_4474,N_4308,N_4224);
nor U4475 (N_4475,N_4344,N_4256);
nor U4476 (N_4476,N_4309,N_4325);
and U4477 (N_4477,N_4354,N_4263);
or U4478 (N_4478,N_4367,N_4203);
nand U4479 (N_4479,N_4379,N_4391);
and U4480 (N_4480,N_4216,N_4352);
nand U4481 (N_4481,N_4388,N_4380);
nor U4482 (N_4482,N_4214,N_4305);
or U4483 (N_4483,N_4330,N_4272);
nor U4484 (N_4484,N_4265,N_4219);
or U4485 (N_4485,N_4372,N_4210);
and U4486 (N_4486,N_4326,N_4283);
and U4487 (N_4487,N_4328,N_4384);
and U4488 (N_4488,N_4215,N_4371);
and U4489 (N_4489,N_4288,N_4286);
and U4490 (N_4490,N_4223,N_4298);
or U4491 (N_4491,N_4335,N_4359);
nor U4492 (N_4492,N_4310,N_4386);
nor U4493 (N_4493,N_4373,N_4375);
nor U4494 (N_4494,N_4260,N_4296);
and U4495 (N_4495,N_4227,N_4275);
and U4496 (N_4496,N_4208,N_4322);
and U4497 (N_4497,N_4357,N_4209);
nand U4498 (N_4498,N_4294,N_4398);
nor U4499 (N_4499,N_4339,N_4229);
or U4500 (N_4500,N_4202,N_4266);
or U4501 (N_4501,N_4306,N_4373);
nor U4502 (N_4502,N_4331,N_4343);
and U4503 (N_4503,N_4224,N_4397);
nand U4504 (N_4504,N_4200,N_4320);
and U4505 (N_4505,N_4293,N_4257);
nor U4506 (N_4506,N_4224,N_4388);
nand U4507 (N_4507,N_4232,N_4297);
nor U4508 (N_4508,N_4257,N_4355);
nand U4509 (N_4509,N_4259,N_4334);
nor U4510 (N_4510,N_4290,N_4368);
nor U4511 (N_4511,N_4380,N_4363);
nor U4512 (N_4512,N_4384,N_4355);
nor U4513 (N_4513,N_4215,N_4330);
nor U4514 (N_4514,N_4348,N_4303);
and U4515 (N_4515,N_4370,N_4338);
or U4516 (N_4516,N_4326,N_4266);
or U4517 (N_4517,N_4238,N_4252);
nor U4518 (N_4518,N_4203,N_4352);
nor U4519 (N_4519,N_4249,N_4305);
nor U4520 (N_4520,N_4262,N_4357);
and U4521 (N_4521,N_4221,N_4333);
and U4522 (N_4522,N_4360,N_4305);
nand U4523 (N_4523,N_4379,N_4327);
nand U4524 (N_4524,N_4215,N_4342);
nor U4525 (N_4525,N_4265,N_4270);
nor U4526 (N_4526,N_4250,N_4289);
nand U4527 (N_4527,N_4363,N_4254);
or U4528 (N_4528,N_4313,N_4366);
or U4529 (N_4529,N_4210,N_4324);
nand U4530 (N_4530,N_4385,N_4366);
nor U4531 (N_4531,N_4205,N_4305);
or U4532 (N_4532,N_4281,N_4273);
nor U4533 (N_4533,N_4391,N_4286);
and U4534 (N_4534,N_4256,N_4395);
or U4535 (N_4535,N_4205,N_4233);
or U4536 (N_4536,N_4207,N_4302);
nor U4537 (N_4537,N_4336,N_4293);
nand U4538 (N_4538,N_4206,N_4276);
and U4539 (N_4539,N_4373,N_4258);
nand U4540 (N_4540,N_4251,N_4239);
nand U4541 (N_4541,N_4323,N_4392);
and U4542 (N_4542,N_4223,N_4338);
or U4543 (N_4543,N_4337,N_4350);
nand U4544 (N_4544,N_4275,N_4287);
or U4545 (N_4545,N_4391,N_4371);
nand U4546 (N_4546,N_4261,N_4290);
nor U4547 (N_4547,N_4244,N_4233);
and U4548 (N_4548,N_4269,N_4266);
and U4549 (N_4549,N_4236,N_4391);
and U4550 (N_4550,N_4235,N_4213);
nand U4551 (N_4551,N_4391,N_4348);
nand U4552 (N_4552,N_4380,N_4361);
and U4553 (N_4553,N_4380,N_4315);
or U4554 (N_4554,N_4364,N_4226);
nor U4555 (N_4555,N_4372,N_4343);
or U4556 (N_4556,N_4214,N_4221);
nor U4557 (N_4557,N_4202,N_4278);
nor U4558 (N_4558,N_4298,N_4228);
nand U4559 (N_4559,N_4221,N_4268);
nand U4560 (N_4560,N_4301,N_4200);
or U4561 (N_4561,N_4379,N_4330);
nor U4562 (N_4562,N_4253,N_4383);
nor U4563 (N_4563,N_4289,N_4377);
nor U4564 (N_4564,N_4220,N_4215);
nor U4565 (N_4565,N_4209,N_4336);
nor U4566 (N_4566,N_4206,N_4349);
and U4567 (N_4567,N_4237,N_4393);
and U4568 (N_4568,N_4376,N_4252);
nand U4569 (N_4569,N_4208,N_4247);
or U4570 (N_4570,N_4260,N_4329);
or U4571 (N_4571,N_4344,N_4333);
or U4572 (N_4572,N_4226,N_4305);
or U4573 (N_4573,N_4377,N_4220);
xnor U4574 (N_4574,N_4377,N_4320);
nor U4575 (N_4575,N_4256,N_4278);
and U4576 (N_4576,N_4307,N_4252);
nand U4577 (N_4577,N_4260,N_4320);
nor U4578 (N_4578,N_4342,N_4388);
or U4579 (N_4579,N_4383,N_4218);
nor U4580 (N_4580,N_4283,N_4214);
nor U4581 (N_4581,N_4266,N_4253);
and U4582 (N_4582,N_4331,N_4245);
nand U4583 (N_4583,N_4244,N_4201);
and U4584 (N_4584,N_4267,N_4389);
nand U4585 (N_4585,N_4286,N_4254);
nand U4586 (N_4586,N_4322,N_4387);
and U4587 (N_4587,N_4361,N_4384);
or U4588 (N_4588,N_4207,N_4220);
and U4589 (N_4589,N_4353,N_4305);
nand U4590 (N_4590,N_4368,N_4284);
nor U4591 (N_4591,N_4346,N_4384);
nor U4592 (N_4592,N_4205,N_4317);
nor U4593 (N_4593,N_4303,N_4242);
or U4594 (N_4594,N_4220,N_4359);
nor U4595 (N_4595,N_4244,N_4313);
nand U4596 (N_4596,N_4380,N_4340);
nand U4597 (N_4597,N_4280,N_4378);
nand U4598 (N_4598,N_4303,N_4231);
and U4599 (N_4599,N_4266,N_4327);
nor U4600 (N_4600,N_4447,N_4505);
nand U4601 (N_4601,N_4514,N_4589);
and U4602 (N_4602,N_4477,N_4592);
and U4603 (N_4603,N_4487,N_4425);
or U4604 (N_4604,N_4462,N_4556);
and U4605 (N_4605,N_4405,N_4433);
and U4606 (N_4606,N_4492,N_4461);
or U4607 (N_4607,N_4407,N_4423);
and U4608 (N_4608,N_4478,N_4580);
xor U4609 (N_4609,N_4403,N_4472);
or U4610 (N_4610,N_4550,N_4490);
nand U4611 (N_4611,N_4553,N_4518);
nand U4612 (N_4612,N_4561,N_4559);
or U4613 (N_4613,N_4460,N_4570);
nor U4614 (N_4614,N_4546,N_4511);
or U4615 (N_4615,N_4568,N_4416);
nand U4616 (N_4616,N_4410,N_4464);
nor U4617 (N_4617,N_4493,N_4577);
xnor U4618 (N_4618,N_4564,N_4434);
nor U4619 (N_4619,N_4418,N_4409);
and U4620 (N_4620,N_4582,N_4566);
and U4621 (N_4621,N_4470,N_4579);
nor U4622 (N_4622,N_4571,N_4507);
nand U4623 (N_4623,N_4541,N_4486);
nor U4624 (N_4624,N_4458,N_4456);
nand U4625 (N_4625,N_4557,N_4465);
nand U4626 (N_4626,N_4598,N_4453);
nand U4627 (N_4627,N_4573,N_4413);
nor U4628 (N_4628,N_4593,N_4414);
and U4629 (N_4629,N_4411,N_4481);
nand U4630 (N_4630,N_4401,N_4536);
nor U4631 (N_4631,N_4599,N_4548);
nand U4632 (N_4632,N_4535,N_4502);
or U4633 (N_4633,N_4545,N_4555);
nor U4634 (N_4634,N_4552,N_4591);
nand U4635 (N_4635,N_4448,N_4578);
and U4636 (N_4636,N_4574,N_4476);
nor U4637 (N_4637,N_4595,N_4585);
nand U4638 (N_4638,N_4499,N_4584);
nand U4639 (N_4639,N_4506,N_4521);
or U4640 (N_4640,N_4430,N_4549);
and U4641 (N_4641,N_4417,N_4594);
and U4642 (N_4642,N_4415,N_4563);
nand U4643 (N_4643,N_4431,N_4451);
or U4644 (N_4644,N_4468,N_4420);
or U4645 (N_4645,N_4404,N_4491);
and U4646 (N_4646,N_4428,N_4586);
or U4647 (N_4647,N_4587,N_4575);
or U4648 (N_4648,N_4479,N_4484);
nand U4649 (N_4649,N_4466,N_4554);
or U4650 (N_4650,N_4443,N_4531);
nor U4651 (N_4651,N_4495,N_4583);
nor U4652 (N_4652,N_4444,N_4565);
and U4653 (N_4653,N_4527,N_4436);
nor U4654 (N_4654,N_4588,N_4560);
or U4655 (N_4655,N_4529,N_4424);
nor U4656 (N_4656,N_4497,N_4569);
and U4657 (N_4657,N_4543,N_4452);
nor U4658 (N_4658,N_4540,N_4526);
nand U4659 (N_4659,N_4515,N_4551);
nand U4660 (N_4660,N_4509,N_4475);
nand U4661 (N_4661,N_4498,N_4567);
nor U4662 (N_4662,N_4525,N_4508);
or U4663 (N_4663,N_4489,N_4441);
nor U4664 (N_4664,N_4520,N_4496);
nand U4665 (N_4665,N_4503,N_4442);
nand U4666 (N_4666,N_4500,N_4422);
nor U4667 (N_4667,N_4547,N_4440);
or U4668 (N_4668,N_4528,N_4412);
or U4669 (N_4669,N_4483,N_4538);
or U4670 (N_4670,N_4519,N_4494);
nor U4671 (N_4671,N_4419,N_4480);
nor U4672 (N_4672,N_4421,N_4473);
nand U4673 (N_4673,N_4469,N_4501);
nand U4674 (N_4674,N_4542,N_4590);
and U4675 (N_4675,N_4534,N_4467);
nand U4676 (N_4676,N_4400,N_4438);
nand U4677 (N_4677,N_4471,N_4510);
nor U4678 (N_4678,N_4539,N_4482);
nand U4679 (N_4679,N_4463,N_4524);
or U4680 (N_4680,N_4485,N_4512);
nand U4681 (N_4681,N_4408,N_4474);
nand U4682 (N_4682,N_4544,N_4459);
or U4683 (N_4683,N_4576,N_4516);
and U4684 (N_4684,N_4504,N_4445);
nor U4685 (N_4685,N_4454,N_4533);
nor U4686 (N_4686,N_4435,N_4432);
and U4687 (N_4687,N_4449,N_4532);
nor U4688 (N_4688,N_4446,N_4455);
nor U4689 (N_4689,N_4426,N_4513);
and U4690 (N_4690,N_4450,N_4596);
or U4691 (N_4691,N_4530,N_4522);
nand U4692 (N_4692,N_4406,N_4439);
nand U4693 (N_4693,N_4402,N_4572);
or U4694 (N_4694,N_4597,N_4488);
and U4695 (N_4695,N_4562,N_4517);
and U4696 (N_4696,N_4457,N_4537);
nand U4697 (N_4697,N_4437,N_4581);
nor U4698 (N_4698,N_4523,N_4427);
nand U4699 (N_4699,N_4558,N_4429);
or U4700 (N_4700,N_4556,N_4478);
nor U4701 (N_4701,N_4440,N_4517);
xnor U4702 (N_4702,N_4471,N_4532);
or U4703 (N_4703,N_4591,N_4565);
nor U4704 (N_4704,N_4450,N_4493);
nand U4705 (N_4705,N_4410,N_4473);
xor U4706 (N_4706,N_4465,N_4420);
nor U4707 (N_4707,N_4560,N_4530);
or U4708 (N_4708,N_4436,N_4513);
xor U4709 (N_4709,N_4592,N_4474);
nor U4710 (N_4710,N_4447,N_4552);
nor U4711 (N_4711,N_4561,N_4404);
and U4712 (N_4712,N_4542,N_4419);
nor U4713 (N_4713,N_4575,N_4504);
nor U4714 (N_4714,N_4426,N_4530);
and U4715 (N_4715,N_4506,N_4592);
and U4716 (N_4716,N_4412,N_4547);
or U4717 (N_4717,N_4540,N_4513);
or U4718 (N_4718,N_4523,N_4555);
or U4719 (N_4719,N_4576,N_4523);
nor U4720 (N_4720,N_4482,N_4557);
nand U4721 (N_4721,N_4563,N_4571);
and U4722 (N_4722,N_4505,N_4430);
and U4723 (N_4723,N_4454,N_4531);
or U4724 (N_4724,N_4544,N_4477);
nand U4725 (N_4725,N_4483,N_4438);
and U4726 (N_4726,N_4494,N_4505);
or U4727 (N_4727,N_4430,N_4473);
or U4728 (N_4728,N_4594,N_4483);
xnor U4729 (N_4729,N_4505,N_4453);
and U4730 (N_4730,N_4564,N_4404);
nand U4731 (N_4731,N_4529,N_4533);
nor U4732 (N_4732,N_4448,N_4435);
or U4733 (N_4733,N_4568,N_4481);
and U4734 (N_4734,N_4526,N_4486);
nand U4735 (N_4735,N_4428,N_4531);
or U4736 (N_4736,N_4503,N_4410);
nand U4737 (N_4737,N_4429,N_4547);
nor U4738 (N_4738,N_4444,N_4563);
nor U4739 (N_4739,N_4545,N_4463);
nor U4740 (N_4740,N_4549,N_4429);
nand U4741 (N_4741,N_4525,N_4460);
or U4742 (N_4742,N_4576,N_4482);
and U4743 (N_4743,N_4464,N_4479);
nor U4744 (N_4744,N_4528,N_4585);
nor U4745 (N_4745,N_4556,N_4593);
or U4746 (N_4746,N_4464,N_4547);
or U4747 (N_4747,N_4421,N_4525);
nand U4748 (N_4748,N_4591,N_4437);
nor U4749 (N_4749,N_4470,N_4400);
nand U4750 (N_4750,N_4586,N_4484);
or U4751 (N_4751,N_4570,N_4493);
and U4752 (N_4752,N_4577,N_4567);
or U4753 (N_4753,N_4494,N_4555);
nand U4754 (N_4754,N_4469,N_4470);
and U4755 (N_4755,N_4573,N_4402);
and U4756 (N_4756,N_4551,N_4527);
xor U4757 (N_4757,N_4474,N_4584);
nand U4758 (N_4758,N_4486,N_4553);
or U4759 (N_4759,N_4525,N_4536);
or U4760 (N_4760,N_4412,N_4480);
nor U4761 (N_4761,N_4506,N_4554);
or U4762 (N_4762,N_4586,N_4541);
and U4763 (N_4763,N_4582,N_4487);
nor U4764 (N_4764,N_4584,N_4467);
nor U4765 (N_4765,N_4551,N_4489);
nor U4766 (N_4766,N_4563,N_4496);
or U4767 (N_4767,N_4544,N_4469);
nand U4768 (N_4768,N_4520,N_4410);
nor U4769 (N_4769,N_4496,N_4457);
or U4770 (N_4770,N_4539,N_4541);
or U4771 (N_4771,N_4521,N_4476);
nor U4772 (N_4772,N_4410,N_4421);
nand U4773 (N_4773,N_4458,N_4467);
nand U4774 (N_4774,N_4416,N_4502);
nand U4775 (N_4775,N_4558,N_4561);
nor U4776 (N_4776,N_4449,N_4474);
or U4777 (N_4777,N_4524,N_4485);
and U4778 (N_4778,N_4450,N_4457);
nor U4779 (N_4779,N_4456,N_4524);
nor U4780 (N_4780,N_4568,N_4584);
nand U4781 (N_4781,N_4452,N_4503);
or U4782 (N_4782,N_4513,N_4529);
nor U4783 (N_4783,N_4519,N_4476);
nor U4784 (N_4784,N_4508,N_4435);
nor U4785 (N_4785,N_4580,N_4476);
nand U4786 (N_4786,N_4502,N_4496);
or U4787 (N_4787,N_4587,N_4509);
nand U4788 (N_4788,N_4411,N_4549);
and U4789 (N_4789,N_4522,N_4579);
and U4790 (N_4790,N_4452,N_4488);
nand U4791 (N_4791,N_4597,N_4471);
or U4792 (N_4792,N_4432,N_4584);
nor U4793 (N_4793,N_4597,N_4551);
and U4794 (N_4794,N_4402,N_4457);
or U4795 (N_4795,N_4438,N_4552);
nor U4796 (N_4796,N_4562,N_4429);
and U4797 (N_4797,N_4512,N_4581);
nand U4798 (N_4798,N_4575,N_4485);
nand U4799 (N_4799,N_4433,N_4506);
nand U4800 (N_4800,N_4755,N_4716);
nor U4801 (N_4801,N_4663,N_4647);
or U4802 (N_4802,N_4637,N_4707);
or U4803 (N_4803,N_4681,N_4727);
nor U4804 (N_4804,N_4714,N_4666);
or U4805 (N_4805,N_4787,N_4679);
or U4806 (N_4806,N_4771,N_4762);
or U4807 (N_4807,N_4708,N_4724);
nor U4808 (N_4808,N_4756,N_4757);
nand U4809 (N_4809,N_4741,N_4743);
and U4810 (N_4810,N_4720,N_4635);
and U4811 (N_4811,N_4703,N_4791);
and U4812 (N_4812,N_4797,N_4618);
nor U4813 (N_4813,N_4626,N_4786);
nand U4814 (N_4814,N_4682,N_4601);
nand U4815 (N_4815,N_4654,N_4646);
nor U4816 (N_4816,N_4617,N_4631);
or U4817 (N_4817,N_4792,N_4783);
nand U4818 (N_4818,N_4701,N_4649);
or U4819 (N_4819,N_4746,N_4697);
and U4820 (N_4820,N_4672,N_4690);
nand U4821 (N_4821,N_4723,N_4713);
or U4822 (N_4822,N_4789,N_4614);
nand U4823 (N_4823,N_4712,N_4625);
and U4824 (N_4824,N_4624,N_4606);
nand U4825 (N_4825,N_4754,N_4760);
nand U4826 (N_4826,N_4655,N_4775);
or U4827 (N_4827,N_4739,N_4653);
nor U4828 (N_4828,N_4761,N_4719);
and U4829 (N_4829,N_4657,N_4639);
and U4830 (N_4830,N_4699,N_4778);
nand U4831 (N_4831,N_4749,N_4620);
or U4832 (N_4832,N_4656,N_4628);
nand U4833 (N_4833,N_4702,N_4600);
and U4834 (N_4834,N_4678,N_4621);
or U4835 (N_4835,N_4717,N_4773);
or U4836 (N_4836,N_4652,N_4742);
nand U4837 (N_4837,N_4684,N_4664);
nand U4838 (N_4838,N_4694,N_4715);
nor U4839 (N_4839,N_4610,N_4732);
or U4840 (N_4840,N_4651,N_4740);
nor U4841 (N_4841,N_4636,N_4602);
nand U4842 (N_4842,N_4634,N_4726);
or U4843 (N_4843,N_4764,N_4765);
nand U4844 (N_4844,N_4766,N_4662);
nand U4845 (N_4845,N_4758,N_4645);
and U4846 (N_4846,N_4680,N_4770);
or U4847 (N_4847,N_4745,N_4613);
nand U4848 (N_4848,N_4648,N_4768);
nand U4849 (N_4849,N_4795,N_4643);
nand U4850 (N_4850,N_4794,N_4733);
nor U4851 (N_4851,N_4661,N_4675);
nand U4852 (N_4852,N_4744,N_4772);
nand U4853 (N_4853,N_4698,N_4706);
nor U4854 (N_4854,N_4734,N_4627);
nand U4855 (N_4855,N_4676,N_4692);
nand U4856 (N_4856,N_4670,N_4659);
nand U4857 (N_4857,N_4780,N_4799);
xor U4858 (N_4858,N_4668,N_4641);
nand U4859 (N_4859,N_4763,N_4777);
nand U4860 (N_4860,N_4753,N_4725);
nand U4861 (N_4861,N_4752,N_4677);
or U4862 (N_4862,N_4750,N_4738);
and U4863 (N_4863,N_4759,N_4779);
or U4864 (N_4864,N_4693,N_4623);
or U4865 (N_4865,N_4671,N_4689);
nor U4866 (N_4866,N_4683,N_4774);
nand U4867 (N_4867,N_4687,N_4711);
and U4868 (N_4868,N_4709,N_4619);
or U4869 (N_4869,N_4607,N_4731);
nand U4870 (N_4870,N_4767,N_4644);
nor U4871 (N_4871,N_4629,N_4695);
or U4872 (N_4872,N_4609,N_4710);
nand U4873 (N_4873,N_4796,N_4630);
nor U4874 (N_4874,N_4665,N_4688);
nand U4875 (N_4875,N_4642,N_4669);
and U4876 (N_4876,N_4776,N_4769);
nor U4877 (N_4877,N_4640,N_4705);
or U4878 (N_4878,N_4660,N_4798);
nand U4879 (N_4879,N_4729,N_4751);
nand U4880 (N_4880,N_4728,N_4632);
or U4881 (N_4881,N_4748,N_4735);
or U4882 (N_4882,N_4686,N_4658);
nor U4883 (N_4883,N_4700,N_4608);
and U4884 (N_4884,N_4782,N_4785);
or U4885 (N_4885,N_4747,N_4612);
and U4886 (N_4886,N_4722,N_4638);
and U4887 (N_4887,N_4615,N_4611);
and U4888 (N_4888,N_4736,N_4788);
nor U4889 (N_4889,N_4781,N_4696);
nor U4890 (N_4890,N_4737,N_4793);
xnor U4891 (N_4891,N_4603,N_4691);
and U4892 (N_4892,N_4622,N_4718);
or U4893 (N_4893,N_4616,N_4633);
and U4894 (N_4894,N_4685,N_4650);
nand U4895 (N_4895,N_4730,N_4784);
and U4896 (N_4896,N_4704,N_4790);
nor U4897 (N_4897,N_4721,N_4605);
or U4898 (N_4898,N_4674,N_4604);
or U4899 (N_4899,N_4673,N_4667);
nor U4900 (N_4900,N_4694,N_4699);
nand U4901 (N_4901,N_4710,N_4798);
nor U4902 (N_4902,N_4721,N_4607);
nor U4903 (N_4903,N_4786,N_4682);
and U4904 (N_4904,N_4685,N_4648);
nor U4905 (N_4905,N_4722,N_4606);
or U4906 (N_4906,N_4685,N_4711);
or U4907 (N_4907,N_4655,N_4732);
and U4908 (N_4908,N_4644,N_4649);
or U4909 (N_4909,N_4635,N_4619);
nand U4910 (N_4910,N_4623,N_4784);
nand U4911 (N_4911,N_4694,N_4739);
nor U4912 (N_4912,N_4699,N_4610);
or U4913 (N_4913,N_4784,N_4728);
nand U4914 (N_4914,N_4610,N_4618);
xor U4915 (N_4915,N_4727,N_4671);
nor U4916 (N_4916,N_4641,N_4710);
or U4917 (N_4917,N_4765,N_4722);
nand U4918 (N_4918,N_4730,N_4654);
or U4919 (N_4919,N_4720,N_4782);
and U4920 (N_4920,N_4669,N_4689);
or U4921 (N_4921,N_4652,N_4637);
and U4922 (N_4922,N_4676,N_4663);
and U4923 (N_4923,N_4681,N_4716);
and U4924 (N_4924,N_4745,N_4744);
nor U4925 (N_4925,N_4680,N_4736);
nand U4926 (N_4926,N_4745,N_4766);
and U4927 (N_4927,N_4602,N_4785);
nor U4928 (N_4928,N_4644,N_4631);
and U4929 (N_4929,N_4637,N_4630);
and U4930 (N_4930,N_4678,N_4669);
or U4931 (N_4931,N_4623,N_4729);
or U4932 (N_4932,N_4727,N_4669);
nor U4933 (N_4933,N_4694,N_4658);
or U4934 (N_4934,N_4655,N_4792);
and U4935 (N_4935,N_4786,N_4722);
and U4936 (N_4936,N_4672,N_4635);
nand U4937 (N_4937,N_4686,N_4629);
nand U4938 (N_4938,N_4772,N_4765);
nor U4939 (N_4939,N_4683,N_4736);
and U4940 (N_4940,N_4765,N_4741);
nor U4941 (N_4941,N_4708,N_4760);
nand U4942 (N_4942,N_4689,N_4719);
and U4943 (N_4943,N_4636,N_4755);
nand U4944 (N_4944,N_4698,N_4611);
nand U4945 (N_4945,N_4728,N_4683);
xnor U4946 (N_4946,N_4686,N_4682);
and U4947 (N_4947,N_4796,N_4615);
and U4948 (N_4948,N_4640,N_4792);
and U4949 (N_4949,N_4765,N_4677);
nand U4950 (N_4950,N_4642,N_4694);
or U4951 (N_4951,N_4605,N_4755);
nor U4952 (N_4952,N_4786,N_4761);
nor U4953 (N_4953,N_4719,N_4694);
nor U4954 (N_4954,N_4606,N_4766);
nor U4955 (N_4955,N_4734,N_4752);
nand U4956 (N_4956,N_4740,N_4724);
nand U4957 (N_4957,N_4705,N_4744);
and U4958 (N_4958,N_4651,N_4679);
or U4959 (N_4959,N_4688,N_4782);
nor U4960 (N_4960,N_4711,N_4738);
or U4961 (N_4961,N_4677,N_4784);
nand U4962 (N_4962,N_4728,N_4775);
and U4963 (N_4963,N_4635,N_4626);
and U4964 (N_4964,N_4600,N_4687);
nor U4965 (N_4965,N_4705,N_4772);
and U4966 (N_4966,N_4612,N_4795);
nor U4967 (N_4967,N_4791,N_4758);
xor U4968 (N_4968,N_4771,N_4634);
nand U4969 (N_4969,N_4741,N_4754);
or U4970 (N_4970,N_4698,N_4780);
or U4971 (N_4971,N_4600,N_4775);
nand U4972 (N_4972,N_4798,N_4604);
or U4973 (N_4973,N_4624,N_4620);
nand U4974 (N_4974,N_4706,N_4796);
nand U4975 (N_4975,N_4606,N_4767);
nor U4976 (N_4976,N_4753,N_4781);
or U4977 (N_4977,N_4740,N_4647);
or U4978 (N_4978,N_4665,N_4721);
and U4979 (N_4979,N_4753,N_4617);
nor U4980 (N_4980,N_4679,N_4722);
nor U4981 (N_4981,N_4793,N_4615);
or U4982 (N_4982,N_4641,N_4691);
nand U4983 (N_4983,N_4658,N_4767);
and U4984 (N_4984,N_4766,N_4636);
nand U4985 (N_4985,N_4789,N_4688);
nor U4986 (N_4986,N_4682,N_4765);
nand U4987 (N_4987,N_4644,N_4742);
nor U4988 (N_4988,N_4737,N_4626);
nor U4989 (N_4989,N_4671,N_4694);
nor U4990 (N_4990,N_4742,N_4637);
or U4991 (N_4991,N_4643,N_4742);
or U4992 (N_4992,N_4754,N_4718);
and U4993 (N_4993,N_4719,N_4705);
nor U4994 (N_4994,N_4777,N_4708);
and U4995 (N_4995,N_4770,N_4781);
nor U4996 (N_4996,N_4628,N_4663);
nand U4997 (N_4997,N_4720,N_4739);
nor U4998 (N_4998,N_4695,N_4643);
and U4999 (N_4999,N_4724,N_4788);
and UO_0 (O_0,N_4879,N_4963);
and UO_1 (O_1,N_4870,N_4903);
nand UO_2 (O_2,N_4966,N_4864);
and UO_3 (O_3,N_4910,N_4956);
xor UO_4 (O_4,N_4824,N_4898);
nand UO_5 (O_5,N_4952,N_4855);
nand UO_6 (O_6,N_4983,N_4920);
nor UO_7 (O_7,N_4816,N_4951);
or UO_8 (O_8,N_4852,N_4974);
and UO_9 (O_9,N_4821,N_4909);
nor UO_10 (O_10,N_4861,N_4978);
or UO_11 (O_11,N_4945,N_4815);
nand UO_12 (O_12,N_4936,N_4817);
nor UO_13 (O_13,N_4930,N_4906);
nand UO_14 (O_14,N_4929,N_4919);
and UO_15 (O_15,N_4986,N_4880);
nand UO_16 (O_16,N_4887,N_4800);
nor UO_17 (O_17,N_4882,N_4829);
or UO_18 (O_18,N_4877,N_4913);
nor UO_19 (O_19,N_4885,N_4865);
xnor UO_20 (O_20,N_4988,N_4976);
and UO_21 (O_21,N_4914,N_4862);
and UO_22 (O_22,N_4933,N_4960);
nand UO_23 (O_23,N_4899,N_4977);
nor UO_24 (O_24,N_4957,N_4999);
and UO_25 (O_25,N_4836,N_4911);
or UO_26 (O_26,N_4912,N_4959);
nor UO_27 (O_27,N_4874,N_4811);
and UO_28 (O_28,N_4840,N_4946);
nor UO_29 (O_29,N_4856,N_4843);
and UO_30 (O_30,N_4834,N_4838);
and UO_31 (O_31,N_4915,N_4812);
nor UO_32 (O_32,N_4828,N_4889);
nand UO_33 (O_33,N_4854,N_4964);
or UO_34 (O_34,N_4878,N_4806);
or UO_35 (O_35,N_4801,N_4975);
nor UO_36 (O_36,N_4979,N_4891);
nand UO_37 (O_37,N_4860,N_4844);
xnor UO_38 (O_38,N_4804,N_4897);
or UO_39 (O_39,N_4851,N_4827);
nor UO_40 (O_40,N_4990,N_4819);
nand UO_41 (O_41,N_4932,N_4872);
or UO_42 (O_42,N_4802,N_4900);
and UO_43 (O_43,N_4892,N_4810);
nand UO_44 (O_44,N_4833,N_4926);
nand UO_45 (O_45,N_4876,N_4907);
and UO_46 (O_46,N_4895,N_4867);
nor UO_47 (O_47,N_4905,N_4995);
nand UO_48 (O_48,N_4841,N_4961);
and UO_49 (O_49,N_4848,N_4808);
nor UO_50 (O_50,N_4928,N_4813);
and UO_51 (O_51,N_4820,N_4883);
nor UO_52 (O_52,N_4871,N_4931);
nand UO_53 (O_53,N_4925,N_4866);
xnor UO_54 (O_54,N_4904,N_4896);
nand UO_55 (O_55,N_4837,N_4832);
nor UO_56 (O_56,N_4980,N_4846);
xnor UO_57 (O_57,N_4849,N_4958);
nor UO_58 (O_58,N_4921,N_4888);
nand UO_59 (O_59,N_4992,N_4868);
and UO_60 (O_60,N_4894,N_4805);
nand UO_61 (O_61,N_4994,N_4917);
nand UO_62 (O_62,N_4941,N_4985);
and UO_63 (O_63,N_4901,N_4949);
nand UO_64 (O_64,N_4916,N_4850);
or UO_65 (O_65,N_4962,N_4902);
nand UO_66 (O_66,N_4845,N_4993);
and UO_67 (O_67,N_4823,N_4981);
nand UO_68 (O_68,N_4942,N_4890);
nor UO_69 (O_69,N_4875,N_4839);
and UO_70 (O_70,N_4881,N_4968);
or UO_71 (O_71,N_4965,N_4922);
nor UO_72 (O_72,N_4873,N_4967);
or UO_73 (O_73,N_4950,N_4818);
nand UO_74 (O_74,N_4982,N_4947);
and UO_75 (O_75,N_4939,N_4908);
nor UO_76 (O_76,N_4927,N_4954);
or UO_77 (O_77,N_4953,N_4842);
nor UO_78 (O_78,N_4948,N_4858);
nor UO_79 (O_79,N_4934,N_4918);
or UO_80 (O_80,N_4998,N_4884);
nor UO_81 (O_81,N_4803,N_4938);
or UO_82 (O_82,N_4935,N_4989);
or UO_83 (O_83,N_4863,N_4923);
nand UO_84 (O_84,N_4853,N_4991);
and UO_85 (O_85,N_4814,N_4970);
nor UO_86 (O_86,N_4826,N_4984);
or UO_87 (O_87,N_4859,N_4987);
nand UO_88 (O_88,N_4893,N_4825);
nor UO_89 (O_89,N_4972,N_4943);
or UO_90 (O_90,N_4822,N_4996);
or UO_91 (O_91,N_4937,N_4847);
xnor UO_92 (O_92,N_4857,N_4997);
and UO_93 (O_93,N_4831,N_4886);
or UO_94 (O_94,N_4971,N_4940);
and UO_95 (O_95,N_4835,N_4869);
and UO_96 (O_96,N_4807,N_4973);
or UO_97 (O_97,N_4830,N_4955);
and UO_98 (O_98,N_4924,N_4969);
and UO_99 (O_99,N_4809,N_4944);
nor UO_100 (O_100,N_4981,N_4903);
and UO_101 (O_101,N_4830,N_4944);
nand UO_102 (O_102,N_4859,N_4852);
and UO_103 (O_103,N_4883,N_4895);
nand UO_104 (O_104,N_4997,N_4951);
and UO_105 (O_105,N_4884,N_4994);
nor UO_106 (O_106,N_4908,N_4827);
nor UO_107 (O_107,N_4939,N_4813);
or UO_108 (O_108,N_4891,N_4901);
nor UO_109 (O_109,N_4894,N_4847);
nand UO_110 (O_110,N_4928,N_4921);
nand UO_111 (O_111,N_4869,N_4812);
or UO_112 (O_112,N_4800,N_4898);
or UO_113 (O_113,N_4813,N_4867);
nand UO_114 (O_114,N_4813,N_4991);
nor UO_115 (O_115,N_4842,N_4880);
nor UO_116 (O_116,N_4933,N_4847);
and UO_117 (O_117,N_4896,N_4805);
nor UO_118 (O_118,N_4804,N_4937);
nand UO_119 (O_119,N_4807,N_4940);
and UO_120 (O_120,N_4884,N_4825);
nor UO_121 (O_121,N_4947,N_4830);
nor UO_122 (O_122,N_4958,N_4991);
nor UO_123 (O_123,N_4962,N_4866);
nand UO_124 (O_124,N_4933,N_4800);
and UO_125 (O_125,N_4972,N_4841);
nand UO_126 (O_126,N_4892,N_4865);
or UO_127 (O_127,N_4813,N_4842);
nor UO_128 (O_128,N_4852,N_4978);
nand UO_129 (O_129,N_4811,N_4852);
or UO_130 (O_130,N_4895,N_4992);
and UO_131 (O_131,N_4977,N_4997);
nand UO_132 (O_132,N_4974,N_4944);
and UO_133 (O_133,N_4857,N_4886);
and UO_134 (O_134,N_4890,N_4956);
nand UO_135 (O_135,N_4834,N_4987);
or UO_136 (O_136,N_4803,N_4886);
nor UO_137 (O_137,N_4992,N_4813);
nand UO_138 (O_138,N_4873,N_4927);
nand UO_139 (O_139,N_4850,N_4872);
nand UO_140 (O_140,N_4817,N_4955);
nand UO_141 (O_141,N_4876,N_4888);
nand UO_142 (O_142,N_4857,N_4845);
or UO_143 (O_143,N_4819,N_4997);
nand UO_144 (O_144,N_4842,N_4955);
and UO_145 (O_145,N_4815,N_4860);
or UO_146 (O_146,N_4905,N_4844);
and UO_147 (O_147,N_4996,N_4951);
nand UO_148 (O_148,N_4859,N_4805);
or UO_149 (O_149,N_4893,N_4947);
and UO_150 (O_150,N_4863,N_4832);
and UO_151 (O_151,N_4951,N_4821);
or UO_152 (O_152,N_4844,N_4979);
nor UO_153 (O_153,N_4928,N_4892);
or UO_154 (O_154,N_4995,N_4903);
nor UO_155 (O_155,N_4894,N_4852);
and UO_156 (O_156,N_4888,N_4920);
nor UO_157 (O_157,N_4937,N_4869);
or UO_158 (O_158,N_4827,N_4841);
or UO_159 (O_159,N_4907,N_4878);
nor UO_160 (O_160,N_4816,N_4829);
and UO_161 (O_161,N_4929,N_4859);
nor UO_162 (O_162,N_4802,N_4985);
nor UO_163 (O_163,N_4909,N_4944);
and UO_164 (O_164,N_4895,N_4927);
nor UO_165 (O_165,N_4991,N_4889);
nor UO_166 (O_166,N_4954,N_4805);
nand UO_167 (O_167,N_4985,N_4913);
nor UO_168 (O_168,N_4914,N_4972);
and UO_169 (O_169,N_4826,N_4918);
nand UO_170 (O_170,N_4949,N_4984);
or UO_171 (O_171,N_4900,N_4863);
and UO_172 (O_172,N_4812,N_4902);
xnor UO_173 (O_173,N_4833,N_4978);
or UO_174 (O_174,N_4862,N_4803);
and UO_175 (O_175,N_4806,N_4844);
nand UO_176 (O_176,N_4997,N_4827);
nand UO_177 (O_177,N_4817,N_4992);
and UO_178 (O_178,N_4914,N_4954);
nand UO_179 (O_179,N_4827,N_4812);
nor UO_180 (O_180,N_4904,N_4981);
or UO_181 (O_181,N_4917,N_4888);
nor UO_182 (O_182,N_4971,N_4842);
nand UO_183 (O_183,N_4979,N_4925);
nor UO_184 (O_184,N_4923,N_4977);
and UO_185 (O_185,N_4942,N_4818);
xor UO_186 (O_186,N_4869,N_4921);
nand UO_187 (O_187,N_4961,N_4993);
nand UO_188 (O_188,N_4884,N_4935);
nand UO_189 (O_189,N_4988,N_4884);
nor UO_190 (O_190,N_4925,N_4915);
nand UO_191 (O_191,N_4959,N_4881);
nor UO_192 (O_192,N_4919,N_4985);
nor UO_193 (O_193,N_4845,N_4878);
or UO_194 (O_194,N_4921,N_4994);
nor UO_195 (O_195,N_4938,N_4911);
nor UO_196 (O_196,N_4876,N_4924);
or UO_197 (O_197,N_4843,N_4889);
nor UO_198 (O_198,N_4832,N_4819);
and UO_199 (O_199,N_4860,N_4897);
nor UO_200 (O_200,N_4931,N_4982);
nor UO_201 (O_201,N_4937,N_4983);
and UO_202 (O_202,N_4858,N_4891);
nand UO_203 (O_203,N_4996,N_4931);
nand UO_204 (O_204,N_4838,N_4973);
or UO_205 (O_205,N_4838,N_4807);
or UO_206 (O_206,N_4902,N_4912);
nand UO_207 (O_207,N_4887,N_4891);
nor UO_208 (O_208,N_4865,N_4908);
or UO_209 (O_209,N_4995,N_4969);
and UO_210 (O_210,N_4849,N_4869);
and UO_211 (O_211,N_4818,N_4874);
nor UO_212 (O_212,N_4817,N_4988);
or UO_213 (O_213,N_4921,N_4898);
and UO_214 (O_214,N_4965,N_4946);
or UO_215 (O_215,N_4991,N_4827);
nor UO_216 (O_216,N_4846,N_4825);
and UO_217 (O_217,N_4887,N_4868);
nand UO_218 (O_218,N_4968,N_4958);
nor UO_219 (O_219,N_4864,N_4950);
nor UO_220 (O_220,N_4935,N_4986);
xor UO_221 (O_221,N_4846,N_4936);
and UO_222 (O_222,N_4835,N_4808);
and UO_223 (O_223,N_4915,N_4847);
or UO_224 (O_224,N_4985,N_4823);
and UO_225 (O_225,N_4898,N_4823);
and UO_226 (O_226,N_4963,N_4855);
and UO_227 (O_227,N_4806,N_4955);
and UO_228 (O_228,N_4886,N_4823);
nor UO_229 (O_229,N_4855,N_4896);
nand UO_230 (O_230,N_4878,N_4986);
nand UO_231 (O_231,N_4934,N_4840);
nor UO_232 (O_232,N_4995,N_4820);
or UO_233 (O_233,N_4888,N_4805);
and UO_234 (O_234,N_4957,N_4878);
nand UO_235 (O_235,N_4896,N_4807);
nand UO_236 (O_236,N_4960,N_4806);
and UO_237 (O_237,N_4976,N_4863);
nand UO_238 (O_238,N_4931,N_4898);
or UO_239 (O_239,N_4977,N_4912);
nor UO_240 (O_240,N_4915,N_4878);
nand UO_241 (O_241,N_4867,N_4912);
or UO_242 (O_242,N_4803,N_4962);
nor UO_243 (O_243,N_4945,N_4967);
or UO_244 (O_244,N_4821,N_4814);
nor UO_245 (O_245,N_4916,N_4987);
nand UO_246 (O_246,N_4893,N_4990);
nand UO_247 (O_247,N_4833,N_4910);
and UO_248 (O_248,N_4811,N_4854);
and UO_249 (O_249,N_4983,N_4944);
and UO_250 (O_250,N_4927,N_4893);
and UO_251 (O_251,N_4806,N_4888);
or UO_252 (O_252,N_4852,N_4907);
nor UO_253 (O_253,N_4948,N_4823);
or UO_254 (O_254,N_4946,N_4857);
or UO_255 (O_255,N_4800,N_4839);
nand UO_256 (O_256,N_4895,N_4806);
or UO_257 (O_257,N_4944,N_4928);
or UO_258 (O_258,N_4806,N_4986);
nand UO_259 (O_259,N_4892,N_4991);
nand UO_260 (O_260,N_4974,N_4820);
or UO_261 (O_261,N_4917,N_4953);
nand UO_262 (O_262,N_4910,N_4995);
and UO_263 (O_263,N_4869,N_4905);
or UO_264 (O_264,N_4936,N_4916);
nand UO_265 (O_265,N_4877,N_4838);
nand UO_266 (O_266,N_4800,N_4926);
nor UO_267 (O_267,N_4953,N_4928);
nand UO_268 (O_268,N_4993,N_4872);
xnor UO_269 (O_269,N_4833,N_4872);
nand UO_270 (O_270,N_4997,N_4996);
nand UO_271 (O_271,N_4898,N_4844);
nor UO_272 (O_272,N_4983,N_4837);
or UO_273 (O_273,N_4989,N_4877);
or UO_274 (O_274,N_4973,N_4997);
or UO_275 (O_275,N_4950,N_4955);
and UO_276 (O_276,N_4816,N_4803);
nand UO_277 (O_277,N_4811,N_4942);
nand UO_278 (O_278,N_4893,N_4997);
nor UO_279 (O_279,N_4864,N_4954);
nand UO_280 (O_280,N_4884,N_4945);
nor UO_281 (O_281,N_4975,N_4901);
and UO_282 (O_282,N_4951,N_4818);
and UO_283 (O_283,N_4957,N_4993);
nand UO_284 (O_284,N_4896,N_4861);
nand UO_285 (O_285,N_4954,N_4944);
and UO_286 (O_286,N_4856,N_4858);
or UO_287 (O_287,N_4941,N_4886);
nor UO_288 (O_288,N_4907,N_4899);
or UO_289 (O_289,N_4835,N_4825);
and UO_290 (O_290,N_4896,N_4946);
nor UO_291 (O_291,N_4989,N_4930);
or UO_292 (O_292,N_4982,N_4848);
nand UO_293 (O_293,N_4917,N_4973);
and UO_294 (O_294,N_4911,N_4985);
nor UO_295 (O_295,N_4945,N_4808);
or UO_296 (O_296,N_4895,N_4926);
and UO_297 (O_297,N_4872,N_4920);
and UO_298 (O_298,N_4932,N_4805);
or UO_299 (O_299,N_4956,N_4983);
and UO_300 (O_300,N_4987,N_4900);
nand UO_301 (O_301,N_4985,N_4877);
nor UO_302 (O_302,N_4898,N_4983);
nor UO_303 (O_303,N_4821,N_4872);
and UO_304 (O_304,N_4872,N_4912);
nor UO_305 (O_305,N_4886,N_4976);
and UO_306 (O_306,N_4902,N_4854);
nand UO_307 (O_307,N_4884,N_4833);
nor UO_308 (O_308,N_4828,N_4957);
and UO_309 (O_309,N_4892,N_4860);
or UO_310 (O_310,N_4854,N_4869);
nand UO_311 (O_311,N_4961,N_4898);
or UO_312 (O_312,N_4948,N_4972);
or UO_313 (O_313,N_4906,N_4958);
nor UO_314 (O_314,N_4915,N_4938);
nand UO_315 (O_315,N_4864,N_4889);
and UO_316 (O_316,N_4823,N_4887);
nor UO_317 (O_317,N_4934,N_4922);
nor UO_318 (O_318,N_4877,N_4930);
nand UO_319 (O_319,N_4895,N_4913);
or UO_320 (O_320,N_4877,N_4840);
and UO_321 (O_321,N_4834,N_4813);
and UO_322 (O_322,N_4912,N_4845);
nor UO_323 (O_323,N_4852,N_4969);
nand UO_324 (O_324,N_4837,N_4907);
or UO_325 (O_325,N_4989,N_4958);
or UO_326 (O_326,N_4900,N_4944);
xnor UO_327 (O_327,N_4849,N_4939);
nor UO_328 (O_328,N_4816,N_4901);
nand UO_329 (O_329,N_4950,N_4873);
or UO_330 (O_330,N_4813,N_4943);
nand UO_331 (O_331,N_4841,N_4873);
nand UO_332 (O_332,N_4815,N_4810);
nor UO_333 (O_333,N_4877,N_4862);
and UO_334 (O_334,N_4992,N_4816);
nor UO_335 (O_335,N_4825,N_4989);
nand UO_336 (O_336,N_4938,N_4834);
or UO_337 (O_337,N_4993,N_4857);
and UO_338 (O_338,N_4952,N_4949);
or UO_339 (O_339,N_4903,N_4935);
nand UO_340 (O_340,N_4872,N_4832);
nand UO_341 (O_341,N_4866,N_4886);
or UO_342 (O_342,N_4874,N_4916);
nand UO_343 (O_343,N_4983,N_4984);
nor UO_344 (O_344,N_4992,N_4864);
nand UO_345 (O_345,N_4868,N_4934);
or UO_346 (O_346,N_4868,N_4944);
or UO_347 (O_347,N_4839,N_4898);
nor UO_348 (O_348,N_4803,N_4963);
and UO_349 (O_349,N_4864,N_4875);
or UO_350 (O_350,N_4952,N_4804);
and UO_351 (O_351,N_4936,N_4845);
or UO_352 (O_352,N_4895,N_4891);
nand UO_353 (O_353,N_4945,N_4858);
xnor UO_354 (O_354,N_4933,N_4953);
nand UO_355 (O_355,N_4864,N_4828);
or UO_356 (O_356,N_4931,N_4912);
and UO_357 (O_357,N_4978,N_4825);
and UO_358 (O_358,N_4941,N_4859);
nor UO_359 (O_359,N_4904,N_4882);
nor UO_360 (O_360,N_4964,N_4931);
and UO_361 (O_361,N_4976,N_4878);
or UO_362 (O_362,N_4822,N_4925);
nand UO_363 (O_363,N_4816,N_4900);
nand UO_364 (O_364,N_4902,N_4809);
or UO_365 (O_365,N_4981,N_4852);
nor UO_366 (O_366,N_4880,N_4988);
or UO_367 (O_367,N_4828,N_4826);
nand UO_368 (O_368,N_4978,N_4967);
nor UO_369 (O_369,N_4927,N_4896);
or UO_370 (O_370,N_4923,N_4925);
nor UO_371 (O_371,N_4934,N_4948);
and UO_372 (O_372,N_4884,N_4981);
nand UO_373 (O_373,N_4807,N_4972);
or UO_374 (O_374,N_4884,N_4894);
nor UO_375 (O_375,N_4911,N_4884);
and UO_376 (O_376,N_4818,N_4836);
nand UO_377 (O_377,N_4997,N_4962);
nor UO_378 (O_378,N_4870,N_4844);
nand UO_379 (O_379,N_4908,N_4841);
nand UO_380 (O_380,N_4842,N_4948);
or UO_381 (O_381,N_4914,N_4993);
nor UO_382 (O_382,N_4934,N_4908);
nor UO_383 (O_383,N_4870,N_4979);
nor UO_384 (O_384,N_4882,N_4983);
nor UO_385 (O_385,N_4991,N_4842);
or UO_386 (O_386,N_4828,N_4825);
nand UO_387 (O_387,N_4887,N_4822);
and UO_388 (O_388,N_4881,N_4827);
nand UO_389 (O_389,N_4983,N_4835);
nand UO_390 (O_390,N_4898,N_4922);
nor UO_391 (O_391,N_4987,N_4885);
nor UO_392 (O_392,N_4941,N_4830);
xor UO_393 (O_393,N_4958,N_4827);
nand UO_394 (O_394,N_4903,N_4977);
and UO_395 (O_395,N_4991,N_4979);
nor UO_396 (O_396,N_4938,N_4888);
nand UO_397 (O_397,N_4923,N_4901);
nand UO_398 (O_398,N_4815,N_4843);
or UO_399 (O_399,N_4842,N_4932);
or UO_400 (O_400,N_4995,N_4978);
nand UO_401 (O_401,N_4859,N_4892);
nand UO_402 (O_402,N_4894,N_4975);
nor UO_403 (O_403,N_4869,N_4897);
or UO_404 (O_404,N_4809,N_4917);
nand UO_405 (O_405,N_4929,N_4956);
nor UO_406 (O_406,N_4956,N_4875);
nand UO_407 (O_407,N_4962,N_4963);
nand UO_408 (O_408,N_4995,N_4857);
or UO_409 (O_409,N_4931,N_4864);
or UO_410 (O_410,N_4809,N_4829);
or UO_411 (O_411,N_4818,N_4806);
or UO_412 (O_412,N_4931,N_4943);
and UO_413 (O_413,N_4801,N_4803);
nand UO_414 (O_414,N_4934,N_4813);
or UO_415 (O_415,N_4897,N_4854);
nand UO_416 (O_416,N_4961,N_4931);
and UO_417 (O_417,N_4812,N_4958);
and UO_418 (O_418,N_4872,N_4847);
nand UO_419 (O_419,N_4992,N_4821);
or UO_420 (O_420,N_4827,N_4937);
nor UO_421 (O_421,N_4998,N_4821);
nor UO_422 (O_422,N_4892,N_4994);
or UO_423 (O_423,N_4911,N_4867);
nand UO_424 (O_424,N_4942,N_4897);
nor UO_425 (O_425,N_4977,N_4837);
nand UO_426 (O_426,N_4802,N_4871);
nor UO_427 (O_427,N_4940,N_4851);
nor UO_428 (O_428,N_4912,N_4934);
or UO_429 (O_429,N_4884,N_4946);
nor UO_430 (O_430,N_4953,N_4900);
nor UO_431 (O_431,N_4835,N_4942);
nor UO_432 (O_432,N_4864,N_4829);
nor UO_433 (O_433,N_4882,N_4824);
or UO_434 (O_434,N_4890,N_4922);
nand UO_435 (O_435,N_4914,N_4804);
and UO_436 (O_436,N_4910,N_4876);
and UO_437 (O_437,N_4912,N_4809);
nor UO_438 (O_438,N_4882,N_4831);
nand UO_439 (O_439,N_4987,N_4892);
and UO_440 (O_440,N_4841,N_4853);
and UO_441 (O_441,N_4934,N_4985);
nand UO_442 (O_442,N_4999,N_4883);
and UO_443 (O_443,N_4925,N_4896);
nand UO_444 (O_444,N_4972,N_4965);
nand UO_445 (O_445,N_4809,N_4945);
nor UO_446 (O_446,N_4963,N_4928);
and UO_447 (O_447,N_4994,N_4841);
or UO_448 (O_448,N_4963,N_4844);
or UO_449 (O_449,N_4880,N_4937);
xnor UO_450 (O_450,N_4884,N_4919);
nor UO_451 (O_451,N_4973,N_4922);
nand UO_452 (O_452,N_4915,N_4822);
or UO_453 (O_453,N_4999,N_4990);
or UO_454 (O_454,N_4971,N_4889);
nor UO_455 (O_455,N_4938,N_4920);
nand UO_456 (O_456,N_4949,N_4968);
and UO_457 (O_457,N_4982,N_4878);
or UO_458 (O_458,N_4906,N_4945);
nand UO_459 (O_459,N_4911,N_4969);
nand UO_460 (O_460,N_4945,N_4879);
nand UO_461 (O_461,N_4959,N_4940);
nor UO_462 (O_462,N_4837,N_4887);
or UO_463 (O_463,N_4970,N_4933);
and UO_464 (O_464,N_4871,N_4981);
nor UO_465 (O_465,N_4814,N_4959);
or UO_466 (O_466,N_4988,N_4807);
and UO_467 (O_467,N_4814,N_4827);
nor UO_468 (O_468,N_4966,N_4955);
nand UO_469 (O_469,N_4882,N_4839);
and UO_470 (O_470,N_4839,N_4925);
and UO_471 (O_471,N_4915,N_4814);
nand UO_472 (O_472,N_4804,N_4866);
nand UO_473 (O_473,N_4968,N_4965);
nand UO_474 (O_474,N_4975,N_4978);
or UO_475 (O_475,N_4975,N_4939);
and UO_476 (O_476,N_4809,N_4852);
nor UO_477 (O_477,N_4897,N_4980);
or UO_478 (O_478,N_4923,N_4917);
nor UO_479 (O_479,N_4926,N_4934);
and UO_480 (O_480,N_4928,N_4923);
nand UO_481 (O_481,N_4981,N_4851);
nand UO_482 (O_482,N_4828,N_4814);
or UO_483 (O_483,N_4852,N_4913);
nand UO_484 (O_484,N_4909,N_4926);
and UO_485 (O_485,N_4852,N_4986);
and UO_486 (O_486,N_4952,N_4874);
and UO_487 (O_487,N_4942,N_4876);
nor UO_488 (O_488,N_4932,N_4870);
and UO_489 (O_489,N_4917,N_4856);
and UO_490 (O_490,N_4902,N_4818);
nor UO_491 (O_491,N_4892,N_4832);
nor UO_492 (O_492,N_4849,N_4998);
and UO_493 (O_493,N_4898,N_4944);
nand UO_494 (O_494,N_4919,N_4843);
and UO_495 (O_495,N_4876,N_4923);
nor UO_496 (O_496,N_4955,N_4967);
nor UO_497 (O_497,N_4976,N_4875);
or UO_498 (O_498,N_4862,N_4957);
nand UO_499 (O_499,N_4846,N_4969);
nand UO_500 (O_500,N_4849,N_4890);
or UO_501 (O_501,N_4940,N_4934);
nand UO_502 (O_502,N_4898,N_4977);
or UO_503 (O_503,N_4846,N_4841);
nand UO_504 (O_504,N_4846,N_4973);
nand UO_505 (O_505,N_4895,N_4842);
and UO_506 (O_506,N_4898,N_4805);
nor UO_507 (O_507,N_4999,N_4976);
and UO_508 (O_508,N_4935,N_4807);
and UO_509 (O_509,N_4889,N_4872);
nand UO_510 (O_510,N_4989,N_4955);
nor UO_511 (O_511,N_4949,N_4808);
nand UO_512 (O_512,N_4898,N_4838);
nor UO_513 (O_513,N_4945,N_4867);
nor UO_514 (O_514,N_4821,N_4948);
and UO_515 (O_515,N_4902,N_4815);
or UO_516 (O_516,N_4931,N_4880);
or UO_517 (O_517,N_4892,N_4895);
nor UO_518 (O_518,N_4997,N_4941);
nor UO_519 (O_519,N_4967,N_4904);
nand UO_520 (O_520,N_4983,N_4930);
nand UO_521 (O_521,N_4854,N_4855);
nor UO_522 (O_522,N_4866,N_4818);
or UO_523 (O_523,N_4863,N_4891);
or UO_524 (O_524,N_4829,N_4918);
nand UO_525 (O_525,N_4915,N_4842);
and UO_526 (O_526,N_4927,N_4981);
and UO_527 (O_527,N_4951,N_4819);
nor UO_528 (O_528,N_4855,N_4953);
nor UO_529 (O_529,N_4995,N_4941);
and UO_530 (O_530,N_4921,N_4993);
or UO_531 (O_531,N_4950,N_4954);
nand UO_532 (O_532,N_4949,N_4833);
and UO_533 (O_533,N_4944,N_4979);
or UO_534 (O_534,N_4805,N_4838);
nand UO_535 (O_535,N_4897,N_4883);
or UO_536 (O_536,N_4946,N_4911);
or UO_537 (O_537,N_4951,N_4804);
nand UO_538 (O_538,N_4811,N_4921);
and UO_539 (O_539,N_4878,N_4989);
nand UO_540 (O_540,N_4961,N_4984);
or UO_541 (O_541,N_4839,N_4910);
nor UO_542 (O_542,N_4926,N_4927);
nor UO_543 (O_543,N_4809,N_4909);
nor UO_544 (O_544,N_4826,N_4873);
nand UO_545 (O_545,N_4904,N_4919);
nor UO_546 (O_546,N_4813,N_4984);
nor UO_547 (O_547,N_4996,N_4885);
or UO_548 (O_548,N_4878,N_4922);
nor UO_549 (O_549,N_4924,N_4973);
nand UO_550 (O_550,N_4967,N_4983);
nand UO_551 (O_551,N_4859,N_4869);
nand UO_552 (O_552,N_4826,N_4802);
nand UO_553 (O_553,N_4964,N_4823);
or UO_554 (O_554,N_4809,N_4885);
or UO_555 (O_555,N_4998,N_4898);
nand UO_556 (O_556,N_4935,N_4848);
nor UO_557 (O_557,N_4876,N_4839);
and UO_558 (O_558,N_4939,N_4819);
nand UO_559 (O_559,N_4876,N_4960);
and UO_560 (O_560,N_4901,N_4950);
nor UO_561 (O_561,N_4941,N_4960);
or UO_562 (O_562,N_4919,N_4889);
nand UO_563 (O_563,N_4851,N_4867);
nor UO_564 (O_564,N_4817,N_4830);
and UO_565 (O_565,N_4996,N_4818);
and UO_566 (O_566,N_4813,N_4828);
or UO_567 (O_567,N_4822,N_4838);
nand UO_568 (O_568,N_4977,N_4916);
nand UO_569 (O_569,N_4936,N_4934);
and UO_570 (O_570,N_4895,N_4928);
or UO_571 (O_571,N_4874,N_4869);
or UO_572 (O_572,N_4833,N_4865);
and UO_573 (O_573,N_4917,N_4965);
nand UO_574 (O_574,N_4853,N_4833);
nor UO_575 (O_575,N_4883,N_4932);
nor UO_576 (O_576,N_4949,N_4973);
or UO_577 (O_577,N_4832,N_4959);
nor UO_578 (O_578,N_4880,N_4833);
and UO_579 (O_579,N_4852,N_4854);
and UO_580 (O_580,N_4837,N_4909);
or UO_581 (O_581,N_4920,N_4903);
and UO_582 (O_582,N_4972,N_4831);
nand UO_583 (O_583,N_4817,N_4859);
nor UO_584 (O_584,N_4939,N_4919);
or UO_585 (O_585,N_4866,N_4972);
or UO_586 (O_586,N_4969,N_4953);
nand UO_587 (O_587,N_4978,N_4817);
nor UO_588 (O_588,N_4851,N_4804);
or UO_589 (O_589,N_4995,N_4937);
nand UO_590 (O_590,N_4891,N_4964);
nor UO_591 (O_591,N_4932,N_4873);
and UO_592 (O_592,N_4980,N_4824);
and UO_593 (O_593,N_4997,N_4938);
and UO_594 (O_594,N_4922,N_4818);
nor UO_595 (O_595,N_4834,N_4823);
or UO_596 (O_596,N_4800,N_4902);
nor UO_597 (O_597,N_4918,N_4849);
nand UO_598 (O_598,N_4877,N_4938);
xnor UO_599 (O_599,N_4965,N_4983);
or UO_600 (O_600,N_4890,N_4923);
nand UO_601 (O_601,N_4971,N_4899);
nor UO_602 (O_602,N_4974,N_4962);
nand UO_603 (O_603,N_4914,N_4888);
xor UO_604 (O_604,N_4825,N_4880);
and UO_605 (O_605,N_4910,N_4838);
or UO_606 (O_606,N_4929,N_4952);
nand UO_607 (O_607,N_4899,N_4915);
nor UO_608 (O_608,N_4830,N_4828);
nand UO_609 (O_609,N_4865,N_4896);
or UO_610 (O_610,N_4858,N_4862);
and UO_611 (O_611,N_4808,N_4924);
nor UO_612 (O_612,N_4934,N_4933);
or UO_613 (O_613,N_4912,N_4964);
nor UO_614 (O_614,N_4910,N_4884);
or UO_615 (O_615,N_4859,N_4860);
or UO_616 (O_616,N_4923,N_4894);
or UO_617 (O_617,N_4899,N_4827);
and UO_618 (O_618,N_4964,N_4945);
and UO_619 (O_619,N_4835,N_4918);
or UO_620 (O_620,N_4825,N_4875);
or UO_621 (O_621,N_4955,N_4867);
nor UO_622 (O_622,N_4817,N_4964);
nand UO_623 (O_623,N_4853,N_4919);
and UO_624 (O_624,N_4971,N_4837);
and UO_625 (O_625,N_4962,N_4863);
nand UO_626 (O_626,N_4884,N_4922);
nor UO_627 (O_627,N_4900,N_4946);
nand UO_628 (O_628,N_4907,N_4921);
and UO_629 (O_629,N_4946,N_4803);
nand UO_630 (O_630,N_4818,N_4895);
and UO_631 (O_631,N_4994,N_4895);
nand UO_632 (O_632,N_4996,N_4858);
or UO_633 (O_633,N_4988,N_4932);
nand UO_634 (O_634,N_4899,N_4856);
xor UO_635 (O_635,N_4938,N_4863);
and UO_636 (O_636,N_4872,N_4981);
nor UO_637 (O_637,N_4800,N_4950);
nor UO_638 (O_638,N_4991,N_4852);
or UO_639 (O_639,N_4937,N_4878);
or UO_640 (O_640,N_4813,N_4881);
nand UO_641 (O_641,N_4957,N_4967);
nor UO_642 (O_642,N_4815,N_4842);
or UO_643 (O_643,N_4940,N_4997);
and UO_644 (O_644,N_4908,N_4890);
and UO_645 (O_645,N_4807,N_4885);
or UO_646 (O_646,N_4800,N_4975);
nand UO_647 (O_647,N_4812,N_4860);
and UO_648 (O_648,N_4812,N_4979);
nor UO_649 (O_649,N_4925,N_4867);
and UO_650 (O_650,N_4840,N_4878);
xnor UO_651 (O_651,N_4895,N_4943);
or UO_652 (O_652,N_4855,N_4812);
and UO_653 (O_653,N_4981,N_4849);
nand UO_654 (O_654,N_4803,N_4841);
nand UO_655 (O_655,N_4955,N_4920);
or UO_656 (O_656,N_4858,N_4982);
nor UO_657 (O_657,N_4899,N_4998);
nor UO_658 (O_658,N_4820,N_4952);
or UO_659 (O_659,N_4810,N_4804);
nor UO_660 (O_660,N_4947,N_4849);
or UO_661 (O_661,N_4969,N_4832);
nand UO_662 (O_662,N_4809,N_4801);
nor UO_663 (O_663,N_4930,N_4873);
nor UO_664 (O_664,N_4823,N_4982);
or UO_665 (O_665,N_4834,N_4933);
nand UO_666 (O_666,N_4941,N_4806);
and UO_667 (O_667,N_4977,N_4913);
or UO_668 (O_668,N_4887,N_4899);
or UO_669 (O_669,N_4854,N_4806);
nand UO_670 (O_670,N_4825,N_4961);
and UO_671 (O_671,N_4802,N_4954);
and UO_672 (O_672,N_4981,N_4997);
nand UO_673 (O_673,N_4873,N_4891);
and UO_674 (O_674,N_4809,N_4864);
nand UO_675 (O_675,N_4991,N_4874);
nand UO_676 (O_676,N_4893,N_4818);
nor UO_677 (O_677,N_4804,N_4832);
nand UO_678 (O_678,N_4877,N_4893);
nand UO_679 (O_679,N_4885,N_4955);
nand UO_680 (O_680,N_4912,N_4861);
and UO_681 (O_681,N_4824,N_4847);
or UO_682 (O_682,N_4915,N_4917);
and UO_683 (O_683,N_4991,N_4975);
nor UO_684 (O_684,N_4913,N_4900);
or UO_685 (O_685,N_4880,N_4949);
nand UO_686 (O_686,N_4992,N_4814);
nand UO_687 (O_687,N_4865,N_4973);
nor UO_688 (O_688,N_4860,N_4982);
and UO_689 (O_689,N_4835,N_4844);
and UO_690 (O_690,N_4809,N_4994);
nand UO_691 (O_691,N_4913,N_4924);
nand UO_692 (O_692,N_4993,N_4806);
and UO_693 (O_693,N_4941,N_4854);
or UO_694 (O_694,N_4834,N_4855);
nor UO_695 (O_695,N_4857,N_4920);
and UO_696 (O_696,N_4990,N_4891);
nand UO_697 (O_697,N_4968,N_4942);
and UO_698 (O_698,N_4951,N_4858);
nand UO_699 (O_699,N_4878,N_4914);
and UO_700 (O_700,N_4821,N_4823);
nand UO_701 (O_701,N_4999,N_4966);
nand UO_702 (O_702,N_4820,N_4814);
nand UO_703 (O_703,N_4950,N_4854);
nor UO_704 (O_704,N_4924,N_4800);
nor UO_705 (O_705,N_4913,N_4920);
and UO_706 (O_706,N_4822,N_4836);
or UO_707 (O_707,N_4826,N_4930);
nor UO_708 (O_708,N_4957,N_4812);
and UO_709 (O_709,N_4818,N_4808);
nand UO_710 (O_710,N_4954,N_4888);
nand UO_711 (O_711,N_4998,N_4890);
and UO_712 (O_712,N_4877,N_4909);
and UO_713 (O_713,N_4838,N_4837);
or UO_714 (O_714,N_4997,N_4937);
and UO_715 (O_715,N_4957,N_4832);
nor UO_716 (O_716,N_4977,N_4993);
nor UO_717 (O_717,N_4920,N_4963);
and UO_718 (O_718,N_4915,N_4937);
or UO_719 (O_719,N_4970,N_4846);
and UO_720 (O_720,N_4830,N_4989);
nand UO_721 (O_721,N_4874,N_4889);
and UO_722 (O_722,N_4919,N_4899);
nor UO_723 (O_723,N_4965,N_4844);
or UO_724 (O_724,N_4969,N_4890);
nand UO_725 (O_725,N_4948,N_4819);
nand UO_726 (O_726,N_4960,N_4977);
or UO_727 (O_727,N_4926,N_4893);
or UO_728 (O_728,N_4871,N_4900);
nor UO_729 (O_729,N_4929,N_4881);
xnor UO_730 (O_730,N_4867,N_4847);
nand UO_731 (O_731,N_4980,N_4959);
nor UO_732 (O_732,N_4911,N_4885);
nand UO_733 (O_733,N_4991,N_4832);
and UO_734 (O_734,N_4877,N_4849);
nor UO_735 (O_735,N_4806,N_4864);
or UO_736 (O_736,N_4846,N_4867);
and UO_737 (O_737,N_4932,N_4990);
nor UO_738 (O_738,N_4883,N_4875);
xor UO_739 (O_739,N_4865,N_4976);
and UO_740 (O_740,N_4929,N_4810);
or UO_741 (O_741,N_4828,N_4906);
and UO_742 (O_742,N_4995,N_4822);
or UO_743 (O_743,N_4852,N_4864);
and UO_744 (O_744,N_4815,N_4861);
or UO_745 (O_745,N_4899,N_4862);
or UO_746 (O_746,N_4907,N_4874);
nand UO_747 (O_747,N_4843,N_4994);
or UO_748 (O_748,N_4958,N_4868);
and UO_749 (O_749,N_4942,N_4855);
or UO_750 (O_750,N_4831,N_4914);
nand UO_751 (O_751,N_4867,N_4899);
or UO_752 (O_752,N_4991,N_4906);
or UO_753 (O_753,N_4931,N_4841);
or UO_754 (O_754,N_4993,N_4941);
or UO_755 (O_755,N_4883,N_4910);
nand UO_756 (O_756,N_4941,N_4977);
or UO_757 (O_757,N_4970,N_4952);
nand UO_758 (O_758,N_4874,N_4891);
or UO_759 (O_759,N_4838,N_4841);
nand UO_760 (O_760,N_4820,N_4861);
nand UO_761 (O_761,N_4921,N_4902);
nand UO_762 (O_762,N_4908,N_4822);
nand UO_763 (O_763,N_4948,N_4844);
or UO_764 (O_764,N_4828,N_4904);
and UO_765 (O_765,N_4959,N_4828);
or UO_766 (O_766,N_4843,N_4893);
nor UO_767 (O_767,N_4991,N_4848);
and UO_768 (O_768,N_4970,N_4913);
and UO_769 (O_769,N_4992,N_4918);
or UO_770 (O_770,N_4950,N_4890);
or UO_771 (O_771,N_4908,N_4967);
and UO_772 (O_772,N_4905,N_4814);
and UO_773 (O_773,N_4914,N_4982);
nand UO_774 (O_774,N_4829,N_4986);
nand UO_775 (O_775,N_4995,N_4855);
and UO_776 (O_776,N_4802,N_4909);
or UO_777 (O_777,N_4896,N_4994);
nor UO_778 (O_778,N_4966,N_4982);
and UO_779 (O_779,N_4847,N_4814);
and UO_780 (O_780,N_4859,N_4896);
and UO_781 (O_781,N_4875,N_4896);
and UO_782 (O_782,N_4888,N_4922);
nor UO_783 (O_783,N_4829,N_4823);
or UO_784 (O_784,N_4921,N_4884);
nor UO_785 (O_785,N_4973,N_4968);
or UO_786 (O_786,N_4939,N_4861);
nand UO_787 (O_787,N_4920,N_4810);
or UO_788 (O_788,N_4977,N_4887);
nand UO_789 (O_789,N_4826,N_4810);
and UO_790 (O_790,N_4873,N_4803);
nand UO_791 (O_791,N_4809,N_4869);
and UO_792 (O_792,N_4812,N_4946);
nand UO_793 (O_793,N_4891,N_4909);
nand UO_794 (O_794,N_4897,N_4983);
nor UO_795 (O_795,N_4864,N_4961);
nor UO_796 (O_796,N_4804,N_4886);
or UO_797 (O_797,N_4812,N_4927);
or UO_798 (O_798,N_4941,N_4934);
nand UO_799 (O_799,N_4809,N_4993);
or UO_800 (O_800,N_4906,N_4964);
and UO_801 (O_801,N_4839,N_4874);
nor UO_802 (O_802,N_4873,N_4937);
or UO_803 (O_803,N_4965,N_4897);
or UO_804 (O_804,N_4818,N_4979);
nor UO_805 (O_805,N_4833,N_4903);
nand UO_806 (O_806,N_4824,N_4994);
nor UO_807 (O_807,N_4954,N_4969);
or UO_808 (O_808,N_4868,N_4876);
and UO_809 (O_809,N_4885,N_4966);
and UO_810 (O_810,N_4918,N_4865);
or UO_811 (O_811,N_4921,N_4990);
or UO_812 (O_812,N_4877,N_4932);
nor UO_813 (O_813,N_4857,N_4854);
and UO_814 (O_814,N_4883,N_4848);
xor UO_815 (O_815,N_4863,N_4903);
nor UO_816 (O_816,N_4846,N_4942);
nor UO_817 (O_817,N_4906,N_4928);
and UO_818 (O_818,N_4921,N_4931);
nor UO_819 (O_819,N_4952,N_4835);
or UO_820 (O_820,N_4815,N_4862);
nor UO_821 (O_821,N_4823,N_4814);
and UO_822 (O_822,N_4877,N_4828);
nor UO_823 (O_823,N_4854,N_4943);
nor UO_824 (O_824,N_4868,N_4816);
or UO_825 (O_825,N_4820,N_4834);
nor UO_826 (O_826,N_4833,N_4907);
or UO_827 (O_827,N_4812,N_4930);
nand UO_828 (O_828,N_4996,N_4995);
and UO_829 (O_829,N_4845,N_4840);
nand UO_830 (O_830,N_4830,N_4962);
and UO_831 (O_831,N_4864,N_4863);
or UO_832 (O_832,N_4862,N_4956);
nor UO_833 (O_833,N_4809,N_4805);
or UO_834 (O_834,N_4881,N_4960);
or UO_835 (O_835,N_4909,N_4804);
nor UO_836 (O_836,N_4978,N_4918);
or UO_837 (O_837,N_4886,N_4929);
nand UO_838 (O_838,N_4914,N_4903);
xor UO_839 (O_839,N_4835,N_4852);
nand UO_840 (O_840,N_4887,N_4856);
and UO_841 (O_841,N_4950,N_4851);
or UO_842 (O_842,N_4969,N_4807);
nand UO_843 (O_843,N_4872,N_4972);
and UO_844 (O_844,N_4896,N_4868);
nor UO_845 (O_845,N_4889,N_4827);
nor UO_846 (O_846,N_4881,N_4987);
and UO_847 (O_847,N_4821,N_4904);
and UO_848 (O_848,N_4950,N_4912);
nor UO_849 (O_849,N_4954,N_4996);
or UO_850 (O_850,N_4988,N_4899);
nor UO_851 (O_851,N_4995,N_4815);
or UO_852 (O_852,N_4902,N_4882);
nand UO_853 (O_853,N_4856,N_4955);
or UO_854 (O_854,N_4933,N_4812);
and UO_855 (O_855,N_4939,N_4979);
nand UO_856 (O_856,N_4929,N_4995);
and UO_857 (O_857,N_4957,N_4955);
nor UO_858 (O_858,N_4839,N_4920);
nor UO_859 (O_859,N_4852,N_4966);
and UO_860 (O_860,N_4956,N_4874);
or UO_861 (O_861,N_4941,N_4974);
nor UO_862 (O_862,N_4813,N_4962);
nand UO_863 (O_863,N_4976,N_4818);
nand UO_864 (O_864,N_4925,N_4984);
nor UO_865 (O_865,N_4870,N_4818);
nand UO_866 (O_866,N_4937,N_4930);
or UO_867 (O_867,N_4897,N_4977);
and UO_868 (O_868,N_4862,N_4977);
or UO_869 (O_869,N_4871,N_4991);
nor UO_870 (O_870,N_4839,N_4939);
nor UO_871 (O_871,N_4966,N_4870);
nand UO_872 (O_872,N_4839,N_4973);
xor UO_873 (O_873,N_4921,N_4984);
nand UO_874 (O_874,N_4919,N_4990);
nand UO_875 (O_875,N_4818,N_4877);
nor UO_876 (O_876,N_4991,N_4928);
and UO_877 (O_877,N_4993,N_4901);
xor UO_878 (O_878,N_4888,N_4813);
nor UO_879 (O_879,N_4863,N_4843);
nor UO_880 (O_880,N_4833,N_4905);
nand UO_881 (O_881,N_4916,N_4820);
or UO_882 (O_882,N_4973,N_4836);
or UO_883 (O_883,N_4931,N_4965);
nor UO_884 (O_884,N_4929,N_4818);
nor UO_885 (O_885,N_4934,N_4846);
and UO_886 (O_886,N_4949,N_4936);
nand UO_887 (O_887,N_4902,N_4820);
or UO_888 (O_888,N_4855,N_4986);
nand UO_889 (O_889,N_4971,N_4967);
nor UO_890 (O_890,N_4959,N_4824);
nor UO_891 (O_891,N_4982,N_4938);
or UO_892 (O_892,N_4876,N_4881);
or UO_893 (O_893,N_4978,N_4988);
or UO_894 (O_894,N_4979,N_4842);
nor UO_895 (O_895,N_4843,N_4804);
nor UO_896 (O_896,N_4998,N_4973);
or UO_897 (O_897,N_4853,N_4889);
nor UO_898 (O_898,N_4807,N_4889);
nor UO_899 (O_899,N_4933,N_4975);
and UO_900 (O_900,N_4959,N_4902);
nand UO_901 (O_901,N_4925,N_4973);
nand UO_902 (O_902,N_4910,N_4971);
nor UO_903 (O_903,N_4873,N_4983);
nand UO_904 (O_904,N_4975,N_4993);
or UO_905 (O_905,N_4858,N_4937);
nor UO_906 (O_906,N_4953,N_4960);
nor UO_907 (O_907,N_4800,N_4923);
nand UO_908 (O_908,N_4974,N_4967);
and UO_909 (O_909,N_4910,N_4894);
and UO_910 (O_910,N_4852,N_4989);
or UO_911 (O_911,N_4817,N_4967);
or UO_912 (O_912,N_4853,N_4900);
nor UO_913 (O_913,N_4850,N_4830);
or UO_914 (O_914,N_4968,N_4840);
nor UO_915 (O_915,N_4906,N_4837);
and UO_916 (O_916,N_4970,N_4955);
or UO_917 (O_917,N_4953,N_4902);
and UO_918 (O_918,N_4857,N_4985);
nand UO_919 (O_919,N_4958,N_4809);
nor UO_920 (O_920,N_4852,N_4970);
and UO_921 (O_921,N_4823,N_4921);
or UO_922 (O_922,N_4842,N_4968);
and UO_923 (O_923,N_4846,N_4855);
or UO_924 (O_924,N_4838,N_4824);
nand UO_925 (O_925,N_4943,N_4879);
and UO_926 (O_926,N_4973,N_4875);
or UO_927 (O_927,N_4800,N_4909);
and UO_928 (O_928,N_4935,N_4882);
and UO_929 (O_929,N_4824,N_4879);
nor UO_930 (O_930,N_4978,N_4925);
and UO_931 (O_931,N_4844,N_4856);
nand UO_932 (O_932,N_4884,N_4930);
nor UO_933 (O_933,N_4802,N_4897);
and UO_934 (O_934,N_4851,N_4912);
and UO_935 (O_935,N_4853,N_4847);
or UO_936 (O_936,N_4960,N_4831);
or UO_937 (O_937,N_4867,N_4900);
and UO_938 (O_938,N_4877,N_4806);
or UO_939 (O_939,N_4993,N_4976);
nor UO_940 (O_940,N_4853,N_4918);
nor UO_941 (O_941,N_4970,N_4882);
nor UO_942 (O_942,N_4827,N_4960);
or UO_943 (O_943,N_4980,N_4866);
xor UO_944 (O_944,N_4836,N_4926);
and UO_945 (O_945,N_4958,N_4911);
and UO_946 (O_946,N_4850,N_4954);
nand UO_947 (O_947,N_4945,N_4847);
nand UO_948 (O_948,N_4979,N_4966);
and UO_949 (O_949,N_4900,N_4801);
and UO_950 (O_950,N_4804,N_4893);
nor UO_951 (O_951,N_4815,N_4811);
or UO_952 (O_952,N_4837,N_4856);
and UO_953 (O_953,N_4887,N_4911);
or UO_954 (O_954,N_4849,N_4961);
or UO_955 (O_955,N_4824,N_4881);
xnor UO_956 (O_956,N_4886,N_4919);
and UO_957 (O_957,N_4953,N_4914);
xnor UO_958 (O_958,N_4904,N_4986);
or UO_959 (O_959,N_4827,N_4879);
nand UO_960 (O_960,N_4858,N_4962);
or UO_961 (O_961,N_4926,N_4813);
nor UO_962 (O_962,N_4868,N_4904);
nor UO_963 (O_963,N_4815,N_4978);
nor UO_964 (O_964,N_4901,N_4933);
nor UO_965 (O_965,N_4877,N_4897);
nor UO_966 (O_966,N_4985,N_4832);
and UO_967 (O_967,N_4974,N_4997);
nor UO_968 (O_968,N_4884,N_4862);
nand UO_969 (O_969,N_4838,N_4980);
nand UO_970 (O_970,N_4945,N_4929);
nor UO_971 (O_971,N_4823,N_4962);
nand UO_972 (O_972,N_4974,N_4943);
nor UO_973 (O_973,N_4996,N_4963);
nor UO_974 (O_974,N_4888,N_4871);
nand UO_975 (O_975,N_4880,N_4812);
nand UO_976 (O_976,N_4984,N_4903);
nand UO_977 (O_977,N_4886,N_4850);
nor UO_978 (O_978,N_4964,N_4875);
or UO_979 (O_979,N_4948,N_4879);
or UO_980 (O_980,N_4882,N_4821);
nor UO_981 (O_981,N_4861,N_4987);
and UO_982 (O_982,N_4982,N_4888);
or UO_983 (O_983,N_4875,N_4966);
or UO_984 (O_984,N_4803,N_4819);
nor UO_985 (O_985,N_4972,N_4806);
nand UO_986 (O_986,N_4919,N_4891);
nor UO_987 (O_987,N_4934,N_4857);
nand UO_988 (O_988,N_4938,N_4864);
nand UO_989 (O_989,N_4805,N_4886);
nand UO_990 (O_990,N_4933,N_4836);
nor UO_991 (O_991,N_4910,N_4855);
or UO_992 (O_992,N_4873,N_4924);
nand UO_993 (O_993,N_4985,N_4895);
and UO_994 (O_994,N_4883,N_4969);
nand UO_995 (O_995,N_4940,N_4870);
nor UO_996 (O_996,N_4807,N_4921);
nor UO_997 (O_997,N_4960,N_4898);
nor UO_998 (O_998,N_4970,N_4827);
and UO_999 (O_999,N_4830,N_4981);
endmodule