module basic_2500_25000_3000_5_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1862,In_2312);
and U1 (N_1,In_829,In_2343);
nand U2 (N_2,In_1970,In_1279);
or U3 (N_3,In_1268,In_1047);
nand U4 (N_4,In_1703,In_2004);
nor U5 (N_5,In_2472,In_91);
nand U6 (N_6,In_533,In_700);
xnor U7 (N_7,In_1372,In_932);
nand U8 (N_8,In_534,In_1820);
or U9 (N_9,In_980,In_181);
nor U10 (N_10,In_163,In_1272);
nand U11 (N_11,In_2393,In_504);
and U12 (N_12,In_1169,In_742);
nor U13 (N_13,In_1219,In_638);
and U14 (N_14,In_253,In_1225);
nand U15 (N_15,In_2308,In_410);
or U16 (N_16,In_2463,In_2261);
and U17 (N_17,In_218,In_1076);
or U18 (N_18,In_654,In_1043);
nand U19 (N_19,In_701,In_1828);
nand U20 (N_20,In_842,In_1863);
or U21 (N_21,In_2056,In_1356);
and U22 (N_22,In_1082,In_399);
or U23 (N_23,In_75,In_1378);
nand U24 (N_24,In_79,In_887);
or U25 (N_25,In_976,In_1083);
nand U26 (N_26,In_865,In_748);
nand U27 (N_27,In_59,In_840);
or U28 (N_28,In_795,In_585);
nor U29 (N_29,In_2286,In_1261);
or U30 (N_30,In_1244,In_2008);
or U31 (N_31,In_1871,In_1445);
nor U32 (N_32,In_1097,In_1945);
nor U33 (N_33,In_1724,In_1202);
and U34 (N_34,In_907,In_150);
nand U35 (N_35,In_867,In_1402);
nand U36 (N_36,In_303,In_162);
and U37 (N_37,In_906,In_728);
nor U38 (N_38,In_2371,In_1699);
and U39 (N_39,In_1514,In_1494);
or U40 (N_40,In_581,In_167);
and U41 (N_41,In_2024,In_1885);
nor U42 (N_42,In_1123,In_1053);
nor U43 (N_43,In_1938,In_1067);
or U44 (N_44,In_1913,In_1957);
and U45 (N_45,In_1236,In_1347);
nor U46 (N_46,In_1231,In_171);
and U47 (N_47,In_1119,In_1636);
nor U48 (N_48,In_506,In_712);
and U49 (N_49,In_574,In_1768);
nor U50 (N_50,In_1249,In_514);
or U51 (N_51,In_995,In_1673);
nor U52 (N_52,In_815,In_622);
or U53 (N_53,In_1095,In_1411);
xor U54 (N_54,In_1031,In_1630);
or U55 (N_55,In_389,In_1438);
or U56 (N_56,In_1847,In_2404);
and U57 (N_57,In_1432,In_10);
or U58 (N_58,In_1985,In_1477);
nor U59 (N_59,In_119,In_1404);
or U60 (N_60,In_1996,In_151);
and U61 (N_61,In_1105,In_1973);
nand U62 (N_62,In_1367,In_838);
nand U63 (N_63,In_407,In_1966);
nand U64 (N_64,In_615,In_1647);
and U65 (N_65,In_612,In_1830);
or U66 (N_66,In_1625,In_108);
nor U67 (N_67,In_1616,In_913);
nand U68 (N_68,In_885,In_383);
and U69 (N_69,In_1998,In_785);
nor U70 (N_70,In_336,In_991);
nor U71 (N_71,In_403,In_99);
or U72 (N_72,In_627,In_244);
nor U73 (N_73,In_1992,In_1653);
nand U74 (N_74,In_1375,In_1574);
or U75 (N_75,In_341,In_539);
nor U76 (N_76,In_2122,In_856);
and U77 (N_77,In_1812,In_1947);
or U78 (N_78,In_1604,In_43);
nor U79 (N_79,In_659,In_203);
nand U80 (N_80,In_1393,In_1486);
nand U81 (N_81,In_1924,In_481);
nand U82 (N_82,In_1192,In_957);
nand U83 (N_83,In_1997,In_454);
or U84 (N_84,In_1296,In_823);
nor U85 (N_85,In_1901,In_740);
nand U86 (N_86,In_1739,In_1104);
or U87 (N_87,In_1805,In_1183);
nand U88 (N_88,In_1191,In_1746);
nor U89 (N_89,In_1651,In_357);
nand U90 (N_90,In_1790,In_625);
nand U91 (N_91,In_2278,In_21);
nand U92 (N_92,In_640,In_658);
or U93 (N_93,In_187,In_1908);
nor U94 (N_94,In_146,In_122);
and U95 (N_95,In_1446,In_1172);
nor U96 (N_96,In_1304,In_1714);
nor U97 (N_97,In_487,In_1029);
nor U98 (N_98,In_2387,In_1363);
or U99 (N_99,In_77,In_2093);
or U100 (N_100,In_1688,In_2285);
nand U101 (N_101,In_2473,In_697);
nand U102 (N_102,In_1388,In_734);
and U103 (N_103,In_1070,In_882);
or U104 (N_104,In_2271,In_193);
and U105 (N_105,In_321,In_2465);
nor U106 (N_106,In_1121,In_918);
nand U107 (N_107,In_880,In_385);
xnor U108 (N_108,In_1934,In_2183);
nand U109 (N_109,In_62,In_103);
nor U110 (N_110,In_820,In_1407);
nor U111 (N_111,In_1107,In_1059);
nand U112 (N_112,In_962,In_1748);
nand U113 (N_113,In_212,In_1253);
or U114 (N_114,In_886,In_1526);
and U115 (N_115,In_183,In_808);
and U116 (N_116,In_1461,In_137);
or U117 (N_117,In_19,In_491);
or U118 (N_118,In_1112,In_1118);
or U119 (N_119,In_173,In_1283);
nor U120 (N_120,In_1403,In_1211);
nand U121 (N_121,In_1979,In_2291);
nand U122 (N_122,In_944,In_1081);
or U123 (N_123,In_2375,In_1889);
or U124 (N_124,In_1334,In_883);
and U125 (N_125,In_617,In_1051);
nor U126 (N_126,In_2200,In_2059);
or U127 (N_127,In_1516,In_2323);
or U128 (N_128,In_161,In_1437);
nor U129 (N_129,In_2170,In_170);
and U130 (N_130,In_1685,In_717);
nor U131 (N_131,In_492,In_2451);
and U132 (N_132,In_607,In_1672);
nand U133 (N_133,In_1556,In_25);
nand U134 (N_134,In_943,In_1116);
nor U135 (N_135,In_2172,In_667);
nor U136 (N_136,In_1887,In_1449);
nand U137 (N_137,In_1852,In_1840);
nand U138 (N_138,In_825,In_806);
and U139 (N_139,In_1565,In_1274);
and U140 (N_140,In_190,In_1988);
and U141 (N_141,In_427,In_1864);
and U142 (N_142,In_1501,In_873);
and U143 (N_143,In_1386,In_1771);
and U144 (N_144,In_1351,In_2042);
or U145 (N_145,In_32,In_971);
and U146 (N_146,In_395,In_778);
nand U147 (N_147,In_993,In_210);
nor U148 (N_148,In_1464,In_1511);
nor U149 (N_149,In_953,In_1902);
or U150 (N_150,In_816,In_2374);
nor U151 (N_151,In_444,In_774);
and U152 (N_152,In_1854,In_1897);
nor U153 (N_153,In_2319,In_269);
nand U154 (N_154,In_2058,In_763);
and U155 (N_155,In_1057,In_165);
nand U156 (N_156,In_1725,In_920);
and U157 (N_157,In_580,In_1727);
or U158 (N_158,In_1346,In_18);
nor U159 (N_159,In_1163,In_1282);
nand U160 (N_160,In_26,In_1472);
nand U161 (N_161,In_827,In_1178);
or U162 (N_162,In_1972,In_1454);
and U163 (N_163,In_2303,In_1702);
or U164 (N_164,In_144,In_967);
or U165 (N_165,In_23,In_339);
and U166 (N_166,In_1350,In_613);
or U167 (N_167,In_546,In_483);
or U168 (N_168,In_1222,In_392);
and U169 (N_169,In_1308,In_922);
nor U170 (N_170,In_1595,In_587);
nand U171 (N_171,In_2203,In_1007);
nor U172 (N_172,In_2388,In_850);
xnor U173 (N_173,In_273,In_837);
and U174 (N_174,In_797,In_1552);
nor U175 (N_175,In_316,In_1482);
nor U176 (N_176,In_2158,In_952);
and U177 (N_177,In_1181,In_964);
and U178 (N_178,In_1553,In_2082);
and U179 (N_179,In_1716,In_1678);
or U180 (N_180,In_1475,In_1692);
or U181 (N_181,In_2031,In_2256);
and U182 (N_182,In_2495,In_985);
or U183 (N_183,In_2259,In_1220);
nand U184 (N_184,In_1020,In_1519);
or U185 (N_185,In_764,In_240);
nor U186 (N_186,In_1661,In_1488);
or U187 (N_187,In_1013,In_1876);
or U188 (N_188,In_2266,In_2152);
and U189 (N_189,In_1370,In_236);
nand U190 (N_190,In_1712,In_1755);
nand U191 (N_191,In_1648,In_156);
and U192 (N_192,In_229,In_1017);
nor U193 (N_193,In_756,In_412);
or U194 (N_194,In_52,In_1807);
nand U195 (N_195,In_9,In_1958);
nor U196 (N_196,In_2089,In_1596);
nand U197 (N_197,In_1237,In_1612);
or U198 (N_198,In_1072,In_180);
and U199 (N_199,In_1615,In_2108);
nor U200 (N_200,In_276,In_1138);
and U201 (N_201,In_1750,In_1117);
nor U202 (N_202,In_1196,In_2146);
or U203 (N_203,In_1773,In_1058);
or U204 (N_204,In_503,In_1780);
or U205 (N_205,In_300,In_1187);
nor U206 (N_206,In_2477,In_2168);
nor U207 (N_207,In_768,In_416);
nand U208 (N_208,In_682,In_1522);
or U209 (N_209,In_490,In_364);
nor U210 (N_210,In_259,In_543);
or U211 (N_211,In_1396,In_458);
xnor U212 (N_212,In_2228,In_46);
nand U213 (N_213,In_349,In_474);
nor U214 (N_214,In_2033,In_552);
nor U215 (N_215,In_1823,In_1336);
nand U216 (N_216,In_1460,In_716);
nand U217 (N_217,In_2432,In_1868);
or U218 (N_218,In_589,In_1280);
nor U219 (N_219,In_2479,In_2464);
nand U220 (N_220,In_2444,In_555);
nor U221 (N_221,In_1663,In_2297);
or U222 (N_222,In_2178,In_1558);
and U223 (N_223,In_1627,In_1801);
or U224 (N_224,In_802,In_1968);
and U225 (N_225,In_1009,In_1817);
nor U226 (N_226,In_2166,In_1259);
nand U227 (N_227,In_2412,In_1867);
and U228 (N_228,In_1835,In_595);
nor U229 (N_229,In_598,In_2358);
and U230 (N_230,In_2173,In_1713);
or U231 (N_231,In_759,In_833);
nor U232 (N_232,In_2486,In_948);
nand U233 (N_233,In_1306,In_1424);
nor U234 (N_234,In_2099,In_2318);
nor U235 (N_235,In_2083,In_94);
or U236 (N_236,In_297,In_1332);
and U237 (N_237,In_1434,In_1664);
and U238 (N_238,In_854,In_354);
xor U239 (N_239,In_689,In_675);
nand U240 (N_240,In_377,In_1641);
nand U241 (N_241,In_1148,In_990);
nor U242 (N_242,In_2287,In_337);
nand U243 (N_243,In_1503,In_835);
xor U244 (N_244,In_649,In_147);
and U245 (N_245,In_1448,In_396);
or U246 (N_246,In_211,In_5);
or U247 (N_247,In_423,In_636);
nor U248 (N_248,In_2025,In_1177);
or U249 (N_249,In_1419,In_1677);
or U250 (N_250,In_2369,In_968);
and U251 (N_251,In_2362,In_1850);
nand U252 (N_252,In_982,In_1915);
nor U253 (N_253,In_1839,In_2013);
or U254 (N_254,In_1610,In_16);
or U255 (N_255,In_2391,In_2225);
or U256 (N_256,In_1459,In_1048);
nor U257 (N_257,In_2484,In_1502);
and U258 (N_258,In_2453,In_1340);
and U259 (N_259,In_558,In_2014);
xnor U260 (N_260,In_1759,In_447);
nor U261 (N_261,In_893,In_745);
or U262 (N_262,In_476,In_2067);
or U263 (N_263,In_2481,In_37);
or U264 (N_264,In_1577,In_2437);
and U265 (N_265,In_1654,In_1490);
and U266 (N_266,In_1978,In_868);
and U267 (N_267,In_2154,In_2100);
nor U268 (N_268,In_934,In_201);
or U269 (N_269,In_1395,In_910);
and U270 (N_270,In_2368,In_1668);
nand U271 (N_271,In_573,In_2068);
and U272 (N_272,In_2349,In_338);
or U273 (N_273,In_2466,In_237);
and U274 (N_274,In_1421,In_2066);
and U275 (N_275,In_1621,In_584);
nor U276 (N_276,In_1320,In_781);
and U277 (N_277,In_2034,In_1015);
nor U278 (N_278,In_1158,In_2348);
nor U279 (N_279,In_2026,In_443);
or U280 (N_280,In_254,In_1783);
nand U281 (N_281,In_2137,In_2037);
nor U282 (N_282,In_1130,In_687);
xnor U283 (N_283,In_1870,In_148);
and U284 (N_284,In_1906,In_790);
and U285 (N_285,In_1377,In_252);
nor U286 (N_286,In_286,In_1731);
nand U287 (N_287,In_1089,In_2499);
xnor U288 (N_288,In_2351,In_1480);
and U289 (N_289,In_448,In_2143);
nand U290 (N_290,In_1929,In_1032);
nand U291 (N_291,In_393,In_2050);
nor U292 (N_292,In_2101,In_22);
nor U293 (N_293,In_1137,In_1646);
nand U294 (N_294,In_1226,In_683);
and U295 (N_295,In_164,In_1715);
and U296 (N_296,In_1875,In_1756);
and U297 (N_297,In_451,In_859);
nand U298 (N_298,In_2195,In_2132);
nor U299 (N_299,In_676,In_1300);
nand U300 (N_300,In_738,In_688);
nor U301 (N_301,In_54,In_516);
nand U302 (N_302,In_60,In_2241);
and U303 (N_303,In_11,In_2096);
nand U304 (N_304,In_1791,In_1085);
nand U305 (N_305,In_2482,In_2324);
and U306 (N_306,In_417,In_757);
or U307 (N_307,In_561,In_1528);
and U308 (N_308,In_846,In_1415);
nor U309 (N_309,In_1623,In_694);
nand U310 (N_310,In_564,In_2142);
nand U311 (N_311,In_2447,In_1951);
nor U312 (N_312,In_1242,In_1591);
or U313 (N_313,In_228,In_769);
xnor U314 (N_314,In_13,In_2065);
and U315 (N_315,In_1605,In_549);
nand U316 (N_316,In_1287,In_557);
nor U317 (N_317,In_196,In_1310);
and U318 (N_318,In_569,In_1986);
nor U319 (N_319,In_360,In_2114);
or U320 (N_320,In_851,In_1977);
nor U321 (N_321,In_308,In_1872);
nand U322 (N_322,In_1321,In_292);
nand U323 (N_323,In_1569,In_1185);
or U324 (N_324,In_2376,In_2251);
and U325 (N_325,In_361,In_974);
nand U326 (N_326,In_586,In_1174);
or U327 (N_327,In_1933,In_1786);
nor U328 (N_328,In_2456,In_1618);
nand U329 (N_329,In_1041,In_1946);
and U330 (N_330,In_789,In_2182);
nand U331 (N_331,In_941,In_325);
nand U332 (N_332,In_1819,In_1531);
or U333 (N_333,In_705,In_2347);
and U334 (N_334,In_1439,In_2010);
or U335 (N_335,In_335,In_27);
or U336 (N_336,In_2053,In_55);
and U337 (N_337,In_965,In_1371);
nand U338 (N_338,In_320,In_1262);
nor U339 (N_339,In_332,In_42);
nand U340 (N_340,In_263,In_2274);
and U341 (N_341,In_1002,In_257);
and U342 (N_342,In_2264,In_1698);
nand U343 (N_343,In_1124,In_2207);
nor U344 (N_344,In_695,In_2433);
or U345 (N_345,In_1940,In_1787);
or U346 (N_346,In_1962,In_1281);
nor U347 (N_347,In_1701,In_1423);
or U348 (N_348,In_1617,In_1145);
nor U349 (N_349,In_1291,In_550);
and U350 (N_350,In_691,In_1642);
nand U351 (N_351,In_1861,In_1066);
nor U352 (N_352,In_2129,In_50);
and U353 (N_353,In_2080,In_2382);
nor U354 (N_354,In_594,In_281);
nand U355 (N_355,In_2430,In_352);
nor U356 (N_356,In_1657,In_57);
xnor U357 (N_357,In_929,In_926);
and U358 (N_358,In_507,In_2284);
or U359 (N_359,In_579,In_2314);
nand U360 (N_360,In_2107,In_1110);
nor U361 (N_361,In_1349,In_810);
or U362 (N_362,In_1252,In_1853);
and U363 (N_363,In_430,In_73);
nand U364 (N_364,In_264,In_853);
nand U365 (N_365,In_2140,In_765);
and U366 (N_366,In_1343,In_665);
nor U367 (N_367,In_2396,In_2153);
and U368 (N_368,In_1011,In_1718);
or U369 (N_369,In_2325,In_895);
and U370 (N_370,In_2036,In_442);
or U371 (N_371,In_1302,In_309);
xor U372 (N_372,In_809,In_1721);
and U373 (N_373,In_1399,In_729);
or U374 (N_374,In_609,In_1880);
xor U375 (N_375,In_736,In_544);
nor U376 (N_376,In_459,In_787);
or U377 (N_377,In_2061,In_1949);
or U378 (N_378,In_1907,In_1342);
and U379 (N_379,In_502,In_235);
nand U380 (N_380,In_317,In_1644);
nor U381 (N_381,In_1587,In_1818);
or U382 (N_382,In_1967,In_1665);
nand U383 (N_383,In_2389,In_551);
or U384 (N_384,In_2454,In_1257);
and U385 (N_385,In_1458,In_1981);
and U386 (N_386,In_1903,In_1042);
and U387 (N_387,In_1214,In_1436);
and U388 (N_388,In_285,In_1675);
or U389 (N_389,In_2399,In_1766);
or U390 (N_390,In_1157,In_2191);
nor U391 (N_391,In_2141,In_2119);
xor U392 (N_392,In_2206,In_2462);
and U393 (N_393,In_1843,In_1781);
nor U394 (N_394,In_696,In_2248);
and U395 (N_395,In_1851,In_2102);
and U396 (N_396,In_1294,In_29);
and U397 (N_397,In_855,In_1418);
nor U398 (N_398,In_2192,In_1330);
nand U399 (N_399,In_637,In_58);
and U400 (N_400,In_2478,In_1896);
nor U401 (N_401,In_256,In_440);
or U402 (N_402,In_128,In_1021);
nor U403 (N_403,In_132,In_1652);
nand U404 (N_404,In_206,In_1466);
or U405 (N_405,In_1373,In_2356);
nand U406 (N_406,In_1659,In_1129);
or U407 (N_407,In_1210,In_470);
and U408 (N_408,In_1570,In_1928);
or U409 (N_409,In_1131,In_1295);
or U410 (N_410,In_266,In_347);
nand U411 (N_411,In_2474,In_784);
nor U412 (N_412,In_426,In_53);
or U413 (N_413,In_817,In_1753);
nand U414 (N_414,In_525,In_279);
nand U415 (N_415,In_274,In_1729);
or U416 (N_416,In_110,In_1133);
or U417 (N_417,In_2295,In_678);
and U418 (N_418,In_106,In_1666);
nand U419 (N_419,In_475,In_1821);
and U420 (N_420,In_1775,In_599);
or U421 (N_421,In_889,In_523);
nand U422 (N_422,In_74,In_1735);
and U423 (N_423,In_2350,In_1926);
or U424 (N_424,In_1856,In_105);
nand U425 (N_425,In_2155,In_1298);
or U426 (N_426,In_2435,In_973);
nand U427 (N_427,In_956,In_391);
and U428 (N_428,In_1892,In_246);
and U429 (N_429,In_1882,In_2103);
nand U430 (N_430,In_63,In_1520);
nor U431 (N_431,In_937,In_1802);
or U432 (N_432,In_2424,In_2339);
or U433 (N_433,In_639,In_663);
nand U434 (N_434,In_1691,In_2431);
xor U435 (N_435,In_2395,In_780);
nor U436 (N_436,In_1171,In_1881);
xor U437 (N_437,In_1359,In_2125);
and U438 (N_438,In_450,In_1662);
nand U439 (N_439,In_1778,In_1782);
nor U440 (N_440,In_2233,In_578);
nor U441 (N_441,In_348,In_1246);
nand U442 (N_442,In_872,In_2230);
and U443 (N_443,In_1136,In_2260);
nor U444 (N_444,In_786,In_2313);
nand U445 (N_445,In_623,In_725);
or U446 (N_446,In_2097,In_2227);
nand U447 (N_447,In_2123,In_511);
nor U448 (N_448,In_901,In_2379);
or U449 (N_449,In_2072,In_1722);
nor U450 (N_450,In_2449,In_1173);
nor U451 (N_451,In_1927,In_1071);
nor U452 (N_452,In_2184,In_1710);
and U453 (N_453,In_2029,In_1200);
nand U454 (N_454,In_31,In_1601);
nand U455 (N_455,In_1877,In_2222);
and U456 (N_456,In_730,In_2087);
or U457 (N_457,In_293,In_1602);
nor U458 (N_458,In_1555,In_2151);
or U459 (N_459,In_81,In_1044);
nand U460 (N_460,In_255,In_722);
nand U461 (N_461,In_102,In_2334);
nor U462 (N_462,In_126,In_44);
and U463 (N_463,In_1470,In_1792);
nor U464 (N_464,In_1626,In_1760);
nand U465 (N_465,In_1498,In_1062);
and U466 (N_466,In_1777,In_2115);
or U467 (N_467,In_2232,In_1218);
or U468 (N_468,In_397,In_2112);
nand U469 (N_469,In_1056,In_814);
or U470 (N_470,In_1216,In_2189);
or U471 (N_471,In_1523,In_460);
or U472 (N_472,In_961,In_2280);
nor U473 (N_473,In_96,In_1765);
or U474 (N_474,In_954,In_532);
nand U475 (N_475,In_1815,In_1260);
or U476 (N_476,In_1538,In_1176);
or U477 (N_477,In_834,In_1740);
and U478 (N_478,In_2018,In_1803);
nand U479 (N_479,In_1763,In_1742);
and U480 (N_480,In_104,In_2335);
and U481 (N_481,In_874,In_2009);
or U482 (N_482,In_415,In_1293);
nand U483 (N_483,In_928,In_750);
nand U484 (N_484,In_1579,In_249);
nor U485 (N_485,In_1960,In_1186);
nand U486 (N_486,In_1205,In_869);
nor U487 (N_487,In_2246,In_1709);
xor U488 (N_488,In_1886,In_2117);
nand U489 (N_489,In_1983,In_2436);
or U490 (N_490,In_78,In_363);
or U491 (N_491,In_1758,In_771);
nand U492 (N_492,In_1785,In_2011);
or U493 (N_493,In_260,In_1263);
or U494 (N_494,In_628,In_0);
or U495 (N_495,In_1719,In_1412);
or U496 (N_496,In_938,In_429);
or U497 (N_497,In_111,In_861);
nor U498 (N_498,In_20,In_1939);
nand U499 (N_499,In_1580,In_2402);
nor U500 (N_500,In_741,In_520);
and U501 (N_501,In_1811,In_811);
or U502 (N_502,In_2150,In_394);
or U503 (N_503,In_1019,In_2492);
nor U504 (N_504,In_381,In_1813);
nor U505 (N_505,In_1273,In_1319);
nor U506 (N_506,In_1098,In_1143);
nor U507 (N_507,In_898,In_2418);
nor U508 (N_508,In_376,In_515);
nor U509 (N_509,In_1800,In_686);
nand U510 (N_510,In_231,In_1738);
nor U511 (N_511,In_311,In_358);
nor U512 (N_512,In_200,In_294);
nor U513 (N_513,In_1540,In_2133);
nand U514 (N_514,In_2483,In_2413);
and U515 (N_515,In_1937,In_2180);
or U516 (N_516,In_1410,In_1122);
and U517 (N_517,In_441,In_897);
nor U518 (N_518,In_1278,In_76);
or U519 (N_519,In_731,In_2398);
and U520 (N_520,In_1447,In_1111);
and U521 (N_521,In_2317,In_2373);
or U522 (N_522,In_315,In_1964);
and U523 (N_523,In_1559,In_970);
or U524 (N_524,In_604,In_1588);
or U525 (N_525,In_153,In_2109);
nand U526 (N_526,In_2095,In_2372);
nand U527 (N_527,In_822,In_979);
or U528 (N_528,In_522,In_2012);
nand U529 (N_529,In_47,In_2120);
nand U530 (N_530,In_1086,In_1451);
or U531 (N_531,In_1799,In_955);
nor U532 (N_532,In_896,In_2270);
nand U533 (N_533,In_205,In_118);
nand U534 (N_534,In_1126,In_2136);
or U535 (N_535,In_2407,In_2434);
nor U536 (N_536,In_1152,In_2370);
or U537 (N_537,In_125,In_2121);
or U538 (N_538,In_1108,In_2054);
and U539 (N_539,In_424,In_326);
and U540 (N_540,In_1422,In_744);
and U541 (N_541,In_866,In_1325);
nor U542 (N_542,In_306,In_2116);
or U543 (N_543,In_1869,In_405);
and U544 (N_544,In_1149,In_97);
nand U545 (N_545,In_2015,In_1542);
and U546 (N_546,In_1414,In_1444);
and U547 (N_547,In_1182,In_267);
nor U548 (N_548,In_509,In_2277);
nor U549 (N_549,In_1266,In_849);
and U550 (N_550,In_2361,In_711);
or U551 (N_551,In_1606,In_340);
nor U552 (N_552,In_120,In_1265);
nor U553 (N_553,In_1571,In_191);
nor U554 (N_554,In_1093,In_699);
nor U555 (N_555,In_39,In_1762);
nand U556 (N_556,In_1567,In_1989);
nand U557 (N_557,In_261,In_1500);
and U558 (N_558,In_1080,In_1468);
nand U559 (N_559,In_702,In_486);
nand U560 (N_560,In_737,In_66);
and U561 (N_561,In_367,In_375);
or U562 (N_562,In_489,In_157);
or U563 (N_563,In_2208,In_1489);
nand U564 (N_564,In_749,In_356);
and U565 (N_565,In_2131,In_2156);
and U566 (N_566,In_2215,In_1380);
nor U567 (N_567,In_1199,In_1165);
nor U568 (N_568,In_2130,In_139);
nor U569 (N_569,In_1164,In_149);
nand U570 (N_570,In_1327,In_1635);
and U571 (N_571,In_719,In_2267);
or U572 (N_572,In_568,In_1338);
or U573 (N_573,In_1991,In_1005);
or U574 (N_574,In_493,In_559);
and U575 (N_575,In_2032,In_2327);
or U576 (N_576,In_1462,In_1554);
nand U577 (N_577,In_560,In_1288);
and U578 (N_578,In_1858,In_596);
xor U579 (N_579,In_1012,In_2217);
nor U580 (N_580,In_1101,In_1090);
nor U581 (N_581,In_2160,In_270);
and U582 (N_582,In_1589,In_681);
and U583 (N_583,In_919,In_1943);
nand U584 (N_584,In_648,In_250);
nor U585 (N_585,In_51,In_1166);
or U586 (N_586,In_468,In_870);
nor U587 (N_587,In_480,In_1491);
nor U588 (N_588,In_88,In_1362);
or U589 (N_589,In_421,In_807);
or U590 (N_590,In_1416,In_726);
and U591 (N_591,In_1368,In_469);
and U592 (N_592,In_1916,In_1473);
nand U593 (N_593,In_312,In_1160);
nor U594 (N_594,In_2144,In_436);
nor U595 (N_595,In_2035,In_84);
nand U596 (N_596,In_857,In_645);
nor U597 (N_597,In_921,In_2385);
or U598 (N_598,In_1674,In_1524);
and U599 (N_599,In_1387,In_1994);
nand U600 (N_600,In_1221,In_1455);
nor U601 (N_601,In_2290,In_1499);
and U602 (N_602,In_652,In_629);
nor U603 (N_603,In_1705,In_1313);
or U604 (N_604,In_2355,In_2177);
and U605 (N_605,In_2110,In_2238);
or U606 (N_606,In_996,In_1240);
nor U607 (N_607,In_127,In_1594);
or U608 (N_608,In_1207,In_1275);
or U609 (N_609,In_1543,In_2386);
or U610 (N_610,In_2229,In_1637);
or U611 (N_611,In_1250,In_330);
nand U612 (N_612,In_508,In_2138);
and U613 (N_613,In_2345,In_1054);
or U614 (N_614,In_2445,In_1736);
or U615 (N_615,In_2383,In_959);
nand U616 (N_616,In_304,In_946);
or U617 (N_617,In_1179,In_1999);
nor U618 (N_618,In_2069,In_891);
nand U619 (N_619,In_2084,In_1643);
and U620 (N_620,In_158,In_2062);
and U621 (N_621,In_2346,In_302);
nor U622 (N_622,In_402,In_1533);
nand U623 (N_623,In_1909,In_1167);
and U624 (N_624,In_1479,In_1796);
and U625 (N_625,In_446,In_2298);
nand U626 (N_626,In_1645,In_1409);
nand U627 (N_627,In_1243,In_655);
or U628 (N_628,In_2187,In_359);
nor U629 (N_629,In_1545,In_1441);
and U630 (N_630,In_2446,In_1329);
nand U631 (N_631,In_753,In_431);
nand U632 (N_632,In_813,In_2357);
or U633 (N_633,In_2197,In_2188);
and U634 (N_634,In_1198,In_1723);
and U635 (N_635,In_2282,In_570);
nor U636 (N_636,In_1035,In_724);
and U637 (N_637,In_2333,In_1267);
and U638 (N_638,In_457,In_331);
nand U639 (N_639,In_1655,In_606);
or U640 (N_640,In_179,In_1038);
nand U641 (N_641,In_1465,In_1752);
nand U642 (N_642,In_904,In_1442);
or U643 (N_643,In_660,In_1530);
or U644 (N_644,In_2470,In_1953);
nor U645 (N_645,In_2423,In_2213);
nor U646 (N_646,In_1671,In_512);
nand U647 (N_647,In_437,In_1001);
or U648 (N_648,In_355,In_145);
or U649 (N_649,In_453,In_2328);
nand U650 (N_650,In_141,In_401);
or U651 (N_651,In_207,In_673);
and U652 (N_652,In_1931,In_2344);
or U653 (N_653,In_7,In_541);
nand U654 (N_654,In_2468,In_1515);
nand U655 (N_655,In_1744,In_762);
nor U656 (N_656,In_121,In_41);
nor U657 (N_657,In_2352,In_2017);
and U658 (N_658,In_1855,In_2145);
and U659 (N_659,In_1798,In_69);
nand U660 (N_660,In_782,In_852);
nand U661 (N_661,In_379,In_1599);
or U662 (N_662,In_1452,In_2091);
xor U663 (N_663,In_1255,In_844);
nor U664 (N_664,In_2212,In_2422);
nor U665 (N_665,In_1134,In_936);
and U666 (N_666,In_277,In_225);
and U667 (N_667,In_2443,In_1471);
nand U668 (N_668,In_1271,In_935);
and U669 (N_669,In_369,In_1217);
nor U670 (N_670,In_1717,In_505);
nand U671 (N_671,In_1073,In_1247);
nand U672 (N_672,In_916,In_291);
nand U673 (N_673,In_535,In_1842);
nand U674 (N_674,In_670,In_592);
nand U675 (N_675,In_1094,In_1239);
nand U676 (N_676,In_1168,In_2421);
and U677 (N_677,In_2293,In_706);
or U678 (N_678,In_1911,In_1607);
and U679 (N_679,In_1687,In_1761);
and U680 (N_680,In_284,In_406);
nor U681 (N_681,In_1061,In_1859);
nand U682 (N_682,In_879,In_2239);
nor U683 (N_683,In_2000,In_620);
and U684 (N_684,In_1695,In_1456);
nor U685 (N_685,In_1064,In_888);
or U686 (N_686,In_2127,In_2147);
or U687 (N_687,In_1233,In_1930);
or U688 (N_688,In_1732,In_2359);
and U689 (N_689,In_1836,In_61);
nor U690 (N_690,In_602,In_746);
or U691 (N_691,In_2193,In_2211);
nor U692 (N_692,In_1003,In_160);
nor U693 (N_693,In_1899,In_565);
or U694 (N_694,In_684,In_1794);
or U695 (N_695,In_1258,In_2092);
nand U696 (N_696,In_832,In_1547);
nor U697 (N_697,In_2007,In_657);
nor U698 (N_698,In_2489,In_2214);
or U699 (N_699,In_1120,In_238);
and U700 (N_700,In_766,In_669);
and U701 (N_701,In_117,In_2253);
and U702 (N_702,In_2003,In_1314);
and U703 (N_703,In_226,In_1284);
nor U704 (N_704,In_479,In_2090);
and U705 (N_705,In_1974,In_1204);
nand U706 (N_706,In_1749,In_1018);
or U707 (N_707,In_1440,In_1987);
or U708 (N_708,In_2409,In_685);
or U709 (N_709,In_1251,In_1629);
and U710 (N_710,In_1976,In_1315);
nor U711 (N_711,In_1077,In_1156);
nand U712 (N_712,In_411,In_334);
nand U713 (N_713,In_1046,In_566);
nand U714 (N_714,In_3,In_2063);
and U715 (N_715,In_2218,In_1353);
or U716 (N_716,In_588,In_112);
or U717 (N_717,In_1532,In_908);
nand U718 (N_718,In_1195,In_2281);
or U719 (N_719,In_1614,In_2366);
nand U720 (N_720,In_1564,In_537);
and U721 (N_721,In_2401,In_2415);
nand U722 (N_722,In_2476,In_1188);
and U723 (N_723,In_499,In_2340);
nor U724 (N_724,In_2363,In_1323);
nand U725 (N_725,In_1023,In_1774);
and U726 (N_726,In_692,In_1045);
nor U727 (N_727,In_2307,In_2074);
or U728 (N_728,In_1517,In_2139);
nor U729 (N_729,In_1925,In_2301);
nand U730 (N_730,In_1797,In_1984);
nand U731 (N_731,In_677,In_318);
nand U732 (N_732,In_821,In_1757);
nand U733 (N_733,In_2330,In_1910);
and U734 (N_734,In_368,In_439);
nor U735 (N_735,In_2475,In_2221);
nor U736 (N_736,In_1682,In_1816);
nand U737 (N_737,In_2006,In_892);
or U738 (N_738,In_1550,In_1303);
nand U739 (N_739,In_1527,In_772);
and U740 (N_740,In_536,In_1316);
nand U741 (N_741,In_538,In_107);
nand U742 (N_742,In_1809,In_1141);
nand U743 (N_743,In_216,In_601);
and U744 (N_744,In_2309,In_48);
or U745 (N_745,In_195,In_994);
and U746 (N_746,In_1788,In_614);
nand U747 (N_747,In_899,In_1450);
or U748 (N_748,In_1376,In_526);
nor U749 (N_749,In_1849,In_1525);
and U750 (N_750,In_1050,In_1175);
nand U751 (N_751,In_2047,In_2186);
nor U752 (N_752,In_1331,In_2043);
and U753 (N_753,In_796,In_1384);
and U754 (N_754,In_1505,In_2493);
or U755 (N_755,In_800,In_1301);
or U756 (N_756,In_80,In_2244);
and U757 (N_757,In_1566,In_455);
nand U758 (N_758,In_251,In_287);
nand U759 (N_759,In_2397,In_222);
or U760 (N_760,In_2380,In_2490);
nor U761 (N_761,In_178,In_945);
nand U762 (N_762,In_1091,In_2076);
and U763 (N_763,In_890,In_1628);
xnor U764 (N_764,In_770,In_438);
and U765 (N_765,In_1720,In_1463);
or U766 (N_766,In_67,In_2403);
nand U767 (N_767,In_836,In_608);
nor U768 (N_768,In_735,In_1624);
and U769 (N_769,In_199,In_1583);
nor U770 (N_770,In_963,In_2073);
nor U771 (N_771,In_1049,In_1784);
and U772 (N_772,In_1529,In_2159);
nand U773 (N_773,In_34,In_577);
and U774 (N_774,In_803,In_1857);
nand U775 (N_775,In_597,In_572);
nor U776 (N_776,In_1694,In_1575);
or U777 (N_777,In_1144,In_720);
nand U778 (N_778,In_871,In_2300);
nor U779 (N_779,In_452,In_1429);
nand U780 (N_780,In_1581,In_1170);
or U781 (N_781,In_1954,In_275);
or U782 (N_782,In_2419,In_2081);
and U783 (N_783,In_1208,In_400);
and U784 (N_784,In_2440,In_1546);
and U785 (N_785,In_1497,In_664);
nor U786 (N_786,In_1289,In_2496);
or U787 (N_787,In_1826,In_2030);
and U788 (N_788,In_1010,In_876);
and U789 (N_789,In_556,In_298);
nand U790 (N_790,In_248,In_1634);
nor U791 (N_791,In_307,In_1474);
or U792 (N_792,In_788,In_989);
nor U793 (N_793,In_2394,In_626);
nand U794 (N_794,In_1328,In_703);
nand U795 (N_795,In_134,In_1900);
nor U796 (N_796,In_2044,In_528);
or U797 (N_797,In_830,In_1069);
and U798 (N_798,In_858,In_258);
or U799 (N_799,In_843,In_2075);
or U800 (N_800,In_1034,In_378);
nor U801 (N_801,In_2,In_1676);
and U802 (N_802,In_828,In_2457);
or U803 (N_803,In_283,In_463);
and U804 (N_804,In_1878,In_2124);
and U805 (N_805,In_1016,In_2064);
nor U806 (N_806,In_804,In_1608);
and U807 (N_807,In_1779,In_217);
nor U808 (N_808,In_1074,In_188);
nand U809 (N_809,In_420,In_1848);
nand U810 (N_810,In_1079,In_1201);
or U811 (N_811,In_1311,In_1369);
nand U812 (N_812,In_1324,In_2171);
nand U813 (N_813,In_295,In_1935);
nor U814 (N_814,In_1087,In_1582);
and U815 (N_815,In_2176,In_1959);
and U816 (N_816,In_1952,In_219);
and U817 (N_817,In_1971,In_718);
and U818 (N_818,In_1613,In_2048);
and U819 (N_819,In_17,In_1844);
or U820 (N_820,In_1689,In_1004);
nand U821 (N_821,In_92,In_245);
nor U822 (N_822,In_445,In_2428);
nand U823 (N_823,In_2448,In_2167);
nand U824 (N_824,In_2216,In_1286);
xnor U825 (N_825,In_35,In_1704);
and U826 (N_826,In_1125,In_2250);
and U827 (N_827,In_1632,In_296);
nor U828 (N_828,In_2360,In_1361);
nor U829 (N_829,In_2311,In_2487);
or U830 (N_830,In_1693,In_1485);
xnor U831 (N_831,In_1609,In_1879);
nor U832 (N_832,In_2485,In_715);
nor U833 (N_833,In_915,In_485);
and U834 (N_834,In_33,In_591);
nand U835 (N_835,In_2181,In_925);
nor U836 (N_836,In_2455,In_732);
nand U837 (N_837,In_243,In_775);
nand U838 (N_838,In_1492,In_2467);
nand U839 (N_839,In_1345,In_831);
or U840 (N_840,In_1433,In_646);
nand U841 (N_841,In_1895,In_1884);
nor U842 (N_842,In_1197,In_386);
nand U843 (N_843,In_1398,In_290);
nor U844 (N_844,In_1649,In_2060);
xnor U845 (N_845,In_2416,In_2111);
nor U846 (N_846,In_215,In_542);
or U847 (N_847,In_1923,In_1557);
nand U848 (N_848,In_2240,In_1845);
and U849 (N_849,In_1726,In_1401);
and U850 (N_850,In_2305,In_818);
nand U851 (N_851,In_1389,In_863);
or U852 (N_852,In_1506,In_571);
and U853 (N_853,In_819,In_322);
nor U854 (N_854,In_999,In_1135);
or U855 (N_855,In_2070,In_619);
and U856 (N_856,In_651,In_1026);
or U857 (N_857,In_2262,In_1052);
nand U858 (N_858,In_927,In_2353);
or U859 (N_859,In_2294,In_214);
or U860 (N_860,In_510,In_739);
and U861 (N_861,In_2016,In_1318);
nand U862 (N_862,In_2236,In_30);
and U863 (N_863,In_495,In_1);
and U864 (N_864,In_848,In_1390);
nand U865 (N_865,In_949,In_1317);
or U866 (N_866,In_2381,In_644);
or U867 (N_867,In_1544,In_1764);
nor U868 (N_868,In_2220,In_902);
nor U869 (N_869,In_2378,In_1322);
nor U870 (N_870,In_83,In_1572);
nor U871 (N_871,In_2005,In_1936);
xnor U872 (N_872,In_656,In_798);
and U873 (N_873,In_1600,In_1620);
or U874 (N_874,In_983,In_2405);
nor U875 (N_875,In_1161,In_1146);
nor U876 (N_876,In_1541,In_2365);
nand U877 (N_877,In_1159,In_2224);
and U878 (N_878,In_1563,In_2077);
nand U879 (N_879,In_969,In_1420);
nor U880 (N_880,In_2237,In_166);
or U881 (N_881,In_278,In_2049);
nor U882 (N_882,In_1223,In_142);
and U883 (N_883,In_690,In_1562);
nor U884 (N_884,In_545,In_2420);
nand U885 (N_885,In_2367,In_1425);
or U886 (N_886,In_647,In_981);
and U887 (N_887,In_708,In_760);
and U888 (N_888,In_1573,In_1770);
nor U889 (N_889,In_2255,In_373);
and U890 (N_890,In_643,In_1707);
or U891 (N_891,In_529,In_1102);
nand U892 (N_892,In_82,In_314);
nand U893 (N_893,In_567,In_1037);
or U894 (N_894,In_2161,In_977);
and U895 (N_895,In_1560,In_2341);
nand U896 (N_896,In_1254,In_824);
nand U897 (N_897,In_366,In_143);
xor U898 (N_898,In_1891,In_845);
xor U899 (N_899,In_1751,In_2185);
or U900 (N_900,In_1975,In_1203);
nor U901 (N_901,In_413,In_1548);
xnor U902 (N_902,In_464,In_1238);
or U903 (N_903,In_1139,In_1834);
nand U904 (N_904,In_631,In_2292);
or U905 (N_905,In_1326,In_343);
nand U906 (N_906,In_473,In_1681);
and U907 (N_907,In_860,In_884);
or U908 (N_908,In_1521,In_1697);
nor U909 (N_909,In_2310,In_909);
and U910 (N_910,In_496,In_2071);
nor U911 (N_911,In_45,In_2400);
nor U912 (N_912,In_2021,In_1213);
nand U913 (N_913,In_1379,In_1030);
or U914 (N_914,In_972,In_1833);
nand U915 (N_915,In_24,In_1358);
and U916 (N_916,In_1063,In_409);
or U917 (N_917,In_1549,In_324);
nand U918 (N_918,In_563,In_2219);
nor U919 (N_919,In_2041,In_2254);
nor U920 (N_920,In_1656,In_224);
nor U921 (N_921,In_2210,In_1065);
and U922 (N_922,In_603,In_1633);
or U923 (N_923,In_2442,In_1394);
nor U924 (N_924,In_1860,In_467);
or U925 (N_925,In_950,In_903);
and U926 (N_926,In_881,In_140);
nor U927 (N_927,In_12,In_1430);
or U928 (N_928,In_2273,In_1443);
and U929 (N_929,In_1980,In_713);
or U930 (N_930,In_1932,In_1806);
nand U931 (N_931,In_582,In_1660);
or U932 (N_932,In_449,In_1597);
and U933 (N_933,In_113,In_1292);
and U934 (N_934,In_562,In_223);
nor U935 (N_935,In_1008,In_527);
and U936 (N_936,In_1743,In_418);
and U937 (N_937,In_1354,In_1982);
nor U938 (N_938,In_1106,In_1679);
nor U939 (N_939,In_1230,In_1961);
or U940 (N_940,In_997,In_2460);
or U941 (N_941,In_1734,In_2040);
or U942 (N_942,In_621,In_1890);
nand U943 (N_943,In_346,In_1212);
or U944 (N_944,In_2164,In_2105);
or U945 (N_945,In_2425,In_194);
or U946 (N_946,In_466,In_992);
nor U947 (N_947,In_930,In_1593);
or U948 (N_948,In_2020,In_2055);
or U949 (N_949,In_342,In_801);
and U950 (N_950,In_71,In_984);
nor U951 (N_951,In_85,In_1917);
and U952 (N_952,In_1686,In_1269);
nor U953 (N_953,In_966,In_1670);
and U954 (N_954,In_1025,In_847);
nand U955 (N_955,In_2190,In_461);
nand U956 (N_956,In_1151,In_2272);
and U957 (N_957,In_169,In_1333);
nand U958 (N_958,In_2002,In_230);
or U959 (N_959,In_2306,In_1383);
nand U960 (N_960,In_2205,In_1706);
or U961 (N_961,In_633,In_2039);
nand U962 (N_962,In_1096,In_2329);
and U963 (N_963,In_2326,In_328);
or U964 (N_964,In_1299,In_1206);
and U965 (N_965,In_531,In_2304);
or U966 (N_966,In_482,In_2332);
and U967 (N_967,In_1590,In_390);
or U968 (N_968,In_666,In_1950);
nand U969 (N_969,In_755,In_299);
nor U970 (N_970,In_547,In_767);
or U971 (N_971,In_14,In_152);
and U972 (N_972,In_1838,In_917);
and U973 (N_973,In_1406,In_1400);
nor U974 (N_974,In_1810,In_1827);
or U975 (N_975,In_864,In_1417);
or U976 (N_976,In_2316,In_2269);
or U977 (N_977,In_679,In_519);
or U978 (N_978,In_2275,In_2247);
xnor U979 (N_979,In_185,In_204);
nand U980 (N_980,In_1075,In_484);
nor U981 (N_981,In_513,In_576);
nor U982 (N_982,In_1995,In_2429);
and U983 (N_983,In_1476,In_616);
nor U984 (N_984,In_184,In_1846);
nor U985 (N_985,In_662,In_1234);
nand U986 (N_986,In_517,In_2174);
nand U987 (N_987,In_2384,In_135);
nor U988 (N_988,In_116,In_1033);
nor U989 (N_989,In_1365,In_548);
nor U990 (N_990,In_435,In_1874);
nor U991 (N_991,In_95,In_2113);
or U992 (N_992,In_380,In_271);
and U993 (N_993,In_488,In_958);
nand U994 (N_994,In_2052,In_743);
nand U995 (N_995,In_1113,In_1730);
nand U996 (N_996,In_680,In_1068);
and U997 (N_997,In_1235,In_2165);
nor U998 (N_998,In_1993,In_1381);
nor U999 (N_999,In_779,In_947);
nand U1000 (N_1000,In_1162,In_2322);
or U1001 (N_1001,In_634,In_434);
and U1002 (N_1002,In_419,In_414);
nor U1003 (N_1003,In_1227,In_2079);
or U1004 (N_1004,In_1507,In_2022);
nand U1005 (N_1005,In_978,In_751);
nor U1006 (N_1006,In_2321,In_1428);
nand U1007 (N_1007,In_2498,In_1215);
nor U1008 (N_1008,In_129,In_433);
or U1009 (N_1009,In_2417,In_2209);
or U1010 (N_1010,In_301,In_1814);
nor U1011 (N_1011,In_362,In_2226);
nor U1012 (N_1012,In_1109,In_1745);
and U1013 (N_1013,In_1922,In_2392);
and U1014 (N_1014,In_761,In_1990);
and U1015 (N_1015,In_553,In_1209);
or U1016 (N_1016,In_2051,In_209);
and U1017 (N_1017,In_1942,In_289);
nor U1018 (N_1018,In_839,In_1228);
nor U1019 (N_1019,In_2252,In_583);
or U1020 (N_1020,In_465,In_707);
nand U1021 (N_1021,In_2302,In_1822);
xor U1022 (N_1022,In_2427,In_1883);
nand U1023 (N_1023,In_1568,In_1535);
nor U1024 (N_1024,In_1824,In_2243);
nor U1025 (N_1025,In_1366,In_721);
nand U1026 (N_1026,In_2390,In_674);
nor U1027 (N_1027,In_2175,In_2249);
or U1028 (N_1028,In_600,In_641);
or U1029 (N_1029,In_2028,In_159);
nand U1030 (N_1030,In_1963,In_305);
nand U1031 (N_1031,In_1405,In_1483);
nor U1032 (N_1032,In_1918,In_875);
or U1033 (N_1033,In_221,In_2098);
or U1034 (N_1034,In_1224,In_841);
nand U1035 (N_1035,In_1578,In_1426);
nand U1036 (N_1036,In_2263,In_2149);
and U1037 (N_1037,In_1690,In_89);
and U1038 (N_1038,In_265,In_2045);
and U1039 (N_1039,In_1551,In_456);
and U1040 (N_1040,In_1586,In_313);
or U1041 (N_1041,In_754,In_2199);
nor U1042 (N_1042,In_227,In_590);
nor U1043 (N_1043,In_2410,In_593);
and U1044 (N_1044,In_1948,In_8);
or U1045 (N_1045,In_1339,In_1808);
and U1046 (N_1046,In_115,In_398);
and U1047 (N_1047,In_1561,In_2471);
nor U1048 (N_1048,In_1508,In_2038);
nand U1049 (N_1049,In_2337,In_727);
nor U1050 (N_1050,In_329,In_1513);
nor U1051 (N_1051,In_1413,In_1006);
nor U1052 (N_1052,In_472,In_900);
xor U1053 (N_1053,In_2299,In_70);
and U1054 (N_1054,In_1696,In_213);
or U1055 (N_1055,In_2046,In_1127);
nand U1056 (N_1056,In_2289,In_1793);
nor U1057 (N_1057,In_202,In_1539);
nand U1058 (N_1058,In_422,In_384);
and U1059 (N_1059,In_610,In_1092);
and U1060 (N_1060,In_1904,In_1382);
and U1061 (N_1061,In_1512,In_1100);
and U1062 (N_1062,In_914,In_387);
or U1063 (N_1063,In_793,In_1084);
and U1064 (N_1064,In_498,In_1099);
and U1065 (N_1065,In_1027,In_101);
nand U1066 (N_1066,In_471,In_758);
nand U1067 (N_1067,In_15,In_862);
nor U1068 (N_1068,In_1427,In_1040);
or U1069 (N_1069,In_540,In_242);
and U1070 (N_1070,In_1737,In_177);
and U1071 (N_1071,In_477,In_1024);
and U1072 (N_1072,In_1592,In_56);
nand U1073 (N_1073,In_2118,In_1355);
nand U1074 (N_1074,In_353,In_494);
nand U1075 (N_1075,In_960,In_2364);
and U1076 (N_1076,In_2202,In_1154);
or U1077 (N_1077,In_333,In_1487);
nand U1078 (N_1078,In_521,In_241);
nor U1079 (N_1079,In_198,In_1140);
and U1080 (N_1080,In_1776,In_1708);
and U1081 (N_1081,In_1344,In_2196);
and U1082 (N_1082,In_186,In_1537);
or U1083 (N_1083,In_1357,In_428);
nand U1084 (N_1084,In_2426,In_345);
nor U1085 (N_1085,In_371,In_1667);
and U1086 (N_1086,In_2480,In_2408);
and U1087 (N_1087,In_1478,In_1841);
and U1088 (N_1088,In_986,In_1297);
nand U1089 (N_1089,In_1036,In_310);
or U1090 (N_1090,In_1000,In_1640);
nor U1091 (N_1091,In_90,In_1534);
and U1092 (N_1092,In_497,In_138);
nand U1093 (N_1093,In_1789,In_1374);
nand U1094 (N_1094,In_1825,In_64);
or U1095 (N_1095,In_1128,In_2204);
or U1096 (N_1096,In_370,In_975);
or U1097 (N_1097,In_1193,In_1638);
nor U1098 (N_1098,In_812,In_175);
nor U1099 (N_1099,In_642,In_1103);
and U1100 (N_1100,In_624,In_611);
and U1101 (N_1101,In_1060,In_1919);
and U1102 (N_1102,In_2452,In_773);
or U1103 (N_1103,In_905,In_2023);
or U1104 (N_1104,In_123,In_1348);
nand U1105 (N_1105,In_1829,In_668);
and U1106 (N_1106,In_1184,In_1155);
or U1107 (N_1107,In_182,In_344);
or U1108 (N_1108,In_1078,In_2441);
nor U1109 (N_1109,In_2497,In_2106);
and U1110 (N_1110,In_2128,In_2414);
or U1111 (N_1111,In_408,In_2163);
or U1112 (N_1112,In_1114,In_1767);
or U1113 (N_1113,In_36,In_2438);
or U1114 (N_1114,In_1190,In_704);
and U1115 (N_1115,In_2086,In_374);
nor U1116 (N_1116,In_1576,In_2342);
xnor U1117 (N_1117,In_432,In_1469);
or U1118 (N_1118,In_1385,In_365);
and U1119 (N_1119,In_2194,In_232);
nand U1120 (N_1120,In_288,In_1194);
and U1121 (N_1121,In_709,In_1639);
nor U1122 (N_1122,In_280,In_1941);
nand U1123 (N_1123,In_2104,In_1147);
and U1124 (N_1124,In_2461,In_234);
or U1125 (N_1125,In_1510,In_1711);
nand U1126 (N_1126,In_1611,In_2488);
nor U1127 (N_1127,In_1920,In_1747);
or U1128 (N_1128,In_124,In_208);
nor U1129 (N_1129,In_425,In_1536);
nand U1130 (N_1130,In_2245,In_136);
nor U1131 (N_1131,In_1088,In_1804);
and U1132 (N_1132,In_2134,In_1733);
or U1133 (N_1133,In_2027,In_462);
nor U1134 (N_1134,In_2336,In_1728);
nor U1135 (N_1135,In_172,In_2078);
or U1136 (N_1136,In_714,In_733);
nand U1137 (N_1137,In_1866,In_1277);
or U1138 (N_1138,In_1669,In_262);
nor U1139 (N_1139,In_1285,In_933);
nand U1140 (N_1140,In_1397,In_1741);
or U1141 (N_1141,In_404,In_2459);
and U1142 (N_1142,In_1408,In_1484);
nor U1143 (N_1143,In_2296,In_575);
nor U1144 (N_1144,In_1837,In_93);
nor U1145 (N_1145,In_1598,In_1956);
or U1146 (N_1146,In_1352,In_1619);
nor U1147 (N_1147,In_2288,In_478);
and U1148 (N_1148,In_518,In_2157);
nor U1149 (N_1149,In_1969,In_826);
nor U1150 (N_1150,In_2279,In_554);
nor U1151 (N_1151,In_987,In_2494);
and U1152 (N_1152,In_1264,In_894);
and U1153 (N_1153,In_1831,In_1229);
and U1154 (N_1154,In_131,In_1290);
nand U1155 (N_1155,In_653,In_1888);
or U1156 (N_1156,In_1309,In_1944);
nand U1157 (N_1157,In_1658,In_693);
and U1158 (N_1158,In_1650,In_1022);
and U1159 (N_1159,In_87,In_2223);
and U1160 (N_1160,In_799,In_630);
xnor U1161 (N_1161,In_372,In_189);
or U1162 (N_1162,In_2085,In_2201);
or U1163 (N_1163,In_878,In_2450);
nand U1164 (N_1164,In_1893,In_777);
nand U1165 (N_1165,In_618,In_877);
and U1166 (N_1166,In_752,In_174);
and U1167 (N_1167,In_1055,In_2242);
nand U1168 (N_1168,In_2094,In_1312);
and U1169 (N_1169,In_2019,In_130);
or U1170 (N_1170,In_1391,In_1457);
nand U1171 (N_1171,In_388,In_176);
nor U1172 (N_1172,In_86,In_1898);
or U1173 (N_1173,In_1622,In_1921);
nor U1174 (N_1174,In_931,In_1453);
nand U1175 (N_1175,In_1754,In_1496);
nor U1176 (N_1176,In_2057,In_1905);
or U1177 (N_1177,In_501,In_28);
and U1178 (N_1178,In_1680,In_632);
or U1179 (N_1179,In_710,In_1683);
or U1180 (N_1180,In_1873,In_912);
and U1181 (N_1181,In_192,In_1245);
nand U1182 (N_1182,In_2231,In_1585);
nor U1183 (N_1183,In_792,In_4);
and U1184 (N_1184,In_1955,In_2198);
or U1185 (N_1185,In_1584,In_1894);
and U1186 (N_1186,In_1307,In_327);
or U1187 (N_1187,In_323,In_1912);
and U1188 (N_1188,In_1467,In_1256);
and U1189 (N_1189,In_98,In_1684);
and U1190 (N_1190,In_1341,In_671);
nand U1191 (N_1191,In_1360,In_1276);
nand U1192 (N_1192,In_1014,In_747);
and U1193 (N_1193,In_1153,In_1028);
or U1194 (N_1194,In_911,In_1832);
and U1195 (N_1195,In_940,In_109);
or U1196 (N_1196,In_1795,In_1435);
nor U1197 (N_1197,In_1865,In_2268);
nand U1198 (N_1198,In_168,In_233);
nand U1199 (N_1199,In_2377,In_2276);
nand U1200 (N_1200,In_2283,In_1772);
nor U1201 (N_1201,In_1180,In_1495);
or U1202 (N_1202,In_1241,In_2235);
nand U1203 (N_1203,In_2001,In_2491);
and U1204 (N_1204,In_1914,In_783);
nor U1205 (N_1205,In_2411,In_672);
nor U1206 (N_1206,In_239,In_1504);
or U1207 (N_1207,In_2179,In_2315);
nor U1208 (N_1208,In_1039,In_2126);
or U1209 (N_1209,In_1115,In_6);
nor U1210 (N_1210,In_350,In_114);
and U1211 (N_1211,In_1270,In_939);
nand U1212 (N_1212,In_2439,In_2135);
and U1213 (N_1213,In_351,In_2088);
and U1214 (N_1214,In_247,In_272);
and U1215 (N_1215,In_2354,In_805);
nor U1216 (N_1216,In_605,In_924);
nand U1217 (N_1217,In_524,In_635);
or U1218 (N_1218,In_1769,In_2469);
and U1219 (N_1219,In_1631,In_988);
nor U1220 (N_1220,In_942,In_951);
xnor U1221 (N_1221,In_49,In_2458);
and U1222 (N_1222,In_794,In_1481);
nand U1223 (N_1223,In_133,In_155);
and U1224 (N_1224,In_1509,In_1493);
nand U1225 (N_1225,In_1603,In_1518);
nor U1226 (N_1226,In_2162,In_2265);
and U1227 (N_1227,In_923,In_998);
and U1228 (N_1228,In_1142,In_1965);
and U1229 (N_1229,In_154,In_791);
and U1230 (N_1230,In_2338,In_197);
nand U1231 (N_1231,In_650,In_382);
or U1232 (N_1232,In_268,In_1132);
nor U1233 (N_1233,In_2331,In_2148);
and U1234 (N_1234,In_776,In_1335);
or U1235 (N_1235,In_2257,In_100);
or U1236 (N_1236,In_1337,In_1150);
or U1237 (N_1237,In_1248,In_282);
or U1238 (N_1238,In_698,In_2169);
or U1239 (N_1239,In_723,In_319);
nand U1240 (N_1240,In_2406,In_1392);
nand U1241 (N_1241,In_220,In_500);
and U1242 (N_1242,In_1700,In_65);
nand U1243 (N_1243,In_2320,In_1364);
nor U1244 (N_1244,In_68,In_661);
nor U1245 (N_1245,In_530,In_40);
xnor U1246 (N_1246,In_72,In_2234);
or U1247 (N_1247,In_2258,In_38);
nor U1248 (N_1248,In_1189,In_1305);
or U1249 (N_1249,In_1431,In_1232);
nand U1250 (N_1250,In_1525,In_2449);
nand U1251 (N_1251,In_811,In_2217);
or U1252 (N_1252,In_1371,In_705);
nand U1253 (N_1253,In_1129,In_602);
nand U1254 (N_1254,In_658,In_1529);
and U1255 (N_1255,In_84,In_1139);
nor U1256 (N_1256,In_324,In_2381);
nand U1257 (N_1257,In_2324,In_1094);
nand U1258 (N_1258,In_606,In_774);
nor U1259 (N_1259,In_900,In_2109);
nor U1260 (N_1260,In_932,In_2116);
nand U1261 (N_1261,In_1857,In_2121);
or U1262 (N_1262,In_142,In_795);
or U1263 (N_1263,In_2135,In_2469);
or U1264 (N_1264,In_743,In_172);
nor U1265 (N_1265,In_2390,In_2113);
or U1266 (N_1266,In_2250,In_1879);
or U1267 (N_1267,In_1775,In_1376);
and U1268 (N_1268,In_1855,In_1556);
nand U1269 (N_1269,In_1690,In_1549);
and U1270 (N_1270,In_761,In_592);
nand U1271 (N_1271,In_2064,In_13);
nand U1272 (N_1272,In_658,In_1497);
xnor U1273 (N_1273,In_767,In_167);
nor U1274 (N_1274,In_738,In_1741);
nor U1275 (N_1275,In_1367,In_1583);
or U1276 (N_1276,In_649,In_1807);
nand U1277 (N_1277,In_1112,In_797);
nand U1278 (N_1278,In_313,In_23);
nand U1279 (N_1279,In_1256,In_1520);
nor U1280 (N_1280,In_1926,In_217);
and U1281 (N_1281,In_1218,In_2405);
or U1282 (N_1282,In_808,In_1646);
nor U1283 (N_1283,In_788,In_1529);
nor U1284 (N_1284,In_844,In_485);
nor U1285 (N_1285,In_1394,In_1545);
nand U1286 (N_1286,In_1199,In_116);
nor U1287 (N_1287,In_482,In_655);
or U1288 (N_1288,In_2420,In_423);
nor U1289 (N_1289,In_905,In_1606);
nor U1290 (N_1290,In_595,In_1800);
nor U1291 (N_1291,In_600,In_2480);
or U1292 (N_1292,In_1999,In_2406);
nor U1293 (N_1293,In_363,In_1239);
and U1294 (N_1294,In_2456,In_1624);
nand U1295 (N_1295,In_1449,In_2217);
or U1296 (N_1296,In_504,In_7);
or U1297 (N_1297,In_2159,In_2061);
nor U1298 (N_1298,In_1865,In_143);
nand U1299 (N_1299,In_377,In_2418);
and U1300 (N_1300,In_2035,In_1425);
and U1301 (N_1301,In_2486,In_2131);
nor U1302 (N_1302,In_692,In_1652);
nor U1303 (N_1303,In_1948,In_1518);
or U1304 (N_1304,In_1764,In_268);
and U1305 (N_1305,In_1972,In_1951);
or U1306 (N_1306,In_1413,In_1769);
and U1307 (N_1307,In_25,In_780);
or U1308 (N_1308,In_988,In_301);
and U1309 (N_1309,In_2307,In_748);
or U1310 (N_1310,In_635,In_1261);
or U1311 (N_1311,In_2188,In_327);
nand U1312 (N_1312,In_180,In_2470);
xor U1313 (N_1313,In_1794,In_973);
or U1314 (N_1314,In_1949,In_1562);
or U1315 (N_1315,In_259,In_1332);
and U1316 (N_1316,In_1276,In_1286);
nand U1317 (N_1317,In_242,In_618);
and U1318 (N_1318,In_1156,In_1289);
xnor U1319 (N_1319,In_157,In_2491);
and U1320 (N_1320,In_2,In_167);
and U1321 (N_1321,In_370,In_1306);
or U1322 (N_1322,In_1878,In_791);
and U1323 (N_1323,In_1205,In_1429);
and U1324 (N_1324,In_1797,In_1155);
nor U1325 (N_1325,In_877,In_554);
nor U1326 (N_1326,In_1619,In_1683);
and U1327 (N_1327,In_520,In_2157);
or U1328 (N_1328,In_1954,In_1636);
nand U1329 (N_1329,In_1109,In_2174);
xnor U1330 (N_1330,In_1228,In_2285);
nand U1331 (N_1331,In_1679,In_1694);
nand U1332 (N_1332,In_2009,In_599);
nand U1333 (N_1333,In_158,In_1371);
and U1334 (N_1334,In_1463,In_625);
and U1335 (N_1335,In_2107,In_727);
and U1336 (N_1336,In_1190,In_687);
or U1337 (N_1337,In_2169,In_1554);
nor U1338 (N_1338,In_186,In_2112);
nand U1339 (N_1339,In_1045,In_1240);
or U1340 (N_1340,In_2339,In_2295);
nand U1341 (N_1341,In_4,In_1424);
nand U1342 (N_1342,In_2157,In_1045);
or U1343 (N_1343,In_812,In_1757);
nand U1344 (N_1344,In_1264,In_633);
nor U1345 (N_1345,In_1337,In_1863);
or U1346 (N_1346,In_631,In_468);
nand U1347 (N_1347,In_208,In_1449);
nand U1348 (N_1348,In_1081,In_136);
or U1349 (N_1349,In_201,In_985);
nor U1350 (N_1350,In_378,In_699);
nand U1351 (N_1351,In_707,In_331);
or U1352 (N_1352,In_1249,In_51);
nand U1353 (N_1353,In_1641,In_2064);
and U1354 (N_1354,In_894,In_2148);
nand U1355 (N_1355,In_2112,In_194);
xor U1356 (N_1356,In_2361,In_1337);
nand U1357 (N_1357,In_1847,In_43);
nand U1358 (N_1358,In_2451,In_447);
nand U1359 (N_1359,In_1608,In_2339);
nor U1360 (N_1360,In_936,In_1824);
nand U1361 (N_1361,In_157,In_1053);
nor U1362 (N_1362,In_497,In_313);
nand U1363 (N_1363,In_496,In_13);
nor U1364 (N_1364,In_2410,In_1883);
xnor U1365 (N_1365,In_1642,In_2387);
nand U1366 (N_1366,In_1001,In_1888);
and U1367 (N_1367,In_206,In_378);
and U1368 (N_1368,In_487,In_1593);
and U1369 (N_1369,In_2375,In_159);
xnor U1370 (N_1370,In_958,In_2068);
or U1371 (N_1371,In_1182,In_1448);
or U1372 (N_1372,In_1511,In_614);
and U1373 (N_1373,In_1435,In_1031);
nand U1374 (N_1374,In_1698,In_194);
or U1375 (N_1375,In_406,In_1691);
nand U1376 (N_1376,In_2006,In_20);
nor U1377 (N_1377,In_2228,In_2106);
nand U1378 (N_1378,In_1977,In_1532);
nand U1379 (N_1379,In_1219,In_2348);
nor U1380 (N_1380,In_2149,In_2232);
nand U1381 (N_1381,In_402,In_1735);
or U1382 (N_1382,In_1277,In_573);
nand U1383 (N_1383,In_2261,In_914);
nand U1384 (N_1384,In_2005,In_1968);
and U1385 (N_1385,In_1437,In_848);
nand U1386 (N_1386,In_913,In_1281);
nor U1387 (N_1387,In_974,In_211);
nand U1388 (N_1388,In_718,In_1610);
xnor U1389 (N_1389,In_2359,In_1749);
nand U1390 (N_1390,In_412,In_895);
nand U1391 (N_1391,In_1035,In_305);
nand U1392 (N_1392,In_2452,In_2172);
and U1393 (N_1393,In_1511,In_865);
nand U1394 (N_1394,In_2374,In_1326);
nor U1395 (N_1395,In_617,In_414);
nand U1396 (N_1396,In_1452,In_531);
and U1397 (N_1397,In_1423,In_28);
and U1398 (N_1398,In_1455,In_204);
nand U1399 (N_1399,In_797,In_1286);
and U1400 (N_1400,In_1942,In_1120);
and U1401 (N_1401,In_1201,In_2093);
or U1402 (N_1402,In_1584,In_1711);
and U1403 (N_1403,In_1393,In_34);
nand U1404 (N_1404,In_1488,In_1952);
nor U1405 (N_1405,In_1748,In_1699);
or U1406 (N_1406,In_966,In_732);
xor U1407 (N_1407,In_1278,In_957);
or U1408 (N_1408,In_405,In_1838);
nor U1409 (N_1409,In_2007,In_1364);
and U1410 (N_1410,In_1060,In_701);
nor U1411 (N_1411,In_2352,In_1280);
nor U1412 (N_1412,In_885,In_1385);
or U1413 (N_1413,In_2461,In_1032);
and U1414 (N_1414,In_1092,In_2447);
nand U1415 (N_1415,In_1222,In_1611);
and U1416 (N_1416,In_271,In_1195);
or U1417 (N_1417,In_1736,In_2464);
nand U1418 (N_1418,In_2271,In_2338);
and U1419 (N_1419,In_1727,In_873);
and U1420 (N_1420,In_481,In_1355);
and U1421 (N_1421,In_1178,In_472);
and U1422 (N_1422,In_414,In_1784);
nor U1423 (N_1423,In_1648,In_554);
and U1424 (N_1424,In_601,In_1876);
nor U1425 (N_1425,In_1195,In_197);
and U1426 (N_1426,In_1482,In_348);
and U1427 (N_1427,In_598,In_367);
or U1428 (N_1428,In_2382,In_1919);
nand U1429 (N_1429,In_1922,In_806);
nand U1430 (N_1430,In_125,In_2047);
and U1431 (N_1431,In_452,In_2206);
nor U1432 (N_1432,In_1351,In_551);
nor U1433 (N_1433,In_194,In_486);
nor U1434 (N_1434,In_2295,In_1906);
or U1435 (N_1435,In_363,In_694);
or U1436 (N_1436,In_847,In_972);
and U1437 (N_1437,In_2363,In_945);
nand U1438 (N_1438,In_59,In_670);
or U1439 (N_1439,In_740,In_1034);
nor U1440 (N_1440,In_595,In_1057);
or U1441 (N_1441,In_1044,In_2441);
or U1442 (N_1442,In_510,In_1024);
and U1443 (N_1443,In_917,In_1895);
or U1444 (N_1444,In_1772,In_1075);
or U1445 (N_1445,In_1604,In_231);
nand U1446 (N_1446,In_2257,In_607);
and U1447 (N_1447,In_240,In_2411);
or U1448 (N_1448,In_1481,In_1610);
and U1449 (N_1449,In_151,In_1553);
and U1450 (N_1450,In_1461,In_543);
and U1451 (N_1451,In_1120,In_1410);
and U1452 (N_1452,In_521,In_983);
and U1453 (N_1453,In_2158,In_214);
nand U1454 (N_1454,In_2204,In_1622);
nor U1455 (N_1455,In_235,In_1695);
nor U1456 (N_1456,In_2265,In_1255);
or U1457 (N_1457,In_120,In_1404);
nand U1458 (N_1458,In_2144,In_518);
nor U1459 (N_1459,In_254,In_1774);
nand U1460 (N_1460,In_1363,In_366);
or U1461 (N_1461,In_1471,In_1635);
or U1462 (N_1462,In_738,In_982);
nor U1463 (N_1463,In_679,In_1006);
or U1464 (N_1464,In_1339,In_625);
and U1465 (N_1465,In_782,In_830);
or U1466 (N_1466,In_1660,In_819);
nand U1467 (N_1467,In_432,In_452);
or U1468 (N_1468,In_387,In_875);
nand U1469 (N_1469,In_2267,In_241);
and U1470 (N_1470,In_862,In_2083);
nor U1471 (N_1471,In_1379,In_1380);
and U1472 (N_1472,In_1083,In_2412);
nand U1473 (N_1473,In_2119,In_1647);
nand U1474 (N_1474,In_1219,In_1811);
and U1475 (N_1475,In_1172,In_102);
or U1476 (N_1476,In_2474,In_667);
xnor U1477 (N_1477,In_1806,In_1074);
and U1478 (N_1478,In_1751,In_762);
nand U1479 (N_1479,In_261,In_694);
nand U1480 (N_1480,In_624,In_1680);
nand U1481 (N_1481,In_682,In_1751);
and U1482 (N_1482,In_1087,In_18);
or U1483 (N_1483,In_338,In_263);
or U1484 (N_1484,In_905,In_84);
nand U1485 (N_1485,In_2499,In_1345);
and U1486 (N_1486,In_2123,In_231);
nor U1487 (N_1487,In_1704,In_1657);
and U1488 (N_1488,In_33,In_589);
and U1489 (N_1489,In_45,In_622);
or U1490 (N_1490,In_1937,In_1562);
nand U1491 (N_1491,In_1845,In_1852);
and U1492 (N_1492,In_1631,In_1233);
or U1493 (N_1493,In_1475,In_2124);
and U1494 (N_1494,In_276,In_1218);
nand U1495 (N_1495,In_1744,In_492);
xor U1496 (N_1496,In_2012,In_2138);
or U1497 (N_1497,In_1434,In_2344);
nand U1498 (N_1498,In_1129,In_1919);
or U1499 (N_1499,In_1818,In_1250);
or U1500 (N_1500,In_375,In_804);
nand U1501 (N_1501,In_1115,In_1345);
or U1502 (N_1502,In_721,In_767);
and U1503 (N_1503,In_2456,In_1676);
or U1504 (N_1504,In_362,In_1200);
or U1505 (N_1505,In_1484,In_2207);
nand U1506 (N_1506,In_858,In_2226);
or U1507 (N_1507,In_2090,In_2376);
and U1508 (N_1508,In_1893,In_2178);
nor U1509 (N_1509,In_2050,In_854);
nand U1510 (N_1510,In_1673,In_851);
nor U1511 (N_1511,In_28,In_2455);
and U1512 (N_1512,In_1321,In_739);
or U1513 (N_1513,In_1759,In_2370);
nand U1514 (N_1514,In_135,In_1196);
or U1515 (N_1515,In_1975,In_1345);
or U1516 (N_1516,In_317,In_2496);
nor U1517 (N_1517,In_1550,In_643);
and U1518 (N_1518,In_951,In_275);
nand U1519 (N_1519,In_1984,In_2400);
or U1520 (N_1520,In_2235,In_2315);
xnor U1521 (N_1521,In_1250,In_2127);
nand U1522 (N_1522,In_719,In_303);
and U1523 (N_1523,In_222,In_652);
xnor U1524 (N_1524,In_1855,In_946);
nor U1525 (N_1525,In_1348,In_1754);
nor U1526 (N_1526,In_1443,In_123);
or U1527 (N_1527,In_2497,In_1653);
and U1528 (N_1528,In_2020,In_841);
or U1529 (N_1529,In_2066,In_470);
nand U1530 (N_1530,In_1808,In_1908);
nand U1531 (N_1531,In_1085,In_1214);
or U1532 (N_1532,In_607,In_1500);
nand U1533 (N_1533,In_126,In_1018);
nand U1534 (N_1534,In_24,In_1731);
and U1535 (N_1535,In_2146,In_1601);
nor U1536 (N_1536,In_732,In_1300);
nand U1537 (N_1537,In_2468,In_1134);
and U1538 (N_1538,In_469,In_1928);
or U1539 (N_1539,In_2405,In_1246);
and U1540 (N_1540,In_1762,In_2480);
and U1541 (N_1541,In_2257,In_310);
or U1542 (N_1542,In_2108,In_952);
nor U1543 (N_1543,In_2488,In_766);
or U1544 (N_1544,In_2359,In_1194);
nor U1545 (N_1545,In_1830,In_1707);
nor U1546 (N_1546,In_611,In_1834);
nor U1547 (N_1547,In_56,In_1425);
nor U1548 (N_1548,In_499,In_872);
or U1549 (N_1549,In_3,In_1192);
or U1550 (N_1550,In_197,In_896);
and U1551 (N_1551,In_312,In_1432);
and U1552 (N_1552,In_258,In_2175);
nand U1553 (N_1553,In_1172,In_95);
nand U1554 (N_1554,In_1623,In_168);
and U1555 (N_1555,In_1035,In_2202);
or U1556 (N_1556,In_1572,In_38);
nor U1557 (N_1557,In_84,In_1726);
xnor U1558 (N_1558,In_1376,In_690);
nor U1559 (N_1559,In_358,In_292);
or U1560 (N_1560,In_1072,In_2222);
nand U1561 (N_1561,In_2374,In_1401);
or U1562 (N_1562,In_640,In_1214);
nor U1563 (N_1563,In_2115,In_1827);
nand U1564 (N_1564,In_1454,In_2474);
and U1565 (N_1565,In_380,In_1693);
and U1566 (N_1566,In_1349,In_1544);
or U1567 (N_1567,In_374,In_2452);
and U1568 (N_1568,In_1273,In_2001);
and U1569 (N_1569,In_2419,In_127);
or U1570 (N_1570,In_306,In_977);
and U1571 (N_1571,In_1706,In_2326);
xor U1572 (N_1572,In_327,In_115);
and U1573 (N_1573,In_281,In_2265);
nand U1574 (N_1574,In_1403,In_1771);
or U1575 (N_1575,In_1246,In_1687);
or U1576 (N_1576,In_228,In_988);
nor U1577 (N_1577,In_2056,In_1852);
nand U1578 (N_1578,In_1724,In_966);
or U1579 (N_1579,In_555,In_1487);
or U1580 (N_1580,In_1666,In_2286);
nand U1581 (N_1581,In_2152,In_391);
xor U1582 (N_1582,In_1052,In_408);
nor U1583 (N_1583,In_1690,In_538);
nand U1584 (N_1584,In_922,In_463);
nand U1585 (N_1585,In_1938,In_437);
nand U1586 (N_1586,In_36,In_427);
or U1587 (N_1587,In_2258,In_667);
and U1588 (N_1588,In_2411,In_2480);
or U1589 (N_1589,In_1930,In_31);
nand U1590 (N_1590,In_498,In_2018);
nor U1591 (N_1591,In_730,In_662);
or U1592 (N_1592,In_1692,In_96);
and U1593 (N_1593,In_2169,In_458);
nand U1594 (N_1594,In_1105,In_976);
and U1595 (N_1595,In_1508,In_1127);
nand U1596 (N_1596,In_55,In_818);
xnor U1597 (N_1597,In_190,In_1478);
nand U1598 (N_1598,In_1177,In_1712);
nor U1599 (N_1599,In_1795,In_1925);
nand U1600 (N_1600,In_1358,In_734);
and U1601 (N_1601,In_1046,In_1919);
nor U1602 (N_1602,In_2073,In_1051);
nor U1603 (N_1603,In_2416,In_2167);
nor U1604 (N_1604,In_175,In_130);
xor U1605 (N_1605,In_2043,In_1236);
or U1606 (N_1606,In_2297,In_1264);
nand U1607 (N_1607,In_657,In_2108);
or U1608 (N_1608,In_562,In_1516);
nor U1609 (N_1609,In_1295,In_1663);
and U1610 (N_1610,In_387,In_1887);
or U1611 (N_1611,In_545,In_620);
and U1612 (N_1612,In_247,In_497);
nor U1613 (N_1613,In_1622,In_1302);
or U1614 (N_1614,In_645,In_311);
xor U1615 (N_1615,In_2457,In_97);
or U1616 (N_1616,In_1362,In_1450);
nand U1617 (N_1617,In_1772,In_184);
and U1618 (N_1618,In_1221,In_1387);
and U1619 (N_1619,In_1313,In_1160);
nor U1620 (N_1620,In_1336,In_1574);
nor U1621 (N_1621,In_82,In_1454);
nor U1622 (N_1622,In_517,In_972);
or U1623 (N_1623,In_396,In_236);
nor U1624 (N_1624,In_2198,In_2404);
or U1625 (N_1625,In_514,In_344);
nor U1626 (N_1626,In_374,In_1241);
nor U1627 (N_1627,In_165,In_2467);
or U1628 (N_1628,In_1226,In_2163);
nor U1629 (N_1629,In_2305,In_1271);
and U1630 (N_1630,In_306,In_378);
nand U1631 (N_1631,In_1177,In_244);
nor U1632 (N_1632,In_415,In_1212);
or U1633 (N_1633,In_1863,In_220);
nor U1634 (N_1634,In_928,In_1256);
or U1635 (N_1635,In_1708,In_1051);
and U1636 (N_1636,In_950,In_2148);
and U1637 (N_1637,In_550,In_457);
or U1638 (N_1638,In_1209,In_793);
nor U1639 (N_1639,In_1038,In_1345);
and U1640 (N_1640,In_1808,In_1878);
nand U1641 (N_1641,In_716,In_1647);
or U1642 (N_1642,In_2341,In_1111);
and U1643 (N_1643,In_2264,In_1130);
nand U1644 (N_1644,In_1146,In_2317);
nor U1645 (N_1645,In_2475,In_506);
and U1646 (N_1646,In_1556,In_1455);
nor U1647 (N_1647,In_1946,In_1868);
or U1648 (N_1648,In_1455,In_1729);
nand U1649 (N_1649,In_46,In_302);
and U1650 (N_1650,In_2220,In_1876);
nand U1651 (N_1651,In_28,In_871);
nor U1652 (N_1652,In_547,In_1563);
nor U1653 (N_1653,In_1211,In_1786);
or U1654 (N_1654,In_1100,In_273);
nand U1655 (N_1655,In_260,In_1677);
and U1656 (N_1656,In_418,In_717);
nor U1657 (N_1657,In_1260,In_1084);
or U1658 (N_1658,In_1357,In_1753);
nor U1659 (N_1659,In_700,In_1380);
nor U1660 (N_1660,In_1682,In_1953);
nand U1661 (N_1661,In_530,In_1820);
and U1662 (N_1662,In_883,In_1963);
or U1663 (N_1663,In_861,In_1966);
xnor U1664 (N_1664,In_1953,In_1320);
xor U1665 (N_1665,In_241,In_1807);
and U1666 (N_1666,In_1642,In_1495);
or U1667 (N_1667,In_973,In_1541);
nand U1668 (N_1668,In_2036,In_1594);
nor U1669 (N_1669,In_2235,In_2021);
nor U1670 (N_1670,In_1108,In_355);
nor U1671 (N_1671,In_930,In_2214);
or U1672 (N_1672,In_1234,In_145);
nand U1673 (N_1673,In_989,In_1783);
xor U1674 (N_1674,In_1080,In_1633);
or U1675 (N_1675,In_1732,In_896);
and U1676 (N_1676,In_1840,In_773);
or U1677 (N_1677,In_375,In_193);
nand U1678 (N_1678,In_521,In_1952);
or U1679 (N_1679,In_132,In_1959);
and U1680 (N_1680,In_752,In_2041);
xor U1681 (N_1681,In_1610,In_310);
nor U1682 (N_1682,In_992,In_511);
nand U1683 (N_1683,In_2420,In_1479);
or U1684 (N_1684,In_2405,In_2188);
or U1685 (N_1685,In_2318,In_1285);
nand U1686 (N_1686,In_2320,In_2339);
nor U1687 (N_1687,In_408,In_1135);
nand U1688 (N_1688,In_337,In_1742);
or U1689 (N_1689,In_1058,In_1284);
nand U1690 (N_1690,In_2300,In_337);
nand U1691 (N_1691,In_1930,In_1337);
nor U1692 (N_1692,In_1845,In_1040);
or U1693 (N_1693,In_986,In_1953);
or U1694 (N_1694,In_467,In_1806);
nor U1695 (N_1695,In_2001,In_584);
nor U1696 (N_1696,In_1710,In_1793);
and U1697 (N_1697,In_1828,In_125);
or U1698 (N_1698,In_639,In_2026);
or U1699 (N_1699,In_1729,In_620);
nor U1700 (N_1700,In_638,In_197);
nand U1701 (N_1701,In_1833,In_907);
nand U1702 (N_1702,In_759,In_969);
and U1703 (N_1703,In_970,In_518);
nor U1704 (N_1704,In_1672,In_2067);
or U1705 (N_1705,In_100,In_1231);
nand U1706 (N_1706,In_696,In_785);
and U1707 (N_1707,In_1611,In_585);
nor U1708 (N_1708,In_1397,In_2210);
nand U1709 (N_1709,In_1429,In_1609);
and U1710 (N_1710,In_1801,In_489);
nor U1711 (N_1711,In_693,In_2193);
and U1712 (N_1712,In_875,In_1932);
and U1713 (N_1713,In_414,In_1691);
nand U1714 (N_1714,In_1885,In_1712);
nand U1715 (N_1715,In_586,In_1445);
or U1716 (N_1716,In_361,In_2174);
nand U1717 (N_1717,In_298,In_2410);
nand U1718 (N_1718,In_41,In_366);
xnor U1719 (N_1719,In_920,In_2183);
or U1720 (N_1720,In_1327,In_236);
or U1721 (N_1721,In_2112,In_2056);
and U1722 (N_1722,In_83,In_2300);
nand U1723 (N_1723,In_1688,In_1585);
or U1724 (N_1724,In_213,In_1639);
nand U1725 (N_1725,In_2145,In_1989);
nand U1726 (N_1726,In_380,In_1334);
nand U1727 (N_1727,In_1277,In_726);
or U1728 (N_1728,In_1528,In_135);
and U1729 (N_1729,In_138,In_87);
and U1730 (N_1730,In_2365,In_2376);
and U1731 (N_1731,In_2282,In_869);
nor U1732 (N_1732,In_865,In_1459);
and U1733 (N_1733,In_642,In_830);
or U1734 (N_1734,In_656,In_2440);
nand U1735 (N_1735,In_2211,In_1242);
or U1736 (N_1736,In_2074,In_2454);
nand U1737 (N_1737,In_514,In_86);
nor U1738 (N_1738,In_1005,In_1269);
or U1739 (N_1739,In_1757,In_1279);
and U1740 (N_1740,In_1668,In_2363);
and U1741 (N_1741,In_335,In_787);
or U1742 (N_1742,In_1718,In_464);
or U1743 (N_1743,In_1032,In_2409);
nand U1744 (N_1744,In_1166,In_1628);
nand U1745 (N_1745,In_2204,In_1348);
nand U1746 (N_1746,In_1058,In_1684);
nor U1747 (N_1747,In_699,In_2379);
and U1748 (N_1748,In_1134,In_1773);
nand U1749 (N_1749,In_718,In_648);
or U1750 (N_1750,In_2437,In_194);
nand U1751 (N_1751,In_1105,In_1857);
nor U1752 (N_1752,In_1456,In_1591);
and U1753 (N_1753,In_564,In_507);
nor U1754 (N_1754,In_93,In_515);
and U1755 (N_1755,In_1231,In_1665);
and U1756 (N_1756,In_1635,In_2289);
or U1757 (N_1757,In_2296,In_1425);
xnor U1758 (N_1758,In_1044,In_568);
and U1759 (N_1759,In_922,In_1135);
or U1760 (N_1760,In_1363,In_685);
nor U1761 (N_1761,In_1108,In_1661);
and U1762 (N_1762,In_2136,In_2420);
or U1763 (N_1763,In_2365,In_1860);
nand U1764 (N_1764,In_269,In_2152);
xnor U1765 (N_1765,In_2183,In_1267);
and U1766 (N_1766,In_931,In_2420);
or U1767 (N_1767,In_869,In_354);
nand U1768 (N_1768,In_2369,In_126);
or U1769 (N_1769,In_1659,In_1718);
nand U1770 (N_1770,In_2013,In_264);
nor U1771 (N_1771,In_1547,In_511);
nor U1772 (N_1772,In_1715,In_1599);
and U1773 (N_1773,In_128,In_2473);
and U1774 (N_1774,In_2112,In_161);
and U1775 (N_1775,In_2148,In_2138);
nor U1776 (N_1776,In_2160,In_66);
and U1777 (N_1777,In_536,In_1163);
nand U1778 (N_1778,In_2275,In_1121);
nor U1779 (N_1779,In_1056,In_1468);
xor U1780 (N_1780,In_153,In_2217);
or U1781 (N_1781,In_403,In_1188);
nor U1782 (N_1782,In_1654,In_1037);
or U1783 (N_1783,In_2082,In_1389);
or U1784 (N_1784,In_1898,In_2428);
nor U1785 (N_1785,In_1441,In_2457);
or U1786 (N_1786,In_141,In_2220);
or U1787 (N_1787,In_2235,In_1666);
nor U1788 (N_1788,In_339,In_1931);
and U1789 (N_1789,In_2023,In_1929);
nand U1790 (N_1790,In_1021,In_462);
nor U1791 (N_1791,In_496,In_2264);
and U1792 (N_1792,In_1008,In_1998);
or U1793 (N_1793,In_1595,In_736);
and U1794 (N_1794,In_245,In_939);
or U1795 (N_1795,In_370,In_982);
and U1796 (N_1796,In_509,In_1621);
or U1797 (N_1797,In_1419,In_1297);
nand U1798 (N_1798,In_2240,In_1488);
nand U1799 (N_1799,In_2280,In_989);
nand U1800 (N_1800,In_211,In_2498);
nor U1801 (N_1801,In_2156,In_850);
nand U1802 (N_1802,In_1952,In_343);
or U1803 (N_1803,In_2030,In_322);
nor U1804 (N_1804,In_995,In_1091);
nand U1805 (N_1805,In_1809,In_2338);
xnor U1806 (N_1806,In_1851,In_1586);
and U1807 (N_1807,In_2091,In_1326);
nand U1808 (N_1808,In_176,In_1807);
nand U1809 (N_1809,In_2228,In_1399);
nand U1810 (N_1810,In_2493,In_1015);
nand U1811 (N_1811,In_1596,In_2232);
or U1812 (N_1812,In_2062,In_5);
nor U1813 (N_1813,In_1943,In_1214);
nor U1814 (N_1814,In_697,In_1493);
or U1815 (N_1815,In_1968,In_872);
nand U1816 (N_1816,In_375,In_1025);
nand U1817 (N_1817,In_919,In_1674);
and U1818 (N_1818,In_666,In_637);
and U1819 (N_1819,In_1490,In_767);
and U1820 (N_1820,In_283,In_764);
or U1821 (N_1821,In_84,In_1503);
and U1822 (N_1822,In_1269,In_218);
nand U1823 (N_1823,In_1571,In_2431);
nor U1824 (N_1824,In_1245,In_41);
nor U1825 (N_1825,In_2282,In_1767);
nand U1826 (N_1826,In_555,In_33);
and U1827 (N_1827,In_100,In_808);
or U1828 (N_1828,In_1088,In_2010);
nand U1829 (N_1829,In_190,In_2322);
or U1830 (N_1830,In_2009,In_1869);
nand U1831 (N_1831,In_1769,In_2278);
or U1832 (N_1832,In_296,In_1036);
and U1833 (N_1833,In_157,In_766);
nor U1834 (N_1834,In_1503,In_1634);
nor U1835 (N_1835,In_2041,In_330);
nand U1836 (N_1836,In_1664,In_2300);
or U1837 (N_1837,In_1661,In_1480);
nand U1838 (N_1838,In_2196,In_1628);
nor U1839 (N_1839,In_1902,In_1912);
nand U1840 (N_1840,In_2383,In_413);
or U1841 (N_1841,In_1844,In_2381);
nand U1842 (N_1842,In_1788,In_1085);
xnor U1843 (N_1843,In_1496,In_1515);
nor U1844 (N_1844,In_1064,In_1914);
or U1845 (N_1845,In_1475,In_1717);
nand U1846 (N_1846,In_664,In_1048);
nand U1847 (N_1847,In_1963,In_401);
or U1848 (N_1848,In_429,In_1854);
nand U1849 (N_1849,In_1121,In_237);
and U1850 (N_1850,In_1183,In_1943);
and U1851 (N_1851,In_2208,In_831);
xor U1852 (N_1852,In_252,In_272);
and U1853 (N_1853,In_298,In_1667);
or U1854 (N_1854,In_1367,In_1928);
or U1855 (N_1855,In_1007,In_719);
or U1856 (N_1856,In_448,In_1435);
or U1857 (N_1857,In_1390,In_1701);
nor U1858 (N_1858,In_64,In_1908);
or U1859 (N_1859,In_1674,In_1564);
and U1860 (N_1860,In_138,In_2374);
nor U1861 (N_1861,In_1153,In_435);
and U1862 (N_1862,In_2213,In_2297);
nor U1863 (N_1863,In_429,In_512);
nand U1864 (N_1864,In_2373,In_635);
nor U1865 (N_1865,In_1326,In_1945);
and U1866 (N_1866,In_1425,In_2139);
nand U1867 (N_1867,In_2215,In_2033);
or U1868 (N_1868,In_1874,In_992);
nor U1869 (N_1869,In_75,In_2475);
and U1870 (N_1870,In_1551,In_2381);
and U1871 (N_1871,In_2074,In_511);
nor U1872 (N_1872,In_2183,In_2027);
or U1873 (N_1873,In_1929,In_1586);
and U1874 (N_1874,In_1315,In_967);
nand U1875 (N_1875,In_2102,In_1428);
nand U1876 (N_1876,In_453,In_17);
or U1877 (N_1877,In_1764,In_2294);
nand U1878 (N_1878,In_1219,In_1696);
and U1879 (N_1879,In_218,In_1434);
or U1880 (N_1880,In_1702,In_472);
nand U1881 (N_1881,In_876,In_1952);
or U1882 (N_1882,In_720,In_1570);
or U1883 (N_1883,In_1366,In_30);
nand U1884 (N_1884,In_664,In_500);
and U1885 (N_1885,In_1217,In_297);
nand U1886 (N_1886,In_742,In_1182);
and U1887 (N_1887,In_2296,In_1856);
nor U1888 (N_1888,In_1596,In_799);
nand U1889 (N_1889,In_209,In_1352);
nor U1890 (N_1890,In_1748,In_827);
or U1891 (N_1891,In_407,In_2284);
and U1892 (N_1892,In_339,In_1690);
nand U1893 (N_1893,In_2243,In_2379);
nand U1894 (N_1894,In_1107,In_1733);
or U1895 (N_1895,In_2458,In_665);
nand U1896 (N_1896,In_2130,In_2365);
nor U1897 (N_1897,In_1854,In_1717);
and U1898 (N_1898,In_468,In_1766);
or U1899 (N_1899,In_1900,In_638);
nor U1900 (N_1900,In_2491,In_2063);
or U1901 (N_1901,In_737,In_1016);
nand U1902 (N_1902,In_244,In_1950);
or U1903 (N_1903,In_167,In_1808);
nor U1904 (N_1904,In_877,In_281);
or U1905 (N_1905,In_580,In_914);
nand U1906 (N_1906,In_295,In_1498);
nor U1907 (N_1907,In_541,In_339);
nor U1908 (N_1908,In_1791,In_1689);
nand U1909 (N_1909,In_1534,In_933);
nor U1910 (N_1910,In_1623,In_2192);
or U1911 (N_1911,In_1645,In_1191);
and U1912 (N_1912,In_1162,In_2498);
nor U1913 (N_1913,In_2406,In_282);
nand U1914 (N_1914,In_42,In_281);
or U1915 (N_1915,In_1338,In_1380);
or U1916 (N_1916,In_2361,In_693);
nand U1917 (N_1917,In_938,In_684);
nand U1918 (N_1918,In_367,In_930);
nor U1919 (N_1919,In_1018,In_2058);
nor U1920 (N_1920,In_2175,In_1354);
or U1921 (N_1921,In_600,In_733);
nor U1922 (N_1922,In_1061,In_1219);
or U1923 (N_1923,In_1083,In_365);
or U1924 (N_1924,In_32,In_1685);
and U1925 (N_1925,In_72,In_1075);
nor U1926 (N_1926,In_314,In_2157);
nand U1927 (N_1927,In_1058,In_1539);
nor U1928 (N_1928,In_1050,In_2112);
nand U1929 (N_1929,In_1623,In_1568);
nor U1930 (N_1930,In_1398,In_1173);
and U1931 (N_1931,In_2254,In_1619);
nor U1932 (N_1932,In_1695,In_2333);
xnor U1933 (N_1933,In_1702,In_2411);
nor U1934 (N_1934,In_2167,In_1588);
nor U1935 (N_1935,In_2348,In_822);
or U1936 (N_1936,In_825,In_58);
nand U1937 (N_1937,In_675,In_47);
nor U1938 (N_1938,In_543,In_823);
nor U1939 (N_1939,In_166,In_1344);
or U1940 (N_1940,In_1688,In_1206);
nor U1941 (N_1941,In_2478,In_1850);
and U1942 (N_1942,In_201,In_539);
and U1943 (N_1943,In_118,In_1296);
nor U1944 (N_1944,In_1323,In_1893);
or U1945 (N_1945,In_1380,In_284);
nor U1946 (N_1946,In_1239,In_1388);
nand U1947 (N_1947,In_703,In_2268);
nand U1948 (N_1948,In_1152,In_956);
nand U1949 (N_1949,In_483,In_624);
or U1950 (N_1950,In_74,In_323);
or U1951 (N_1951,In_1967,In_2113);
nor U1952 (N_1952,In_167,In_1843);
nor U1953 (N_1953,In_1384,In_793);
and U1954 (N_1954,In_2051,In_161);
nor U1955 (N_1955,In_2351,In_1718);
or U1956 (N_1956,In_2243,In_1334);
and U1957 (N_1957,In_1262,In_252);
nor U1958 (N_1958,In_2071,In_1463);
or U1959 (N_1959,In_2209,In_2373);
nand U1960 (N_1960,In_1235,In_1681);
and U1961 (N_1961,In_1851,In_509);
nor U1962 (N_1962,In_1321,In_94);
nor U1963 (N_1963,In_2352,In_575);
and U1964 (N_1964,In_954,In_2006);
nor U1965 (N_1965,In_1366,In_88);
or U1966 (N_1966,In_1301,In_2003);
nand U1967 (N_1967,In_1439,In_1410);
nor U1968 (N_1968,In_212,In_1719);
and U1969 (N_1969,In_833,In_344);
or U1970 (N_1970,In_2251,In_33);
nand U1971 (N_1971,In_1106,In_784);
nand U1972 (N_1972,In_516,In_553);
nand U1973 (N_1973,In_2033,In_1700);
or U1974 (N_1974,In_594,In_388);
or U1975 (N_1975,In_2089,In_2071);
and U1976 (N_1976,In_1158,In_28);
nand U1977 (N_1977,In_551,In_559);
and U1978 (N_1978,In_26,In_44);
or U1979 (N_1979,In_1597,In_1756);
nor U1980 (N_1980,In_1366,In_1375);
nor U1981 (N_1981,In_195,In_630);
and U1982 (N_1982,In_1837,In_1395);
nor U1983 (N_1983,In_2380,In_2376);
nand U1984 (N_1984,In_458,In_2181);
xor U1985 (N_1985,In_2059,In_1502);
or U1986 (N_1986,In_1848,In_292);
and U1987 (N_1987,In_266,In_33);
nor U1988 (N_1988,In_2124,In_1646);
and U1989 (N_1989,In_370,In_1720);
nand U1990 (N_1990,In_1243,In_1495);
nor U1991 (N_1991,In_1678,In_302);
and U1992 (N_1992,In_890,In_428);
or U1993 (N_1993,In_1857,In_2093);
xor U1994 (N_1994,In_745,In_1299);
and U1995 (N_1995,In_917,In_2049);
or U1996 (N_1996,In_2197,In_236);
nor U1997 (N_1997,In_820,In_564);
or U1998 (N_1998,In_96,In_609);
nor U1999 (N_1999,In_564,In_69);
xnor U2000 (N_2000,In_2499,In_378);
nor U2001 (N_2001,In_589,In_775);
and U2002 (N_2002,In_764,In_630);
and U2003 (N_2003,In_69,In_834);
nor U2004 (N_2004,In_458,In_1753);
or U2005 (N_2005,In_1248,In_2246);
and U2006 (N_2006,In_1714,In_618);
nor U2007 (N_2007,In_948,In_960);
or U2008 (N_2008,In_2288,In_2218);
nand U2009 (N_2009,In_996,In_784);
nand U2010 (N_2010,In_2194,In_1194);
xor U2011 (N_2011,In_822,In_355);
xnor U2012 (N_2012,In_1343,In_1261);
nor U2013 (N_2013,In_2370,In_136);
nand U2014 (N_2014,In_1432,In_1787);
nor U2015 (N_2015,In_1123,In_185);
nand U2016 (N_2016,In_363,In_2287);
nor U2017 (N_2017,In_469,In_2200);
and U2018 (N_2018,In_2283,In_1692);
nand U2019 (N_2019,In_1525,In_1355);
and U2020 (N_2020,In_1876,In_2145);
nand U2021 (N_2021,In_360,In_1543);
nand U2022 (N_2022,In_2496,In_2276);
and U2023 (N_2023,In_152,In_1921);
nand U2024 (N_2024,In_1677,In_2486);
xor U2025 (N_2025,In_1693,In_1581);
or U2026 (N_2026,In_1977,In_1378);
or U2027 (N_2027,In_1024,In_551);
nand U2028 (N_2028,In_294,In_154);
and U2029 (N_2029,In_625,In_1529);
and U2030 (N_2030,In_1738,In_1488);
nor U2031 (N_2031,In_2117,In_2044);
nor U2032 (N_2032,In_1704,In_2144);
nand U2033 (N_2033,In_833,In_1292);
or U2034 (N_2034,In_798,In_1173);
nand U2035 (N_2035,In_1873,In_224);
and U2036 (N_2036,In_1924,In_2260);
nor U2037 (N_2037,In_2486,In_1434);
nand U2038 (N_2038,In_2200,In_1228);
xor U2039 (N_2039,In_708,In_2190);
nor U2040 (N_2040,In_214,In_2196);
and U2041 (N_2041,In_789,In_1144);
nor U2042 (N_2042,In_37,In_2064);
or U2043 (N_2043,In_583,In_1784);
nand U2044 (N_2044,In_1349,In_268);
or U2045 (N_2045,In_890,In_1640);
or U2046 (N_2046,In_1814,In_85);
or U2047 (N_2047,In_1131,In_1404);
or U2048 (N_2048,In_1460,In_755);
nor U2049 (N_2049,In_143,In_2057);
and U2050 (N_2050,In_402,In_416);
and U2051 (N_2051,In_1856,In_1286);
or U2052 (N_2052,In_1324,In_570);
and U2053 (N_2053,In_1566,In_362);
or U2054 (N_2054,In_1380,In_433);
nor U2055 (N_2055,In_1805,In_2043);
nand U2056 (N_2056,In_1581,In_1649);
or U2057 (N_2057,In_248,In_1657);
or U2058 (N_2058,In_989,In_979);
nand U2059 (N_2059,In_980,In_2347);
or U2060 (N_2060,In_2307,In_8);
nand U2061 (N_2061,In_80,In_1196);
nand U2062 (N_2062,In_1554,In_2317);
xnor U2063 (N_2063,In_1273,In_970);
or U2064 (N_2064,In_2288,In_1103);
nor U2065 (N_2065,In_1992,In_694);
nor U2066 (N_2066,In_1267,In_783);
or U2067 (N_2067,In_1552,In_95);
nand U2068 (N_2068,In_236,In_1847);
nand U2069 (N_2069,In_946,In_44);
or U2070 (N_2070,In_945,In_2370);
or U2071 (N_2071,In_884,In_727);
and U2072 (N_2072,In_544,In_2308);
or U2073 (N_2073,In_809,In_768);
nor U2074 (N_2074,In_883,In_898);
nand U2075 (N_2075,In_1782,In_1518);
nand U2076 (N_2076,In_1285,In_515);
nand U2077 (N_2077,In_958,In_1286);
and U2078 (N_2078,In_905,In_1641);
nor U2079 (N_2079,In_1785,In_2077);
or U2080 (N_2080,In_2462,In_1029);
or U2081 (N_2081,In_1480,In_1848);
and U2082 (N_2082,In_1839,In_1387);
nand U2083 (N_2083,In_403,In_953);
and U2084 (N_2084,In_959,In_1278);
and U2085 (N_2085,In_2093,In_2478);
xnor U2086 (N_2086,In_63,In_108);
or U2087 (N_2087,In_734,In_1812);
and U2088 (N_2088,In_761,In_1096);
or U2089 (N_2089,In_2009,In_1786);
and U2090 (N_2090,In_1626,In_1916);
and U2091 (N_2091,In_651,In_1895);
nand U2092 (N_2092,In_222,In_840);
nor U2093 (N_2093,In_623,In_1169);
or U2094 (N_2094,In_55,In_1854);
or U2095 (N_2095,In_2478,In_2425);
and U2096 (N_2096,In_2134,In_1654);
or U2097 (N_2097,In_2038,In_378);
and U2098 (N_2098,In_2090,In_1448);
nor U2099 (N_2099,In_641,In_2101);
nor U2100 (N_2100,In_1564,In_276);
nor U2101 (N_2101,In_1719,In_2062);
or U2102 (N_2102,In_1127,In_1825);
or U2103 (N_2103,In_1619,In_386);
nand U2104 (N_2104,In_1569,In_438);
or U2105 (N_2105,In_2377,In_1616);
nor U2106 (N_2106,In_1420,In_465);
and U2107 (N_2107,In_1329,In_2422);
and U2108 (N_2108,In_2248,In_484);
nor U2109 (N_2109,In_1756,In_1454);
or U2110 (N_2110,In_1846,In_1935);
or U2111 (N_2111,In_215,In_1595);
nor U2112 (N_2112,In_2237,In_1353);
nand U2113 (N_2113,In_2260,In_1297);
nor U2114 (N_2114,In_62,In_2077);
nand U2115 (N_2115,In_1921,In_110);
nand U2116 (N_2116,In_1620,In_1578);
nor U2117 (N_2117,In_498,In_1853);
nor U2118 (N_2118,In_2145,In_2226);
and U2119 (N_2119,In_558,In_215);
nand U2120 (N_2120,In_2391,In_2123);
and U2121 (N_2121,In_319,In_1656);
or U2122 (N_2122,In_399,In_1289);
nor U2123 (N_2123,In_128,In_402);
nor U2124 (N_2124,In_1431,In_701);
nand U2125 (N_2125,In_904,In_401);
nand U2126 (N_2126,In_1617,In_2171);
and U2127 (N_2127,In_663,In_359);
and U2128 (N_2128,In_1428,In_1950);
nor U2129 (N_2129,In_105,In_1974);
or U2130 (N_2130,In_2289,In_245);
and U2131 (N_2131,In_2432,In_218);
and U2132 (N_2132,In_2421,In_277);
and U2133 (N_2133,In_1703,In_3);
or U2134 (N_2134,In_1730,In_1958);
nand U2135 (N_2135,In_2442,In_406);
or U2136 (N_2136,In_779,In_1868);
nand U2137 (N_2137,In_934,In_442);
or U2138 (N_2138,In_2460,In_296);
xnor U2139 (N_2139,In_1492,In_1286);
nor U2140 (N_2140,In_1921,In_1236);
or U2141 (N_2141,In_1814,In_1930);
and U2142 (N_2142,In_682,In_1570);
nand U2143 (N_2143,In_885,In_1434);
nor U2144 (N_2144,In_1714,In_2144);
or U2145 (N_2145,In_1252,In_540);
nor U2146 (N_2146,In_1767,In_1488);
nor U2147 (N_2147,In_2143,In_1140);
and U2148 (N_2148,In_550,In_756);
nor U2149 (N_2149,In_98,In_1480);
and U2150 (N_2150,In_1097,In_1764);
nand U2151 (N_2151,In_24,In_2255);
and U2152 (N_2152,In_603,In_2064);
and U2153 (N_2153,In_823,In_607);
nor U2154 (N_2154,In_1782,In_284);
nand U2155 (N_2155,In_2474,In_147);
or U2156 (N_2156,In_912,In_1268);
and U2157 (N_2157,In_1113,In_2072);
nor U2158 (N_2158,In_562,In_1839);
and U2159 (N_2159,In_1938,In_15);
or U2160 (N_2160,In_1623,In_1109);
nand U2161 (N_2161,In_673,In_1856);
and U2162 (N_2162,In_672,In_658);
nand U2163 (N_2163,In_1456,In_1453);
nand U2164 (N_2164,In_78,In_39);
and U2165 (N_2165,In_1768,In_2200);
nor U2166 (N_2166,In_815,In_65);
or U2167 (N_2167,In_1259,In_2030);
nand U2168 (N_2168,In_1308,In_1711);
and U2169 (N_2169,In_507,In_1676);
nand U2170 (N_2170,In_1963,In_744);
or U2171 (N_2171,In_1223,In_2411);
nor U2172 (N_2172,In_569,In_89);
or U2173 (N_2173,In_2057,In_2426);
nor U2174 (N_2174,In_2375,In_1939);
or U2175 (N_2175,In_1438,In_1118);
nand U2176 (N_2176,In_1495,In_714);
or U2177 (N_2177,In_952,In_1472);
or U2178 (N_2178,In_14,In_1157);
nand U2179 (N_2179,In_1291,In_869);
nor U2180 (N_2180,In_2252,In_454);
nand U2181 (N_2181,In_1697,In_1494);
or U2182 (N_2182,In_1639,In_729);
or U2183 (N_2183,In_308,In_1403);
nor U2184 (N_2184,In_2102,In_1323);
or U2185 (N_2185,In_979,In_85);
nor U2186 (N_2186,In_349,In_1799);
or U2187 (N_2187,In_625,In_2042);
nand U2188 (N_2188,In_765,In_965);
and U2189 (N_2189,In_1440,In_1590);
nand U2190 (N_2190,In_1049,In_140);
nand U2191 (N_2191,In_604,In_594);
nor U2192 (N_2192,In_2095,In_1994);
or U2193 (N_2193,In_1216,In_1480);
or U2194 (N_2194,In_1837,In_864);
nand U2195 (N_2195,In_1826,In_264);
nor U2196 (N_2196,In_396,In_2244);
nor U2197 (N_2197,In_1527,In_288);
nor U2198 (N_2198,In_593,In_1831);
and U2199 (N_2199,In_1578,In_1456);
and U2200 (N_2200,In_1539,In_312);
nor U2201 (N_2201,In_401,In_318);
and U2202 (N_2202,In_879,In_728);
nor U2203 (N_2203,In_768,In_1906);
xor U2204 (N_2204,In_2314,In_604);
nor U2205 (N_2205,In_137,In_1759);
nor U2206 (N_2206,In_2256,In_2085);
nand U2207 (N_2207,In_1797,In_486);
or U2208 (N_2208,In_618,In_2392);
or U2209 (N_2209,In_951,In_1454);
nor U2210 (N_2210,In_591,In_1776);
or U2211 (N_2211,In_236,In_1382);
and U2212 (N_2212,In_1240,In_876);
nand U2213 (N_2213,In_2370,In_246);
or U2214 (N_2214,In_1234,In_1686);
and U2215 (N_2215,In_329,In_2404);
or U2216 (N_2216,In_2061,In_1828);
and U2217 (N_2217,In_929,In_2447);
nand U2218 (N_2218,In_1959,In_2278);
and U2219 (N_2219,In_844,In_2475);
nor U2220 (N_2220,In_626,In_798);
nand U2221 (N_2221,In_2313,In_1830);
or U2222 (N_2222,In_2092,In_515);
and U2223 (N_2223,In_1415,In_1528);
or U2224 (N_2224,In_329,In_389);
nand U2225 (N_2225,In_2091,In_1681);
nand U2226 (N_2226,In_1037,In_1584);
or U2227 (N_2227,In_1063,In_1713);
or U2228 (N_2228,In_299,In_1680);
nand U2229 (N_2229,In_1353,In_305);
or U2230 (N_2230,In_2024,In_346);
nand U2231 (N_2231,In_2299,In_597);
nand U2232 (N_2232,In_1412,In_102);
and U2233 (N_2233,In_2310,In_100);
nor U2234 (N_2234,In_1588,In_986);
or U2235 (N_2235,In_2314,In_729);
nand U2236 (N_2236,In_1632,In_2217);
or U2237 (N_2237,In_2271,In_350);
nor U2238 (N_2238,In_2205,In_456);
and U2239 (N_2239,In_1867,In_1815);
nand U2240 (N_2240,In_668,In_2203);
and U2241 (N_2241,In_2077,In_1890);
and U2242 (N_2242,In_695,In_533);
nand U2243 (N_2243,In_1702,In_1782);
and U2244 (N_2244,In_2207,In_1012);
and U2245 (N_2245,In_1684,In_280);
and U2246 (N_2246,In_1916,In_1255);
nor U2247 (N_2247,In_2188,In_2024);
xnor U2248 (N_2248,In_412,In_2031);
and U2249 (N_2249,In_1293,In_668);
or U2250 (N_2250,In_1287,In_894);
nand U2251 (N_2251,In_141,In_1019);
nor U2252 (N_2252,In_2393,In_868);
nand U2253 (N_2253,In_1851,In_1091);
or U2254 (N_2254,In_2266,In_507);
and U2255 (N_2255,In_1319,In_1850);
nor U2256 (N_2256,In_1898,In_1865);
nor U2257 (N_2257,In_658,In_2429);
and U2258 (N_2258,In_1634,In_893);
nor U2259 (N_2259,In_2302,In_7);
nor U2260 (N_2260,In_1666,In_1183);
nor U2261 (N_2261,In_1570,In_2265);
or U2262 (N_2262,In_2168,In_823);
or U2263 (N_2263,In_2208,In_2072);
xnor U2264 (N_2264,In_1422,In_2118);
and U2265 (N_2265,In_1853,In_1318);
or U2266 (N_2266,In_2048,In_2289);
nor U2267 (N_2267,In_1623,In_1715);
or U2268 (N_2268,In_1341,In_1446);
xnor U2269 (N_2269,In_2086,In_57);
nor U2270 (N_2270,In_330,In_553);
or U2271 (N_2271,In_520,In_1591);
nand U2272 (N_2272,In_243,In_659);
and U2273 (N_2273,In_639,In_688);
nand U2274 (N_2274,In_210,In_1697);
xnor U2275 (N_2275,In_1798,In_835);
or U2276 (N_2276,In_813,In_756);
nand U2277 (N_2277,In_1026,In_1841);
and U2278 (N_2278,In_487,In_2412);
or U2279 (N_2279,In_1325,In_1208);
nand U2280 (N_2280,In_312,In_1750);
or U2281 (N_2281,In_1567,In_1891);
nor U2282 (N_2282,In_451,In_2261);
and U2283 (N_2283,In_2421,In_526);
and U2284 (N_2284,In_712,In_2304);
or U2285 (N_2285,In_1140,In_1428);
nand U2286 (N_2286,In_665,In_2323);
and U2287 (N_2287,In_404,In_2324);
or U2288 (N_2288,In_1245,In_926);
or U2289 (N_2289,In_789,In_424);
nand U2290 (N_2290,In_1083,In_2399);
and U2291 (N_2291,In_190,In_1448);
or U2292 (N_2292,In_2070,In_2288);
and U2293 (N_2293,In_748,In_1181);
nor U2294 (N_2294,In_36,In_1505);
or U2295 (N_2295,In_984,In_520);
or U2296 (N_2296,In_1423,In_672);
nand U2297 (N_2297,In_2290,In_758);
or U2298 (N_2298,In_54,In_1370);
or U2299 (N_2299,In_1088,In_618);
nand U2300 (N_2300,In_343,In_2071);
and U2301 (N_2301,In_2492,In_2052);
nor U2302 (N_2302,In_2428,In_1106);
or U2303 (N_2303,In_630,In_173);
or U2304 (N_2304,In_2083,In_1422);
nand U2305 (N_2305,In_136,In_156);
nor U2306 (N_2306,In_2000,In_1467);
nor U2307 (N_2307,In_544,In_1969);
nor U2308 (N_2308,In_269,In_337);
nor U2309 (N_2309,In_1091,In_1100);
nand U2310 (N_2310,In_901,In_2130);
nor U2311 (N_2311,In_2230,In_939);
nor U2312 (N_2312,In_2346,In_27);
or U2313 (N_2313,In_1434,In_533);
nand U2314 (N_2314,In_521,In_1623);
nand U2315 (N_2315,In_2414,In_280);
xnor U2316 (N_2316,In_2497,In_1352);
nand U2317 (N_2317,In_1372,In_1820);
nor U2318 (N_2318,In_623,In_2157);
nand U2319 (N_2319,In_1699,In_688);
and U2320 (N_2320,In_2202,In_1714);
and U2321 (N_2321,In_1379,In_1182);
nor U2322 (N_2322,In_1768,In_263);
nor U2323 (N_2323,In_788,In_864);
and U2324 (N_2324,In_2183,In_1705);
xnor U2325 (N_2325,In_357,In_395);
and U2326 (N_2326,In_649,In_1639);
and U2327 (N_2327,In_612,In_836);
or U2328 (N_2328,In_966,In_1441);
or U2329 (N_2329,In_2195,In_969);
and U2330 (N_2330,In_2067,In_928);
nand U2331 (N_2331,In_1095,In_1624);
nor U2332 (N_2332,In_1279,In_1292);
or U2333 (N_2333,In_1001,In_2243);
nand U2334 (N_2334,In_2108,In_508);
nor U2335 (N_2335,In_2067,In_396);
nand U2336 (N_2336,In_1856,In_1642);
nor U2337 (N_2337,In_1369,In_1352);
and U2338 (N_2338,In_178,In_1559);
nand U2339 (N_2339,In_1299,In_377);
nor U2340 (N_2340,In_1934,In_721);
and U2341 (N_2341,In_100,In_2448);
nand U2342 (N_2342,In_606,In_1539);
nor U2343 (N_2343,In_1282,In_718);
and U2344 (N_2344,In_1783,In_2225);
nor U2345 (N_2345,In_86,In_1927);
nand U2346 (N_2346,In_2019,In_2176);
nand U2347 (N_2347,In_1436,In_1985);
or U2348 (N_2348,In_1301,In_1907);
or U2349 (N_2349,In_1274,In_2249);
nand U2350 (N_2350,In_2069,In_427);
nor U2351 (N_2351,In_1040,In_419);
nor U2352 (N_2352,In_41,In_1335);
nor U2353 (N_2353,In_50,In_2097);
nand U2354 (N_2354,In_616,In_751);
nand U2355 (N_2355,In_650,In_325);
nor U2356 (N_2356,In_2175,In_1478);
nand U2357 (N_2357,In_614,In_1749);
nand U2358 (N_2358,In_2102,In_474);
or U2359 (N_2359,In_1944,In_443);
nand U2360 (N_2360,In_2036,In_896);
and U2361 (N_2361,In_1396,In_1156);
and U2362 (N_2362,In_2349,In_649);
or U2363 (N_2363,In_1901,In_1964);
xnor U2364 (N_2364,In_1862,In_612);
nand U2365 (N_2365,In_740,In_1780);
and U2366 (N_2366,In_304,In_1785);
xor U2367 (N_2367,In_1477,In_713);
nor U2368 (N_2368,In_2008,In_393);
and U2369 (N_2369,In_1578,In_2306);
nor U2370 (N_2370,In_1109,In_707);
or U2371 (N_2371,In_1132,In_255);
and U2372 (N_2372,In_510,In_2440);
or U2373 (N_2373,In_1471,In_121);
and U2374 (N_2374,In_1901,In_1395);
nand U2375 (N_2375,In_2216,In_1384);
or U2376 (N_2376,In_423,In_1008);
or U2377 (N_2377,In_128,In_503);
and U2378 (N_2378,In_1955,In_1723);
or U2379 (N_2379,In_1815,In_947);
nand U2380 (N_2380,In_1666,In_1435);
nor U2381 (N_2381,In_1032,In_2427);
nand U2382 (N_2382,In_76,In_1956);
nand U2383 (N_2383,In_217,In_1403);
or U2384 (N_2384,In_2345,In_1680);
nor U2385 (N_2385,In_1302,In_1271);
nor U2386 (N_2386,In_1262,In_25);
nor U2387 (N_2387,In_1410,In_930);
nand U2388 (N_2388,In_2418,In_136);
or U2389 (N_2389,In_2008,In_1905);
or U2390 (N_2390,In_129,In_968);
and U2391 (N_2391,In_8,In_404);
nand U2392 (N_2392,In_104,In_430);
and U2393 (N_2393,In_1051,In_2322);
nand U2394 (N_2394,In_121,In_86);
nand U2395 (N_2395,In_985,In_1016);
and U2396 (N_2396,In_293,In_901);
nor U2397 (N_2397,In_66,In_412);
nand U2398 (N_2398,In_929,In_629);
or U2399 (N_2399,In_994,In_2213);
nand U2400 (N_2400,In_1132,In_551);
xnor U2401 (N_2401,In_825,In_140);
nand U2402 (N_2402,In_817,In_307);
or U2403 (N_2403,In_1311,In_2210);
or U2404 (N_2404,In_1416,In_224);
nor U2405 (N_2405,In_2340,In_1617);
nor U2406 (N_2406,In_888,In_1459);
or U2407 (N_2407,In_798,In_136);
or U2408 (N_2408,In_207,In_1862);
nor U2409 (N_2409,In_2216,In_1998);
and U2410 (N_2410,In_2185,In_885);
nand U2411 (N_2411,In_248,In_1286);
nand U2412 (N_2412,In_477,In_53);
and U2413 (N_2413,In_423,In_880);
and U2414 (N_2414,In_27,In_1387);
xor U2415 (N_2415,In_526,In_532);
nand U2416 (N_2416,In_1064,In_1786);
and U2417 (N_2417,In_1217,In_1536);
nor U2418 (N_2418,In_1217,In_1401);
and U2419 (N_2419,In_1374,In_2252);
nor U2420 (N_2420,In_983,In_883);
nor U2421 (N_2421,In_266,In_1131);
or U2422 (N_2422,In_1412,In_1900);
or U2423 (N_2423,In_2333,In_1573);
and U2424 (N_2424,In_1514,In_1423);
and U2425 (N_2425,In_1014,In_48);
and U2426 (N_2426,In_1300,In_0);
nand U2427 (N_2427,In_2487,In_597);
or U2428 (N_2428,In_2359,In_1590);
nand U2429 (N_2429,In_762,In_1300);
or U2430 (N_2430,In_643,In_1892);
nand U2431 (N_2431,In_2024,In_1893);
nand U2432 (N_2432,In_1547,In_1618);
and U2433 (N_2433,In_697,In_278);
or U2434 (N_2434,In_399,In_1993);
or U2435 (N_2435,In_1105,In_2181);
and U2436 (N_2436,In_2374,In_894);
nand U2437 (N_2437,In_525,In_303);
or U2438 (N_2438,In_1247,In_1547);
and U2439 (N_2439,In_1866,In_2358);
and U2440 (N_2440,In_1362,In_1197);
and U2441 (N_2441,In_402,In_2416);
nor U2442 (N_2442,In_1213,In_250);
nand U2443 (N_2443,In_1965,In_507);
or U2444 (N_2444,In_861,In_721);
nor U2445 (N_2445,In_1951,In_2094);
and U2446 (N_2446,In_1313,In_1138);
or U2447 (N_2447,In_1664,In_425);
or U2448 (N_2448,In_351,In_1444);
nor U2449 (N_2449,In_51,In_2476);
nor U2450 (N_2450,In_2091,In_770);
nor U2451 (N_2451,In_1968,In_798);
or U2452 (N_2452,In_2302,In_345);
nor U2453 (N_2453,In_697,In_2281);
nand U2454 (N_2454,In_1261,In_1920);
or U2455 (N_2455,In_347,In_1385);
nor U2456 (N_2456,In_619,In_1618);
nor U2457 (N_2457,In_726,In_206);
nand U2458 (N_2458,In_688,In_359);
and U2459 (N_2459,In_194,In_1809);
nor U2460 (N_2460,In_1286,In_764);
and U2461 (N_2461,In_302,In_463);
nand U2462 (N_2462,In_1149,In_2171);
nor U2463 (N_2463,In_1954,In_1751);
and U2464 (N_2464,In_1289,In_1058);
nand U2465 (N_2465,In_1831,In_1310);
and U2466 (N_2466,In_1851,In_1159);
nor U2467 (N_2467,In_524,In_520);
nand U2468 (N_2468,In_1056,In_2193);
nand U2469 (N_2469,In_881,In_849);
or U2470 (N_2470,In_122,In_941);
nor U2471 (N_2471,In_181,In_440);
and U2472 (N_2472,In_1677,In_1028);
or U2473 (N_2473,In_1817,In_907);
nor U2474 (N_2474,In_1141,In_1331);
xnor U2475 (N_2475,In_951,In_837);
or U2476 (N_2476,In_258,In_573);
nand U2477 (N_2477,In_886,In_1881);
nor U2478 (N_2478,In_1428,In_1080);
nor U2479 (N_2479,In_559,In_1938);
nor U2480 (N_2480,In_2196,In_481);
nand U2481 (N_2481,In_1869,In_159);
and U2482 (N_2482,In_1136,In_1781);
nor U2483 (N_2483,In_121,In_1049);
or U2484 (N_2484,In_1893,In_762);
and U2485 (N_2485,In_1367,In_404);
and U2486 (N_2486,In_375,In_1351);
and U2487 (N_2487,In_2182,In_2063);
and U2488 (N_2488,In_128,In_1017);
and U2489 (N_2489,In_2201,In_1035);
nand U2490 (N_2490,In_19,In_737);
nor U2491 (N_2491,In_1954,In_2473);
nand U2492 (N_2492,In_381,In_415);
or U2493 (N_2493,In_1768,In_1231);
xor U2494 (N_2494,In_840,In_2191);
nor U2495 (N_2495,In_851,In_372);
nand U2496 (N_2496,In_594,In_1416);
or U2497 (N_2497,In_1288,In_1977);
nor U2498 (N_2498,In_601,In_425);
and U2499 (N_2499,In_1126,In_438);
and U2500 (N_2500,In_1195,In_1156);
or U2501 (N_2501,In_1662,In_2317);
xnor U2502 (N_2502,In_837,In_849);
and U2503 (N_2503,In_920,In_2404);
nor U2504 (N_2504,In_178,In_475);
nand U2505 (N_2505,In_769,In_252);
nor U2506 (N_2506,In_1192,In_116);
and U2507 (N_2507,In_1274,In_1024);
and U2508 (N_2508,In_618,In_99);
or U2509 (N_2509,In_1823,In_1149);
and U2510 (N_2510,In_223,In_2331);
or U2511 (N_2511,In_2160,In_1825);
and U2512 (N_2512,In_374,In_183);
nand U2513 (N_2513,In_1235,In_2412);
nor U2514 (N_2514,In_421,In_1742);
nor U2515 (N_2515,In_1164,In_2273);
nand U2516 (N_2516,In_2362,In_1515);
or U2517 (N_2517,In_1244,In_1769);
or U2518 (N_2518,In_1319,In_2015);
and U2519 (N_2519,In_646,In_1224);
nor U2520 (N_2520,In_362,In_2293);
nand U2521 (N_2521,In_186,In_1143);
and U2522 (N_2522,In_272,In_441);
nand U2523 (N_2523,In_2433,In_2117);
nand U2524 (N_2524,In_295,In_1592);
nor U2525 (N_2525,In_1829,In_556);
and U2526 (N_2526,In_2107,In_1676);
nor U2527 (N_2527,In_2356,In_1065);
or U2528 (N_2528,In_1893,In_2155);
or U2529 (N_2529,In_605,In_596);
nor U2530 (N_2530,In_974,In_464);
and U2531 (N_2531,In_1310,In_2007);
and U2532 (N_2532,In_1987,In_264);
and U2533 (N_2533,In_2042,In_24);
nor U2534 (N_2534,In_668,In_839);
nand U2535 (N_2535,In_93,In_690);
nand U2536 (N_2536,In_1660,In_2024);
nor U2537 (N_2537,In_648,In_2445);
nand U2538 (N_2538,In_83,In_342);
nand U2539 (N_2539,In_829,In_1654);
and U2540 (N_2540,In_413,In_1248);
nor U2541 (N_2541,In_1949,In_1776);
and U2542 (N_2542,In_473,In_2205);
and U2543 (N_2543,In_2021,In_2207);
nand U2544 (N_2544,In_1309,In_562);
and U2545 (N_2545,In_52,In_91);
and U2546 (N_2546,In_534,In_1499);
and U2547 (N_2547,In_1356,In_672);
and U2548 (N_2548,In_1435,In_2031);
and U2549 (N_2549,In_194,In_2263);
nand U2550 (N_2550,In_2404,In_2456);
or U2551 (N_2551,In_1884,In_2397);
or U2552 (N_2552,In_638,In_651);
or U2553 (N_2553,In_2226,In_1944);
nor U2554 (N_2554,In_2285,In_274);
and U2555 (N_2555,In_988,In_1379);
nor U2556 (N_2556,In_1622,In_2413);
and U2557 (N_2557,In_812,In_2277);
nand U2558 (N_2558,In_742,In_146);
and U2559 (N_2559,In_1505,In_185);
or U2560 (N_2560,In_2004,In_2418);
or U2561 (N_2561,In_2364,In_2104);
nand U2562 (N_2562,In_2126,In_2080);
or U2563 (N_2563,In_609,In_1694);
or U2564 (N_2564,In_1456,In_11);
nor U2565 (N_2565,In_2127,In_1949);
or U2566 (N_2566,In_1155,In_2491);
nor U2567 (N_2567,In_624,In_2267);
and U2568 (N_2568,In_445,In_504);
nor U2569 (N_2569,In_52,In_2195);
and U2570 (N_2570,In_753,In_2259);
nand U2571 (N_2571,In_2308,In_2485);
xnor U2572 (N_2572,In_936,In_2361);
nand U2573 (N_2573,In_1252,In_1756);
or U2574 (N_2574,In_1554,In_449);
and U2575 (N_2575,In_623,In_687);
or U2576 (N_2576,In_2099,In_345);
or U2577 (N_2577,In_688,In_112);
nor U2578 (N_2578,In_2422,In_692);
xor U2579 (N_2579,In_1617,In_171);
and U2580 (N_2580,In_1068,In_602);
nor U2581 (N_2581,In_223,In_2158);
nand U2582 (N_2582,In_1051,In_512);
or U2583 (N_2583,In_569,In_2285);
and U2584 (N_2584,In_1694,In_2299);
nor U2585 (N_2585,In_1130,In_513);
or U2586 (N_2586,In_1498,In_438);
or U2587 (N_2587,In_2156,In_1892);
nand U2588 (N_2588,In_2125,In_2213);
nand U2589 (N_2589,In_2416,In_1866);
and U2590 (N_2590,In_982,In_1146);
nand U2591 (N_2591,In_1669,In_194);
nand U2592 (N_2592,In_1059,In_301);
and U2593 (N_2593,In_1895,In_2319);
and U2594 (N_2594,In_2006,In_1758);
nand U2595 (N_2595,In_1498,In_1948);
or U2596 (N_2596,In_926,In_835);
nand U2597 (N_2597,In_1503,In_1286);
and U2598 (N_2598,In_684,In_2371);
nor U2599 (N_2599,In_2291,In_941);
nor U2600 (N_2600,In_593,In_1756);
nor U2601 (N_2601,In_21,In_2019);
nor U2602 (N_2602,In_1377,In_754);
nor U2603 (N_2603,In_398,In_907);
nand U2604 (N_2604,In_401,In_1096);
and U2605 (N_2605,In_2457,In_1919);
nand U2606 (N_2606,In_1925,In_1368);
or U2607 (N_2607,In_2287,In_888);
nor U2608 (N_2608,In_2158,In_2335);
nand U2609 (N_2609,In_2387,In_330);
and U2610 (N_2610,In_126,In_738);
nand U2611 (N_2611,In_2223,In_2215);
nor U2612 (N_2612,In_1936,In_299);
and U2613 (N_2613,In_214,In_2161);
and U2614 (N_2614,In_638,In_1191);
and U2615 (N_2615,In_1967,In_1432);
nand U2616 (N_2616,In_589,In_1496);
or U2617 (N_2617,In_574,In_1714);
or U2618 (N_2618,In_1719,In_264);
nand U2619 (N_2619,In_97,In_1579);
nor U2620 (N_2620,In_936,In_2246);
or U2621 (N_2621,In_111,In_899);
or U2622 (N_2622,In_848,In_878);
and U2623 (N_2623,In_359,In_443);
nor U2624 (N_2624,In_1715,In_1446);
nand U2625 (N_2625,In_34,In_73);
nor U2626 (N_2626,In_2325,In_1593);
nor U2627 (N_2627,In_1093,In_855);
nand U2628 (N_2628,In_683,In_2279);
nor U2629 (N_2629,In_433,In_1256);
nor U2630 (N_2630,In_515,In_583);
nor U2631 (N_2631,In_1312,In_648);
nand U2632 (N_2632,In_26,In_1721);
nand U2633 (N_2633,In_11,In_2376);
and U2634 (N_2634,In_109,In_2101);
or U2635 (N_2635,In_1790,In_1056);
and U2636 (N_2636,In_248,In_913);
nand U2637 (N_2637,In_1515,In_1078);
nand U2638 (N_2638,In_1805,In_851);
nand U2639 (N_2639,In_1973,In_1070);
nor U2640 (N_2640,In_121,In_1825);
nor U2641 (N_2641,In_567,In_2076);
and U2642 (N_2642,In_690,In_1872);
nor U2643 (N_2643,In_1200,In_1861);
or U2644 (N_2644,In_110,In_2414);
nor U2645 (N_2645,In_1408,In_1793);
nor U2646 (N_2646,In_2089,In_1046);
or U2647 (N_2647,In_316,In_2149);
and U2648 (N_2648,In_1951,In_2398);
and U2649 (N_2649,In_177,In_1335);
nor U2650 (N_2650,In_567,In_1892);
and U2651 (N_2651,In_154,In_898);
and U2652 (N_2652,In_1382,In_1283);
and U2653 (N_2653,In_1757,In_64);
and U2654 (N_2654,In_2336,In_258);
or U2655 (N_2655,In_371,In_695);
and U2656 (N_2656,In_1907,In_2084);
nor U2657 (N_2657,In_2291,In_1267);
nand U2658 (N_2658,In_1935,In_1363);
and U2659 (N_2659,In_975,In_1831);
and U2660 (N_2660,In_856,In_1028);
nor U2661 (N_2661,In_1099,In_1203);
and U2662 (N_2662,In_178,In_391);
and U2663 (N_2663,In_1975,In_407);
or U2664 (N_2664,In_1054,In_775);
nor U2665 (N_2665,In_1670,In_1872);
and U2666 (N_2666,In_994,In_802);
nor U2667 (N_2667,In_705,In_2065);
nand U2668 (N_2668,In_2246,In_1662);
nor U2669 (N_2669,In_80,In_996);
nor U2670 (N_2670,In_2243,In_2256);
xor U2671 (N_2671,In_921,In_971);
nand U2672 (N_2672,In_1484,In_1094);
nand U2673 (N_2673,In_873,In_1375);
nand U2674 (N_2674,In_801,In_1437);
and U2675 (N_2675,In_953,In_1186);
and U2676 (N_2676,In_2446,In_1149);
or U2677 (N_2677,In_1166,In_169);
and U2678 (N_2678,In_2474,In_490);
and U2679 (N_2679,In_618,In_672);
or U2680 (N_2680,In_744,In_1394);
and U2681 (N_2681,In_2194,In_1745);
nand U2682 (N_2682,In_2390,In_1918);
or U2683 (N_2683,In_928,In_1258);
nor U2684 (N_2684,In_693,In_741);
nand U2685 (N_2685,In_2148,In_1272);
and U2686 (N_2686,In_1601,In_165);
nand U2687 (N_2687,In_1709,In_2065);
nand U2688 (N_2688,In_497,In_854);
or U2689 (N_2689,In_878,In_1668);
and U2690 (N_2690,In_743,In_236);
or U2691 (N_2691,In_641,In_933);
or U2692 (N_2692,In_1791,In_64);
nor U2693 (N_2693,In_238,In_336);
and U2694 (N_2694,In_1287,In_637);
nor U2695 (N_2695,In_429,In_1180);
nand U2696 (N_2696,In_883,In_1773);
nor U2697 (N_2697,In_2035,In_2290);
nor U2698 (N_2698,In_1458,In_1431);
or U2699 (N_2699,In_961,In_1056);
nor U2700 (N_2700,In_342,In_1859);
or U2701 (N_2701,In_853,In_2054);
nor U2702 (N_2702,In_622,In_57);
xnor U2703 (N_2703,In_294,In_1713);
nand U2704 (N_2704,In_1493,In_1377);
or U2705 (N_2705,In_1585,In_31);
and U2706 (N_2706,In_569,In_1510);
xnor U2707 (N_2707,In_1907,In_1036);
and U2708 (N_2708,In_241,In_979);
nor U2709 (N_2709,In_1611,In_367);
nand U2710 (N_2710,In_1836,In_2465);
and U2711 (N_2711,In_1108,In_2195);
or U2712 (N_2712,In_1873,In_2305);
nor U2713 (N_2713,In_1857,In_1813);
nand U2714 (N_2714,In_490,In_1551);
and U2715 (N_2715,In_678,In_1297);
nor U2716 (N_2716,In_1413,In_2011);
or U2717 (N_2717,In_371,In_4);
and U2718 (N_2718,In_1716,In_1552);
and U2719 (N_2719,In_2424,In_1247);
nand U2720 (N_2720,In_1638,In_1247);
and U2721 (N_2721,In_778,In_2110);
nand U2722 (N_2722,In_621,In_987);
nand U2723 (N_2723,In_1009,In_93);
and U2724 (N_2724,In_1770,In_1876);
and U2725 (N_2725,In_1756,In_1871);
xnor U2726 (N_2726,In_457,In_1443);
nand U2727 (N_2727,In_470,In_512);
nor U2728 (N_2728,In_1847,In_2032);
and U2729 (N_2729,In_563,In_455);
and U2730 (N_2730,In_935,In_2366);
nand U2731 (N_2731,In_2440,In_1159);
or U2732 (N_2732,In_2024,In_1771);
or U2733 (N_2733,In_337,In_178);
and U2734 (N_2734,In_189,In_1485);
and U2735 (N_2735,In_736,In_1456);
or U2736 (N_2736,In_931,In_2125);
nand U2737 (N_2737,In_2298,In_335);
nand U2738 (N_2738,In_825,In_1593);
nand U2739 (N_2739,In_2206,In_790);
nand U2740 (N_2740,In_1483,In_2187);
and U2741 (N_2741,In_928,In_1152);
or U2742 (N_2742,In_1644,In_210);
or U2743 (N_2743,In_2254,In_2130);
nand U2744 (N_2744,In_1532,In_1579);
and U2745 (N_2745,In_2388,In_1727);
nand U2746 (N_2746,In_2345,In_1410);
nand U2747 (N_2747,In_772,In_1162);
and U2748 (N_2748,In_2169,In_1245);
nand U2749 (N_2749,In_55,In_2148);
or U2750 (N_2750,In_2100,In_1248);
xor U2751 (N_2751,In_1198,In_1460);
nor U2752 (N_2752,In_430,In_532);
nor U2753 (N_2753,In_223,In_2087);
nand U2754 (N_2754,In_1178,In_2166);
nand U2755 (N_2755,In_1595,In_483);
xor U2756 (N_2756,In_1589,In_2074);
xnor U2757 (N_2757,In_1407,In_608);
nor U2758 (N_2758,In_1457,In_226);
nor U2759 (N_2759,In_2244,In_325);
or U2760 (N_2760,In_520,In_481);
nand U2761 (N_2761,In_1395,In_1943);
or U2762 (N_2762,In_1863,In_609);
nor U2763 (N_2763,In_1178,In_583);
nand U2764 (N_2764,In_2496,In_1914);
nand U2765 (N_2765,In_724,In_2154);
and U2766 (N_2766,In_498,In_760);
or U2767 (N_2767,In_1096,In_2036);
and U2768 (N_2768,In_2259,In_527);
nand U2769 (N_2769,In_31,In_1554);
or U2770 (N_2770,In_510,In_1786);
and U2771 (N_2771,In_1950,In_770);
and U2772 (N_2772,In_1426,In_1620);
nor U2773 (N_2773,In_1155,In_1163);
or U2774 (N_2774,In_38,In_1428);
or U2775 (N_2775,In_2083,In_2005);
and U2776 (N_2776,In_1859,In_1172);
nor U2777 (N_2777,In_2179,In_1043);
xor U2778 (N_2778,In_2151,In_456);
or U2779 (N_2779,In_825,In_885);
nor U2780 (N_2780,In_2036,In_664);
or U2781 (N_2781,In_2051,In_376);
or U2782 (N_2782,In_1943,In_2253);
and U2783 (N_2783,In_179,In_123);
nand U2784 (N_2784,In_1356,In_1810);
nand U2785 (N_2785,In_166,In_814);
and U2786 (N_2786,In_1409,In_791);
nor U2787 (N_2787,In_515,In_1747);
or U2788 (N_2788,In_1744,In_288);
xnor U2789 (N_2789,In_385,In_2331);
or U2790 (N_2790,In_252,In_1619);
nor U2791 (N_2791,In_626,In_989);
or U2792 (N_2792,In_1049,In_390);
nor U2793 (N_2793,In_336,In_1230);
nor U2794 (N_2794,In_2480,In_823);
nor U2795 (N_2795,In_914,In_2222);
nor U2796 (N_2796,In_2122,In_1920);
or U2797 (N_2797,In_1742,In_1158);
or U2798 (N_2798,In_82,In_1245);
and U2799 (N_2799,In_2249,In_2112);
xor U2800 (N_2800,In_845,In_1089);
or U2801 (N_2801,In_66,In_2041);
nor U2802 (N_2802,In_1621,In_1003);
and U2803 (N_2803,In_582,In_1508);
or U2804 (N_2804,In_197,In_1903);
xnor U2805 (N_2805,In_98,In_1566);
nand U2806 (N_2806,In_1615,In_1271);
and U2807 (N_2807,In_2498,In_2049);
nor U2808 (N_2808,In_325,In_41);
and U2809 (N_2809,In_2086,In_826);
and U2810 (N_2810,In_1753,In_2224);
nand U2811 (N_2811,In_415,In_549);
nand U2812 (N_2812,In_1849,In_217);
nand U2813 (N_2813,In_1558,In_631);
and U2814 (N_2814,In_1373,In_1380);
nor U2815 (N_2815,In_2459,In_735);
nor U2816 (N_2816,In_2109,In_1444);
nor U2817 (N_2817,In_1268,In_459);
or U2818 (N_2818,In_1684,In_995);
or U2819 (N_2819,In_1370,In_1801);
and U2820 (N_2820,In_1429,In_2120);
or U2821 (N_2821,In_222,In_368);
nand U2822 (N_2822,In_2063,In_565);
nor U2823 (N_2823,In_371,In_938);
or U2824 (N_2824,In_1486,In_2179);
nor U2825 (N_2825,In_84,In_2397);
nor U2826 (N_2826,In_1372,In_665);
nand U2827 (N_2827,In_626,In_2132);
and U2828 (N_2828,In_273,In_2043);
nand U2829 (N_2829,In_743,In_1406);
nand U2830 (N_2830,In_2107,In_1723);
nor U2831 (N_2831,In_916,In_1402);
and U2832 (N_2832,In_1802,In_1670);
or U2833 (N_2833,In_2057,In_803);
or U2834 (N_2834,In_1148,In_2185);
or U2835 (N_2835,In_552,In_1073);
or U2836 (N_2836,In_1489,In_1353);
nor U2837 (N_2837,In_754,In_2360);
or U2838 (N_2838,In_484,In_1387);
nand U2839 (N_2839,In_732,In_538);
nor U2840 (N_2840,In_1769,In_1979);
nor U2841 (N_2841,In_412,In_2101);
nor U2842 (N_2842,In_552,In_1416);
nor U2843 (N_2843,In_367,In_1612);
nand U2844 (N_2844,In_1630,In_385);
or U2845 (N_2845,In_1660,In_452);
nor U2846 (N_2846,In_1943,In_1747);
nor U2847 (N_2847,In_2107,In_1468);
nor U2848 (N_2848,In_2134,In_1730);
or U2849 (N_2849,In_1282,In_2062);
nor U2850 (N_2850,In_414,In_1177);
or U2851 (N_2851,In_1240,In_910);
or U2852 (N_2852,In_1538,In_354);
and U2853 (N_2853,In_444,In_1496);
nor U2854 (N_2854,In_1265,In_822);
or U2855 (N_2855,In_713,In_1410);
nand U2856 (N_2856,In_2163,In_1517);
and U2857 (N_2857,In_524,In_937);
and U2858 (N_2858,In_1229,In_1506);
nor U2859 (N_2859,In_1990,In_2363);
or U2860 (N_2860,In_2413,In_292);
or U2861 (N_2861,In_1260,In_1613);
nand U2862 (N_2862,In_394,In_1784);
nand U2863 (N_2863,In_2028,In_293);
or U2864 (N_2864,In_1323,In_748);
nand U2865 (N_2865,In_1715,In_303);
or U2866 (N_2866,In_2456,In_10);
nor U2867 (N_2867,In_58,In_1096);
or U2868 (N_2868,In_988,In_2148);
xnor U2869 (N_2869,In_692,In_550);
nand U2870 (N_2870,In_1881,In_753);
nor U2871 (N_2871,In_120,In_1833);
or U2872 (N_2872,In_1082,In_825);
nand U2873 (N_2873,In_1816,In_1135);
and U2874 (N_2874,In_443,In_29);
nor U2875 (N_2875,In_399,In_2310);
nand U2876 (N_2876,In_1601,In_2400);
or U2877 (N_2877,In_1338,In_91);
and U2878 (N_2878,In_579,In_844);
or U2879 (N_2879,In_98,In_1218);
xor U2880 (N_2880,In_1753,In_2025);
or U2881 (N_2881,In_2188,In_265);
and U2882 (N_2882,In_1032,In_1611);
nand U2883 (N_2883,In_725,In_884);
nand U2884 (N_2884,In_1264,In_1469);
and U2885 (N_2885,In_741,In_1204);
or U2886 (N_2886,In_1896,In_407);
and U2887 (N_2887,In_1429,In_673);
nor U2888 (N_2888,In_833,In_1265);
nand U2889 (N_2889,In_1254,In_276);
and U2890 (N_2890,In_569,In_1856);
nor U2891 (N_2891,In_1463,In_1304);
and U2892 (N_2892,In_919,In_1376);
nor U2893 (N_2893,In_1087,In_2299);
or U2894 (N_2894,In_2486,In_1387);
nand U2895 (N_2895,In_2457,In_2302);
or U2896 (N_2896,In_1985,In_2081);
or U2897 (N_2897,In_8,In_49);
nand U2898 (N_2898,In_963,In_71);
nand U2899 (N_2899,In_136,In_1759);
nand U2900 (N_2900,In_2359,In_640);
nand U2901 (N_2901,In_2177,In_1142);
and U2902 (N_2902,In_529,In_2018);
or U2903 (N_2903,In_2241,In_1580);
nor U2904 (N_2904,In_728,In_1391);
xor U2905 (N_2905,In_1129,In_2414);
and U2906 (N_2906,In_2431,In_1236);
and U2907 (N_2907,In_530,In_1376);
or U2908 (N_2908,In_1531,In_2441);
or U2909 (N_2909,In_1150,In_618);
nand U2910 (N_2910,In_309,In_1322);
and U2911 (N_2911,In_1150,In_219);
or U2912 (N_2912,In_685,In_2153);
nor U2913 (N_2913,In_1850,In_331);
and U2914 (N_2914,In_1877,In_1267);
nand U2915 (N_2915,In_726,In_2313);
nand U2916 (N_2916,In_1058,In_1532);
or U2917 (N_2917,In_19,In_451);
nor U2918 (N_2918,In_858,In_494);
and U2919 (N_2919,In_914,In_1971);
xor U2920 (N_2920,In_330,In_190);
nor U2921 (N_2921,In_1745,In_1493);
xnor U2922 (N_2922,In_927,In_196);
and U2923 (N_2923,In_2423,In_1652);
nand U2924 (N_2924,In_1438,In_2396);
and U2925 (N_2925,In_1840,In_1742);
nor U2926 (N_2926,In_1126,In_2434);
nand U2927 (N_2927,In_635,In_1125);
and U2928 (N_2928,In_1799,In_29);
and U2929 (N_2929,In_2063,In_627);
xnor U2930 (N_2930,In_539,In_1519);
xnor U2931 (N_2931,In_858,In_358);
or U2932 (N_2932,In_612,In_1721);
nor U2933 (N_2933,In_1068,In_1330);
xor U2934 (N_2934,In_1463,In_1668);
nand U2935 (N_2935,In_877,In_1911);
xnor U2936 (N_2936,In_901,In_2236);
nand U2937 (N_2937,In_1170,In_2138);
and U2938 (N_2938,In_1473,In_8);
or U2939 (N_2939,In_2253,In_594);
and U2940 (N_2940,In_2141,In_507);
or U2941 (N_2941,In_1581,In_931);
and U2942 (N_2942,In_2233,In_1130);
or U2943 (N_2943,In_1420,In_1536);
and U2944 (N_2944,In_1997,In_110);
nor U2945 (N_2945,In_1733,In_290);
nor U2946 (N_2946,In_1547,In_1456);
nand U2947 (N_2947,In_1565,In_1892);
nor U2948 (N_2948,In_863,In_1833);
or U2949 (N_2949,In_61,In_1769);
nand U2950 (N_2950,In_2443,In_1379);
nor U2951 (N_2951,In_1967,In_2281);
or U2952 (N_2952,In_1837,In_2339);
nor U2953 (N_2953,In_1219,In_1934);
nand U2954 (N_2954,In_1010,In_2036);
nor U2955 (N_2955,In_7,In_183);
nand U2956 (N_2956,In_568,In_865);
and U2957 (N_2957,In_1676,In_658);
nor U2958 (N_2958,In_1440,In_78);
nor U2959 (N_2959,In_1686,In_98);
or U2960 (N_2960,In_133,In_332);
or U2961 (N_2961,In_271,In_541);
or U2962 (N_2962,In_2274,In_1092);
or U2963 (N_2963,In_204,In_1387);
nand U2964 (N_2964,In_613,In_2249);
or U2965 (N_2965,In_619,In_1934);
nor U2966 (N_2966,In_2250,In_1291);
or U2967 (N_2967,In_775,In_1586);
nand U2968 (N_2968,In_1638,In_1695);
nor U2969 (N_2969,In_1579,In_1740);
nand U2970 (N_2970,In_590,In_796);
or U2971 (N_2971,In_463,In_487);
and U2972 (N_2972,In_1262,In_2113);
and U2973 (N_2973,In_831,In_2262);
and U2974 (N_2974,In_118,In_299);
nor U2975 (N_2975,In_1603,In_2351);
xnor U2976 (N_2976,In_2353,In_390);
nor U2977 (N_2977,In_172,In_1227);
nor U2978 (N_2978,In_2345,In_839);
nand U2979 (N_2979,In_1505,In_529);
and U2980 (N_2980,In_1599,In_1696);
nand U2981 (N_2981,In_2174,In_32);
or U2982 (N_2982,In_1974,In_1871);
and U2983 (N_2983,In_1454,In_1397);
nand U2984 (N_2984,In_1999,In_315);
nand U2985 (N_2985,In_814,In_363);
and U2986 (N_2986,In_587,In_855);
or U2987 (N_2987,In_1719,In_270);
xnor U2988 (N_2988,In_1460,In_425);
and U2989 (N_2989,In_1929,In_100);
nor U2990 (N_2990,In_2341,In_980);
or U2991 (N_2991,In_2093,In_1529);
and U2992 (N_2992,In_1396,In_639);
and U2993 (N_2993,In_2134,In_816);
nand U2994 (N_2994,In_1089,In_2196);
nor U2995 (N_2995,In_290,In_1638);
or U2996 (N_2996,In_814,In_1961);
nor U2997 (N_2997,In_1417,In_2253);
or U2998 (N_2998,In_2175,In_4);
and U2999 (N_2999,In_1237,In_1708);
nor U3000 (N_3000,In_522,In_1729);
or U3001 (N_3001,In_935,In_1771);
nand U3002 (N_3002,In_1784,In_2312);
nor U3003 (N_3003,In_1132,In_307);
or U3004 (N_3004,In_1606,In_1576);
nor U3005 (N_3005,In_823,In_549);
nand U3006 (N_3006,In_303,In_1319);
nor U3007 (N_3007,In_1198,In_595);
nand U3008 (N_3008,In_553,In_801);
nand U3009 (N_3009,In_1099,In_311);
and U3010 (N_3010,In_1238,In_2188);
nor U3011 (N_3011,In_1721,In_417);
and U3012 (N_3012,In_1169,In_402);
or U3013 (N_3013,In_989,In_498);
and U3014 (N_3014,In_1185,In_840);
nand U3015 (N_3015,In_1616,In_721);
and U3016 (N_3016,In_991,In_1948);
nand U3017 (N_3017,In_1016,In_1789);
nor U3018 (N_3018,In_1421,In_2327);
or U3019 (N_3019,In_2401,In_407);
nand U3020 (N_3020,In_1291,In_2246);
xnor U3021 (N_3021,In_762,In_1042);
or U3022 (N_3022,In_853,In_622);
nor U3023 (N_3023,In_815,In_86);
and U3024 (N_3024,In_394,In_1380);
nor U3025 (N_3025,In_1154,In_1313);
nor U3026 (N_3026,In_955,In_963);
nand U3027 (N_3027,In_1788,In_1021);
and U3028 (N_3028,In_126,In_1425);
or U3029 (N_3029,In_2090,In_686);
or U3030 (N_3030,In_478,In_2138);
or U3031 (N_3031,In_772,In_1583);
or U3032 (N_3032,In_2080,In_782);
nand U3033 (N_3033,In_1863,In_567);
nor U3034 (N_3034,In_1076,In_2322);
or U3035 (N_3035,In_1653,In_2006);
and U3036 (N_3036,In_1639,In_36);
or U3037 (N_3037,In_1368,In_1726);
or U3038 (N_3038,In_2148,In_1263);
nor U3039 (N_3039,In_375,In_1684);
nor U3040 (N_3040,In_2254,In_1189);
or U3041 (N_3041,In_1675,In_1648);
nand U3042 (N_3042,In_2237,In_1555);
or U3043 (N_3043,In_235,In_1256);
nor U3044 (N_3044,In_2307,In_1721);
or U3045 (N_3045,In_1332,In_923);
and U3046 (N_3046,In_80,In_1850);
and U3047 (N_3047,In_1758,In_379);
nand U3048 (N_3048,In_1185,In_51);
or U3049 (N_3049,In_204,In_1745);
and U3050 (N_3050,In_1432,In_388);
and U3051 (N_3051,In_413,In_1036);
and U3052 (N_3052,In_2388,In_1796);
or U3053 (N_3053,In_2258,In_88);
or U3054 (N_3054,In_392,In_677);
and U3055 (N_3055,In_1439,In_674);
xor U3056 (N_3056,In_999,In_845);
nor U3057 (N_3057,In_242,In_1959);
or U3058 (N_3058,In_104,In_538);
nand U3059 (N_3059,In_514,In_371);
nand U3060 (N_3060,In_2296,In_930);
nor U3061 (N_3061,In_818,In_2194);
or U3062 (N_3062,In_678,In_314);
and U3063 (N_3063,In_2237,In_452);
xor U3064 (N_3064,In_1880,In_628);
or U3065 (N_3065,In_2299,In_1839);
and U3066 (N_3066,In_1317,In_1580);
and U3067 (N_3067,In_563,In_2110);
nand U3068 (N_3068,In_1430,In_1573);
nand U3069 (N_3069,In_1126,In_1495);
nor U3070 (N_3070,In_835,In_2288);
nand U3071 (N_3071,In_186,In_599);
nor U3072 (N_3072,In_956,In_960);
xnor U3073 (N_3073,In_1956,In_792);
and U3074 (N_3074,In_206,In_734);
nand U3075 (N_3075,In_2100,In_1610);
nor U3076 (N_3076,In_2014,In_1512);
nor U3077 (N_3077,In_1869,In_762);
nand U3078 (N_3078,In_1996,In_1413);
nor U3079 (N_3079,In_184,In_1161);
nor U3080 (N_3080,In_649,In_2338);
and U3081 (N_3081,In_729,In_1179);
nand U3082 (N_3082,In_1839,In_2262);
or U3083 (N_3083,In_2130,In_2243);
and U3084 (N_3084,In_276,In_1663);
nand U3085 (N_3085,In_768,In_2113);
and U3086 (N_3086,In_1016,In_1511);
nor U3087 (N_3087,In_1475,In_508);
and U3088 (N_3088,In_913,In_2463);
and U3089 (N_3089,In_2049,In_2190);
nand U3090 (N_3090,In_191,In_1048);
and U3091 (N_3091,In_2256,In_772);
and U3092 (N_3092,In_1001,In_460);
nor U3093 (N_3093,In_1854,In_1563);
or U3094 (N_3094,In_1335,In_2045);
and U3095 (N_3095,In_1600,In_1750);
and U3096 (N_3096,In_2075,In_1160);
or U3097 (N_3097,In_956,In_678);
or U3098 (N_3098,In_50,In_2003);
and U3099 (N_3099,In_2032,In_461);
and U3100 (N_3100,In_2417,In_322);
or U3101 (N_3101,In_1356,In_1997);
and U3102 (N_3102,In_1123,In_1277);
and U3103 (N_3103,In_714,In_1152);
nand U3104 (N_3104,In_1530,In_1500);
or U3105 (N_3105,In_2313,In_680);
and U3106 (N_3106,In_854,In_1456);
nand U3107 (N_3107,In_1905,In_2183);
or U3108 (N_3108,In_1635,In_1294);
and U3109 (N_3109,In_1408,In_2070);
nor U3110 (N_3110,In_1199,In_973);
nand U3111 (N_3111,In_2155,In_435);
and U3112 (N_3112,In_953,In_389);
nand U3113 (N_3113,In_1988,In_2468);
nand U3114 (N_3114,In_1439,In_1825);
or U3115 (N_3115,In_526,In_416);
nand U3116 (N_3116,In_1958,In_1684);
nand U3117 (N_3117,In_2372,In_1443);
and U3118 (N_3118,In_595,In_279);
and U3119 (N_3119,In_436,In_312);
nand U3120 (N_3120,In_2274,In_876);
or U3121 (N_3121,In_187,In_1381);
nor U3122 (N_3122,In_1332,In_890);
or U3123 (N_3123,In_2021,In_1289);
and U3124 (N_3124,In_2102,In_922);
nor U3125 (N_3125,In_53,In_2224);
nand U3126 (N_3126,In_2336,In_746);
nand U3127 (N_3127,In_563,In_667);
nor U3128 (N_3128,In_1355,In_585);
and U3129 (N_3129,In_1512,In_481);
and U3130 (N_3130,In_663,In_2306);
or U3131 (N_3131,In_39,In_1428);
or U3132 (N_3132,In_1606,In_1326);
nor U3133 (N_3133,In_14,In_1941);
or U3134 (N_3134,In_1123,In_352);
nand U3135 (N_3135,In_1750,In_1562);
and U3136 (N_3136,In_887,In_2207);
and U3137 (N_3137,In_2145,In_1395);
nor U3138 (N_3138,In_2127,In_1575);
and U3139 (N_3139,In_1,In_852);
or U3140 (N_3140,In_688,In_1028);
or U3141 (N_3141,In_584,In_2064);
nand U3142 (N_3142,In_802,In_337);
nand U3143 (N_3143,In_504,In_1133);
or U3144 (N_3144,In_740,In_968);
and U3145 (N_3145,In_985,In_2278);
or U3146 (N_3146,In_374,In_229);
nor U3147 (N_3147,In_2351,In_871);
nand U3148 (N_3148,In_1350,In_770);
and U3149 (N_3149,In_2250,In_2405);
or U3150 (N_3150,In_1031,In_1673);
nand U3151 (N_3151,In_790,In_88);
or U3152 (N_3152,In_481,In_1256);
and U3153 (N_3153,In_1728,In_2326);
nand U3154 (N_3154,In_1237,In_1735);
or U3155 (N_3155,In_332,In_369);
nand U3156 (N_3156,In_302,In_2024);
or U3157 (N_3157,In_329,In_2114);
nor U3158 (N_3158,In_28,In_744);
nand U3159 (N_3159,In_1601,In_1634);
or U3160 (N_3160,In_505,In_646);
or U3161 (N_3161,In_317,In_837);
nor U3162 (N_3162,In_120,In_1756);
and U3163 (N_3163,In_150,In_1148);
nand U3164 (N_3164,In_1246,In_2053);
nand U3165 (N_3165,In_227,In_938);
or U3166 (N_3166,In_139,In_1530);
or U3167 (N_3167,In_258,In_2168);
or U3168 (N_3168,In_2031,In_1589);
or U3169 (N_3169,In_2131,In_2272);
nand U3170 (N_3170,In_2091,In_515);
or U3171 (N_3171,In_1421,In_796);
nand U3172 (N_3172,In_2023,In_196);
nor U3173 (N_3173,In_437,In_530);
or U3174 (N_3174,In_423,In_482);
nand U3175 (N_3175,In_2062,In_1060);
and U3176 (N_3176,In_501,In_385);
and U3177 (N_3177,In_2268,In_2241);
xor U3178 (N_3178,In_1122,In_826);
nand U3179 (N_3179,In_691,In_172);
or U3180 (N_3180,In_37,In_1451);
nand U3181 (N_3181,In_1223,In_9);
nor U3182 (N_3182,In_476,In_374);
or U3183 (N_3183,In_2363,In_1114);
nand U3184 (N_3184,In_274,In_1745);
nand U3185 (N_3185,In_968,In_71);
nand U3186 (N_3186,In_2028,In_2042);
nand U3187 (N_3187,In_847,In_616);
and U3188 (N_3188,In_1619,In_1957);
or U3189 (N_3189,In_1683,In_252);
nand U3190 (N_3190,In_493,In_1481);
nor U3191 (N_3191,In_1594,In_1053);
and U3192 (N_3192,In_1275,In_212);
nor U3193 (N_3193,In_2063,In_1632);
nor U3194 (N_3194,In_575,In_1563);
nand U3195 (N_3195,In_1559,In_2493);
xnor U3196 (N_3196,In_970,In_2002);
or U3197 (N_3197,In_311,In_1097);
and U3198 (N_3198,In_178,In_1281);
nand U3199 (N_3199,In_1998,In_1286);
nor U3200 (N_3200,In_1133,In_1631);
xnor U3201 (N_3201,In_1371,In_2353);
nor U3202 (N_3202,In_127,In_615);
and U3203 (N_3203,In_673,In_2370);
nand U3204 (N_3204,In_1658,In_486);
nor U3205 (N_3205,In_1258,In_2211);
or U3206 (N_3206,In_855,In_603);
nand U3207 (N_3207,In_2436,In_1240);
nand U3208 (N_3208,In_723,In_85);
nor U3209 (N_3209,In_866,In_647);
or U3210 (N_3210,In_1584,In_2153);
xnor U3211 (N_3211,In_199,In_1780);
nand U3212 (N_3212,In_1840,In_588);
nand U3213 (N_3213,In_756,In_520);
nand U3214 (N_3214,In_2433,In_1590);
and U3215 (N_3215,In_1905,In_705);
xor U3216 (N_3216,In_2449,In_932);
and U3217 (N_3217,In_1158,In_625);
and U3218 (N_3218,In_47,In_1155);
and U3219 (N_3219,In_1995,In_1309);
or U3220 (N_3220,In_2397,In_70);
nor U3221 (N_3221,In_1434,In_237);
nand U3222 (N_3222,In_324,In_988);
or U3223 (N_3223,In_730,In_461);
or U3224 (N_3224,In_1875,In_757);
nor U3225 (N_3225,In_80,In_1272);
or U3226 (N_3226,In_667,In_174);
nor U3227 (N_3227,In_472,In_170);
and U3228 (N_3228,In_1607,In_675);
nor U3229 (N_3229,In_1869,In_1549);
or U3230 (N_3230,In_1725,In_397);
and U3231 (N_3231,In_2300,In_198);
and U3232 (N_3232,In_877,In_1365);
or U3233 (N_3233,In_664,In_1252);
and U3234 (N_3234,In_1077,In_945);
nand U3235 (N_3235,In_1661,In_93);
xnor U3236 (N_3236,In_835,In_5);
or U3237 (N_3237,In_2236,In_841);
or U3238 (N_3238,In_1502,In_2291);
or U3239 (N_3239,In_2376,In_463);
or U3240 (N_3240,In_299,In_1505);
or U3241 (N_3241,In_1270,In_1307);
nor U3242 (N_3242,In_964,In_1593);
and U3243 (N_3243,In_131,In_732);
or U3244 (N_3244,In_581,In_189);
and U3245 (N_3245,In_2469,In_1678);
nand U3246 (N_3246,In_1161,In_1010);
nand U3247 (N_3247,In_2187,In_1728);
nand U3248 (N_3248,In_1354,In_799);
and U3249 (N_3249,In_2301,In_149);
xnor U3250 (N_3250,In_518,In_208);
nor U3251 (N_3251,In_623,In_1641);
and U3252 (N_3252,In_586,In_1598);
nor U3253 (N_3253,In_1895,In_230);
nand U3254 (N_3254,In_242,In_895);
or U3255 (N_3255,In_1564,In_1274);
or U3256 (N_3256,In_657,In_2354);
nor U3257 (N_3257,In_1432,In_650);
nand U3258 (N_3258,In_407,In_1164);
nor U3259 (N_3259,In_393,In_60);
and U3260 (N_3260,In_1769,In_23);
or U3261 (N_3261,In_392,In_557);
xor U3262 (N_3262,In_328,In_1209);
nand U3263 (N_3263,In_2321,In_368);
nand U3264 (N_3264,In_1922,In_644);
or U3265 (N_3265,In_2440,In_1628);
and U3266 (N_3266,In_1543,In_2425);
nor U3267 (N_3267,In_2211,In_1581);
and U3268 (N_3268,In_2414,In_8);
or U3269 (N_3269,In_1522,In_420);
nor U3270 (N_3270,In_321,In_990);
and U3271 (N_3271,In_1472,In_713);
nor U3272 (N_3272,In_1687,In_2462);
and U3273 (N_3273,In_1887,In_632);
nand U3274 (N_3274,In_1368,In_1435);
or U3275 (N_3275,In_2433,In_1171);
and U3276 (N_3276,In_1551,In_2278);
and U3277 (N_3277,In_172,In_2285);
nor U3278 (N_3278,In_1048,In_2216);
and U3279 (N_3279,In_979,In_1824);
and U3280 (N_3280,In_849,In_1629);
nand U3281 (N_3281,In_498,In_1266);
or U3282 (N_3282,In_853,In_166);
or U3283 (N_3283,In_1531,In_1530);
nand U3284 (N_3284,In_90,In_2446);
or U3285 (N_3285,In_1959,In_2288);
nor U3286 (N_3286,In_1681,In_2218);
and U3287 (N_3287,In_2384,In_826);
and U3288 (N_3288,In_1194,In_1608);
nor U3289 (N_3289,In_1111,In_411);
nor U3290 (N_3290,In_1262,In_35);
nor U3291 (N_3291,In_132,In_1298);
xor U3292 (N_3292,In_200,In_2068);
nand U3293 (N_3293,In_1296,In_1117);
and U3294 (N_3294,In_1813,In_1647);
nand U3295 (N_3295,In_204,In_442);
and U3296 (N_3296,In_1670,In_350);
nor U3297 (N_3297,In_1901,In_1822);
or U3298 (N_3298,In_570,In_14);
and U3299 (N_3299,In_1838,In_1813);
and U3300 (N_3300,In_1788,In_1102);
nand U3301 (N_3301,In_1942,In_1967);
or U3302 (N_3302,In_1742,In_701);
or U3303 (N_3303,In_70,In_817);
nand U3304 (N_3304,In_1852,In_99);
and U3305 (N_3305,In_93,In_103);
nand U3306 (N_3306,In_961,In_1675);
and U3307 (N_3307,In_1909,In_1113);
nor U3308 (N_3308,In_435,In_1651);
nand U3309 (N_3309,In_871,In_185);
nand U3310 (N_3310,In_427,In_363);
nor U3311 (N_3311,In_314,In_1721);
and U3312 (N_3312,In_32,In_1952);
and U3313 (N_3313,In_1177,In_1497);
or U3314 (N_3314,In_1911,In_1909);
and U3315 (N_3315,In_2198,In_1521);
nor U3316 (N_3316,In_1004,In_88);
and U3317 (N_3317,In_1894,In_894);
nor U3318 (N_3318,In_804,In_397);
or U3319 (N_3319,In_544,In_1918);
nand U3320 (N_3320,In_1958,In_527);
and U3321 (N_3321,In_2081,In_949);
nand U3322 (N_3322,In_2019,In_2272);
and U3323 (N_3323,In_411,In_156);
and U3324 (N_3324,In_954,In_914);
and U3325 (N_3325,In_2203,In_690);
nand U3326 (N_3326,In_1099,In_275);
or U3327 (N_3327,In_199,In_924);
nor U3328 (N_3328,In_1067,In_1139);
or U3329 (N_3329,In_1148,In_779);
nor U3330 (N_3330,In_458,In_475);
nor U3331 (N_3331,In_1622,In_498);
or U3332 (N_3332,In_2184,In_1870);
and U3333 (N_3333,In_285,In_383);
and U3334 (N_3334,In_745,In_246);
nor U3335 (N_3335,In_2404,In_991);
or U3336 (N_3336,In_1636,In_1508);
nand U3337 (N_3337,In_2062,In_2146);
nand U3338 (N_3338,In_211,In_1190);
nand U3339 (N_3339,In_2052,In_1022);
nor U3340 (N_3340,In_2080,In_2);
nand U3341 (N_3341,In_1726,In_2159);
and U3342 (N_3342,In_523,In_278);
nor U3343 (N_3343,In_125,In_1767);
xnor U3344 (N_3344,In_1269,In_683);
nand U3345 (N_3345,In_1249,In_2283);
or U3346 (N_3346,In_2275,In_448);
xor U3347 (N_3347,In_118,In_2127);
nand U3348 (N_3348,In_2174,In_1290);
and U3349 (N_3349,In_2027,In_1108);
nor U3350 (N_3350,In_2055,In_323);
and U3351 (N_3351,In_2155,In_384);
nand U3352 (N_3352,In_1227,In_112);
and U3353 (N_3353,In_721,In_2270);
and U3354 (N_3354,In_2294,In_307);
or U3355 (N_3355,In_2141,In_1290);
and U3356 (N_3356,In_2446,In_2350);
and U3357 (N_3357,In_1002,In_2055);
nand U3358 (N_3358,In_1386,In_1420);
and U3359 (N_3359,In_1041,In_2421);
or U3360 (N_3360,In_372,In_26);
or U3361 (N_3361,In_2062,In_430);
xnor U3362 (N_3362,In_1926,In_2072);
nor U3363 (N_3363,In_1465,In_507);
and U3364 (N_3364,In_32,In_967);
or U3365 (N_3365,In_1648,In_933);
nor U3366 (N_3366,In_1509,In_1808);
nand U3367 (N_3367,In_775,In_543);
or U3368 (N_3368,In_1728,In_704);
nor U3369 (N_3369,In_537,In_1151);
nor U3370 (N_3370,In_416,In_2122);
nand U3371 (N_3371,In_1624,In_2372);
and U3372 (N_3372,In_2270,In_2034);
or U3373 (N_3373,In_1852,In_2169);
nor U3374 (N_3374,In_1261,In_2395);
nand U3375 (N_3375,In_857,In_497);
nor U3376 (N_3376,In_827,In_1729);
or U3377 (N_3377,In_1625,In_1158);
or U3378 (N_3378,In_665,In_201);
xor U3379 (N_3379,In_1459,In_2480);
nand U3380 (N_3380,In_2036,In_784);
or U3381 (N_3381,In_1740,In_1033);
and U3382 (N_3382,In_1142,In_2498);
nor U3383 (N_3383,In_314,In_500);
nand U3384 (N_3384,In_1656,In_2297);
or U3385 (N_3385,In_847,In_1538);
and U3386 (N_3386,In_711,In_379);
or U3387 (N_3387,In_1863,In_2193);
and U3388 (N_3388,In_1354,In_1446);
and U3389 (N_3389,In_577,In_814);
nand U3390 (N_3390,In_2329,In_2145);
or U3391 (N_3391,In_910,In_340);
or U3392 (N_3392,In_1727,In_70);
or U3393 (N_3393,In_189,In_1167);
nand U3394 (N_3394,In_1478,In_1001);
and U3395 (N_3395,In_171,In_2351);
nand U3396 (N_3396,In_382,In_1423);
and U3397 (N_3397,In_277,In_623);
nand U3398 (N_3398,In_1469,In_2182);
nand U3399 (N_3399,In_1383,In_920);
nor U3400 (N_3400,In_1448,In_619);
nand U3401 (N_3401,In_1497,In_261);
nor U3402 (N_3402,In_1338,In_307);
and U3403 (N_3403,In_1802,In_2410);
nand U3404 (N_3404,In_979,In_1521);
and U3405 (N_3405,In_1253,In_571);
nor U3406 (N_3406,In_652,In_1408);
or U3407 (N_3407,In_1536,In_184);
or U3408 (N_3408,In_604,In_1047);
and U3409 (N_3409,In_849,In_1118);
and U3410 (N_3410,In_2151,In_1275);
and U3411 (N_3411,In_839,In_2150);
nand U3412 (N_3412,In_386,In_920);
and U3413 (N_3413,In_88,In_1007);
or U3414 (N_3414,In_93,In_1621);
xor U3415 (N_3415,In_558,In_2216);
or U3416 (N_3416,In_1229,In_520);
or U3417 (N_3417,In_541,In_1947);
or U3418 (N_3418,In_2273,In_1265);
and U3419 (N_3419,In_2116,In_2283);
nand U3420 (N_3420,In_665,In_757);
and U3421 (N_3421,In_1735,In_257);
nor U3422 (N_3422,In_2133,In_853);
nand U3423 (N_3423,In_1572,In_1202);
or U3424 (N_3424,In_1974,In_1000);
and U3425 (N_3425,In_43,In_2325);
xor U3426 (N_3426,In_1970,In_1100);
nor U3427 (N_3427,In_2054,In_861);
and U3428 (N_3428,In_2266,In_2099);
nor U3429 (N_3429,In_2279,In_1688);
nand U3430 (N_3430,In_1522,In_1750);
or U3431 (N_3431,In_1091,In_1434);
or U3432 (N_3432,In_582,In_1765);
or U3433 (N_3433,In_856,In_2128);
and U3434 (N_3434,In_1735,In_739);
or U3435 (N_3435,In_101,In_632);
nor U3436 (N_3436,In_460,In_775);
and U3437 (N_3437,In_1619,In_1652);
and U3438 (N_3438,In_2160,In_50);
nand U3439 (N_3439,In_2421,In_2127);
and U3440 (N_3440,In_935,In_1093);
or U3441 (N_3441,In_1635,In_2319);
nor U3442 (N_3442,In_410,In_999);
nor U3443 (N_3443,In_2232,In_969);
nand U3444 (N_3444,In_813,In_1305);
nand U3445 (N_3445,In_2371,In_844);
and U3446 (N_3446,In_423,In_1636);
nand U3447 (N_3447,In_1825,In_1375);
or U3448 (N_3448,In_397,In_244);
nor U3449 (N_3449,In_637,In_2337);
nand U3450 (N_3450,In_1633,In_2336);
nand U3451 (N_3451,In_997,In_371);
and U3452 (N_3452,In_459,In_967);
nand U3453 (N_3453,In_982,In_1236);
and U3454 (N_3454,In_449,In_2008);
nor U3455 (N_3455,In_1116,In_414);
nor U3456 (N_3456,In_840,In_1397);
nor U3457 (N_3457,In_1207,In_1227);
and U3458 (N_3458,In_691,In_855);
nor U3459 (N_3459,In_392,In_902);
nand U3460 (N_3460,In_1981,In_1692);
and U3461 (N_3461,In_518,In_1941);
nor U3462 (N_3462,In_2311,In_1762);
nor U3463 (N_3463,In_1274,In_850);
or U3464 (N_3464,In_1564,In_1977);
nor U3465 (N_3465,In_858,In_2434);
nand U3466 (N_3466,In_2122,In_1534);
or U3467 (N_3467,In_872,In_2320);
nand U3468 (N_3468,In_2422,In_1320);
or U3469 (N_3469,In_889,In_233);
nor U3470 (N_3470,In_2157,In_119);
nor U3471 (N_3471,In_1842,In_1364);
nor U3472 (N_3472,In_629,In_1455);
nor U3473 (N_3473,In_766,In_1154);
or U3474 (N_3474,In_1132,In_2081);
and U3475 (N_3475,In_1741,In_1843);
or U3476 (N_3476,In_908,In_639);
or U3477 (N_3477,In_317,In_108);
or U3478 (N_3478,In_34,In_1098);
and U3479 (N_3479,In_131,In_2024);
and U3480 (N_3480,In_411,In_390);
or U3481 (N_3481,In_683,In_1556);
or U3482 (N_3482,In_2076,In_1552);
and U3483 (N_3483,In_1219,In_23);
nor U3484 (N_3484,In_658,In_2086);
or U3485 (N_3485,In_2390,In_1818);
and U3486 (N_3486,In_2410,In_309);
nand U3487 (N_3487,In_1397,In_1420);
nand U3488 (N_3488,In_2155,In_2001);
nor U3489 (N_3489,In_2168,In_2384);
xor U3490 (N_3490,In_902,In_140);
or U3491 (N_3491,In_176,In_860);
or U3492 (N_3492,In_729,In_1286);
and U3493 (N_3493,In_2180,In_1736);
nor U3494 (N_3494,In_227,In_995);
or U3495 (N_3495,In_2444,In_1338);
xnor U3496 (N_3496,In_2494,In_431);
nor U3497 (N_3497,In_270,In_2339);
nor U3498 (N_3498,In_2060,In_1264);
nand U3499 (N_3499,In_939,In_1663);
nor U3500 (N_3500,In_2241,In_2254);
nor U3501 (N_3501,In_816,In_1158);
and U3502 (N_3502,In_1222,In_1157);
and U3503 (N_3503,In_845,In_1939);
nor U3504 (N_3504,In_1493,In_1652);
nand U3505 (N_3505,In_2057,In_2137);
and U3506 (N_3506,In_1660,In_1652);
nor U3507 (N_3507,In_501,In_2492);
nor U3508 (N_3508,In_2477,In_528);
and U3509 (N_3509,In_2333,In_129);
nor U3510 (N_3510,In_1934,In_39);
and U3511 (N_3511,In_1806,In_2459);
nand U3512 (N_3512,In_2226,In_752);
and U3513 (N_3513,In_1943,In_103);
nor U3514 (N_3514,In_1846,In_1753);
or U3515 (N_3515,In_1282,In_92);
nor U3516 (N_3516,In_1779,In_2114);
nand U3517 (N_3517,In_1742,In_1214);
and U3518 (N_3518,In_1499,In_834);
or U3519 (N_3519,In_1613,In_1424);
nand U3520 (N_3520,In_539,In_2385);
nor U3521 (N_3521,In_2102,In_1326);
or U3522 (N_3522,In_1452,In_1370);
and U3523 (N_3523,In_179,In_1949);
or U3524 (N_3524,In_120,In_549);
or U3525 (N_3525,In_1796,In_723);
nor U3526 (N_3526,In_1314,In_638);
nor U3527 (N_3527,In_2322,In_732);
nor U3528 (N_3528,In_2037,In_1624);
nand U3529 (N_3529,In_2468,In_1427);
nand U3530 (N_3530,In_1365,In_1702);
nand U3531 (N_3531,In_1180,In_2067);
and U3532 (N_3532,In_478,In_2044);
and U3533 (N_3533,In_2131,In_1424);
nand U3534 (N_3534,In_1920,In_1559);
nand U3535 (N_3535,In_1437,In_2357);
nor U3536 (N_3536,In_1597,In_711);
or U3537 (N_3537,In_1722,In_75);
xor U3538 (N_3538,In_1762,In_1549);
xor U3539 (N_3539,In_514,In_817);
xor U3540 (N_3540,In_1012,In_343);
or U3541 (N_3541,In_2299,In_1858);
and U3542 (N_3542,In_941,In_890);
nand U3543 (N_3543,In_2178,In_811);
nor U3544 (N_3544,In_2426,In_1267);
nand U3545 (N_3545,In_810,In_972);
or U3546 (N_3546,In_1878,In_1572);
nand U3547 (N_3547,In_252,In_1466);
nor U3548 (N_3548,In_1831,In_2323);
nor U3549 (N_3549,In_208,In_1855);
and U3550 (N_3550,In_111,In_958);
nor U3551 (N_3551,In_1816,In_1835);
nor U3552 (N_3552,In_1270,In_661);
and U3553 (N_3553,In_1778,In_998);
or U3554 (N_3554,In_1250,In_1680);
nand U3555 (N_3555,In_288,In_1096);
nor U3556 (N_3556,In_162,In_1547);
and U3557 (N_3557,In_931,In_81);
nor U3558 (N_3558,In_153,In_1468);
nand U3559 (N_3559,In_262,In_1125);
nor U3560 (N_3560,In_1200,In_222);
and U3561 (N_3561,In_993,In_1861);
or U3562 (N_3562,In_1053,In_2479);
xor U3563 (N_3563,In_654,In_309);
or U3564 (N_3564,In_1657,In_1157);
nor U3565 (N_3565,In_191,In_102);
nor U3566 (N_3566,In_1143,In_2128);
nor U3567 (N_3567,In_1087,In_920);
nor U3568 (N_3568,In_1875,In_1659);
or U3569 (N_3569,In_1618,In_344);
nor U3570 (N_3570,In_2151,In_714);
nand U3571 (N_3571,In_281,In_2116);
xnor U3572 (N_3572,In_2075,In_1487);
or U3573 (N_3573,In_2263,In_1233);
nor U3574 (N_3574,In_2487,In_430);
nor U3575 (N_3575,In_779,In_56);
nor U3576 (N_3576,In_1311,In_506);
and U3577 (N_3577,In_854,In_70);
nor U3578 (N_3578,In_914,In_2443);
or U3579 (N_3579,In_501,In_1665);
nor U3580 (N_3580,In_510,In_1397);
or U3581 (N_3581,In_1727,In_445);
nand U3582 (N_3582,In_516,In_1907);
or U3583 (N_3583,In_669,In_522);
nor U3584 (N_3584,In_355,In_2268);
nand U3585 (N_3585,In_172,In_1725);
nand U3586 (N_3586,In_1342,In_654);
nor U3587 (N_3587,In_362,In_1812);
nand U3588 (N_3588,In_2269,In_2256);
or U3589 (N_3589,In_601,In_1438);
or U3590 (N_3590,In_908,In_1644);
and U3591 (N_3591,In_932,In_1136);
or U3592 (N_3592,In_1693,In_842);
or U3593 (N_3593,In_54,In_2486);
nand U3594 (N_3594,In_1965,In_1362);
nand U3595 (N_3595,In_627,In_2248);
and U3596 (N_3596,In_310,In_55);
and U3597 (N_3597,In_2209,In_2080);
and U3598 (N_3598,In_337,In_2141);
nor U3599 (N_3599,In_229,In_1921);
and U3600 (N_3600,In_1100,In_1643);
or U3601 (N_3601,In_920,In_460);
nand U3602 (N_3602,In_263,In_1826);
xnor U3603 (N_3603,In_2314,In_192);
or U3604 (N_3604,In_463,In_637);
and U3605 (N_3605,In_184,In_2341);
nor U3606 (N_3606,In_2427,In_1044);
or U3607 (N_3607,In_1564,In_1203);
or U3608 (N_3608,In_1447,In_1605);
nor U3609 (N_3609,In_284,In_183);
nand U3610 (N_3610,In_352,In_2081);
nor U3611 (N_3611,In_949,In_711);
and U3612 (N_3612,In_1650,In_598);
or U3613 (N_3613,In_1989,In_836);
and U3614 (N_3614,In_1005,In_2478);
and U3615 (N_3615,In_2382,In_220);
nor U3616 (N_3616,In_646,In_2090);
nand U3617 (N_3617,In_1726,In_2052);
nor U3618 (N_3618,In_1949,In_1638);
and U3619 (N_3619,In_729,In_2236);
nor U3620 (N_3620,In_1058,In_99);
nand U3621 (N_3621,In_1625,In_1293);
nor U3622 (N_3622,In_252,In_947);
and U3623 (N_3623,In_2353,In_809);
and U3624 (N_3624,In_1720,In_442);
nor U3625 (N_3625,In_1350,In_1188);
or U3626 (N_3626,In_1469,In_703);
and U3627 (N_3627,In_1415,In_1604);
or U3628 (N_3628,In_141,In_1950);
or U3629 (N_3629,In_504,In_1226);
nor U3630 (N_3630,In_1896,In_2133);
or U3631 (N_3631,In_783,In_2172);
or U3632 (N_3632,In_1961,In_267);
nand U3633 (N_3633,In_499,In_1651);
nand U3634 (N_3634,In_2005,In_658);
or U3635 (N_3635,In_166,In_54);
and U3636 (N_3636,In_975,In_1562);
or U3637 (N_3637,In_520,In_1245);
nor U3638 (N_3638,In_2133,In_163);
or U3639 (N_3639,In_1222,In_1167);
nand U3640 (N_3640,In_819,In_2414);
and U3641 (N_3641,In_1513,In_2371);
nand U3642 (N_3642,In_1692,In_1616);
nand U3643 (N_3643,In_518,In_785);
or U3644 (N_3644,In_561,In_101);
or U3645 (N_3645,In_394,In_569);
or U3646 (N_3646,In_2308,In_1777);
nand U3647 (N_3647,In_533,In_2451);
nand U3648 (N_3648,In_317,In_2151);
or U3649 (N_3649,In_133,In_1616);
xor U3650 (N_3650,In_329,In_1457);
or U3651 (N_3651,In_2121,In_1572);
nor U3652 (N_3652,In_648,In_1339);
nand U3653 (N_3653,In_1273,In_34);
nor U3654 (N_3654,In_876,In_1021);
and U3655 (N_3655,In_1776,In_1682);
nor U3656 (N_3656,In_326,In_1991);
nand U3657 (N_3657,In_12,In_413);
nand U3658 (N_3658,In_1280,In_2015);
or U3659 (N_3659,In_652,In_1361);
nand U3660 (N_3660,In_1250,In_2163);
nor U3661 (N_3661,In_1486,In_260);
nand U3662 (N_3662,In_2314,In_1094);
nand U3663 (N_3663,In_2187,In_1715);
nor U3664 (N_3664,In_338,In_1025);
nand U3665 (N_3665,In_269,In_1438);
nand U3666 (N_3666,In_2079,In_1356);
and U3667 (N_3667,In_1436,In_2140);
or U3668 (N_3668,In_710,In_1760);
nand U3669 (N_3669,In_2386,In_2272);
and U3670 (N_3670,In_719,In_1977);
nor U3671 (N_3671,In_1514,In_2074);
nand U3672 (N_3672,In_2481,In_274);
nor U3673 (N_3673,In_130,In_984);
or U3674 (N_3674,In_522,In_451);
nand U3675 (N_3675,In_1013,In_2067);
nor U3676 (N_3676,In_1534,In_1039);
nor U3677 (N_3677,In_1280,In_195);
or U3678 (N_3678,In_1692,In_463);
or U3679 (N_3679,In_997,In_1458);
or U3680 (N_3680,In_231,In_239);
nand U3681 (N_3681,In_164,In_545);
and U3682 (N_3682,In_1493,In_841);
xnor U3683 (N_3683,In_344,In_1380);
nand U3684 (N_3684,In_882,In_2279);
and U3685 (N_3685,In_549,In_2313);
nor U3686 (N_3686,In_825,In_592);
nor U3687 (N_3687,In_829,In_202);
or U3688 (N_3688,In_1374,In_1166);
or U3689 (N_3689,In_1165,In_251);
nand U3690 (N_3690,In_28,In_143);
and U3691 (N_3691,In_2243,In_1689);
or U3692 (N_3692,In_2401,In_1810);
nor U3693 (N_3693,In_1431,In_2280);
or U3694 (N_3694,In_508,In_732);
nor U3695 (N_3695,In_2020,In_2358);
nor U3696 (N_3696,In_538,In_679);
nor U3697 (N_3697,In_971,In_1070);
and U3698 (N_3698,In_1163,In_2481);
nor U3699 (N_3699,In_625,In_240);
and U3700 (N_3700,In_985,In_1217);
nor U3701 (N_3701,In_1847,In_1830);
or U3702 (N_3702,In_725,In_609);
nand U3703 (N_3703,In_1534,In_2165);
nor U3704 (N_3704,In_1920,In_995);
and U3705 (N_3705,In_1186,In_2498);
and U3706 (N_3706,In_1347,In_1282);
and U3707 (N_3707,In_994,In_251);
or U3708 (N_3708,In_2079,In_198);
nand U3709 (N_3709,In_360,In_2399);
nor U3710 (N_3710,In_833,In_2313);
nand U3711 (N_3711,In_1010,In_2205);
nand U3712 (N_3712,In_2325,In_1876);
nand U3713 (N_3713,In_1355,In_1233);
nor U3714 (N_3714,In_1892,In_897);
nand U3715 (N_3715,In_98,In_799);
nand U3716 (N_3716,In_1276,In_2364);
and U3717 (N_3717,In_1134,In_1524);
or U3718 (N_3718,In_1381,In_925);
and U3719 (N_3719,In_674,In_1230);
and U3720 (N_3720,In_2490,In_149);
and U3721 (N_3721,In_1564,In_79);
or U3722 (N_3722,In_2172,In_2150);
nor U3723 (N_3723,In_1775,In_2288);
nand U3724 (N_3724,In_516,In_2202);
or U3725 (N_3725,In_691,In_1539);
nand U3726 (N_3726,In_2410,In_2185);
or U3727 (N_3727,In_1573,In_2194);
or U3728 (N_3728,In_247,In_2042);
and U3729 (N_3729,In_1494,In_2217);
and U3730 (N_3730,In_63,In_1362);
or U3731 (N_3731,In_2115,In_450);
nor U3732 (N_3732,In_1619,In_2197);
nand U3733 (N_3733,In_1557,In_426);
nand U3734 (N_3734,In_967,In_2338);
or U3735 (N_3735,In_1723,In_2458);
nor U3736 (N_3736,In_1486,In_552);
nor U3737 (N_3737,In_931,In_1584);
or U3738 (N_3738,In_779,In_1569);
nor U3739 (N_3739,In_1617,In_2135);
nand U3740 (N_3740,In_1189,In_1309);
nor U3741 (N_3741,In_2460,In_1542);
and U3742 (N_3742,In_2215,In_1950);
or U3743 (N_3743,In_1150,In_2042);
and U3744 (N_3744,In_254,In_618);
nand U3745 (N_3745,In_1636,In_362);
nand U3746 (N_3746,In_856,In_142);
and U3747 (N_3747,In_1160,In_940);
nand U3748 (N_3748,In_87,In_2151);
or U3749 (N_3749,In_2347,In_1696);
nor U3750 (N_3750,In_1578,In_315);
nor U3751 (N_3751,In_2020,In_731);
and U3752 (N_3752,In_2285,In_2428);
nor U3753 (N_3753,In_1245,In_542);
and U3754 (N_3754,In_1720,In_1960);
nand U3755 (N_3755,In_616,In_836);
or U3756 (N_3756,In_452,In_1355);
and U3757 (N_3757,In_259,In_1174);
and U3758 (N_3758,In_1773,In_1595);
xnor U3759 (N_3759,In_2035,In_23);
nor U3760 (N_3760,In_2227,In_2247);
or U3761 (N_3761,In_1701,In_342);
and U3762 (N_3762,In_198,In_2473);
or U3763 (N_3763,In_752,In_399);
nand U3764 (N_3764,In_99,In_2355);
nor U3765 (N_3765,In_971,In_1278);
nor U3766 (N_3766,In_1985,In_291);
nand U3767 (N_3767,In_2087,In_1464);
and U3768 (N_3768,In_1920,In_393);
nor U3769 (N_3769,In_1563,In_1597);
and U3770 (N_3770,In_751,In_1338);
and U3771 (N_3771,In_1192,In_2477);
nor U3772 (N_3772,In_2340,In_1770);
or U3773 (N_3773,In_45,In_950);
and U3774 (N_3774,In_185,In_624);
nand U3775 (N_3775,In_2455,In_366);
and U3776 (N_3776,In_2017,In_2001);
nor U3777 (N_3777,In_821,In_623);
or U3778 (N_3778,In_571,In_2031);
nor U3779 (N_3779,In_573,In_2366);
nor U3780 (N_3780,In_1665,In_1651);
nand U3781 (N_3781,In_1166,In_321);
or U3782 (N_3782,In_2035,In_367);
or U3783 (N_3783,In_617,In_775);
and U3784 (N_3784,In_733,In_628);
and U3785 (N_3785,In_1027,In_1816);
nand U3786 (N_3786,In_786,In_822);
and U3787 (N_3787,In_922,In_179);
or U3788 (N_3788,In_955,In_410);
nor U3789 (N_3789,In_740,In_1272);
and U3790 (N_3790,In_1191,In_1011);
or U3791 (N_3791,In_669,In_256);
nand U3792 (N_3792,In_1480,In_1360);
and U3793 (N_3793,In_1,In_1459);
nor U3794 (N_3794,In_748,In_2362);
nor U3795 (N_3795,In_1758,In_1960);
and U3796 (N_3796,In_2360,In_1291);
and U3797 (N_3797,In_1233,In_1906);
or U3798 (N_3798,In_531,In_1954);
or U3799 (N_3799,In_892,In_2246);
nor U3800 (N_3800,In_331,In_302);
and U3801 (N_3801,In_876,In_311);
nor U3802 (N_3802,In_1959,In_1796);
nor U3803 (N_3803,In_2024,In_1222);
or U3804 (N_3804,In_1864,In_2137);
and U3805 (N_3805,In_1462,In_1230);
nand U3806 (N_3806,In_1393,In_507);
nand U3807 (N_3807,In_2386,In_1249);
nand U3808 (N_3808,In_2269,In_896);
or U3809 (N_3809,In_1188,In_13);
or U3810 (N_3810,In_130,In_716);
or U3811 (N_3811,In_1132,In_111);
or U3812 (N_3812,In_499,In_2361);
and U3813 (N_3813,In_1929,In_50);
nand U3814 (N_3814,In_985,In_1953);
or U3815 (N_3815,In_1110,In_939);
and U3816 (N_3816,In_148,In_142);
nand U3817 (N_3817,In_1720,In_15);
nand U3818 (N_3818,In_442,In_1289);
and U3819 (N_3819,In_2218,In_1980);
nand U3820 (N_3820,In_2177,In_1827);
and U3821 (N_3821,In_51,In_2449);
nor U3822 (N_3822,In_922,In_1717);
nor U3823 (N_3823,In_1612,In_1082);
or U3824 (N_3824,In_2188,In_1214);
nand U3825 (N_3825,In_2338,In_2266);
or U3826 (N_3826,In_151,In_2082);
and U3827 (N_3827,In_2158,In_1866);
nand U3828 (N_3828,In_1488,In_2239);
nand U3829 (N_3829,In_2352,In_258);
or U3830 (N_3830,In_1329,In_1800);
or U3831 (N_3831,In_2303,In_1858);
or U3832 (N_3832,In_2499,In_1536);
or U3833 (N_3833,In_1214,In_1425);
nor U3834 (N_3834,In_2222,In_358);
nand U3835 (N_3835,In_1612,In_61);
nor U3836 (N_3836,In_62,In_1694);
or U3837 (N_3837,In_308,In_1921);
and U3838 (N_3838,In_316,In_2305);
nand U3839 (N_3839,In_821,In_1997);
nor U3840 (N_3840,In_201,In_974);
nand U3841 (N_3841,In_1544,In_653);
nor U3842 (N_3842,In_2215,In_534);
nor U3843 (N_3843,In_782,In_368);
xnor U3844 (N_3844,In_1007,In_1886);
nand U3845 (N_3845,In_1346,In_2452);
nor U3846 (N_3846,In_2217,In_2345);
and U3847 (N_3847,In_1062,In_259);
and U3848 (N_3848,In_843,In_2237);
nor U3849 (N_3849,In_855,In_103);
or U3850 (N_3850,In_1411,In_1036);
or U3851 (N_3851,In_963,In_2000);
and U3852 (N_3852,In_1888,In_2252);
nand U3853 (N_3853,In_510,In_1851);
nor U3854 (N_3854,In_1287,In_846);
and U3855 (N_3855,In_145,In_692);
or U3856 (N_3856,In_2052,In_1288);
nand U3857 (N_3857,In_734,In_200);
or U3858 (N_3858,In_1580,In_619);
nor U3859 (N_3859,In_535,In_1166);
or U3860 (N_3860,In_925,In_1662);
and U3861 (N_3861,In_2250,In_2138);
and U3862 (N_3862,In_20,In_2023);
and U3863 (N_3863,In_475,In_681);
nor U3864 (N_3864,In_1691,In_1220);
or U3865 (N_3865,In_1208,In_252);
nand U3866 (N_3866,In_1222,In_1354);
nand U3867 (N_3867,In_1458,In_2124);
and U3868 (N_3868,In_758,In_526);
nand U3869 (N_3869,In_2192,In_527);
or U3870 (N_3870,In_2093,In_459);
nor U3871 (N_3871,In_1700,In_2462);
nand U3872 (N_3872,In_2347,In_1554);
and U3873 (N_3873,In_965,In_1568);
nand U3874 (N_3874,In_977,In_774);
or U3875 (N_3875,In_281,In_779);
and U3876 (N_3876,In_930,In_1154);
or U3877 (N_3877,In_562,In_1056);
nor U3878 (N_3878,In_1299,In_2482);
nor U3879 (N_3879,In_2219,In_2067);
and U3880 (N_3880,In_1257,In_2320);
nor U3881 (N_3881,In_918,In_2099);
and U3882 (N_3882,In_1070,In_568);
nor U3883 (N_3883,In_626,In_806);
nor U3884 (N_3884,In_633,In_1467);
or U3885 (N_3885,In_1745,In_2264);
nand U3886 (N_3886,In_1707,In_1172);
and U3887 (N_3887,In_1675,In_2477);
nor U3888 (N_3888,In_1791,In_1384);
nor U3889 (N_3889,In_1012,In_378);
or U3890 (N_3890,In_1727,In_907);
nor U3891 (N_3891,In_1541,In_819);
nand U3892 (N_3892,In_1081,In_1721);
and U3893 (N_3893,In_2167,In_2462);
nand U3894 (N_3894,In_1660,In_2493);
xnor U3895 (N_3895,In_811,In_1288);
nand U3896 (N_3896,In_2074,In_2268);
nand U3897 (N_3897,In_777,In_2177);
or U3898 (N_3898,In_1425,In_357);
or U3899 (N_3899,In_1151,In_1175);
nand U3900 (N_3900,In_2027,In_347);
nor U3901 (N_3901,In_1476,In_1805);
and U3902 (N_3902,In_1567,In_1881);
nand U3903 (N_3903,In_1993,In_988);
or U3904 (N_3904,In_1155,In_570);
nor U3905 (N_3905,In_485,In_1241);
or U3906 (N_3906,In_284,In_1366);
or U3907 (N_3907,In_200,In_1389);
nor U3908 (N_3908,In_824,In_1921);
or U3909 (N_3909,In_363,In_1540);
nor U3910 (N_3910,In_1036,In_1894);
or U3911 (N_3911,In_2021,In_1398);
nand U3912 (N_3912,In_808,In_911);
and U3913 (N_3913,In_882,In_623);
and U3914 (N_3914,In_285,In_1229);
nor U3915 (N_3915,In_1913,In_2446);
nand U3916 (N_3916,In_210,In_501);
and U3917 (N_3917,In_517,In_2319);
nor U3918 (N_3918,In_354,In_1636);
or U3919 (N_3919,In_542,In_310);
nand U3920 (N_3920,In_42,In_2004);
nor U3921 (N_3921,In_607,In_1781);
or U3922 (N_3922,In_1426,In_2388);
and U3923 (N_3923,In_833,In_1096);
nor U3924 (N_3924,In_2392,In_2489);
nor U3925 (N_3925,In_2013,In_61);
or U3926 (N_3926,In_700,In_1984);
nand U3927 (N_3927,In_2142,In_281);
or U3928 (N_3928,In_2114,In_868);
nand U3929 (N_3929,In_2031,In_2186);
nor U3930 (N_3930,In_1108,In_2499);
nor U3931 (N_3931,In_174,In_1567);
or U3932 (N_3932,In_1379,In_1869);
nand U3933 (N_3933,In_1187,In_1014);
nor U3934 (N_3934,In_1051,In_878);
nor U3935 (N_3935,In_444,In_1271);
and U3936 (N_3936,In_2235,In_88);
nand U3937 (N_3937,In_1571,In_1647);
and U3938 (N_3938,In_321,In_644);
nor U3939 (N_3939,In_807,In_2016);
or U3940 (N_3940,In_686,In_7);
and U3941 (N_3941,In_1002,In_1177);
nand U3942 (N_3942,In_1639,In_1397);
nand U3943 (N_3943,In_918,In_74);
and U3944 (N_3944,In_1627,In_2008);
nor U3945 (N_3945,In_138,In_2252);
xnor U3946 (N_3946,In_1737,In_2216);
or U3947 (N_3947,In_2075,In_1095);
nor U3948 (N_3948,In_2449,In_702);
nor U3949 (N_3949,In_364,In_553);
nand U3950 (N_3950,In_1308,In_774);
and U3951 (N_3951,In_1297,In_2042);
nand U3952 (N_3952,In_574,In_63);
or U3953 (N_3953,In_763,In_399);
nor U3954 (N_3954,In_1938,In_616);
nor U3955 (N_3955,In_1405,In_2491);
nand U3956 (N_3956,In_2405,In_946);
or U3957 (N_3957,In_554,In_2384);
nor U3958 (N_3958,In_2180,In_1386);
nand U3959 (N_3959,In_1499,In_266);
nor U3960 (N_3960,In_2270,In_1619);
nor U3961 (N_3961,In_72,In_496);
or U3962 (N_3962,In_1346,In_2496);
nand U3963 (N_3963,In_566,In_1207);
or U3964 (N_3964,In_1247,In_110);
and U3965 (N_3965,In_2007,In_997);
nand U3966 (N_3966,In_1884,In_2105);
nand U3967 (N_3967,In_221,In_1245);
nor U3968 (N_3968,In_279,In_2192);
nor U3969 (N_3969,In_1834,In_1849);
or U3970 (N_3970,In_2364,In_764);
nand U3971 (N_3971,In_627,In_1747);
nand U3972 (N_3972,In_590,In_122);
or U3973 (N_3973,In_1179,In_1376);
or U3974 (N_3974,In_1835,In_2310);
nor U3975 (N_3975,In_969,In_997);
or U3976 (N_3976,In_2054,In_2430);
nor U3977 (N_3977,In_549,In_2045);
or U3978 (N_3978,In_1677,In_1199);
nor U3979 (N_3979,In_2107,In_845);
nand U3980 (N_3980,In_802,In_1350);
nor U3981 (N_3981,In_1516,In_881);
and U3982 (N_3982,In_287,In_1826);
and U3983 (N_3983,In_2005,In_314);
or U3984 (N_3984,In_2206,In_1549);
nand U3985 (N_3985,In_1706,In_344);
or U3986 (N_3986,In_1178,In_121);
xor U3987 (N_3987,In_1676,In_1308);
nor U3988 (N_3988,In_1939,In_1193);
nor U3989 (N_3989,In_483,In_119);
or U3990 (N_3990,In_828,In_1233);
and U3991 (N_3991,In_138,In_1628);
and U3992 (N_3992,In_1208,In_1510);
nand U3993 (N_3993,In_1425,In_1782);
and U3994 (N_3994,In_1656,In_1775);
nand U3995 (N_3995,In_2220,In_1500);
nor U3996 (N_3996,In_1036,In_1250);
nor U3997 (N_3997,In_953,In_303);
nor U3998 (N_3998,In_678,In_1833);
nand U3999 (N_3999,In_1965,In_2097);
or U4000 (N_4000,In_649,In_780);
nor U4001 (N_4001,In_24,In_1616);
and U4002 (N_4002,In_2396,In_644);
nand U4003 (N_4003,In_1443,In_287);
and U4004 (N_4004,In_768,In_728);
and U4005 (N_4005,In_2443,In_1851);
and U4006 (N_4006,In_384,In_42);
nand U4007 (N_4007,In_2187,In_298);
and U4008 (N_4008,In_942,In_503);
nor U4009 (N_4009,In_2282,In_722);
nor U4010 (N_4010,In_2133,In_405);
nor U4011 (N_4011,In_865,In_231);
nor U4012 (N_4012,In_2197,In_2462);
nand U4013 (N_4013,In_987,In_1771);
or U4014 (N_4014,In_147,In_2004);
nand U4015 (N_4015,In_517,In_1285);
nor U4016 (N_4016,In_1881,In_1394);
nand U4017 (N_4017,In_344,In_604);
and U4018 (N_4018,In_74,In_223);
or U4019 (N_4019,In_1156,In_2352);
nand U4020 (N_4020,In_888,In_160);
and U4021 (N_4021,In_1936,In_2188);
and U4022 (N_4022,In_309,In_487);
or U4023 (N_4023,In_347,In_838);
nor U4024 (N_4024,In_259,In_702);
nor U4025 (N_4025,In_2300,In_425);
or U4026 (N_4026,In_288,In_1164);
and U4027 (N_4027,In_1553,In_464);
nor U4028 (N_4028,In_1192,In_1546);
and U4029 (N_4029,In_181,In_2472);
and U4030 (N_4030,In_230,In_1832);
or U4031 (N_4031,In_1297,In_1465);
and U4032 (N_4032,In_1809,In_79);
nor U4033 (N_4033,In_1351,In_514);
nand U4034 (N_4034,In_571,In_393);
or U4035 (N_4035,In_1774,In_1647);
and U4036 (N_4036,In_503,In_1089);
and U4037 (N_4037,In_1107,In_2390);
or U4038 (N_4038,In_1970,In_135);
nand U4039 (N_4039,In_1972,In_454);
and U4040 (N_4040,In_391,In_1035);
nor U4041 (N_4041,In_1020,In_2185);
and U4042 (N_4042,In_783,In_584);
and U4043 (N_4043,In_949,In_880);
nand U4044 (N_4044,In_2186,In_540);
or U4045 (N_4045,In_2493,In_473);
nand U4046 (N_4046,In_2017,In_2298);
nor U4047 (N_4047,In_636,In_1507);
or U4048 (N_4048,In_2470,In_598);
or U4049 (N_4049,In_2317,In_76);
nand U4050 (N_4050,In_113,In_990);
nor U4051 (N_4051,In_394,In_1030);
nand U4052 (N_4052,In_211,In_857);
and U4053 (N_4053,In_1069,In_2481);
xnor U4054 (N_4054,In_1199,In_1552);
and U4055 (N_4055,In_91,In_1474);
nor U4056 (N_4056,In_1390,In_350);
nor U4057 (N_4057,In_2153,In_269);
and U4058 (N_4058,In_1412,In_57);
nor U4059 (N_4059,In_346,In_1402);
or U4060 (N_4060,In_458,In_369);
nor U4061 (N_4061,In_1658,In_241);
nand U4062 (N_4062,In_705,In_1028);
nand U4063 (N_4063,In_2322,In_2286);
or U4064 (N_4064,In_2287,In_741);
and U4065 (N_4065,In_860,In_355);
nor U4066 (N_4066,In_212,In_660);
nand U4067 (N_4067,In_709,In_786);
nor U4068 (N_4068,In_2323,In_2066);
nand U4069 (N_4069,In_1296,In_2218);
or U4070 (N_4070,In_273,In_1069);
nand U4071 (N_4071,In_1598,In_1049);
nor U4072 (N_4072,In_398,In_134);
xnor U4073 (N_4073,In_447,In_401);
or U4074 (N_4074,In_1412,In_86);
nand U4075 (N_4075,In_1848,In_1598);
or U4076 (N_4076,In_1341,In_458);
and U4077 (N_4077,In_2481,In_1707);
or U4078 (N_4078,In_1473,In_1886);
nor U4079 (N_4079,In_1245,In_675);
nor U4080 (N_4080,In_2354,In_458);
nand U4081 (N_4081,In_1818,In_2335);
nor U4082 (N_4082,In_380,In_1223);
or U4083 (N_4083,In_1217,In_2192);
nor U4084 (N_4084,In_905,In_272);
or U4085 (N_4085,In_623,In_905);
nand U4086 (N_4086,In_1529,In_1565);
or U4087 (N_4087,In_2216,In_596);
nor U4088 (N_4088,In_916,In_2361);
nor U4089 (N_4089,In_1592,In_2169);
nor U4090 (N_4090,In_1566,In_2155);
nand U4091 (N_4091,In_2155,In_1289);
and U4092 (N_4092,In_1093,In_702);
nand U4093 (N_4093,In_180,In_719);
and U4094 (N_4094,In_1708,In_1345);
or U4095 (N_4095,In_2460,In_1179);
nand U4096 (N_4096,In_438,In_765);
nand U4097 (N_4097,In_25,In_2296);
nor U4098 (N_4098,In_595,In_823);
nor U4099 (N_4099,In_454,In_2016);
and U4100 (N_4100,In_1168,In_1270);
or U4101 (N_4101,In_1063,In_967);
nor U4102 (N_4102,In_2467,In_1252);
nor U4103 (N_4103,In_880,In_1623);
nand U4104 (N_4104,In_2353,In_746);
and U4105 (N_4105,In_2396,In_256);
nand U4106 (N_4106,In_1248,In_2141);
nand U4107 (N_4107,In_2458,In_1250);
nand U4108 (N_4108,In_411,In_1053);
nand U4109 (N_4109,In_506,In_2148);
and U4110 (N_4110,In_2271,In_1850);
nand U4111 (N_4111,In_1451,In_1914);
and U4112 (N_4112,In_328,In_1856);
or U4113 (N_4113,In_652,In_1507);
and U4114 (N_4114,In_431,In_1435);
and U4115 (N_4115,In_2145,In_2187);
xnor U4116 (N_4116,In_3,In_1755);
nand U4117 (N_4117,In_1296,In_2327);
and U4118 (N_4118,In_743,In_587);
and U4119 (N_4119,In_219,In_1097);
nand U4120 (N_4120,In_1984,In_110);
or U4121 (N_4121,In_890,In_1981);
nor U4122 (N_4122,In_2372,In_921);
xnor U4123 (N_4123,In_1095,In_572);
xor U4124 (N_4124,In_1442,In_1768);
nor U4125 (N_4125,In_1283,In_2370);
xnor U4126 (N_4126,In_212,In_1096);
and U4127 (N_4127,In_218,In_2347);
nor U4128 (N_4128,In_388,In_1587);
and U4129 (N_4129,In_867,In_1010);
nor U4130 (N_4130,In_917,In_1701);
nand U4131 (N_4131,In_2358,In_1080);
and U4132 (N_4132,In_2307,In_1947);
or U4133 (N_4133,In_2206,In_1083);
nand U4134 (N_4134,In_1140,In_1358);
nand U4135 (N_4135,In_478,In_2119);
nand U4136 (N_4136,In_1610,In_954);
nor U4137 (N_4137,In_2351,In_1014);
or U4138 (N_4138,In_2391,In_1070);
nand U4139 (N_4139,In_205,In_931);
nor U4140 (N_4140,In_1911,In_227);
and U4141 (N_4141,In_1602,In_798);
and U4142 (N_4142,In_1486,In_322);
and U4143 (N_4143,In_1326,In_1899);
nand U4144 (N_4144,In_917,In_454);
nand U4145 (N_4145,In_1494,In_846);
nand U4146 (N_4146,In_689,In_1871);
and U4147 (N_4147,In_2099,In_406);
nor U4148 (N_4148,In_937,In_1489);
nor U4149 (N_4149,In_1900,In_793);
and U4150 (N_4150,In_1158,In_324);
or U4151 (N_4151,In_2030,In_2164);
nand U4152 (N_4152,In_543,In_1283);
or U4153 (N_4153,In_1232,In_1164);
nand U4154 (N_4154,In_1596,In_177);
and U4155 (N_4155,In_878,In_1573);
nand U4156 (N_4156,In_2455,In_1651);
xnor U4157 (N_4157,In_191,In_289);
nor U4158 (N_4158,In_70,In_696);
and U4159 (N_4159,In_1664,In_1803);
and U4160 (N_4160,In_823,In_1714);
or U4161 (N_4161,In_1022,In_244);
or U4162 (N_4162,In_1130,In_340);
nand U4163 (N_4163,In_261,In_645);
nor U4164 (N_4164,In_44,In_1104);
and U4165 (N_4165,In_1554,In_2031);
xor U4166 (N_4166,In_18,In_252);
nand U4167 (N_4167,In_1840,In_632);
or U4168 (N_4168,In_797,In_1818);
nand U4169 (N_4169,In_2315,In_2495);
or U4170 (N_4170,In_2042,In_1197);
nor U4171 (N_4171,In_2493,In_2178);
nor U4172 (N_4172,In_738,In_1630);
or U4173 (N_4173,In_1890,In_2272);
and U4174 (N_4174,In_398,In_1412);
and U4175 (N_4175,In_509,In_781);
or U4176 (N_4176,In_440,In_1511);
nor U4177 (N_4177,In_2162,In_694);
nor U4178 (N_4178,In_109,In_1396);
nand U4179 (N_4179,In_1448,In_430);
or U4180 (N_4180,In_920,In_1056);
nor U4181 (N_4181,In_740,In_1842);
nand U4182 (N_4182,In_2126,In_1199);
or U4183 (N_4183,In_1594,In_2066);
nand U4184 (N_4184,In_1599,In_1337);
nor U4185 (N_4185,In_2226,In_547);
nand U4186 (N_4186,In_1301,In_340);
nor U4187 (N_4187,In_1743,In_2320);
nor U4188 (N_4188,In_1199,In_155);
xnor U4189 (N_4189,In_340,In_1720);
or U4190 (N_4190,In_1001,In_1000);
and U4191 (N_4191,In_1332,In_2188);
or U4192 (N_4192,In_2315,In_1102);
and U4193 (N_4193,In_697,In_1065);
or U4194 (N_4194,In_1463,In_722);
nand U4195 (N_4195,In_1360,In_1828);
and U4196 (N_4196,In_302,In_1649);
nand U4197 (N_4197,In_956,In_2292);
xor U4198 (N_4198,In_628,In_592);
nor U4199 (N_4199,In_665,In_906);
or U4200 (N_4200,In_1071,In_2181);
nor U4201 (N_4201,In_2391,In_1704);
and U4202 (N_4202,In_1920,In_1072);
nor U4203 (N_4203,In_644,In_339);
and U4204 (N_4204,In_331,In_179);
or U4205 (N_4205,In_510,In_326);
nor U4206 (N_4206,In_1356,In_1053);
nor U4207 (N_4207,In_900,In_1807);
nand U4208 (N_4208,In_876,In_1106);
nand U4209 (N_4209,In_2450,In_2330);
nor U4210 (N_4210,In_1492,In_1578);
and U4211 (N_4211,In_125,In_1728);
or U4212 (N_4212,In_2377,In_405);
nor U4213 (N_4213,In_1367,In_353);
and U4214 (N_4214,In_31,In_1787);
or U4215 (N_4215,In_828,In_1400);
nand U4216 (N_4216,In_191,In_703);
nand U4217 (N_4217,In_1789,In_1568);
or U4218 (N_4218,In_2198,In_635);
and U4219 (N_4219,In_1182,In_1500);
and U4220 (N_4220,In_1654,In_1218);
or U4221 (N_4221,In_2021,In_1359);
and U4222 (N_4222,In_174,In_2493);
nand U4223 (N_4223,In_314,In_2322);
or U4224 (N_4224,In_2349,In_1417);
nand U4225 (N_4225,In_799,In_1100);
nor U4226 (N_4226,In_218,In_1282);
nand U4227 (N_4227,In_1572,In_1406);
and U4228 (N_4228,In_1308,In_495);
and U4229 (N_4229,In_884,In_1055);
nor U4230 (N_4230,In_292,In_1567);
xnor U4231 (N_4231,In_1213,In_1986);
and U4232 (N_4232,In_482,In_1111);
or U4233 (N_4233,In_1518,In_962);
and U4234 (N_4234,In_1001,In_2202);
nor U4235 (N_4235,In_1218,In_947);
nand U4236 (N_4236,In_834,In_2040);
or U4237 (N_4237,In_901,In_890);
and U4238 (N_4238,In_1026,In_2368);
or U4239 (N_4239,In_806,In_515);
nor U4240 (N_4240,In_1101,In_1286);
nand U4241 (N_4241,In_403,In_1744);
and U4242 (N_4242,In_1890,In_1209);
nor U4243 (N_4243,In_2276,In_949);
and U4244 (N_4244,In_2450,In_1478);
nor U4245 (N_4245,In_1102,In_298);
nor U4246 (N_4246,In_1483,In_947);
and U4247 (N_4247,In_2159,In_1934);
and U4248 (N_4248,In_237,In_1064);
nor U4249 (N_4249,In_1668,In_241);
nor U4250 (N_4250,In_564,In_1899);
or U4251 (N_4251,In_403,In_1468);
nand U4252 (N_4252,In_1525,In_788);
or U4253 (N_4253,In_813,In_318);
nor U4254 (N_4254,In_1934,In_408);
nor U4255 (N_4255,In_1817,In_951);
nand U4256 (N_4256,In_887,In_289);
and U4257 (N_4257,In_256,In_86);
or U4258 (N_4258,In_1333,In_690);
nor U4259 (N_4259,In_2435,In_2396);
or U4260 (N_4260,In_1268,In_1433);
or U4261 (N_4261,In_1701,In_1690);
and U4262 (N_4262,In_1021,In_1517);
xnor U4263 (N_4263,In_2415,In_1967);
nand U4264 (N_4264,In_420,In_1934);
nand U4265 (N_4265,In_2032,In_737);
and U4266 (N_4266,In_1564,In_2420);
or U4267 (N_4267,In_1767,In_158);
nand U4268 (N_4268,In_412,In_394);
nand U4269 (N_4269,In_490,In_327);
nor U4270 (N_4270,In_1948,In_1837);
nor U4271 (N_4271,In_929,In_833);
or U4272 (N_4272,In_244,In_249);
nor U4273 (N_4273,In_2155,In_402);
nor U4274 (N_4274,In_1893,In_1320);
nand U4275 (N_4275,In_276,In_956);
nor U4276 (N_4276,In_779,In_578);
nor U4277 (N_4277,In_25,In_223);
nor U4278 (N_4278,In_2003,In_1148);
nand U4279 (N_4279,In_2238,In_1220);
or U4280 (N_4280,In_1569,In_1602);
or U4281 (N_4281,In_490,In_1010);
xor U4282 (N_4282,In_2440,In_214);
nand U4283 (N_4283,In_2170,In_2281);
and U4284 (N_4284,In_183,In_698);
nor U4285 (N_4285,In_695,In_921);
and U4286 (N_4286,In_620,In_415);
nand U4287 (N_4287,In_2293,In_1024);
or U4288 (N_4288,In_2101,In_901);
and U4289 (N_4289,In_1785,In_1375);
and U4290 (N_4290,In_214,In_1376);
and U4291 (N_4291,In_1568,In_634);
or U4292 (N_4292,In_1810,In_116);
nand U4293 (N_4293,In_2040,In_1471);
nand U4294 (N_4294,In_1480,In_733);
nor U4295 (N_4295,In_1197,In_901);
nand U4296 (N_4296,In_1056,In_1300);
nor U4297 (N_4297,In_1774,In_1752);
nor U4298 (N_4298,In_2359,In_2287);
nor U4299 (N_4299,In_1644,In_1243);
nor U4300 (N_4300,In_2102,In_1680);
nand U4301 (N_4301,In_884,In_1863);
and U4302 (N_4302,In_1190,In_1474);
and U4303 (N_4303,In_332,In_59);
nor U4304 (N_4304,In_2465,In_318);
or U4305 (N_4305,In_2371,In_80);
or U4306 (N_4306,In_204,In_2291);
or U4307 (N_4307,In_2448,In_2010);
and U4308 (N_4308,In_2340,In_475);
and U4309 (N_4309,In_2043,In_1456);
or U4310 (N_4310,In_1745,In_309);
or U4311 (N_4311,In_2101,In_1873);
nand U4312 (N_4312,In_1835,In_1919);
nor U4313 (N_4313,In_1765,In_2170);
or U4314 (N_4314,In_191,In_1921);
and U4315 (N_4315,In_2126,In_2116);
xor U4316 (N_4316,In_1898,In_1976);
and U4317 (N_4317,In_1137,In_1022);
nand U4318 (N_4318,In_167,In_1863);
or U4319 (N_4319,In_2389,In_916);
nand U4320 (N_4320,In_919,In_1298);
nand U4321 (N_4321,In_559,In_686);
or U4322 (N_4322,In_870,In_2286);
or U4323 (N_4323,In_312,In_24);
and U4324 (N_4324,In_1263,In_338);
nand U4325 (N_4325,In_74,In_1526);
nand U4326 (N_4326,In_952,In_1522);
and U4327 (N_4327,In_881,In_298);
nand U4328 (N_4328,In_1625,In_847);
or U4329 (N_4329,In_1524,In_1806);
or U4330 (N_4330,In_344,In_87);
and U4331 (N_4331,In_518,In_1982);
or U4332 (N_4332,In_1483,In_2093);
or U4333 (N_4333,In_851,In_860);
and U4334 (N_4334,In_1582,In_921);
and U4335 (N_4335,In_2491,In_128);
nor U4336 (N_4336,In_123,In_1150);
nand U4337 (N_4337,In_322,In_474);
and U4338 (N_4338,In_2320,In_317);
or U4339 (N_4339,In_2474,In_356);
nor U4340 (N_4340,In_256,In_1890);
or U4341 (N_4341,In_1887,In_2306);
nor U4342 (N_4342,In_74,In_438);
and U4343 (N_4343,In_1833,In_2212);
nor U4344 (N_4344,In_1879,In_726);
nor U4345 (N_4345,In_1349,In_812);
xnor U4346 (N_4346,In_945,In_385);
or U4347 (N_4347,In_1301,In_2134);
nand U4348 (N_4348,In_2432,In_1636);
or U4349 (N_4349,In_1012,In_394);
nand U4350 (N_4350,In_1707,In_1100);
or U4351 (N_4351,In_1712,In_152);
or U4352 (N_4352,In_1884,In_1561);
nor U4353 (N_4353,In_2476,In_330);
nand U4354 (N_4354,In_1138,In_2299);
or U4355 (N_4355,In_242,In_1741);
nor U4356 (N_4356,In_766,In_417);
or U4357 (N_4357,In_270,In_2263);
and U4358 (N_4358,In_1350,In_1178);
and U4359 (N_4359,In_1100,In_1329);
and U4360 (N_4360,In_582,In_1767);
or U4361 (N_4361,In_1723,In_2328);
and U4362 (N_4362,In_1972,In_2228);
xor U4363 (N_4363,In_1848,In_731);
or U4364 (N_4364,In_1355,In_1057);
or U4365 (N_4365,In_270,In_597);
or U4366 (N_4366,In_1412,In_2355);
nand U4367 (N_4367,In_1135,In_1166);
or U4368 (N_4368,In_1091,In_67);
or U4369 (N_4369,In_204,In_1986);
xor U4370 (N_4370,In_943,In_606);
nor U4371 (N_4371,In_1863,In_1174);
nor U4372 (N_4372,In_2055,In_2169);
nand U4373 (N_4373,In_723,In_1082);
and U4374 (N_4374,In_1116,In_2198);
nor U4375 (N_4375,In_810,In_955);
nor U4376 (N_4376,In_1852,In_540);
nor U4377 (N_4377,In_791,In_2129);
or U4378 (N_4378,In_1267,In_54);
and U4379 (N_4379,In_91,In_2242);
or U4380 (N_4380,In_1517,In_430);
and U4381 (N_4381,In_2257,In_1702);
and U4382 (N_4382,In_2295,In_2112);
nor U4383 (N_4383,In_1395,In_1487);
and U4384 (N_4384,In_2108,In_1802);
and U4385 (N_4385,In_2394,In_728);
nor U4386 (N_4386,In_1384,In_385);
or U4387 (N_4387,In_546,In_602);
nand U4388 (N_4388,In_2125,In_633);
nand U4389 (N_4389,In_320,In_921);
and U4390 (N_4390,In_272,In_992);
or U4391 (N_4391,In_454,In_764);
or U4392 (N_4392,In_516,In_1134);
nor U4393 (N_4393,In_321,In_329);
nand U4394 (N_4394,In_1772,In_1898);
and U4395 (N_4395,In_658,In_2238);
and U4396 (N_4396,In_1979,In_1870);
or U4397 (N_4397,In_1693,In_1678);
or U4398 (N_4398,In_418,In_78);
nor U4399 (N_4399,In_796,In_1164);
nor U4400 (N_4400,In_1781,In_746);
and U4401 (N_4401,In_1611,In_94);
nor U4402 (N_4402,In_1755,In_2006);
or U4403 (N_4403,In_1130,In_2217);
nand U4404 (N_4404,In_197,In_59);
or U4405 (N_4405,In_733,In_119);
nand U4406 (N_4406,In_1012,In_1727);
nor U4407 (N_4407,In_225,In_1021);
nand U4408 (N_4408,In_646,In_1615);
nand U4409 (N_4409,In_1091,In_1000);
and U4410 (N_4410,In_1989,In_2329);
and U4411 (N_4411,In_1149,In_594);
and U4412 (N_4412,In_2001,In_2200);
and U4413 (N_4413,In_2482,In_1161);
and U4414 (N_4414,In_1252,In_68);
nand U4415 (N_4415,In_1861,In_750);
or U4416 (N_4416,In_2076,In_701);
and U4417 (N_4417,In_1137,In_540);
or U4418 (N_4418,In_1688,In_2263);
or U4419 (N_4419,In_957,In_132);
or U4420 (N_4420,In_809,In_1560);
nor U4421 (N_4421,In_174,In_1827);
nand U4422 (N_4422,In_1397,In_479);
and U4423 (N_4423,In_885,In_1906);
or U4424 (N_4424,In_1930,In_170);
nand U4425 (N_4425,In_860,In_2153);
nand U4426 (N_4426,In_1285,In_1371);
nand U4427 (N_4427,In_1537,In_190);
and U4428 (N_4428,In_959,In_1818);
nor U4429 (N_4429,In_2175,In_2318);
nand U4430 (N_4430,In_2406,In_1247);
nand U4431 (N_4431,In_1416,In_633);
nor U4432 (N_4432,In_1692,In_1449);
or U4433 (N_4433,In_2114,In_1163);
or U4434 (N_4434,In_1392,In_329);
and U4435 (N_4435,In_2155,In_1368);
or U4436 (N_4436,In_2481,In_332);
or U4437 (N_4437,In_774,In_1853);
nand U4438 (N_4438,In_1585,In_412);
or U4439 (N_4439,In_453,In_2004);
and U4440 (N_4440,In_141,In_1511);
xnor U4441 (N_4441,In_913,In_69);
nor U4442 (N_4442,In_249,In_2428);
and U4443 (N_4443,In_951,In_1315);
or U4444 (N_4444,In_477,In_88);
nor U4445 (N_4445,In_1363,In_1759);
nor U4446 (N_4446,In_2016,In_604);
nand U4447 (N_4447,In_1034,In_1674);
xnor U4448 (N_4448,In_1287,In_2081);
and U4449 (N_4449,In_803,In_673);
nor U4450 (N_4450,In_168,In_1067);
or U4451 (N_4451,In_692,In_716);
nor U4452 (N_4452,In_1915,In_533);
nand U4453 (N_4453,In_1298,In_1909);
nor U4454 (N_4454,In_1129,In_2465);
nand U4455 (N_4455,In_2259,In_1511);
nor U4456 (N_4456,In_563,In_2388);
or U4457 (N_4457,In_1355,In_1666);
and U4458 (N_4458,In_1611,In_1135);
or U4459 (N_4459,In_2355,In_1310);
xor U4460 (N_4460,In_1005,In_1358);
or U4461 (N_4461,In_163,In_827);
nor U4462 (N_4462,In_2058,In_1303);
nand U4463 (N_4463,In_877,In_1039);
xnor U4464 (N_4464,In_1120,In_2454);
or U4465 (N_4465,In_1350,In_1715);
and U4466 (N_4466,In_629,In_1916);
nand U4467 (N_4467,In_504,In_598);
and U4468 (N_4468,In_936,In_1677);
nor U4469 (N_4469,In_2328,In_1990);
or U4470 (N_4470,In_470,In_1136);
nand U4471 (N_4471,In_761,In_309);
or U4472 (N_4472,In_899,In_1416);
nand U4473 (N_4473,In_1692,In_1946);
nand U4474 (N_4474,In_366,In_1880);
nand U4475 (N_4475,In_1080,In_1115);
and U4476 (N_4476,In_2081,In_1158);
nor U4477 (N_4477,In_2027,In_1479);
nand U4478 (N_4478,In_1971,In_6);
and U4479 (N_4479,In_1013,In_949);
and U4480 (N_4480,In_2340,In_676);
or U4481 (N_4481,In_2315,In_1579);
and U4482 (N_4482,In_769,In_521);
nand U4483 (N_4483,In_2195,In_1893);
nand U4484 (N_4484,In_46,In_791);
nor U4485 (N_4485,In_507,In_131);
or U4486 (N_4486,In_450,In_803);
nand U4487 (N_4487,In_1604,In_1761);
and U4488 (N_4488,In_2427,In_285);
nand U4489 (N_4489,In_979,In_533);
or U4490 (N_4490,In_2496,In_2414);
and U4491 (N_4491,In_2286,In_303);
or U4492 (N_4492,In_2370,In_49);
nand U4493 (N_4493,In_946,In_480);
nand U4494 (N_4494,In_593,In_1911);
nor U4495 (N_4495,In_2199,In_601);
and U4496 (N_4496,In_185,In_1059);
nand U4497 (N_4497,In_777,In_791);
nand U4498 (N_4498,In_2433,In_2455);
xor U4499 (N_4499,In_1561,In_753);
or U4500 (N_4500,In_1937,In_2341);
and U4501 (N_4501,In_2296,In_766);
nand U4502 (N_4502,In_701,In_1419);
nor U4503 (N_4503,In_1826,In_1673);
or U4504 (N_4504,In_204,In_1059);
and U4505 (N_4505,In_1894,In_1566);
or U4506 (N_4506,In_2028,In_871);
nor U4507 (N_4507,In_1190,In_1984);
nor U4508 (N_4508,In_181,In_2396);
and U4509 (N_4509,In_974,In_849);
or U4510 (N_4510,In_1339,In_2233);
and U4511 (N_4511,In_1074,In_2459);
nor U4512 (N_4512,In_452,In_1649);
or U4513 (N_4513,In_2046,In_1568);
nor U4514 (N_4514,In_314,In_1542);
nor U4515 (N_4515,In_374,In_1851);
xnor U4516 (N_4516,In_422,In_2400);
or U4517 (N_4517,In_608,In_1896);
and U4518 (N_4518,In_1848,In_823);
or U4519 (N_4519,In_1844,In_828);
nor U4520 (N_4520,In_554,In_375);
nor U4521 (N_4521,In_1449,In_1087);
nand U4522 (N_4522,In_1920,In_1229);
or U4523 (N_4523,In_977,In_656);
nor U4524 (N_4524,In_266,In_1495);
or U4525 (N_4525,In_1002,In_1963);
or U4526 (N_4526,In_43,In_1327);
and U4527 (N_4527,In_1049,In_581);
and U4528 (N_4528,In_760,In_1487);
nor U4529 (N_4529,In_580,In_62);
nor U4530 (N_4530,In_564,In_460);
nor U4531 (N_4531,In_1289,In_488);
or U4532 (N_4532,In_1829,In_1724);
nor U4533 (N_4533,In_2333,In_2305);
and U4534 (N_4534,In_2086,In_1699);
nand U4535 (N_4535,In_338,In_1300);
nor U4536 (N_4536,In_66,In_1626);
and U4537 (N_4537,In_330,In_2397);
or U4538 (N_4538,In_337,In_1393);
or U4539 (N_4539,In_1144,In_1089);
nand U4540 (N_4540,In_795,In_1585);
nand U4541 (N_4541,In_2235,In_592);
nor U4542 (N_4542,In_1653,In_6);
or U4543 (N_4543,In_1069,In_1254);
or U4544 (N_4544,In_541,In_1899);
nor U4545 (N_4545,In_2318,In_438);
and U4546 (N_4546,In_317,In_202);
nand U4547 (N_4547,In_139,In_2377);
and U4548 (N_4548,In_34,In_203);
nand U4549 (N_4549,In_1986,In_534);
and U4550 (N_4550,In_1941,In_2310);
and U4551 (N_4551,In_716,In_854);
or U4552 (N_4552,In_1511,In_1326);
or U4553 (N_4553,In_1731,In_1882);
nor U4554 (N_4554,In_1405,In_2145);
or U4555 (N_4555,In_721,In_573);
or U4556 (N_4556,In_158,In_383);
xnor U4557 (N_4557,In_1023,In_1135);
and U4558 (N_4558,In_1691,In_1831);
or U4559 (N_4559,In_1954,In_473);
or U4560 (N_4560,In_177,In_913);
nand U4561 (N_4561,In_730,In_476);
nor U4562 (N_4562,In_423,In_2185);
nor U4563 (N_4563,In_845,In_419);
nor U4564 (N_4564,In_1365,In_1198);
nor U4565 (N_4565,In_145,In_1757);
nor U4566 (N_4566,In_1802,In_1777);
xor U4567 (N_4567,In_867,In_1354);
nand U4568 (N_4568,In_61,In_645);
or U4569 (N_4569,In_1515,In_1700);
or U4570 (N_4570,In_463,In_2304);
and U4571 (N_4571,In_573,In_1651);
nand U4572 (N_4572,In_41,In_2092);
nand U4573 (N_4573,In_2017,In_1263);
nand U4574 (N_4574,In_524,In_1767);
nor U4575 (N_4575,In_542,In_620);
nand U4576 (N_4576,In_1148,In_2213);
nand U4577 (N_4577,In_2420,In_1083);
nor U4578 (N_4578,In_711,In_1090);
and U4579 (N_4579,In_1004,In_2298);
and U4580 (N_4580,In_659,In_1590);
nor U4581 (N_4581,In_1340,In_465);
nor U4582 (N_4582,In_702,In_2050);
and U4583 (N_4583,In_1827,In_1536);
nor U4584 (N_4584,In_545,In_2243);
and U4585 (N_4585,In_1978,In_1781);
or U4586 (N_4586,In_103,In_159);
nor U4587 (N_4587,In_2482,In_660);
nand U4588 (N_4588,In_847,In_2498);
and U4589 (N_4589,In_857,In_516);
nor U4590 (N_4590,In_786,In_36);
or U4591 (N_4591,In_2204,In_1374);
nand U4592 (N_4592,In_1014,In_694);
nand U4593 (N_4593,In_1312,In_534);
nand U4594 (N_4594,In_1164,In_1894);
nand U4595 (N_4595,In_1624,In_1706);
nand U4596 (N_4596,In_71,In_2179);
nand U4597 (N_4597,In_357,In_1117);
and U4598 (N_4598,In_923,In_2232);
nor U4599 (N_4599,In_604,In_299);
and U4600 (N_4600,In_2444,In_423);
or U4601 (N_4601,In_1697,In_1469);
nand U4602 (N_4602,In_2334,In_615);
nand U4603 (N_4603,In_1929,In_734);
nand U4604 (N_4604,In_603,In_2319);
or U4605 (N_4605,In_802,In_1209);
nand U4606 (N_4606,In_460,In_95);
nor U4607 (N_4607,In_2481,In_1511);
nand U4608 (N_4608,In_623,In_1432);
nand U4609 (N_4609,In_197,In_860);
nor U4610 (N_4610,In_437,In_1100);
and U4611 (N_4611,In_1105,In_2010);
or U4612 (N_4612,In_1446,In_1295);
or U4613 (N_4613,In_1288,In_2196);
nor U4614 (N_4614,In_2394,In_678);
nand U4615 (N_4615,In_1348,In_684);
nand U4616 (N_4616,In_169,In_108);
and U4617 (N_4617,In_738,In_1528);
nand U4618 (N_4618,In_2240,In_1770);
and U4619 (N_4619,In_2059,In_690);
nor U4620 (N_4620,In_1446,In_2020);
and U4621 (N_4621,In_1893,In_588);
and U4622 (N_4622,In_2225,In_2357);
and U4623 (N_4623,In_1357,In_1536);
nor U4624 (N_4624,In_1784,In_636);
and U4625 (N_4625,In_647,In_2174);
nor U4626 (N_4626,In_1901,In_726);
nor U4627 (N_4627,In_2287,In_1802);
nor U4628 (N_4628,In_482,In_1808);
and U4629 (N_4629,In_1173,In_2248);
and U4630 (N_4630,In_1898,In_634);
and U4631 (N_4631,In_1913,In_818);
or U4632 (N_4632,In_740,In_2262);
nor U4633 (N_4633,In_2474,In_1914);
nand U4634 (N_4634,In_1536,In_96);
nand U4635 (N_4635,In_1495,In_1447);
and U4636 (N_4636,In_2276,In_720);
and U4637 (N_4637,In_1772,In_556);
and U4638 (N_4638,In_1162,In_1495);
nor U4639 (N_4639,In_2488,In_1444);
nor U4640 (N_4640,In_1478,In_2009);
nor U4641 (N_4641,In_287,In_1278);
and U4642 (N_4642,In_1048,In_1247);
nand U4643 (N_4643,In_2197,In_336);
nor U4644 (N_4644,In_1570,In_1353);
nand U4645 (N_4645,In_1943,In_1671);
or U4646 (N_4646,In_1576,In_1868);
or U4647 (N_4647,In_2467,In_2256);
nor U4648 (N_4648,In_1967,In_2215);
or U4649 (N_4649,In_2196,In_1193);
or U4650 (N_4650,In_1044,In_504);
or U4651 (N_4651,In_66,In_2119);
nor U4652 (N_4652,In_1848,In_2014);
and U4653 (N_4653,In_597,In_418);
nor U4654 (N_4654,In_1604,In_503);
and U4655 (N_4655,In_1432,In_435);
nor U4656 (N_4656,In_1942,In_2131);
nand U4657 (N_4657,In_256,In_1687);
nand U4658 (N_4658,In_395,In_1983);
nand U4659 (N_4659,In_1462,In_809);
and U4660 (N_4660,In_1888,In_2091);
and U4661 (N_4661,In_1649,In_2201);
nand U4662 (N_4662,In_202,In_2070);
nand U4663 (N_4663,In_134,In_126);
or U4664 (N_4664,In_166,In_2308);
xnor U4665 (N_4665,In_1096,In_1707);
and U4666 (N_4666,In_2323,In_2129);
or U4667 (N_4667,In_1380,In_569);
or U4668 (N_4668,In_77,In_2094);
nor U4669 (N_4669,In_1397,In_2088);
or U4670 (N_4670,In_1935,In_1359);
or U4671 (N_4671,In_1665,In_893);
nand U4672 (N_4672,In_2225,In_1837);
nand U4673 (N_4673,In_2326,In_734);
nand U4674 (N_4674,In_904,In_1245);
and U4675 (N_4675,In_465,In_2475);
nand U4676 (N_4676,In_2334,In_998);
and U4677 (N_4677,In_2264,In_813);
or U4678 (N_4678,In_1770,In_935);
nand U4679 (N_4679,In_1497,In_2240);
nand U4680 (N_4680,In_500,In_899);
and U4681 (N_4681,In_2353,In_2146);
nor U4682 (N_4682,In_115,In_1157);
and U4683 (N_4683,In_1310,In_2033);
nand U4684 (N_4684,In_1239,In_921);
and U4685 (N_4685,In_414,In_1917);
nor U4686 (N_4686,In_2499,In_1517);
or U4687 (N_4687,In_1063,In_300);
nor U4688 (N_4688,In_1177,In_299);
nand U4689 (N_4689,In_1659,In_772);
nand U4690 (N_4690,In_1107,In_374);
and U4691 (N_4691,In_1159,In_485);
nand U4692 (N_4692,In_1022,In_2284);
or U4693 (N_4693,In_54,In_794);
nand U4694 (N_4694,In_1960,In_813);
nor U4695 (N_4695,In_129,In_1720);
or U4696 (N_4696,In_761,In_2361);
nor U4697 (N_4697,In_1413,In_1922);
nor U4698 (N_4698,In_1329,In_1053);
and U4699 (N_4699,In_518,In_872);
or U4700 (N_4700,In_1592,In_1446);
nand U4701 (N_4701,In_1807,In_1768);
nand U4702 (N_4702,In_1687,In_2431);
or U4703 (N_4703,In_1240,In_2196);
nand U4704 (N_4704,In_468,In_576);
or U4705 (N_4705,In_2070,In_2031);
nor U4706 (N_4706,In_1162,In_1028);
nand U4707 (N_4707,In_1422,In_1725);
and U4708 (N_4708,In_1138,In_2421);
or U4709 (N_4709,In_1125,In_2434);
or U4710 (N_4710,In_2432,In_2312);
and U4711 (N_4711,In_1137,In_112);
nor U4712 (N_4712,In_2424,In_1963);
nand U4713 (N_4713,In_39,In_731);
and U4714 (N_4714,In_218,In_425);
nand U4715 (N_4715,In_2423,In_2235);
nand U4716 (N_4716,In_1170,In_2041);
and U4717 (N_4717,In_1681,In_1414);
or U4718 (N_4718,In_541,In_1397);
nand U4719 (N_4719,In_1391,In_251);
nand U4720 (N_4720,In_131,In_1068);
or U4721 (N_4721,In_1657,In_635);
nor U4722 (N_4722,In_110,In_1823);
nor U4723 (N_4723,In_1944,In_1368);
and U4724 (N_4724,In_2274,In_1659);
or U4725 (N_4725,In_1720,In_249);
and U4726 (N_4726,In_177,In_1274);
nand U4727 (N_4727,In_369,In_220);
nand U4728 (N_4728,In_1722,In_1262);
and U4729 (N_4729,In_1658,In_2067);
nand U4730 (N_4730,In_2372,In_401);
or U4731 (N_4731,In_547,In_2402);
nand U4732 (N_4732,In_1164,In_1549);
and U4733 (N_4733,In_1420,In_2163);
nor U4734 (N_4734,In_2140,In_1856);
or U4735 (N_4735,In_2400,In_2290);
and U4736 (N_4736,In_1763,In_82);
nand U4737 (N_4737,In_1040,In_2199);
nor U4738 (N_4738,In_476,In_128);
nor U4739 (N_4739,In_1277,In_478);
and U4740 (N_4740,In_568,In_1445);
nor U4741 (N_4741,In_2013,In_1217);
and U4742 (N_4742,In_2378,In_481);
or U4743 (N_4743,In_107,In_2048);
or U4744 (N_4744,In_2116,In_1559);
or U4745 (N_4745,In_1747,In_1623);
nand U4746 (N_4746,In_2384,In_249);
nand U4747 (N_4747,In_638,In_1304);
or U4748 (N_4748,In_267,In_2470);
nand U4749 (N_4749,In_863,In_2471);
nand U4750 (N_4750,In_1070,In_1708);
nand U4751 (N_4751,In_1453,In_631);
nor U4752 (N_4752,In_599,In_1643);
nand U4753 (N_4753,In_2332,In_1968);
or U4754 (N_4754,In_2057,In_1595);
nand U4755 (N_4755,In_2169,In_781);
xnor U4756 (N_4756,In_1558,In_869);
nor U4757 (N_4757,In_652,In_1841);
nand U4758 (N_4758,In_507,In_1739);
nor U4759 (N_4759,In_2222,In_115);
and U4760 (N_4760,In_1761,In_2475);
nor U4761 (N_4761,In_2272,In_928);
xnor U4762 (N_4762,In_2350,In_217);
nand U4763 (N_4763,In_2214,In_426);
and U4764 (N_4764,In_120,In_772);
nand U4765 (N_4765,In_2067,In_331);
and U4766 (N_4766,In_1216,In_1898);
and U4767 (N_4767,In_442,In_762);
nand U4768 (N_4768,In_2339,In_2328);
and U4769 (N_4769,In_1133,In_1196);
or U4770 (N_4770,In_330,In_348);
or U4771 (N_4771,In_2075,In_391);
nand U4772 (N_4772,In_594,In_269);
or U4773 (N_4773,In_1483,In_1629);
or U4774 (N_4774,In_2496,In_1865);
nand U4775 (N_4775,In_862,In_1159);
or U4776 (N_4776,In_53,In_36);
nand U4777 (N_4777,In_2453,In_499);
nor U4778 (N_4778,In_1469,In_1395);
or U4779 (N_4779,In_483,In_1294);
and U4780 (N_4780,In_1362,In_1826);
nor U4781 (N_4781,In_1567,In_382);
nand U4782 (N_4782,In_62,In_1185);
nor U4783 (N_4783,In_956,In_324);
nor U4784 (N_4784,In_2212,In_1661);
and U4785 (N_4785,In_1353,In_1818);
nand U4786 (N_4786,In_3,In_1224);
xnor U4787 (N_4787,In_1998,In_1311);
and U4788 (N_4788,In_1512,In_1682);
and U4789 (N_4789,In_2345,In_591);
or U4790 (N_4790,In_190,In_1301);
or U4791 (N_4791,In_345,In_748);
nand U4792 (N_4792,In_2309,In_2286);
or U4793 (N_4793,In_744,In_1202);
or U4794 (N_4794,In_203,In_165);
and U4795 (N_4795,In_1027,In_1072);
nand U4796 (N_4796,In_1029,In_2189);
nor U4797 (N_4797,In_1565,In_2159);
nand U4798 (N_4798,In_358,In_87);
nor U4799 (N_4799,In_396,In_2101);
and U4800 (N_4800,In_1451,In_2492);
and U4801 (N_4801,In_2468,In_1020);
and U4802 (N_4802,In_2464,In_1486);
nand U4803 (N_4803,In_1693,In_612);
nand U4804 (N_4804,In_255,In_1772);
and U4805 (N_4805,In_2003,In_250);
nand U4806 (N_4806,In_654,In_970);
nand U4807 (N_4807,In_1740,In_1820);
nand U4808 (N_4808,In_1210,In_595);
nor U4809 (N_4809,In_1191,In_98);
xnor U4810 (N_4810,In_2408,In_2474);
and U4811 (N_4811,In_2009,In_2296);
or U4812 (N_4812,In_42,In_1307);
or U4813 (N_4813,In_749,In_420);
nand U4814 (N_4814,In_2255,In_1115);
nand U4815 (N_4815,In_1498,In_1809);
nand U4816 (N_4816,In_1963,In_592);
and U4817 (N_4817,In_982,In_1812);
and U4818 (N_4818,In_127,In_1928);
or U4819 (N_4819,In_2219,In_887);
and U4820 (N_4820,In_971,In_897);
or U4821 (N_4821,In_1108,In_1297);
and U4822 (N_4822,In_2064,In_1529);
and U4823 (N_4823,In_686,In_145);
and U4824 (N_4824,In_2098,In_892);
or U4825 (N_4825,In_1236,In_2088);
nor U4826 (N_4826,In_1606,In_1451);
or U4827 (N_4827,In_2255,In_679);
nor U4828 (N_4828,In_1180,In_1551);
nor U4829 (N_4829,In_1944,In_246);
or U4830 (N_4830,In_1841,In_894);
or U4831 (N_4831,In_91,In_1303);
or U4832 (N_4832,In_1970,In_2478);
or U4833 (N_4833,In_2130,In_2201);
and U4834 (N_4834,In_1307,In_414);
and U4835 (N_4835,In_1783,In_1357);
nor U4836 (N_4836,In_1877,In_1723);
nand U4837 (N_4837,In_1188,In_112);
nand U4838 (N_4838,In_1822,In_2078);
and U4839 (N_4839,In_1136,In_889);
or U4840 (N_4840,In_2367,In_845);
and U4841 (N_4841,In_489,In_132);
nand U4842 (N_4842,In_2447,In_1782);
nand U4843 (N_4843,In_255,In_822);
or U4844 (N_4844,In_1794,In_313);
nand U4845 (N_4845,In_2087,In_1739);
nor U4846 (N_4846,In_719,In_734);
nand U4847 (N_4847,In_480,In_64);
or U4848 (N_4848,In_1334,In_1063);
nand U4849 (N_4849,In_1271,In_989);
nor U4850 (N_4850,In_849,In_1892);
nand U4851 (N_4851,In_379,In_1907);
and U4852 (N_4852,In_646,In_177);
or U4853 (N_4853,In_437,In_2026);
nand U4854 (N_4854,In_426,In_524);
or U4855 (N_4855,In_1912,In_1583);
nor U4856 (N_4856,In_1600,In_1611);
and U4857 (N_4857,In_648,In_2364);
and U4858 (N_4858,In_1960,In_174);
or U4859 (N_4859,In_1965,In_306);
or U4860 (N_4860,In_406,In_83);
nor U4861 (N_4861,In_1614,In_1416);
nand U4862 (N_4862,In_1945,In_219);
nor U4863 (N_4863,In_1094,In_1038);
nor U4864 (N_4864,In_828,In_2467);
and U4865 (N_4865,In_51,In_1295);
or U4866 (N_4866,In_1767,In_1881);
or U4867 (N_4867,In_780,In_1703);
or U4868 (N_4868,In_715,In_387);
nand U4869 (N_4869,In_222,In_580);
nor U4870 (N_4870,In_938,In_847);
xor U4871 (N_4871,In_65,In_1602);
or U4872 (N_4872,In_1059,In_708);
and U4873 (N_4873,In_1417,In_427);
and U4874 (N_4874,In_1426,In_26);
and U4875 (N_4875,In_325,In_714);
and U4876 (N_4876,In_1717,In_1062);
nor U4877 (N_4877,In_808,In_323);
and U4878 (N_4878,In_686,In_656);
nand U4879 (N_4879,In_817,In_170);
or U4880 (N_4880,In_1383,In_2219);
and U4881 (N_4881,In_25,In_1255);
nand U4882 (N_4882,In_539,In_984);
nor U4883 (N_4883,In_240,In_1422);
and U4884 (N_4884,In_325,In_1211);
and U4885 (N_4885,In_1231,In_483);
nand U4886 (N_4886,In_397,In_1151);
nand U4887 (N_4887,In_2472,In_1193);
nand U4888 (N_4888,In_2392,In_554);
nor U4889 (N_4889,In_576,In_1130);
nor U4890 (N_4890,In_1216,In_465);
nor U4891 (N_4891,In_1637,In_800);
and U4892 (N_4892,In_4,In_635);
and U4893 (N_4893,In_2475,In_1501);
nand U4894 (N_4894,In_194,In_1173);
nor U4895 (N_4895,In_838,In_1402);
nor U4896 (N_4896,In_224,In_641);
nand U4897 (N_4897,In_1638,In_942);
xnor U4898 (N_4898,In_1381,In_974);
or U4899 (N_4899,In_2370,In_338);
nand U4900 (N_4900,In_2358,In_2132);
and U4901 (N_4901,In_1420,In_1298);
xnor U4902 (N_4902,In_1710,In_538);
and U4903 (N_4903,In_1271,In_1109);
and U4904 (N_4904,In_2428,In_2203);
and U4905 (N_4905,In_2122,In_801);
nand U4906 (N_4906,In_872,In_202);
nand U4907 (N_4907,In_566,In_713);
or U4908 (N_4908,In_656,In_1015);
nand U4909 (N_4909,In_1042,In_174);
or U4910 (N_4910,In_1989,In_482);
nor U4911 (N_4911,In_2254,In_560);
nor U4912 (N_4912,In_506,In_1155);
and U4913 (N_4913,In_780,In_1501);
nand U4914 (N_4914,In_2377,In_1624);
nor U4915 (N_4915,In_2003,In_566);
nor U4916 (N_4916,In_147,In_1577);
and U4917 (N_4917,In_1393,In_889);
nor U4918 (N_4918,In_1904,In_1572);
nand U4919 (N_4919,In_926,In_1238);
nor U4920 (N_4920,In_822,In_2392);
xnor U4921 (N_4921,In_2299,In_2274);
nor U4922 (N_4922,In_274,In_495);
and U4923 (N_4923,In_1843,In_882);
xnor U4924 (N_4924,In_39,In_666);
or U4925 (N_4925,In_981,In_2039);
or U4926 (N_4926,In_2304,In_1694);
nand U4927 (N_4927,In_603,In_2035);
and U4928 (N_4928,In_737,In_704);
nor U4929 (N_4929,In_2118,In_538);
nor U4930 (N_4930,In_890,In_723);
or U4931 (N_4931,In_1421,In_305);
nor U4932 (N_4932,In_1423,In_1124);
or U4933 (N_4933,In_696,In_1744);
nand U4934 (N_4934,In_1472,In_674);
nand U4935 (N_4935,In_644,In_65);
or U4936 (N_4936,In_9,In_1126);
nor U4937 (N_4937,In_929,In_2429);
or U4938 (N_4938,In_2137,In_351);
nand U4939 (N_4939,In_2005,In_938);
and U4940 (N_4940,In_335,In_2082);
or U4941 (N_4941,In_842,In_2065);
and U4942 (N_4942,In_215,In_1908);
or U4943 (N_4943,In_1148,In_1213);
nand U4944 (N_4944,In_1368,In_1585);
and U4945 (N_4945,In_827,In_1738);
and U4946 (N_4946,In_1291,In_442);
or U4947 (N_4947,In_942,In_264);
nand U4948 (N_4948,In_73,In_1973);
xor U4949 (N_4949,In_783,In_2364);
nand U4950 (N_4950,In_1870,In_1993);
or U4951 (N_4951,In_1938,In_4);
nand U4952 (N_4952,In_114,In_2314);
or U4953 (N_4953,In_304,In_2445);
and U4954 (N_4954,In_505,In_1537);
nor U4955 (N_4955,In_1576,In_1032);
nor U4956 (N_4956,In_479,In_1404);
xor U4957 (N_4957,In_1850,In_704);
nor U4958 (N_4958,In_2008,In_2007);
and U4959 (N_4959,In_2146,In_2227);
nand U4960 (N_4960,In_1117,In_1277);
or U4961 (N_4961,In_1361,In_2426);
nand U4962 (N_4962,In_2439,In_726);
and U4963 (N_4963,In_483,In_1455);
nand U4964 (N_4964,In_1371,In_672);
nor U4965 (N_4965,In_1256,In_2116);
and U4966 (N_4966,In_996,In_579);
nand U4967 (N_4967,In_879,In_697);
and U4968 (N_4968,In_478,In_1723);
nor U4969 (N_4969,In_400,In_2380);
nand U4970 (N_4970,In_2126,In_2);
nand U4971 (N_4971,In_1516,In_1848);
nor U4972 (N_4972,In_2020,In_833);
or U4973 (N_4973,In_965,In_1326);
xor U4974 (N_4974,In_2447,In_912);
and U4975 (N_4975,In_2254,In_615);
nand U4976 (N_4976,In_79,In_2230);
or U4977 (N_4977,In_2179,In_2147);
xnor U4978 (N_4978,In_2428,In_969);
or U4979 (N_4979,In_840,In_2169);
nand U4980 (N_4980,In_1521,In_1760);
and U4981 (N_4981,In_2145,In_2118);
or U4982 (N_4982,In_349,In_2248);
and U4983 (N_4983,In_1352,In_1914);
nand U4984 (N_4984,In_911,In_440);
nor U4985 (N_4985,In_1461,In_537);
and U4986 (N_4986,In_1598,In_1948);
nor U4987 (N_4987,In_2267,In_1519);
nand U4988 (N_4988,In_2330,In_1656);
and U4989 (N_4989,In_132,In_1991);
nand U4990 (N_4990,In_879,In_750);
and U4991 (N_4991,In_1072,In_246);
or U4992 (N_4992,In_2176,In_158);
xnor U4993 (N_4993,In_2430,In_169);
and U4994 (N_4994,In_1591,In_1181);
nand U4995 (N_4995,In_2113,In_811);
nor U4996 (N_4996,In_2028,In_926);
xor U4997 (N_4997,In_1820,In_2483);
and U4998 (N_4998,In_798,In_1270);
and U4999 (N_4999,In_715,In_1032);
nand U5000 (N_5000,N_2098,N_3474);
or U5001 (N_5001,N_1344,N_3487);
nand U5002 (N_5002,N_610,N_2706);
xnor U5003 (N_5003,N_999,N_4202);
nor U5004 (N_5004,N_4080,N_2390);
nand U5005 (N_5005,N_1660,N_3924);
xor U5006 (N_5006,N_1051,N_4010);
nor U5007 (N_5007,N_3630,N_1274);
xnor U5008 (N_5008,N_2040,N_2104);
nor U5009 (N_5009,N_2264,N_2058);
nor U5010 (N_5010,N_3661,N_404);
or U5011 (N_5011,N_3446,N_3510);
or U5012 (N_5012,N_1960,N_1722);
or U5013 (N_5013,N_1101,N_3895);
nor U5014 (N_5014,N_4078,N_1597);
nand U5015 (N_5015,N_27,N_1943);
or U5016 (N_5016,N_1777,N_2421);
and U5017 (N_5017,N_4687,N_1911);
and U5018 (N_5018,N_4669,N_2169);
and U5019 (N_5019,N_4882,N_2784);
nand U5020 (N_5020,N_3909,N_745);
and U5021 (N_5021,N_3766,N_4626);
nor U5022 (N_5022,N_2577,N_3231);
or U5023 (N_5023,N_640,N_2090);
nand U5024 (N_5024,N_3550,N_1673);
and U5025 (N_5025,N_2665,N_574);
nor U5026 (N_5026,N_3005,N_914);
and U5027 (N_5027,N_4243,N_1255);
nor U5028 (N_5028,N_2267,N_1538);
or U5029 (N_5029,N_1359,N_1225);
nand U5030 (N_5030,N_3320,N_3761);
nand U5031 (N_5031,N_4329,N_4814);
nor U5032 (N_5032,N_2762,N_4156);
and U5033 (N_5033,N_571,N_3720);
nand U5034 (N_5034,N_1298,N_1886);
or U5035 (N_5035,N_3544,N_418);
nor U5036 (N_5036,N_1581,N_118);
and U5037 (N_5037,N_957,N_1682);
nor U5038 (N_5038,N_4664,N_4510);
and U5039 (N_5039,N_464,N_635);
or U5040 (N_5040,N_3883,N_1366);
nor U5041 (N_5041,N_4710,N_4379);
nand U5042 (N_5042,N_3095,N_4138);
and U5043 (N_5043,N_4601,N_383);
nand U5044 (N_5044,N_1213,N_2233);
or U5045 (N_5045,N_3438,N_3684);
nand U5046 (N_5046,N_1358,N_1445);
and U5047 (N_5047,N_4954,N_3532);
and U5048 (N_5048,N_1750,N_3113);
nand U5049 (N_5049,N_3567,N_741);
or U5050 (N_5050,N_1927,N_3491);
and U5051 (N_5051,N_4246,N_155);
nand U5052 (N_5052,N_2862,N_2603);
and U5053 (N_5053,N_805,N_1820);
or U5054 (N_5054,N_221,N_4830);
nand U5055 (N_5055,N_1281,N_750);
or U5056 (N_5056,N_644,N_3069);
or U5057 (N_5057,N_4424,N_1015);
or U5058 (N_5058,N_1694,N_2349);
and U5059 (N_5059,N_2580,N_301);
nor U5060 (N_5060,N_1243,N_2883);
nor U5061 (N_5061,N_3391,N_4183);
or U5062 (N_5062,N_1419,N_4220);
and U5063 (N_5063,N_3549,N_3979);
and U5064 (N_5064,N_3017,N_1356);
xnor U5065 (N_5065,N_3019,N_1007);
and U5066 (N_5066,N_3706,N_4725);
nand U5067 (N_5067,N_2332,N_2326);
or U5068 (N_5068,N_3132,N_3203);
nand U5069 (N_5069,N_2864,N_2994);
or U5070 (N_5070,N_3792,N_2944);
or U5071 (N_5071,N_1476,N_1185);
or U5072 (N_5072,N_2286,N_708);
and U5073 (N_5073,N_1981,N_334);
nand U5074 (N_5074,N_3899,N_1202);
and U5075 (N_5075,N_2441,N_1577);
nor U5076 (N_5076,N_2813,N_237);
nor U5077 (N_5077,N_3617,N_4477);
nand U5078 (N_5078,N_658,N_1721);
and U5079 (N_5079,N_2247,N_385);
and U5080 (N_5080,N_1057,N_1043);
or U5081 (N_5081,N_2878,N_1761);
nand U5082 (N_5082,N_2561,N_1124);
nor U5083 (N_5083,N_3667,N_2625);
nor U5084 (N_5084,N_3837,N_4630);
nand U5085 (N_5085,N_3219,N_1730);
nand U5086 (N_5086,N_216,N_4497);
nand U5087 (N_5087,N_2088,N_1751);
and U5088 (N_5088,N_2036,N_993);
nor U5089 (N_5089,N_1606,N_1857);
nor U5090 (N_5090,N_3879,N_833);
or U5091 (N_5091,N_2719,N_1936);
nand U5092 (N_5092,N_3647,N_423);
and U5093 (N_5093,N_886,N_1004);
nor U5094 (N_5094,N_365,N_4457);
and U5095 (N_5095,N_2854,N_4742);
or U5096 (N_5096,N_3568,N_3271);
or U5097 (N_5097,N_3977,N_2427);
nand U5098 (N_5098,N_1883,N_2263);
and U5099 (N_5099,N_4124,N_3200);
nand U5100 (N_5100,N_3065,N_1129);
nor U5101 (N_5101,N_3082,N_1576);
nor U5102 (N_5102,N_2016,N_375);
nand U5103 (N_5103,N_187,N_1764);
and U5104 (N_5104,N_1700,N_4828);
and U5105 (N_5105,N_2544,N_3664);
nand U5106 (N_5106,N_4875,N_63);
or U5107 (N_5107,N_4729,N_1279);
nand U5108 (N_5108,N_4170,N_579);
nor U5109 (N_5109,N_871,N_1338);
or U5110 (N_5110,N_2078,N_3620);
or U5111 (N_5111,N_3289,N_4652);
nor U5112 (N_5112,N_2428,N_1687);
nand U5113 (N_5113,N_1210,N_4499);
nand U5114 (N_5114,N_2904,N_1941);
nor U5115 (N_5115,N_1417,N_3870);
or U5116 (N_5116,N_1413,N_2395);
nor U5117 (N_5117,N_3756,N_3989);
and U5118 (N_5118,N_1148,N_2309);
or U5119 (N_5119,N_784,N_2193);
and U5120 (N_5120,N_3497,N_620);
nand U5121 (N_5121,N_2621,N_4863);
and U5122 (N_5122,N_169,N_1157);
or U5123 (N_5123,N_1420,N_3830);
nor U5124 (N_5124,N_4118,N_1931);
or U5125 (N_5125,N_3364,N_2844);
nor U5126 (N_5126,N_2879,N_523);
nor U5127 (N_5127,N_3535,N_2414);
or U5128 (N_5128,N_1240,N_4825);
nor U5129 (N_5129,N_4537,N_3359);
nand U5130 (N_5130,N_3418,N_1830);
nand U5131 (N_5131,N_4256,N_2458);
nand U5132 (N_5132,N_539,N_1234);
nor U5133 (N_5133,N_4889,N_1187);
or U5134 (N_5134,N_1042,N_2257);
or U5135 (N_5135,N_2785,N_3758);
nor U5136 (N_5136,N_2492,N_1474);
and U5137 (N_5137,N_1945,N_1726);
nand U5138 (N_5138,N_894,N_4341);
nand U5139 (N_5139,N_2005,N_2516);
and U5140 (N_5140,N_807,N_605);
nor U5141 (N_5141,N_4689,N_3938);
or U5142 (N_5142,N_2092,N_843);
nor U5143 (N_5143,N_1592,N_4273);
nand U5144 (N_5144,N_2687,N_1360);
nand U5145 (N_5145,N_4451,N_1220);
nand U5146 (N_5146,N_3217,N_4475);
or U5147 (N_5147,N_3596,N_1746);
or U5148 (N_5148,N_1778,N_4168);
nand U5149 (N_5149,N_3960,N_577);
nand U5150 (N_5150,N_431,N_3365);
or U5151 (N_5151,N_2788,N_4888);
xor U5152 (N_5152,N_4673,N_4821);
nand U5153 (N_5153,N_1647,N_4539);
and U5154 (N_5154,N_1551,N_3026);
nand U5155 (N_5155,N_1123,N_2117);
or U5156 (N_5156,N_4921,N_1423);
or U5157 (N_5157,N_3945,N_4844);
nand U5158 (N_5158,N_4059,N_3304);
or U5159 (N_5159,N_2979,N_2359);
and U5160 (N_5160,N_119,N_1229);
nand U5161 (N_5161,N_3844,N_535);
nand U5162 (N_5162,N_1033,N_1006);
nand U5163 (N_5163,N_3123,N_4439);
nand U5164 (N_5164,N_2748,N_4019);
and U5165 (N_5165,N_973,N_2314);
nor U5166 (N_5166,N_3441,N_2564);
nor U5167 (N_5167,N_4406,N_1491);
nor U5168 (N_5168,N_1913,N_2658);
xnor U5169 (N_5169,N_2705,N_3654);
nor U5170 (N_5170,N_735,N_3463);
or U5171 (N_5171,N_2137,N_1986);
and U5172 (N_5172,N_508,N_2235);
nand U5173 (N_5173,N_1587,N_4727);
or U5174 (N_5174,N_1780,N_1070);
nor U5175 (N_5175,N_4684,N_585);
and U5176 (N_5176,N_4074,N_1885);
and U5177 (N_5177,N_4883,N_3936);
nor U5178 (N_5178,N_2221,N_3882);
and U5179 (N_5179,N_1457,N_850);
or U5180 (N_5180,N_2899,N_4224);
and U5181 (N_5181,N_2791,N_2674);
or U5182 (N_5182,N_2560,N_1416);
nand U5183 (N_5183,N_3384,N_4544);
nor U5184 (N_5184,N_4775,N_1675);
and U5185 (N_5185,N_1291,N_2799);
and U5186 (N_5186,N_3975,N_2815);
nand U5187 (N_5187,N_4733,N_2639);
nor U5188 (N_5188,N_4219,N_2446);
nor U5189 (N_5189,N_2150,N_3032);
nor U5190 (N_5190,N_562,N_3609);
nand U5191 (N_5191,N_4274,N_4267);
nand U5192 (N_5192,N_1757,N_4460);
or U5193 (N_5193,N_4798,N_1224);
nand U5194 (N_5194,N_359,N_2623);
and U5195 (N_5195,N_46,N_2211);
nor U5196 (N_5196,N_3054,N_622);
and U5197 (N_5197,N_1030,N_4075);
or U5198 (N_5198,N_3188,N_3686);
or U5199 (N_5199,N_2397,N_2461);
nor U5200 (N_5200,N_3395,N_205);
and U5201 (N_5201,N_3416,N_2311);
nor U5202 (N_5202,N_2959,N_878);
nor U5203 (N_5203,N_1045,N_2281);
and U5204 (N_5204,N_3229,N_4643);
nor U5205 (N_5205,N_21,N_695);
nor U5206 (N_5206,N_507,N_2415);
nand U5207 (N_5207,N_288,N_2858);
and U5208 (N_5208,N_4752,N_1353);
and U5209 (N_5209,N_2357,N_1855);
nor U5210 (N_5210,N_1209,N_2116);
or U5211 (N_5211,N_1345,N_3243);
nor U5212 (N_5212,N_3691,N_504);
nand U5213 (N_5213,N_1071,N_2481);
and U5214 (N_5214,N_922,N_1377);
or U5215 (N_5215,N_2283,N_4038);
nor U5216 (N_5216,N_151,N_3230);
nand U5217 (N_5217,N_672,N_3845);
or U5218 (N_5218,N_3457,N_428);
nand U5219 (N_5219,N_236,N_1824);
nand U5220 (N_5220,N_2124,N_302);
nand U5221 (N_5221,N_2042,N_981);
nand U5222 (N_5222,N_4667,N_3294);
or U5223 (N_5223,N_4430,N_2069);
xnor U5224 (N_5224,N_4396,N_3049);
and U5225 (N_5225,N_515,N_76);
nor U5226 (N_5226,N_2228,N_2751);
xnor U5227 (N_5227,N_1912,N_4744);
and U5228 (N_5228,N_4190,N_253);
or U5229 (N_5229,N_797,N_3759);
and U5230 (N_5230,N_3619,N_4618);
nand U5231 (N_5231,N_4125,N_4845);
or U5232 (N_5232,N_3305,N_1284);
nand U5233 (N_5233,N_177,N_454);
or U5234 (N_5234,N_1142,N_701);
nor U5235 (N_5235,N_42,N_1072);
nor U5236 (N_5236,N_2569,N_3744);
nand U5237 (N_5237,N_446,N_4528);
and U5238 (N_5238,N_2523,N_3934);
nor U5239 (N_5239,N_2918,N_4739);
xnor U5240 (N_5240,N_636,N_214);
nor U5241 (N_5241,N_3947,N_3990);
nor U5242 (N_5242,N_2158,N_1181);
nor U5243 (N_5243,N_4975,N_1866);
nand U5244 (N_5244,N_737,N_2012);
nand U5245 (N_5245,N_171,N_4226);
nand U5246 (N_5246,N_4732,N_2726);
or U5247 (N_5247,N_4992,N_3774);
or U5248 (N_5248,N_2660,N_4134);
nor U5249 (N_5249,N_1381,N_4550);
or U5250 (N_5250,N_615,N_3927);
nor U5251 (N_5251,N_4536,N_3861);
or U5252 (N_5252,N_3961,N_4015);
and U5253 (N_5253,N_3907,N_2304);
nand U5254 (N_5254,N_1816,N_2070);
nor U5255 (N_5255,N_4867,N_2472);
nor U5256 (N_5256,N_2554,N_2373);
or U5257 (N_5257,N_1590,N_2491);
and U5258 (N_5258,N_4769,N_40);
xor U5259 (N_5259,N_3075,N_4611);
nand U5260 (N_5260,N_1292,N_4913);
or U5261 (N_5261,N_486,N_3660);
nor U5262 (N_5262,N_3878,N_3555);
nand U5263 (N_5263,N_1488,N_1792);
and U5264 (N_5264,N_2614,N_1485);
or U5265 (N_5265,N_4011,N_4456);
xor U5266 (N_5266,N_4209,N_2924);
nor U5267 (N_5267,N_3712,N_2974);
nand U5268 (N_5268,N_324,N_1343);
nor U5269 (N_5269,N_4301,N_2379);
nor U5270 (N_5270,N_433,N_4143);
or U5271 (N_5271,N_3740,N_4068);
or U5272 (N_5272,N_1075,N_1900);
nand U5273 (N_5273,N_4187,N_2175);
and U5274 (N_5274,N_4440,N_378);
and U5275 (N_5275,N_2853,N_4251);
nor U5276 (N_5276,N_3378,N_3625);
nand U5277 (N_5277,N_597,N_624);
nor U5278 (N_5278,N_4325,N_2723);
or U5279 (N_5279,N_0,N_4351);
nand U5280 (N_5280,N_2619,N_1283);
and U5281 (N_5281,N_4496,N_3454);
nand U5282 (N_5282,N_4271,N_4278);
or U5283 (N_5283,N_3949,N_2778);
nand U5284 (N_5284,N_3502,N_1953);
nor U5285 (N_5285,N_3914,N_958);
nor U5286 (N_5286,N_2123,N_3615);
nand U5287 (N_5287,N_4280,N_2287);
and U5288 (N_5288,N_4487,N_2322);
or U5289 (N_5289,N_1670,N_1002);
xor U5290 (N_5290,N_657,N_2195);
nand U5291 (N_5291,N_2252,N_3876);
or U5292 (N_5292,N_3117,N_2896);
nor U5293 (N_5293,N_4816,N_50);
or U5294 (N_5294,N_3853,N_1685);
or U5295 (N_5295,N_2488,N_942);
nor U5296 (N_5296,N_2900,N_3077);
nand U5297 (N_5297,N_3473,N_890);
nand U5298 (N_5298,N_348,N_2120);
or U5299 (N_5299,N_592,N_1989);
and U5300 (N_5300,N_1511,N_3517);
nand U5301 (N_5301,N_3492,N_2850);
and U5302 (N_5302,N_799,N_1863);
nor U5303 (N_5303,N_678,N_2889);
and U5304 (N_5304,N_1378,N_1973);
nor U5305 (N_5305,N_4211,N_275);
nor U5306 (N_5306,N_2769,N_566);
nand U5307 (N_5307,N_4859,N_1658);
and U5308 (N_5308,N_1979,N_4270);
or U5309 (N_5309,N_1742,N_2023);
nor U5310 (N_5310,N_4257,N_3437);
and U5311 (N_5311,N_2021,N_3786);
and U5312 (N_5312,N_1138,N_2581);
and U5313 (N_5313,N_1846,N_1582);
nor U5314 (N_5314,N_3632,N_2392);
nor U5315 (N_5315,N_903,N_3805);
nand U5316 (N_5316,N_1957,N_2295);
or U5317 (N_5317,N_606,N_3973);
nor U5318 (N_5318,N_1354,N_1003);
nand U5319 (N_5319,N_2125,N_1940);
or U5320 (N_5320,N_4206,N_3081);
or U5321 (N_5321,N_2672,N_1087);
nor U5322 (N_5322,N_3920,N_800);
nand U5323 (N_5323,N_2893,N_2503);
nand U5324 (N_5324,N_1231,N_1479);
nor U5325 (N_5325,N_1781,N_4425);
or U5326 (N_5326,N_927,N_959);
nand U5327 (N_5327,N_2310,N_1013);
nand U5328 (N_5328,N_645,N_1517);
nor U5329 (N_5329,N_2215,N_2616);
or U5330 (N_5330,N_744,N_4833);
nand U5331 (N_5331,N_400,N_1654);
or U5332 (N_5332,N_4861,N_3445);
nor U5333 (N_5333,N_2184,N_3571);
xor U5334 (N_5334,N_35,N_3925);
and U5335 (N_5335,N_2777,N_3121);
nor U5336 (N_5336,N_4149,N_4549);
nor U5337 (N_5337,N_1390,N_4616);
and U5338 (N_5338,N_4355,N_3963);
nand U5339 (N_5339,N_182,N_2056);
or U5340 (N_5340,N_338,N_3149);
and U5341 (N_5341,N_3577,N_341);
and U5342 (N_5342,N_3295,N_3504);
or U5343 (N_5343,N_3701,N_4057);
or U5344 (N_5344,N_145,N_2370);
nor U5345 (N_5345,N_1336,N_4344);
nand U5346 (N_5346,N_2,N_3073);
nand U5347 (N_5347,N_3103,N_1162);
or U5348 (N_5348,N_3164,N_1672);
nand U5349 (N_5349,N_2970,N_70);
nand U5350 (N_5350,N_3591,N_361);
nor U5351 (N_5351,N_4512,N_3828);
nor U5352 (N_5352,N_4426,N_3213);
nor U5353 (N_5353,N_3848,N_4455);
and U5354 (N_5354,N_4965,N_4051);
or U5355 (N_5355,N_2948,N_1559);
and U5356 (N_5356,N_4926,N_720);
and U5357 (N_5357,N_3275,N_1106);
and U5358 (N_5358,N_4395,N_4552);
or U5359 (N_5359,N_505,N_3223);
and U5360 (N_5360,N_3102,N_3602);
or U5361 (N_5361,N_4304,N_3776);
nand U5362 (N_5362,N_2266,N_1405);
xor U5363 (N_5363,N_1332,N_1422);
and U5364 (N_5364,N_1659,N_3150);
nor U5365 (N_5365,N_474,N_4297);
nand U5366 (N_5366,N_1314,N_4158);
or U5367 (N_5367,N_671,N_2216);
nor U5368 (N_5368,N_3037,N_791);
and U5369 (N_5369,N_2693,N_38);
nor U5370 (N_5370,N_4152,N_4827);
nand U5371 (N_5371,N_3721,N_242);
nor U5372 (N_5372,N_1618,N_2207);
or U5373 (N_5373,N_1619,N_4824);
nand U5374 (N_5374,N_4576,N_3478);
or U5375 (N_5375,N_291,N_2246);
and U5376 (N_5376,N_1621,N_2647);
nand U5377 (N_5377,N_3593,N_126);
nor U5378 (N_5378,N_2841,N_2015);
or U5379 (N_5379,N_2008,N_4698);
nor U5380 (N_5380,N_772,N_1341);
and U5381 (N_5381,N_1199,N_1985);
and U5382 (N_5382,N_2499,N_4398);
nor U5383 (N_5383,N_2327,N_49);
nand U5384 (N_5384,N_4945,N_1990);
and U5385 (N_5385,N_103,N_2411);
or U5386 (N_5386,N_4334,N_4951);
nor U5387 (N_5387,N_482,N_1882);
nor U5388 (N_5388,N_1014,N_1056);
or U5389 (N_5389,N_4041,N_1444);
nand U5390 (N_5390,N_686,N_4592);
nor U5391 (N_5391,N_3493,N_4392);
or U5392 (N_5392,N_3906,N_2869);
nand U5393 (N_5393,N_3042,N_1270);
nor U5394 (N_5394,N_1130,N_1200);
or U5395 (N_5395,N_638,N_3433);
nor U5396 (N_5396,N_2405,N_2248);
nor U5397 (N_5397,N_4638,N_4035);
or U5398 (N_5398,N_4708,N_274);
or U5399 (N_5399,N_3682,N_4786);
and U5400 (N_5400,N_1260,N_1723);
nor U5401 (N_5401,N_4350,N_2294);
or U5402 (N_5402,N_891,N_1430);
and U5403 (N_5403,N_699,N_3405);
nand U5404 (N_5404,N_3900,N_1891);
nor U5405 (N_5405,N_2757,N_556);
or U5406 (N_5406,N_3018,N_918);
and U5407 (N_5407,N_163,N_80);
and U5408 (N_5408,N_3827,N_4409);
xnor U5409 (N_5409,N_1942,N_2060);
nand U5410 (N_5410,N_2431,N_3672);
or U5411 (N_5411,N_4373,N_3783);
and U5412 (N_5412,N_971,N_1712);
nand U5413 (N_5413,N_3265,N_4346);
and U5414 (N_5414,N_2825,N_2513);
and U5415 (N_5415,N_1546,N_1005);
xnor U5416 (N_5416,N_3133,N_905);
nor U5417 (N_5417,N_1790,N_292);
nand U5418 (N_5418,N_2276,N_2102);
and U5419 (N_5419,N_94,N_2548);
and U5420 (N_5420,N_239,N_2677);
or U5421 (N_5421,N_2911,N_3059);
and U5422 (N_5422,N_3051,N_3980);
nor U5423 (N_5423,N_2832,N_803);
nand U5424 (N_5424,N_3542,N_2562);
nor U5425 (N_5425,N_3987,N_223);
nor U5426 (N_5426,N_3892,N_1939);
nor U5427 (N_5427,N_3604,N_1203);
nand U5428 (N_5428,N_3588,N_4122);
nand U5429 (N_5429,N_2097,N_412);
and U5430 (N_5430,N_3551,N_4879);
or U5431 (N_5431,N_945,N_4320);
xnor U5432 (N_5432,N_4826,N_4466);
xor U5433 (N_5433,N_3525,N_4383);
nand U5434 (N_5434,N_2836,N_3125);
and U5435 (N_5435,N_321,N_950);
nand U5436 (N_5436,N_1897,N_2131);
nor U5437 (N_5437,N_3109,N_688);
or U5438 (N_5438,N_848,N_4401);
nor U5439 (N_5439,N_3965,N_3107);
nor U5440 (N_5440,N_3098,N_4144);
or U5441 (N_5441,N_3689,N_600);
nand U5442 (N_5442,N_2775,N_4255);
nand U5443 (N_5443,N_246,N_1921);
and U5444 (N_5444,N_2100,N_3386);
and U5445 (N_5445,N_3880,N_3648);
nor U5446 (N_5446,N_254,N_2676);
nand U5447 (N_5447,N_923,N_628);
nand U5448 (N_5448,N_1829,N_1835);
or U5449 (N_5449,N_757,N_1902);
or U5450 (N_5450,N_3262,N_1168);
and U5451 (N_5451,N_55,N_4785);
and U5452 (N_5452,N_1278,N_1585);
xnor U5453 (N_5453,N_4995,N_4461);
and U5454 (N_5454,N_4422,N_661);
and U5455 (N_5455,N_3376,N_2149);
nand U5456 (N_5456,N_676,N_3822);
nor U5457 (N_5457,N_4818,N_4088);
and U5458 (N_5458,N_3206,N_3523);
nand U5459 (N_5459,N_3291,N_4612);
or U5460 (N_5460,N_3972,N_4864);
or U5461 (N_5461,N_4868,N_3351);
or U5462 (N_5462,N_2052,N_832);
or U5463 (N_5463,N_2934,N_824);
nor U5464 (N_5464,N_430,N_4751);
nor U5465 (N_5465,N_441,N_1348);
xor U5466 (N_5466,N_2200,N_4071);
nand U5467 (N_5467,N_4145,N_1331);
and U5468 (N_5468,N_4628,N_1550);
nor U5469 (N_5469,N_3940,N_1612);
and U5470 (N_5470,N_866,N_1076);
nand U5471 (N_5471,N_4121,N_892);
nor U5472 (N_5472,N_4623,N_1428);
and U5473 (N_5473,N_1692,N_3736);
nor U5474 (N_5474,N_1770,N_1650);
nor U5475 (N_5475,N_1347,N_473);
or U5476 (N_5476,N_1704,N_1561);
nand U5477 (N_5477,N_435,N_1055);
or U5478 (N_5478,N_1481,N_4666);
and U5479 (N_5479,N_874,N_2921);
or U5480 (N_5480,N_1140,N_32);
and U5481 (N_5481,N_3015,N_2291);
nor U5482 (N_5482,N_2133,N_829);
or U5483 (N_5483,N_3572,N_3310);
nand U5484 (N_5484,N_4159,N_4822);
and U5485 (N_5485,N_448,N_3997);
nand U5486 (N_5486,N_2394,N_1452);
and U5487 (N_5487,N_1933,N_1321);
nor U5488 (N_5488,N_912,N_1465);
nor U5489 (N_5489,N_1048,N_2227);
or U5490 (N_5490,N_2801,N_444);
and U5491 (N_5491,N_178,N_329);
or U5492 (N_5492,N_1573,N_1806);
or U5493 (N_5493,N_2075,N_4047);
or U5494 (N_5494,N_1242,N_2375);
nand U5495 (N_5495,N_1178,N_818);
and U5496 (N_5496,N_1988,N_4902);
or U5497 (N_5497,N_4791,N_170);
or U5498 (N_5498,N_3426,N_4268);
nor U5499 (N_5499,N_4363,N_1808);
nand U5500 (N_5500,N_2447,N_61);
or U5501 (N_5501,N_1424,N_4558);
nand U5502 (N_5502,N_3515,N_255);
and U5503 (N_5503,N_4369,N_3599);
or U5504 (N_5504,N_4186,N_1272);
or U5505 (N_5505,N_325,N_1276);
xor U5506 (N_5506,N_573,N_4155);
and U5507 (N_5507,N_2416,N_2508);
nand U5508 (N_5508,N_1901,N_96);
nand U5509 (N_5509,N_1873,N_2781);
or U5510 (N_5510,N_1850,N_4343);
nand U5511 (N_5511,N_1991,N_339);
nand U5512 (N_5512,N_3236,N_2527);
and U5513 (N_5513,N_2826,N_2789);
nand U5514 (N_5514,N_1614,N_2681);
or U5515 (N_5515,N_2939,N_3890);
nor U5516 (N_5516,N_3677,N_1477);
nor U5517 (N_5517,N_3247,N_1074);
and U5518 (N_5518,N_687,N_4543);
nand U5519 (N_5519,N_3272,N_3919);
nand U5520 (N_5520,N_4520,N_1096);
nand U5521 (N_5521,N_1807,N_390);
nor U5522 (N_5522,N_3719,N_2689);
and U5523 (N_5523,N_2337,N_3613);
nor U5524 (N_5524,N_2312,N_4624);
or U5525 (N_5525,N_2296,N_1545);
nor U5526 (N_5526,N_4709,N_2967);
nand U5527 (N_5527,N_4681,N_2540);
nand U5528 (N_5528,N_1066,N_2958);
and U5529 (N_5529,N_2897,N_436);
nand U5530 (N_5530,N_2507,N_2145);
and U5531 (N_5531,N_1357,N_3586);
or U5532 (N_5532,N_2086,N_194);
nor U5533 (N_5533,N_2685,N_1475);
or U5534 (N_5534,N_3791,N_4016);
and U5535 (N_5535,N_2521,N_4087);
xor U5536 (N_5536,N_4738,N_2340);
and U5537 (N_5537,N_419,N_3855);
or U5538 (N_5538,N_3872,N_2985);
xor U5539 (N_5539,N_117,N_703);
nand U5540 (N_5540,N_1399,N_4541);
xor U5541 (N_5541,N_4629,N_1400);
or U5542 (N_5542,N_3450,N_1251);
xor U5543 (N_5543,N_955,N_3420);
nor U5544 (N_5544,N_2196,N_1152);
or U5545 (N_5545,N_4340,N_3939);
or U5546 (N_5546,N_279,N_3499);
or U5547 (N_5547,N_634,N_2001);
nor U5548 (N_5548,N_1163,N_3464);
or U5549 (N_5549,N_1232,N_3190);
nand U5550 (N_5550,N_3142,N_4571);
or U5551 (N_5551,N_2057,N_2420);
and U5552 (N_5552,N_1832,N_4869);
or U5553 (N_5553,N_3244,N_3519);
nor U5554 (N_5554,N_4846,N_3000);
or U5555 (N_5555,N_4436,N_4419);
or U5556 (N_5556,N_4820,N_598);
nor U5557 (N_5557,N_4476,N_2803);
nand U5558 (N_5558,N_2444,N_3531);
nand U5559 (N_5559,N_651,N_2122);
and U5560 (N_5560,N_518,N_4655);
and U5561 (N_5561,N_1728,N_3157);
and U5562 (N_5562,N_1489,N_1306);
nor U5563 (N_5563,N_232,N_3564);
nor U5564 (N_5564,N_1646,N_2456);
or U5565 (N_5565,N_3085,N_2535);
nand U5566 (N_5566,N_1001,N_2018);
nand U5567 (N_5567,N_4631,N_1916);
and U5568 (N_5568,N_2747,N_1480);
nor U5569 (N_5569,N_1190,N_4091);
nor U5570 (N_5570,N_377,N_459);
or U5571 (N_5571,N_533,N_2584);
or U5572 (N_5572,N_4956,N_4500);
or U5573 (N_5573,N_2663,N_1035);
nor U5574 (N_5574,N_1880,N_4702);
and U5575 (N_5575,N_4117,N_2118);
nand U5576 (N_5576,N_322,N_777);
and U5577 (N_5577,N_1233,N_3657);
nor U5578 (N_5578,N_1340,N_1024);
and U5579 (N_5579,N_3444,N_2429);
nand U5580 (N_5580,N_3352,N_3723);
nand U5581 (N_5581,N_3024,N_528);
and U5582 (N_5582,N_3253,N_2720);
or U5583 (N_5583,N_3583,N_4384);
or U5584 (N_5584,N_207,N_3483);
and U5585 (N_5585,N_3545,N_2599);
nand U5586 (N_5586,N_1814,N_2729);
nand U5587 (N_5587,N_3226,N_732);
nand U5588 (N_5588,N_2376,N_1460);
or U5589 (N_5589,N_3214,N_4431);
nand U5590 (N_5590,N_1161,N_1403);
nor U5591 (N_5591,N_296,N_3366);
xor U5592 (N_5592,N_4692,N_2352);
and U5593 (N_5593,N_1890,N_1164);
and U5594 (N_5594,N_2710,N_4388);
and U5595 (N_5595,N_780,N_1724);
nand U5596 (N_5596,N_4916,N_1908);
and U5597 (N_5597,N_1553,N_189);
nand U5598 (N_5598,N_583,N_1745);
nand U5599 (N_5599,N_764,N_2998);
and U5600 (N_5600,N_1826,N_3179);
nor U5601 (N_5601,N_2319,N_406);
nor U5602 (N_5602,N_1392,N_519);
nor U5603 (N_5603,N_3600,N_452);
nand U5604 (N_5604,N_3933,N_3823);
and U5605 (N_5605,N_2237,N_789);
nand U5606 (N_5606,N_2372,N_66);
or U5607 (N_5607,N_1391,N_4627);
or U5608 (N_5608,N_873,N_4311);
and U5609 (N_5609,N_1666,N_1552);
and U5610 (N_5610,N_3715,N_2992);
and U5611 (N_5611,N_921,N_2163);
and U5612 (N_5612,N_1729,N_1818);
nand U5613 (N_5613,N_2511,N_1868);
and U5614 (N_5614,N_3072,N_907);
or U5615 (N_5615,N_3948,N_1668);
and U5616 (N_5616,N_4399,N_4967);
or U5617 (N_5617,N_29,N_370);
nor U5618 (N_5618,N_1305,N_4728);
or U5619 (N_5619,N_623,N_4778);
nand U5620 (N_5620,N_1128,N_2793);
nand U5621 (N_5621,N_14,N_2270);
and U5622 (N_5622,N_1793,N_4313);
and U5623 (N_5623,N_771,N_1875);
xnor U5624 (N_5624,N_3280,N_2205);
or U5625 (N_5625,N_3982,N_3857);
nor U5626 (N_5626,N_4195,N_2419);
or U5627 (N_5627,N_1257,N_4260);
nand U5628 (N_5628,N_3607,N_2528);
nand U5629 (N_5629,N_367,N_3419);
nor U5630 (N_5630,N_4377,N_3813);
nor U5631 (N_5631,N_3831,N_1368);
nand U5632 (N_5632,N_4222,N_1259);
nor U5633 (N_5633,N_1246,N_3821);
nor U5634 (N_5634,N_4575,N_991);
and U5635 (N_5635,N_1955,N_4939);
or U5636 (N_5636,N_3374,N_1333);
and U5637 (N_5637,N_3193,N_3518);
or U5638 (N_5638,N_3699,N_3528);
nand U5639 (N_5639,N_839,N_3292);
nor U5640 (N_5640,N_2568,N_391);
nand U5641 (N_5641,N_1789,N_2526);
nor U5642 (N_5642,N_3184,N_2017);
nand U5643 (N_5643,N_4375,N_277);
or U5644 (N_5644,N_4971,N_3658);
nand U5645 (N_5645,N_1113,N_1895);
nor U5646 (N_5646,N_4238,N_3700);
nor U5647 (N_5647,N_2978,N_4447);
or U5648 (N_5648,N_3237,N_884);
or U5649 (N_5649,N_362,N_17);
and U5650 (N_5650,N_2643,N_2324);
nand U5651 (N_5651,N_4443,N_3057);
or U5652 (N_5652,N_272,N_88);
nand U5653 (N_5653,N_1827,N_887);
and U5654 (N_5654,N_3479,N_3239);
nand U5655 (N_5655,N_57,N_1533);
nand U5656 (N_5656,N_4730,N_3768);
and U5657 (N_5657,N_337,N_4694);
and U5658 (N_5658,N_4448,N_2305);
and U5659 (N_5659,N_2068,N_3091);
or U5660 (N_5660,N_2880,N_4890);
nand U5661 (N_5661,N_608,N_512);
xor U5662 (N_5662,N_2635,N_4205);
nand U5663 (N_5663,N_395,N_698);
and U5664 (N_5664,N_1586,N_3313);
and U5665 (N_5665,N_217,N_3401);
nor U5666 (N_5666,N_4175,N_2204);
nand U5667 (N_5667,N_1851,N_352);
and U5668 (N_5668,N_4482,N_3299);
nor U5669 (N_5669,N_4050,N_3178);
nor U5670 (N_5670,N_2545,N_54);
nand U5671 (N_5671,N_3819,N_2358);
nand U5672 (N_5672,N_809,N_3833);
or U5673 (N_5673,N_2675,N_4342);
nand U5674 (N_5674,N_2460,N_3516);
or U5675 (N_5675,N_3290,N_1068);
and U5676 (N_5676,N_2838,N_294);
or U5677 (N_5677,N_2301,N_4855);
and U5678 (N_5678,N_3735,N_555);
or U5679 (N_5679,N_1570,N_1389);
or U5680 (N_5680,N_2566,N_984);
and U5681 (N_5681,N_897,N_4298);
nor U5682 (N_5682,N_1756,N_3155);
or U5683 (N_5683,N_75,N_3012);
nand U5684 (N_5684,N_1227,N_2082);
or U5685 (N_5685,N_1296,N_3603);
nand U5686 (N_5686,N_4173,N_1714);
nor U5687 (N_5687,N_2901,N_664);
or U5688 (N_5688,N_184,N_1174);
xor U5689 (N_5689,N_1387,N_4840);
or U5690 (N_5690,N_1616,N_4160);
xor U5691 (N_5691,N_1644,N_2667);
or U5692 (N_5692,N_4044,N_305);
nor U5693 (N_5693,N_3199,N_295);
or U5694 (N_5694,N_4005,N_1059);
or U5695 (N_5695,N_2275,N_4107);
or U5696 (N_5696,N_4464,N_4411);
nor U5697 (N_5697,N_3707,N_4668);
nand U5698 (N_5698,N_2489,N_2400);
and U5699 (N_5699,N_3152,N_1282);
and U5700 (N_5700,N_4474,N_4417);
and U5701 (N_5701,N_1342,N_2336);
nand U5702 (N_5702,N_3676,N_4641);
nand U5703 (N_5703,N_175,N_1547);
and U5704 (N_5704,N_2550,N_2750);
or U5705 (N_5705,N_3110,N_604);
nor U5706 (N_5706,N_115,N_3796);
or U5707 (N_5707,N_2525,N_2615);
nand U5708 (N_5708,N_161,N_2320);
nor U5709 (N_5709,N_4854,N_2538);
nand U5710 (N_5710,N_1633,N_1450);
nand U5711 (N_5711,N_2651,N_3811);
xor U5712 (N_5712,N_3637,N_172);
nor U5713 (N_5713,N_4262,N_4228);
nor U5714 (N_5714,N_3175,N_1145);
nor U5715 (N_5715,N_4527,N_1679);
and U5716 (N_5716,N_1084,N_4067);
and U5717 (N_5717,N_4999,N_20);
and U5718 (N_5718,N_3202,N_2847);
nand U5719 (N_5719,N_3639,N_2572);
or U5720 (N_5720,N_557,N_2172);
nand U5721 (N_5721,N_3536,N_763);
xor U5722 (N_5722,N_2463,N_593);
xnor U5723 (N_5723,N_3453,N_795);
nor U5724 (N_5724,N_2920,N_3449);
and U5725 (N_5725,N_4053,N_1126);
nand U5726 (N_5726,N_1996,N_2870);
nor U5727 (N_5727,N_1774,N_1948);
and U5728 (N_5728,N_3340,N_1849);
nor U5729 (N_5729,N_251,N_4385);
or U5730 (N_5730,N_1791,N_102);
nand U5731 (N_5731,N_3903,N_466);
xnor U5732 (N_5732,N_106,N_4101);
and U5733 (N_5733,N_3146,N_770);
and U5734 (N_5734,N_985,N_712);
and U5735 (N_5735,N_785,N_3252);
nand U5736 (N_5736,N_4737,N_660);
nand U5737 (N_5737,N_1135,N_1280);
and U5738 (N_5738,N_531,N_2085);
nor U5739 (N_5739,N_3489,N_601);
or U5740 (N_5740,N_159,N_4848);
nand U5741 (N_5741,N_3598,N_898);
and U5742 (N_5742,N_4715,N_2515);
or U5743 (N_5743,N_2081,N_537);
or U5744 (N_5744,N_1924,N_522);
nor U5745 (N_5745,N_1786,N_2160);
and U5746 (N_5746,N_1301,N_1469);
or U5747 (N_5747,N_2741,N_919);
and U5748 (N_5748,N_4289,N_4352);
or U5749 (N_5749,N_966,N_4521);
or U5750 (N_5750,N_1036,N_739);
nand U5751 (N_5751,N_62,N_4072);
or U5752 (N_5752,N_4171,N_691);
and U5753 (N_5753,N_4887,N_1809);
nor U5754 (N_5754,N_4347,N_3812);
nand U5755 (N_5755,N_2154,N_4567);
or U5756 (N_5756,N_1881,N_849);
nand U5757 (N_5757,N_2684,N_2776);
and U5758 (N_5758,N_2721,N_1934);
nand U5759 (N_5759,N_4030,N_1134);
nand U5760 (N_5760,N_3045,N_2454);
nor U5761 (N_5761,N_3260,N_1765);
xnor U5762 (N_5762,N_4265,N_127);
nand U5763 (N_5763,N_1512,N_1684);
nor U5764 (N_5764,N_206,N_1468);
nand U5765 (N_5765,N_1019,N_345);
nand U5766 (N_5766,N_2148,N_4557);
and U5767 (N_5767,N_529,N_2077);
nor U5768 (N_5768,N_3801,N_2485);
and U5769 (N_5769,N_1917,N_2424);
and U5770 (N_5770,N_4565,N_4648);
or U5771 (N_5771,N_1248,N_869);
nand U5772 (N_5772,N_3908,N_3498);
nand U5773 (N_5773,N_4841,N_1810);
or U5774 (N_5774,N_1133,N_468);
nand U5775 (N_5775,N_2144,N_2367);
nand U5776 (N_5776,N_3988,N_186);
nor U5777 (N_5777,N_1295,N_3156);
and U5778 (N_5778,N_1334,N_3459);
or U5779 (N_5779,N_4547,N_877);
or U5780 (N_5780,N_796,N_2072);
and U5781 (N_5781,N_1579,N_4261);
nand U5782 (N_5782,N_3322,N_3553);
or U5783 (N_5783,N_213,N_4858);
or U5784 (N_5784,N_1995,N_1267);
nand U5785 (N_5785,N_4018,N_641);
nand U5786 (N_5786,N_1402,N_388);
nand U5787 (N_5787,N_3610,N_4244);
and U5788 (N_5788,N_4163,N_4985);
xor U5789 (N_5789,N_1064,N_3056);
nor U5790 (N_5790,N_1734,N_411);
or U5791 (N_5791,N_821,N_4192);
nor U5792 (N_5792,N_4930,N_3047);
and U5793 (N_5793,N_1086,N_56);
or U5794 (N_5794,N_1976,N_1852);
xnor U5795 (N_5795,N_402,N_3622);
or U5796 (N_5796,N_4063,N_933);
nand U5797 (N_5797,N_1884,N_2830);
and U5798 (N_5798,N_4803,N_1732);
nor U5799 (N_5799,N_4315,N_1877);
and U5800 (N_5800,N_2543,N_1099);
nand U5801 (N_5801,N_2197,N_1799);
or U5802 (N_5802,N_3669,N_2051);
or U5803 (N_5803,N_1182,N_2013);
nand U5804 (N_5804,N_1530,N_1194);
or U5805 (N_5805,N_1067,N_1275);
nor U5806 (N_5806,N_2849,N_2299);
nor U5807 (N_5807,N_3181,N_1686);
and U5808 (N_5808,N_4136,N_3554);
and U5809 (N_5809,N_1523,N_546);
and U5810 (N_5810,N_3066,N_2961);
nor U5811 (N_5811,N_3624,N_1186);
nor U5812 (N_5812,N_2833,N_2576);
nor U5813 (N_5813,N_2110,N_1600);
nand U5814 (N_5814,N_3039,N_2565);
and U5815 (N_5815,N_1738,N_3434);
nand U5816 (N_5816,N_4811,N_1047);
nand U5817 (N_5817,N_4866,N_3527);
and U5818 (N_5818,N_3480,N_1000);
nand U5819 (N_5819,N_3331,N_1589);
nand U5820 (N_5820,N_511,N_2063);
nor U5821 (N_5821,N_2868,N_3135);
xor U5822 (N_5822,N_2274,N_4538);
nand U5823 (N_5823,N_3488,N_3404);
nor U5824 (N_5824,N_3342,N_2430);
nand U5825 (N_5825,N_3346,N_2344);
nor U5826 (N_5826,N_258,N_3127);
or U5827 (N_5827,N_2374,N_4745);
or U5828 (N_5828,N_3785,N_3079);
nand U5829 (N_5829,N_1028,N_4777);
and U5830 (N_5830,N_124,N_3732);
and U5831 (N_5831,N_1495,N_1708);
and U5832 (N_5832,N_4001,N_1077);
and U5833 (N_5833,N_4693,N_1693);
and U5834 (N_5834,N_2073,N_4194);
and U5835 (N_5835,N_736,N_2514);
or U5836 (N_5836,N_2654,N_3456);
nor U5837 (N_5837,N_2963,N_1888);
and U5838 (N_5838,N_3318,N_4766);
nand U5839 (N_5839,N_4052,N_1379);
or U5840 (N_5840,N_3189,N_4003);
or U5841 (N_5841,N_1150,N_847);
nor U5842 (N_5842,N_2714,N_3216);
nand U5843 (N_5843,N_4333,N_3034);
nand U5844 (N_5844,N_24,N_3089);
and U5845 (N_5845,N_753,N_4353);
and U5846 (N_5846,N_4906,N_1893);
nand U5847 (N_5847,N_3038,N_3905);
and U5848 (N_5848,N_3274,N_1598);
nand U5849 (N_5849,N_3777,N_455);
nor U5850 (N_5850,N_2906,N_1226);
or U5851 (N_5851,N_4179,N_2383);
or U5852 (N_5852,N_1563,N_4459);
or U5853 (N_5853,N_4093,N_3606);
or U5854 (N_5854,N_1173,N_2417);
nand U5855 (N_5855,N_3846,N_495);
xnor U5856 (N_5856,N_1768,N_1591);
and U5857 (N_5857,N_677,N_4254);
nand U5858 (N_5858,N_2730,N_3731);
nor U5859 (N_5859,N_4905,N_200);
or U5860 (N_5860,N_148,N_1892);
xnor U5861 (N_5861,N_2530,N_872);
nand U5862 (N_5862,N_3636,N_4942);
nand U5863 (N_5863,N_1741,N_4711);
nand U5864 (N_5864,N_1180,N_1376);
nand U5865 (N_5865,N_3286,N_4515);
nor U5866 (N_5866,N_3028,N_1510);
or U5867 (N_5867,N_180,N_328);
or U5868 (N_5868,N_494,N_526);
or U5869 (N_5869,N_4247,N_3704);
or U5870 (N_5870,N_881,N_1798);
and U5871 (N_5871,N_3321,N_1397);
and U5872 (N_5872,N_3968,N_2582);
nand U5873 (N_5873,N_2298,N_2807);
nand U5874 (N_5874,N_4762,N_2214);
nand U5875 (N_5875,N_4444,N_4332);
and U5876 (N_5876,N_3344,N_1992);
and U5877 (N_5877,N_4522,N_3263);
nor U5878 (N_5878,N_451,N_4530);
nor U5879 (N_5879,N_1862,N_1965);
and U5880 (N_5880,N_790,N_3741);
nand U5881 (N_5881,N_4605,N_2517);
and U5882 (N_5882,N_1574,N_2155);
nor U5883 (N_5883,N_3443,N_4435);
nand U5884 (N_5884,N_82,N_2925);
nor U5885 (N_5885,N_2321,N_3967);
and U5886 (N_5886,N_1642,N_4797);
or U5887 (N_5887,N_4922,N_2736);
and U5888 (N_5888,N_93,N_4504);
and U5889 (N_5889,N_4400,N_3114);
or U5890 (N_5890,N_4843,N_563);
or U5891 (N_5891,N_3076,N_3061);
and U5892 (N_5892,N_2254,N_2923);
and U5893 (N_5893,N_4469,N_316);
nor U5894 (N_5894,N_3501,N_4452);
and U5895 (N_5895,N_4172,N_1968);
and U5896 (N_5896,N_3379,N_939);
nand U5897 (N_5897,N_1817,N_289);
and U5898 (N_5898,N_1762,N_952);
and U5899 (N_5899,N_4914,N_4119);
nor U5900 (N_5900,N_3264,N_3966);
nand U5901 (N_5901,N_3888,N_748);
and U5902 (N_5902,N_3978,N_520);
nand U5903 (N_5903,N_2497,N_3584);
nor U5904 (N_5904,N_394,N_212);
nor U5905 (N_5905,N_90,N_4193);
or U5906 (N_5906,N_1615,N_1747);
and U5907 (N_5907,N_2244,N_3645);
or U5908 (N_5908,N_1566,N_4572);
or U5909 (N_5909,N_2671,N_4305);
nor U5910 (N_5910,N_3071,N_2575);
or U5911 (N_5911,N_144,N_838);
nor U5912 (N_5912,N_2239,N_332);
or U5913 (N_5913,N_3653,N_1717);
or U5914 (N_5914,N_60,N_3339);
nor U5915 (N_5915,N_1304,N_4948);
nor U5916 (N_5916,N_2126,N_586);
and U5917 (N_5917,N_1440,N_1216);
or U5918 (N_5918,N_2887,N_2702);
or U5919 (N_5919,N_4291,N_4819);
nor U5920 (N_5920,N_4659,N_1701);
or U5921 (N_5921,N_2952,N_590);
nand U5922 (N_5922,N_3576,N_2903);
and U5923 (N_5923,N_1524,N_1608);
or U5924 (N_5924,N_4348,N_2709);
or U5925 (N_5925,N_4776,N_3356);
nor U5926 (N_5926,N_2698,N_3918);
nand U5927 (N_5927,N_4894,N_4199);
nor U5928 (N_5928,N_3116,N_2604);
nand U5929 (N_5929,N_2435,N_343);
and U5930 (N_5930,N_2534,N_2824);
nor U5931 (N_5931,N_4847,N_3623);
nor U5932 (N_5932,N_1053,N_2679);
or U5933 (N_5933,N_1599,N_4759);
nand U5934 (N_5934,N_2997,N_414);
and U5935 (N_5935,N_2134,N_1796);
nor U5936 (N_5936,N_467,N_1874);
nand U5937 (N_5937,N_1287,N_2065);
nor U5938 (N_5938,N_3324,N_4962);
nand U5939 (N_5939,N_440,N_2725);
and U5940 (N_5940,N_3308,N_26);
nor U5941 (N_5941,N_4513,N_1253);
nand U5942 (N_5942,N_1362,N_2546);
or U5943 (N_5943,N_1492,N_4893);
nor U5944 (N_5944,N_4564,N_2877);
nand U5945 (N_5945,N_2265,N_2895);
or U5946 (N_5946,N_642,N_883);
or U5947 (N_5947,N_2520,N_1617);
nor U5948 (N_5948,N_3627,N_4740);
nor U5949 (N_5949,N_4407,N_1998);
or U5950 (N_5950,N_3894,N_902);
or U5951 (N_5951,N_762,N_1394);
or U5952 (N_5952,N_2034,N_450);
and U5953 (N_5953,N_1235,N_2591);
nand U5954 (N_5954,N_3820,N_475);
nand U5955 (N_5955,N_3772,N_4782);
xnor U5956 (N_5956,N_655,N_4660);
or U5957 (N_5957,N_1011,N_4753);
or U5958 (N_5958,N_3267,N_1427);
nor U5959 (N_5959,N_1183,N_3194);
xnor U5960 (N_5960,N_4749,N_2280);
or U5961 (N_5961,N_2931,N_3422);
and U5962 (N_5962,N_3326,N_4680);
or U5963 (N_5963,N_2398,N_3007);
or U5964 (N_5964,N_4695,N_759);
or U5965 (N_5965,N_1537,N_2464);
nand U5966 (N_5966,N_778,N_3245);
and U5967 (N_5967,N_2157,N_4479);
or U5968 (N_5968,N_2855,N_382);
nor U5969 (N_5969,N_4765,N_4829);
or U5970 (N_5970,N_4442,N_4569);
or U5971 (N_5971,N_977,N_2111);
and U5972 (N_5972,N_4473,N_743);
or U5973 (N_5973,N_2033,N_4580);
nand U5974 (N_5974,N_2364,N_4253);
nor U5975 (N_5975,N_4153,N_4090);
nor U5976 (N_5976,N_2496,N_1560);
nand U5977 (N_5977,N_2382,N_3010);
or U5978 (N_5978,N_1330,N_4368);
or U5979 (N_5979,N_768,N_2541);
and U5980 (N_5980,N_48,N_3641);
nor U5981 (N_5981,N_726,N_280);
and U5982 (N_5982,N_2927,N_4004);
nand U5983 (N_5983,N_1797,N_857);
and U5984 (N_5984,N_2744,N_417);
nand U5985 (N_5985,N_2536,N_2798);
nor U5986 (N_5986,N_4650,N_2003);
nor U5987 (N_5987,N_1034,N_1172);
nand U5988 (N_5988,N_904,N_4405);
nand U5989 (N_5989,N_2938,N_1567);
and U5990 (N_5990,N_3235,N_4276);
and U5991 (N_5991,N_756,N_3662);
nor U5992 (N_5992,N_4635,N_2161);
and U5993 (N_5993,N_168,N_3521);
nand U5994 (N_5994,N_3902,N_2241);
nand U5995 (N_5995,N_3382,N_4314);
nor U5996 (N_5996,N_4164,N_2213);
and U5997 (N_5997,N_3250,N_1665);
nor U5998 (N_5998,N_4774,N_1602);
nand U5999 (N_5999,N_4263,N_4637);
nor U6000 (N_6000,N_3136,N_188);
nand U6001 (N_6001,N_2153,N_2650);
or U6002 (N_6002,N_4339,N_2542);
nand U6003 (N_6003,N_480,N_989);
or U6004 (N_6004,N_2014,N_3889);
or U6005 (N_6005,N_1804,N_540);
nor U6006 (N_6006,N_3471,N_4690);
and U6007 (N_6007,N_4113,N_1794);
or U6008 (N_6008,N_723,N_3904);
or U6009 (N_6009,N_3025,N_499);
and U6010 (N_6010,N_78,N_398);
nand U6011 (N_6011,N_1514,N_4801);
xnor U6012 (N_6012,N_2432,N_4613);
nand U6013 (N_6013,N_1447,N_618);
and U6014 (N_6014,N_1041,N_6);
and U6015 (N_6015,N_4089,N_4984);
nand U6016 (N_6016,N_729,N_1458);
and U6017 (N_6017,N_930,N_3447);
or U6018 (N_6018,N_2930,N_1063);
nand U6019 (N_6019,N_3509,N_4976);
nand U6020 (N_6020,N_167,N_3407);
nand U6021 (N_6021,N_1758,N_1801);
nand U6022 (N_6022,N_1870,N_2602);
and U6023 (N_6023,N_3143,N_683);
nor U6024 (N_6024,N_407,N_2814);
or U6025 (N_6025,N_1785,N_1993);
and U6026 (N_6026,N_1191,N_3257);
and U6027 (N_6027,N_1739,N_2048);
nor U6028 (N_6028,N_4585,N_1842);
and U6029 (N_6029,N_3871,N_3655);
nand U6030 (N_6030,N_4006,N_457);
xor U6031 (N_6031,N_1151,N_2594);
or U6032 (N_6032,N_2600,N_3460);
or U6033 (N_6033,N_1878,N_4054);
or U6034 (N_6034,N_4594,N_252);
or U6035 (N_6035,N_932,N_3703);
or U6036 (N_6036,N_3705,N_3601);
nand U6037 (N_6037,N_3233,N_4294);
or U6038 (N_6038,N_1914,N_3974);
or U6039 (N_6039,N_408,N_4237);
or U6040 (N_6040,N_3552,N_300);
nand U6041 (N_6041,N_2004,N_3765);
and U6042 (N_6042,N_3222,N_3580);
and U6043 (N_6043,N_868,N_4116);
and U6044 (N_6044,N_2386,N_273);
or U6045 (N_6045,N_3165,N_4123);
nor U6046 (N_6046,N_4242,N_3524);
or U6047 (N_6047,N_3952,N_4997);
xor U6048 (N_6048,N_7,N_2809);
nor U6049 (N_6049,N_3442,N_1596);
nand U6050 (N_6050,N_650,N_2509);
or U6051 (N_6051,N_3718,N_2223);
nand U6052 (N_6052,N_2629,N_954);
nand U6053 (N_6053,N_3663,N_1222);
or U6054 (N_6054,N_1269,N_2179);
nand U6055 (N_6055,N_1264,N_3539);
or U6056 (N_6056,N_4157,N_89);
and U6057 (N_6057,N_4617,N_3742);
nor U6058 (N_6058,N_183,N_928);
or U6059 (N_6059,N_2132,N_4987);
or U6060 (N_6060,N_3755,N_4106);
nand U6061 (N_6061,N_3794,N_4852);
nor U6062 (N_6062,N_4309,N_1153);
nor U6063 (N_6063,N_3052,N_210);
and U6064 (N_6064,N_724,N_4895);
and U6065 (N_6065,N_1097,N_1046);
or U6066 (N_6066,N_1490,N_2245);
or U6067 (N_6067,N_690,N_4252);
or U6068 (N_6068,N_2024,N_3120);
xnor U6069 (N_6069,N_4832,N_1098);
or U6070 (N_6070,N_3868,N_852);
or U6071 (N_6071,N_2074,N_153);
xnor U6072 (N_6072,N_3162,N_3547);
nor U6073 (N_6073,N_2688,N_700);
and U6074 (N_6074,N_3508,N_3874);
nor U6075 (N_6075,N_834,N_2401);
or U6076 (N_6076,N_570,N_4958);
and U6077 (N_6077,N_738,N_4586);
and U6078 (N_6078,N_4046,N_1925);
and U6079 (N_6079,N_648,N_2916);
nor U6080 (N_6080,N_704,N_752);
nand U6081 (N_6081,N_1604,N_2162);
nor U6082 (N_6082,N_3173,N_3417);
nand U6083 (N_6083,N_3205,N_2039);
nand U6084 (N_6084,N_4842,N_2636);
or U6085 (N_6085,N_3992,N_3323);
or U6086 (N_6086,N_3465,N_2170);
nand U6087 (N_6087,N_2646,N_2735);
or U6088 (N_6088,N_2106,N_209);
and U6089 (N_6089,N_116,N_1923);
or U6090 (N_6090,N_1308,N_1307);
nand U6091 (N_6091,N_2378,N_1388);
nand U6092 (N_6092,N_1266,N_1906);
or U6093 (N_6093,N_1539,N_3074);
and U6094 (N_6094,N_3824,N_3537);
xor U6095 (N_6095,N_1094,N_1984);
nor U6096 (N_6096,N_1207,N_774);
nand U6097 (N_6097,N_197,N_3273);
or U6098 (N_6098,N_749,N_2041);
and U6099 (N_6099,N_4525,N_3198);
and U6100 (N_6100,N_4658,N_1156);
and U6101 (N_6101,N_4857,N_416);
or U6102 (N_6102,N_3469,N_2780);
nor U6103 (N_6103,N_1104,N_4102);
nor U6104 (N_6104,N_2329,N_2362);
nand U6105 (N_6105,N_2302,N_4608);
and U6106 (N_6106,N_140,N_944);
nand U6107 (N_6107,N_4897,N_1412);
or U6108 (N_6108,N_1154,N_2529);
and U6109 (N_6109,N_3004,N_333);
nand U6110 (N_6110,N_1974,N_4441);
nor U6111 (N_6111,N_2549,N_2187);
nor U6112 (N_6112,N_4429,N_4364);
or U6113 (N_6113,N_2555,N_2760);
or U6114 (N_6114,N_4097,N_3795);
xnor U6115 (N_6115,N_2505,N_1978);
and U6116 (N_6116,N_559,N_1525);
nor U6117 (N_6117,N_314,N_9);
xor U6118 (N_6118,N_4446,N_2843);
nor U6119 (N_6119,N_1211,N_3950);
nand U6120 (N_6120,N_830,N_1926);
and U6121 (N_6121,N_4099,N_1813);
nand U6122 (N_6122,N_980,N_77);
nand U6123 (N_6123,N_3728,N_2605);
nand U6124 (N_6124,N_3931,N_4542);
or U6125 (N_6125,N_4128,N_595);
nor U6126 (N_6126,N_2945,N_1903);
nor U6127 (N_6127,N_2445,N_233);
and U6128 (N_6128,N_551,N_313);
and U6129 (N_6129,N_3020,N_2552);
or U6130 (N_6130,N_222,N_3105);
nor U6131 (N_6131,N_1535,N_3126);
or U6132 (N_6132,N_2573,N_2819);
nand U6133 (N_6133,N_1466,N_596);
and U6134 (N_6134,N_1840,N_4458);
nor U6135 (N_6135,N_3370,N_4810);
or U6136 (N_6136,N_675,N_853);
nor U6137 (N_6137,N_2229,N_4404);
and U6138 (N_6138,N_825,N_3494);
and U6139 (N_6139,N_2828,N_4964);
nor U6140 (N_6140,N_426,N_4714);
or U6141 (N_6141,N_1371,N_1667);
and U6142 (N_6142,N_2422,N_4998);
nor U6143 (N_6143,N_1027,N_4239);
nand U6144 (N_6144,N_2774,N_1703);
nor U6145 (N_6145,N_1373,N_547);
and U6146 (N_6146,N_4823,N_2330);
or U6147 (N_6147,N_2152,N_4165);
nand U6148 (N_6148,N_3986,N_3666);
nand U6149 (N_6149,N_4073,N_4639);
or U6150 (N_6150,N_2189,N_3285);
nand U6151 (N_6151,N_4972,N_865);
or U6152 (N_6152,N_854,N_2335);
nand U6153 (N_6153,N_1165,N_2218);
nand U6154 (N_6154,N_4028,N_425);
nand U6155 (N_6155,N_1230,N_2586);
nor U6156 (N_6156,N_542,N_1176);
or U6157 (N_6157,N_1652,N_4688);
and U6158 (N_6158,N_2084,N_4647);
or U6159 (N_6159,N_1856,N_1737);
or U6160 (N_6160,N_2975,N_4634);
and U6161 (N_6161,N_4566,N_1626);
and U6162 (N_6162,N_3083,N_4114);
or U6163 (N_6163,N_2112,N_1206);
and U6164 (N_6164,N_2669,N_3565);
xnor U6165 (N_6165,N_1837,N_1309);
and U6166 (N_6166,N_1223,N_727);
nor U6167 (N_6167,N_2673,N_4656);
and U6168 (N_6168,N_4927,N_1558);
and U6169 (N_6169,N_107,N_83);
and U6170 (N_6170,N_3412,N_192);
nand U6171 (N_6171,N_3710,N_31);
or U6172 (N_6172,N_393,N_3084);
or U6173 (N_6173,N_1073,N_1335);
nor U6174 (N_6174,N_4100,N_3424);
xor U6175 (N_6175,N_2053,N_3377);
and U6176 (N_6176,N_3916,N_1610);
and U6177 (N_6177,N_1404,N_2164);
nor U6178 (N_6178,N_2763,N_2632);
and U6179 (N_6179,N_4978,N_33);
nor U6180 (N_6180,N_2009,N_1975);
or U6181 (N_6181,N_1175,N_4366);
nor U6182 (N_6182,N_4034,N_3067);
nand U6183 (N_6183,N_3048,N_73);
or U6184 (N_6184,N_1502,N_4214);
nand U6185 (N_6185,N_371,N_1127);
or U6186 (N_6186,N_472,N_1613);
nor U6187 (N_6187,N_3760,N_3787);
or U6188 (N_6188,N_589,N_4208);
or U6189 (N_6189,N_3041,N_1093);
or U6190 (N_6190,N_1238,N_4578);
or U6191 (N_6191,N_2066,N_481);
nand U6192 (N_6192,N_3131,N_2700);
and U6193 (N_6193,N_304,N_1634);
nor U6194 (N_6194,N_4717,N_2457);
nand U6195 (N_6195,N_1092,N_1787);
nor U6196 (N_6196,N_681,N_4794);
and U6197 (N_6197,N_4463,N_4277);
nor U6198 (N_6198,N_1518,N_3635);
nor U6199 (N_6199,N_4095,N_662);
nor U6200 (N_6200,N_157,N_52);
nor U6201 (N_6201,N_220,N_935);
and U6202 (N_6202,N_2437,N_4198);
or U6203 (N_6203,N_4802,N_1811);
nand U6204 (N_6204,N_1905,N_544);
xnor U6205 (N_6205,N_568,N_2779);
nor U6206 (N_6206,N_248,N_4177);
nand U6207 (N_6207,N_4,N_765);
and U6208 (N_6208,N_1625,N_2451);
or U6209 (N_6209,N_179,N_1117);
nand U6210 (N_6210,N_3093,N_1118);
nor U6211 (N_6211,N_3333,N_386);
and U6212 (N_6212,N_3611,N_802);
nand U6213 (N_6213,N_1681,N_4837);
nor U6214 (N_6214,N_3976,N_4915);
or U6215 (N_6215,N_340,N_2147);
nand U6216 (N_6216,N_1325,N_2914);
and U6217 (N_6217,N_808,N_3080);
nand U6218 (N_6218,N_2557,N_3158);
or U6219 (N_6219,N_4236,N_2969);
nand U6220 (N_6220,N_4336,N_3725);
or U6221 (N_6221,N_438,N_1782);
or U6222 (N_6222,N_1372,N_1622);
nor U6223 (N_6223,N_3797,N_4959);
nand U6224 (N_6224,N_2589,N_1091);
or U6225 (N_6225,N_3278,N_484);
nor U6226 (N_6226,N_315,N_3336);
or U6227 (N_6227,N_3981,N_1421);
and U6228 (N_6228,N_2238,N_342);
or U6229 (N_6229,N_3543,N_4185);
and U6230 (N_6230,N_893,N_2995);
nand U6231 (N_6231,N_1100,N_4853);
nor U6232 (N_6232,N_4176,N_2532);
nor U6233 (N_6233,N_2559,N_2307);
and U6234 (N_6234,N_1839,N_4596);
and U6235 (N_6235,N_4950,N_2177);
and U6236 (N_6236,N_2738,N_2442);
nand U6237 (N_6237,N_1972,N_351);
xnor U6238 (N_6238,N_3347,N_719);
nand U6239 (N_6239,N_3697,N_1025);
nor U6240 (N_6240,N_4755,N_2377);
nor U6241 (N_6241,N_1879,N_1261);
xnor U6242 (N_6242,N_4449,N_982);
or U6243 (N_6243,N_1311,N_2861);
nand U6244 (N_6244,N_1409,N_1247);
or U6245 (N_6245,N_2128,N_4319);
and U6246 (N_6246,N_1958,N_483);
or U6247 (N_6247,N_2453,N_4620);
nor U6248 (N_6248,N_3680,N_885);
nor U6249 (N_6249,N_4562,N_2093);
nand U6250 (N_6250,N_2500,N_1382);
nor U6251 (N_6251,N_3690,N_4969);
xor U6252 (N_6252,N_2740,N_4633);
nor U6253 (N_6253,N_4662,N_1472);
nand U6254 (N_6254,N_4773,N_536);
nand U6255 (N_6255,N_4968,N_1326);
nor U6256 (N_6256,N_3829,N_1828);
and U6257 (N_6257,N_4492,N_1406);
and U6258 (N_6258,N_2232,N_4112);
or U6259 (N_6259,N_4700,N_3186);
and U6260 (N_6260,N_3029,N_629);
and U6261 (N_6261,N_4625,N_2874);
nor U6262 (N_6262,N_2038,N_929);
and U6263 (N_6263,N_2942,N_4903);
or U6264 (N_6264,N_3296,N_4065);
nand U6265 (N_6265,N_2202,N_3512);
nor U6266 (N_6266,N_3490,N_2011);
nand U6267 (N_6267,N_2231,N_1744);
nor U6268 (N_6268,N_4581,N_1970);
nand U6269 (N_6269,N_227,N_3293);
nor U6270 (N_6270,N_4110,N_2999);
xnor U6271 (N_6271,N_2210,N_1434);
nor U6272 (N_6272,N_4699,N_917);
nand U6273 (N_6273,N_575,N_2334);
and U6274 (N_6274,N_1664,N_2662);
nand U6275 (N_6275,N_689,N_2704);
nor U6276 (N_6276,N_3090,N_2976);
and U6277 (N_6277,N_4491,N_1876);
nor U6278 (N_6278,N_2872,N_1896);
or U6279 (N_6279,N_335,N_1638);
and U6280 (N_6280,N_3141,N_4000);
nor U6281 (N_6281,N_4108,N_3695);
nor U6282 (N_6282,N_3448,N_2032);
nand U6283 (N_6283,N_2404,N_3177);
nand U6284 (N_6284,N_401,N_1710);
nand U6285 (N_6285,N_3764,N_4245);
nand U6286 (N_6286,N_2316,N_4007);
and U6287 (N_6287,N_290,N_1116);
nand U6288 (N_6288,N_988,N_4337);
nor U6289 (N_6289,N_3802,N_2964);
or U6290 (N_6290,N_1715,N_353);
nor U6291 (N_6291,N_1499,N_1904);
nor U6292 (N_6292,N_86,N_104);
or U6293 (N_6293,N_1204,N_4317);
or U6294 (N_6294,N_4955,N_2805);
or U6295 (N_6295,N_1556,N_1743);
nor U6296 (N_6296,N_1779,N_3656);
nand U6297 (N_6297,N_2138,N_2356);
and U6298 (N_6298,N_514,N_1937);
and U6299 (N_6299,N_3885,N_421);
nand U6300 (N_6300,N_3917,N_3818);
and U6301 (N_6301,N_621,N_936);
nor U6302 (N_6302,N_3800,N_4880);
and U6303 (N_6303,N_308,N_1515);
and U6304 (N_6304,N_4873,N_3212);
nor U6305 (N_6305,N_99,N_1844);
and U6306 (N_6306,N_320,N_1706);
nand U6307 (N_6307,N_372,N_1620);
nand U6308 (N_6308,N_3566,N_4507);
nor U6309 (N_6309,N_1102,N_2139);
nand U6310 (N_6310,N_355,N_895);
nor U6311 (N_6311,N_1364,N_2191);
and U6312 (N_6312,N_4258,N_4851);
and U6313 (N_6313,N_4345,N_1899);
or U6314 (N_6314,N_3228,N_3994);
or U6315 (N_6315,N_4805,N_3569);
and U6316 (N_6316,N_3288,N_4508);
xor U6317 (N_6317,N_3838,N_4746);
or U6318 (N_6318,N_3174,N_978);
nand U6319 (N_6319,N_1601,N_3139);
nor U6320 (N_6320,N_3842,N_4402);
or U6321 (N_6321,N_3023,N_3688);
nand U6322 (N_6322,N_564,N_1867);
nand U6323 (N_6323,N_1534,N_2371);
nor U6324 (N_6324,N_656,N_4809);
and U6325 (N_6325,N_3261,N_4014);
or U6326 (N_6326,N_4269,N_725);
and U6327 (N_6327,N_3534,N_541);
and U6328 (N_6328,N_637,N_2255);
or U6329 (N_6329,N_2450,N_4240);
nand U6330 (N_6330,N_3452,N_4718);
nor U6331 (N_6331,N_906,N_968);
and U6332 (N_6332,N_2842,N_1653);
or U6333 (N_6333,N_665,N_3530);
xnor U6334 (N_6334,N_1595,N_3616);
and U6335 (N_6335,N_1775,N_970);
or U6336 (N_6336,N_3484,N_1017);
and U6337 (N_6337,N_3282,N_3597);
or U6338 (N_6338,N_862,N_122);
and U6339 (N_6339,N_2465,N_2553);
or U6340 (N_6340,N_447,N_3343);
xor U6341 (N_6341,N_3241,N_2617);
or U6342 (N_6342,N_4941,N_134);
nor U6343 (N_6343,N_961,N_2989);
or U6344 (N_6344,N_4812,N_822);
xnor U6345 (N_6345,N_4632,N_3476);
nor U6346 (N_6346,N_4568,N_1339);
or U6347 (N_6347,N_2668,N_1214);
and U6348 (N_6348,N_3495,N_3302);
or U6349 (N_6349,N_2292,N_1483);
or U6350 (N_6350,N_1503,N_4607);
nand U6351 (N_6351,N_4062,N_3238);
nor U6352 (N_6352,N_733,N_2022);
nand U6353 (N_6353,N_4654,N_946);
and U6354 (N_6354,N_4670,N_828);
nor U6355 (N_6355,N_1215,N_2770);
or U6356 (N_6356,N_4033,N_453);
nand U6357 (N_6357,N_2440,N_1451);
nor U6358 (N_6358,N_123,N_69);
nor U6359 (N_6359,N_4083,N_2845);
nand U6360 (N_6360,N_264,N_2907);
nor U6361 (N_6361,N_1448,N_3030);
or U6362 (N_6362,N_3100,N_2049);
nand U6363 (N_6363,N_2360,N_2890);
nand U6364 (N_6364,N_2061,N_4232);
and U6365 (N_6365,N_429,N_909);
or U6366 (N_6366,N_100,N_2278);
or U6367 (N_6367,N_4671,N_751);
and U6368 (N_6368,N_3612,N_1393);
nor U6369 (N_6369,N_3560,N_3832);
and U6370 (N_6370,N_4389,N_3033);
and U6371 (N_6371,N_2758,N_2610);
nand U6372 (N_6372,N_3390,N_3375);
nor U6373 (N_6373,N_2756,N_4529);
or U6374 (N_6374,N_3036,N_1208);
nor U6375 (N_6375,N_3594,N_3353);
nand U6376 (N_6376,N_195,N_354);
nand U6377 (N_6377,N_166,N_611);
and U6378 (N_6378,N_3850,N_2183);
nand U6379 (N_6379,N_2423,N_2655);
or U6380 (N_6380,N_3839,N_2338);
and U6381 (N_6381,N_2396,N_1624);
or U6382 (N_6382,N_2409,N_1212);
nand U6383 (N_6383,N_3301,N_3763);
and U6384 (N_6384,N_1889,N_3500);
and U6385 (N_6385,N_2345,N_2300);
nand U6386 (N_6386,N_1323,N_2181);
or U6387 (N_6387,N_4870,N_1865);
xor U6388 (N_6388,N_3869,N_603);
and U6389 (N_6389,N_3849,N_2644);
or U6390 (N_6390,N_2563,N_2611);
nand U6391 (N_6391,N_2802,N_3481);
and U6392 (N_6392,N_4382,N_4498);
xor U6393 (N_6393,N_2888,N_2363);
and U6394 (N_6394,N_4908,N_2099);
or U6395 (N_6395,N_524,N_47);
and U6396 (N_6396,N_2987,N_4316);
or U6397 (N_6397,N_3541,N_3408);
nor U6398 (N_6398,N_3807,N_4058);
nand U6399 (N_6399,N_4212,N_1149);
nand U6400 (N_6400,N_4534,N_3389);
nand U6401 (N_6401,N_3893,N_4284);
or U6402 (N_6402,N_2613,N_682);
nand U6403 (N_6403,N_3817,N_1707);
nor U6404 (N_6404,N_323,N_4077);
nand U6405 (N_6405,N_349,N_1337);
nand U6406 (N_6406,N_1095,N_3991);
nor U6407 (N_6407,N_4836,N_3788);
or U6408 (N_6408,N_3749,N_4535);
or U6409 (N_6409,N_1050,N_3315);
nor U6410 (N_6410,N_3319,N_4523);
or U6411 (N_6411,N_1894,N_1244);
and U6412 (N_6412,N_2829,N_1473);
and U6413 (N_6413,N_680,N_1631);
nor U6414 (N_6414,N_2108,N_143);
or U6415 (N_6415,N_3031,N_2754);
nor U6416 (N_6416,N_4761,N_3790);
nor U6417 (N_6417,N_4302,N_4076);
nand U6418 (N_6418,N_3727,N_4928);
nor U6419 (N_6419,N_2361,N_4591);
nor U6420 (N_6420,N_3234,N_2587);
nor U6421 (N_6421,N_817,N_2174);
and U6422 (N_6422,N_1583,N_2391);
nand U6423 (N_6423,N_2167,N_3284);
nor U6424 (N_6424,N_4056,N_4323);
and U6425 (N_6425,N_4174,N_298);
or U6426 (N_6426,N_4064,N_363);
or U6427 (N_6427,N_1090,N_4509);
nand U6428 (N_6428,N_1239,N_4979);
nand U6429 (N_6429,N_489,N_4288);
nand U6430 (N_6430,N_4993,N_4724);
nand U6431 (N_6431,N_4661,N_1286);
or U6432 (N_6432,N_1549,N_4790);
nand U6433 (N_6433,N_381,N_2875);
and U6434 (N_6434,N_4166,N_98);
nor U6435 (N_6435,N_1478,N_2166);
xnor U6436 (N_6436,N_1543,N_3144);
and U6437 (N_6437,N_2297,N_41);
or U6438 (N_6438,N_3297,N_4713);
nand U6439 (N_6439,N_4907,N_1864);
or U6440 (N_6440,N_845,N_1627);
nor U6441 (N_6441,N_844,N_4996);
and U6442 (N_6442,N_2224,N_670);
nor U6443 (N_6443,N_1763,N_2151);
or U6444 (N_6444,N_1455,N_2608);
nor U6445 (N_6445,N_3145,N_616);
nor U6446 (N_6446,N_1008,N_2664);
and U6447 (N_6447,N_4891,N_1365);
or U6448 (N_6448,N_3160,N_2230);
nor U6449 (N_6449,N_806,N_3854);
xnor U6450 (N_6450,N_766,N_3999);
nor U6451 (N_6451,N_3793,N_594);
nand U6452 (N_6452,N_1464,N_940);
or U6453 (N_6453,N_84,N_4081);
and U6454 (N_6454,N_1964,N_4428);
xor U6455 (N_6455,N_2983,N_2910);
nand U6456 (N_6456,N_1401,N_4800);
nand U6457 (N_6457,N_4920,N_4275);
or U6458 (N_6458,N_4636,N_565);
and U6459 (N_6459,N_584,N_3215);
nor U6460 (N_6460,N_1136,N_1061);
and U6461 (N_6461,N_4040,N_427);
or U6462 (N_6462,N_4360,N_2064);
xor U6463 (N_6463,N_496,N_2025);
and U6464 (N_6464,N_3276,N_4705);
or U6465 (N_6465,N_3503,N_1554);
or U6466 (N_6466,N_1317,N_1121);
xnor U6467 (N_6467,N_1825,N_3640);
and U6468 (N_6468,N_1812,N_1909);
nor U6469 (N_6469,N_2369,N_1698);
and U6470 (N_6470,N_4574,N_2913);
nand U6471 (N_6471,N_503,N_2201);
or U6472 (N_6472,N_4126,N_68);
and U6473 (N_6473,N_713,N_326);
nand U6474 (N_6474,N_1355,N_3063);
nand U6475 (N_6475,N_1137,N_1623);
or U6476 (N_6476,N_2666,N_2225);
or U6477 (N_6477,N_2313,N_3287);
or U6478 (N_6478,N_4380,N_5);
nor U6479 (N_6479,N_819,N_2129);
or U6480 (N_6480,N_3670,N_578);
nor U6481 (N_6481,N_3087,N_4532);
or U6482 (N_6482,N_4619,N_1188);
nand U6483 (N_6483,N_2570,N_346);
nor U6484 (N_6484,N_2722,N_3659);
and U6485 (N_6485,N_1109,N_1588);
nand U6486 (N_6486,N_23,N_4963);
nor U6487 (N_6487,N_3022,N_3119);
nand U6488 (N_6488,N_1249,N_249);
or U6489 (N_6489,N_1954,N_4413);
nand U6490 (N_6490,N_4679,N_2524);
or U6491 (N_6491,N_4579,N_2408);
nand U6492 (N_6492,N_4197,N_1346);
xnor U6493 (N_6493,N_479,N_4234);
nor U6494 (N_6494,N_2574,N_2957);
and U6495 (N_6495,N_1303,N_3224);
nand U6496 (N_6496,N_2727,N_4560);
or U6497 (N_6497,N_4386,N_2094);
and U6498 (N_6498,N_3937,N_3574);
nand U6499 (N_6499,N_798,N_2653);
or U6500 (N_6500,N_549,N_1641);
nor U6501 (N_6501,N_1695,N_3529);
nand U6502 (N_6502,N_4503,N_3316);
nand U6503 (N_6503,N_2277,N_4296);
nor U6504 (N_6504,N_543,N_3929);
nor U6505 (N_6505,N_649,N_2510);
or U6506 (N_6506,N_259,N_2637);
nor U6507 (N_6507,N_4146,N_3096);
nand U6508 (N_6508,N_1396,N_34);
or U6509 (N_6509,N_1315,N_722);
nand U6510 (N_6510,N_4932,N_3477);
nand U6511 (N_6511,N_3775,N_471);
nor U6512 (N_6512,N_2062,N_158);
or U6513 (N_6513,N_4416,N_4885);
nor U6514 (N_6514,N_731,N_4938);
nor U6515 (N_6515,N_3702,N_4470);
and U6516 (N_6516,N_841,N_2260);
and U6517 (N_6517,N_4983,N_3470);
nand U6518 (N_6518,N_3638,N_3357);
nand U6519 (N_6519,N_4685,N_773);
and U6520 (N_6520,N_3505,N_3383);
nor U6521 (N_6521,N_3866,N_2343);
nor U6522 (N_6522,N_1350,N_22);
nand U6523 (N_6523,N_1869,N_996);
nand U6524 (N_6524,N_2010,N_4060);
or U6525 (N_6525,N_4665,N_3099);
or U6526 (N_6526,N_855,N_4086);
or U6527 (N_6527,N_4012,N_831);
nor U6528 (N_6528,N_3643,N_3159);
and U6529 (N_6529,N_2708,N_135);
and U6530 (N_6530,N_4838,N_4142);
nor U6531 (N_6531,N_1575,N_717);
or U6532 (N_6532,N_938,N_3928);
nand U6533 (N_6533,N_1426,N_3006);
nor U6534 (N_6534,N_4281,N_837);
or U6535 (N_6535,N_1456,N_4306);
or U6536 (N_6536,N_4454,N_2821);
and U6537 (N_6537,N_4167,N_2027);
nor U6538 (N_6538,N_3124,N_3332);
and U6539 (N_6539,N_4973,N_4312);
or U6540 (N_6540,N_4210,N_1166);
and U6541 (N_6541,N_2317,N_2996);
nand U6542 (N_6542,N_2339,N_238);
nand U6543 (N_6543,N_1755,N_4009);
or U6544 (N_6544,N_1504,N_3590);
and U6545 (N_6545,N_2955,N_4595);
nor U6546 (N_6546,N_718,N_3248);
or U6547 (N_6547,N_2269,N_112);
and U6548 (N_6548,N_4526,N_2622);
or U6549 (N_6549,N_3246,N_4953);
or U6550 (N_6550,N_3115,N_3752);
or U6551 (N_6551,N_3726,N_674);
nor U6552 (N_6552,N_1236,N_2493);
or U6553 (N_6553,N_1263,N_120);
and U6554 (N_6554,N_755,N_1022);
nor U6555 (N_6555,N_2645,N_1449);
and U6556 (N_6556,N_2127,N_2936);
nor U6557 (N_6557,N_1221,N_424);
xor U6558 (N_6558,N_3897,N_3360);
and U6559 (N_6559,N_37,N_4771);
nand U6560 (N_6560,N_139,N_647);
or U6561 (N_6561,N_1997,N_125);
or U6562 (N_6562,N_1967,N_920);
nor U6563 (N_6563,N_2764,N_1370);
and U6564 (N_6564,N_612,N_1383);
nand U6565 (N_6565,N_497,N_2898);
nor U6566 (N_6566,N_1783,N_4150);
nand U6567 (N_6567,N_224,N_4241);
or U6568 (N_6568,N_1661,N_4374);
or U6569 (N_6569,N_3482,N_1380);
nor U6570 (N_6570,N_2902,N_3969);
or U6571 (N_6571,N_2348,N_3808);
or U6572 (N_6572,N_3649,N_3130);
or U6573 (N_6573,N_992,N_3650);
nand U6574 (N_6574,N_229,N_3851);
and U6575 (N_6575,N_1407,N_2468);
nor U6576 (N_6576,N_3251,N_3971);
nor U6577 (N_6577,N_2273,N_728);
and U6578 (N_6578,N_4943,N_4990);
or U6579 (N_6579,N_1928,N_734);
or U6580 (N_6580,N_3402,N_2823);
nand U6581 (N_6581,N_3913,N_2818);
nor U6582 (N_6582,N_1322,N_4381);
and U6583 (N_6583,N_916,N_4609);
nor U6584 (N_6584,N_3708,N_4488);
nor U6585 (N_6585,N_3396,N_4259);
nor U6586 (N_6586,N_3891,N_4871);
or U6587 (N_6587,N_2991,N_2477);
or U6588 (N_6588,N_2113,N_3782);
nor U6589 (N_6589,N_2425,N_1277);
nor U6590 (N_6590,N_3392,N_3863);
or U6591 (N_6591,N_706,N_1318);
nand U6592 (N_6592,N_2080,N_3767);
nand U6593 (N_6593,N_2840,N_2180);
nand U6594 (N_6594,N_4590,N_1147);
nor U6595 (N_6595,N_2249,N_4468);
or U6596 (N_6596,N_3134,N_4519);
and U6597 (N_6597,N_769,N_2752);
nand U6598 (N_6598,N_1784,N_3614);
or U6599 (N_6599,N_2947,N_1669);
or U6600 (N_6600,N_614,N_3208);
nor U6601 (N_6601,N_3166,N_2701);
or U6602 (N_6602,N_3522,N_3711);
xor U6603 (N_6603,N_1629,N_4937);
nand U6604 (N_6604,N_13,N_1861);
nor U6605 (N_6605,N_1605,N_366);
or U6606 (N_6606,N_3784,N_3930);
nor U6607 (N_6607,N_1938,N_4701);
nor U6608 (N_6608,N_3932,N_1678);
nor U6609 (N_6609,N_1446,N_3472);
and U6610 (N_6610,N_413,N_3277);
nand U6611 (N_6611,N_4328,N_3575);
or U6612 (N_6612,N_2703,N_3415);
nand U6613 (N_6613,N_1773,N_4672);
or U6614 (N_6614,N_458,N_910);
and U6615 (N_6615,N_3730,N_2119);
nor U6616 (N_6616,N_3169,N_3486);
nor U6617 (N_6617,N_943,N_2827);
nor U6618 (N_6618,N_3496,N_4290);
nand U6619 (N_6619,N_4189,N_2315);
and U6620 (N_6620,N_2486,N_3862);
or U6621 (N_6621,N_4850,N_3540);
or U6622 (N_6622,N_3055,N_4213);
nand U6623 (N_6623,N_4048,N_44);
or U6624 (N_6624,N_1351,N_2031);
nand U6625 (N_6625,N_2217,N_858);
nor U6626 (N_6626,N_4390,N_2028);
and U6627 (N_6627,N_3201,N_602);
or U6628 (N_6628,N_4554,N_1952);
and U6629 (N_6629,N_150,N_2135);
xor U6630 (N_6630,N_4720,N_4233);
or U6631 (N_6631,N_2782,N_1860);
and U6632 (N_6632,N_3147,N_3780);
and U6633 (N_6633,N_4763,N_3810);
nand U6634 (N_6634,N_312,N_4584);
and U6635 (N_6635,N_498,N_3187);
nand U6636 (N_6636,N_3148,N_1594);
nor U6637 (N_6637,N_3335,N_10);
nand U6638 (N_6638,N_3317,N_2755);
nand U6639 (N_6639,N_2426,N_318);
or U6640 (N_6640,N_4977,N_4421);
and U6641 (N_6641,N_4204,N_4622);
nor U6642 (N_6642,N_2350,N_191);
nor U6643 (N_6643,N_1689,N_2630);
nand U6644 (N_6644,N_4061,N_399);
and U6645 (N_6645,N_199,N_1411);
and U6646 (N_6646,N_3209,N_101);
nand U6647 (N_6647,N_4221,N_461);
or U6648 (N_6648,N_1956,N_1189);
nand U6649 (N_6649,N_3865,N_1994);
nor U6650 (N_6650,N_3358,N_3714);
nand U6651 (N_6651,N_2919,N_2479);
and U6652 (N_6652,N_4865,N_2406);
nand U6653 (N_6653,N_4981,N_3520);
nand U6654 (N_6654,N_4540,N_4949);
nor U6655 (N_6655,N_1299,N_3582);
and U6656 (N_6656,N_4683,N_1112);
or U6657 (N_6657,N_3354,N_1122);
xor U6658 (N_6658,N_2501,N_1932);
nand U6659 (N_6659,N_4485,N_3896);
nor U6660 (N_6660,N_4279,N_4248);
nor U6661 (N_6661,N_1143,N_1432);
and U6662 (N_6662,N_3747,N_2766);
nor U6663 (N_6663,N_3984,N_2474);
nor U6664 (N_6664,N_3128,N_2402);
nor U6665 (N_6665,N_1078,N_1532);
or U6666 (N_6666,N_132,N_2467);
nand U6667 (N_6667,N_742,N_1674);
or U6668 (N_6668,N_3646,N_747);
nor U6669 (N_6669,N_1640,N_3922);
nor U6670 (N_6670,N_1526,N_1327);
or U6671 (N_6671,N_532,N_4511);
or U6672 (N_6672,N_2649,N_4925);
nand U6673 (N_6673,N_3345,N_3154);
or U6674 (N_6674,N_2007,N_3673);
nand U6675 (N_6675,N_685,N_794);
nand U6676 (N_6676,N_4372,N_630);
and U6677 (N_6677,N_814,N_3692);
and U6678 (N_6678,N_3799,N_2288);
or U6679 (N_6679,N_1177,N_811);
and U6680 (N_6680,N_3185,N_3923);
nor U6681 (N_6681,N_3858,N_4787);
nand U6682 (N_6682,N_1982,N_267);
nand U6683 (N_6683,N_1312,N_202);
and U6684 (N_6684,N_4235,N_2256);
xor U6685 (N_6685,N_3397,N_405);
or U6686 (N_6686,N_4649,N_1501);
or U6687 (N_6687,N_2892,N_4598);
or U6688 (N_6688,N_4960,N_4593);
and U6689 (N_6689,N_823,N_4286);
nand U6690 (N_6690,N_2773,N_3681);
or U6691 (N_6691,N_3425,N_631);
nor U6692 (N_6692,N_2578,N_4486);
and U6693 (N_6693,N_2452,N_2403);
and U6694 (N_6694,N_554,N_3062);
nor U6695 (N_6695,N_2020,N_4741);
nor U6696 (N_6696,N_4877,N_4874);
nor U6697 (N_6697,N_396,N_3197);
nand U6698 (N_6698,N_3398,N_1505);
nor U6699 (N_6699,N_193,N_4292);
and U6700 (N_6700,N_3008,N_2800);
or U6701 (N_6701,N_4266,N_1702);
nand U6702 (N_6702,N_1920,N_4021);
and U6703 (N_6703,N_4767,N_3348);
and U6704 (N_6704,N_1319,N_4602);
and U6705 (N_6705,N_3314,N_1572);
or U6706 (N_6706,N_775,N_3514);
and U6707 (N_6707,N_3717,N_4899);
or U6708 (N_6708,N_2487,N_357);
nor U6709 (N_6709,N_4516,N_4911);
nor U6710 (N_6710,N_516,N_2262);
and U6711 (N_6711,N_3204,N_1527);
and U6712 (N_6712,N_1120,N_3009);
nand U6713 (N_6713,N_128,N_11);
or U6714 (N_6714,N_4045,N_1369);
and U6715 (N_6715,N_576,N_4293);
or U6716 (N_6716,N_4726,N_4770);
nand U6717 (N_6717,N_3232,N_3097);
nor U6718 (N_6718,N_1039,N_4783);
nor U6719 (N_6719,N_2933,N_2812);
or U6720 (N_6720,N_3011,N_403);
nand U6721 (N_6721,N_3840,N_130);
nand U6722 (N_6722,N_108,N_3778);
nor U6723 (N_6723,N_4483,N_152);
nand U6724 (N_6724,N_241,N_2871);
or U6725 (N_6725,N_4151,N_4272);
nand U6726 (N_6726,N_1966,N_4982);
nand U6727 (N_6727,N_4331,N_2087);
or U6728 (N_6728,N_4531,N_2882);
and U6729 (N_6729,N_863,N_2518);
and U6730 (N_6730,N_3675,N_715);
or U6731 (N_6731,N_2739,N_310);
xnor U6732 (N_6732,N_2732,N_3170);
nand U6733 (N_6733,N_1769,N_3826);
and U6734 (N_6734,N_587,N_4132);
nand U6735 (N_6735,N_113,N_1159);
or U6736 (N_6736,N_1329,N_4606);
or U6737 (N_6737,N_3381,N_105);
nor U6738 (N_6738,N_3168,N_793);
and U6739 (N_6739,N_469,N_3266);
or U6740 (N_6740,N_2101,N_3556);
nand U6741 (N_6741,N_2121,N_4924);
and U6742 (N_6742,N_3002,N_4703);
or U6743 (N_6743,N_2387,N_2856);
or U6744 (N_6744,N_1459,N_4283);
and U6745 (N_6745,N_4722,N_2863);
and U6746 (N_6746,N_226,N_2333);
nor U6747 (N_6747,N_4141,N_3713);
nor U6748 (N_6748,N_1959,N_684);
nand U6749 (N_6749,N_3935,N_1699);
or U6750 (N_6750,N_1571,N_2476);
and U6751 (N_6751,N_4651,N_1788);
or U6752 (N_6752,N_347,N_162);
or U6753 (N_6753,N_293,N_979);
nand U6754 (N_6754,N_2130,N_2626);
or U6755 (N_6755,N_3694,N_456);
nand U6756 (N_6756,N_859,N_2712);
nand U6757 (N_6757,N_1980,N_3050);
nor U6758 (N_6758,N_4359,N_820);
nor U6759 (N_6759,N_3970,N_501);
and U6760 (N_6760,N_1398,N_2186);
or U6761 (N_6761,N_730,N_4104);
or U6762 (N_6762,N_4561,N_3559);
nand U6763 (N_6763,N_4223,N_97);
or U6764 (N_6764,N_2290,N_1454);
or U6765 (N_6765,N_369,N_1496);
xor U6766 (N_6766,N_4335,N_2571);
and U6767 (N_6767,N_1155,N_3430);
or U6768 (N_6768,N_947,N_827);
or U6769 (N_6769,N_1568,N_1951);
nor U6770 (N_6770,N_3745,N_3957);
or U6771 (N_6771,N_443,N_3312);
and U6772 (N_6772,N_3633,N_2753);
and U6773 (N_6773,N_915,N_3101);
nand U6774 (N_6774,N_1736,N_2866);
nand U6775 (N_6775,N_3716,N_2289);
nand U6776 (N_6776,N_4098,N_3771);
nand U6777 (N_6777,N_3138,N_1105);
or U6778 (N_6778,N_2822,N_3373);
nand U6779 (N_6779,N_1771,N_2966);
and U6780 (N_6780,N_1179,N_3595);
nand U6781 (N_6781,N_2045,N_668);
and U6782 (N_6782,N_2716,N_3773);
or U6783 (N_6783,N_1578,N_2981);
nand U6784 (N_6784,N_3325,N_3956);
or U6785 (N_6785,N_2695,N_513);
nand U6786 (N_6786,N_2439,N_270);
and U6787 (N_6787,N_3436,N_4196);
and U6788 (N_6788,N_397,N_1696);
nor U6789 (N_6789,N_174,N_1115);
and U6790 (N_6790,N_245,N_956);
nand U6791 (N_6791,N_4570,N_1297);
nor U6792 (N_6792,N_1192,N_4989);
nand U6793 (N_6793,N_1821,N_71);
or U6794 (N_6794,N_3218,N_1506);
nor U6795 (N_6795,N_2258,N_4039);
xor U6796 (N_6796,N_4022,N_327);
nor U6797 (N_6797,N_4365,N_4229);
nand U6798 (N_6798,N_3432,N_129);
nor U6799 (N_6799,N_311,N_4161);
or U6800 (N_6800,N_4663,N_1823);
nand U6801 (N_6801,N_3118,N_3877);
nand U6802 (N_6802,N_445,N_389);
xnor U6803 (N_6803,N_2734,N_2699);
nand U6804 (N_6804,N_792,N_3281);
or U6805 (N_6805,N_131,N_509);
and U6806 (N_6806,N_4467,N_3330);
nand U6807 (N_6807,N_488,N_1749);
nand U6808 (N_6808,N_364,N_4789);
nand U6809 (N_6809,N_1012,N_4704);
or U6810 (N_6810,N_2083,N_3196);
nor U6811 (N_6811,N_2480,N_4815);
and U6812 (N_6812,N_74,N_2618);
and U6813 (N_6813,N_4587,N_4563);
nand U6814 (N_6814,N_3746,N_3581);
and U6815 (N_6815,N_1841,N_3259);
nand U6816 (N_6816,N_2198,N_1089);
nand U6817 (N_6817,N_2659,N_2226);
or U6818 (N_6818,N_669,N_3954);
nor U6819 (N_6819,N_3995,N_1201);
or U6820 (N_6820,N_2539,N_4024);
nor U6821 (N_6821,N_2656,N_2715);
nand U6822 (N_6822,N_2680,N_1141);
or U6823 (N_6823,N_1040,N_2531);
nor U6824 (N_6824,N_4445,N_2816);
nand U6825 (N_6825,N_3183,N_4856);
nor U6826 (N_6826,N_3016,N_476);
xnor U6827 (N_6827,N_4037,N_30);
nand U6828 (N_6828,N_2728,N_2873);
nor U6829 (N_6829,N_1520,N_1498);
nand U6830 (N_6830,N_3804,N_3328);
nand U6831 (N_6831,N_319,N_941);
nor U6832 (N_6832,N_3592,N_2707);
nor U6833 (N_6833,N_81,N_3249);
nor U6834 (N_6834,N_2951,N_880);
nor U6835 (N_6835,N_3867,N_867);
nand U6836 (N_6836,N_1442,N_4370);
nand U6837 (N_6837,N_1285,N_1361);
nand U6838 (N_6838,N_500,N_4675);
or U6839 (N_6839,N_710,N_4397);
or U6840 (N_6840,N_2285,N_3431);
nand U6841 (N_6841,N_4750,N_4716);
or U6842 (N_6842,N_4831,N_3468);
nand U6843 (N_6843,N_3192,N_2640);
and U6844 (N_6844,N_2718,N_201);
and U6845 (N_6845,N_2284,N_4931);
or U6846 (N_6846,N_1081,N_4808);
nand U6847 (N_6847,N_4231,N_3001);
or U6848 (N_6848,N_2043,N_1971);
and U6849 (N_6849,N_2973,N_1429);
nor U6850 (N_6850,N_3875,N_2176);
nand U6851 (N_6851,N_4501,N_4308);
nand U6852 (N_6852,N_659,N_1548);
and U6853 (N_6853,N_4135,N_2820);
or U6854 (N_6854,N_3843,N_3361);
or U6855 (N_6855,N_3068,N_1021);
nor U6856 (N_6856,N_3070,N_2696);
nor U6857 (N_6857,N_3751,N_4980);
and U6858 (N_6858,N_1029,N_1217);
nand U6859 (N_6859,N_1643,N_4674);
or U6860 (N_6860,N_3225,N_3242);
and U6861 (N_6861,N_1754,N_4394);
nand U6862 (N_6862,N_1907,N_2876);
and U6863 (N_6863,N_2365,N_525);
nand U6864 (N_6864,N_4412,N_2328);
nand U6865 (N_6865,N_2711,N_219);
or U6866 (N_6866,N_4300,N_3254);
nor U6867 (N_6867,N_782,N_1146);
and U6868 (N_6868,N_3962,N_3);
nand U6869 (N_6869,N_2950,N_1603);
nor U6870 (N_6870,N_4599,N_3942);
or U6871 (N_6871,N_2792,N_2368);
or U6872 (N_6872,N_4799,N_4588);
nor U6873 (N_6873,N_812,N_3809);
nand U6874 (N_6874,N_1847,N_3910);
nand U6875 (N_6875,N_1584,N_4070);
and U6876 (N_6876,N_2076,N_3309);
and U6877 (N_6877,N_1218,N_2860);
or U6878 (N_6878,N_4013,N_2977);
nor U6879 (N_6879,N_1961,N_3088);
or U6880 (N_6880,N_607,N_1848);
and U6881 (N_6881,N_2470,N_4147);
or U6882 (N_6882,N_235,N_3847);
nand U6883 (N_6883,N_1026,N_4849);
or U6884 (N_6884,N_2046,N_373);
or U6885 (N_6885,N_4055,N_109);
or U6886 (N_6886,N_204,N_1436);
or U6887 (N_6887,N_1910,N_1691);
nand U6888 (N_6888,N_2194,N_208);
or U6889 (N_6889,N_1709,N_4148);
nor U6890 (N_6890,N_2960,N_3461);
nor U6891 (N_6891,N_740,N_4321);
or U6892 (N_6892,N_1049,N_4084);
or U6893 (N_6893,N_705,N_1544);
or U6894 (N_6894,N_4505,N_4203);
and U6895 (N_6895,N_4502,N_626);
and U6896 (N_6896,N_211,N_987);
or U6897 (N_6897,N_111,N_137);
nor U6898 (N_6898,N_3955,N_2648);
nor U6899 (N_6899,N_1310,N_786);
and U6900 (N_6900,N_2691,N_3814);
and U6901 (N_6901,N_1740,N_3137);
nand U6902 (N_6902,N_896,N_3983);
nor U6903 (N_6903,N_2837,N_2438);
or U6904 (N_6904,N_2282,N_3451);
nor U6905 (N_6905,N_4111,N_1487);
or U6906 (N_6906,N_3570,N_25);
nor U6907 (N_6907,N_1930,N_2484);
nand U6908 (N_6908,N_1528,N_4307);
or U6909 (N_6909,N_3380,N_4162);
nor U6910 (N_6910,N_3629,N_1470);
nor U6911 (N_6911,N_265,N_4677);
and U6912 (N_6912,N_1167,N_934);
or U6913 (N_6913,N_1759,N_4788);
or U6914 (N_6914,N_1838,N_1795);
nand U6915 (N_6915,N_4338,N_697);
or U6916 (N_6916,N_284,N_4282);
or U6917 (N_6917,N_2765,N_1037);
nor U6918 (N_6918,N_4768,N_2612);
nand U6919 (N_6919,N_1639,N_3211);
xnor U6920 (N_6920,N_2787,N_3926);
and U6921 (N_6921,N_3411,N_4719);
nor U6922 (N_6922,N_3369,N_716);
and U6923 (N_6923,N_4986,N_2199);
and U6924 (N_6924,N_986,N_420);
nor U6925 (N_6925,N_2030,N_1871);
and U6926 (N_6926,N_879,N_2743);
and U6927 (N_6927,N_4437,N_176);
nand U6928 (N_6928,N_1854,N_1632);
or U6929 (N_6929,N_3191,N_3750);
xnor U6930 (N_6930,N_1845,N_4184);
nand U6931 (N_6931,N_85,N_4582);
and U6932 (N_6932,N_1819,N_2436);
nand U6933 (N_6933,N_4934,N_2342);
or U6934 (N_6934,N_164,N_779);
xnor U6935 (N_6935,N_4901,N_3685);
nor U6936 (N_6936,N_1080,N_2551);
and U6937 (N_6937,N_931,N_12);
nor U6938 (N_6938,N_967,N_2661);
and U6939 (N_6939,N_1772,N_591);
nand U6940 (N_6940,N_1410,N_1197);
and U6941 (N_6941,N_714,N_4933);
nor U6942 (N_6942,N_4249,N_1463);
nand U6943 (N_6943,N_2006,N_4109);
nand U6944 (N_6944,N_2050,N_2002);
or U6945 (N_6945,N_3060,N_1018);
nor U6946 (N_6946,N_4957,N_3548);
nand U6947 (N_6947,N_1607,N_1753);
or U6948 (N_6948,N_2388,N_4551);
nand U6949 (N_6949,N_4120,N_4415);
and U6950 (N_6950,N_1963,N_2188);
nand U6951 (N_6951,N_581,N_4127);
nand U6952 (N_6952,N_3270,N_3409);
nor U6953 (N_6953,N_3993,N_2717);
nor U6954 (N_6954,N_2293,N_303);
and U6955 (N_6955,N_4735,N_2982);
nor U6956 (N_6956,N_3887,N_376);
and U6957 (N_6957,N_1630,N_1593);
and U6958 (N_6958,N_317,N_3734);
and U6959 (N_6959,N_2713,N_1999);
nand U6960 (N_6960,N_4376,N_1054);
nand U6961 (N_6961,N_2915,N_3852);
nand U6962 (N_6962,N_2203,N_2846);
nand U6963 (N_6963,N_787,N_8);
nand U6964 (N_6964,N_3176,N_3044);
or U6965 (N_6965,N_558,N_4217);
nand U6966 (N_6966,N_1946,N_2795);
nor U6967 (N_6967,N_3743,N_709);
and U6968 (N_6968,N_2954,N_4910);
and U6969 (N_6969,N_3210,N_1110);
and U6970 (N_6970,N_3944,N_4140);
nor U6971 (N_6971,N_1425,N_2583);
nor U6972 (N_6972,N_913,N_2935);
nor U6973 (N_6973,N_3912,N_663);
or U6974 (N_6974,N_2243,N_4556);
nand U6975 (N_6975,N_240,N_813);
nand U6976 (N_6976,N_1023,N_2606);
or U6977 (N_6977,N_1649,N_181);
or U6978 (N_6978,N_2579,N_3207);
and U6979 (N_6979,N_1935,N_4423);
nor U6980 (N_6980,N_3687,N_1193);
nand U6981 (N_6981,N_2448,N_2558);
nand U6982 (N_6982,N_983,N_1467);
nor U6983 (N_6983,N_4462,N_1009);
or U6984 (N_6984,N_3941,N_3153);
nor U6985 (N_6985,N_2731,N_1562);
or U6986 (N_6986,N_1636,N_2459);
or U6987 (N_6987,N_4577,N_439);
nor U6988 (N_6988,N_4872,N_1083);
or U6989 (N_6989,N_4909,N_667);
nor U6990 (N_6990,N_2035,N_4597);
and U6991 (N_6991,N_2054,N_3435);
nor U6992 (N_6992,N_3798,N_4079);
and U6993 (N_6993,N_972,N_4069);
nor U6994 (N_6994,N_141,N_1461);
and U6995 (N_6995,N_3538,N_960);
nor U6996 (N_6996,N_548,N_215);
nor U6997 (N_6997,N_2029,N_2494);
and U6998 (N_6998,N_4025,N_3733);
and U6999 (N_6999,N_2859,N_4731);
and U7000 (N_7000,N_4137,N_2797);
nor U7001 (N_7001,N_856,N_2353);
nand U7002 (N_7002,N_2990,N_1637);
nor U7003 (N_7003,N_2306,N_801);
nor U7004 (N_7004,N_4573,N_1060);
nand U7005 (N_7005,N_4418,N_1987);
nor U7006 (N_7006,N_4676,N_3674);
or U7007 (N_7007,N_2026,N_1484);
or U7008 (N_7008,N_3921,N_3388);
nor U7009 (N_7009,N_2109,N_4303);
or U7010 (N_7010,N_2808,N_45);
nand U7011 (N_7011,N_379,N_234);
and U7012 (N_7012,N_1822,N_1733);
or U7013 (N_7013,N_2932,N_269);
nand U7014 (N_7014,N_1271,N_4621);
nand U7015 (N_7015,N_2434,N_4546);
nand U7016 (N_7016,N_2498,N_3151);
or U7017 (N_7017,N_4002,N_2212);
or U7018 (N_7018,N_1836,N_2694);
and U7019 (N_7019,N_2271,N_4031);
nand U7020 (N_7020,N_4026,N_1418);
and U7021 (N_7021,N_4974,N_2000);
nor U7022 (N_7022,N_2279,N_3911);
or U7023 (N_7023,N_3769,N_2347);
nand U7024 (N_7024,N_4779,N_746);
nor U7025 (N_7025,N_2980,N_783);
or U7026 (N_7026,N_3172,N_4707);
nor U7027 (N_7027,N_2686,N_846);
nand U7028 (N_7028,N_1044,N_3311);
nand U7029 (N_7029,N_3429,N_4834);
or U7030 (N_7030,N_4358,N_4721);
nand U7031 (N_7031,N_1433,N_3108);
nand U7032 (N_7032,N_3003,N_2886);
nor U7033 (N_7033,N_3779,N_2171);
or U7034 (N_7034,N_900,N_1536);
nor U7035 (N_7035,N_969,N_4657);
or U7036 (N_7036,N_4795,N_3511);
and U7037 (N_7037,N_1,N_4453);
nand U7038 (N_7038,N_3860,N_3427);
nand U7039 (N_7039,N_864,N_963);
and U7040 (N_7040,N_4427,N_2641);
nor U7041 (N_7041,N_4792,N_2251);
and U7042 (N_7042,N_3709,N_3698);
and U7043 (N_7043,N_875,N_2851);
nand U7044 (N_7044,N_4092,N_1853);
nand U7045 (N_7045,N_4545,N_3946);
nor U7046 (N_7046,N_79,N_1131);
or U7047 (N_7047,N_3651,N_949);
nand U7048 (N_7048,N_1500,N_1262);
or U7049 (N_7049,N_4493,N_1531);
xnor U7050 (N_7050,N_4480,N_876);
nor U7051 (N_7051,N_2834,N_173);
and U7052 (N_7052,N_4178,N_59);
nor U7053 (N_7053,N_1408,N_2682);
or U7054 (N_7054,N_1521,N_1062);
nand U7055 (N_7055,N_2943,N_3466);
nand U7056 (N_7056,N_2482,N_633);
or U7057 (N_7057,N_1079,N_3748);
and U7058 (N_7058,N_3337,N_2473);
nor U7059 (N_7059,N_51,N_3722);
and U7060 (N_7060,N_3996,N_4946);
or U7061 (N_7061,N_4299,N_1697);
or U7062 (N_7062,N_3092,N_1725);
nor U7063 (N_7063,N_3458,N_3881);
or U7064 (N_7064,N_4105,N_2634);
and U7065 (N_7065,N_2206,N_1887);
nand U7066 (N_7066,N_4784,N_4169);
nor U7067 (N_7067,N_2055,N_4181);
nor U7068 (N_7068,N_2794,N_91);
nor U7069 (N_7069,N_534,N_2346);
and U7070 (N_7070,N_2817,N_3413);
nor U7071 (N_7071,N_4878,N_3058);
and U7072 (N_7072,N_410,N_281);
nand U7073 (N_7073,N_4420,N_4944);
nand U7074 (N_7074,N_3671,N_925);
nor U7075 (N_7075,N_3421,N_2114);
or U7076 (N_7076,N_2234,N_250);
nor U7077 (N_7077,N_2642,N_4438);
nand U7078 (N_7078,N_4216,N_3578);
nand U7079 (N_7079,N_3683,N_449);
or U7080 (N_7080,N_4361,N_2867);
or U7081 (N_7081,N_1858,N_3605);
nor U7082 (N_7082,N_3985,N_2790);
and U7083 (N_7083,N_4604,N_3628);
nor U7084 (N_7084,N_3563,N_4640);
nand U7085 (N_7085,N_4615,N_3729);
nand U7086 (N_7086,N_4327,N_3943);
and U7087 (N_7087,N_4410,N_4904);
and U7088 (N_7088,N_4645,N_2590);
nand U7089 (N_7089,N_889,N_2490);
nand U7090 (N_7090,N_1611,N_1671);
or U7091 (N_7091,N_4471,N_1494);
nor U7092 (N_7092,N_2136,N_694);
or U7093 (N_7093,N_4806,N_4495);
or U7094 (N_7094,N_1766,N_39);
nor U7095 (N_7095,N_4780,N_3334);
or U7096 (N_7096,N_490,N_133);
or U7097 (N_7097,N_1088,N_87);
or U7098 (N_7098,N_4367,N_3665);
or U7099 (N_7099,N_64,N_3255);
nor U7100 (N_7100,N_860,N_3256);
nor U7101 (N_7101,N_1438,N_4043);
nand U7102 (N_7102,N_609,N_4371);
nand U7103 (N_7103,N_4524,N_3046);
xor U7104 (N_7104,N_1683,N_4860);
and U7105 (N_7105,N_1919,N_4758);
nor U7106 (N_7106,N_2929,N_3013);
nor U7107 (N_7107,N_4712,N_3859);
nor U7108 (N_7108,N_2595,N_2355);
nor U7109 (N_7109,N_4188,N_2483);
or U7110 (N_7110,N_1663,N_1805);
nand U7111 (N_7111,N_1949,N_2620);
nor U7112 (N_7112,N_3467,N_538);
and U7113 (N_7113,N_1228,N_842);
and U7114 (N_7114,N_2478,N_1290);
nand U7115 (N_7115,N_3355,N_3898);
nor U7116 (N_7116,N_4201,N_1713);
nand U7117 (N_7117,N_4484,N_4961);
nor U7118 (N_7118,N_4723,N_2941);
and U7119 (N_7119,N_3816,N_506);
nor U7120 (N_7120,N_1082,N_2399);
nand U7121 (N_7121,N_2609,N_2737);
nor U7122 (N_7122,N_1507,N_3951);
or U7123 (N_7123,N_2724,N_2410);
or U7124 (N_7124,N_2522,N_392);
and U7125 (N_7125,N_1522,N_3587);
nor U7126 (N_7126,N_2103,N_888);
nor U7127 (N_7127,N_1677,N_2909);
and U7128 (N_7128,N_776,N_4610);
nand U7129 (N_7129,N_225,N_4036);
nor U7130 (N_7130,N_4696,N_4250);
or U7131 (N_7131,N_3371,N_422);
or U7132 (N_7132,N_1171,N_4603);
nand U7133 (N_7133,N_580,N_2443);
nor U7134 (N_7134,N_1352,N_4747);
nor U7135 (N_7135,N_2091,N_297);
and U7136 (N_7136,N_2354,N_2592);
nand U7137 (N_7137,N_2037,N_4465);
nor U7138 (N_7138,N_3739,N_4191);
nand U7139 (N_7139,N_3428,N_3958);
or U7140 (N_7140,N_3835,N_788);
or U7141 (N_7141,N_4154,N_3372);
nor U7142 (N_7142,N_3781,N_4085);
or U7143 (N_7143,N_654,N_3642);
nand U7144 (N_7144,N_344,N_2831);
and U7145 (N_7145,N_4489,N_2768);
nor U7146 (N_7146,N_4772,N_4356);
nor U7147 (N_7147,N_826,N_2986);
xnor U7148 (N_7148,N_1676,N_1439);
and U7149 (N_7149,N_901,N_851);
nor U7150 (N_7150,N_1052,N_994);
nand U7151 (N_7151,N_3106,N_4813);
nand U7152 (N_7152,N_2761,N_619);
nand U7153 (N_7153,N_3462,N_707);
nand U7154 (N_7154,N_3679,N_2657);
nor U7155 (N_7155,N_2323,N_2115);
and U7156 (N_7156,N_1471,N_1265);
or U7157 (N_7157,N_2182,N_835);
nor U7158 (N_7158,N_3455,N_3507);
or U7159 (N_7159,N_1437,N_1542);
nand U7160 (N_7160,N_1375,N_121);
nor U7161 (N_7161,N_409,N_2697);
or U7162 (N_7162,N_3770,N_2926);
and U7163 (N_7163,N_4644,N_1288);
or U7164 (N_7164,N_2308,N_815);
nand U7165 (N_7165,N_502,N_4349);
and U7166 (N_7166,N_965,N_2141);
nor U7167 (N_7167,N_2767,N_1205);
nor U7168 (N_7168,N_545,N_4994);
nand U7169 (N_7169,N_2593,N_282);
nor U7170 (N_7170,N_4862,N_4553);
and U7171 (N_7171,N_1158,N_3329);
and U7172 (N_7172,N_2380,N_3171);
or U7173 (N_7173,N_2341,N_2905);
nand U7174 (N_7174,N_1947,N_3608);
or U7175 (N_7175,N_2219,N_4614);
and U7176 (N_7176,N_1108,N_3367);
nand U7177 (N_7177,N_1125,N_387);
nor U7178 (N_7178,N_1803,N_1395);
nand U7179 (N_7179,N_4970,N_2413);
nand U7180 (N_7180,N_190,N_4131);
and U7181 (N_7181,N_2381,N_4324);
and U7182 (N_7182,N_3111,N_2598);
nand U7183 (N_7183,N_3589,N_3738);
nor U7184 (N_7184,N_4378,N_465);
and U7185 (N_7185,N_65,N_4514);
nand U7186 (N_7186,N_974,N_4481);
and U7187 (N_7187,N_1160,N_666);
nor U7188 (N_7188,N_4876,N_2471);
nor U7189 (N_7189,N_4130,N_1760);
or U7190 (N_7190,N_1119,N_3400);
nor U7191 (N_7191,N_1680,N_2537);
or U7192 (N_7192,N_4020,N_2891);
nand U7193 (N_7193,N_1497,N_3724);
and U7194 (N_7194,N_861,N_3021);
or U7195 (N_7195,N_3557,N_3104);
or U7196 (N_7196,N_2894,N_2146);
xor U7197 (N_7197,N_231,N_3306);
xnor U7198 (N_7198,N_2462,N_1414);
or U7199 (N_7199,N_2089,N_2140);
and U7200 (N_7200,N_4952,N_4264);
nand U7201 (N_7201,N_4697,N_2588);
and U7202 (N_7202,N_2079,N_3393);
xnor U7203 (N_7203,N_4936,N_653);
nand U7204 (N_7204,N_1802,N_3269);
and U7205 (N_7205,N_1294,N_3268);
or U7206 (N_7206,N_4839,N_4642);
nand U7207 (N_7207,N_2449,N_1103);
nor U7208 (N_7208,N_3526,N_1872);
nand U7209 (N_7209,N_3349,N_3043);
or U7210 (N_7210,N_1564,N_2168);
nor U7211 (N_7211,N_840,N_2912);
nand U7212 (N_7212,N_816,N_368);
or U7213 (N_7213,N_613,N_58);
nor U7214 (N_7214,N_962,N_3014);
nor U7215 (N_7215,N_4947,N_1431);
and U7216 (N_7216,N_1254,N_572);
nor U7217 (N_7217,N_2156,N_492);
nand U7218 (N_7218,N_2835,N_1859);
nand U7219 (N_7219,N_72,N_3403);
nor U7220 (N_7220,N_1922,N_487);
xnor U7221 (N_7221,N_951,N_2142);
and U7222 (N_7222,N_4898,N_976);
nand U7223 (N_7223,N_3618,N_3220);
and U7224 (N_7224,N_1415,N_3362);
nand U7225 (N_7225,N_3182,N_4391);
or U7226 (N_7226,N_3035,N_4318);
nand U7227 (N_7227,N_4354,N_1519);
nor U7228 (N_7228,N_964,N_4686);
nand U7229 (N_7229,N_2624,N_3387);
or U7230 (N_7230,N_1557,N_1302);
and U7231 (N_7231,N_198,N_1719);
nor U7232 (N_7232,N_4691,N_110);
and U7233 (N_7233,N_2096,N_1349);
and U7234 (N_7234,N_1767,N_4966);
nor U7235 (N_7235,N_1635,N_196);
nand U7236 (N_7236,N_4517,N_2418);
and U7237 (N_7237,N_16,N_3122);
nand U7238 (N_7238,N_415,N_2165);
or U7239 (N_7239,N_899,N_95);
nand U7240 (N_7240,N_4706,N_2384);
nand U7241 (N_7241,N_1198,N_1950);
nor U7242 (N_7242,N_4029,N_2533);
or U7243 (N_7243,N_4230,N_4988);
xnor U7244 (N_7244,N_67,N_627);
nor U7245 (N_7245,N_268,N_3129);
xor U7246 (N_7246,N_4518,N_882);
nand U7247 (N_7247,N_374,N_1252);
nand U7248 (N_7248,N_2178,N_3631);
and U7249 (N_7249,N_2631,N_4923);
and U7250 (N_7250,N_4393,N_1363);
or U7251 (N_7251,N_4357,N_561);
or U7252 (N_7252,N_1245,N_3506);
or U7253 (N_7253,N_4403,N_521);
nand U7254 (N_7254,N_2389,N_4918);
nor U7255 (N_7255,N_2733,N_244);
nand U7256 (N_7256,N_307,N_1569);
and U7257 (N_7257,N_1915,N_4295);
nand U7258 (N_7258,N_2627,N_2692);
and U7259 (N_7259,N_3327,N_4432);
nor U7260 (N_7260,N_2547,N_4133);
and U7261 (N_7261,N_1111,N_1720);
or U7262 (N_7262,N_2222,N_2810);
and U7263 (N_7263,N_4678,N_721);
nand U7264 (N_7264,N_2965,N_154);
nand U7265 (N_7265,N_4682,N_4807);
xnor U7266 (N_7266,N_360,N_4760);
or U7267 (N_7267,N_2331,N_3086);
nand U7268 (N_7268,N_2940,N_4330);
and U7269 (N_7269,N_4646,N_228);
nand U7270 (N_7270,N_2811,N_3341);
and U7271 (N_7271,N_995,N_3841);
or U7272 (N_7272,N_758,N_1727);
nand U7273 (N_7273,N_552,N_4433);
and U7274 (N_7274,N_4748,N_203);
nand U7275 (N_7275,N_3094,N_43);
nor U7276 (N_7276,N_1834,N_2956);
or U7277 (N_7277,N_3399,N_4218);
or U7278 (N_7278,N_3078,N_3815);
nand U7279 (N_7279,N_1580,N_434);
nand U7280 (N_7280,N_2192,N_2601);
nor U7281 (N_7281,N_588,N_4900);
or U7282 (N_7282,N_460,N_3298);
xor U7283 (N_7283,N_1386,N_1139);
nor U7284 (N_7284,N_92,N_2993);
nand U7285 (N_7285,N_4287,N_4362);
or U7286 (N_7286,N_2455,N_3864);
nor U7287 (N_7287,N_1898,N_3338);
nor U7288 (N_7288,N_2261,N_4207);
nor U7289 (N_7289,N_3753,N_4533);
or U7290 (N_7290,N_3836,N_560);
nor U7291 (N_7291,N_1540,N_437);
or U7292 (N_7292,N_1367,N_2059);
and U7293 (N_7293,N_1716,N_2949);
nand U7294 (N_7294,N_1833,N_3626);
nor U7295 (N_7295,N_1114,N_463);
nand U7296 (N_7296,N_3363,N_632);
nor U7297 (N_7297,N_1289,N_1662);
or U7298 (N_7298,N_3834,N_2917);
nor U7299 (N_7299,N_2937,N_3279);
or U7300 (N_7300,N_1058,N_1453);
and U7301 (N_7301,N_3873,N_470);
and U7302 (N_7302,N_3040,N_4049);
xor U7303 (N_7303,N_147,N_2393);
or U7304 (N_7304,N_1977,N_4743);
or U7305 (N_7305,N_2796,N_1555);
nand U7306 (N_7306,N_3161,N_3112);
nor U7307 (N_7307,N_998,N_1628);
or U7308 (N_7308,N_4559,N_19);
and U7309 (N_7309,N_1462,N_1929);
or U7310 (N_7310,N_358,N_1831);
nor U7311 (N_7311,N_2839,N_2466);
nand U7312 (N_7312,N_2268,N_1328);
nand U7313 (N_7313,N_2502,N_2107);
and U7314 (N_7314,N_4506,N_4082);
nor U7315 (N_7315,N_2922,N_4835);
or U7316 (N_7316,N_3140,N_2208);
and U7317 (N_7317,N_3053,N_3195);
or U7318 (N_7318,N_4008,N_2272);
or U7319 (N_7319,N_4408,N_3546);
nor U7320 (N_7320,N_3475,N_1690);
and U7321 (N_7321,N_1800,N_4548);
or U7322 (N_7322,N_1144,N_1241);
and U7323 (N_7323,N_4892,N_4115);
nor U7324 (N_7324,N_1645,N_3440);
nand U7325 (N_7325,N_1219,N_330);
nor U7326 (N_7326,N_2804,N_781);
nor U7327 (N_7327,N_696,N_1169);
or U7328 (N_7328,N_136,N_3825);
and U7329 (N_7329,N_3064,N_1509);
nor U7330 (N_7330,N_3163,N_1195);
nand U7331 (N_7331,N_1320,N_442);
nor U7332 (N_7332,N_3585,N_2857);
nor U7333 (N_7333,N_4929,N_230);
nor U7334 (N_7334,N_3573,N_1250);
nand U7335 (N_7335,N_4884,N_1032);
nand U7336 (N_7336,N_260,N_3368);
nand U7337 (N_7337,N_306,N_477);
and U7338 (N_7338,N_2407,N_517);
or U7339 (N_7339,N_652,N_2159);
nor U7340 (N_7340,N_356,N_2928);
nor U7341 (N_7341,N_2019,N_3998);
nand U7342 (N_7342,N_4414,N_2742);
nor U7343 (N_7343,N_4450,N_553);
nor U7344 (N_7344,N_2173,N_3562);
nor U7345 (N_7345,N_1069,N_1293);
nor U7346 (N_7346,N_1441,N_4180);
or U7347 (N_7347,N_146,N_810);
xor U7348 (N_7348,N_643,N_4326);
nand U7349 (N_7349,N_1313,N_2852);
nor U7350 (N_7350,N_4940,N_1268);
or U7351 (N_7351,N_1273,N_3221);
or U7352 (N_7352,N_2884,N_4736);
and U7353 (N_7353,N_550,N_28);
and U7354 (N_7354,N_3167,N_1258);
nand U7355 (N_7355,N_462,N_4793);
and U7356 (N_7356,N_3406,N_3307);
and U7357 (N_7357,N_767,N_2412);
and U7358 (N_7358,N_2506,N_3227);
nand U7359 (N_7359,N_2972,N_218);
nor U7360 (N_7360,N_4096,N_2504);
nor U7361 (N_7361,N_331,N_4589);
nor U7362 (N_7362,N_990,N_276);
and U7363 (N_7363,N_2670,N_2746);
or U7364 (N_7364,N_1031,N_1316);
xor U7365 (N_7365,N_1748,N_2143);
nor U7366 (N_7366,N_3240,N_261);
nor U7367 (N_7367,N_18,N_761);
or U7368 (N_7368,N_2683,N_2351);
nand U7369 (N_7369,N_36,N_4757);
and U7370 (N_7370,N_299,N_3678);
nor U7371 (N_7371,N_1815,N_263);
nor U7372 (N_7372,N_2519,N_4881);
or U7373 (N_7373,N_1983,N_3513);
or U7374 (N_7374,N_2678,N_4103);
or U7375 (N_7375,N_4129,N_639);
nor U7376 (N_7376,N_243,N_646);
or U7377 (N_7377,N_1513,N_3856);
or U7378 (N_7378,N_2968,N_997);
nor U7379 (N_7379,N_2633,N_4781);
xor U7380 (N_7380,N_1010,N_4796);
or U7381 (N_7381,N_1516,N_2607);
and U7382 (N_7382,N_2067,N_4139);
or U7383 (N_7383,N_530,N_2690);
or U7384 (N_7384,N_1385,N_625);
and U7385 (N_7385,N_1541,N_870);
or U7386 (N_7386,N_926,N_567);
nand U7387 (N_7387,N_2044,N_1705);
or U7388 (N_7388,N_692,N_1565);
and U7389 (N_7389,N_2209,N_3757);
nor U7390 (N_7390,N_2240,N_4472);
nor U7391 (N_7391,N_350,N_2495);
nor U7392 (N_7392,N_4912,N_3803);
nand U7393 (N_7393,N_257,N_693);
and U7394 (N_7394,N_2469,N_1107);
or U7395 (N_7395,N_1016,N_3668);
and U7396 (N_7396,N_432,N_4023);
and U7397 (N_7397,N_1486,N_2638);
or U7398 (N_7398,N_953,N_4225);
and U7399 (N_7399,N_3558,N_3959);
or U7400 (N_7400,N_1508,N_247);
nand U7401 (N_7401,N_1969,N_4896);
nor U7402 (N_7402,N_2303,N_3737);
and U7403 (N_7403,N_2962,N_3180);
nor U7404 (N_7404,N_2220,N_2325);
nand U7405 (N_7405,N_3439,N_2885);
nor U7406 (N_7406,N_3964,N_384);
and U7407 (N_7407,N_278,N_1065);
nor U7408 (N_7408,N_760,N_2806);
nor U7409 (N_7409,N_2848,N_2047);
and U7410 (N_7410,N_2946,N_3027);
or U7411 (N_7411,N_673,N_3561);
and U7412 (N_7412,N_1655,N_599);
nor U7413 (N_7413,N_2783,N_4066);
and U7414 (N_7414,N_2786,N_1711);
and U7415 (N_7415,N_569,N_1443);
nor U7416 (N_7416,N_1656,N_2881);
nand U7417 (N_7417,N_3621,N_380);
nand U7418 (N_7418,N_804,N_3414);
and U7419 (N_7419,N_1482,N_1918);
or U7420 (N_7420,N_2095,N_2596);
nand U7421 (N_7421,N_160,N_1020);
and U7422 (N_7422,N_924,N_1237);
nand U7423 (N_7423,N_4917,N_4494);
nor U7424 (N_7424,N_2628,N_4027);
and U7425 (N_7425,N_286,N_1256);
and U7426 (N_7426,N_165,N_4919);
nand U7427 (N_7427,N_754,N_2105);
nand U7428 (N_7428,N_937,N_1688);
or U7429 (N_7429,N_3303,N_3394);
or U7430 (N_7430,N_2556,N_309);
or U7431 (N_7431,N_3806,N_3652);
nor U7432 (N_7432,N_478,N_493);
and U7433 (N_7433,N_4387,N_911);
or U7434 (N_7434,N_2385,N_2433);
and U7435 (N_7435,N_271,N_2071);
and U7436 (N_7436,N_4991,N_3696);
and U7437 (N_7437,N_1718,N_2250);
and U7438 (N_7438,N_4653,N_2190);
or U7439 (N_7439,N_2366,N_4200);
or U7440 (N_7440,N_4764,N_1962);
and U7441 (N_7441,N_4734,N_702);
nand U7442 (N_7442,N_3423,N_287);
xnor U7443 (N_7443,N_4555,N_2185);
or U7444 (N_7444,N_2759,N_142);
nor U7445 (N_7445,N_1196,N_3789);
nand U7446 (N_7446,N_4804,N_2512);
nand U7447 (N_7447,N_2236,N_4310);
and U7448 (N_7448,N_3953,N_2585);
or U7449 (N_7449,N_4032,N_3579);
nor U7450 (N_7450,N_4094,N_138);
nor U7451 (N_7451,N_1735,N_1038);
and U7452 (N_7452,N_1132,N_975);
nand U7453 (N_7453,N_256,N_491);
and U7454 (N_7454,N_4182,N_485);
and U7455 (N_7455,N_4434,N_3634);
xor U7456 (N_7456,N_3410,N_1651);
xnor U7457 (N_7457,N_1657,N_2749);
or U7458 (N_7458,N_4285,N_1752);
xnor U7459 (N_7459,N_948,N_3762);
nand U7460 (N_7460,N_3901,N_3886);
or U7461 (N_7461,N_3385,N_4754);
nand U7462 (N_7462,N_149,N_3300);
nor U7463 (N_7463,N_1843,N_2953);
and U7464 (N_7464,N_1184,N_2242);
nand U7465 (N_7465,N_2318,N_2971);
or U7466 (N_7466,N_114,N_4600);
nor U7467 (N_7467,N_679,N_2567);
nand U7468 (N_7468,N_1384,N_156);
or U7469 (N_7469,N_2771,N_3283);
and U7470 (N_7470,N_53,N_4756);
nand U7471 (N_7471,N_2908,N_1300);
nand U7472 (N_7472,N_2652,N_617);
and U7473 (N_7473,N_185,N_1731);
or U7474 (N_7474,N_2865,N_2259);
nand U7475 (N_7475,N_908,N_285);
nand U7476 (N_7476,N_1648,N_3485);
nor U7477 (N_7477,N_15,N_4478);
and U7478 (N_7478,N_2988,N_262);
nor U7479 (N_7479,N_1435,N_2475);
nand U7480 (N_7480,N_1609,N_4215);
and U7481 (N_7481,N_336,N_1324);
nor U7482 (N_7482,N_3884,N_582);
or U7483 (N_7483,N_3754,N_3915);
nand U7484 (N_7484,N_3533,N_510);
nand U7485 (N_7485,N_4935,N_1493);
nor U7486 (N_7486,N_4017,N_4042);
nor U7487 (N_7487,N_3350,N_4322);
nand U7488 (N_7488,N_1085,N_1944);
or U7489 (N_7489,N_266,N_4490);
or U7490 (N_7490,N_4227,N_2597);
nand U7491 (N_7491,N_3644,N_836);
or U7492 (N_7492,N_4886,N_283);
nor U7493 (N_7493,N_2745,N_2253);
nand U7494 (N_7494,N_2984,N_527);
xnor U7495 (N_7495,N_1529,N_4583);
and U7496 (N_7496,N_1374,N_711);
nand U7497 (N_7497,N_3258,N_4817);
nor U7498 (N_7498,N_1776,N_2772);
nand U7499 (N_7499,N_1170,N_3693);
or U7500 (N_7500,N_1788,N_3967);
nand U7501 (N_7501,N_4409,N_2952);
nor U7502 (N_7502,N_2702,N_4468);
nand U7503 (N_7503,N_1007,N_1652);
and U7504 (N_7504,N_629,N_1865);
nor U7505 (N_7505,N_1746,N_4654);
and U7506 (N_7506,N_3840,N_3692);
nand U7507 (N_7507,N_1930,N_960);
nand U7508 (N_7508,N_2641,N_1601);
nand U7509 (N_7509,N_3787,N_3133);
nand U7510 (N_7510,N_600,N_428);
nand U7511 (N_7511,N_3185,N_3755);
or U7512 (N_7512,N_4182,N_4432);
nor U7513 (N_7513,N_2477,N_4312);
nor U7514 (N_7514,N_234,N_1281);
nor U7515 (N_7515,N_2656,N_1373);
and U7516 (N_7516,N_3552,N_1748);
and U7517 (N_7517,N_210,N_4186);
and U7518 (N_7518,N_2461,N_1637);
and U7519 (N_7519,N_1102,N_3733);
or U7520 (N_7520,N_3489,N_2695);
nand U7521 (N_7521,N_2261,N_3085);
nand U7522 (N_7522,N_1143,N_133);
and U7523 (N_7523,N_1693,N_3906);
and U7524 (N_7524,N_4996,N_1056);
or U7525 (N_7525,N_700,N_2153);
or U7526 (N_7526,N_4257,N_676);
nand U7527 (N_7527,N_2693,N_1135);
nand U7528 (N_7528,N_1325,N_1660);
nand U7529 (N_7529,N_1229,N_777);
nand U7530 (N_7530,N_3598,N_705);
or U7531 (N_7531,N_1412,N_1301);
nor U7532 (N_7532,N_631,N_4649);
nand U7533 (N_7533,N_3250,N_3329);
nand U7534 (N_7534,N_1673,N_4892);
or U7535 (N_7535,N_1947,N_468);
and U7536 (N_7536,N_2168,N_1254);
nand U7537 (N_7537,N_4068,N_4519);
and U7538 (N_7538,N_461,N_4568);
nand U7539 (N_7539,N_1889,N_4679);
nor U7540 (N_7540,N_4754,N_1660);
or U7541 (N_7541,N_1794,N_4138);
and U7542 (N_7542,N_3431,N_1937);
nand U7543 (N_7543,N_3755,N_2095);
and U7544 (N_7544,N_1957,N_2049);
nand U7545 (N_7545,N_1119,N_1547);
or U7546 (N_7546,N_378,N_842);
nand U7547 (N_7547,N_4548,N_4416);
or U7548 (N_7548,N_544,N_4057);
or U7549 (N_7549,N_2230,N_3039);
nor U7550 (N_7550,N_2582,N_3700);
or U7551 (N_7551,N_1149,N_136);
nand U7552 (N_7552,N_3446,N_528);
or U7553 (N_7553,N_1569,N_3014);
nand U7554 (N_7554,N_4228,N_2885);
xor U7555 (N_7555,N_2563,N_1873);
nand U7556 (N_7556,N_4078,N_1334);
nand U7557 (N_7557,N_1526,N_451);
or U7558 (N_7558,N_4465,N_1541);
and U7559 (N_7559,N_3228,N_2);
and U7560 (N_7560,N_806,N_3730);
nand U7561 (N_7561,N_4110,N_1516);
or U7562 (N_7562,N_790,N_2755);
and U7563 (N_7563,N_3887,N_2474);
nor U7564 (N_7564,N_2282,N_2435);
nor U7565 (N_7565,N_4815,N_3431);
nand U7566 (N_7566,N_2521,N_2462);
or U7567 (N_7567,N_870,N_1186);
or U7568 (N_7568,N_2553,N_1099);
nor U7569 (N_7569,N_743,N_740);
or U7570 (N_7570,N_1111,N_1834);
nand U7571 (N_7571,N_1195,N_2984);
or U7572 (N_7572,N_2888,N_3368);
and U7573 (N_7573,N_64,N_1840);
or U7574 (N_7574,N_3417,N_4931);
and U7575 (N_7575,N_53,N_1132);
nor U7576 (N_7576,N_2392,N_2743);
xnor U7577 (N_7577,N_4916,N_2204);
and U7578 (N_7578,N_3891,N_4543);
xnor U7579 (N_7579,N_1560,N_2486);
and U7580 (N_7580,N_1859,N_3602);
and U7581 (N_7581,N_1615,N_750);
nor U7582 (N_7582,N_4339,N_3546);
or U7583 (N_7583,N_3761,N_2029);
xnor U7584 (N_7584,N_845,N_1308);
or U7585 (N_7585,N_3861,N_476);
nand U7586 (N_7586,N_1170,N_2079);
and U7587 (N_7587,N_302,N_3055);
nand U7588 (N_7588,N_2760,N_558);
nand U7589 (N_7589,N_1524,N_2139);
nand U7590 (N_7590,N_329,N_371);
or U7591 (N_7591,N_2542,N_4964);
and U7592 (N_7592,N_1753,N_90);
nand U7593 (N_7593,N_4762,N_4765);
or U7594 (N_7594,N_4017,N_3837);
nor U7595 (N_7595,N_113,N_851);
nor U7596 (N_7596,N_3495,N_3297);
or U7597 (N_7597,N_1021,N_3489);
or U7598 (N_7598,N_2589,N_4633);
or U7599 (N_7599,N_2427,N_4391);
nor U7600 (N_7600,N_2482,N_2026);
or U7601 (N_7601,N_2785,N_941);
or U7602 (N_7602,N_535,N_4972);
nand U7603 (N_7603,N_2819,N_3165);
or U7604 (N_7604,N_3702,N_1034);
nor U7605 (N_7605,N_3999,N_2344);
and U7606 (N_7606,N_1973,N_3527);
or U7607 (N_7607,N_668,N_4999);
nor U7608 (N_7608,N_2487,N_4549);
and U7609 (N_7609,N_2199,N_1254);
and U7610 (N_7610,N_2353,N_771);
nand U7611 (N_7611,N_823,N_3411);
or U7612 (N_7612,N_2335,N_985);
or U7613 (N_7613,N_35,N_1806);
or U7614 (N_7614,N_2161,N_3429);
or U7615 (N_7615,N_4799,N_4406);
or U7616 (N_7616,N_944,N_3263);
nand U7617 (N_7617,N_730,N_41);
nand U7618 (N_7618,N_1661,N_1857);
and U7619 (N_7619,N_2593,N_3057);
or U7620 (N_7620,N_4437,N_281);
and U7621 (N_7621,N_1331,N_672);
nor U7622 (N_7622,N_1226,N_1584);
and U7623 (N_7623,N_3653,N_647);
or U7624 (N_7624,N_3399,N_3484);
nor U7625 (N_7625,N_4935,N_3915);
or U7626 (N_7626,N_1074,N_4863);
or U7627 (N_7627,N_959,N_4983);
nand U7628 (N_7628,N_4637,N_3944);
or U7629 (N_7629,N_3711,N_1830);
nor U7630 (N_7630,N_4896,N_374);
or U7631 (N_7631,N_4273,N_1537);
or U7632 (N_7632,N_2063,N_889);
and U7633 (N_7633,N_2238,N_1705);
or U7634 (N_7634,N_849,N_3076);
nand U7635 (N_7635,N_2405,N_1622);
and U7636 (N_7636,N_4354,N_3040);
nor U7637 (N_7637,N_2164,N_3413);
nor U7638 (N_7638,N_1687,N_2761);
and U7639 (N_7639,N_1303,N_4072);
nand U7640 (N_7640,N_2288,N_2839);
nand U7641 (N_7641,N_1901,N_3218);
or U7642 (N_7642,N_83,N_4282);
or U7643 (N_7643,N_2578,N_2933);
and U7644 (N_7644,N_207,N_4929);
nand U7645 (N_7645,N_4253,N_1971);
nor U7646 (N_7646,N_2013,N_4346);
nor U7647 (N_7647,N_2774,N_3070);
or U7648 (N_7648,N_3246,N_2551);
and U7649 (N_7649,N_382,N_4279);
or U7650 (N_7650,N_3068,N_949);
and U7651 (N_7651,N_4072,N_144);
or U7652 (N_7652,N_1743,N_3870);
or U7653 (N_7653,N_2362,N_3921);
nand U7654 (N_7654,N_1257,N_999);
nor U7655 (N_7655,N_3726,N_2766);
nor U7656 (N_7656,N_3985,N_3186);
or U7657 (N_7657,N_2345,N_4514);
nand U7658 (N_7658,N_2475,N_3745);
and U7659 (N_7659,N_2749,N_1848);
nand U7660 (N_7660,N_2773,N_2559);
nor U7661 (N_7661,N_1103,N_4071);
nor U7662 (N_7662,N_4417,N_2143);
nor U7663 (N_7663,N_56,N_519);
xnor U7664 (N_7664,N_4935,N_2461);
or U7665 (N_7665,N_502,N_4892);
or U7666 (N_7666,N_130,N_3128);
nand U7667 (N_7667,N_508,N_4437);
and U7668 (N_7668,N_2251,N_2778);
nand U7669 (N_7669,N_580,N_805);
and U7670 (N_7670,N_4392,N_2013);
nor U7671 (N_7671,N_3316,N_3144);
nand U7672 (N_7672,N_1942,N_1978);
nor U7673 (N_7673,N_532,N_1476);
and U7674 (N_7674,N_4052,N_2546);
nor U7675 (N_7675,N_2258,N_4915);
or U7676 (N_7676,N_4841,N_3521);
and U7677 (N_7677,N_3788,N_1931);
nor U7678 (N_7678,N_3958,N_2334);
xnor U7679 (N_7679,N_2942,N_3994);
nor U7680 (N_7680,N_4256,N_4647);
nand U7681 (N_7681,N_3610,N_4900);
nand U7682 (N_7682,N_4153,N_3391);
nand U7683 (N_7683,N_358,N_4526);
and U7684 (N_7684,N_1125,N_2501);
nor U7685 (N_7685,N_3994,N_3481);
or U7686 (N_7686,N_1199,N_2225);
and U7687 (N_7687,N_1604,N_2413);
and U7688 (N_7688,N_298,N_1719);
and U7689 (N_7689,N_4945,N_191);
or U7690 (N_7690,N_1597,N_2279);
nor U7691 (N_7691,N_2007,N_1931);
or U7692 (N_7692,N_3881,N_4833);
and U7693 (N_7693,N_3627,N_2683);
nand U7694 (N_7694,N_2560,N_4373);
and U7695 (N_7695,N_421,N_4336);
nor U7696 (N_7696,N_4511,N_3231);
and U7697 (N_7697,N_423,N_4164);
and U7698 (N_7698,N_4428,N_3523);
nor U7699 (N_7699,N_3168,N_531);
or U7700 (N_7700,N_3977,N_3917);
nor U7701 (N_7701,N_302,N_2954);
nand U7702 (N_7702,N_4990,N_4601);
nor U7703 (N_7703,N_4649,N_2303);
or U7704 (N_7704,N_2545,N_1303);
and U7705 (N_7705,N_3710,N_3507);
nor U7706 (N_7706,N_3506,N_507);
nor U7707 (N_7707,N_3948,N_551);
nor U7708 (N_7708,N_4920,N_2904);
and U7709 (N_7709,N_1061,N_2030);
and U7710 (N_7710,N_4868,N_577);
or U7711 (N_7711,N_3301,N_4352);
and U7712 (N_7712,N_1337,N_3897);
nand U7713 (N_7713,N_691,N_1159);
nor U7714 (N_7714,N_1123,N_3042);
nor U7715 (N_7715,N_2129,N_1160);
nor U7716 (N_7716,N_3758,N_1104);
nand U7717 (N_7717,N_2740,N_2974);
and U7718 (N_7718,N_2433,N_115);
nor U7719 (N_7719,N_391,N_254);
nand U7720 (N_7720,N_1558,N_4690);
nor U7721 (N_7721,N_1035,N_347);
and U7722 (N_7722,N_1437,N_2602);
nor U7723 (N_7723,N_4,N_1159);
nor U7724 (N_7724,N_2574,N_4148);
xor U7725 (N_7725,N_3547,N_43);
or U7726 (N_7726,N_1137,N_3704);
or U7727 (N_7727,N_2846,N_1986);
and U7728 (N_7728,N_4720,N_2941);
nand U7729 (N_7729,N_4821,N_220);
and U7730 (N_7730,N_2837,N_3554);
or U7731 (N_7731,N_57,N_3936);
nand U7732 (N_7732,N_1279,N_2861);
nand U7733 (N_7733,N_4509,N_1510);
nor U7734 (N_7734,N_1411,N_1711);
nor U7735 (N_7735,N_2163,N_1168);
nor U7736 (N_7736,N_4594,N_2586);
nor U7737 (N_7737,N_648,N_4685);
or U7738 (N_7738,N_787,N_3546);
nor U7739 (N_7739,N_1769,N_2035);
and U7740 (N_7740,N_3521,N_4284);
and U7741 (N_7741,N_3851,N_1345);
nand U7742 (N_7742,N_2839,N_3769);
nor U7743 (N_7743,N_1083,N_3264);
or U7744 (N_7744,N_2909,N_1021);
or U7745 (N_7745,N_127,N_1451);
nand U7746 (N_7746,N_2308,N_336);
and U7747 (N_7747,N_1496,N_2574);
nand U7748 (N_7748,N_276,N_4175);
or U7749 (N_7749,N_2464,N_3600);
nand U7750 (N_7750,N_3479,N_4908);
nand U7751 (N_7751,N_1524,N_960);
nor U7752 (N_7752,N_4616,N_2597);
nand U7753 (N_7753,N_4032,N_4270);
and U7754 (N_7754,N_3098,N_2603);
and U7755 (N_7755,N_3789,N_4904);
or U7756 (N_7756,N_4147,N_98);
and U7757 (N_7757,N_1600,N_677);
nor U7758 (N_7758,N_3863,N_694);
and U7759 (N_7759,N_4504,N_2003);
or U7760 (N_7760,N_1347,N_2905);
nand U7761 (N_7761,N_856,N_4995);
nor U7762 (N_7762,N_2432,N_1263);
or U7763 (N_7763,N_4410,N_3226);
nor U7764 (N_7764,N_4933,N_456);
nor U7765 (N_7765,N_4006,N_2213);
or U7766 (N_7766,N_1856,N_1959);
nand U7767 (N_7767,N_1158,N_4111);
or U7768 (N_7768,N_1332,N_3661);
or U7769 (N_7769,N_2604,N_122);
and U7770 (N_7770,N_665,N_1131);
and U7771 (N_7771,N_79,N_898);
and U7772 (N_7772,N_4315,N_1585);
or U7773 (N_7773,N_3260,N_3698);
or U7774 (N_7774,N_3713,N_1014);
and U7775 (N_7775,N_521,N_4453);
nand U7776 (N_7776,N_173,N_3960);
nand U7777 (N_7777,N_1788,N_4294);
nor U7778 (N_7778,N_4064,N_4285);
nand U7779 (N_7779,N_4228,N_4293);
and U7780 (N_7780,N_4716,N_4739);
nand U7781 (N_7781,N_2696,N_339);
and U7782 (N_7782,N_2715,N_2513);
nand U7783 (N_7783,N_4857,N_3841);
or U7784 (N_7784,N_1037,N_1348);
xnor U7785 (N_7785,N_3849,N_3177);
xnor U7786 (N_7786,N_2012,N_2530);
xor U7787 (N_7787,N_2053,N_3757);
nand U7788 (N_7788,N_3359,N_127);
nand U7789 (N_7789,N_143,N_2433);
and U7790 (N_7790,N_2760,N_1444);
nand U7791 (N_7791,N_3373,N_2559);
nor U7792 (N_7792,N_3369,N_4384);
and U7793 (N_7793,N_4768,N_2025);
and U7794 (N_7794,N_2120,N_4719);
nand U7795 (N_7795,N_4304,N_192);
nand U7796 (N_7796,N_4379,N_4544);
nand U7797 (N_7797,N_2135,N_641);
and U7798 (N_7798,N_1823,N_182);
and U7799 (N_7799,N_400,N_3283);
nor U7800 (N_7800,N_3997,N_4505);
nor U7801 (N_7801,N_2862,N_2296);
and U7802 (N_7802,N_2992,N_242);
nor U7803 (N_7803,N_106,N_183);
and U7804 (N_7804,N_4221,N_3438);
nor U7805 (N_7805,N_4605,N_4630);
or U7806 (N_7806,N_3160,N_367);
nor U7807 (N_7807,N_1472,N_3177);
nand U7808 (N_7808,N_4572,N_4749);
nor U7809 (N_7809,N_1102,N_4176);
nor U7810 (N_7810,N_4835,N_8);
or U7811 (N_7811,N_233,N_3171);
xnor U7812 (N_7812,N_2977,N_1505);
nand U7813 (N_7813,N_4049,N_3999);
or U7814 (N_7814,N_4091,N_2269);
or U7815 (N_7815,N_3427,N_4111);
or U7816 (N_7816,N_2376,N_1715);
and U7817 (N_7817,N_1929,N_4559);
or U7818 (N_7818,N_175,N_4477);
nand U7819 (N_7819,N_725,N_3806);
or U7820 (N_7820,N_3629,N_3525);
or U7821 (N_7821,N_138,N_1688);
or U7822 (N_7822,N_1103,N_3011);
nor U7823 (N_7823,N_3593,N_4693);
and U7824 (N_7824,N_375,N_2440);
and U7825 (N_7825,N_4264,N_3995);
or U7826 (N_7826,N_2412,N_1535);
nand U7827 (N_7827,N_4049,N_711);
nand U7828 (N_7828,N_1789,N_4425);
and U7829 (N_7829,N_2051,N_2524);
xnor U7830 (N_7830,N_1408,N_4326);
and U7831 (N_7831,N_771,N_729);
nor U7832 (N_7832,N_2886,N_3122);
nand U7833 (N_7833,N_4785,N_1033);
nor U7834 (N_7834,N_735,N_2032);
or U7835 (N_7835,N_2188,N_3306);
or U7836 (N_7836,N_4117,N_880);
or U7837 (N_7837,N_4086,N_738);
or U7838 (N_7838,N_2344,N_974);
nor U7839 (N_7839,N_3080,N_3487);
or U7840 (N_7840,N_1458,N_2997);
and U7841 (N_7841,N_3582,N_2028);
nor U7842 (N_7842,N_3274,N_4515);
nor U7843 (N_7843,N_1977,N_3359);
and U7844 (N_7844,N_1497,N_2812);
or U7845 (N_7845,N_161,N_1564);
nand U7846 (N_7846,N_4722,N_2816);
or U7847 (N_7847,N_744,N_4399);
and U7848 (N_7848,N_1849,N_4309);
nor U7849 (N_7849,N_4828,N_2595);
or U7850 (N_7850,N_4941,N_3591);
or U7851 (N_7851,N_2152,N_3501);
or U7852 (N_7852,N_4099,N_1449);
nor U7853 (N_7853,N_1806,N_4210);
nand U7854 (N_7854,N_2912,N_4042);
or U7855 (N_7855,N_1465,N_2282);
and U7856 (N_7856,N_995,N_907);
nor U7857 (N_7857,N_1771,N_85);
nand U7858 (N_7858,N_216,N_3856);
and U7859 (N_7859,N_4799,N_1137);
and U7860 (N_7860,N_833,N_600);
or U7861 (N_7861,N_4523,N_3890);
and U7862 (N_7862,N_4680,N_2418);
nand U7863 (N_7863,N_432,N_3207);
nand U7864 (N_7864,N_1106,N_3241);
nand U7865 (N_7865,N_679,N_1740);
nand U7866 (N_7866,N_808,N_1021);
or U7867 (N_7867,N_3953,N_1597);
nor U7868 (N_7868,N_3431,N_2176);
nor U7869 (N_7869,N_4946,N_3038);
and U7870 (N_7870,N_3979,N_3431);
nor U7871 (N_7871,N_3495,N_2201);
or U7872 (N_7872,N_875,N_1726);
nor U7873 (N_7873,N_1402,N_4242);
nor U7874 (N_7874,N_4559,N_4703);
or U7875 (N_7875,N_262,N_228);
nand U7876 (N_7876,N_2657,N_4724);
or U7877 (N_7877,N_4005,N_4722);
nor U7878 (N_7878,N_3587,N_2306);
or U7879 (N_7879,N_2341,N_2171);
nor U7880 (N_7880,N_1129,N_3922);
nand U7881 (N_7881,N_401,N_2462);
nand U7882 (N_7882,N_2578,N_97);
or U7883 (N_7883,N_1567,N_652);
or U7884 (N_7884,N_853,N_674);
and U7885 (N_7885,N_4634,N_45);
nor U7886 (N_7886,N_560,N_4295);
nand U7887 (N_7887,N_2062,N_1641);
nand U7888 (N_7888,N_4265,N_4523);
nor U7889 (N_7889,N_1819,N_4456);
xnor U7890 (N_7890,N_3892,N_3467);
nand U7891 (N_7891,N_3450,N_874);
nand U7892 (N_7892,N_4020,N_2591);
nor U7893 (N_7893,N_1015,N_2516);
xnor U7894 (N_7894,N_23,N_3885);
or U7895 (N_7895,N_3822,N_4488);
nor U7896 (N_7896,N_199,N_4493);
nand U7897 (N_7897,N_2549,N_3357);
xor U7898 (N_7898,N_2088,N_2717);
nor U7899 (N_7899,N_4654,N_672);
and U7900 (N_7900,N_1332,N_4734);
or U7901 (N_7901,N_44,N_235);
and U7902 (N_7902,N_1016,N_608);
and U7903 (N_7903,N_3753,N_1847);
nor U7904 (N_7904,N_2503,N_3399);
nand U7905 (N_7905,N_1754,N_2655);
nor U7906 (N_7906,N_2658,N_2619);
nor U7907 (N_7907,N_2408,N_3717);
nor U7908 (N_7908,N_201,N_1708);
and U7909 (N_7909,N_709,N_4007);
or U7910 (N_7910,N_3238,N_961);
or U7911 (N_7911,N_2035,N_3878);
or U7912 (N_7912,N_985,N_1079);
xnor U7913 (N_7913,N_1632,N_4933);
or U7914 (N_7914,N_583,N_4632);
nand U7915 (N_7915,N_1098,N_956);
or U7916 (N_7916,N_3438,N_2076);
and U7917 (N_7917,N_4463,N_1348);
and U7918 (N_7918,N_3650,N_4380);
nand U7919 (N_7919,N_4607,N_1508);
nor U7920 (N_7920,N_2920,N_2922);
nand U7921 (N_7921,N_3200,N_1022);
or U7922 (N_7922,N_2494,N_3060);
or U7923 (N_7923,N_2840,N_3809);
or U7924 (N_7924,N_3590,N_3764);
nor U7925 (N_7925,N_3576,N_4044);
nand U7926 (N_7926,N_3665,N_1964);
nand U7927 (N_7927,N_2988,N_4520);
xnor U7928 (N_7928,N_4061,N_1792);
nor U7929 (N_7929,N_395,N_1559);
and U7930 (N_7930,N_689,N_2138);
and U7931 (N_7931,N_2422,N_402);
nor U7932 (N_7932,N_2656,N_3988);
nor U7933 (N_7933,N_366,N_909);
and U7934 (N_7934,N_392,N_1989);
and U7935 (N_7935,N_717,N_1449);
or U7936 (N_7936,N_2469,N_1887);
xnor U7937 (N_7937,N_2305,N_1317);
or U7938 (N_7938,N_801,N_4965);
and U7939 (N_7939,N_1757,N_3508);
xnor U7940 (N_7940,N_730,N_1617);
and U7941 (N_7941,N_2997,N_3334);
and U7942 (N_7942,N_915,N_840);
or U7943 (N_7943,N_2384,N_278);
nand U7944 (N_7944,N_892,N_2736);
or U7945 (N_7945,N_2209,N_4895);
and U7946 (N_7946,N_363,N_4189);
and U7947 (N_7947,N_58,N_1862);
or U7948 (N_7948,N_1173,N_2516);
or U7949 (N_7949,N_3703,N_2222);
or U7950 (N_7950,N_2637,N_4415);
or U7951 (N_7951,N_586,N_996);
or U7952 (N_7952,N_2813,N_1107);
nand U7953 (N_7953,N_2579,N_2783);
and U7954 (N_7954,N_44,N_93);
or U7955 (N_7955,N_3185,N_1379);
or U7956 (N_7956,N_2779,N_1802);
nand U7957 (N_7957,N_51,N_1274);
or U7958 (N_7958,N_1742,N_2160);
nor U7959 (N_7959,N_948,N_1317);
nand U7960 (N_7960,N_4724,N_4564);
or U7961 (N_7961,N_3125,N_942);
nand U7962 (N_7962,N_1105,N_4314);
or U7963 (N_7963,N_4808,N_3788);
nand U7964 (N_7964,N_4156,N_2191);
nor U7965 (N_7965,N_3208,N_123);
or U7966 (N_7966,N_3120,N_2788);
and U7967 (N_7967,N_646,N_2565);
or U7968 (N_7968,N_4011,N_4424);
nor U7969 (N_7969,N_3065,N_2165);
and U7970 (N_7970,N_3268,N_4598);
and U7971 (N_7971,N_1159,N_1692);
nor U7972 (N_7972,N_4174,N_1193);
and U7973 (N_7973,N_1661,N_3996);
and U7974 (N_7974,N_2335,N_1944);
or U7975 (N_7975,N_1886,N_3164);
nor U7976 (N_7976,N_38,N_1340);
or U7977 (N_7977,N_4550,N_1325);
nor U7978 (N_7978,N_3910,N_1813);
or U7979 (N_7979,N_3709,N_3070);
or U7980 (N_7980,N_437,N_6);
xor U7981 (N_7981,N_3468,N_1645);
or U7982 (N_7982,N_1240,N_1237);
nand U7983 (N_7983,N_4728,N_911);
nand U7984 (N_7984,N_3505,N_1654);
nand U7985 (N_7985,N_3059,N_1274);
nor U7986 (N_7986,N_3413,N_773);
nand U7987 (N_7987,N_4438,N_407);
xor U7988 (N_7988,N_251,N_2447);
nor U7989 (N_7989,N_2800,N_2070);
or U7990 (N_7990,N_3540,N_3189);
nor U7991 (N_7991,N_1813,N_2634);
and U7992 (N_7992,N_4254,N_220);
nand U7993 (N_7993,N_2499,N_3375);
or U7994 (N_7994,N_3332,N_4496);
and U7995 (N_7995,N_3376,N_646);
and U7996 (N_7996,N_4134,N_1818);
nand U7997 (N_7997,N_4009,N_4523);
or U7998 (N_7998,N_3773,N_4343);
or U7999 (N_7999,N_1579,N_3232);
or U8000 (N_8000,N_4299,N_4971);
nor U8001 (N_8001,N_700,N_4241);
nand U8002 (N_8002,N_1617,N_1219);
nor U8003 (N_8003,N_3805,N_4155);
nor U8004 (N_8004,N_3449,N_2761);
and U8005 (N_8005,N_4263,N_4471);
nor U8006 (N_8006,N_402,N_3857);
or U8007 (N_8007,N_532,N_769);
nand U8008 (N_8008,N_456,N_366);
or U8009 (N_8009,N_1744,N_1644);
or U8010 (N_8010,N_3359,N_2223);
nor U8011 (N_8011,N_2400,N_1548);
nor U8012 (N_8012,N_4913,N_914);
and U8013 (N_8013,N_1139,N_2627);
nand U8014 (N_8014,N_544,N_2136);
nand U8015 (N_8015,N_396,N_3792);
nor U8016 (N_8016,N_2895,N_2777);
nor U8017 (N_8017,N_3238,N_3347);
xnor U8018 (N_8018,N_3681,N_415);
and U8019 (N_8019,N_4029,N_2301);
nor U8020 (N_8020,N_112,N_4638);
or U8021 (N_8021,N_815,N_4960);
nand U8022 (N_8022,N_1086,N_209);
and U8023 (N_8023,N_4304,N_2937);
nand U8024 (N_8024,N_1839,N_1713);
nand U8025 (N_8025,N_1976,N_4171);
nor U8026 (N_8026,N_2175,N_1995);
and U8027 (N_8027,N_1375,N_2267);
or U8028 (N_8028,N_4523,N_955);
nor U8029 (N_8029,N_2248,N_3611);
or U8030 (N_8030,N_3510,N_3363);
or U8031 (N_8031,N_2874,N_2909);
and U8032 (N_8032,N_1695,N_206);
or U8033 (N_8033,N_2804,N_1709);
nor U8034 (N_8034,N_4196,N_516);
nand U8035 (N_8035,N_2094,N_1728);
nand U8036 (N_8036,N_1735,N_3011);
or U8037 (N_8037,N_1710,N_3643);
and U8038 (N_8038,N_271,N_1503);
and U8039 (N_8039,N_792,N_4700);
nand U8040 (N_8040,N_2189,N_4013);
and U8041 (N_8041,N_3344,N_3188);
and U8042 (N_8042,N_2615,N_1946);
nand U8043 (N_8043,N_4187,N_3918);
nor U8044 (N_8044,N_2984,N_4906);
and U8045 (N_8045,N_3613,N_1381);
and U8046 (N_8046,N_789,N_2830);
nor U8047 (N_8047,N_2357,N_1151);
nand U8048 (N_8048,N_2927,N_150);
and U8049 (N_8049,N_16,N_349);
or U8050 (N_8050,N_2909,N_2753);
or U8051 (N_8051,N_2422,N_2941);
nand U8052 (N_8052,N_1209,N_632);
and U8053 (N_8053,N_1091,N_2708);
nor U8054 (N_8054,N_3129,N_4940);
nand U8055 (N_8055,N_1856,N_1302);
or U8056 (N_8056,N_3700,N_3581);
and U8057 (N_8057,N_3269,N_3170);
or U8058 (N_8058,N_1790,N_1666);
nor U8059 (N_8059,N_448,N_2762);
nor U8060 (N_8060,N_1445,N_87);
and U8061 (N_8061,N_1551,N_4549);
and U8062 (N_8062,N_1117,N_1065);
and U8063 (N_8063,N_4566,N_2769);
and U8064 (N_8064,N_3940,N_555);
nor U8065 (N_8065,N_2615,N_2239);
nand U8066 (N_8066,N_1691,N_4614);
and U8067 (N_8067,N_2995,N_3675);
nand U8068 (N_8068,N_2040,N_2218);
nand U8069 (N_8069,N_181,N_4223);
or U8070 (N_8070,N_1250,N_766);
nor U8071 (N_8071,N_2752,N_93);
or U8072 (N_8072,N_806,N_3642);
or U8073 (N_8073,N_3870,N_3002);
nand U8074 (N_8074,N_1742,N_4408);
nand U8075 (N_8075,N_4803,N_1960);
and U8076 (N_8076,N_1039,N_2067);
xnor U8077 (N_8077,N_1292,N_3);
or U8078 (N_8078,N_997,N_3566);
nand U8079 (N_8079,N_2564,N_2099);
and U8080 (N_8080,N_1805,N_3079);
nand U8081 (N_8081,N_517,N_175);
xnor U8082 (N_8082,N_501,N_686);
nand U8083 (N_8083,N_3475,N_2146);
nand U8084 (N_8084,N_4374,N_2908);
or U8085 (N_8085,N_486,N_3831);
nor U8086 (N_8086,N_3198,N_3385);
nand U8087 (N_8087,N_57,N_4986);
or U8088 (N_8088,N_4508,N_3020);
and U8089 (N_8089,N_1942,N_3864);
or U8090 (N_8090,N_3873,N_4746);
and U8091 (N_8091,N_2478,N_131);
nand U8092 (N_8092,N_2053,N_3790);
nor U8093 (N_8093,N_1534,N_1381);
nand U8094 (N_8094,N_4556,N_3135);
and U8095 (N_8095,N_617,N_2054);
and U8096 (N_8096,N_3896,N_4489);
nor U8097 (N_8097,N_4778,N_4493);
nor U8098 (N_8098,N_2666,N_662);
nand U8099 (N_8099,N_1425,N_1511);
nand U8100 (N_8100,N_2227,N_1571);
or U8101 (N_8101,N_2947,N_4317);
nor U8102 (N_8102,N_650,N_3737);
nor U8103 (N_8103,N_94,N_4165);
or U8104 (N_8104,N_385,N_3790);
nand U8105 (N_8105,N_2088,N_2471);
or U8106 (N_8106,N_3799,N_4630);
or U8107 (N_8107,N_415,N_2879);
nor U8108 (N_8108,N_679,N_4977);
and U8109 (N_8109,N_4655,N_406);
or U8110 (N_8110,N_4591,N_1330);
nand U8111 (N_8111,N_1724,N_3645);
nand U8112 (N_8112,N_3595,N_3899);
nor U8113 (N_8113,N_4871,N_293);
or U8114 (N_8114,N_1037,N_943);
nand U8115 (N_8115,N_4467,N_4623);
or U8116 (N_8116,N_3131,N_4748);
and U8117 (N_8117,N_860,N_598);
nor U8118 (N_8118,N_1201,N_48);
or U8119 (N_8119,N_2204,N_2746);
nor U8120 (N_8120,N_1035,N_3782);
and U8121 (N_8121,N_2285,N_2716);
nand U8122 (N_8122,N_1329,N_4374);
nand U8123 (N_8123,N_3678,N_2665);
nor U8124 (N_8124,N_200,N_2943);
and U8125 (N_8125,N_4434,N_2631);
nor U8126 (N_8126,N_14,N_2656);
nand U8127 (N_8127,N_3125,N_2937);
nand U8128 (N_8128,N_2631,N_3987);
or U8129 (N_8129,N_1359,N_976);
or U8130 (N_8130,N_2333,N_4519);
nor U8131 (N_8131,N_3117,N_3309);
xor U8132 (N_8132,N_1721,N_4942);
or U8133 (N_8133,N_1505,N_1591);
xor U8134 (N_8134,N_2040,N_1961);
and U8135 (N_8135,N_1037,N_1679);
nor U8136 (N_8136,N_1068,N_2553);
nand U8137 (N_8137,N_299,N_3327);
and U8138 (N_8138,N_1620,N_2239);
or U8139 (N_8139,N_4905,N_4065);
and U8140 (N_8140,N_4508,N_4737);
and U8141 (N_8141,N_3406,N_840);
nor U8142 (N_8142,N_4451,N_3664);
nor U8143 (N_8143,N_339,N_1750);
nor U8144 (N_8144,N_4717,N_2124);
or U8145 (N_8145,N_1626,N_2554);
nor U8146 (N_8146,N_3423,N_4653);
nor U8147 (N_8147,N_808,N_61);
nand U8148 (N_8148,N_1735,N_2699);
and U8149 (N_8149,N_1960,N_2769);
and U8150 (N_8150,N_183,N_3973);
nand U8151 (N_8151,N_4282,N_205);
and U8152 (N_8152,N_3864,N_2479);
and U8153 (N_8153,N_2358,N_1402);
or U8154 (N_8154,N_132,N_1522);
and U8155 (N_8155,N_2444,N_1751);
and U8156 (N_8156,N_1159,N_4797);
nand U8157 (N_8157,N_2495,N_1561);
and U8158 (N_8158,N_2167,N_3727);
nand U8159 (N_8159,N_3635,N_3494);
and U8160 (N_8160,N_859,N_3425);
or U8161 (N_8161,N_2452,N_4224);
or U8162 (N_8162,N_577,N_4263);
or U8163 (N_8163,N_486,N_918);
nand U8164 (N_8164,N_662,N_3316);
nand U8165 (N_8165,N_1268,N_2819);
or U8166 (N_8166,N_4424,N_1876);
or U8167 (N_8167,N_2343,N_2995);
and U8168 (N_8168,N_4490,N_1133);
and U8169 (N_8169,N_4069,N_4550);
or U8170 (N_8170,N_4206,N_4828);
and U8171 (N_8171,N_583,N_3560);
nor U8172 (N_8172,N_4164,N_2372);
or U8173 (N_8173,N_2713,N_3072);
nor U8174 (N_8174,N_2392,N_1701);
nand U8175 (N_8175,N_1798,N_479);
or U8176 (N_8176,N_2669,N_1444);
or U8177 (N_8177,N_1039,N_172);
and U8178 (N_8178,N_2874,N_3489);
and U8179 (N_8179,N_4339,N_452);
or U8180 (N_8180,N_3302,N_453);
or U8181 (N_8181,N_3652,N_1796);
and U8182 (N_8182,N_1466,N_3757);
nor U8183 (N_8183,N_1604,N_4696);
nand U8184 (N_8184,N_3044,N_1836);
and U8185 (N_8185,N_332,N_3978);
or U8186 (N_8186,N_923,N_794);
nor U8187 (N_8187,N_2780,N_1108);
or U8188 (N_8188,N_809,N_2008);
and U8189 (N_8189,N_3537,N_1173);
nor U8190 (N_8190,N_2681,N_1790);
nor U8191 (N_8191,N_3303,N_4204);
nand U8192 (N_8192,N_3413,N_922);
nor U8193 (N_8193,N_2288,N_3322);
or U8194 (N_8194,N_1336,N_1124);
nor U8195 (N_8195,N_534,N_435);
xor U8196 (N_8196,N_2359,N_2704);
or U8197 (N_8197,N_4450,N_1833);
nand U8198 (N_8198,N_1816,N_3562);
nand U8199 (N_8199,N_4874,N_283);
nand U8200 (N_8200,N_4339,N_1744);
or U8201 (N_8201,N_4175,N_1871);
nor U8202 (N_8202,N_1389,N_1526);
nand U8203 (N_8203,N_2794,N_3666);
and U8204 (N_8204,N_3562,N_822);
xor U8205 (N_8205,N_3832,N_373);
nor U8206 (N_8206,N_1863,N_1510);
and U8207 (N_8207,N_2470,N_4784);
and U8208 (N_8208,N_290,N_2693);
or U8209 (N_8209,N_3242,N_1296);
and U8210 (N_8210,N_2120,N_1075);
nand U8211 (N_8211,N_1844,N_1787);
nor U8212 (N_8212,N_4115,N_621);
or U8213 (N_8213,N_3039,N_3167);
or U8214 (N_8214,N_3283,N_4652);
and U8215 (N_8215,N_2284,N_991);
or U8216 (N_8216,N_3830,N_3608);
or U8217 (N_8217,N_3772,N_1337);
nor U8218 (N_8218,N_405,N_2021);
and U8219 (N_8219,N_1655,N_4264);
nand U8220 (N_8220,N_4265,N_220);
nand U8221 (N_8221,N_4652,N_1618);
or U8222 (N_8222,N_4075,N_4689);
or U8223 (N_8223,N_1884,N_3500);
nand U8224 (N_8224,N_4730,N_3462);
or U8225 (N_8225,N_2428,N_2389);
nor U8226 (N_8226,N_4934,N_349);
or U8227 (N_8227,N_4746,N_3102);
nand U8228 (N_8228,N_2679,N_2064);
or U8229 (N_8229,N_887,N_800);
nand U8230 (N_8230,N_4302,N_2187);
and U8231 (N_8231,N_782,N_3367);
nor U8232 (N_8232,N_707,N_762);
nor U8233 (N_8233,N_142,N_4241);
nor U8234 (N_8234,N_3402,N_4672);
nand U8235 (N_8235,N_3835,N_2980);
nor U8236 (N_8236,N_4608,N_2774);
nand U8237 (N_8237,N_244,N_3722);
and U8238 (N_8238,N_708,N_2093);
xnor U8239 (N_8239,N_822,N_2986);
and U8240 (N_8240,N_4097,N_2573);
or U8241 (N_8241,N_292,N_3902);
nand U8242 (N_8242,N_3307,N_3494);
and U8243 (N_8243,N_2848,N_4826);
nand U8244 (N_8244,N_3545,N_3682);
xnor U8245 (N_8245,N_3212,N_3101);
and U8246 (N_8246,N_3143,N_2753);
nor U8247 (N_8247,N_855,N_1536);
and U8248 (N_8248,N_9,N_218);
nand U8249 (N_8249,N_2134,N_945);
or U8250 (N_8250,N_1495,N_2636);
nor U8251 (N_8251,N_3902,N_4325);
nand U8252 (N_8252,N_3774,N_4297);
nor U8253 (N_8253,N_4880,N_681);
or U8254 (N_8254,N_2248,N_1188);
and U8255 (N_8255,N_2338,N_2316);
nor U8256 (N_8256,N_1670,N_2811);
nand U8257 (N_8257,N_4446,N_3305);
or U8258 (N_8258,N_1523,N_2512);
nor U8259 (N_8259,N_4855,N_1700);
nand U8260 (N_8260,N_3461,N_3544);
nor U8261 (N_8261,N_227,N_1055);
and U8262 (N_8262,N_4745,N_1461);
nor U8263 (N_8263,N_92,N_3123);
nor U8264 (N_8264,N_1248,N_3856);
nor U8265 (N_8265,N_3432,N_1502);
nand U8266 (N_8266,N_2914,N_3639);
and U8267 (N_8267,N_2472,N_718);
or U8268 (N_8268,N_582,N_4511);
and U8269 (N_8269,N_422,N_4023);
or U8270 (N_8270,N_4454,N_1050);
and U8271 (N_8271,N_4622,N_4201);
nand U8272 (N_8272,N_1073,N_2105);
nor U8273 (N_8273,N_4597,N_876);
nor U8274 (N_8274,N_3563,N_363);
and U8275 (N_8275,N_2105,N_1440);
and U8276 (N_8276,N_3682,N_1110);
nand U8277 (N_8277,N_1730,N_39);
nand U8278 (N_8278,N_190,N_958);
or U8279 (N_8279,N_1517,N_1634);
or U8280 (N_8280,N_3853,N_258);
nor U8281 (N_8281,N_719,N_2887);
nor U8282 (N_8282,N_1021,N_297);
nor U8283 (N_8283,N_1392,N_4207);
and U8284 (N_8284,N_2794,N_1869);
nand U8285 (N_8285,N_4427,N_4025);
or U8286 (N_8286,N_1147,N_2857);
nor U8287 (N_8287,N_3984,N_4335);
nand U8288 (N_8288,N_3236,N_3963);
nand U8289 (N_8289,N_1017,N_3491);
or U8290 (N_8290,N_2256,N_3292);
and U8291 (N_8291,N_3767,N_1032);
nor U8292 (N_8292,N_4848,N_2466);
nand U8293 (N_8293,N_4555,N_1935);
nor U8294 (N_8294,N_3427,N_4443);
or U8295 (N_8295,N_584,N_3997);
nand U8296 (N_8296,N_2687,N_2202);
or U8297 (N_8297,N_1288,N_2593);
nor U8298 (N_8298,N_1102,N_1428);
or U8299 (N_8299,N_2452,N_3101);
or U8300 (N_8300,N_1996,N_315);
and U8301 (N_8301,N_506,N_1851);
nor U8302 (N_8302,N_3398,N_3211);
or U8303 (N_8303,N_1109,N_2945);
nand U8304 (N_8304,N_4464,N_3961);
nand U8305 (N_8305,N_3560,N_154);
nor U8306 (N_8306,N_837,N_1644);
nor U8307 (N_8307,N_925,N_3197);
or U8308 (N_8308,N_4004,N_77);
and U8309 (N_8309,N_1748,N_2977);
nor U8310 (N_8310,N_1205,N_1257);
and U8311 (N_8311,N_2192,N_3772);
or U8312 (N_8312,N_1952,N_1751);
and U8313 (N_8313,N_6,N_2956);
nand U8314 (N_8314,N_2989,N_1875);
or U8315 (N_8315,N_2366,N_3791);
or U8316 (N_8316,N_3691,N_2600);
and U8317 (N_8317,N_135,N_3769);
and U8318 (N_8318,N_769,N_300);
nand U8319 (N_8319,N_211,N_4533);
and U8320 (N_8320,N_750,N_1679);
and U8321 (N_8321,N_4360,N_1289);
or U8322 (N_8322,N_1134,N_261);
nor U8323 (N_8323,N_645,N_2474);
nand U8324 (N_8324,N_856,N_4585);
nand U8325 (N_8325,N_2078,N_526);
and U8326 (N_8326,N_1497,N_4896);
nor U8327 (N_8327,N_3252,N_1656);
nand U8328 (N_8328,N_3639,N_2699);
nand U8329 (N_8329,N_3653,N_3189);
or U8330 (N_8330,N_4929,N_4990);
and U8331 (N_8331,N_265,N_3606);
nand U8332 (N_8332,N_2764,N_4423);
nand U8333 (N_8333,N_97,N_2742);
or U8334 (N_8334,N_978,N_2509);
or U8335 (N_8335,N_4321,N_1116);
and U8336 (N_8336,N_3090,N_1257);
nor U8337 (N_8337,N_2220,N_4275);
or U8338 (N_8338,N_697,N_2119);
and U8339 (N_8339,N_1800,N_3603);
and U8340 (N_8340,N_1352,N_1901);
or U8341 (N_8341,N_1276,N_1061);
nor U8342 (N_8342,N_1831,N_606);
and U8343 (N_8343,N_4018,N_801);
or U8344 (N_8344,N_1257,N_2945);
and U8345 (N_8345,N_1823,N_41);
or U8346 (N_8346,N_2660,N_1317);
xnor U8347 (N_8347,N_1866,N_1183);
or U8348 (N_8348,N_2702,N_2450);
or U8349 (N_8349,N_3568,N_2576);
nor U8350 (N_8350,N_1566,N_2496);
and U8351 (N_8351,N_4675,N_3476);
or U8352 (N_8352,N_4299,N_3201);
and U8353 (N_8353,N_342,N_2143);
and U8354 (N_8354,N_1102,N_3494);
and U8355 (N_8355,N_858,N_556);
and U8356 (N_8356,N_2531,N_1919);
nand U8357 (N_8357,N_298,N_2725);
nor U8358 (N_8358,N_3084,N_4845);
nor U8359 (N_8359,N_3833,N_1626);
nor U8360 (N_8360,N_1105,N_964);
nor U8361 (N_8361,N_3911,N_770);
and U8362 (N_8362,N_4778,N_1404);
or U8363 (N_8363,N_3034,N_1605);
nor U8364 (N_8364,N_2092,N_1495);
and U8365 (N_8365,N_2319,N_3832);
nor U8366 (N_8366,N_1374,N_3556);
or U8367 (N_8367,N_1887,N_492);
nand U8368 (N_8368,N_1167,N_695);
nand U8369 (N_8369,N_4764,N_4684);
and U8370 (N_8370,N_2301,N_1260);
nand U8371 (N_8371,N_3442,N_877);
nand U8372 (N_8372,N_4574,N_4705);
nor U8373 (N_8373,N_4953,N_2121);
nand U8374 (N_8374,N_4263,N_3983);
xnor U8375 (N_8375,N_2489,N_321);
xor U8376 (N_8376,N_3072,N_3484);
nor U8377 (N_8377,N_2051,N_4851);
and U8378 (N_8378,N_1522,N_2983);
nor U8379 (N_8379,N_2313,N_1561);
nor U8380 (N_8380,N_682,N_1732);
nand U8381 (N_8381,N_1897,N_1943);
and U8382 (N_8382,N_4616,N_442);
and U8383 (N_8383,N_1850,N_4766);
nor U8384 (N_8384,N_2557,N_3973);
and U8385 (N_8385,N_128,N_283);
or U8386 (N_8386,N_1929,N_2128);
and U8387 (N_8387,N_550,N_78);
and U8388 (N_8388,N_1127,N_426);
nand U8389 (N_8389,N_2927,N_3276);
nand U8390 (N_8390,N_3876,N_789);
xnor U8391 (N_8391,N_3650,N_3435);
xor U8392 (N_8392,N_1891,N_833);
and U8393 (N_8393,N_3480,N_4810);
or U8394 (N_8394,N_2982,N_4183);
or U8395 (N_8395,N_4245,N_4240);
and U8396 (N_8396,N_2209,N_1468);
and U8397 (N_8397,N_23,N_197);
or U8398 (N_8398,N_478,N_883);
nand U8399 (N_8399,N_4268,N_3904);
nand U8400 (N_8400,N_280,N_4243);
nor U8401 (N_8401,N_256,N_3768);
and U8402 (N_8402,N_320,N_4560);
nand U8403 (N_8403,N_3992,N_525);
nand U8404 (N_8404,N_2592,N_1992);
and U8405 (N_8405,N_1529,N_2082);
nor U8406 (N_8406,N_1474,N_4490);
nand U8407 (N_8407,N_4006,N_757);
nor U8408 (N_8408,N_4197,N_438);
or U8409 (N_8409,N_1488,N_320);
and U8410 (N_8410,N_2178,N_212);
and U8411 (N_8411,N_485,N_1201);
and U8412 (N_8412,N_1126,N_216);
or U8413 (N_8413,N_987,N_4163);
or U8414 (N_8414,N_200,N_466);
and U8415 (N_8415,N_3471,N_2329);
and U8416 (N_8416,N_3216,N_4600);
or U8417 (N_8417,N_2476,N_4288);
nor U8418 (N_8418,N_4769,N_3558);
nor U8419 (N_8419,N_2945,N_832);
or U8420 (N_8420,N_4375,N_1872);
nor U8421 (N_8421,N_4326,N_2287);
or U8422 (N_8422,N_3763,N_153);
and U8423 (N_8423,N_4129,N_2741);
and U8424 (N_8424,N_3037,N_2147);
nand U8425 (N_8425,N_3107,N_4160);
or U8426 (N_8426,N_3615,N_3159);
nor U8427 (N_8427,N_2556,N_1926);
nand U8428 (N_8428,N_988,N_4910);
nor U8429 (N_8429,N_2299,N_1983);
or U8430 (N_8430,N_2076,N_2138);
nand U8431 (N_8431,N_499,N_606);
or U8432 (N_8432,N_2850,N_4098);
nor U8433 (N_8433,N_1767,N_4964);
and U8434 (N_8434,N_2134,N_4502);
or U8435 (N_8435,N_1018,N_4773);
nor U8436 (N_8436,N_1081,N_4799);
or U8437 (N_8437,N_1585,N_3208);
and U8438 (N_8438,N_3623,N_4364);
and U8439 (N_8439,N_3596,N_1373);
nor U8440 (N_8440,N_2057,N_4577);
nor U8441 (N_8441,N_2294,N_4844);
nor U8442 (N_8442,N_451,N_3465);
nand U8443 (N_8443,N_4368,N_2223);
nor U8444 (N_8444,N_3878,N_4812);
nand U8445 (N_8445,N_224,N_4080);
nand U8446 (N_8446,N_2709,N_1992);
nor U8447 (N_8447,N_2793,N_184);
and U8448 (N_8448,N_1655,N_2148);
or U8449 (N_8449,N_2632,N_983);
and U8450 (N_8450,N_2055,N_4033);
nor U8451 (N_8451,N_786,N_4174);
nand U8452 (N_8452,N_4066,N_2065);
or U8453 (N_8453,N_1777,N_1932);
nand U8454 (N_8454,N_393,N_4708);
nor U8455 (N_8455,N_3328,N_4352);
nand U8456 (N_8456,N_3756,N_917);
nor U8457 (N_8457,N_2272,N_4709);
nand U8458 (N_8458,N_2015,N_2684);
nor U8459 (N_8459,N_2635,N_1129);
nand U8460 (N_8460,N_4811,N_779);
or U8461 (N_8461,N_3730,N_4938);
nor U8462 (N_8462,N_1296,N_2599);
nor U8463 (N_8463,N_4974,N_1649);
nor U8464 (N_8464,N_1631,N_531);
nor U8465 (N_8465,N_923,N_169);
and U8466 (N_8466,N_1673,N_3207);
nand U8467 (N_8467,N_847,N_4635);
and U8468 (N_8468,N_4599,N_4689);
nand U8469 (N_8469,N_1022,N_2079);
and U8470 (N_8470,N_2582,N_1869);
nand U8471 (N_8471,N_627,N_488);
and U8472 (N_8472,N_3890,N_1439);
and U8473 (N_8473,N_4722,N_3090);
or U8474 (N_8474,N_2486,N_3878);
nand U8475 (N_8475,N_2827,N_3893);
nand U8476 (N_8476,N_394,N_2888);
and U8477 (N_8477,N_3143,N_4119);
and U8478 (N_8478,N_239,N_697);
nand U8479 (N_8479,N_3520,N_3243);
nand U8480 (N_8480,N_3784,N_3722);
or U8481 (N_8481,N_1571,N_793);
or U8482 (N_8482,N_2156,N_123);
nor U8483 (N_8483,N_1610,N_193);
and U8484 (N_8484,N_3776,N_4586);
nand U8485 (N_8485,N_2839,N_4634);
or U8486 (N_8486,N_429,N_3759);
nand U8487 (N_8487,N_968,N_2287);
nor U8488 (N_8488,N_3600,N_4898);
or U8489 (N_8489,N_3246,N_2354);
nor U8490 (N_8490,N_486,N_3234);
and U8491 (N_8491,N_3560,N_3006);
and U8492 (N_8492,N_4358,N_4349);
and U8493 (N_8493,N_2293,N_860);
and U8494 (N_8494,N_54,N_745);
or U8495 (N_8495,N_304,N_4858);
and U8496 (N_8496,N_1006,N_882);
nor U8497 (N_8497,N_4017,N_585);
or U8498 (N_8498,N_3460,N_3275);
and U8499 (N_8499,N_4157,N_1383);
xor U8500 (N_8500,N_1258,N_3817);
nor U8501 (N_8501,N_946,N_211);
or U8502 (N_8502,N_4052,N_2267);
and U8503 (N_8503,N_1046,N_2858);
or U8504 (N_8504,N_2613,N_4805);
and U8505 (N_8505,N_3094,N_2395);
or U8506 (N_8506,N_333,N_3804);
nand U8507 (N_8507,N_4828,N_111);
nand U8508 (N_8508,N_3937,N_1998);
or U8509 (N_8509,N_4025,N_1892);
or U8510 (N_8510,N_382,N_799);
nand U8511 (N_8511,N_3967,N_175);
nor U8512 (N_8512,N_1791,N_2509);
and U8513 (N_8513,N_3598,N_3589);
nand U8514 (N_8514,N_4828,N_3416);
or U8515 (N_8515,N_4609,N_729);
and U8516 (N_8516,N_1226,N_1918);
nor U8517 (N_8517,N_4154,N_4601);
or U8518 (N_8518,N_2479,N_2650);
nor U8519 (N_8519,N_2830,N_1336);
nor U8520 (N_8520,N_109,N_4871);
and U8521 (N_8521,N_4857,N_3139);
and U8522 (N_8522,N_4408,N_3777);
or U8523 (N_8523,N_364,N_1368);
and U8524 (N_8524,N_2870,N_4178);
and U8525 (N_8525,N_1346,N_710);
nand U8526 (N_8526,N_8,N_2536);
or U8527 (N_8527,N_1871,N_734);
and U8528 (N_8528,N_1265,N_1942);
nor U8529 (N_8529,N_2935,N_1594);
or U8530 (N_8530,N_2622,N_2231);
and U8531 (N_8531,N_1710,N_1806);
nor U8532 (N_8532,N_1496,N_941);
nand U8533 (N_8533,N_3142,N_2);
nand U8534 (N_8534,N_2188,N_2679);
nor U8535 (N_8535,N_1487,N_1633);
or U8536 (N_8536,N_1166,N_81);
and U8537 (N_8537,N_1328,N_2592);
or U8538 (N_8538,N_1774,N_2681);
or U8539 (N_8539,N_2435,N_3053);
and U8540 (N_8540,N_1826,N_2771);
nor U8541 (N_8541,N_617,N_3446);
nand U8542 (N_8542,N_2356,N_2303);
or U8543 (N_8543,N_699,N_1743);
xor U8544 (N_8544,N_3093,N_4746);
nand U8545 (N_8545,N_2909,N_3901);
or U8546 (N_8546,N_1207,N_4953);
and U8547 (N_8547,N_2850,N_3130);
nand U8548 (N_8548,N_2143,N_794);
nand U8549 (N_8549,N_1046,N_3640);
nand U8550 (N_8550,N_3773,N_1181);
nand U8551 (N_8551,N_880,N_921);
xor U8552 (N_8552,N_2923,N_2626);
nand U8553 (N_8553,N_2542,N_1472);
or U8554 (N_8554,N_280,N_2499);
or U8555 (N_8555,N_679,N_403);
or U8556 (N_8556,N_1595,N_2034);
and U8557 (N_8557,N_3851,N_4364);
nor U8558 (N_8558,N_430,N_1036);
nor U8559 (N_8559,N_762,N_1249);
or U8560 (N_8560,N_2747,N_686);
or U8561 (N_8561,N_30,N_2962);
nor U8562 (N_8562,N_1286,N_494);
nand U8563 (N_8563,N_3273,N_3619);
or U8564 (N_8564,N_1900,N_2508);
nor U8565 (N_8565,N_3249,N_3494);
or U8566 (N_8566,N_57,N_2571);
or U8567 (N_8567,N_4617,N_3612);
nor U8568 (N_8568,N_1507,N_19);
and U8569 (N_8569,N_4530,N_542);
and U8570 (N_8570,N_1882,N_3327);
nor U8571 (N_8571,N_510,N_853);
nor U8572 (N_8572,N_259,N_1484);
and U8573 (N_8573,N_4019,N_2647);
nor U8574 (N_8574,N_2993,N_1833);
xnor U8575 (N_8575,N_3683,N_3188);
and U8576 (N_8576,N_2489,N_2028);
or U8577 (N_8577,N_2766,N_78);
nand U8578 (N_8578,N_1380,N_4771);
and U8579 (N_8579,N_2418,N_4238);
or U8580 (N_8580,N_4898,N_155);
or U8581 (N_8581,N_3857,N_76);
nor U8582 (N_8582,N_145,N_2727);
or U8583 (N_8583,N_3794,N_3450);
nand U8584 (N_8584,N_928,N_2050);
nor U8585 (N_8585,N_435,N_1611);
nor U8586 (N_8586,N_4975,N_826);
nand U8587 (N_8587,N_1866,N_568);
nor U8588 (N_8588,N_2878,N_3971);
or U8589 (N_8589,N_1686,N_702);
nor U8590 (N_8590,N_1686,N_4159);
nand U8591 (N_8591,N_3092,N_1526);
nand U8592 (N_8592,N_2541,N_4529);
nand U8593 (N_8593,N_1278,N_4704);
nand U8594 (N_8594,N_4320,N_3067);
nand U8595 (N_8595,N_1278,N_1940);
or U8596 (N_8596,N_3646,N_558);
nand U8597 (N_8597,N_1620,N_1525);
and U8598 (N_8598,N_290,N_151);
or U8599 (N_8599,N_3655,N_833);
nor U8600 (N_8600,N_4060,N_4455);
or U8601 (N_8601,N_2283,N_2531);
nor U8602 (N_8602,N_3178,N_3820);
nand U8603 (N_8603,N_3440,N_4308);
nor U8604 (N_8604,N_3167,N_846);
and U8605 (N_8605,N_4968,N_1124);
and U8606 (N_8606,N_857,N_110);
nand U8607 (N_8607,N_3960,N_3424);
and U8608 (N_8608,N_1417,N_2440);
xor U8609 (N_8609,N_3079,N_4279);
or U8610 (N_8610,N_1892,N_1526);
nor U8611 (N_8611,N_3206,N_1736);
xnor U8612 (N_8612,N_4190,N_1281);
and U8613 (N_8613,N_3431,N_2522);
and U8614 (N_8614,N_612,N_2450);
or U8615 (N_8615,N_2246,N_228);
and U8616 (N_8616,N_3723,N_2250);
and U8617 (N_8617,N_163,N_4544);
and U8618 (N_8618,N_473,N_2474);
and U8619 (N_8619,N_103,N_253);
nand U8620 (N_8620,N_90,N_2424);
and U8621 (N_8621,N_1981,N_353);
or U8622 (N_8622,N_1886,N_1599);
nand U8623 (N_8623,N_3482,N_2519);
nand U8624 (N_8624,N_3783,N_1509);
xnor U8625 (N_8625,N_1131,N_3222);
and U8626 (N_8626,N_2481,N_3331);
or U8627 (N_8627,N_3511,N_2229);
or U8628 (N_8628,N_32,N_1045);
or U8629 (N_8629,N_3497,N_2753);
nand U8630 (N_8630,N_3236,N_2215);
nor U8631 (N_8631,N_1086,N_1213);
nand U8632 (N_8632,N_4568,N_34);
and U8633 (N_8633,N_4667,N_2943);
nor U8634 (N_8634,N_4043,N_986);
nand U8635 (N_8635,N_4829,N_4015);
nor U8636 (N_8636,N_3743,N_33);
or U8637 (N_8637,N_535,N_3594);
nor U8638 (N_8638,N_19,N_4203);
xnor U8639 (N_8639,N_2859,N_3199);
nor U8640 (N_8640,N_4644,N_681);
and U8641 (N_8641,N_1345,N_3032);
and U8642 (N_8642,N_1720,N_955);
or U8643 (N_8643,N_2481,N_2535);
nor U8644 (N_8644,N_743,N_4905);
or U8645 (N_8645,N_3893,N_2789);
nor U8646 (N_8646,N_524,N_71);
and U8647 (N_8647,N_2332,N_4396);
or U8648 (N_8648,N_2731,N_3792);
and U8649 (N_8649,N_1389,N_4038);
and U8650 (N_8650,N_4434,N_1038);
or U8651 (N_8651,N_3985,N_371);
nand U8652 (N_8652,N_312,N_4952);
nor U8653 (N_8653,N_2053,N_362);
nand U8654 (N_8654,N_1219,N_3981);
nand U8655 (N_8655,N_2132,N_4693);
nor U8656 (N_8656,N_3387,N_2);
and U8657 (N_8657,N_55,N_2904);
or U8658 (N_8658,N_2634,N_368);
nand U8659 (N_8659,N_3473,N_3260);
nor U8660 (N_8660,N_747,N_1719);
or U8661 (N_8661,N_4943,N_4799);
nor U8662 (N_8662,N_1605,N_108);
or U8663 (N_8663,N_4699,N_1357);
or U8664 (N_8664,N_4153,N_1645);
and U8665 (N_8665,N_2302,N_2623);
and U8666 (N_8666,N_1869,N_2277);
or U8667 (N_8667,N_3771,N_3662);
nor U8668 (N_8668,N_1606,N_4439);
or U8669 (N_8669,N_228,N_4446);
and U8670 (N_8670,N_1143,N_3638);
or U8671 (N_8671,N_2852,N_3246);
and U8672 (N_8672,N_3999,N_229);
or U8673 (N_8673,N_985,N_4585);
or U8674 (N_8674,N_3963,N_360);
and U8675 (N_8675,N_3169,N_4550);
or U8676 (N_8676,N_3041,N_4603);
nand U8677 (N_8677,N_1323,N_1801);
or U8678 (N_8678,N_633,N_257);
nor U8679 (N_8679,N_2893,N_2748);
and U8680 (N_8680,N_3183,N_1442);
and U8681 (N_8681,N_3008,N_3090);
and U8682 (N_8682,N_4834,N_3518);
nand U8683 (N_8683,N_3245,N_700);
nand U8684 (N_8684,N_736,N_1244);
nand U8685 (N_8685,N_633,N_3534);
nand U8686 (N_8686,N_328,N_3216);
and U8687 (N_8687,N_4034,N_2040);
or U8688 (N_8688,N_2259,N_4111);
and U8689 (N_8689,N_430,N_4379);
nor U8690 (N_8690,N_4627,N_4077);
and U8691 (N_8691,N_750,N_694);
nand U8692 (N_8692,N_4545,N_1167);
or U8693 (N_8693,N_25,N_4422);
nor U8694 (N_8694,N_1334,N_442);
or U8695 (N_8695,N_1711,N_3287);
or U8696 (N_8696,N_2382,N_3377);
and U8697 (N_8697,N_1505,N_2060);
nand U8698 (N_8698,N_1379,N_916);
and U8699 (N_8699,N_3767,N_1992);
nand U8700 (N_8700,N_1516,N_4650);
nand U8701 (N_8701,N_1676,N_573);
xnor U8702 (N_8702,N_3433,N_4692);
nor U8703 (N_8703,N_881,N_672);
or U8704 (N_8704,N_2457,N_1951);
nand U8705 (N_8705,N_604,N_482);
nand U8706 (N_8706,N_2932,N_865);
nor U8707 (N_8707,N_793,N_3050);
nand U8708 (N_8708,N_1904,N_729);
or U8709 (N_8709,N_3984,N_2744);
nand U8710 (N_8710,N_1755,N_2121);
and U8711 (N_8711,N_4742,N_2722);
nor U8712 (N_8712,N_2404,N_3628);
or U8713 (N_8713,N_222,N_2392);
nand U8714 (N_8714,N_4832,N_3157);
or U8715 (N_8715,N_1865,N_4712);
or U8716 (N_8716,N_2900,N_2339);
nand U8717 (N_8717,N_4302,N_1469);
nand U8718 (N_8718,N_3609,N_2116);
or U8719 (N_8719,N_1751,N_3718);
nor U8720 (N_8720,N_4214,N_2814);
nand U8721 (N_8721,N_2738,N_3179);
or U8722 (N_8722,N_2635,N_1338);
or U8723 (N_8723,N_4049,N_4409);
and U8724 (N_8724,N_348,N_3859);
xor U8725 (N_8725,N_1337,N_3221);
nand U8726 (N_8726,N_3636,N_3233);
or U8727 (N_8727,N_4483,N_3681);
nor U8728 (N_8728,N_3832,N_2126);
or U8729 (N_8729,N_1537,N_640);
and U8730 (N_8730,N_2956,N_3794);
or U8731 (N_8731,N_3683,N_3537);
nand U8732 (N_8732,N_2848,N_2530);
and U8733 (N_8733,N_4053,N_2140);
nand U8734 (N_8734,N_798,N_4381);
nand U8735 (N_8735,N_3989,N_1438);
nor U8736 (N_8736,N_742,N_4864);
and U8737 (N_8737,N_1840,N_1895);
nand U8738 (N_8738,N_932,N_615);
and U8739 (N_8739,N_2288,N_1259);
or U8740 (N_8740,N_4414,N_4302);
or U8741 (N_8741,N_4835,N_2981);
nand U8742 (N_8742,N_1406,N_2338);
or U8743 (N_8743,N_4529,N_3510);
and U8744 (N_8744,N_4883,N_4110);
or U8745 (N_8745,N_3392,N_161);
nor U8746 (N_8746,N_2794,N_2077);
or U8747 (N_8747,N_2544,N_524);
xor U8748 (N_8748,N_1324,N_3092);
xor U8749 (N_8749,N_1855,N_3043);
nand U8750 (N_8750,N_2066,N_3083);
xnor U8751 (N_8751,N_307,N_3213);
nand U8752 (N_8752,N_3927,N_530);
or U8753 (N_8753,N_2865,N_3290);
nor U8754 (N_8754,N_2916,N_47);
nor U8755 (N_8755,N_3531,N_4284);
nor U8756 (N_8756,N_673,N_1566);
and U8757 (N_8757,N_4891,N_515);
nand U8758 (N_8758,N_3765,N_2018);
nor U8759 (N_8759,N_2053,N_4908);
and U8760 (N_8760,N_4794,N_2196);
nand U8761 (N_8761,N_373,N_4631);
nor U8762 (N_8762,N_4264,N_486);
or U8763 (N_8763,N_4377,N_202);
nand U8764 (N_8764,N_2781,N_1187);
nand U8765 (N_8765,N_3597,N_3828);
nor U8766 (N_8766,N_2528,N_4202);
nand U8767 (N_8767,N_2356,N_319);
or U8768 (N_8768,N_3675,N_4336);
nor U8769 (N_8769,N_27,N_3421);
nor U8770 (N_8770,N_3708,N_1187);
and U8771 (N_8771,N_1788,N_1602);
or U8772 (N_8772,N_3652,N_4848);
and U8773 (N_8773,N_2599,N_4802);
or U8774 (N_8774,N_293,N_1386);
nor U8775 (N_8775,N_149,N_1366);
or U8776 (N_8776,N_3051,N_3795);
and U8777 (N_8777,N_2447,N_1147);
nand U8778 (N_8778,N_2759,N_4113);
and U8779 (N_8779,N_1505,N_884);
or U8780 (N_8780,N_3037,N_3504);
nor U8781 (N_8781,N_2544,N_1327);
and U8782 (N_8782,N_912,N_2498);
nand U8783 (N_8783,N_3612,N_3415);
and U8784 (N_8784,N_1203,N_700);
nand U8785 (N_8785,N_1901,N_3643);
or U8786 (N_8786,N_4606,N_3502);
nand U8787 (N_8787,N_1635,N_3257);
nor U8788 (N_8788,N_2134,N_413);
nand U8789 (N_8789,N_887,N_2586);
nor U8790 (N_8790,N_3573,N_241);
or U8791 (N_8791,N_469,N_1463);
or U8792 (N_8792,N_3481,N_1591);
or U8793 (N_8793,N_4307,N_3821);
nor U8794 (N_8794,N_3642,N_4427);
and U8795 (N_8795,N_4436,N_3276);
nand U8796 (N_8796,N_4260,N_4337);
nand U8797 (N_8797,N_1626,N_2919);
and U8798 (N_8798,N_2079,N_2367);
nand U8799 (N_8799,N_1686,N_3035);
nand U8800 (N_8800,N_4018,N_1325);
and U8801 (N_8801,N_491,N_3045);
nand U8802 (N_8802,N_4704,N_2405);
and U8803 (N_8803,N_483,N_2562);
nand U8804 (N_8804,N_3340,N_1147);
nor U8805 (N_8805,N_4659,N_927);
or U8806 (N_8806,N_1164,N_643);
or U8807 (N_8807,N_3258,N_1713);
or U8808 (N_8808,N_3385,N_3422);
and U8809 (N_8809,N_3195,N_1890);
and U8810 (N_8810,N_3209,N_2278);
xnor U8811 (N_8811,N_1460,N_1672);
and U8812 (N_8812,N_3065,N_3797);
and U8813 (N_8813,N_4314,N_4684);
or U8814 (N_8814,N_1793,N_174);
nand U8815 (N_8815,N_375,N_4477);
nand U8816 (N_8816,N_2636,N_616);
nand U8817 (N_8817,N_2808,N_1839);
and U8818 (N_8818,N_3350,N_3235);
xnor U8819 (N_8819,N_2756,N_4263);
nor U8820 (N_8820,N_4085,N_3061);
or U8821 (N_8821,N_2330,N_4515);
or U8822 (N_8822,N_4259,N_636);
and U8823 (N_8823,N_2419,N_1098);
nor U8824 (N_8824,N_4895,N_258);
and U8825 (N_8825,N_4313,N_2066);
xnor U8826 (N_8826,N_2808,N_4483);
nor U8827 (N_8827,N_3303,N_3556);
or U8828 (N_8828,N_3867,N_3322);
or U8829 (N_8829,N_427,N_2873);
and U8830 (N_8830,N_1837,N_2262);
nand U8831 (N_8831,N_2710,N_2166);
nor U8832 (N_8832,N_1120,N_4564);
nand U8833 (N_8833,N_3115,N_3678);
or U8834 (N_8834,N_2495,N_2806);
or U8835 (N_8835,N_848,N_3373);
nand U8836 (N_8836,N_4852,N_900);
and U8837 (N_8837,N_4942,N_2749);
or U8838 (N_8838,N_3450,N_3349);
or U8839 (N_8839,N_2658,N_2059);
nor U8840 (N_8840,N_2816,N_2969);
nor U8841 (N_8841,N_2888,N_1050);
or U8842 (N_8842,N_4654,N_4593);
and U8843 (N_8843,N_1467,N_4250);
and U8844 (N_8844,N_1795,N_861);
or U8845 (N_8845,N_3339,N_2686);
and U8846 (N_8846,N_4054,N_2104);
nand U8847 (N_8847,N_1085,N_1868);
or U8848 (N_8848,N_3771,N_1971);
nand U8849 (N_8849,N_3724,N_3818);
nor U8850 (N_8850,N_960,N_4756);
and U8851 (N_8851,N_1159,N_744);
or U8852 (N_8852,N_1810,N_4097);
nand U8853 (N_8853,N_4429,N_1040);
nor U8854 (N_8854,N_1700,N_2030);
nand U8855 (N_8855,N_3964,N_684);
and U8856 (N_8856,N_690,N_1697);
nand U8857 (N_8857,N_117,N_650);
and U8858 (N_8858,N_862,N_1585);
or U8859 (N_8859,N_4672,N_164);
and U8860 (N_8860,N_114,N_628);
xnor U8861 (N_8861,N_1269,N_3661);
or U8862 (N_8862,N_2936,N_4769);
and U8863 (N_8863,N_27,N_742);
nand U8864 (N_8864,N_932,N_1109);
nand U8865 (N_8865,N_2341,N_4305);
nand U8866 (N_8866,N_1217,N_1043);
or U8867 (N_8867,N_4895,N_1857);
nand U8868 (N_8868,N_2220,N_2840);
and U8869 (N_8869,N_3344,N_731);
and U8870 (N_8870,N_2087,N_335);
nand U8871 (N_8871,N_1115,N_2134);
nand U8872 (N_8872,N_181,N_2877);
nor U8873 (N_8873,N_278,N_2749);
nand U8874 (N_8874,N_3717,N_949);
nand U8875 (N_8875,N_208,N_2790);
and U8876 (N_8876,N_2160,N_190);
nand U8877 (N_8877,N_3985,N_3683);
nand U8878 (N_8878,N_1223,N_4762);
or U8879 (N_8879,N_2921,N_1897);
nand U8880 (N_8880,N_4038,N_1985);
or U8881 (N_8881,N_3704,N_115);
nor U8882 (N_8882,N_772,N_2388);
or U8883 (N_8883,N_4726,N_2954);
or U8884 (N_8884,N_2965,N_1993);
and U8885 (N_8885,N_3714,N_3431);
and U8886 (N_8886,N_862,N_3208);
nor U8887 (N_8887,N_3147,N_3985);
and U8888 (N_8888,N_3439,N_4085);
nor U8889 (N_8889,N_960,N_832);
and U8890 (N_8890,N_2293,N_1430);
nor U8891 (N_8891,N_4651,N_3179);
nand U8892 (N_8892,N_2218,N_903);
and U8893 (N_8893,N_2753,N_4867);
nand U8894 (N_8894,N_1053,N_1748);
and U8895 (N_8895,N_3053,N_164);
or U8896 (N_8896,N_1177,N_1287);
and U8897 (N_8897,N_2155,N_3711);
nand U8898 (N_8898,N_2358,N_1045);
nand U8899 (N_8899,N_2393,N_2151);
and U8900 (N_8900,N_2126,N_4808);
and U8901 (N_8901,N_3018,N_1435);
nand U8902 (N_8902,N_1811,N_1237);
nor U8903 (N_8903,N_325,N_3870);
and U8904 (N_8904,N_3769,N_148);
nor U8905 (N_8905,N_3697,N_1635);
and U8906 (N_8906,N_4573,N_2998);
and U8907 (N_8907,N_799,N_2632);
or U8908 (N_8908,N_3734,N_682);
or U8909 (N_8909,N_2812,N_500);
nand U8910 (N_8910,N_1818,N_4882);
or U8911 (N_8911,N_2383,N_4634);
xnor U8912 (N_8912,N_417,N_4085);
nand U8913 (N_8913,N_4561,N_2980);
and U8914 (N_8914,N_823,N_4386);
and U8915 (N_8915,N_3073,N_110);
or U8916 (N_8916,N_2935,N_1051);
nor U8917 (N_8917,N_4198,N_610);
nand U8918 (N_8918,N_3652,N_982);
nand U8919 (N_8919,N_3781,N_1137);
and U8920 (N_8920,N_2033,N_3438);
and U8921 (N_8921,N_2634,N_278);
and U8922 (N_8922,N_2884,N_2983);
or U8923 (N_8923,N_578,N_1834);
nor U8924 (N_8924,N_3954,N_1682);
nor U8925 (N_8925,N_1663,N_2173);
and U8926 (N_8926,N_138,N_4427);
nor U8927 (N_8927,N_1169,N_2113);
nor U8928 (N_8928,N_185,N_1398);
or U8929 (N_8929,N_4680,N_4273);
nor U8930 (N_8930,N_645,N_4831);
nor U8931 (N_8931,N_1463,N_4359);
and U8932 (N_8932,N_785,N_2119);
nand U8933 (N_8933,N_4467,N_319);
or U8934 (N_8934,N_4336,N_2118);
and U8935 (N_8935,N_744,N_2488);
and U8936 (N_8936,N_1043,N_1193);
nor U8937 (N_8937,N_4567,N_3106);
or U8938 (N_8938,N_2806,N_4622);
nand U8939 (N_8939,N_3962,N_1853);
nor U8940 (N_8940,N_699,N_1653);
and U8941 (N_8941,N_2152,N_4472);
or U8942 (N_8942,N_2072,N_4997);
nand U8943 (N_8943,N_3414,N_4440);
nand U8944 (N_8944,N_3210,N_2991);
and U8945 (N_8945,N_943,N_3934);
and U8946 (N_8946,N_3616,N_827);
nand U8947 (N_8947,N_1866,N_1483);
nand U8948 (N_8948,N_3264,N_4690);
xnor U8949 (N_8949,N_2620,N_3137);
and U8950 (N_8950,N_255,N_1343);
nand U8951 (N_8951,N_2719,N_2704);
nor U8952 (N_8952,N_4252,N_4440);
nor U8953 (N_8953,N_1794,N_3614);
nand U8954 (N_8954,N_3411,N_2868);
nand U8955 (N_8955,N_591,N_3305);
nand U8956 (N_8956,N_3279,N_3868);
nand U8957 (N_8957,N_815,N_1929);
and U8958 (N_8958,N_3977,N_4965);
and U8959 (N_8959,N_2742,N_4346);
nor U8960 (N_8960,N_3845,N_938);
or U8961 (N_8961,N_3647,N_4486);
nor U8962 (N_8962,N_1326,N_445);
nor U8963 (N_8963,N_2305,N_2703);
or U8964 (N_8964,N_1136,N_4645);
or U8965 (N_8965,N_1017,N_3480);
nand U8966 (N_8966,N_4022,N_4263);
nand U8967 (N_8967,N_478,N_4614);
or U8968 (N_8968,N_4311,N_1289);
and U8969 (N_8969,N_4792,N_3199);
and U8970 (N_8970,N_2058,N_4174);
or U8971 (N_8971,N_4286,N_4721);
or U8972 (N_8972,N_4107,N_2896);
and U8973 (N_8973,N_3987,N_1988);
nand U8974 (N_8974,N_1717,N_3396);
or U8975 (N_8975,N_3,N_2739);
or U8976 (N_8976,N_537,N_5);
and U8977 (N_8977,N_3293,N_965);
nor U8978 (N_8978,N_1271,N_2983);
and U8979 (N_8979,N_2483,N_447);
and U8980 (N_8980,N_2794,N_4436);
nor U8981 (N_8981,N_1548,N_2368);
or U8982 (N_8982,N_2227,N_1547);
nand U8983 (N_8983,N_2255,N_1731);
and U8984 (N_8984,N_1133,N_3630);
nor U8985 (N_8985,N_796,N_4609);
and U8986 (N_8986,N_1265,N_4285);
nor U8987 (N_8987,N_3765,N_3528);
and U8988 (N_8988,N_392,N_3033);
nor U8989 (N_8989,N_1857,N_778);
xnor U8990 (N_8990,N_525,N_1825);
or U8991 (N_8991,N_875,N_305);
nor U8992 (N_8992,N_579,N_3868);
and U8993 (N_8993,N_3601,N_2319);
nor U8994 (N_8994,N_2132,N_2039);
nor U8995 (N_8995,N_4427,N_467);
nand U8996 (N_8996,N_3009,N_2311);
nor U8997 (N_8997,N_3968,N_513);
and U8998 (N_8998,N_4721,N_3951);
or U8999 (N_8999,N_938,N_3558);
and U9000 (N_9000,N_3386,N_2098);
and U9001 (N_9001,N_1384,N_2551);
nand U9002 (N_9002,N_2289,N_4417);
or U9003 (N_9003,N_2480,N_4674);
nand U9004 (N_9004,N_1261,N_4498);
or U9005 (N_9005,N_3288,N_626);
or U9006 (N_9006,N_3247,N_2958);
nand U9007 (N_9007,N_4351,N_948);
nor U9008 (N_9008,N_1970,N_1137);
nor U9009 (N_9009,N_3228,N_2080);
or U9010 (N_9010,N_2081,N_3690);
nor U9011 (N_9011,N_1146,N_3372);
or U9012 (N_9012,N_1778,N_1706);
nor U9013 (N_9013,N_1062,N_272);
nor U9014 (N_9014,N_4133,N_4180);
and U9015 (N_9015,N_2400,N_1370);
nand U9016 (N_9016,N_994,N_824);
nor U9017 (N_9017,N_1439,N_3355);
and U9018 (N_9018,N_3999,N_2473);
and U9019 (N_9019,N_1336,N_4673);
nand U9020 (N_9020,N_4842,N_424);
nor U9021 (N_9021,N_2996,N_4838);
nand U9022 (N_9022,N_3608,N_3308);
and U9023 (N_9023,N_725,N_122);
nand U9024 (N_9024,N_4898,N_1900);
nor U9025 (N_9025,N_230,N_2790);
or U9026 (N_9026,N_2655,N_1191);
nand U9027 (N_9027,N_3559,N_4934);
or U9028 (N_9028,N_3599,N_4856);
and U9029 (N_9029,N_1124,N_478);
nand U9030 (N_9030,N_1589,N_4036);
or U9031 (N_9031,N_3158,N_231);
and U9032 (N_9032,N_1202,N_3433);
and U9033 (N_9033,N_686,N_2603);
or U9034 (N_9034,N_3321,N_4735);
and U9035 (N_9035,N_2796,N_4318);
and U9036 (N_9036,N_222,N_3619);
nor U9037 (N_9037,N_1067,N_2370);
nand U9038 (N_9038,N_226,N_3134);
xnor U9039 (N_9039,N_342,N_1099);
nand U9040 (N_9040,N_2006,N_3015);
nand U9041 (N_9041,N_3385,N_1928);
nand U9042 (N_9042,N_3356,N_3714);
nand U9043 (N_9043,N_4503,N_399);
nand U9044 (N_9044,N_4928,N_1162);
or U9045 (N_9045,N_2331,N_1399);
nand U9046 (N_9046,N_3173,N_2692);
and U9047 (N_9047,N_2169,N_80);
nor U9048 (N_9048,N_1504,N_489);
nand U9049 (N_9049,N_2506,N_87);
or U9050 (N_9050,N_4903,N_1346);
nand U9051 (N_9051,N_742,N_2341);
and U9052 (N_9052,N_2423,N_760);
and U9053 (N_9053,N_2696,N_4044);
and U9054 (N_9054,N_310,N_2260);
or U9055 (N_9055,N_4281,N_3807);
or U9056 (N_9056,N_3074,N_2689);
and U9057 (N_9057,N_1255,N_1896);
or U9058 (N_9058,N_3022,N_2358);
nor U9059 (N_9059,N_4732,N_283);
nor U9060 (N_9060,N_4577,N_1999);
nor U9061 (N_9061,N_4289,N_1426);
nand U9062 (N_9062,N_872,N_3519);
nand U9063 (N_9063,N_1105,N_4161);
or U9064 (N_9064,N_1445,N_231);
nor U9065 (N_9065,N_2475,N_4226);
or U9066 (N_9066,N_3935,N_1676);
nor U9067 (N_9067,N_536,N_1917);
nand U9068 (N_9068,N_4604,N_2752);
or U9069 (N_9069,N_352,N_651);
nor U9070 (N_9070,N_987,N_4804);
and U9071 (N_9071,N_896,N_3733);
or U9072 (N_9072,N_21,N_4166);
or U9073 (N_9073,N_4754,N_3736);
or U9074 (N_9074,N_3729,N_3022);
nor U9075 (N_9075,N_4165,N_1706);
nor U9076 (N_9076,N_2724,N_708);
nor U9077 (N_9077,N_3905,N_533);
nor U9078 (N_9078,N_626,N_877);
nand U9079 (N_9079,N_4929,N_5);
and U9080 (N_9080,N_2225,N_520);
nand U9081 (N_9081,N_3804,N_3016);
nand U9082 (N_9082,N_1488,N_4296);
or U9083 (N_9083,N_4223,N_1492);
nor U9084 (N_9084,N_1885,N_3018);
or U9085 (N_9085,N_175,N_4983);
or U9086 (N_9086,N_4131,N_3650);
xor U9087 (N_9087,N_2403,N_2225);
or U9088 (N_9088,N_693,N_3329);
nand U9089 (N_9089,N_3796,N_268);
and U9090 (N_9090,N_3517,N_2140);
nand U9091 (N_9091,N_1245,N_4541);
nor U9092 (N_9092,N_1031,N_1341);
and U9093 (N_9093,N_4353,N_2737);
or U9094 (N_9094,N_3291,N_482);
and U9095 (N_9095,N_1804,N_2713);
and U9096 (N_9096,N_955,N_974);
nor U9097 (N_9097,N_3820,N_1988);
or U9098 (N_9098,N_4086,N_3383);
nand U9099 (N_9099,N_4330,N_1659);
nand U9100 (N_9100,N_3873,N_3200);
nand U9101 (N_9101,N_3208,N_112);
or U9102 (N_9102,N_2357,N_1257);
nand U9103 (N_9103,N_3733,N_2968);
or U9104 (N_9104,N_4962,N_92);
or U9105 (N_9105,N_2118,N_125);
nand U9106 (N_9106,N_1469,N_3463);
nor U9107 (N_9107,N_3285,N_2713);
nand U9108 (N_9108,N_1833,N_1136);
nor U9109 (N_9109,N_4004,N_4212);
nor U9110 (N_9110,N_366,N_4523);
nand U9111 (N_9111,N_3886,N_1853);
or U9112 (N_9112,N_4307,N_423);
and U9113 (N_9113,N_53,N_1018);
and U9114 (N_9114,N_3138,N_3845);
xor U9115 (N_9115,N_603,N_1567);
or U9116 (N_9116,N_4361,N_3009);
or U9117 (N_9117,N_1585,N_2652);
nand U9118 (N_9118,N_3019,N_4937);
and U9119 (N_9119,N_2732,N_1192);
nor U9120 (N_9120,N_4707,N_3817);
and U9121 (N_9121,N_882,N_3938);
nand U9122 (N_9122,N_2742,N_4283);
or U9123 (N_9123,N_4760,N_1092);
xnor U9124 (N_9124,N_1635,N_1103);
nand U9125 (N_9125,N_3630,N_3474);
or U9126 (N_9126,N_2524,N_622);
nor U9127 (N_9127,N_1300,N_2425);
or U9128 (N_9128,N_1898,N_1264);
nor U9129 (N_9129,N_415,N_495);
nor U9130 (N_9130,N_296,N_2809);
or U9131 (N_9131,N_758,N_756);
nor U9132 (N_9132,N_1391,N_2829);
nand U9133 (N_9133,N_4035,N_4832);
nor U9134 (N_9134,N_4756,N_614);
or U9135 (N_9135,N_3570,N_1936);
and U9136 (N_9136,N_3251,N_1047);
and U9137 (N_9137,N_956,N_146);
nand U9138 (N_9138,N_2895,N_1698);
nand U9139 (N_9139,N_4824,N_1689);
or U9140 (N_9140,N_3795,N_3505);
nand U9141 (N_9141,N_916,N_2518);
or U9142 (N_9142,N_777,N_3044);
and U9143 (N_9143,N_4698,N_4486);
nand U9144 (N_9144,N_4616,N_4543);
nor U9145 (N_9145,N_2866,N_4601);
and U9146 (N_9146,N_2056,N_593);
or U9147 (N_9147,N_3640,N_873);
nor U9148 (N_9148,N_3971,N_352);
or U9149 (N_9149,N_1745,N_4561);
and U9150 (N_9150,N_499,N_4192);
nor U9151 (N_9151,N_1739,N_4163);
nand U9152 (N_9152,N_3491,N_3713);
nor U9153 (N_9153,N_1309,N_2581);
or U9154 (N_9154,N_3567,N_1500);
nand U9155 (N_9155,N_4789,N_4930);
nor U9156 (N_9156,N_3688,N_1282);
nand U9157 (N_9157,N_3776,N_1422);
or U9158 (N_9158,N_493,N_876);
or U9159 (N_9159,N_652,N_2814);
nand U9160 (N_9160,N_1337,N_3079);
or U9161 (N_9161,N_4206,N_991);
nand U9162 (N_9162,N_4381,N_1468);
or U9163 (N_9163,N_2739,N_1285);
nor U9164 (N_9164,N_463,N_2597);
nor U9165 (N_9165,N_4708,N_2002);
nor U9166 (N_9166,N_883,N_1245);
nor U9167 (N_9167,N_2928,N_4618);
nand U9168 (N_9168,N_3923,N_175);
and U9169 (N_9169,N_2893,N_1815);
and U9170 (N_9170,N_3908,N_3692);
nand U9171 (N_9171,N_431,N_1933);
nor U9172 (N_9172,N_3985,N_673);
and U9173 (N_9173,N_4758,N_2334);
nor U9174 (N_9174,N_3174,N_4972);
and U9175 (N_9175,N_3894,N_4056);
or U9176 (N_9176,N_2909,N_247);
nand U9177 (N_9177,N_4722,N_3841);
or U9178 (N_9178,N_3013,N_4454);
or U9179 (N_9179,N_4703,N_537);
and U9180 (N_9180,N_4408,N_443);
xnor U9181 (N_9181,N_404,N_3755);
or U9182 (N_9182,N_2194,N_4911);
nand U9183 (N_9183,N_3807,N_600);
xor U9184 (N_9184,N_2389,N_2124);
or U9185 (N_9185,N_4970,N_4323);
or U9186 (N_9186,N_3092,N_4968);
nor U9187 (N_9187,N_3420,N_1007);
and U9188 (N_9188,N_1562,N_4055);
and U9189 (N_9189,N_4062,N_1799);
nor U9190 (N_9190,N_530,N_373);
nor U9191 (N_9191,N_2176,N_140);
nor U9192 (N_9192,N_3909,N_4197);
nand U9193 (N_9193,N_3803,N_3138);
xor U9194 (N_9194,N_2497,N_4491);
nor U9195 (N_9195,N_3818,N_4332);
nand U9196 (N_9196,N_3772,N_2005);
or U9197 (N_9197,N_507,N_4491);
nor U9198 (N_9198,N_2739,N_4736);
and U9199 (N_9199,N_481,N_4650);
and U9200 (N_9200,N_4489,N_2810);
or U9201 (N_9201,N_3259,N_2313);
nor U9202 (N_9202,N_2692,N_3680);
nand U9203 (N_9203,N_2162,N_4545);
nor U9204 (N_9204,N_4780,N_481);
or U9205 (N_9205,N_2176,N_234);
or U9206 (N_9206,N_802,N_1935);
nor U9207 (N_9207,N_1787,N_1212);
or U9208 (N_9208,N_1328,N_4691);
nor U9209 (N_9209,N_182,N_1750);
or U9210 (N_9210,N_3161,N_3384);
and U9211 (N_9211,N_2546,N_3944);
and U9212 (N_9212,N_1085,N_4018);
nand U9213 (N_9213,N_4151,N_1215);
and U9214 (N_9214,N_4096,N_2770);
or U9215 (N_9215,N_618,N_1999);
nor U9216 (N_9216,N_3748,N_1857);
and U9217 (N_9217,N_823,N_2068);
or U9218 (N_9218,N_857,N_1389);
nor U9219 (N_9219,N_369,N_3723);
nand U9220 (N_9220,N_3230,N_4502);
and U9221 (N_9221,N_1666,N_4804);
nor U9222 (N_9222,N_2930,N_2736);
and U9223 (N_9223,N_2792,N_965);
or U9224 (N_9224,N_744,N_3338);
nor U9225 (N_9225,N_4551,N_2896);
and U9226 (N_9226,N_1851,N_1506);
nor U9227 (N_9227,N_3882,N_1632);
or U9228 (N_9228,N_2530,N_625);
nor U9229 (N_9229,N_2236,N_2449);
nand U9230 (N_9230,N_1070,N_390);
or U9231 (N_9231,N_3236,N_3559);
nand U9232 (N_9232,N_4660,N_4442);
nand U9233 (N_9233,N_4685,N_187);
or U9234 (N_9234,N_849,N_787);
and U9235 (N_9235,N_2168,N_1932);
and U9236 (N_9236,N_4897,N_4309);
or U9237 (N_9237,N_342,N_1096);
nor U9238 (N_9238,N_4885,N_253);
or U9239 (N_9239,N_3743,N_2164);
and U9240 (N_9240,N_427,N_1122);
nor U9241 (N_9241,N_510,N_4438);
or U9242 (N_9242,N_2622,N_2689);
nand U9243 (N_9243,N_3801,N_12);
or U9244 (N_9244,N_4292,N_546);
nor U9245 (N_9245,N_670,N_263);
nand U9246 (N_9246,N_1152,N_3216);
nand U9247 (N_9247,N_609,N_3836);
xnor U9248 (N_9248,N_3781,N_2280);
and U9249 (N_9249,N_4700,N_2425);
nand U9250 (N_9250,N_4775,N_506);
nor U9251 (N_9251,N_631,N_3856);
or U9252 (N_9252,N_4556,N_1626);
nand U9253 (N_9253,N_1606,N_2523);
and U9254 (N_9254,N_454,N_3159);
nand U9255 (N_9255,N_2612,N_2821);
nand U9256 (N_9256,N_1814,N_902);
or U9257 (N_9257,N_3709,N_4561);
nand U9258 (N_9258,N_4030,N_1709);
nor U9259 (N_9259,N_3543,N_881);
nor U9260 (N_9260,N_4063,N_2237);
or U9261 (N_9261,N_3413,N_776);
xnor U9262 (N_9262,N_160,N_4867);
and U9263 (N_9263,N_1405,N_4565);
nor U9264 (N_9264,N_3134,N_4432);
or U9265 (N_9265,N_2673,N_2727);
nand U9266 (N_9266,N_4894,N_4155);
or U9267 (N_9267,N_1424,N_3637);
and U9268 (N_9268,N_2849,N_3486);
nor U9269 (N_9269,N_2003,N_4187);
or U9270 (N_9270,N_113,N_4923);
and U9271 (N_9271,N_2745,N_1575);
and U9272 (N_9272,N_1059,N_3672);
nand U9273 (N_9273,N_4209,N_2596);
and U9274 (N_9274,N_1726,N_2266);
or U9275 (N_9275,N_462,N_312);
or U9276 (N_9276,N_4336,N_3980);
xnor U9277 (N_9277,N_4034,N_722);
and U9278 (N_9278,N_3136,N_2655);
or U9279 (N_9279,N_3781,N_2327);
nor U9280 (N_9280,N_1035,N_3242);
nor U9281 (N_9281,N_361,N_2089);
nor U9282 (N_9282,N_29,N_1308);
nor U9283 (N_9283,N_2956,N_1192);
nor U9284 (N_9284,N_2773,N_2142);
or U9285 (N_9285,N_4616,N_1588);
nand U9286 (N_9286,N_3171,N_2113);
nor U9287 (N_9287,N_2886,N_2685);
nand U9288 (N_9288,N_3980,N_1762);
nor U9289 (N_9289,N_95,N_4179);
nor U9290 (N_9290,N_3327,N_841);
nor U9291 (N_9291,N_1827,N_2945);
and U9292 (N_9292,N_742,N_3667);
nand U9293 (N_9293,N_2634,N_871);
or U9294 (N_9294,N_1751,N_858);
nand U9295 (N_9295,N_317,N_2636);
and U9296 (N_9296,N_805,N_946);
or U9297 (N_9297,N_712,N_1878);
or U9298 (N_9298,N_1494,N_4226);
nor U9299 (N_9299,N_1101,N_4679);
or U9300 (N_9300,N_1980,N_323);
nand U9301 (N_9301,N_1230,N_4054);
nor U9302 (N_9302,N_3458,N_1628);
and U9303 (N_9303,N_3611,N_2419);
nor U9304 (N_9304,N_3335,N_3403);
nand U9305 (N_9305,N_97,N_662);
xnor U9306 (N_9306,N_1076,N_3866);
nand U9307 (N_9307,N_77,N_3354);
or U9308 (N_9308,N_656,N_1650);
nand U9309 (N_9309,N_3734,N_4143);
nor U9310 (N_9310,N_4409,N_1298);
and U9311 (N_9311,N_814,N_294);
nand U9312 (N_9312,N_2426,N_3761);
or U9313 (N_9313,N_1768,N_1837);
or U9314 (N_9314,N_3629,N_1955);
nand U9315 (N_9315,N_466,N_2997);
nand U9316 (N_9316,N_3471,N_3249);
or U9317 (N_9317,N_4644,N_4099);
nor U9318 (N_9318,N_283,N_1297);
and U9319 (N_9319,N_499,N_3972);
and U9320 (N_9320,N_3880,N_3929);
nand U9321 (N_9321,N_4193,N_1739);
nand U9322 (N_9322,N_1521,N_508);
nand U9323 (N_9323,N_1068,N_1822);
nand U9324 (N_9324,N_4248,N_3780);
or U9325 (N_9325,N_2578,N_4195);
or U9326 (N_9326,N_3019,N_689);
nand U9327 (N_9327,N_4341,N_4243);
and U9328 (N_9328,N_3972,N_1782);
nor U9329 (N_9329,N_3010,N_343);
or U9330 (N_9330,N_3330,N_3720);
and U9331 (N_9331,N_2542,N_2707);
and U9332 (N_9332,N_281,N_2336);
and U9333 (N_9333,N_2255,N_3435);
and U9334 (N_9334,N_3903,N_1767);
or U9335 (N_9335,N_1487,N_2397);
xnor U9336 (N_9336,N_1334,N_4874);
and U9337 (N_9337,N_788,N_370);
nand U9338 (N_9338,N_1296,N_3007);
nor U9339 (N_9339,N_864,N_4428);
and U9340 (N_9340,N_3831,N_2867);
nand U9341 (N_9341,N_4037,N_2498);
nand U9342 (N_9342,N_3994,N_2582);
or U9343 (N_9343,N_1991,N_898);
or U9344 (N_9344,N_3309,N_4855);
nor U9345 (N_9345,N_4318,N_1076);
nand U9346 (N_9346,N_6,N_4757);
nand U9347 (N_9347,N_1232,N_1437);
nor U9348 (N_9348,N_1318,N_4611);
and U9349 (N_9349,N_3366,N_1739);
or U9350 (N_9350,N_4739,N_2699);
and U9351 (N_9351,N_2366,N_4421);
and U9352 (N_9352,N_3179,N_1789);
and U9353 (N_9353,N_4270,N_3977);
or U9354 (N_9354,N_2165,N_3442);
xor U9355 (N_9355,N_3852,N_2900);
or U9356 (N_9356,N_3544,N_283);
or U9357 (N_9357,N_142,N_950);
nor U9358 (N_9358,N_3412,N_3320);
nand U9359 (N_9359,N_2899,N_2354);
or U9360 (N_9360,N_499,N_262);
or U9361 (N_9361,N_581,N_4157);
or U9362 (N_9362,N_3525,N_1366);
nor U9363 (N_9363,N_1923,N_4352);
nand U9364 (N_9364,N_696,N_3992);
or U9365 (N_9365,N_223,N_707);
xor U9366 (N_9366,N_41,N_2915);
or U9367 (N_9367,N_1349,N_2290);
nand U9368 (N_9368,N_1786,N_4112);
nor U9369 (N_9369,N_1953,N_4885);
xor U9370 (N_9370,N_2429,N_1178);
and U9371 (N_9371,N_3149,N_4865);
or U9372 (N_9372,N_3098,N_3617);
nand U9373 (N_9373,N_4965,N_4661);
nand U9374 (N_9374,N_2907,N_1958);
and U9375 (N_9375,N_2799,N_119);
xnor U9376 (N_9376,N_1742,N_3344);
nor U9377 (N_9377,N_4052,N_4629);
nor U9378 (N_9378,N_4249,N_440);
xor U9379 (N_9379,N_3763,N_2434);
or U9380 (N_9380,N_4591,N_290);
nand U9381 (N_9381,N_2779,N_1904);
or U9382 (N_9382,N_1148,N_3579);
nor U9383 (N_9383,N_2823,N_598);
nor U9384 (N_9384,N_4225,N_3913);
nor U9385 (N_9385,N_1906,N_4344);
or U9386 (N_9386,N_2141,N_599);
nand U9387 (N_9387,N_3601,N_756);
and U9388 (N_9388,N_208,N_2347);
and U9389 (N_9389,N_4002,N_3157);
or U9390 (N_9390,N_2406,N_101);
nor U9391 (N_9391,N_3725,N_4845);
and U9392 (N_9392,N_911,N_4280);
or U9393 (N_9393,N_4207,N_3636);
or U9394 (N_9394,N_1486,N_1436);
nor U9395 (N_9395,N_2799,N_2984);
and U9396 (N_9396,N_600,N_2323);
nand U9397 (N_9397,N_3181,N_2969);
nor U9398 (N_9398,N_895,N_1337);
nand U9399 (N_9399,N_1668,N_2025);
and U9400 (N_9400,N_4217,N_2520);
nand U9401 (N_9401,N_4688,N_4418);
nor U9402 (N_9402,N_4640,N_10);
and U9403 (N_9403,N_1734,N_3190);
nand U9404 (N_9404,N_2465,N_777);
and U9405 (N_9405,N_2348,N_477);
nor U9406 (N_9406,N_2928,N_4340);
and U9407 (N_9407,N_1997,N_836);
and U9408 (N_9408,N_21,N_3488);
nand U9409 (N_9409,N_3026,N_3491);
nor U9410 (N_9410,N_2012,N_4946);
nor U9411 (N_9411,N_93,N_2688);
nor U9412 (N_9412,N_4517,N_4167);
nor U9413 (N_9413,N_1820,N_4009);
or U9414 (N_9414,N_4909,N_421);
or U9415 (N_9415,N_2377,N_3461);
or U9416 (N_9416,N_152,N_4109);
and U9417 (N_9417,N_356,N_4476);
or U9418 (N_9418,N_2632,N_2817);
and U9419 (N_9419,N_3833,N_2502);
xnor U9420 (N_9420,N_2772,N_2041);
nand U9421 (N_9421,N_1493,N_3661);
nor U9422 (N_9422,N_2350,N_2484);
or U9423 (N_9423,N_3495,N_1350);
or U9424 (N_9424,N_881,N_1983);
and U9425 (N_9425,N_2612,N_1723);
or U9426 (N_9426,N_4046,N_1379);
nand U9427 (N_9427,N_260,N_119);
nor U9428 (N_9428,N_2853,N_3760);
and U9429 (N_9429,N_2823,N_816);
nor U9430 (N_9430,N_1522,N_3519);
nor U9431 (N_9431,N_3989,N_2202);
nand U9432 (N_9432,N_1289,N_1500);
nand U9433 (N_9433,N_4713,N_3671);
nand U9434 (N_9434,N_4481,N_3075);
or U9435 (N_9435,N_2122,N_4342);
and U9436 (N_9436,N_4802,N_4328);
nor U9437 (N_9437,N_2990,N_780);
or U9438 (N_9438,N_4067,N_3179);
nor U9439 (N_9439,N_936,N_3846);
and U9440 (N_9440,N_1549,N_939);
nor U9441 (N_9441,N_1724,N_1836);
nor U9442 (N_9442,N_859,N_182);
nand U9443 (N_9443,N_4812,N_2645);
nor U9444 (N_9444,N_4336,N_337);
or U9445 (N_9445,N_1940,N_1203);
and U9446 (N_9446,N_3962,N_2281);
and U9447 (N_9447,N_4936,N_3750);
nand U9448 (N_9448,N_3394,N_4791);
and U9449 (N_9449,N_2281,N_4728);
nand U9450 (N_9450,N_4135,N_4064);
and U9451 (N_9451,N_3652,N_1681);
nor U9452 (N_9452,N_765,N_3589);
nor U9453 (N_9453,N_2983,N_2911);
or U9454 (N_9454,N_1085,N_2127);
and U9455 (N_9455,N_3116,N_971);
or U9456 (N_9456,N_843,N_3308);
and U9457 (N_9457,N_1684,N_493);
nand U9458 (N_9458,N_127,N_1663);
and U9459 (N_9459,N_1021,N_1995);
nand U9460 (N_9460,N_1947,N_979);
or U9461 (N_9461,N_736,N_4087);
and U9462 (N_9462,N_3913,N_3836);
nor U9463 (N_9463,N_2041,N_1301);
or U9464 (N_9464,N_4673,N_3733);
nand U9465 (N_9465,N_1756,N_2626);
nor U9466 (N_9466,N_3752,N_4936);
nand U9467 (N_9467,N_893,N_974);
nand U9468 (N_9468,N_1020,N_2196);
and U9469 (N_9469,N_2354,N_1718);
nand U9470 (N_9470,N_3144,N_1737);
nand U9471 (N_9471,N_2207,N_1995);
nand U9472 (N_9472,N_3245,N_4711);
nor U9473 (N_9473,N_1424,N_2118);
and U9474 (N_9474,N_4409,N_1494);
or U9475 (N_9475,N_1729,N_4516);
nor U9476 (N_9476,N_2776,N_1703);
nand U9477 (N_9477,N_1954,N_3775);
or U9478 (N_9478,N_4105,N_1227);
and U9479 (N_9479,N_3855,N_2892);
or U9480 (N_9480,N_2226,N_433);
nor U9481 (N_9481,N_689,N_599);
or U9482 (N_9482,N_362,N_2829);
or U9483 (N_9483,N_3632,N_1744);
and U9484 (N_9484,N_2459,N_2058);
and U9485 (N_9485,N_4655,N_2944);
nor U9486 (N_9486,N_3795,N_3393);
and U9487 (N_9487,N_2543,N_4032);
xnor U9488 (N_9488,N_3934,N_1937);
or U9489 (N_9489,N_4879,N_4187);
or U9490 (N_9490,N_1731,N_3892);
nor U9491 (N_9491,N_4988,N_4829);
nand U9492 (N_9492,N_805,N_3097);
xnor U9493 (N_9493,N_3706,N_3728);
nand U9494 (N_9494,N_1825,N_1643);
nor U9495 (N_9495,N_3938,N_2812);
and U9496 (N_9496,N_2082,N_3752);
xor U9497 (N_9497,N_1930,N_740);
nor U9498 (N_9498,N_3181,N_4606);
and U9499 (N_9499,N_4346,N_840);
xor U9500 (N_9500,N_2217,N_2773);
nand U9501 (N_9501,N_4914,N_247);
nand U9502 (N_9502,N_2186,N_654);
nor U9503 (N_9503,N_3250,N_1539);
or U9504 (N_9504,N_492,N_3216);
nor U9505 (N_9505,N_1667,N_3405);
nor U9506 (N_9506,N_875,N_955);
and U9507 (N_9507,N_309,N_1587);
nand U9508 (N_9508,N_457,N_3932);
or U9509 (N_9509,N_3740,N_1279);
nand U9510 (N_9510,N_807,N_1105);
and U9511 (N_9511,N_779,N_1336);
or U9512 (N_9512,N_336,N_160);
or U9513 (N_9513,N_187,N_1494);
nand U9514 (N_9514,N_4496,N_460);
and U9515 (N_9515,N_1427,N_508);
nand U9516 (N_9516,N_12,N_3504);
or U9517 (N_9517,N_317,N_359);
and U9518 (N_9518,N_321,N_3647);
nand U9519 (N_9519,N_2890,N_2039);
nand U9520 (N_9520,N_575,N_1107);
and U9521 (N_9521,N_342,N_4327);
nor U9522 (N_9522,N_2257,N_1752);
and U9523 (N_9523,N_2609,N_1849);
nor U9524 (N_9524,N_3438,N_1910);
or U9525 (N_9525,N_2658,N_1323);
nand U9526 (N_9526,N_79,N_3073);
nor U9527 (N_9527,N_325,N_3889);
or U9528 (N_9528,N_3170,N_2798);
nor U9529 (N_9529,N_320,N_2275);
or U9530 (N_9530,N_3172,N_2487);
or U9531 (N_9531,N_3242,N_2316);
or U9532 (N_9532,N_3442,N_4357);
and U9533 (N_9533,N_4921,N_789);
nor U9534 (N_9534,N_1836,N_1859);
and U9535 (N_9535,N_1827,N_2623);
or U9536 (N_9536,N_4644,N_2741);
nor U9537 (N_9537,N_834,N_675);
or U9538 (N_9538,N_1353,N_2493);
and U9539 (N_9539,N_2403,N_3935);
nor U9540 (N_9540,N_568,N_2688);
or U9541 (N_9541,N_3512,N_1845);
and U9542 (N_9542,N_1583,N_2595);
nor U9543 (N_9543,N_4016,N_2831);
nor U9544 (N_9544,N_2602,N_2639);
nor U9545 (N_9545,N_1311,N_3566);
nor U9546 (N_9546,N_2198,N_3245);
and U9547 (N_9547,N_4210,N_557);
and U9548 (N_9548,N_3097,N_1299);
nor U9549 (N_9549,N_1352,N_4159);
nand U9550 (N_9550,N_1912,N_2078);
nand U9551 (N_9551,N_470,N_2351);
nand U9552 (N_9552,N_2882,N_3869);
and U9553 (N_9553,N_3589,N_1835);
nor U9554 (N_9554,N_1665,N_3059);
or U9555 (N_9555,N_3640,N_4007);
and U9556 (N_9556,N_3453,N_1734);
or U9557 (N_9557,N_3836,N_816);
and U9558 (N_9558,N_4658,N_1524);
and U9559 (N_9559,N_1565,N_4957);
and U9560 (N_9560,N_495,N_4208);
and U9561 (N_9561,N_2274,N_3705);
nor U9562 (N_9562,N_344,N_4063);
and U9563 (N_9563,N_3244,N_1243);
nand U9564 (N_9564,N_2051,N_4937);
nand U9565 (N_9565,N_815,N_2393);
and U9566 (N_9566,N_311,N_2244);
nor U9567 (N_9567,N_2405,N_2194);
nand U9568 (N_9568,N_2248,N_2364);
nor U9569 (N_9569,N_4461,N_4047);
and U9570 (N_9570,N_3553,N_1816);
and U9571 (N_9571,N_2864,N_792);
nor U9572 (N_9572,N_1051,N_2971);
and U9573 (N_9573,N_1111,N_3460);
or U9574 (N_9574,N_1613,N_2115);
or U9575 (N_9575,N_2033,N_1416);
or U9576 (N_9576,N_2180,N_837);
nand U9577 (N_9577,N_4544,N_5);
nor U9578 (N_9578,N_3895,N_3420);
and U9579 (N_9579,N_1449,N_3760);
nor U9580 (N_9580,N_57,N_2240);
or U9581 (N_9581,N_447,N_2049);
and U9582 (N_9582,N_687,N_3263);
nand U9583 (N_9583,N_1695,N_4757);
nand U9584 (N_9584,N_3501,N_206);
or U9585 (N_9585,N_4618,N_2195);
nor U9586 (N_9586,N_17,N_2153);
or U9587 (N_9587,N_686,N_654);
nor U9588 (N_9588,N_1217,N_1001);
nand U9589 (N_9589,N_66,N_1847);
or U9590 (N_9590,N_2506,N_3263);
nor U9591 (N_9591,N_1522,N_555);
nand U9592 (N_9592,N_465,N_1567);
and U9593 (N_9593,N_3145,N_2704);
nor U9594 (N_9594,N_613,N_3973);
nor U9595 (N_9595,N_1443,N_4495);
or U9596 (N_9596,N_2882,N_2095);
nor U9597 (N_9597,N_3919,N_4754);
and U9598 (N_9598,N_4341,N_3653);
xnor U9599 (N_9599,N_1506,N_3416);
or U9600 (N_9600,N_2757,N_2892);
and U9601 (N_9601,N_4456,N_3684);
xnor U9602 (N_9602,N_2236,N_2750);
nand U9603 (N_9603,N_3230,N_425);
nand U9604 (N_9604,N_1425,N_4482);
and U9605 (N_9605,N_841,N_3188);
nand U9606 (N_9606,N_4176,N_4043);
nand U9607 (N_9607,N_3836,N_2233);
nor U9608 (N_9608,N_1504,N_3777);
nand U9609 (N_9609,N_956,N_3694);
and U9610 (N_9610,N_3887,N_2519);
nor U9611 (N_9611,N_1003,N_4222);
nand U9612 (N_9612,N_1717,N_1110);
and U9613 (N_9613,N_2398,N_4678);
and U9614 (N_9614,N_298,N_3722);
nand U9615 (N_9615,N_194,N_2112);
nor U9616 (N_9616,N_618,N_2243);
and U9617 (N_9617,N_3214,N_4511);
nand U9618 (N_9618,N_4915,N_3905);
nor U9619 (N_9619,N_4782,N_1918);
nor U9620 (N_9620,N_4781,N_1698);
nor U9621 (N_9621,N_105,N_1686);
or U9622 (N_9622,N_4295,N_203);
or U9623 (N_9623,N_3569,N_1799);
nor U9624 (N_9624,N_2419,N_682);
nand U9625 (N_9625,N_593,N_4424);
or U9626 (N_9626,N_3907,N_61);
or U9627 (N_9627,N_1197,N_3070);
or U9628 (N_9628,N_2384,N_3541);
nor U9629 (N_9629,N_3640,N_2689);
or U9630 (N_9630,N_2771,N_3804);
nand U9631 (N_9631,N_3659,N_2835);
and U9632 (N_9632,N_4876,N_1089);
or U9633 (N_9633,N_3282,N_383);
nor U9634 (N_9634,N_1375,N_4587);
nor U9635 (N_9635,N_3548,N_2289);
nor U9636 (N_9636,N_1344,N_982);
or U9637 (N_9637,N_3566,N_2323);
and U9638 (N_9638,N_3028,N_1434);
nand U9639 (N_9639,N_2104,N_3629);
nor U9640 (N_9640,N_2062,N_4013);
nand U9641 (N_9641,N_660,N_2409);
nor U9642 (N_9642,N_1764,N_1052);
nand U9643 (N_9643,N_3021,N_893);
xnor U9644 (N_9644,N_4887,N_2427);
nor U9645 (N_9645,N_4230,N_247);
or U9646 (N_9646,N_2786,N_3179);
nor U9647 (N_9647,N_552,N_2480);
xor U9648 (N_9648,N_2427,N_440);
nor U9649 (N_9649,N_687,N_2328);
or U9650 (N_9650,N_1314,N_1804);
or U9651 (N_9651,N_3004,N_1542);
nand U9652 (N_9652,N_4154,N_645);
xor U9653 (N_9653,N_3772,N_340);
or U9654 (N_9654,N_178,N_762);
and U9655 (N_9655,N_993,N_3957);
nand U9656 (N_9656,N_1138,N_578);
nand U9657 (N_9657,N_3877,N_3242);
nand U9658 (N_9658,N_3823,N_2572);
or U9659 (N_9659,N_675,N_1346);
nor U9660 (N_9660,N_4730,N_582);
nor U9661 (N_9661,N_1662,N_3013);
nor U9662 (N_9662,N_4676,N_4527);
or U9663 (N_9663,N_4375,N_3832);
nand U9664 (N_9664,N_2928,N_201);
and U9665 (N_9665,N_4607,N_2835);
or U9666 (N_9666,N_1264,N_1889);
and U9667 (N_9667,N_2426,N_4232);
and U9668 (N_9668,N_2153,N_3286);
or U9669 (N_9669,N_1004,N_3255);
and U9670 (N_9670,N_4507,N_2585);
nand U9671 (N_9671,N_2771,N_2720);
nand U9672 (N_9672,N_3500,N_3644);
nand U9673 (N_9673,N_1275,N_256);
nor U9674 (N_9674,N_3963,N_1072);
and U9675 (N_9675,N_2258,N_2122);
or U9676 (N_9676,N_4921,N_3202);
and U9677 (N_9677,N_2849,N_4323);
nor U9678 (N_9678,N_4364,N_2966);
nand U9679 (N_9679,N_3615,N_571);
nand U9680 (N_9680,N_3491,N_4514);
or U9681 (N_9681,N_4404,N_1252);
or U9682 (N_9682,N_4171,N_3699);
or U9683 (N_9683,N_1423,N_1291);
and U9684 (N_9684,N_1524,N_1223);
or U9685 (N_9685,N_4823,N_1651);
nor U9686 (N_9686,N_3090,N_1003);
and U9687 (N_9687,N_473,N_4625);
nand U9688 (N_9688,N_3138,N_1923);
nor U9689 (N_9689,N_1931,N_2764);
and U9690 (N_9690,N_1223,N_1259);
nand U9691 (N_9691,N_3118,N_2500);
and U9692 (N_9692,N_3879,N_2500);
and U9693 (N_9693,N_2048,N_248);
nor U9694 (N_9694,N_3397,N_4291);
nand U9695 (N_9695,N_3706,N_4089);
nand U9696 (N_9696,N_821,N_4532);
and U9697 (N_9697,N_4231,N_426);
nand U9698 (N_9698,N_1721,N_1398);
and U9699 (N_9699,N_4306,N_4077);
or U9700 (N_9700,N_1253,N_2879);
nand U9701 (N_9701,N_2570,N_3324);
xnor U9702 (N_9702,N_3447,N_3492);
or U9703 (N_9703,N_537,N_3375);
or U9704 (N_9704,N_3178,N_3867);
nand U9705 (N_9705,N_2290,N_4735);
or U9706 (N_9706,N_2024,N_3174);
xnor U9707 (N_9707,N_1954,N_3726);
nand U9708 (N_9708,N_746,N_3133);
and U9709 (N_9709,N_4696,N_1321);
nor U9710 (N_9710,N_274,N_4386);
or U9711 (N_9711,N_1884,N_3256);
nor U9712 (N_9712,N_354,N_3015);
and U9713 (N_9713,N_4308,N_867);
xor U9714 (N_9714,N_3582,N_1392);
nor U9715 (N_9715,N_2531,N_2121);
or U9716 (N_9716,N_465,N_2063);
nand U9717 (N_9717,N_683,N_846);
or U9718 (N_9718,N_1792,N_1322);
nor U9719 (N_9719,N_1058,N_549);
nand U9720 (N_9720,N_3851,N_528);
nand U9721 (N_9721,N_3835,N_1307);
and U9722 (N_9722,N_143,N_1007);
and U9723 (N_9723,N_28,N_3876);
and U9724 (N_9724,N_1559,N_3096);
or U9725 (N_9725,N_3199,N_2094);
and U9726 (N_9726,N_4599,N_4890);
and U9727 (N_9727,N_466,N_173);
or U9728 (N_9728,N_4429,N_1198);
nand U9729 (N_9729,N_1296,N_4252);
nor U9730 (N_9730,N_2169,N_2946);
or U9731 (N_9731,N_37,N_1610);
nand U9732 (N_9732,N_160,N_530);
and U9733 (N_9733,N_1217,N_4816);
or U9734 (N_9734,N_4443,N_3841);
or U9735 (N_9735,N_2806,N_1247);
and U9736 (N_9736,N_3729,N_3696);
and U9737 (N_9737,N_1350,N_1555);
nor U9738 (N_9738,N_253,N_1358);
nand U9739 (N_9739,N_3397,N_585);
nor U9740 (N_9740,N_3688,N_1799);
and U9741 (N_9741,N_3426,N_880);
and U9742 (N_9742,N_4049,N_99);
or U9743 (N_9743,N_2567,N_3614);
and U9744 (N_9744,N_2275,N_2877);
and U9745 (N_9745,N_3407,N_2239);
nand U9746 (N_9746,N_3555,N_570);
and U9747 (N_9747,N_3821,N_988);
or U9748 (N_9748,N_4469,N_2290);
nor U9749 (N_9749,N_2745,N_3602);
nor U9750 (N_9750,N_4633,N_4744);
nor U9751 (N_9751,N_3347,N_667);
and U9752 (N_9752,N_4720,N_997);
or U9753 (N_9753,N_2079,N_53);
nor U9754 (N_9754,N_3104,N_4498);
nor U9755 (N_9755,N_3520,N_4437);
nor U9756 (N_9756,N_1978,N_2444);
xnor U9757 (N_9757,N_474,N_2297);
or U9758 (N_9758,N_1030,N_4849);
nand U9759 (N_9759,N_916,N_77);
nand U9760 (N_9760,N_869,N_2935);
nand U9761 (N_9761,N_871,N_4310);
or U9762 (N_9762,N_4777,N_489);
nand U9763 (N_9763,N_4086,N_1741);
and U9764 (N_9764,N_1480,N_4994);
and U9765 (N_9765,N_1215,N_3220);
nor U9766 (N_9766,N_4441,N_4717);
or U9767 (N_9767,N_1238,N_2687);
or U9768 (N_9768,N_4576,N_2604);
nand U9769 (N_9769,N_2054,N_1431);
or U9770 (N_9770,N_3758,N_1910);
nor U9771 (N_9771,N_2151,N_3100);
xor U9772 (N_9772,N_258,N_3440);
xnor U9773 (N_9773,N_1245,N_3425);
or U9774 (N_9774,N_1422,N_2827);
nand U9775 (N_9775,N_383,N_2650);
nor U9776 (N_9776,N_330,N_1055);
or U9777 (N_9777,N_399,N_4100);
and U9778 (N_9778,N_2393,N_346);
and U9779 (N_9779,N_786,N_1124);
nand U9780 (N_9780,N_608,N_1965);
nand U9781 (N_9781,N_4018,N_1956);
nor U9782 (N_9782,N_3822,N_2107);
or U9783 (N_9783,N_4315,N_3214);
or U9784 (N_9784,N_624,N_395);
and U9785 (N_9785,N_1156,N_965);
and U9786 (N_9786,N_4330,N_2704);
and U9787 (N_9787,N_3846,N_1807);
and U9788 (N_9788,N_3331,N_4129);
or U9789 (N_9789,N_198,N_17);
and U9790 (N_9790,N_39,N_4092);
or U9791 (N_9791,N_4807,N_4409);
nor U9792 (N_9792,N_3352,N_345);
nor U9793 (N_9793,N_171,N_3287);
or U9794 (N_9794,N_2038,N_3338);
nor U9795 (N_9795,N_2695,N_615);
nand U9796 (N_9796,N_2172,N_4451);
nor U9797 (N_9797,N_4937,N_1034);
and U9798 (N_9798,N_3737,N_2469);
or U9799 (N_9799,N_426,N_2987);
nand U9800 (N_9800,N_2062,N_1742);
or U9801 (N_9801,N_3967,N_2957);
nand U9802 (N_9802,N_3149,N_613);
nor U9803 (N_9803,N_3169,N_1464);
nand U9804 (N_9804,N_898,N_4500);
nand U9805 (N_9805,N_3359,N_848);
nand U9806 (N_9806,N_2654,N_1969);
or U9807 (N_9807,N_3799,N_4278);
and U9808 (N_9808,N_3708,N_452);
or U9809 (N_9809,N_3313,N_1927);
and U9810 (N_9810,N_1450,N_168);
nand U9811 (N_9811,N_3387,N_1263);
nand U9812 (N_9812,N_1686,N_1705);
and U9813 (N_9813,N_2932,N_3044);
nor U9814 (N_9814,N_1558,N_4616);
nand U9815 (N_9815,N_2639,N_4442);
nor U9816 (N_9816,N_3858,N_273);
and U9817 (N_9817,N_1673,N_1512);
nand U9818 (N_9818,N_2628,N_3477);
and U9819 (N_9819,N_4925,N_1454);
and U9820 (N_9820,N_91,N_89);
and U9821 (N_9821,N_3790,N_3297);
nor U9822 (N_9822,N_1712,N_4276);
or U9823 (N_9823,N_2312,N_2432);
and U9824 (N_9824,N_1688,N_4088);
nand U9825 (N_9825,N_3973,N_377);
and U9826 (N_9826,N_1533,N_154);
nor U9827 (N_9827,N_2671,N_3205);
xnor U9828 (N_9828,N_1802,N_785);
nor U9829 (N_9829,N_4212,N_4383);
nand U9830 (N_9830,N_2450,N_309);
xnor U9831 (N_9831,N_2486,N_726);
and U9832 (N_9832,N_3433,N_3846);
or U9833 (N_9833,N_3864,N_4828);
nor U9834 (N_9834,N_2315,N_2569);
nand U9835 (N_9835,N_3614,N_2839);
and U9836 (N_9836,N_4162,N_9);
nor U9837 (N_9837,N_2735,N_1629);
and U9838 (N_9838,N_4415,N_4577);
nor U9839 (N_9839,N_2624,N_608);
nor U9840 (N_9840,N_4507,N_1028);
nor U9841 (N_9841,N_2984,N_3260);
or U9842 (N_9842,N_3798,N_2562);
and U9843 (N_9843,N_1036,N_3553);
and U9844 (N_9844,N_3365,N_4914);
nor U9845 (N_9845,N_3194,N_3007);
nor U9846 (N_9846,N_1038,N_3592);
and U9847 (N_9847,N_438,N_2621);
nand U9848 (N_9848,N_380,N_1668);
and U9849 (N_9849,N_1742,N_2207);
or U9850 (N_9850,N_2653,N_2738);
and U9851 (N_9851,N_1454,N_3576);
and U9852 (N_9852,N_2877,N_3221);
or U9853 (N_9853,N_2991,N_2111);
or U9854 (N_9854,N_2453,N_1133);
nand U9855 (N_9855,N_3366,N_459);
nand U9856 (N_9856,N_2119,N_1108);
and U9857 (N_9857,N_1855,N_1424);
nand U9858 (N_9858,N_2200,N_3479);
nor U9859 (N_9859,N_3945,N_624);
or U9860 (N_9860,N_4030,N_1151);
and U9861 (N_9861,N_3372,N_1552);
or U9862 (N_9862,N_2816,N_3811);
or U9863 (N_9863,N_3100,N_1062);
nand U9864 (N_9864,N_2040,N_3884);
or U9865 (N_9865,N_3173,N_4009);
and U9866 (N_9866,N_4674,N_1068);
nor U9867 (N_9867,N_4447,N_3478);
nand U9868 (N_9868,N_4876,N_3919);
nand U9869 (N_9869,N_1654,N_3931);
nand U9870 (N_9870,N_1076,N_4332);
and U9871 (N_9871,N_3916,N_2952);
nor U9872 (N_9872,N_697,N_2903);
nor U9873 (N_9873,N_3973,N_1458);
or U9874 (N_9874,N_2486,N_2810);
or U9875 (N_9875,N_2265,N_3996);
and U9876 (N_9876,N_1916,N_1292);
nor U9877 (N_9877,N_999,N_3294);
nand U9878 (N_9878,N_3532,N_3315);
nand U9879 (N_9879,N_1347,N_2385);
and U9880 (N_9880,N_1398,N_2339);
or U9881 (N_9881,N_211,N_3836);
nand U9882 (N_9882,N_3514,N_2667);
and U9883 (N_9883,N_3377,N_2844);
nor U9884 (N_9884,N_3775,N_1213);
nand U9885 (N_9885,N_2388,N_3223);
nand U9886 (N_9886,N_3941,N_1814);
and U9887 (N_9887,N_327,N_4678);
and U9888 (N_9888,N_2493,N_1437);
or U9889 (N_9889,N_4466,N_4528);
nand U9890 (N_9890,N_4348,N_4622);
nand U9891 (N_9891,N_2496,N_539);
nor U9892 (N_9892,N_743,N_3511);
or U9893 (N_9893,N_1870,N_449);
nor U9894 (N_9894,N_3497,N_4972);
nand U9895 (N_9895,N_4858,N_991);
nor U9896 (N_9896,N_2545,N_498);
nand U9897 (N_9897,N_4029,N_2906);
and U9898 (N_9898,N_4729,N_869);
or U9899 (N_9899,N_2242,N_3171);
nor U9900 (N_9900,N_227,N_500);
nand U9901 (N_9901,N_2621,N_2248);
nor U9902 (N_9902,N_2086,N_4090);
nor U9903 (N_9903,N_4919,N_3450);
or U9904 (N_9904,N_1265,N_4067);
nor U9905 (N_9905,N_2273,N_3980);
nand U9906 (N_9906,N_1940,N_1383);
nor U9907 (N_9907,N_2254,N_2527);
nor U9908 (N_9908,N_803,N_992);
nor U9909 (N_9909,N_3936,N_4589);
nand U9910 (N_9910,N_2144,N_4568);
nand U9911 (N_9911,N_2047,N_3142);
and U9912 (N_9912,N_2946,N_2387);
nand U9913 (N_9913,N_1899,N_3382);
nor U9914 (N_9914,N_1661,N_91);
nor U9915 (N_9915,N_3279,N_2304);
nand U9916 (N_9916,N_4346,N_4413);
and U9917 (N_9917,N_3295,N_4522);
nand U9918 (N_9918,N_4198,N_3598);
or U9919 (N_9919,N_2208,N_3835);
and U9920 (N_9920,N_1813,N_24);
nand U9921 (N_9921,N_1139,N_4906);
and U9922 (N_9922,N_327,N_1014);
nand U9923 (N_9923,N_2406,N_421);
nor U9924 (N_9924,N_565,N_1526);
nand U9925 (N_9925,N_4673,N_4982);
nor U9926 (N_9926,N_2079,N_1036);
or U9927 (N_9927,N_203,N_1535);
nor U9928 (N_9928,N_1800,N_3844);
or U9929 (N_9929,N_3512,N_829);
and U9930 (N_9930,N_4715,N_4409);
nor U9931 (N_9931,N_482,N_474);
and U9932 (N_9932,N_691,N_2440);
and U9933 (N_9933,N_4260,N_1168);
nand U9934 (N_9934,N_2644,N_2104);
or U9935 (N_9935,N_1947,N_2592);
nand U9936 (N_9936,N_2724,N_1540);
nand U9937 (N_9937,N_3022,N_4517);
nor U9938 (N_9938,N_3741,N_594);
nor U9939 (N_9939,N_2560,N_2537);
xnor U9940 (N_9940,N_876,N_4196);
xor U9941 (N_9941,N_186,N_373);
nor U9942 (N_9942,N_380,N_4265);
and U9943 (N_9943,N_3343,N_3431);
or U9944 (N_9944,N_4973,N_1845);
and U9945 (N_9945,N_3820,N_1259);
xnor U9946 (N_9946,N_2367,N_2245);
nor U9947 (N_9947,N_1935,N_1470);
and U9948 (N_9948,N_1667,N_2937);
nor U9949 (N_9949,N_4115,N_1084);
or U9950 (N_9950,N_636,N_1359);
or U9951 (N_9951,N_4132,N_1559);
and U9952 (N_9952,N_848,N_3777);
or U9953 (N_9953,N_4435,N_1420);
nor U9954 (N_9954,N_1097,N_2317);
or U9955 (N_9955,N_1890,N_2685);
nand U9956 (N_9956,N_3827,N_1012);
or U9957 (N_9957,N_87,N_4876);
nand U9958 (N_9958,N_1352,N_4160);
or U9959 (N_9959,N_2337,N_1606);
or U9960 (N_9960,N_632,N_2860);
nor U9961 (N_9961,N_3942,N_4758);
nor U9962 (N_9962,N_1107,N_4844);
nor U9963 (N_9963,N_4929,N_1772);
or U9964 (N_9964,N_225,N_2107);
nor U9965 (N_9965,N_315,N_1311);
and U9966 (N_9966,N_3410,N_3910);
or U9967 (N_9967,N_3748,N_2179);
nor U9968 (N_9968,N_3936,N_4932);
nor U9969 (N_9969,N_896,N_4612);
and U9970 (N_9970,N_4358,N_486);
or U9971 (N_9971,N_117,N_3125);
or U9972 (N_9972,N_2450,N_1429);
or U9973 (N_9973,N_3067,N_2182);
and U9974 (N_9974,N_2989,N_4215);
and U9975 (N_9975,N_826,N_2058);
nor U9976 (N_9976,N_2692,N_415);
nand U9977 (N_9977,N_646,N_3543);
nand U9978 (N_9978,N_1408,N_3660);
nor U9979 (N_9979,N_3964,N_2210);
nor U9980 (N_9980,N_4441,N_757);
or U9981 (N_9981,N_1767,N_3057);
nand U9982 (N_9982,N_3733,N_2187);
nor U9983 (N_9983,N_536,N_2188);
or U9984 (N_9984,N_4035,N_4132);
xnor U9985 (N_9985,N_3327,N_1782);
and U9986 (N_9986,N_1638,N_4776);
and U9987 (N_9987,N_3172,N_2753);
and U9988 (N_9988,N_578,N_4406);
nor U9989 (N_9989,N_1483,N_855);
or U9990 (N_9990,N_4611,N_3619);
nor U9991 (N_9991,N_681,N_550);
nand U9992 (N_9992,N_1806,N_3631);
nand U9993 (N_9993,N_318,N_4047);
or U9994 (N_9994,N_3850,N_2737);
nor U9995 (N_9995,N_3375,N_2143);
and U9996 (N_9996,N_3377,N_1148);
or U9997 (N_9997,N_2054,N_3251);
nor U9998 (N_9998,N_3766,N_1527);
nor U9999 (N_9999,N_1236,N_1607);
xor U10000 (N_10000,N_7507,N_9868);
nand U10001 (N_10001,N_9209,N_9346);
nand U10002 (N_10002,N_5818,N_6078);
nor U10003 (N_10003,N_8087,N_9797);
nor U10004 (N_10004,N_9656,N_5293);
nor U10005 (N_10005,N_6392,N_9618);
nor U10006 (N_10006,N_8163,N_8833);
xor U10007 (N_10007,N_8721,N_5905);
and U10008 (N_10008,N_7020,N_8762);
and U10009 (N_10009,N_8118,N_5536);
or U10010 (N_10010,N_9224,N_7904);
nor U10011 (N_10011,N_5459,N_9244);
nor U10012 (N_10012,N_5550,N_5594);
and U10013 (N_10013,N_7070,N_6575);
nand U10014 (N_10014,N_9768,N_8270);
or U10015 (N_10015,N_7099,N_8634);
and U10016 (N_10016,N_6811,N_9642);
nand U10017 (N_10017,N_5815,N_9643);
nor U10018 (N_10018,N_9315,N_5476);
xnor U10019 (N_10019,N_7515,N_8298);
nor U10020 (N_10020,N_7999,N_7236);
and U10021 (N_10021,N_7519,N_5682);
nand U10022 (N_10022,N_8048,N_5795);
and U10023 (N_10023,N_5745,N_7976);
or U10024 (N_10024,N_5358,N_7528);
or U10025 (N_10025,N_9197,N_6063);
nor U10026 (N_10026,N_7531,N_9969);
and U10027 (N_10027,N_6974,N_9192);
xor U10028 (N_10028,N_7693,N_9886);
nand U10029 (N_10029,N_6466,N_6071);
nand U10030 (N_10030,N_5457,N_9329);
nor U10031 (N_10031,N_6668,N_7392);
or U10032 (N_10032,N_8247,N_9143);
or U10033 (N_10033,N_5100,N_9781);
or U10034 (N_10034,N_8815,N_7607);
nor U10035 (N_10035,N_5284,N_9906);
nor U10036 (N_10036,N_7382,N_5409);
and U10037 (N_10037,N_5396,N_7019);
and U10038 (N_10038,N_6124,N_9857);
and U10039 (N_10039,N_5556,N_6039);
nand U10040 (N_10040,N_8290,N_9903);
or U10041 (N_10041,N_6086,N_5881);
nand U10042 (N_10042,N_8932,N_9021);
or U10043 (N_10043,N_6253,N_6195);
nand U10044 (N_10044,N_6228,N_8486);
or U10045 (N_10045,N_5047,N_7104);
and U10046 (N_10046,N_5912,N_8489);
nand U10047 (N_10047,N_9310,N_6970);
nor U10048 (N_10048,N_9740,N_8205);
or U10049 (N_10049,N_5207,N_9974);
xnor U10050 (N_10050,N_6802,N_8312);
or U10051 (N_10051,N_9145,N_8481);
or U10052 (N_10052,N_6881,N_6284);
or U10053 (N_10053,N_6452,N_5346);
nand U10054 (N_10054,N_8672,N_9045);
and U10055 (N_10055,N_7297,N_7932);
or U10056 (N_10056,N_5723,N_6153);
and U10057 (N_10057,N_8367,N_9251);
and U10058 (N_10058,N_8374,N_5640);
nor U10059 (N_10059,N_8222,N_9882);
or U10060 (N_10060,N_8111,N_8327);
nor U10061 (N_10061,N_8835,N_5230);
nand U10062 (N_10062,N_6029,N_9478);
and U10063 (N_10063,N_9975,N_7597);
and U10064 (N_10064,N_8477,N_6088);
and U10065 (N_10065,N_9535,N_5634);
xnor U10066 (N_10066,N_7547,N_5338);
nor U10067 (N_10067,N_7919,N_8994);
and U10068 (N_10068,N_6880,N_9429);
and U10069 (N_10069,N_7439,N_7734);
nand U10070 (N_10070,N_5874,N_8878);
nand U10071 (N_10071,N_6479,N_6994);
and U10072 (N_10072,N_5071,N_9439);
and U10073 (N_10073,N_7376,N_7827);
nand U10074 (N_10074,N_7492,N_6131);
nand U10075 (N_10075,N_5502,N_9074);
and U10076 (N_10076,N_6354,N_8902);
nand U10077 (N_10077,N_8403,N_6254);
or U10078 (N_10078,N_5810,N_8010);
or U10079 (N_10079,N_5208,N_6788);
or U10080 (N_10080,N_7645,N_6932);
or U10081 (N_10081,N_8814,N_9304);
nor U10082 (N_10082,N_8873,N_5929);
or U10083 (N_10083,N_7961,N_7143);
and U10084 (N_10084,N_8775,N_5983);
nand U10085 (N_10085,N_7161,N_9409);
nand U10086 (N_10086,N_7270,N_5703);
nand U10087 (N_10087,N_6281,N_7227);
nor U10088 (N_10088,N_9722,N_9313);
nor U10089 (N_10089,N_5057,N_9621);
or U10090 (N_10090,N_7307,N_9416);
or U10091 (N_10091,N_9543,N_6931);
nand U10092 (N_10092,N_9606,N_5359);
xnor U10093 (N_10093,N_6004,N_9691);
or U10094 (N_10094,N_8852,N_7621);
and U10095 (N_10095,N_8934,N_7466);
nor U10096 (N_10096,N_5177,N_9807);
and U10097 (N_10097,N_5577,N_9255);
nor U10098 (N_10098,N_5507,N_5258);
and U10099 (N_10099,N_7012,N_6859);
and U10100 (N_10100,N_9909,N_8246);
or U10101 (N_10101,N_5834,N_5781);
or U10102 (N_10102,N_9679,N_6112);
and U10103 (N_10103,N_7430,N_6629);
nand U10104 (N_10104,N_6902,N_7811);
or U10105 (N_10105,N_6398,N_9619);
or U10106 (N_10106,N_5835,N_8889);
and U10107 (N_10107,N_7194,N_5349);
and U10108 (N_10108,N_5618,N_8777);
or U10109 (N_10109,N_5959,N_9765);
xnor U10110 (N_10110,N_6965,N_5751);
nand U10111 (N_10111,N_7577,N_5650);
and U10112 (N_10112,N_9908,N_6408);
and U10113 (N_10113,N_9250,N_6335);
nor U10114 (N_10114,N_7663,N_8953);
and U10115 (N_10115,N_8514,N_6337);
nand U10116 (N_10116,N_9047,N_7184);
and U10117 (N_10117,N_8359,N_5218);
or U10118 (N_10118,N_6765,N_8865);
and U10119 (N_10119,N_7209,N_6371);
nor U10120 (N_10120,N_8068,N_5360);
nand U10121 (N_10121,N_8159,N_8664);
or U10122 (N_10122,N_9595,N_5681);
nand U10123 (N_10123,N_6106,N_5001);
and U10124 (N_10124,N_7578,N_5078);
and U10125 (N_10125,N_8871,N_6600);
and U10126 (N_10126,N_6935,N_6647);
nor U10127 (N_10127,N_7892,N_8131);
nand U10128 (N_10128,N_7694,N_8513);
nand U10129 (N_10129,N_8862,N_5730);
nor U10130 (N_10130,N_7896,N_8002);
nand U10131 (N_10131,N_8909,N_8135);
or U10132 (N_10132,N_7302,N_6735);
nand U10133 (N_10133,N_9476,N_6971);
and U10134 (N_10134,N_8425,N_5309);
xnor U10135 (N_10135,N_6294,N_7927);
and U10136 (N_10136,N_8348,N_9944);
and U10137 (N_10137,N_7698,N_9907);
nor U10138 (N_10138,N_6576,N_7167);
nor U10139 (N_10139,N_5471,N_5626);
or U10140 (N_10140,N_5696,N_9718);
nor U10141 (N_10141,N_6197,N_6766);
and U10142 (N_10142,N_7922,N_9484);
and U10143 (N_10143,N_7786,N_6486);
and U10144 (N_10144,N_5739,N_9075);
or U10145 (N_10145,N_9587,N_5320);
nand U10146 (N_10146,N_7991,N_5060);
or U10147 (N_10147,N_9692,N_8504);
and U10148 (N_10148,N_9261,N_7342);
nor U10149 (N_10149,N_9319,N_7863);
nand U10150 (N_10150,N_6906,N_5294);
nand U10151 (N_10151,N_5203,N_9254);
and U10152 (N_10152,N_8628,N_5805);
nor U10153 (N_10153,N_5165,N_6706);
or U10154 (N_10154,N_8987,N_7052);
or U10155 (N_10155,N_5351,N_9537);
and U10156 (N_10156,N_7110,N_9294);
nand U10157 (N_10157,N_5375,N_6862);
nor U10158 (N_10158,N_8299,N_9381);
nor U10159 (N_10159,N_5106,N_7848);
nand U10160 (N_10160,N_9242,N_9308);
nor U10161 (N_10161,N_7544,N_6885);
and U10162 (N_10162,N_7906,N_9811);
nor U10163 (N_10163,N_8611,N_6440);
nor U10164 (N_10164,N_5576,N_9555);
nand U10165 (N_10165,N_7898,N_6443);
or U10166 (N_10166,N_6105,N_6526);
and U10167 (N_10167,N_6055,N_6665);
or U10168 (N_10168,N_8378,N_9931);
or U10169 (N_10169,N_7945,N_6857);
or U10170 (N_10170,N_6879,N_8686);
or U10171 (N_10171,N_6468,N_5825);
nor U10172 (N_10172,N_5738,N_7047);
and U10173 (N_10173,N_7969,N_9675);
or U10174 (N_10174,N_7217,N_5123);
or U10175 (N_10175,N_8052,N_7650);
nand U10176 (N_10176,N_7814,N_9227);
or U10177 (N_10177,N_9672,N_7196);
nand U10178 (N_10178,N_6980,N_5121);
or U10179 (N_10179,N_7718,N_5092);
nor U10180 (N_10180,N_5603,N_5010);
and U10181 (N_10181,N_6239,N_9876);
nand U10182 (N_10182,N_6400,N_7576);
and U10183 (N_10183,N_8322,N_6410);
or U10184 (N_10184,N_9548,N_8960);
or U10185 (N_10185,N_5674,N_7114);
and U10186 (N_10186,N_5002,N_7797);
and U10187 (N_10187,N_7452,N_6393);
nor U10188 (N_10188,N_6651,N_7843);
nor U10189 (N_10189,N_5924,N_6381);
or U10190 (N_10190,N_8980,N_6843);
and U10191 (N_10191,N_5018,N_9785);
and U10192 (N_10192,N_9126,N_5153);
nor U10193 (N_10193,N_8985,N_5679);
and U10194 (N_10194,N_8619,N_8482);
nand U10195 (N_10195,N_7781,N_5026);
nand U10196 (N_10196,N_6511,N_7000);
nand U10197 (N_10197,N_5788,N_5257);
and U10198 (N_10198,N_8394,N_5438);
nand U10199 (N_10199,N_9165,N_7008);
or U10200 (N_10200,N_9370,N_8066);
nand U10201 (N_10201,N_8726,N_9398);
and U10202 (N_10202,N_6134,N_7353);
and U10203 (N_10203,N_9965,N_7890);
and U10204 (N_10204,N_8910,N_5544);
or U10205 (N_10205,N_6867,N_7418);
nand U10206 (N_10206,N_8062,N_7238);
or U10207 (N_10207,N_5567,N_5006);
or U10208 (N_10208,N_9096,N_8741);
nand U10209 (N_10209,N_6723,N_9832);
nor U10210 (N_10210,N_5316,N_9467);
nand U10211 (N_10211,N_5098,N_9554);
and U10212 (N_10212,N_5128,N_5821);
or U10213 (N_10213,N_7351,N_5385);
nor U10214 (N_10214,N_5566,N_7673);
and U10215 (N_10215,N_9497,N_7431);
and U10216 (N_10216,N_9879,N_9410);
nor U10217 (N_10217,N_8340,N_9697);
and U10218 (N_10218,N_7958,N_8140);
nand U10219 (N_10219,N_9479,N_5202);
or U10220 (N_10220,N_6672,N_6169);
or U10221 (N_10221,N_6663,N_8714);
nor U10222 (N_10222,N_5324,N_6758);
or U10223 (N_10223,N_8832,N_8461);
and U10224 (N_10224,N_5042,N_5247);
and U10225 (N_10225,N_5491,N_9446);
and U10226 (N_10226,N_5523,N_5132);
and U10227 (N_10227,N_7970,N_7281);
nand U10228 (N_10228,N_6151,N_5463);
or U10229 (N_10229,N_6777,N_7593);
nand U10230 (N_10230,N_8644,N_6907);
and U10231 (N_10231,N_6554,N_7579);
nor U10232 (N_10232,N_5210,N_7442);
or U10233 (N_10233,N_9359,N_6127);
nand U10234 (N_10234,N_9996,N_9744);
nor U10235 (N_10235,N_9417,N_8373);
and U10236 (N_10236,N_5704,N_7674);
xnor U10237 (N_10237,N_6451,N_9150);
and U10238 (N_10238,N_7926,N_7423);
or U10239 (N_10239,N_5557,N_6904);
and U10240 (N_10240,N_6241,N_5558);
nand U10241 (N_10241,N_6545,N_9085);
xor U10242 (N_10242,N_5472,N_6051);
nor U10243 (N_10243,N_7975,N_7344);
xor U10244 (N_10244,N_6525,N_9542);
nor U10245 (N_10245,N_6014,N_5740);
nand U10246 (N_10246,N_9508,N_8153);
and U10247 (N_10247,N_8596,N_6924);
nand U10248 (N_10248,N_6521,N_5794);
nand U10249 (N_10249,N_6805,N_5447);
or U10250 (N_10250,N_7195,N_7461);
xor U10251 (N_10251,N_7352,N_7659);
nand U10252 (N_10252,N_8931,N_9930);
or U10253 (N_10253,N_9447,N_7875);
nor U10254 (N_10254,N_6459,N_8470);
and U10255 (N_10255,N_6341,N_5407);
and U10256 (N_10256,N_7065,N_5149);
nor U10257 (N_10257,N_6161,N_6616);
xnor U10258 (N_10258,N_5148,N_5382);
and U10259 (N_10259,N_7913,N_7733);
nor U10260 (N_10260,N_7299,N_9959);
nor U10261 (N_10261,N_9659,N_6117);
nand U10262 (N_10262,N_8090,N_8431);
nor U10263 (N_10263,N_6181,N_9665);
nand U10264 (N_10264,N_5999,N_8521);
nand U10265 (N_10265,N_8665,N_5553);
nor U10266 (N_10266,N_5446,N_8105);
or U10267 (N_10267,N_9057,N_5237);
nor U10268 (N_10268,N_6588,N_7974);
nor U10269 (N_10269,N_8620,N_8998);
and U10270 (N_10270,N_5778,N_6355);
or U10271 (N_10271,N_7883,N_8175);
nor U10272 (N_10272,N_6952,N_5226);
nand U10273 (N_10273,N_8187,N_6707);
xor U10274 (N_10274,N_8297,N_7041);
nor U10275 (N_10275,N_7822,N_9772);
or U10276 (N_10276,N_8911,N_7518);
and U10277 (N_10277,N_7247,N_5125);
and U10278 (N_10278,N_7244,N_8345);
and U10279 (N_10279,N_6348,N_5314);
nor U10280 (N_10280,N_6426,N_8165);
nor U10281 (N_10281,N_5059,N_6065);
and U10282 (N_10282,N_9574,N_5055);
nand U10283 (N_10283,N_8724,N_5198);
and U10284 (N_10284,N_6139,N_9490);
or U10285 (N_10285,N_8447,N_7510);
or U10286 (N_10286,N_9133,N_8767);
or U10287 (N_10287,N_7998,N_9644);
and U10288 (N_10288,N_8974,N_5624);
or U10289 (N_10289,N_8778,N_5496);
nand U10290 (N_10290,N_7754,N_8361);
nand U10291 (N_10291,N_9204,N_5058);
nand U10292 (N_10292,N_5790,N_8480);
nand U10293 (N_10293,N_5233,N_8209);
nor U10294 (N_10294,N_7385,N_7314);
or U10295 (N_10295,N_5942,N_6028);
nor U10296 (N_10296,N_7657,N_5901);
nand U10297 (N_10297,N_5819,N_8914);
nor U10298 (N_10298,N_8988,N_5570);
nand U10299 (N_10299,N_6357,N_6512);
or U10300 (N_10300,N_7661,N_7941);
and U10301 (N_10301,N_5973,N_6091);
and U10302 (N_10302,N_7695,N_8956);
nand U10303 (N_10303,N_8208,N_7769);
nor U10304 (N_10304,N_6048,N_5826);
or U10305 (N_10305,N_9966,N_6547);
or U10306 (N_10306,N_6611,N_6298);
and U10307 (N_10307,N_8607,N_5986);
or U10308 (N_10308,N_5285,N_5486);
nand U10309 (N_10309,N_5242,N_6598);
nor U10310 (N_10310,N_9711,N_6058);
nor U10311 (N_10311,N_7018,N_9696);
or U10312 (N_10312,N_7648,N_7766);
nand U10313 (N_10313,N_6009,N_5525);
and U10314 (N_10314,N_7933,N_8490);
or U10315 (N_10315,N_8530,N_8785);
nor U10316 (N_10316,N_5381,N_7680);
nand U10317 (N_10317,N_6311,N_7756);
nand U10318 (N_10318,N_9229,N_9688);
nand U10319 (N_10319,N_7239,N_8696);
nand U10320 (N_10320,N_5114,N_7497);
and U10321 (N_10321,N_7292,N_5076);
nand U10322 (N_10322,N_9686,N_6043);
and U10323 (N_10323,N_9101,N_6945);
xnor U10324 (N_10324,N_8275,N_8642);
nor U10325 (N_10325,N_5526,N_7658);
nor U10326 (N_10326,N_7949,N_8540);
nand U10327 (N_10327,N_8827,N_8751);
nor U10328 (N_10328,N_5948,N_6995);
nor U10329 (N_10329,N_9915,N_9088);
or U10330 (N_10330,N_6810,N_7714);
or U10331 (N_10331,N_7152,N_5261);
nor U10332 (N_10332,N_8983,N_5880);
and U10333 (N_10333,N_9758,N_6478);
nand U10334 (N_10334,N_5764,N_6428);
nor U10335 (N_10335,N_5155,N_8479);
and U10336 (N_10336,N_6204,N_5754);
nand U10337 (N_10337,N_6615,N_9211);
nand U10338 (N_10338,N_5717,N_5775);
nor U10339 (N_10339,N_7044,N_7048);
nand U10340 (N_10340,N_5994,N_6539);
nor U10341 (N_10341,N_9703,N_9993);
and U10342 (N_10342,N_9431,N_6309);
or U10343 (N_10343,N_5938,N_6352);
or U10344 (N_10344,N_8615,N_6940);
or U10345 (N_10345,N_5964,N_6081);
or U10346 (N_10346,N_9015,N_5926);
nand U10347 (N_10347,N_8176,N_6704);
and U10348 (N_10348,N_9817,N_8429);
and U10349 (N_10349,N_7891,N_7634);
nor U10350 (N_10350,N_7076,N_6774);
or U10351 (N_10351,N_5753,N_9103);
and U10352 (N_10352,N_9199,N_8734);
and U10353 (N_10353,N_9342,N_9472);
and U10354 (N_10354,N_8973,N_9598);
nor U10355 (N_10355,N_8574,N_5801);
nand U10356 (N_10356,N_8263,N_7681);
and U10357 (N_10357,N_5737,N_7583);
nand U10358 (N_10358,N_5061,N_8295);
nor U10359 (N_10359,N_8346,N_5464);
or U10360 (N_10360,N_7463,N_8905);
and U10361 (N_10361,N_9335,N_9233);
and U10362 (N_10362,N_6515,N_6760);
or U10363 (N_10363,N_7062,N_5399);
nor U10364 (N_10364,N_6927,N_6771);
and U10365 (N_10365,N_5126,N_8660);
xor U10366 (N_10366,N_8203,N_8915);
nand U10367 (N_10367,N_5402,N_7264);
nand U10368 (N_10368,N_5229,N_9955);
xnor U10369 (N_10369,N_8921,N_6420);
or U10370 (N_10370,N_7642,N_5777);
or U10371 (N_10371,N_6892,N_6250);
nor U10372 (N_10372,N_6780,N_8635);
or U10373 (N_10373,N_9059,N_8935);
nand U10374 (N_10374,N_6514,N_9037);
nand U10375 (N_10375,N_9583,N_8793);
nand U10376 (N_10376,N_5990,N_7130);
nor U10377 (N_10377,N_5003,N_8602);
or U10378 (N_10378,N_9815,N_6506);
and U10379 (N_10379,N_7042,N_8089);
nand U10380 (N_10380,N_5363,N_6087);
and U10381 (N_10381,N_8899,N_8957);
nor U10382 (N_10382,N_8586,N_6888);
and U10383 (N_10383,N_7046,N_7889);
nor U10384 (N_10384,N_7436,N_9989);
nor U10385 (N_10385,N_6226,N_6943);
and U10386 (N_10386,N_9248,N_7815);
nand U10387 (N_10387,N_9161,N_7273);
or U10388 (N_10388,N_9658,N_6808);
and U10389 (N_10389,N_7987,N_5272);
nor U10390 (N_10390,N_8325,N_7837);
nor U10391 (N_10391,N_6411,N_6263);
and U10392 (N_10392,N_9475,N_6283);
nor U10393 (N_10393,N_6336,N_7066);
xnor U10394 (N_10394,N_6293,N_5063);
or U10395 (N_10395,N_5761,N_5503);
nand U10396 (N_10396,N_7940,N_5984);
or U10397 (N_10397,N_5043,N_6669);
or U10398 (N_10398,N_6445,N_9881);
nand U10399 (N_10399,N_5291,N_7780);
xnor U10400 (N_10400,N_7955,N_6987);
or U10401 (N_10401,N_8007,N_9917);
nand U10402 (N_10402,N_8241,N_5112);
xnor U10403 (N_10403,N_8301,N_5303);
and U10404 (N_10404,N_7592,N_9384);
and U10405 (N_10405,N_8593,N_5283);
nand U10406 (N_10406,N_9337,N_8109);
or U10407 (N_10407,N_8830,N_9585);
or U10408 (N_10408,N_6351,N_6017);
nor U10409 (N_10409,N_6449,N_6310);
or U10410 (N_10410,N_5392,N_9312);
or U10411 (N_10411,N_8508,N_7054);
and U10412 (N_10412,N_9284,N_8004);
nor U10413 (N_10413,N_9182,N_5473);
nor U10414 (N_10414,N_6244,N_9121);
nor U10415 (N_10415,N_5008,N_8310);
and U10416 (N_10416,N_9040,N_9473);
nor U10417 (N_10417,N_6848,N_6789);
nor U10418 (N_10418,N_9998,N_8377);
nor U10419 (N_10419,N_8923,N_7284);
nand U10420 (N_10420,N_7983,N_9592);
and U10421 (N_10421,N_9138,N_6018);
nor U10422 (N_10422,N_9393,N_5231);
and U10423 (N_10423,N_6366,N_8146);
or U10424 (N_10424,N_7487,N_5528);
xor U10425 (N_10425,N_8582,N_7666);
nand U10426 (N_10426,N_5904,N_8903);
or U10427 (N_10427,N_5105,N_5840);
nand U10428 (N_10428,N_9838,N_7458);
nor U10429 (N_10429,N_8167,N_8344);
and U10430 (N_10430,N_5541,N_8006);
or U10431 (N_10431,N_5094,N_7034);
nor U10432 (N_10432,N_9952,N_6214);
nor U10433 (N_10433,N_5522,N_6076);
nor U10434 (N_10434,N_5041,N_9043);
and U10435 (N_10435,N_7986,N_5312);
or U10436 (N_10436,N_6962,N_7910);
and U10437 (N_10437,N_8698,N_7834);
nor U10438 (N_10438,N_7445,N_6713);
nand U10439 (N_10439,N_5434,N_6077);
nand U10440 (N_10440,N_9385,N_6147);
nand U10441 (N_10441,N_8730,N_7801);
nor U10442 (N_10442,N_6080,N_5920);
or U10443 (N_10443,N_8787,N_5050);
or U10444 (N_10444,N_6699,N_9260);
nor U10445 (N_10445,N_9546,N_7628);
and U10446 (N_10446,N_6075,N_5131);
nand U10447 (N_10447,N_6527,N_8423);
nor U10448 (N_10448,N_5605,N_7616);
or U10449 (N_10449,N_9424,N_8776);
nor U10450 (N_10450,N_5833,N_7015);
nand U10451 (N_10451,N_7635,N_9159);
and U10452 (N_10452,N_9935,N_6860);
or U10453 (N_10453,N_5658,N_5930);
or U10454 (N_10454,N_7512,N_7334);
nor U10455 (N_10455,N_8129,N_9185);
or U10456 (N_10456,N_7071,N_5000);
and U10457 (N_10457,N_9347,N_9742);
and U10458 (N_10458,N_8836,N_6031);
nor U10459 (N_10459,N_8880,N_8594);
and U10460 (N_10460,N_6435,N_6308);
and U10461 (N_10461,N_8166,N_9982);
nand U10462 (N_10462,N_9395,N_6865);
nand U10463 (N_10463,N_9871,N_9883);
and U10464 (N_10464,N_6436,N_9400);
and U10465 (N_10465,N_7032,N_5096);
and U10466 (N_10466,N_7391,N_6701);
nand U10467 (N_10467,N_9375,N_9506);
nand U10468 (N_10468,N_6054,N_8376);
nand U10469 (N_10469,N_9243,N_6377);
and U10470 (N_10470,N_8227,N_5489);
or U10471 (N_10471,N_7809,N_7760);
nand U10472 (N_10472,N_8571,N_6567);
nor U10473 (N_10473,N_8224,N_6194);
and U10474 (N_10474,N_7771,N_7994);
and U10475 (N_10475,N_6316,N_5118);
nand U10476 (N_10476,N_6296,N_9788);
and U10477 (N_10477,N_7946,N_9977);
nor U10478 (N_10478,N_7453,N_8700);
or U10479 (N_10479,N_8210,N_6834);
or U10480 (N_10480,N_8761,N_7085);
and U10481 (N_10481,N_6417,N_8306);
nand U10482 (N_10482,N_5933,N_7493);
nand U10483 (N_10483,N_8800,N_5729);
nor U10484 (N_10484,N_6406,N_6422);
or U10485 (N_10485,N_5326,N_8712);
or U10486 (N_10486,N_9983,N_7660);
or U10487 (N_10487,N_5823,N_7559);
nand U10488 (N_10488,N_6231,N_6674);
xnor U10489 (N_10489,N_7918,N_7477);
and U10490 (N_10490,N_7371,N_9822);
and U10491 (N_10491,N_6564,N_9468);
nand U10492 (N_10492,N_6794,N_5670);
and U10493 (N_10493,N_6661,N_9941);
nor U10494 (N_10494,N_9352,N_9669);
nand U10495 (N_10495,N_8856,N_5638);
nand U10496 (N_10496,N_5398,N_7909);
nand U10497 (N_10497,N_8013,N_7142);
nand U10498 (N_10498,N_6198,N_7981);
nand U10499 (N_10499,N_8936,N_9591);
nor U10500 (N_10500,N_5164,N_5054);
nor U10501 (N_10501,N_8413,N_5333);
nor U10502 (N_10502,N_9076,N_6957);
nor U10503 (N_10503,N_9338,N_7805);
and U10504 (N_10504,N_6991,N_9900);
nor U10505 (N_10505,N_8435,N_6968);
nor U10506 (N_10506,N_7524,N_5592);
nor U10507 (N_10507,N_9302,N_9089);
and U10508 (N_10508,N_5292,N_5200);
nor U10509 (N_10509,N_8536,N_5537);
nand U10510 (N_10510,N_6222,N_7644);
xor U10511 (N_10511,N_7268,N_7870);
nor U10512 (N_10512,N_5019,N_7736);
or U10513 (N_10513,N_9787,N_5174);
and U10514 (N_10514,N_8211,N_9252);
nand U10515 (N_10515,N_6235,N_6887);
nand U10516 (N_10516,N_6209,N_9274);
nand U10517 (N_10517,N_7826,N_5913);
nor U10518 (N_10518,N_8546,N_5066);
or U10519 (N_10519,N_6635,N_8317);
nor U10520 (N_10520,N_7216,N_7122);
nor U10521 (N_10521,N_7043,N_5957);
nor U10522 (N_10522,N_6257,N_5797);
and U10523 (N_10523,N_9623,N_7366);
and U10524 (N_10524,N_6981,N_5240);
and U10525 (N_10525,N_6856,N_6480);
or U10526 (N_10526,N_7120,N_8600);
nand U10527 (N_10527,N_8952,N_8419);
and U10528 (N_10528,N_9867,N_6565);
and U10529 (N_10529,N_7447,N_6684);
or U10530 (N_10530,N_7556,N_8485);
and U10531 (N_10531,N_5871,N_7516);
or U10532 (N_10532,N_8946,N_8439);
and U10533 (N_10533,N_8891,N_9379);
and U10534 (N_10534,N_7428,N_8537);
and U10535 (N_10535,N_9873,N_8967);
and U10536 (N_10536,N_6557,N_8585);
or U10537 (N_10537,N_8040,N_6550);
and U10538 (N_10538,N_9652,N_7717);
nor U10539 (N_10539,N_7586,N_5470);
or U10540 (N_10540,N_6773,N_8829);
or U10541 (N_10541,N_5456,N_7846);
or U10542 (N_10542,N_6040,N_9034);
nand U10543 (N_10543,N_7265,N_9418);
nand U10544 (N_10544,N_8202,N_9693);
nor U10545 (N_10545,N_8239,N_8502);
nor U10546 (N_10546,N_7288,N_9938);
nand U10547 (N_10547,N_6249,N_7884);
nand U10548 (N_10548,N_7171,N_8618);
nor U10549 (N_10549,N_9147,N_5757);
nor U10550 (N_10550,N_8190,N_9282);
and U10551 (N_10551,N_7369,N_8784);
nand U10552 (N_10552,N_8742,N_5374);
and U10553 (N_10553,N_9741,N_7878);
nor U10554 (N_10554,N_8193,N_8874);
and U10555 (N_10555,N_7482,N_9466);
or U10556 (N_10556,N_9754,N_5803);
and U10557 (N_10557,N_5531,N_6152);
nand U10558 (N_10558,N_7191,N_5588);
nand U10559 (N_10559,N_5280,N_5822);
and U10560 (N_10560,N_7857,N_7943);
nand U10561 (N_10561,N_8898,N_9709);
nor U10562 (N_10562,N_8242,N_8441);
and U10563 (N_10563,N_9639,N_9193);
nor U10564 (N_10564,N_9191,N_6424);
nand U10565 (N_10565,N_9918,N_6993);
or U10566 (N_10566,N_8869,N_9816);
nand U10567 (N_10567,N_7189,N_6929);
or U10568 (N_10568,N_9636,N_8755);
or U10569 (N_10569,N_5263,N_6650);
nand U10570 (N_10570,N_6485,N_6524);
and U10571 (N_10571,N_7929,N_8693);
nor U10572 (N_10572,N_9611,N_9256);
or U10573 (N_10573,N_5453,N_7160);
nor U10574 (N_10574,N_9025,N_6916);
or U10575 (N_10575,N_5318,N_8789);
and U10576 (N_10576,N_9171,N_7877);
nand U10577 (N_10577,N_7598,N_9009);
nor U10578 (N_10578,N_5864,N_6264);
nand U10579 (N_10579,N_9766,N_9664);
nand U10580 (N_10580,N_6913,N_7553);
nand U10581 (N_10581,N_7327,N_7093);
nor U10582 (N_10582,N_6985,N_6399);
nand U10583 (N_10583,N_7254,N_7704);
nand U10584 (N_10584,N_5005,N_9571);
and U10585 (N_10585,N_8992,N_9023);
nand U10586 (N_10586,N_9596,N_7276);
nor U10587 (N_10587,N_6960,N_5953);
or U10588 (N_10588,N_7619,N_9230);
nor U10589 (N_10589,N_7350,N_6438);
nand U10590 (N_10590,N_9861,N_6340);
and U10591 (N_10591,N_8752,N_6384);
and U10592 (N_10592,N_8955,N_6083);
nor U10593 (N_10593,N_9538,N_5715);
or U10594 (N_10594,N_8305,N_7689);
nor U10595 (N_10595,N_9855,N_7231);
nand U10596 (N_10596,N_6516,N_9663);
or U10597 (N_10597,N_5661,N_9719);
or U10598 (N_10598,N_7115,N_8556);
nand U10599 (N_10599,N_5136,N_7803);
or U10600 (N_10600,N_5633,N_6596);
nor U10601 (N_10601,N_7851,N_9728);
or U10602 (N_10602,N_9705,N_7608);
and U10603 (N_10603,N_5270,N_9607);
and U10604 (N_10604,N_6103,N_8288);
or U10605 (N_10605,N_6900,N_6403);
or U10606 (N_10606,N_6597,N_5878);
xor U10607 (N_10607,N_6431,N_6624);
xor U10608 (N_10608,N_7321,N_6279);
nand U10609 (N_10609,N_5030,N_9770);
or U10610 (N_10610,N_6429,N_9083);
nand U10611 (N_10611,N_7424,N_5073);
xnor U10612 (N_10612,N_7149,N_7058);
or U10613 (N_10613,N_7500,N_6786);
and U10614 (N_10614,N_6130,N_7699);
and U10615 (N_10615,N_9661,N_9942);
nor U10616 (N_10616,N_8251,N_9856);
and U10617 (N_10617,N_7169,N_7179);
and U10618 (N_10618,N_6110,N_6477);
and U10619 (N_10619,N_9155,N_9763);
or U10620 (N_10620,N_5147,N_7102);
and U10621 (N_10621,N_6005,N_8001);
and U10622 (N_10622,N_5007,N_9806);
xor U10623 (N_10623,N_9834,N_6394);
and U10624 (N_10624,N_5279,N_5477);
nand U10625 (N_10625,N_7995,N_6333);
nor U10626 (N_10626,N_6140,N_6367);
nand U10627 (N_10627,N_6414,N_7711);
nor U10628 (N_10628,N_9028,N_5461);
and U10629 (N_10629,N_8801,N_8529);
or U10630 (N_10630,N_6812,N_7491);
nand U10631 (N_10631,N_8970,N_9559);
nor U10632 (N_10632,N_8888,N_6421);
or U10633 (N_10633,N_9819,N_5278);
nor U10634 (N_10634,N_7494,N_9474);
nor U10635 (N_10635,N_9102,N_6292);
and U10636 (N_10636,N_9190,N_8771);
and U10637 (N_10637,N_9968,N_9281);
and U10638 (N_10638,N_6656,N_7923);
nor U10639 (N_10639,N_6767,N_9866);
and U10640 (N_10640,N_6893,N_6711);
nor U10641 (N_10641,N_7655,N_7197);
nand U10642 (N_10642,N_9860,N_5304);
nor U10643 (N_10643,N_8631,N_5345);
nand U10644 (N_10644,N_5412,N_7903);
or U10645 (N_10645,N_9704,N_6248);
or U10646 (N_10646,N_5836,N_5273);
or U10647 (N_10647,N_5917,N_8831);
nand U10648 (N_10648,N_6282,N_6496);
nand U10649 (N_10649,N_9810,N_5639);
nand U10650 (N_10650,N_5615,N_5702);
nor U10651 (N_10651,N_8408,N_7033);
nand U10652 (N_10652,N_7778,N_8112);
nand U10653 (N_10653,N_6033,N_7021);
and U10654 (N_10654,N_6804,N_7407);
nand U10655 (N_10655,N_9378,N_8884);
nor U10656 (N_10656,N_7091,N_5350);
nand U10657 (N_10657,N_6079,N_8311);
and U10658 (N_10658,N_6158,N_8358);
nor U10659 (N_10659,N_5691,N_6725);
or U10660 (N_10660,N_5462,N_5571);
nand U10661 (N_10661,N_8701,N_8517);
nand U10662 (N_10662,N_6693,N_7035);
nand U10663 (N_10663,N_5533,N_8018);
and U10664 (N_10664,N_7464,N_8382);
nand U10665 (N_10665,N_5698,N_9510);
and U10666 (N_10666,N_5296,N_6645);
nand U10667 (N_10667,N_6680,N_6630);
or U10668 (N_10668,N_7223,N_7098);
nand U10669 (N_10669,N_8280,N_8750);
nor U10670 (N_10670,N_9053,N_9752);
or U10671 (N_10671,N_9253,N_5535);
xor U10672 (N_10672,N_6819,N_9210);
nand U10673 (N_10673,N_6905,N_6177);
and U10674 (N_10674,N_8472,N_6895);
or U10675 (N_10675,N_6455,N_7722);
nor U10676 (N_10676,N_5510,N_7310);
and U10677 (N_10677,N_8182,N_7745);
nand U10678 (N_10678,N_9603,N_7092);
or U10679 (N_10679,N_6732,N_5628);
and U10680 (N_10680,N_7335,N_9540);
nor U10681 (N_10681,N_7762,N_8879);
nand U10682 (N_10682,N_8454,N_8578);
and U10683 (N_10683,N_9203,N_9033);
nand U10684 (N_10684,N_5625,N_8969);
nand U10685 (N_10685,N_6067,N_7075);
nand U10686 (N_10686,N_7282,N_9826);
nor U10687 (N_10687,N_8120,N_9973);
nor U10688 (N_10688,N_7031,N_5667);
or U10689 (N_10689,N_9630,N_6500);
or U10690 (N_10690,N_6331,N_5425);
nand U10691 (N_10691,N_6548,N_5719);
or U10692 (N_10692,N_5201,N_9051);
nor U10693 (N_10693,N_8663,N_6863);
or U10694 (N_10694,N_6495,N_5655);
or U10695 (N_10695,N_8675,N_7654);
and U10696 (N_10696,N_9392,N_5606);
nand U10697 (N_10697,N_9824,N_5420);
or U10698 (N_10698,N_9561,N_6096);
and U10699 (N_10699,N_9245,N_8940);
nor U10700 (N_10700,N_8872,N_8262);
and U10701 (N_10701,N_6433,N_5950);
and U10702 (N_10702,N_5561,N_8838);
nand U10703 (N_10703,N_8959,N_9802);
nand U10704 (N_10704,N_8293,N_5602);
and U10705 (N_10705,N_5460,N_6499);
or U10706 (N_10706,N_9434,N_7721);
or U10707 (N_10707,N_6413,N_9620);
and U10708 (N_10708,N_8729,N_6679);
or U10709 (N_10709,N_6196,N_9492);
xnor U10710 (N_10710,N_6136,N_8387);
nand U10711 (N_10711,N_5978,N_9188);
nand U10712 (N_10712,N_7383,N_5743);
and U10713 (N_10713,N_6829,N_8859);
nor U10714 (N_10714,N_9481,N_7220);
nand U10715 (N_10715,N_7425,N_6275);
nor U10716 (N_10716,N_6979,N_8558);
nor U10717 (N_10717,N_6397,N_7212);
xnor U10718 (N_10718,N_6783,N_9545);
nor U10719 (N_10719,N_6769,N_7627);
and U10720 (N_10720,N_6474,N_8848);
and U10721 (N_10721,N_8632,N_5652);
and U10722 (N_10722,N_8749,N_8725);
nand U10723 (N_10723,N_8674,N_7455);
nand U10724 (N_10724,N_8853,N_9683);
or U10725 (N_10725,N_5171,N_5741);
nor U10726 (N_10726,N_5262,N_6070);
nand U10727 (N_10727,N_8025,N_7591);
or U10728 (N_10728,N_6391,N_8650);
and U10729 (N_10729,N_7700,N_6148);
nor U10730 (N_10730,N_9421,N_7481);
nor U10731 (N_10731,N_8488,N_5474);
nand U10732 (N_10732,N_8279,N_6059);
xor U10733 (N_10733,N_8255,N_8551);
and U10734 (N_10734,N_8860,N_5894);
or U10735 (N_10735,N_8524,N_8892);
nand U10736 (N_10736,N_6685,N_5689);
nand U10737 (N_10737,N_7633,N_7920);
and U10738 (N_10738,N_8799,N_8575);
nand U10739 (N_10739,N_9776,N_7448);
nand U10740 (N_10740,N_8989,N_5190);
nand U10741 (N_10741,N_9613,N_9813);
nand U10742 (N_10742,N_9262,N_7419);
or U10743 (N_10743,N_6488,N_6188);
xor U10744 (N_10744,N_5540,N_7045);
or U10745 (N_10745,N_8047,N_6089);
nand U10746 (N_10746,N_8964,N_9647);
nand U10747 (N_10747,N_7939,N_9444);
nor U10748 (N_10748,N_6750,N_7077);
nor U10749 (N_10749,N_8291,N_9577);
and U10750 (N_10750,N_7588,N_6967);
or U10751 (N_10751,N_5172,N_6217);
and U10752 (N_10752,N_6736,N_6705);
xor U10753 (N_10753,N_5820,N_9030);
xnor U10754 (N_10754,N_9163,N_8221);
and U10755 (N_10755,N_5196,N_8583);
or U10756 (N_10756,N_9563,N_9924);
nor U10757 (N_10757,N_7899,N_5384);
nor U10758 (N_10758,N_9298,N_7200);
nor U10759 (N_10759,N_9366,N_9213);
or U10760 (N_10760,N_7330,N_6655);
nor U10761 (N_10761,N_9239,N_7174);
xor U10762 (N_10762,N_9362,N_9753);
or U10763 (N_10763,N_9004,N_5455);
nor U10764 (N_10764,N_5587,N_6584);
and U10765 (N_10765,N_9678,N_7858);
or U10766 (N_10766,N_5065,N_9780);
or U10767 (N_10767,N_7542,N_9990);
nor U10768 (N_10768,N_5839,N_7687);
nand U10769 (N_10769,N_6207,N_8401);
nand U10770 (N_10770,N_8128,N_6060);
nand U10771 (N_10771,N_5093,N_5583);
or U10772 (N_10772,N_9014,N_6874);
nor U10773 (N_10773,N_7651,N_6798);
and U10774 (N_10774,N_9277,N_9594);
or U10775 (N_10775,N_7763,N_5976);
or U10776 (N_10776,N_8243,N_7682);
and U10777 (N_10777,N_5339,N_5724);
or U10778 (N_10778,N_9721,N_7207);
and U10779 (N_10779,N_7752,N_9588);
nor U10780 (N_10780,N_9953,N_9828);
or U10781 (N_10781,N_5879,N_5676);
nor U10782 (N_10782,N_6082,N_7400);
nand U10783 (N_10783,N_7397,N_8220);
or U10784 (N_10784,N_8099,N_8851);
nor U10785 (N_10785,N_5750,N_8084);
nor U10786 (N_10786,N_6210,N_8824);
nand U10787 (N_10787,N_6692,N_9280);
nor U10788 (N_10788,N_7818,N_6821);
nand U10789 (N_10789,N_6350,N_6619);
and U10790 (N_10790,N_5194,N_8999);
nand U10791 (N_10791,N_6742,N_6509);
and U10792 (N_10792,N_8039,N_8133);
nand U10793 (N_10793,N_7213,N_7005);
nor U10794 (N_10794,N_5221,N_8181);
nor U10795 (N_10795,N_8158,N_7847);
or U10796 (N_10796,N_9365,N_7526);
nor U10797 (N_10797,N_7649,N_9237);
nor U10798 (N_10798,N_7845,N_5934);
and U10799 (N_10799,N_9293,N_6579);
or U10800 (N_10800,N_8231,N_8850);
nor U10801 (N_10801,N_6016,N_5575);
nand U10802 (N_10802,N_9695,N_8337);
nand U10803 (N_10803,N_9648,N_6458);
and U10804 (N_10804,N_5708,N_9617);
and U10805 (N_10805,N_7758,N_8038);
nand U10806 (N_10806,N_8503,N_8391);
or U10807 (N_10807,N_9685,N_7724);
nor U10808 (N_10808,N_7414,N_9862);
and U10809 (N_10809,N_5366,N_6415);
and U10810 (N_10810,N_8626,N_9287);
xor U10811 (N_10811,N_5154,N_8493);
and U10812 (N_10812,N_7090,N_7109);
nor U10813 (N_10813,N_6300,N_6795);
nor U10814 (N_10814,N_8939,N_7232);
nor U10815 (N_10815,N_9804,N_6702);
and U10816 (N_10816,N_8240,N_8277);
or U10817 (N_10817,N_6364,N_6562);
or U10818 (N_10818,N_8720,N_8442);
nand U10819 (N_10819,N_7600,N_6386);
nor U10820 (N_10820,N_8415,N_6191);
or U10821 (N_10821,N_5214,N_7963);
and U10822 (N_10822,N_8792,N_5543);
or U10823 (N_10823,N_6050,N_5909);
or U10824 (N_10824,N_6602,N_7835);
or U10825 (N_10825,N_8913,N_5612);
and U10826 (N_10826,N_9141,N_5259);
and U10827 (N_10827,N_9386,N_5791);
or U10828 (N_10828,N_8533,N_5785);
and U10829 (N_10829,N_6587,N_9522);
and U10830 (N_10830,N_8154,N_8796);
and U10831 (N_10831,N_6637,N_8828);
and U10832 (N_10832,N_6825,N_7716);
or U10833 (N_10833,N_5872,N_6276);
nand U10834 (N_10834,N_6833,N_6928);
nor U10835 (N_10835,N_7541,N_5097);
nor U10836 (N_10836,N_7697,N_6094);
nor U10837 (N_10837,N_6503,N_5875);
nor U10838 (N_10838,N_8212,N_9641);
nand U10839 (N_10839,N_8573,N_7962);
nor U10840 (N_10840,N_5900,N_7656);
nor U10841 (N_10841,N_5012,N_9928);
xnor U10842 (N_10842,N_8522,N_9258);
or U10843 (N_10843,N_8766,N_5016);
and U10844 (N_10844,N_7537,N_8846);
nor U10845 (N_10845,N_9301,N_6746);
and U10846 (N_10846,N_7703,N_8136);
and U10847 (N_10847,N_8991,N_9414);
or U10848 (N_10848,N_9894,N_6126);
nor U10849 (N_10849,N_8802,N_5673);
and U10850 (N_10850,N_6437,N_9082);
nand U10851 (N_10851,N_7444,N_6463);
and U10852 (N_10852,N_5082,N_7079);
nand U10853 (N_10853,N_6376,N_9638);
nor U10854 (N_10854,N_9503,N_8844);
nand U10855 (N_10855,N_8092,N_9622);
or U10856 (N_10856,N_7796,N_7006);
and U10857 (N_10857,N_9307,N_5664);
nand U10858 (N_10858,N_9368,N_6781);
nor U10859 (N_10859,N_6446,N_5952);
and U10860 (N_10860,N_6036,N_5241);
xnor U10861 (N_10861,N_7748,N_8947);
nand U10862 (N_10862,N_5167,N_8150);
or U10863 (N_10863,N_8688,N_6013);
or U10864 (N_10864,N_6729,N_7309);
and U10865 (N_10865,N_6508,N_8214);
nand U10866 (N_10866,N_5569,N_8169);
and U10867 (N_10867,N_7121,N_7287);
nand U10868 (N_10868,N_5083,N_5307);
nand U10869 (N_10869,N_8307,N_8468);
or U10870 (N_10870,N_5965,N_6113);
or U10871 (N_10871,N_8961,N_5947);
or U10872 (N_10872,N_7315,N_6592);
nor U10873 (N_10873,N_7233,N_8498);
and U10874 (N_10874,N_6473,N_6984);
nor U10875 (N_10875,N_7905,N_6097);
nand U10876 (N_10876,N_8807,N_8806);
nor U10877 (N_10877,N_8757,N_5124);
nand U10878 (N_10878,N_6419,N_7128);
or U10879 (N_10879,N_6277,N_9269);
nand U10880 (N_10880,N_7839,N_9422);
or U10881 (N_10881,N_9323,N_9864);
and U10882 (N_10882,N_6618,N_5331);
or U10883 (N_10883,N_9220,N_8887);
and U10884 (N_10884,N_8417,N_7381);
or U10885 (N_10885,N_9505,N_9714);
and U10886 (N_10886,N_9325,N_8610);
or U10887 (N_10887,N_7535,N_9095);
nor U10888 (N_10888,N_7560,N_8564);
and U10889 (N_10889,N_5529,N_5029);
nand U10890 (N_10890,N_9616,N_8737);
nand U10891 (N_10891,N_8282,N_5939);
or U10892 (N_10892,N_7916,N_9995);
nand U10893 (N_10893,N_5415,N_6926);
or U10894 (N_10894,N_6327,N_6444);
nor U10895 (N_10895,N_8185,N_6038);
nand U10896 (N_10896,N_9205,N_7741);
and U10897 (N_10897,N_8303,N_9633);
nand U10898 (N_10898,N_9232,N_9129);
or U10899 (N_10899,N_6073,N_9764);
or U10900 (N_10900,N_9509,N_7816);
nand U10901 (N_10901,N_6832,N_5509);
nor U10902 (N_10902,N_8951,N_6305);
nand U10903 (N_10903,N_6574,N_5787);
nor U10904 (N_10904,N_5520,N_6163);
and U10905 (N_10905,N_5993,N_8300);
nor U10906 (N_10906,N_6258,N_6032);
or U10907 (N_10907,N_9132,N_6375);
or U10908 (N_10908,N_7040,N_7671);
nand U10909 (N_10909,N_8444,N_7615);
or U10910 (N_10910,N_6121,N_9461);
or U10911 (N_10911,N_8950,N_8562);
nor U10912 (N_10912,N_8907,N_9438);
nand U10913 (N_10913,N_8769,N_8671);
or U10914 (N_10914,N_9814,N_8706);
and U10915 (N_10915,N_6749,N_9738);
nor U10916 (N_10916,N_7384,N_9118);
and U10917 (N_10917,N_9646,N_5627);
or U10918 (N_10918,N_6726,N_8681);
or U10919 (N_10919,N_9212,N_9332);
nor U10920 (N_10920,N_5260,N_6467);
and U10921 (N_10921,N_6269,N_8061);
nand U10922 (N_10922,N_9451,N_7930);
or U10923 (N_10923,N_6011,N_5809);
and U10924 (N_10924,N_8137,N_9169);
or U10925 (N_10925,N_7570,N_5927);
or U10926 (N_10926,N_8637,N_6775);
and U10927 (N_10927,N_7263,N_9701);
or U10928 (N_10928,N_9125,N_7272);
nand U10929 (N_10929,N_7379,N_9922);
and U10930 (N_10930,N_7036,N_9783);
nand U10931 (N_10931,N_8478,N_6199);
nor U10932 (N_10932,N_7504,N_5256);
xnor U10933 (N_10933,N_6510,N_7367);
or U10934 (N_10934,N_9809,N_6329);
and U10935 (N_10935,N_8855,N_8123);
nor U10936 (N_10936,N_5863,N_6814);
and U10937 (N_10937,N_7417,N_8079);
nor U10938 (N_10938,N_8051,N_7973);
and U10939 (N_10939,N_6370,N_6313);
and U10940 (N_10940,N_7406,N_6062);
or U10941 (N_10941,N_7785,N_7457);
or U10942 (N_10942,N_6183,N_5045);
or U10943 (N_10943,N_9877,N_7168);
nor U10944 (N_10944,N_7485,N_5701);
nand U10945 (N_10945,N_9609,N_7190);
or U10946 (N_10946,N_7505,N_7552);
and U10947 (N_10947,N_7301,N_6690);
or U10948 (N_10948,N_7880,N_7951);
nor U10949 (N_10949,N_5653,N_5620);
or U10950 (N_10950,N_6314,N_9673);
or U10951 (N_10951,N_5498,N_5772);
or U10952 (N_10952,N_9099,N_5383);
and U10953 (N_10953,N_6362,N_9158);
or U10954 (N_10954,N_8786,N_8196);
and U10955 (N_10955,N_6291,N_9087);
nand U10956 (N_10956,N_7513,N_7473);
and U10957 (N_10957,N_8858,N_6838);
nor U10958 (N_10958,N_6747,N_8434);
or U10959 (N_10959,N_5250,N_5417);
nor U10960 (N_10960,N_8825,N_5690);
or U10961 (N_10961,N_9808,N_5183);
nor U10962 (N_10962,N_6439,N_8031);
nor U10963 (N_10963,N_6844,N_8226);
or U10964 (N_10964,N_7675,N_5141);
and U10965 (N_10965,N_9305,N_7938);
nand U10966 (N_10966,N_9175,N_9391);
and U10967 (N_10967,N_6740,N_5254);
nor U10968 (N_10968,N_5433,N_5746);
or U10969 (N_10969,N_5022,N_9453);
or U10970 (N_10970,N_5157,N_6764);
and U10971 (N_10971,N_7250,N_9837);
nand U10972 (N_10972,N_9353,N_5554);
nand U10973 (N_10973,N_6664,N_5393);
or U10974 (N_10974,N_8795,N_8958);
and U10975 (N_10975,N_8719,N_8278);
and U10976 (N_10976,N_8711,N_9425);
or U10977 (N_10977,N_8612,N_5160);
and U10978 (N_10978,N_9778,N_6205);
and U10979 (N_10979,N_6846,N_5792);
or U10980 (N_10980,N_6379,N_5829);
nor U10981 (N_10981,N_6776,N_7317);
or U10982 (N_10982,N_6796,N_8591);
or U10983 (N_10983,N_8427,N_5107);
or U10984 (N_10984,N_6243,N_6135);
and U10985 (N_10985,N_6658,N_9318);
or U10986 (N_10986,N_6156,N_6741);
nor U10987 (N_10987,N_9666,N_6830);
or U10988 (N_10988,N_6008,N_5432);
nor U10989 (N_10989,N_6015,N_9130);
or U10990 (N_10990,N_6517,N_8805);
and U10991 (N_10991,N_7612,N_6167);
and U10992 (N_10992,N_6108,N_7543);
and U10993 (N_10993,N_8963,N_9978);
nand U10994 (N_10994,N_5405,N_5075);
nor U10995 (N_10995,N_7713,N_8289);
and U10996 (N_10996,N_8922,N_8354);
and U10997 (N_10997,N_7498,N_7235);
xnor U10998 (N_10998,N_7779,N_9708);
nand U10999 (N_10999,N_9850,N_7611);
nor U11000 (N_11000,N_7267,N_9945);
or U11001 (N_11001,N_7456,N_6380);
or U11002 (N_11002,N_9552,N_9218);
nand U11003 (N_11003,N_6470,N_9904);
or U11004 (N_11004,N_8342,N_7789);
nand U11005 (N_11005,N_7337,N_6884);
nand U11006 (N_11006,N_7411,N_8545);
nand U11007 (N_11007,N_7433,N_8995);
and U11008 (N_11008,N_5357,N_5032);
nor U11009 (N_11009,N_8822,N_5400);
nand U11010 (N_11010,N_7359,N_9062);
nor U11011 (N_11011,N_8876,N_9751);
and U11012 (N_11012,N_7132,N_9231);
nor U11013 (N_11013,N_8285,N_6552);
nor U11014 (N_11014,N_8535,N_7057);
nor U11015 (N_11015,N_8385,N_7324);
or U11016 (N_11016,N_7480,N_5129);
or U11017 (N_11017,N_7777,N_7587);
nor U11018 (N_11018,N_6064,N_9303);
nor U11019 (N_11019,N_7055,N_8206);
nor U11020 (N_11020,N_8849,N_7810);
and U11021 (N_11021,N_5828,N_5884);
nor U11022 (N_11022,N_6784,N_5418);
or U11023 (N_11023,N_7813,N_5549);
and U11024 (N_11024,N_7709,N_5513);
nand U11025 (N_11025,N_9279,N_9735);
and U11026 (N_11026,N_9437,N_5662);
nand U11027 (N_11027,N_8331,N_8499);
or U11028 (N_11028,N_5300,N_8067);
or U11029 (N_11029,N_6387,N_6569);
nor U11030 (N_11030,N_6807,N_6986);
nor U11031 (N_11031,N_5666,N_8024);
and U11032 (N_11032,N_5475,N_6529);
xor U11033 (N_11033,N_5062,N_6585);
nor U11034 (N_11034,N_5120,N_6737);
nor U11035 (N_11035,N_5494,N_6487);
and U11036 (N_11036,N_9536,N_6654);
or U11037 (N_11037,N_6165,N_9569);
nor U11038 (N_11038,N_7306,N_7915);
or U11039 (N_11039,N_6941,N_7532);
or U11040 (N_11040,N_7214,N_9164);
nor U11041 (N_11041,N_5598,N_9372);
or U11042 (N_11042,N_9275,N_7224);
nor U11043 (N_11043,N_9901,N_7467);
nor U11044 (N_11044,N_5322,N_5782);
nor U11045 (N_11045,N_7861,N_6708);
nand U11046 (N_11046,N_8445,N_5416);
nor U11047 (N_11047,N_9488,N_7097);
and U11048 (N_11048,N_9799,N_6836);
nand U11049 (N_11049,N_8679,N_8371);
nand U11050 (N_11050,N_7865,N_8560);
nor U11051 (N_11051,N_7825,N_7278);
nor U11052 (N_11052,N_7502,N_9448);
nand U11053 (N_11053,N_6827,N_5072);
nand U11054 (N_11054,N_5113,N_7271);
nor U11055 (N_11055,N_7002,N_8143);
or U11056 (N_11056,N_9796,N_7470);
nor U11057 (N_11057,N_6869,N_8033);
nand U11058 (N_11058,N_8443,N_7427);
and U11059 (N_11059,N_9612,N_6373);
or U11060 (N_11060,N_9360,N_5034);
or U11061 (N_11061,N_6770,N_6427);
nor U11062 (N_11062,N_6910,N_9972);
nand U11063 (N_11063,N_8928,N_5842);
nand U11064 (N_11064,N_6102,N_9747);
nor U11065 (N_11065,N_9667,N_5087);
nand U11066 (N_11066,N_7774,N_8017);
nand U11067 (N_11067,N_6123,N_9593);
and U11068 (N_11068,N_6259,N_7409);
and U11069 (N_11069,N_9905,N_8997);
or U11070 (N_11070,N_5565,N_6320);
nor U11071 (N_11071,N_9640,N_8321);
nor U11072 (N_11072,N_8177,N_8680);
and U11073 (N_11073,N_9949,N_5817);
nand U11074 (N_11074,N_8057,N_7582);
or U11075 (N_11075,N_8446,N_7087);
or U11076 (N_11076,N_8432,N_8058);
or U11077 (N_11077,N_8816,N_7368);
or U11078 (N_11078,N_7730,N_6657);
nand U11079 (N_11079,N_9156,N_8539);
or U11080 (N_11080,N_7180,N_8438);
nor U11081 (N_11081,N_6631,N_8094);
nor U11082 (N_11082,N_7253,N_5249);
nand U11083 (N_11083,N_9092,N_7868);
or U11084 (N_11084,N_6441,N_6533);
or U11085 (N_11085,N_8405,N_7775);
and U11086 (N_11086,N_7696,N_9523);
or U11087 (N_11087,N_9657,N_5914);
or U11088 (N_11088,N_9035,N_5137);
nor U11089 (N_11089,N_7921,N_9104);
and U11090 (N_11090,N_9296,N_9635);
xnor U11091 (N_11091,N_9749,N_9676);
nor U11092 (N_11092,N_5130,N_9097);
nand U11093 (N_11093,N_8471,N_9825);
nor U11094 (N_11094,N_5319,N_7283);
nand U11095 (N_11095,N_8324,N_6476);
nor U11096 (N_11096,N_7211,N_9061);
and U11097 (N_11097,N_5584,N_9225);
and U11098 (N_11098,N_7415,N_9330);
and U11099 (N_11099,N_7303,N_8821);
and U11100 (N_11100,N_5354,N_6026);
nor U11101 (N_11101,N_6883,N_6858);
or U11102 (N_11102,N_6721,N_8254);
and U11103 (N_11103,N_6176,N_5267);
or U11104 (N_11104,N_5430,N_9011);
or U11105 (N_11105,N_8703,N_9888);
nor U11106 (N_11106,N_6272,N_7050);
nor U11107 (N_11107,N_6047,N_7117);
and U11108 (N_11108,N_6144,N_6675);
or U11109 (N_11109,N_8739,N_8102);
nor U11110 (N_11110,N_6678,N_5958);
or U11111 (N_11111,N_8036,N_7037);
nor U11112 (N_11112,N_6395,N_5919);
or U11113 (N_11113,N_7201,N_8333);
nand U11114 (N_11114,N_5467,N_5156);
and U11115 (N_11115,N_9180,N_8895);
nand U11116 (N_11116,N_6914,N_8597);
nor U11117 (N_11117,N_8646,N_6639);
nor U11118 (N_11118,N_7137,N_6107);
nor U11119 (N_11119,N_5725,N_9207);
nor U11120 (N_11120,N_5923,N_7013);
nor U11121 (N_11121,N_9098,N_5982);
nor U11122 (N_11122,N_6453,N_6155);
and U11123 (N_11123,N_7118,N_8171);
nand U11124 (N_11124,N_9142,N_5538);
and U11125 (N_11125,N_9962,N_5732);
and U11126 (N_11126,N_5187,N_6505);
nor U11127 (N_11127,N_5501,N_5334);
or U11128 (N_11128,N_7984,N_9649);
and U11129 (N_11129,N_9456,N_6171);
nor U11130 (N_11130,N_8668,N_6989);
xor U11131 (N_11131,N_8754,N_6286);
and U11132 (N_11132,N_8809,N_6852);
or U11133 (N_11133,N_8421,N_5414);
or U11134 (N_11134,N_5271,N_7677);
nor U11135 (N_11135,N_8519,N_9729);
or U11136 (N_11136,N_9402,N_5786);
and U11137 (N_11137,N_8791,N_6744);
nor U11138 (N_11138,N_5867,N_6556);
and U11139 (N_11139,N_7313,N_9202);
and U11140 (N_11140,N_9580,N_8689);
and U11141 (N_11141,N_5011,N_9629);
nand U11142 (N_11142,N_8072,N_6586);
and U11143 (N_11143,N_7640,N_5117);
or U11144 (N_11144,N_7176,N_5372);
or U11145 (N_11145,N_6632,N_6182);
nor U11146 (N_11146,N_5980,N_5413);
nor U11147 (N_11147,N_9743,N_6344);
or U11148 (N_11148,N_7343,N_9173);
nor U11149 (N_11149,N_6933,N_5560);
nor U11150 (N_11150,N_9297,N_6288);
and U11151 (N_11151,N_5601,N_7864);
or U11152 (N_11152,N_6622,N_9511);
and U11153 (N_11153,N_7454,N_7398);
nor U11154 (N_11154,N_7738,N_5450);
nor U11155 (N_11155,N_5552,N_6211);
and U11156 (N_11156,N_8151,N_8122);
or U11157 (N_11157,N_8592,N_7246);
or U11158 (N_11158,N_8457,N_5579);
nor U11159 (N_11159,N_6202,N_8309);
nor U11160 (N_11160,N_8433,N_9584);
nor U11161 (N_11161,N_5110,N_9194);
or U11162 (N_11162,N_6688,N_7953);
and U11163 (N_11163,N_6240,N_9048);
and U11164 (N_11164,N_5895,N_8707);
and U11165 (N_11165,N_7038,N_6307);
and U11166 (N_11166,N_7725,N_5876);
or U11167 (N_11167,N_6695,N_7508);
or U11168 (N_11168,N_5145,N_6150);
and U11169 (N_11169,N_9339,N_5678);
nand U11170 (N_11170,N_7226,N_5426);
and U11171 (N_11171,N_6594,N_9820);
nor U11172 (N_11172,N_5440,N_8424);
nand U11173 (N_11173,N_9746,N_8684);
and U11174 (N_11174,N_5910,N_7141);
or U11175 (N_11175,N_5376,N_6137);
nor U11176 (N_11176,N_7010,N_9334);
nand U11177 (N_11177,N_8191,N_5362);
nand U11178 (N_11178,N_8032,N_7490);
nand U11179 (N_11179,N_6899,N_9800);
nand U11180 (N_11180,N_7051,N_5669);
nor U11181 (N_11181,N_9005,N_9899);
nand U11182 (N_11182,N_9272,N_5971);
and U11183 (N_11183,N_9249,N_9131);
or U11184 (N_11184,N_6220,N_7603);
or U11185 (N_11185,N_9777,N_7630);
nand U11186 (N_11186,N_5763,N_8156);
or U11187 (N_11187,N_5049,N_6227);
or U11188 (N_11188,N_5936,N_8496);
nand U11189 (N_11189,N_7465,N_7824);
or U11190 (N_11190,N_5586,N_5677);
nand U11191 (N_11191,N_7336,N_9976);
nand U11192 (N_11192,N_5395,N_5642);
nand U11193 (N_11193,N_7787,N_5946);
nor U11194 (N_11194,N_7893,N_9271);
nand U11195 (N_11195,N_5851,N_9668);
nor U11196 (N_11196,N_9936,N_8966);
or U11197 (N_11197,N_7746,N_6687);
nor U11198 (N_11198,N_5804,N_6159);
nand U11199 (N_11199,N_7449,N_9960);
nand U11200 (N_11200,N_9306,N_9206);
nand U11201 (N_11201,N_5176,N_9920);
nor U11202 (N_11202,N_7243,N_5811);
nand U11203 (N_11203,N_5865,N_8326);
or U11204 (N_11204,N_6216,N_9361);
nand U11205 (N_11205,N_9528,N_9299);
or U11206 (N_11206,N_8584,N_8839);
xnor U11207 (N_11207,N_5340,N_5807);
nor U11208 (N_11208,N_6751,N_6580);
nor U11209 (N_11209,N_5368,N_8975);
or U11210 (N_11210,N_7257,N_9712);
and U11211 (N_11211,N_9739,N_7164);
or U11212 (N_11212,N_5188,N_7561);
and U11213 (N_11213,N_7966,N_9550);
nor U11214 (N_11214,N_9032,N_9300);
xnor U11215 (N_11215,N_7061,N_9779);
or U11216 (N_11216,N_5955,N_5197);
nand U11217 (N_11217,N_7073,N_7665);
nand U11218 (N_11218,N_8469,N_7274);
and U11219 (N_11219,N_5539,N_6471);
nor U11220 (N_11220,N_5080,N_5281);
and U11221 (N_11221,N_8037,N_5944);
and U11222 (N_11222,N_9002,N_6698);
or U11223 (N_11223,N_6959,N_9390);
nand U11224 (N_11224,N_5313,N_8990);
nand U11225 (N_11225,N_6261,N_6409);
nand U11226 (N_11226,N_7358,N_6583);
and U11227 (N_11227,N_6234,N_6247);
nor U11228 (N_11228,N_6595,N_5518);
nand U11229 (N_11229,N_8201,N_6012);
and U11230 (N_11230,N_8511,N_8065);
or U11231 (N_11231,N_8842,N_8904);
or U11232 (N_11232,N_5422,N_9179);
or U11233 (N_11233,N_9154,N_6875);
and U11234 (N_11234,N_5966,N_5928);
nand U11235 (N_11235,N_6560,N_9500);
nor U11236 (N_11236,N_8993,N_5493);
or U11237 (N_11237,N_9458,N_6218);
or U11238 (N_11238,N_5935,N_8097);
or U11239 (N_11239,N_7363,N_5134);
or U11240 (N_11240,N_9333,N_8811);
and U11241 (N_11241,N_6052,N_5095);
nor U11242 (N_11242,N_5330,N_9435);
nand U11243 (N_11243,N_7242,N_6612);
and U11244 (N_11244,N_8819,N_9677);
nand U11245 (N_11245,N_6897,N_7989);
nor U11246 (N_11246,N_8657,N_5873);
or U11247 (N_11247,N_9412,N_6950);
and U11248 (N_11248,N_9292,N_6315);
xnor U11249 (N_11249,N_5680,N_6743);
nor U11250 (N_11250,N_6034,N_6390);
nand U11251 (N_11251,N_8568,N_9979);
and U11252 (N_11252,N_9520,N_6372);
nand U11253 (N_11253,N_6098,N_5580);
and U11254 (N_11254,N_7108,N_5115);
or U11255 (N_11255,N_5033,N_9166);
nand U11256 (N_11256,N_6189,N_8296);
or U11257 (N_11257,N_7203,N_7218);
nor U11258 (N_11258,N_5328,N_6304);
nor U11259 (N_11259,N_9113,N_5889);
nand U11260 (N_11260,N_7626,N_6911);
and U11261 (N_11261,N_6483,N_9408);
or U11262 (N_11262,N_5053,N_8271);
nor U11263 (N_11263,N_7866,N_6019);
nand U11264 (N_11264,N_9181,N_8581);
or U11265 (N_11265,N_5232,N_5317);
nand U11266 (N_11266,N_9058,N_8073);
nor U11267 (N_11267,N_8229,N_8713);
nand U11268 (N_11268,N_6145,N_7605);
nand U11269 (N_11269,N_7731,N_5675);
or U11270 (N_11270,N_7229,N_5466);
nand U11271 (N_11271,N_5512,N_9265);
or U11272 (N_11272,N_8000,N_6603);
nand U11273 (N_11273,N_5379,N_6638);
nand U11274 (N_11274,N_6649,N_8658);
nand U11275 (N_11275,N_6535,N_7739);
and U11276 (N_11276,N_7003,N_5776);
nor U11277 (N_11277,N_8124,N_5173);
and U11278 (N_11278,N_8183,N_5643);
and U11279 (N_11279,N_7147,N_5848);
or U11280 (N_11280,N_9507,N_9404);
and U11281 (N_11281,N_6570,N_5013);
nand U11282 (N_11282,N_5243,N_5862);
and U11283 (N_11283,N_6342,N_8138);
nand U11284 (N_11284,N_9836,N_7808);
or U11285 (N_11285,N_8518,N_5854);
nand U11286 (N_11286,N_7182,N_8818);
and U11287 (N_11287,N_5265,N_8702);
and U11288 (N_11288,N_5356,N_6854);
or U11289 (N_11289,N_9144,N_5151);
nand U11290 (N_11290,N_5515,N_9426);
nand U11291 (N_11291,N_6001,N_9148);
nor U11292 (N_11292,N_8389,N_6757);
or U11293 (N_11293,N_8845,N_6731);
and U11294 (N_11294,N_5555,N_6432);
nor U11295 (N_11295,N_9991,N_8386);
and U11296 (N_11296,N_6608,N_8576);
or U11297 (N_11297,N_5744,N_5428);
nand U11298 (N_11298,N_8449,N_5758);
nor U11299 (N_11299,N_9003,N_5490);
and U11300 (N_11300,N_5688,N_8238);
nor U11301 (N_11301,N_8753,N_5747);
and U11302 (N_11302,N_9499,N_5505);
and U11303 (N_11303,N_9316,N_9558);
and U11304 (N_11304,N_7804,N_9050);
or U11305 (N_11305,N_6229,N_7838);
nand U11306 (N_11306,N_9449,N_8651);
and U11307 (N_11307,N_5175,N_6694);
nand U11308 (N_11308,N_8565,N_6578);
or U11309 (N_11309,N_5610,N_5977);
or U11310 (N_11310,N_9263,N_9529);
nand U11311 (N_11311,N_6886,N_9184);
nand U11312 (N_11312,N_9268,N_9858);
nor U11313 (N_11313,N_7800,N_7429);
and U11314 (N_11314,N_7275,N_9396);
nand U11315 (N_11315,N_9653,N_8349);
nand U11316 (N_11316,N_7589,N_6132);
nor U11317 (N_11317,N_9963,N_7744);
nor U11318 (N_11318,N_5025,N_6319);
or U11319 (N_11319,N_6779,N_9913);
and U11320 (N_11320,N_5127,N_7533);
or U11321 (N_11321,N_7146,N_6238);
nand U11322 (N_11322,N_9351,N_9849);
or U11323 (N_11323,N_8082,N_7581);
nand U11324 (N_11324,N_6866,N_8740);
nand U11325 (N_11325,N_7860,N_5969);
and U11326 (N_11326,N_8590,N_8798);
nor U11327 (N_11327,N_5517,N_5389);
nand U11328 (N_11328,N_5573,N_9525);
and U11329 (N_11329,N_6072,N_9572);
nand U11330 (N_11330,N_6686,N_5888);
nor U11331 (N_11331,N_8284,N_6734);
nor U11332 (N_11332,N_7131,N_7869);
or U11333 (N_11333,N_9736,N_6454);
or U11334 (N_11334,N_7924,N_6146);
xor U11335 (N_11335,N_5940,N_8213);
or U11336 (N_11336,N_8267,N_6700);
and U11337 (N_11337,N_8944,N_7511);
or U11338 (N_11338,N_7679,N_5814);
or U11339 (N_11339,N_7806,N_9645);
nor U11340 (N_11340,N_5500,N_6507);
nand U11341 (N_11341,N_8738,N_5448);
or U11342 (N_11342,N_8292,N_6324);
and U11343 (N_11343,N_7821,N_8355);
nor U11344 (N_11344,N_5616,N_9687);
nor U11345 (N_11345,N_8782,N_9937);
and U11346 (N_11346,N_5244,N_8035);
nand U11347 (N_11347,N_9413,N_6803);
and U11348 (N_11348,N_8765,N_6301);
nand U11349 (N_11349,N_8866,N_7039);
nor U11350 (N_11350,N_8982,N_5274);
or U11351 (N_11351,N_6689,N_8130);
or U11352 (N_11352,N_9767,N_9846);
or U11353 (N_11353,N_7964,N_8843);
and U11354 (N_11354,N_7375,N_5534);
nand U11355 (N_11355,N_8216,N_9759);
nor U11356 (N_11356,N_8075,N_9793);
or U11357 (N_11357,N_5542,N_6818);
nor U11358 (N_11358,N_8929,N_5355);
and U11359 (N_11359,N_7931,N_8256);
or U11360 (N_11360,N_5941,N_5907);
and U11361 (N_11361,N_6538,N_9331);
or U11362 (N_11362,N_6360,N_5182);
nor U11363 (N_11363,N_9541,N_9755);
and U11364 (N_11364,N_9423,N_6025);
nand U11365 (N_11365,N_9356,N_7637);
and U11366 (N_11366,N_7129,N_8670);
or U11367 (N_11367,N_7885,N_6365);
or U11368 (N_11368,N_9236,N_6321);
nor U11369 (N_11369,N_7438,N_5135);
nor U11370 (N_11370,N_6100,N_6976);
or U11371 (N_11371,N_9823,N_8746);
and U11372 (N_11372,N_7080,N_6754);
nand U11373 (N_11373,N_8404,N_9311);
nor U11374 (N_11374,N_9007,N_7936);
nor U11375 (N_11375,N_9487,N_6345);
nor U11376 (N_11376,N_5646,N_5212);
and U11377 (N_11377,N_5524,N_7434);
xnor U11378 (N_11378,N_9320,N_5454);
nor U11379 (N_11379,N_9355,N_5837);
nand U11380 (N_11380,N_8372,N_8942);
or U11381 (N_11381,N_7653,N_8555);
or U11382 (N_11382,N_5239,N_9187);
nand U11383 (N_11383,N_8570,N_9997);
and U11384 (N_11384,N_9276,N_5546);
nor U11385 (N_11385,N_7900,N_6180);
or U11386 (N_11386,N_6710,N_7088);
nor U11387 (N_11387,N_6356,N_6839);
nor U11388 (N_11388,N_5660,N_6280);
or U11389 (N_11389,N_6546,N_6972);
or U11390 (N_11390,N_7403,N_9235);
and U11391 (N_11391,N_6447,N_7240);
nand U11392 (N_11392,N_7145,N_5287);
and U11393 (N_11393,N_8768,N_9290);
and U11394 (N_11394,N_9844,N_6828);
and U11395 (N_11395,N_7228,N_8937);
or U11396 (N_11396,N_8813,N_9798);
or U11397 (N_11397,N_9586,N_9502);
nand U11398 (N_11398,N_6010,N_7622);
nor U11399 (N_11399,N_5436,N_7960);
or U11400 (N_11400,N_6697,N_9388);
nand U11401 (N_11401,N_9562,N_5562);
nand U11402 (N_11402,N_9859,N_9682);
or U11403 (N_11403,N_8599,N_6659);
nand U11404 (N_11404,N_8142,N_5590);
nor U11405 (N_11405,N_5086,N_9367);
xnor U11406 (N_11406,N_9433,N_5850);
or U11407 (N_11407,N_9885,N_7793);
nor U11408 (N_11408,N_9382,N_8569);
or U11409 (N_11409,N_9521,N_5623);
xnor U11410 (N_11410,N_5853,N_6949);
and U11411 (N_11411,N_9027,N_6346);
or U11412 (N_11412,N_5692,N_5798);
or U11413 (N_11413,N_6917,N_7165);
and U11414 (N_11414,N_9531,N_8132);
or U11415 (N_11415,N_7617,N_6334);
or U11416 (N_11416,N_8329,N_9394);
nand U11417 (N_11417,N_8881,N_5885);
and U11418 (N_11418,N_9012,N_8339);
nor U11419 (N_11419,N_6530,N_8005);
or U11420 (N_11420,N_6568,N_8070);
nand U11421 (N_11421,N_5347,N_9146);
or U11422 (N_11422,N_9878,N_5992);
or U11423 (N_11423,N_5298,N_5180);
nor U11424 (N_11424,N_5866,N_5611);
or U11425 (N_11425,N_7765,N_7396);
nor U11426 (N_11426,N_6628,N_9471);
nand U11427 (N_11427,N_5377,N_9835);
and U11428 (N_11428,N_7595,N_9013);
or U11429 (N_11429,N_9625,N_9605);
nand U11430 (N_11430,N_9240,N_8465);
nand U11431 (N_11431,N_6878,N_8717);
nor U11432 (N_11432,N_8548,N_8316);
nor U11433 (N_11433,N_5158,N_7879);
nor U11434 (N_11434,N_6142,N_9557);
and U11435 (N_11435,N_6709,N_7277);
xnor U11436 (N_11436,N_5783,N_6299);
nor U11437 (N_11437,N_8074,N_5713);
and U11438 (N_11438,N_5401,N_9286);
nand U11439 (N_11439,N_7204,N_8260);
nand U11440 (N_11440,N_5632,N_6003);
nand U11441 (N_11441,N_9874,N_7163);
or U11442 (N_11442,N_5711,N_5578);
nand U11443 (N_11443,N_9950,N_8894);
and U11444 (N_11444,N_7841,N_6988);
nor U11445 (N_11445,N_9518,N_7664);
nor U11446 (N_11446,N_8343,N_8379);
and U11447 (N_11447,N_6206,N_6918);
nand U11448 (N_11448,N_6265,N_6604);
or U11449 (N_11449,N_9578,N_5547);
or U11450 (N_11450,N_9840,N_9340);
nand U11451 (N_11451,N_8718,N_6958);
nand U11452 (N_11452,N_9322,N_9600);
or U11453 (N_11453,N_9789,N_8170);
nand U11454 (N_11454,N_8897,N_8356);
or U11455 (N_11455,N_9238,N_6727);
and U11456 (N_11456,N_9226,N_6791);
and U11457 (N_11457,N_8516,N_5998);
and U11458 (N_11458,N_9177,N_9782);
and U11459 (N_11459,N_7399,N_8475);
or U11460 (N_11460,N_6640,N_5070);
nor U11461 (N_11461,N_5246,N_6192);
or U11462 (N_11462,N_5987,N_5727);
or U11463 (N_11463,N_5325,N_5348);
and U11464 (N_11464,N_6378,N_8608);
and U11465 (N_11465,N_8589,N_8360);
or U11466 (N_11466,N_7527,N_6369);
nor U11467 (N_11467,N_6513,N_9892);
or U11468 (N_11468,N_5600,N_5268);
nand U11469 (N_11469,N_5189,N_9706);
or U11470 (N_11470,N_7355,N_9769);
or U11471 (N_11471,N_8756,N_5897);
or U11472 (N_11472,N_7853,N_8920);
or U11473 (N_11473,N_7727,N_5282);
and U11474 (N_11474,N_8225,N_9775);
and U11475 (N_11475,N_5038,N_8250);
nand U11476 (N_11476,N_6203,N_6997);
nor U11477 (N_11477,N_9112,N_6049);
or U11478 (N_11478,N_6797,N_7820);
nor U11479 (N_11479,N_6787,N_5800);
and U11480 (N_11480,N_7867,N_6571);
and U11481 (N_11481,N_9801,N_8630);
and U11482 (N_11482,N_9854,N_9515);
nor U11483 (N_11483,N_8466,N_9851);
nand U11484 (N_11484,N_7862,N_5397);
nand U11485 (N_11485,N_9589,N_8402);
or U11486 (N_11486,N_6682,N_6312);
nand U11487 (N_11487,N_5449,N_8636);
and U11488 (N_11488,N_6566,N_7387);
and U11489 (N_11489,N_5388,N_7749);
or U11490 (N_11490,N_9018,N_8979);
or U11491 (N_11491,N_9485,N_9610);
or U11492 (N_11492,N_7876,N_9183);
and U11493 (N_11493,N_6864,N_9671);
nor U11494 (N_11494,N_9094,N_7568);
or U11495 (N_11495,N_7856,N_7221);
or U11496 (N_11496,N_6221,N_7280);
and U11497 (N_11497,N_6268,N_8022);
nand U11498 (N_11498,N_7641,N_9153);
and U11499 (N_11499,N_6817,N_8235);
nand U11500 (N_11500,N_8925,N_5235);
nand U11501 (N_11501,N_5222,N_8487);
nand U11502 (N_11502,N_6670,N_5184);
or U11503 (N_11503,N_7170,N_9726);
nor U11504 (N_11504,N_9196,N_6733);
and U11505 (N_11505,N_5619,N_5364);
nor U11506 (N_11506,N_9919,N_5090);
nor U11507 (N_11507,N_5766,N_5845);
nor U11508 (N_11508,N_8365,N_9690);
or U11509 (N_11509,N_6418,N_8204);
nor U11510 (N_11510,N_8640,N_8020);
or U11511 (N_11511,N_8148,N_9650);
or U11512 (N_11512,N_6978,N_7740);
nor U11513 (N_11513,N_9670,N_5067);
or U11514 (N_11514,N_5609,N_6617);
nand U11515 (N_11515,N_8567,N_9994);
nor U11516 (N_11516,N_5707,N_8351);
nor U11517 (N_11517,N_8287,N_5089);
nor U11518 (N_11518,N_7972,N_9178);
xnor U11519 (N_11519,N_7631,N_6000);
nor U11520 (N_11520,N_8563,N_7618);
nand U11521 (N_11521,N_5099,N_9116);
nor U11522 (N_11522,N_9189,N_9078);
nor U11523 (N_11523,N_9430,N_7064);
or U11524 (N_11524,N_6223,N_6806);
nor U11525 (N_11525,N_6101,N_7416);
nand U11526 (N_11526,N_8127,N_9140);
nand U11527 (N_11527,N_9397,N_9114);
nor U11528 (N_11528,N_7022,N_6593);
and U11529 (N_11529,N_5762,N_6620);
and U11530 (N_11530,N_9006,N_9818);
and U11531 (N_11531,N_5697,N_8986);
nor U11532 (N_11532,N_5937,N_9463);
nand U11533 (N_11533,N_5192,N_8722);
nor U11534 (N_11534,N_5521,N_5150);
or U11535 (N_11535,N_9684,N_5411);
nand U11536 (N_11536,N_6104,N_9440);
nand U11537 (N_11537,N_8758,N_7198);
nand U11538 (N_11538,N_7550,N_6671);
and U11539 (N_11539,N_6681,N_9512);
or U11540 (N_11540,N_8334,N_7319);
nor U11541 (N_11541,N_5119,N_9570);
nand U11542 (N_11542,N_6484,N_9482);
nand U11543 (N_11543,N_7669,N_9827);
nand U11544 (N_11544,N_7715,N_6720);
nand U11545 (N_11545,N_8252,N_6919);
nand U11546 (N_11546,N_6212,N_8091);
nand U11547 (N_11547,N_9582,N_7193);
nand U11548 (N_11548,N_7978,N_8676);
nor U11549 (N_11549,N_5631,N_5824);
or U11550 (N_11550,N_8972,N_8406);
and U11551 (N_11551,N_7988,N_9999);
or U11552 (N_11552,N_6273,N_9328);
and U11553 (N_11553,N_9891,N_9134);
and U11554 (N_11554,N_7293,N_5139);
or U11555 (N_11555,N_8731,N_9805);
and U11556 (N_11556,N_9848,N_6278);
or U11557 (N_11557,N_7124,N_6519);
or U11558 (N_11558,N_6572,N_7551);
nor U11559 (N_11559,N_5574,N_9601);
and U11560 (N_11560,N_8172,N_7056);
nand U11561 (N_11561,N_6691,N_8095);
or U11562 (N_11562,N_7017,N_8735);
and U11563 (N_11563,N_6066,N_8218);
nand U11564 (N_11564,N_8553,N_7405);
or U11565 (N_11565,N_7817,N_8320);
and U11566 (N_11566,N_5665,N_5683);
nand U11567 (N_11567,N_8198,N_9036);
nor U11568 (N_11568,N_5991,N_9427);
or U11569 (N_11569,N_8501,N_7125);
and U11570 (N_11570,N_6738,N_6061);
nor U11571 (N_11571,N_7157,N_5581);
and U11572 (N_11572,N_9136,N_9160);
and U11573 (N_11573,N_6930,N_8900);
nand U11574 (N_11574,N_8954,N_8507);
and U11575 (N_11575,N_7549,N_9761);
nor U11576 (N_11576,N_6850,N_8223);
nand U11577 (N_11577,N_8669,N_6224);
nand U11578 (N_11578,N_5211,N_5423);
nor U11579 (N_11579,N_6173,N_7753);
or U11580 (N_11580,N_9790,N_8603);
or U11581 (N_11581,N_9285,N_6085);
and U11582 (N_11582,N_9516,N_9940);
and U11583 (N_11583,N_9228,N_8179);
nor U11584 (N_11584,N_5236,N_7446);
nor U11585 (N_11585,N_6361,N_7565);
nor U11586 (N_11586,N_7601,N_8532);
and U11587 (N_11587,N_7346,N_8266);
and U11588 (N_11588,N_7100,N_6936);
nand U11589 (N_11589,N_8259,N_9715);
or U11590 (N_11590,N_9662,N_5868);
or U11591 (N_11591,N_8621,N_6339);
nor U11592 (N_11592,N_9713,N_8407);
nor U11593 (N_11593,N_6270,N_7386);
nand U11594 (N_11594,N_9750,N_8015);
nor U11595 (N_11595,N_8237,N_9737);
nor U11596 (N_11596,N_8462,N_6166);
nor U11597 (N_11597,N_9925,N_5564);
and U11598 (N_11598,N_5299,N_6908);
and U11599 (N_11599,N_6037,N_5442);
nand U11600 (N_11600,N_5767,N_6642);
or U11601 (N_11601,N_6589,N_9551);
and U11602 (N_11602,N_5403,N_7580);
or U11603 (N_11603,N_8232,N_6260);
or U11604 (N_11604,N_6896,N_9655);
nor U11605 (N_11605,N_6790,N_7548);
nand U11606 (N_11606,N_7728,N_9278);
nor U11607 (N_11607,N_9527,N_6536);
and U11608 (N_11608,N_8467,N_6287);
and U11609 (N_11609,N_8483,N_5645);
and U11610 (N_11610,N_6172,N_5315);
nand U11611 (N_11611,N_7985,N_9575);
and U11612 (N_11612,N_9221,N_7520);
and U11613 (N_11613,N_7234,N_6745);
and U11614 (N_11614,N_7374,N_8008);
nand U11615 (N_11615,N_5234,N_5755);
nor U11616 (N_11616,N_8641,N_9106);
nand U11617 (N_11617,N_9547,N_6035);
nand U11618 (N_11618,N_6966,N_5813);
and U11619 (N_11619,N_5048,N_8249);
and U11620 (N_11620,N_6045,N_7594);
nand U11621 (N_11621,N_7222,N_7401);
or U11622 (N_11622,N_6799,N_7496);
nor U11623 (N_11623,N_7735,N_8662);
nand U11624 (N_11624,N_5995,N_8523);
or U11625 (N_11625,N_5796,N_8160);
nand U11626 (N_11626,N_7072,N_5663);
and U11627 (N_11627,N_5644,N_7688);
nand U11628 (N_11628,N_5140,N_7895);
or U11629 (N_11629,N_7027,N_8893);
nand U11630 (N_11630,N_5954,N_7881);
or U11631 (N_11631,N_7202,N_7574);
nand U11632 (N_11632,N_7486,N_5802);
and U11633 (N_11633,N_8448,N_6621);
nand U11634 (N_11634,N_7590,N_5488);
and U11635 (N_11635,N_9698,N_8544);
or U11636 (N_11636,N_5902,N_6840);
nor U11637 (N_11637,N_5424,N_7347);
nand U11638 (N_11638,N_7613,N_7410);
and U11639 (N_11639,N_9403,N_7370);
nor U11640 (N_11640,N_8195,N_5255);
and U11641 (N_11641,N_8313,N_6374);
nor U11642 (N_11642,N_6497,N_7083);
nand U11643 (N_11643,N_7112,N_9247);
and U11644 (N_11644,N_7183,N_5431);
nor U11645 (N_11645,N_7333,N_9350);
or U11646 (N_11646,N_7349,N_5228);
nor U11647 (N_11647,N_6947,N_9872);
nand U11648 (N_11648,N_9259,N_7668);
nand U11649 (N_11649,N_5159,N_7676);
nand U11650 (N_11650,N_5069,N_7928);
nor U11651 (N_11651,N_5479,N_8335);
or U11652 (N_11652,N_6890,N_8338);
nor U11653 (N_11653,N_6561,N_9086);
and U11654 (N_11654,N_9223,N_6023);
nor U11655 (N_11655,N_9241,N_5899);
and U11656 (N_11656,N_7210,N_6763);
or U11657 (N_11657,N_7572,N_9597);
nor U11658 (N_11658,N_5441,N_7440);
nor U11659 (N_11659,N_6871,N_9627);
nand U11660 (N_11660,N_8430,N_7360);
nand U11661 (N_11661,N_6831,N_7888);
and U11662 (N_11662,N_5961,N_7501);
and U11663 (N_11663,N_6401,N_7742);
xor U11664 (N_11664,N_9852,N_8943);
and U11665 (N_11665,N_6465,N_7323);
nor U11666 (N_11666,N_5918,N_6537);
nand U11667 (N_11667,N_7529,N_9795);
and U11668 (N_11668,N_9399,N_9052);
and U11669 (N_11669,N_8197,N_6753);
or U11670 (N_11670,N_9530,N_7802);
and U11671 (N_11671,N_5908,N_5290);
or U11672 (N_11672,N_9631,N_9450);
or U11673 (N_11673,N_7341,N_6826);
and U11674 (N_11674,N_5310,N_6898);
or U11675 (N_11675,N_8059,N_5144);
and U11676 (N_11676,N_7377,N_7420);
and U11677 (N_11677,N_6363,N_5036);
or U11678 (N_11678,N_5979,N_5185);
xor U11679 (N_11679,N_5252,N_7632);
and U11680 (N_11680,N_6920,N_6396);
or U11681 (N_11681,N_8347,N_6816);
and U11682 (N_11682,N_8534,N_8315);
or U11683 (N_11683,N_8606,N_7258);
nor U11684 (N_11684,N_5248,N_6297);
or U11685 (N_11685,N_8763,N_7150);
nor U11686 (N_11686,N_8622,N_9774);
and U11687 (N_11687,N_8268,N_7956);
nand U11688 (N_11688,N_6877,N_7534);
or U11689 (N_11689,N_8810,N_8412);
nand U11690 (N_11690,N_7474,N_9831);
or U11691 (N_11691,N_7127,N_9055);
nor U11692 (N_11692,N_8234,N_5482);
and U11693 (N_11693,N_5191,N_8028);
and U11694 (N_11694,N_7389,N_8996);
or U11695 (N_11695,N_8117,N_8526);
and U11696 (N_11696,N_6606,N_8078);
nor U11697 (N_11697,N_9733,N_7245);
nand U11698 (N_11698,N_8045,N_9896);
and U11699 (N_11699,N_8352,N_5694);
nor U11700 (N_11700,N_9895,N_9454);
nand U11701 (N_11701,N_8244,N_7773);
and U11702 (N_11702,N_6955,N_5217);
nor U11703 (N_11703,N_5654,N_5714);
nor U11704 (N_11704,N_8086,N_8538);
nand U11705 (N_11705,N_5527,N_5238);
and U11706 (N_11706,N_7747,N_8854);
xnor U11707 (N_11707,N_8655,N_5056);
and U11708 (N_11708,N_9452,N_8192);
and U11709 (N_11709,N_9821,N_5445);
and U11710 (N_11710,N_6290,N_6909);
nand U11711 (N_11711,N_7935,N_8528);
nor U11712 (N_11712,N_5726,N_6613);
or U11713 (N_11713,N_9039,N_6332);
and U11714 (N_11714,N_5215,N_6128);
nor U11715 (N_11715,N_9309,N_5404);
xor U11716 (N_11716,N_6457,N_5844);
and U11717 (N_11717,N_5286,N_7158);
and U11718 (N_11718,N_8009,N_7832);
nand U11719 (N_11719,N_9151,N_9214);
and U11720 (N_11720,N_5329,N_8699);
nor U11721 (N_11721,N_9717,N_8264);
and U11722 (N_11722,N_7539,N_8308);
and U11723 (N_11723,N_8691,N_5219);
nand U11724 (N_11724,N_5088,N_7957);
nand U11725 (N_11725,N_8023,N_8161);
nor U11726 (N_11726,N_9483,N_8927);
and U11727 (N_11727,N_7162,N_7882);
and U11728 (N_11728,N_5506,N_7525);
and U11729 (N_11729,N_8189,N_8180);
nor U11730 (N_11730,N_5887,N_5302);
or U11731 (N_11731,N_9067,N_7304);
nor U11732 (N_11732,N_5988,N_7829);
nand U11733 (N_11733,N_7610,N_8494);
nor U11734 (N_11734,N_5799,N_5074);
nor U11735 (N_11735,N_6481,N_6041);
nand U11736 (N_11736,N_8506,N_7237);
nand U11737 (N_11737,N_8042,N_6660);
nand U11738 (N_11738,N_9730,N_9343);
nor U11739 (N_11739,N_8281,N_7291);
and U11740 (N_11740,N_7028,N_6542);
nand U11741 (N_11741,N_8145,N_5492);
nor U11742 (N_11742,N_6577,N_8916);
nor U11743 (N_11743,N_5352,N_7723);
nand U11744 (N_11744,N_8901,N_5387);
nand U11745 (N_11745,N_5808,N_9833);
nor U11746 (N_11746,N_8505,N_6215);
or U11747 (N_11747,N_9495,N_6090);
nor U11748 (N_11748,N_5742,N_8812);
and U11749 (N_11749,N_7325,N_5410);
or U11750 (N_11750,N_7606,N_7279);
nand U11751 (N_11751,N_7133,N_5997);
and U11752 (N_11752,N_5769,N_9890);
nor U11753 (N_11753,N_5780,N_8076);
nand U11754 (N_11754,N_9407,N_6502);
and U11755 (N_11755,N_8542,N_5922);
nor U11756 (N_11756,N_9401,N_7545);
and U11757 (N_11757,N_7476,N_7831);
or U11758 (N_11758,N_5031,N_6225);
nor U11759 (N_11759,N_7390,N_8629);
and U11760 (N_11760,N_7764,N_9091);
or U11761 (N_11761,N_9257,N_5656);
nand U11762 (N_11762,N_5608,N_8774);
nand U11763 (N_11763,N_7691,N_8877);
nor U11764 (N_11764,N_7584,N_6813);
and U11765 (N_11765,N_9460,N_6498);
nor U11766 (N_11766,N_5308,N_7643);
and U11767 (N_11767,N_8080,N_5311);
and U11768 (N_11768,N_8396,N_8257);
nand U11769 (N_11769,N_7672,N_6162);
nor U11770 (N_11770,N_8380,N_6030);
and U11771 (N_11771,N_5483,N_6450);
xnor U11772 (N_11772,N_8687,N_5551);
or U11773 (N_11773,N_8949,N_5336);
nand U11774 (N_11774,N_8119,N_8783);
xor U11775 (N_11775,N_5068,N_6923);
nor U11776 (N_11776,N_8748,N_6752);
and U11777 (N_11777,N_6472,N_5353);
and U11778 (N_11778,N_9344,N_7911);
nor U11779 (N_11779,N_8890,N_5648);
nand U11780 (N_11780,N_7706,N_9135);
nand U11781 (N_11781,N_8149,N_7007);
nor U11782 (N_11782,N_9628,N_6636);
and U11783 (N_11783,N_5595,N_6493);
nand U11784 (N_11784,N_7624,N_6492);
nor U11785 (N_11785,N_6236,N_7081);
nor U11786 (N_11786,N_9470,N_8302);
nor U11787 (N_11787,N_7365,N_8984);
and U11788 (N_11788,N_7737,N_9590);
nor U11789 (N_11789,N_6951,N_8125);
and U11790 (N_11790,N_8841,N_7996);
and U11791 (N_11791,N_5945,N_5668);
and U11792 (N_11792,N_9869,N_7063);
or U11793 (N_11793,N_6230,N_8525);
nand U11794 (N_11794,N_6242,N_9792);
or U11795 (N_11795,N_9581,N_9288);
and U11796 (N_11796,N_8697,N_7432);
or U11797 (N_11797,N_6111,N_6343);
and U11798 (N_11798,N_6118,N_5102);
nor U11799 (N_11799,N_5593,N_7854);
and U11800 (N_11800,N_5380,N_8863);
nor U11801 (N_11801,N_5163,N_9947);
nand U11802 (N_11802,N_7181,N_9745);
and U11803 (N_11803,N_8614,N_8867);
nor U11804 (N_11804,N_9295,N_7435);
nand U11805 (N_11805,N_7629,N_8598);
nor U11806 (N_11806,N_5027,N_8837);
and U11807 (N_11807,N_9724,N_9870);
nor U11808 (N_11808,N_6652,N_6338);
or U11809 (N_11809,N_7573,N_7690);
nand U11810 (N_11810,N_7225,N_9049);
nand U11811 (N_11811,N_5168,N_9513);
nand U11812 (N_11812,N_7684,N_8912);
nor U11813 (N_11813,N_7126,N_7563);
nand U11814 (N_11814,N_7901,N_7106);
and U11815 (N_11815,N_7523,N_8977);
and U11816 (N_11816,N_8041,N_8088);
or U11817 (N_11817,N_6349,N_8027);
nor U11818 (N_11818,N_9517,N_8695);
nand U11819 (N_11819,N_6541,N_6792);
or U11820 (N_11820,N_9681,N_6847);
nand U11821 (N_11821,N_9090,N_8780);
or U11822 (N_11822,N_7208,N_7426);
and U11823 (N_11823,N_5179,N_6703);
nand U11824 (N_11824,N_8393,N_5035);
nand U11825 (N_11825,N_9491,N_8919);
nand U11826 (N_11826,N_9283,N_8779);
and U11827 (N_11827,N_8826,N_8760);
and U11828 (N_11828,N_6201,N_8083);
nand U11829 (N_11829,N_7067,N_9411);
and U11830 (N_11830,N_9533,N_5974);
or U11831 (N_11831,N_6006,N_8685);
and U11832 (N_11832,N_9457,N_9902);
or U11833 (N_11833,N_5956,N_7026);
nand U11834 (N_11834,N_8272,N_8588);
nand U11835 (N_11835,N_6074,N_8572);
nor U11836 (N_11836,N_5647,N_9345);
xnor U11837 (N_11837,N_5178,N_9843);
nor U11838 (N_11838,N_7702,N_5369);
nand U11839 (N_11839,N_7478,N_7354);
nand U11840 (N_11840,N_6174,N_9921);
and U11841 (N_11841,N_5972,N_5793);
nor U11842 (N_11842,N_5699,N_6129);
nor U11843 (N_11843,N_6504,N_7001);
nand U11844 (N_11844,N_9415,N_7850);
or U11845 (N_11845,N_8759,N_9459);
or U11846 (N_11846,N_6520,N_7107);
nand U11847 (N_11847,N_7113,N_5548);
and U11848 (N_11848,N_6295,N_5931);
and U11849 (N_11849,N_7322,N_8276);
and U11850 (N_11850,N_9700,N_5855);
or U11851 (N_11851,N_6903,N_5365);
or U11852 (N_11852,N_7886,N_8885);
xnor U11853 (N_11853,N_7852,N_7609);
and U11854 (N_11854,N_7393,N_9980);
and U11855 (N_11855,N_6138,N_7557);
nor U11856 (N_11856,N_8019,N_6056);
nand U11857 (N_11857,N_8723,N_8797);
xnor U11858 (N_11858,N_7828,N_6460);
xnor U11859 (N_11859,N_6266,N_5572);
nor U11860 (N_11860,N_6582,N_5516);
or U11861 (N_11861,N_6662,N_7794);
xor U11862 (N_11862,N_9732,N_7011);
and U11863 (N_11863,N_7134,N_5712);
xor U11864 (N_11864,N_7316,N_6518);
nor U11865 (N_11865,N_8817,N_6416);
nor U11866 (N_11866,N_5224,N_7812);
or U11867 (N_11867,N_6544,N_8474);
nor U11868 (N_11868,N_9707,N_8948);
or U11869 (N_11869,N_5275,N_8659);
nor U11870 (N_11870,N_9501,N_7249);
nor U11871 (N_11871,N_5733,N_6841);
or U11872 (N_11872,N_6412,N_5896);
nor U11873 (N_11873,N_8625,N_8500);
nand U11874 (N_11874,N_6109,N_8426);
or U11875 (N_11875,N_7086,N_5321);
and U11876 (N_11876,N_9951,N_9016);
nand U11877 (N_11877,N_9137,N_6133);
and U11878 (N_11878,N_7555,N_8370);
or U11879 (N_11879,N_6590,N_6772);
nand U11880 (N_11880,N_6549,N_5869);
and U11881 (N_11881,N_7421,N_9198);
or U11882 (N_11882,N_5693,N_7156);
nor U11883 (N_11883,N_9219,N_9929);
nand U11884 (N_11884,N_7506,N_6501);
and U11885 (N_11885,N_9762,N_9567);
or U11886 (N_11886,N_6262,N_7772);
nand U11887 (N_11887,N_6448,N_7947);
and U11888 (N_11888,N_6461,N_9363);
or U11889 (N_11889,N_7755,N_7348);
nor U11890 (N_11890,N_5975,N_5816);
and U11891 (N_11891,N_6759,N_5734);
or U11892 (N_11892,N_8453,N_9923);
nor U11893 (N_11893,N_8044,N_5091);
or U11894 (N_11894,N_9934,N_8541);
or U11895 (N_11895,N_9469,N_9791);
and U11896 (N_11896,N_6024,N_5519);
or U11897 (N_11897,N_5305,N_8808);
or U11898 (N_11898,N_8116,N_8704);
nor U11899 (N_11899,N_9486,N_7571);
and U11900 (N_11900,N_7968,N_8463);
nand U11901 (N_11901,N_5161,N_7783);
nand U11902 (N_11902,N_9149,N_6179);
nor U11903 (N_11903,N_8609,N_9689);
or U11904 (N_11904,N_7260,N_7364);
nor U11905 (N_11905,N_5858,N_9077);
or U11906 (N_11906,N_5373,N_5591);
and U11907 (N_11907,N_9100,N_7701);
nand U11908 (N_11908,N_8459,N_5585);
nand U11909 (N_11909,N_7604,N_5731);
nor U11910 (N_11910,N_5361,N_5883);
nor U11911 (N_11911,N_6961,N_5419);
nand U11912 (N_11912,N_5722,N_6388);
or U11913 (N_11913,N_9893,N_5774);
xor U11914 (N_11914,N_7305,N_5451);
nor U11915 (N_11915,N_9022,N_7514);
and U11916 (N_11916,N_6149,N_5849);
nand U11917 (N_11917,N_9364,N_6717);
and U11918 (N_11918,N_5079,N_6423);
nand U11919 (N_11919,N_6425,N_6434);
nand U11920 (N_11920,N_9604,N_7295);
or U11921 (N_11921,N_6116,N_6475);
or U11922 (N_11922,N_9405,N_7925);
and U11923 (N_11923,N_7959,N_7460);
and U11924 (N_11924,N_7096,N_5635);
nor U11925 (N_11925,N_7443,N_6861);
and U11926 (N_11926,N_6894,N_8100);
and U11927 (N_11927,N_8673,N_6274);
nor U11928 (N_11928,N_7489,N_8054);
and U11929 (N_11929,N_8790,N_9208);
nand U11930 (N_11930,N_6643,N_8861);
or U11931 (N_11931,N_5133,N_8745);
or U11932 (N_11932,N_7751,N_9327);
nand U11933 (N_11933,N_5020,N_9270);
nor U11934 (N_11934,N_9357,N_6141);
and U11935 (N_11935,N_9624,N_8554);
xor U11936 (N_11936,N_6125,N_9986);
nor U11937 (N_11937,N_7950,N_6801);
or U11938 (N_11938,N_8440,N_7016);
or U11939 (N_11939,N_6007,N_8654);
or U11940 (N_11940,N_5597,N_5295);
nand U11941 (N_11941,N_7345,N_6800);
nand U11942 (N_11942,N_9760,N_9534);
nand U11943 (N_11943,N_8101,N_8978);
nand U11944 (N_11944,N_9956,N_9992);
or U11945 (N_11945,N_8587,N_7558);
nand U11946 (N_11946,N_7422,N_8605);
or U11947 (N_11947,N_7546,N_5335);
or U11948 (N_11948,N_9734,N_7902);
nand U11949 (N_11949,N_7620,N_8126);
nand U11950 (N_11950,N_5478,N_7874);
nor U11951 (N_11951,N_9071,N_8579);
or U11952 (N_11952,N_6271,N_9699);
nand U11953 (N_11953,N_6627,N_7503);
or U11954 (N_11954,N_6383,N_8416);
and U11955 (N_11955,N_5341,N_8174);
nor U11956 (N_11956,N_5077,N_5458);
or U11957 (N_11957,N_9803,N_6551);
and U11958 (N_11958,N_9072,N_5206);
nor U11959 (N_11959,N_9066,N_7308);
nor U11960 (N_11960,N_9374,N_8883);
nand U11961 (N_11961,N_8510,N_6184);
nand U11962 (N_11962,N_7849,N_9026);
nor U11963 (N_11963,N_9927,N_9694);
or U11964 (N_11964,N_9317,N_5760);
nand U11965 (N_11965,N_9336,N_8945);
nor U11966 (N_11966,N_8258,N_6719);
and U11967 (N_11967,N_8604,N_8690);
and U11968 (N_11968,N_9010,N_6822);
and U11969 (N_11969,N_8577,N_5838);
nand U11970 (N_11970,N_6673,N_6728);
or U11971 (N_11971,N_7712,N_9933);
and U11972 (N_11972,N_6256,N_5370);
or U11973 (N_11973,N_7499,N_8773);
xnor U11974 (N_11974,N_6407,N_6591);
and U11975 (N_11975,N_9128,N_9884);
nand U11976 (N_11976,N_5951,N_6555);
nor U11977 (N_11977,N_8357,N_7942);
nand U11978 (N_11978,N_9608,N_5288);
or U11979 (N_11979,N_8509,N_9354);
or U11980 (N_11980,N_6022,N_5204);
or U11981 (N_11981,N_9549,N_6809);
nand U11982 (N_11982,N_5004,N_7175);
or U11983 (N_11983,N_8184,N_5103);
xnor U11984 (N_11984,N_7979,N_9157);
nand U11985 (N_11985,N_6490,N_6683);
nor U11986 (N_11986,N_9984,N_9376);
and U11987 (N_11987,N_6237,N_8381);
nor U11988 (N_11988,N_7252,N_5152);
nand U11989 (N_11989,N_6722,N_7567);
or U11990 (N_11990,N_8736,N_9264);
nand U11991 (N_11991,N_8021,N_5138);
and U11992 (N_11992,N_5015,N_8464);
and U11993 (N_11993,N_7084,N_9674);
and U11994 (N_11994,N_5903,N_6969);
nor U11995 (N_11995,N_6782,N_5225);
nand U11996 (N_11996,N_5687,N_7318);
nand U11997 (N_11997,N_5511,N_9847);
or U11998 (N_11998,N_9504,N_8110);
or U11999 (N_11999,N_6876,N_9079);
nor U12000 (N_12000,N_9170,N_9957);
or U12001 (N_12001,N_8366,N_5765);
nor U12002 (N_12002,N_7907,N_7014);
and U12003 (N_12003,N_6353,N_5582);
nand U12004 (N_12004,N_6306,N_5251);
nor U12005 (N_12005,N_8484,N_9000);
or U12006 (N_12006,N_7729,N_8616);
or U12007 (N_12007,N_8981,N_9373);
or U12008 (N_12008,N_6322,N_7719);
nand U12009 (N_12009,N_7776,N_9981);
and U12010 (N_12010,N_8627,N_5752);
and U12011 (N_12011,N_5028,N_9084);
or U12012 (N_12012,N_5843,N_7230);
and U12013 (N_12013,N_6998,N_7101);
nor U12014 (N_12014,N_6190,N_7708);
nand U12015 (N_12015,N_7484,N_8077);
xnor U12016 (N_12016,N_8868,N_6021);
and U12017 (N_12017,N_5629,N_6835);
nand U12018 (N_12018,N_8794,N_8053);
or U12019 (N_12019,N_7408,N_9532);
or U12020 (N_12020,N_8069,N_7667);
and U12021 (N_12021,N_6922,N_8857);
and U12022 (N_12022,N_8864,N_6948);
or U12023 (N_12023,N_9369,N_5044);
and U12024 (N_12024,N_6882,N_8046);
nor U12025 (N_12025,N_5846,N_8173);
and U12026 (N_12026,N_6068,N_7872);
and U12027 (N_12027,N_7599,N_5963);
nand U12028 (N_12028,N_5831,N_5452);
nor U12029 (N_12029,N_8261,N_8162);
nand U12030 (N_12030,N_9123,N_9911);
nand U12031 (N_12031,N_8495,N_6042);
nand U12032 (N_12032,N_6402,N_5779);
or U12033 (N_12033,N_7329,N_9948);
xnor U12034 (N_12034,N_7248,N_6069);
or U12035 (N_12035,N_5181,N_9442);
nand U12036 (N_12036,N_8188,N_8081);
nor U12037 (N_12037,N_7692,N_6285);
nor U12038 (N_12038,N_8144,N_7340);
nand U12039 (N_12039,N_8747,N_8515);
nor U12040 (N_12040,N_9428,N_7298);
nand U12041 (N_12041,N_6873,N_8064);
or U12042 (N_12042,N_6605,N_7361);
and U12043 (N_12043,N_8744,N_5877);
or U12044 (N_12044,N_6002,N_5545);
nor U12045 (N_12045,N_7992,N_7178);
nor U12046 (N_12046,N_7536,N_8456);
nand U12047 (N_12047,N_5532,N_8353);
and U12048 (N_12048,N_5716,N_8350);
and U12049 (N_12049,N_8803,N_7154);
nand U12050 (N_12050,N_6964,N_9498);
nor U12051 (N_12051,N_8147,N_6718);
nor U12052 (N_12052,N_6715,N_8624);
nand U12053 (N_12053,N_8870,N_8178);
and U12054 (N_12054,N_7908,N_9599);
nand U12055 (N_12055,N_7554,N_5637);
nand U12056 (N_12056,N_9812,N_9651);
nand U12057 (N_12057,N_5297,N_7705);
nor U12058 (N_12058,N_6851,N_9139);
nand U12059 (N_12059,N_9560,N_6164);
and U12060 (N_12060,N_9916,N_5841);
or U12061 (N_12061,N_5830,N_6641);
nor U12062 (N_12062,N_7269,N_6289);
or U12063 (N_12063,N_7205,N_7188);
and U12064 (N_12064,N_8492,N_5468);
and U12065 (N_12065,N_9024,N_6044);
nand U12066 (N_12066,N_9326,N_8896);
or U12067 (N_12067,N_9794,N_6178);
nand U12068 (N_12068,N_7024,N_8473);
or U12069 (N_12069,N_8633,N_6442);
and U12070 (N_12070,N_5672,N_6469);
and U12071 (N_12071,N_6901,N_7840);
nand U12072 (N_12072,N_5391,N_6219);
nand U12073 (N_12073,N_7639,N_5081);
and U12074 (N_12074,N_8886,N_6175);
or U12075 (N_12075,N_7338,N_5882);
and U12076 (N_12076,N_9038,N_6532);
nand U12077 (N_12077,N_7166,N_8029);
nor U12078 (N_12078,N_5949,N_9771);
or U12079 (N_12079,N_6330,N_5695);
or U12080 (N_12080,N_9480,N_8155);
and U12081 (N_12081,N_7767,N_7111);
and U12082 (N_12082,N_9195,N_5367);
nor U12083 (N_12083,N_5962,N_6186);
xnor U12084 (N_12084,N_7798,N_8330);
nand U12085 (N_12085,N_6653,N_5170);
and U12086 (N_12086,N_9115,N_8733);
nand U12087 (N_12087,N_6937,N_9070);
nor U12088 (N_12088,N_7373,N_8230);
nor U12089 (N_12089,N_9946,N_6559);
or U12090 (N_12090,N_9419,N_5812);
and U12091 (N_12091,N_9615,N_9958);
and U12092 (N_12092,N_7625,N_7934);
nor U12093 (N_12093,N_9566,N_7331);
and U12094 (N_12094,N_8595,N_6716);
or U12095 (N_12095,N_9654,N_7339);
and U12096 (N_12096,N_7029,N_9081);
nand U12097 (N_12097,N_8656,N_6154);
and U12098 (N_12098,N_9389,N_5343);
or U12099 (N_12099,N_7138,N_6601);
and U12100 (N_12100,N_5890,N_6187);
nor U12101 (N_12101,N_6494,N_5216);
nor U12102 (N_12102,N_7471,N_5710);
and U12103 (N_12103,N_8194,N_6522);
nor U12104 (N_12104,N_7378,N_9853);
xnor U12105 (N_12105,N_7871,N_9524);
nand U12106 (N_12106,N_7119,N_6246);
and U12107 (N_12107,N_5046,N_8265);
or U12108 (N_12108,N_5051,N_6714);
nor U12109 (N_12109,N_5891,N_7873);
xnor U12110 (N_12110,N_9875,N_8071);
nand U12111 (N_12111,N_6925,N_6267);
nor U12112 (N_12112,N_8661,N_8834);
nand U12113 (N_12113,N_7990,N_8314);
xor U12114 (N_12114,N_7602,N_7726);
nand U12115 (N_12115,N_7469,N_5371);
nor U12116 (N_12116,N_6623,N_9967);
or U12117 (N_12117,N_8638,N_8245);
and U12118 (N_12118,N_9702,N_8011);
or U12119 (N_12119,N_7562,N_7285);
or U12120 (N_12120,N_9716,N_5568);
or U12121 (N_12121,N_7049,N_8383);
or U12122 (N_12122,N_6326,N_9117);
nand U12123 (N_12123,N_9680,N_7185);
nand U12124 (N_12124,N_8294,N_7261);
nor U12125 (N_12125,N_5981,N_8375);
and U12126 (N_12126,N_5996,N_5916);
or U12127 (N_12127,N_8971,N_9441);
nand U12128 (N_12128,N_8107,N_5622);
and U12129 (N_12129,N_9068,N_5671);
or U12130 (N_12130,N_8400,N_6768);
nor U12131 (N_12131,N_9065,N_8318);
nor U12132 (N_12132,N_7488,N_7855);
xnor U12133 (N_12133,N_7894,N_8217);
or U12134 (N_12134,N_6644,N_8368);
and U12135 (N_12135,N_7683,N_7148);
nand U12136 (N_12136,N_7759,N_5504);
nor U12137 (N_12137,N_8286,N_9961);
nand U12138 (N_12138,N_8715,N_8362);
nand U12139 (N_12139,N_9167,N_6953);
and U12140 (N_12140,N_9019,N_7025);
or U12141 (N_12141,N_5009,N_9477);
and U12142 (N_12142,N_6977,N_6302);
nor U12143 (N_12143,N_6677,N_7136);
nand U12144 (N_12144,N_5223,N_9564);
nor U12145 (N_12145,N_7380,N_9348);
or U12146 (N_12146,N_7952,N_9044);
or U12147 (N_12147,N_7412,N_9069);
or U12148 (N_12148,N_9579,N_6607);
or U12149 (N_12149,N_6382,N_5497);
nand U12150 (N_12150,N_6837,N_9514);
nand U12151 (N_12151,N_7495,N_5651);
nand U12152 (N_12152,N_8772,N_7842);
and U12153 (N_12153,N_7053,N_5706);
and U12154 (N_12154,N_8968,N_7459);
nand U12155 (N_12155,N_9119,N_6553);
nor U12156 (N_12156,N_5659,N_9324);
nand U12157 (N_12157,N_7320,N_5342);
and U12158 (N_12158,N_5378,N_9406);
nor U12159 (N_12159,N_7312,N_9215);
nor U12160 (N_12160,N_7967,N_6213);
and U12161 (N_12161,N_5444,N_7192);
nor U12162 (N_12162,N_8388,N_9544);
xor U12163 (N_12163,N_5116,N_9314);
and U12164 (N_12164,N_8274,N_5443);
nor U12165 (N_12165,N_5989,N_5641);
or U12166 (N_12166,N_7332,N_9786);
and U12167 (N_12167,N_8580,N_5253);
and U12168 (N_12168,N_7836,N_8452);
nor U12169 (N_12169,N_8164,N_6303);
nor U12170 (N_12170,N_5925,N_6160);
nor U12171 (N_12171,N_8328,N_9267);
nor U12172 (N_12172,N_6868,N_5827);
and U12173 (N_12173,N_5289,N_8543);
nand U12174 (N_12174,N_8547,N_6558);
nor U12175 (N_12175,N_6696,N_9727);
nor U12176 (N_12176,N_6232,N_9757);
xnor U12177 (N_12177,N_7623,N_5636);
and U12178 (N_12178,N_5429,N_6573);
nand U12179 (N_12179,N_6944,N_7095);
nor U12180 (N_12180,N_7937,N_6119);
nand U12181 (N_12181,N_5748,N_7636);
or U12182 (N_12182,N_6185,N_8395);
or U12183 (N_12183,N_7830,N_5220);
and U12184 (N_12184,N_6531,N_9120);
and U12185 (N_12185,N_7914,N_9377);
nor U12186 (N_12186,N_8491,N_8050);
nand U12187 (N_12187,N_5735,N_8093);
nor U12188 (N_12188,N_5427,N_5039);
nand U12189 (N_12189,N_5269,N_7670);
nor U12190 (N_12190,N_7944,N_5406);
nor U12191 (N_12191,N_5111,N_8199);
nor U12192 (N_12192,N_9174,N_9939);
nor U12193 (N_12193,N_9110,N_7251);
and U12194 (N_12194,N_5146,N_7678);
and U12195 (N_12195,N_9246,N_7977);
nand U12196 (N_12196,N_5921,N_8764);
or U12197 (N_12197,N_6093,N_5213);
or U12198 (N_12198,N_6855,N_5487);
or U12199 (N_12199,N_7707,N_5344);
or U12200 (N_12200,N_8134,N_8823);
or U12201 (N_12201,N_7153,N_5856);
nand U12202 (N_12202,N_6778,N_5227);
nand U12203 (N_12203,N_5040,N_9573);
or U12204 (N_12204,N_5337,N_8694);
and U12205 (N_12205,N_6842,N_6815);
nand U12206 (N_12206,N_6404,N_9539);
and U12207 (N_12207,N_8397,N_8926);
and U12208 (N_12208,N_5771,N_8962);
nand U12209 (N_12209,N_9988,N_6385);
nand U12210 (N_12210,N_8398,N_9932);
or U12211 (N_12211,N_7395,N_5162);
or U12212 (N_12212,N_6633,N_8364);
or U12213 (N_12213,N_7139,N_5773);
nor U12214 (N_12214,N_9200,N_8683);
nand U12215 (N_12215,N_5408,N_5832);
nand U12216 (N_12216,N_7206,N_8422);
nor U12217 (N_12217,N_7362,N_8392);
and U12218 (N_12218,N_8336,N_8908);
or U12219 (N_12219,N_9266,N_6092);
and U12220 (N_12220,N_7078,N_9383);
or U12221 (N_12221,N_5327,N_7462);
or U12222 (N_12222,N_5480,N_5108);
nand U12223 (N_12223,N_8319,N_5861);
nor U12224 (N_12224,N_7638,N_9865);
xnor U12225 (N_12225,N_8115,N_5469);
or U12226 (N_12226,N_7199,N_8152);
or U12227 (N_12227,N_7788,N_5789);
nand U12228 (N_12228,N_8788,N_7965);
and U12229 (N_12229,N_7172,N_5142);
or U12230 (N_12230,N_9291,N_8186);
or U12231 (N_12231,N_8414,N_7479);
xnor U12232 (N_12232,N_5847,N_5705);
nor U12233 (N_12233,N_6761,N_9008);
or U12234 (N_12234,N_5718,N_8215);
or U12235 (N_12235,N_5143,N_7652);
and U12236 (N_12236,N_8436,N_8930);
or U12237 (N_12237,N_9273,N_6762);
and U12238 (N_12238,N_5596,N_6389);
nor U12239 (N_12239,N_5685,N_7897);
nand U12240 (N_12240,N_7792,N_7782);
nor U12241 (N_12241,N_9845,N_6996);
and U12242 (N_12242,N_9926,N_5514);
nand U12243 (N_12243,N_7646,N_5784);
and U12244 (N_12244,N_6999,N_9321);
nor U12245 (N_12245,N_6200,N_5970);
nor U12246 (N_12246,N_8106,N_5195);
nor U12247 (N_12247,N_8055,N_8428);
and U12248 (N_12248,N_9234,N_5915);
and U12249 (N_12249,N_7757,N_5893);
nor U12250 (N_12250,N_9462,N_7468);
nor U12251 (N_12251,N_8840,N_6625);
nand U12252 (N_12252,N_7790,N_8384);
and U12253 (N_12253,N_8323,N_9358);
and U12254 (N_12254,N_6120,N_5621);
nand U12255 (N_12255,N_9289,N_5892);
nand U12256 (N_12256,N_6793,N_9710);
nand U12257 (N_12257,N_9387,N_8168);
and U12258 (N_12258,N_5024,N_5684);
nor U12259 (N_12259,N_6534,N_6456);
or U12260 (N_12260,N_7105,N_5686);
xnor U12261 (N_12261,N_9201,N_7116);
nor U12262 (N_12262,N_8601,N_7585);
nand U12263 (N_12263,N_8708,N_7451);
or U12264 (N_12264,N_5770,N_7388);
nor U12265 (N_12265,N_6318,N_9109);
nand U12266 (N_12266,N_7259,N_8108);
nand U12267 (N_12267,N_8228,N_5721);
or U12268 (N_12268,N_8639,N_5386);
nor U12269 (N_12269,N_5017,N_8781);
and U12270 (N_12270,N_5481,N_8030);
and U12271 (N_12271,N_5421,N_7954);
nand U12272 (N_12272,N_6170,N_8409);
and U12273 (N_12273,N_6921,N_8410);
or U12274 (N_12274,N_8557,N_5484);
and U12275 (N_12275,N_6626,N_7123);
nor U12276 (N_12276,N_7483,N_5205);
xnor U12277 (N_12277,N_9489,N_9108);
or U12278 (N_12278,N_5630,N_8647);
or U12279 (N_12279,N_9556,N_5749);
and U12280 (N_12280,N_9060,N_6845);
and U12281 (N_12281,N_7685,N_8341);
nand U12282 (N_12282,N_9842,N_7290);
and U12283 (N_12283,N_6934,N_5101);
nor U12284 (N_12284,N_8682,N_8399);
or U12285 (N_12285,N_6609,N_5266);
nor U12286 (N_12286,N_9602,N_6634);
xor U12287 (N_12287,N_6610,N_8770);
and U12288 (N_12288,N_5911,N_7187);
or U12289 (N_12289,N_6464,N_9105);
and U12290 (N_12290,N_5607,N_7372);
nor U12291 (N_12291,N_5465,N_8043);
and U12292 (N_12292,N_6912,N_5599);
and U12293 (N_12293,N_7140,N_5906);
and U12294 (N_12294,N_8304,N_5021);
and U12295 (N_12295,N_7823,N_7068);
or U12296 (N_12296,N_6143,N_5613);
nor U12297 (N_12297,N_9020,N_8283);
nor U12298 (N_12298,N_8034,N_6405);
and U12299 (N_12299,N_6462,N_7538);
nor U12300 (N_12300,N_8369,N_5968);
nand U12301 (N_12301,N_7566,N_6251);
nand U12302 (N_12302,N_7887,N_9371);
or U12303 (N_12303,N_8692,N_9637);
nor U12304 (N_12304,N_6245,N_7094);
or U12305 (N_12305,N_7241,N_9841);
nor U12306 (N_12306,N_7807,N_7596);
nand U12307 (N_12307,N_5014,N_7743);
and U12308 (N_12308,N_7004,N_9046);
and U12309 (N_12309,N_8906,N_7357);
or U12310 (N_12310,N_6489,N_6599);
nor U12311 (N_12311,N_5985,N_5485);
and U12312 (N_12312,N_9176,N_7413);
nor U12313 (N_12313,N_6233,N_5064);
and U12314 (N_12314,N_8527,N_6676);
nand U12315 (N_12315,N_9168,N_9349);
and U12316 (N_12316,N_5857,N_8219);
and U12317 (N_12317,N_8104,N_6057);
or U12318 (N_12318,N_8727,N_9063);
nand U12319 (N_12319,N_9111,N_7402);
nor U12320 (N_12320,N_8273,N_9443);
and U12321 (N_12321,N_7173,N_8924);
and U12322 (N_12322,N_5306,N_7159);
and U12323 (N_12323,N_7472,N_6724);
nand U12324 (N_12324,N_9127,N_5870);
and U12325 (N_12325,N_6963,N_7296);
nor U12326 (N_12326,N_7103,N_6823);
nor U12327 (N_12327,N_8332,N_9731);
or U12328 (N_12328,N_5604,N_6581);
nand U12329 (N_12329,N_8060,N_8363);
nor U12330 (N_12330,N_8705,N_7289);
or U12331 (N_12331,N_9565,N_9748);
or U12332 (N_12332,N_6956,N_7262);
or U12333 (N_12333,N_6982,N_7356);
or U12334 (N_12334,N_7844,N_6648);
nor U12335 (N_12335,N_8056,N_5859);
nand U12336 (N_12336,N_8063,N_7732);
nor U12337 (N_12337,N_5614,N_6990);
nor U12338 (N_12338,N_6563,N_8617);
and U12339 (N_12339,N_8649,N_8476);
nor U12340 (N_12340,N_9954,N_8096);
nor U12341 (N_12341,N_5657,N_9432);
nor U12342 (N_12342,N_6748,N_8411);
nor U12343 (N_12343,N_8531,N_8820);
nand U12344 (N_12344,N_5301,N_5530);
nand U12345 (N_12345,N_9031,N_8460);
nor U12346 (N_12346,N_7784,N_9568);
nand U12347 (N_12347,N_6323,N_8559);
and U12348 (N_12348,N_6646,N_9080);
nor U12349 (N_12349,N_8420,N_5499);
and U12350 (N_12350,N_7521,N_7256);
and U12351 (N_12351,N_6359,N_8667);
or U12352 (N_12352,N_5852,N_5508);
or U12353 (N_12353,N_9898,N_9186);
and U12354 (N_12354,N_7564,N_5390);
or U12355 (N_12355,N_9519,N_6975);
nand U12356 (N_12356,N_6973,N_8561);
nor U12357 (N_12357,N_9042,N_5264);
and U12358 (N_12358,N_7186,N_8458);
or U12359 (N_12359,N_9124,N_8652);
nand U12360 (N_12360,N_7710,N_9720);
nor U12361 (N_12361,N_7404,N_5023);
nand U12362 (N_12362,N_7177,N_8098);
and U12363 (N_12363,N_8566,N_6942);
nand U12364 (N_12364,N_7089,N_9172);
or U12365 (N_12365,N_6358,N_9222);
and U12366 (N_12366,N_7509,N_8014);
nor U12367 (N_12367,N_9987,N_9614);
or U12368 (N_12368,N_6020,N_8253);
nand U12369 (N_12369,N_8918,N_6992);
or U12370 (N_12370,N_8732,N_5736);
or U12371 (N_12371,N_6756,N_6193);
or U12372 (N_12372,N_8512,N_8677);
and U12373 (N_12373,N_7082,N_9464);
nor U12374 (N_12374,N_7971,N_7575);
or U12375 (N_12375,N_7993,N_9122);
and U12376 (N_12376,N_8716,N_6666);
nand U12377 (N_12377,N_7997,N_5109);
nor U12378 (N_12378,N_8103,N_6870);
or U12379 (N_12379,N_7030,N_7219);
or U12380 (N_12380,N_7750,N_8200);
nor U12381 (N_12381,N_7023,N_9784);
nand U12382 (N_12382,N_9162,N_6491);
nor U12383 (N_12383,N_6824,N_9217);
xnor U12384 (N_12384,N_8269,N_8520);
and U12385 (N_12385,N_6053,N_7686);
and U12386 (N_12386,N_5932,N_5122);
and U12387 (N_12387,N_8085,N_7614);
nand U12388 (N_12388,N_6739,N_9493);
or U12389 (N_12389,N_7859,N_8550);
nor U12390 (N_12390,N_5085,N_8236);
and U12391 (N_12391,N_9970,N_6523);
nand U12392 (N_12392,N_8552,N_9634);
xor U12393 (N_12393,N_8437,N_9887);
nor U12394 (N_12394,N_5435,N_6755);
nand U12395 (N_12395,N_6946,N_9839);
or U12396 (N_12396,N_6347,N_5437);
and U12397 (N_12397,N_5960,N_6328);
and U12398 (N_12398,N_7328,N_9889);
xor U12399 (N_12399,N_8847,N_5332);
nand U12400 (N_12400,N_9073,N_7770);
nand U12401 (N_12401,N_5967,N_5768);
or U12402 (N_12402,N_7441,N_7791);
nand U12403 (N_12403,N_9897,N_6528);
nor U12404 (N_12404,N_8003,N_7647);
nand U12405 (N_12405,N_5166,N_6540);
and U12406 (N_12406,N_9632,N_5860);
and U12407 (N_12407,N_9054,N_8418);
nor U12408 (N_12408,N_5589,N_8026);
or U12409 (N_12409,N_7768,N_7266);
nor U12410 (N_12410,N_8207,N_8549);
nor U12411 (N_12411,N_6872,N_8653);
or U12412 (N_12412,N_7300,N_7530);
nand U12413 (N_12413,N_8666,N_5052);
nor U12414 (N_12414,N_9830,N_8114);
or U12415 (N_12415,N_8882,N_5276);
xnor U12416 (N_12416,N_9863,N_9526);
nand U12417 (N_12417,N_6115,N_9985);
nand U12418 (N_12418,N_7982,N_7522);
or U12419 (N_12419,N_7074,N_8645);
or U12420 (N_12420,N_8121,N_6938);
or U12421 (N_12421,N_5186,N_7450);
or U12422 (N_12422,N_6095,N_6168);
nand U12423 (N_12423,N_9093,N_5199);
or U12424 (N_12424,N_5886,N_8623);
or U12425 (N_12425,N_6084,N_6889);
or U12426 (N_12426,N_5245,N_5759);
nand U12427 (N_12427,N_9152,N_6325);
and U12428 (N_12428,N_9056,N_7720);
nand U12429 (N_12429,N_6317,N_7917);
and U12430 (N_12430,N_9626,N_5277);
or U12431 (N_12431,N_7326,N_5700);
nand U12432 (N_12432,N_7569,N_7294);
and U12433 (N_12433,N_6939,N_5495);
nand U12434 (N_12434,N_8613,N_9910);
nor U12435 (N_12435,N_9380,N_7069);
or U12436 (N_12436,N_5943,N_8941);
nand U12437 (N_12437,N_7948,N_8248);
nand U12438 (N_12438,N_6430,N_8139);
xor U12439 (N_12439,N_5104,N_6891);
and U12440 (N_12440,N_8976,N_7437);
or U12441 (N_12441,N_7060,N_8451);
nand U12442 (N_12442,N_6954,N_6853);
nand U12443 (N_12443,N_9943,N_7912);
nor U12444 (N_12444,N_6122,N_6543);
or U12445 (N_12445,N_7540,N_6046);
nor U12446 (N_12446,N_6820,N_7833);
or U12447 (N_12447,N_6368,N_8016);
nand U12448 (N_12448,N_9064,N_9494);
or U12449 (N_12449,N_7059,N_9107);
nor U12450 (N_12450,N_9756,N_9971);
xor U12451 (N_12451,N_8390,N_5084);
and U12452 (N_12452,N_7009,N_5756);
nor U12453 (N_12453,N_5394,N_5193);
and U12454 (N_12454,N_6730,N_9436);
and U12455 (N_12455,N_5649,N_6849);
or U12456 (N_12456,N_5806,N_9914);
xor U12457 (N_12457,N_6614,N_9455);
nand U12458 (N_12458,N_7215,N_8455);
and U12459 (N_12459,N_6252,N_7135);
nand U12460 (N_12460,N_6915,N_7151);
nor U12461 (N_12461,N_7311,N_6027);
nor U12462 (N_12462,N_8643,N_8917);
or U12463 (N_12463,N_7819,N_9880);
or U12464 (N_12464,N_9964,N_7155);
and U12465 (N_12465,N_8233,N_9041);
and U12466 (N_12466,N_6482,N_7517);
nand U12467 (N_12467,N_8710,N_6712);
nand U12468 (N_12468,N_5323,N_8049);
or U12469 (N_12469,N_9341,N_7394);
and U12470 (N_12470,N_9912,N_9029);
nand U12471 (N_12471,N_8450,N_7980);
nor U12472 (N_12472,N_5720,N_8678);
and U12473 (N_12473,N_8648,N_7761);
and U12474 (N_12474,N_7795,N_5617);
or U12475 (N_12475,N_6099,N_8938);
nor U12476 (N_12476,N_5169,N_9723);
nor U12477 (N_12477,N_6157,N_8497);
and U12478 (N_12478,N_8141,N_9017);
nor U12479 (N_12479,N_8113,N_5563);
or U12480 (N_12480,N_7475,N_8709);
or U12481 (N_12481,N_8965,N_9465);
and U12482 (N_12482,N_8157,N_7255);
and U12483 (N_12483,N_7286,N_8728);
or U12484 (N_12484,N_9660,N_5559);
nand U12485 (N_12485,N_7144,N_5209);
and U12486 (N_12486,N_9725,N_5709);
nor U12487 (N_12487,N_9445,N_9829);
or U12488 (N_12488,N_9576,N_8875);
nand U12489 (N_12489,N_7662,N_9496);
nor U12490 (N_12490,N_7799,N_8804);
nor U12491 (N_12491,N_9420,N_6255);
nand U12492 (N_12492,N_5037,N_8933);
nor U12493 (N_12493,N_6667,N_9773);
or U12494 (N_12494,N_9553,N_9216);
nand U12495 (N_12495,N_5439,N_9001);
or U12496 (N_12496,N_5728,N_5898);
nand U12497 (N_12497,N_6983,N_6785);
nor U12498 (N_12498,N_6114,N_8012);
nor U12499 (N_12499,N_8743,N_6208);
and U12500 (N_12500,N_7045,N_8134);
and U12501 (N_12501,N_7188,N_7373);
nor U12502 (N_12502,N_8238,N_5987);
nand U12503 (N_12503,N_9913,N_7023);
and U12504 (N_12504,N_7661,N_5265);
nor U12505 (N_12505,N_7246,N_7252);
nor U12506 (N_12506,N_8572,N_7421);
nor U12507 (N_12507,N_7587,N_9783);
nor U12508 (N_12508,N_6595,N_6180);
nor U12509 (N_12509,N_6455,N_5698);
and U12510 (N_12510,N_7464,N_7552);
and U12511 (N_12511,N_9494,N_9397);
or U12512 (N_12512,N_5224,N_8864);
nand U12513 (N_12513,N_6900,N_8404);
or U12514 (N_12514,N_9326,N_5774);
xor U12515 (N_12515,N_7665,N_7015);
nor U12516 (N_12516,N_9411,N_5877);
nor U12517 (N_12517,N_5125,N_6602);
and U12518 (N_12518,N_9812,N_6808);
nor U12519 (N_12519,N_9513,N_5792);
and U12520 (N_12520,N_8580,N_8832);
nand U12521 (N_12521,N_6558,N_9253);
nor U12522 (N_12522,N_6860,N_7076);
xor U12523 (N_12523,N_5628,N_9257);
and U12524 (N_12524,N_8272,N_6203);
or U12525 (N_12525,N_8930,N_5461);
nand U12526 (N_12526,N_5693,N_7221);
and U12527 (N_12527,N_5105,N_7356);
nor U12528 (N_12528,N_6367,N_8677);
nor U12529 (N_12529,N_5216,N_6889);
nor U12530 (N_12530,N_8558,N_5887);
xnor U12531 (N_12531,N_5479,N_9443);
nor U12532 (N_12532,N_6928,N_8078);
and U12533 (N_12533,N_5252,N_8346);
and U12534 (N_12534,N_6084,N_7960);
or U12535 (N_12535,N_9477,N_8158);
and U12536 (N_12536,N_8816,N_9216);
and U12537 (N_12537,N_7630,N_9818);
nor U12538 (N_12538,N_8764,N_7382);
xnor U12539 (N_12539,N_8799,N_7541);
and U12540 (N_12540,N_5572,N_8578);
nor U12541 (N_12541,N_7289,N_7793);
nand U12542 (N_12542,N_5514,N_9664);
nor U12543 (N_12543,N_9877,N_6796);
and U12544 (N_12544,N_8812,N_7077);
and U12545 (N_12545,N_8095,N_9954);
nand U12546 (N_12546,N_9593,N_9633);
and U12547 (N_12547,N_7408,N_7664);
xor U12548 (N_12548,N_7632,N_8714);
nor U12549 (N_12549,N_6282,N_9676);
or U12550 (N_12550,N_9904,N_8968);
nand U12551 (N_12551,N_5978,N_7162);
or U12552 (N_12552,N_5373,N_5681);
nand U12553 (N_12553,N_7210,N_9300);
nor U12554 (N_12554,N_7515,N_7144);
xor U12555 (N_12555,N_9061,N_9077);
or U12556 (N_12556,N_8259,N_5545);
nor U12557 (N_12557,N_7863,N_9958);
xnor U12558 (N_12558,N_8257,N_8108);
and U12559 (N_12559,N_9830,N_9128);
or U12560 (N_12560,N_5359,N_6153);
xnor U12561 (N_12561,N_5298,N_6138);
nor U12562 (N_12562,N_7967,N_6033);
and U12563 (N_12563,N_5985,N_8999);
nor U12564 (N_12564,N_8178,N_7837);
nand U12565 (N_12565,N_9133,N_6538);
and U12566 (N_12566,N_9543,N_5541);
nand U12567 (N_12567,N_8141,N_8771);
and U12568 (N_12568,N_9622,N_7653);
nand U12569 (N_12569,N_5857,N_8761);
xor U12570 (N_12570,N_6872,N_8499);
or U12571 (N_12571,N_9285,N_6273);
nor U12572 (N_12572,N_9891,N_6182);
xor U12573 (N_12573,N_6316,N_7192);
nand U12574 (N_12574,N_7170,N_6304);
or U12575 (N_12575,N_7463,N_9240);
and U12576 (N_12576,N_6477,N_9654);
nor U12577 (N_12577,N_9465,N_8092);
nor U12578 (N_12578,N_7901,N_7594);
and U12579 (N_12579,N_5773,N_9848);
and U12580 (N_12580,N_6582,N_5632);
xor U12581 (N_12581,N_7642,N_8913);
or U12582 (N_12582,N_7698,N_7471);
nor U12583 (N_12583,N_6931,N_8747);
or U12584 (N_12584,N_9408,N_6484);
nand U12585 (N_12585,N_8173,N_7987);
nand U12586 (N_12586,N_5337,N_8855);
or U12587 (N_12587,N_8017,N_9360);
nor U12588 (N_12588,N_8773,N_9997);
and U12589 (N_12589,N_8349,N_9813);
or U12590 (N_12590,N_7486,N_6119);
and U12591 (N_12591,N_7241,N_9130);
nor U12592 (N_12592,N_5458,N_5542);
nand U12593 (N_12593,N_7852,N_5461);
or U12594 (N_12594,N_6829,N_9024);
nor U12595 (N_12595,N_6839,N_8542);
or U12596 (N_12596,N_8060,N_5174);
nor U12597 (N_12597,N_9660,N_5661);
xor U12598 (N_12598,N_7859,N_6551);
and U12599 (N_12599,N_9858,N_7114);
or U12600 (N_12600,N_8919,N_7043);
nand U12601 (N_12601,N_5685,N_6133);
nand U12602 (N_12602,N_7572,N_7231);
nand U12603 (N_12603,N_7560,N_5508);
nand U12604 (N_12604,N_6281,N_8369);
nand U12605 (N_12605,N_6340,N_5982);
nand U12606 (N_12606,N_5962,N_6017);
and U12607 (N_12607,N_9200,N_6926);
and U12608 (N_12608,N_6833,N_5692);
or U12609 (N_12609,N_9892,N_6627);
and U12610 (N_12610,N_8437,N_9723);
or U12611 (N_12611,N_6384,N_9520);
nand U12612 (N_12612,N_7403,N_9862);
nor U12613 (N_12613,N_6770,N_8469);
and U12614 (N_12614,N_6666,N_9652);
or U12615 (N_12615,N_5754,N_7149);
or U12616 (N_12616,N_7088,N_6796);
nand U12617 (N_12617,N_6840,N_7930);
nand U12618 (N_12618,N_5411,N_9506);
and U12619 (N_12619,N_6216,N_9730);
or U12620 (N_12620,N_9320,N_7242);
nor U12621 (N_12621,N_9277,N_8995);
or U12622 (N_12622,N_9956,N_6627);
nor U12623 (N_12623,N_8678,N_5004);
and U12624 (N_12624,N_9630,N_5158);
nand U12625 (N_12625,N_9247,N_7533);
or U12626 (N_12626,N_8821,N_7296);
nand U12627 (N_12627,N_6833,N_6321);
and U12628 (N_12628,N_7460,N_8536);
nand U12629 (N_12629,N_8274,N_8205);
or U12630 (N_12630,N_8997,N_5201);
nand U12631 (N_12631,N_7317,N_7713);
and U12632 (N_12632,N_7180,N_5337);
nor U12633 (N_12633,N_6142,N_9026);
or U12634 (N_12634,N_7204,N_7932);
or U12635 (N_12635,N_5645,N_8267);
and U12636 (N_12636,N_7450,N_9706);
and U12637 (N_12637,N_7526,N_6238);
and U12638 (N_12638,N_9252,N_6160);
or U12639 (N_12639,N_8123,N_9283);
and U12640 (N_12640,N_8711,N_8544);
and U12641 (N_12641,N_8951,N_8865);
nor U12642 (N_12642,N_7707,N_9107);
nor U12643 (N_12643,N_8768,N_6040);
or U12644 (N_12644,N_7497,N_8179);
or U12645 (N_12645,N_8501,N_5991);
nor U12646 (N_12646,N_5980,N_7875);
or U12647 (N_12647,N_6781,N_7070);
nand U12648 (N_12648,N_6668,N_5826);
or U12649 (N_12649,N_9363,N_7248);
and U12650 (N_12650,N_6923,N_9999);
and U12651 (N_12651,N_6134,N_5579);
nor U12652 (N_12652,N_8255,N_7475);
xor U12653 (N_12653,N_5408,N_6108);
or U12654 (N_12654,N_6860,N_9926);
nor U12655 (N_12655,N_5566,N_8089);
and U12656 (N_12656,N_5356,N_9454);
and U12657 (N_12657,N_6475,N_5689);
nor U12658 (N_12658,N_6930,N_8755);
and U12659 (N_12659,N_9399,N_7404);
and U12660 (N_12660,N_7126,N_8631);
and U12661 (N_12661,N_8938,N_9515);
nand U12662 (N_12662,N_9948,N_6393);
nand U12663 (N_12663,N_6984,N_9861);
and U12664 (N_12664,N_5579,N_5139);
and U12665 (N_12665,N_5465,N_5890);
or U12666 (N_12666,N_9851,N_6164);
and U12667 (N_12667,N_7461,N_9189);
and U12668 (N_12668,N_5234,N_7306);
nand U12669 (N_12669,N_6003,N_5538);
nand U12670 (N_12670,N_7208,N_9706);
and U12671 (N_12671,N_8052,N_5223);
or U12672 (N_12672,N_7373,N_8313);
nor U12673 (N_12673,N_5846,N_8520);
nand U12674 (N_12674,N_8809,N_5028);
nor U12675 (N_12675,N_8026,N_7080);
nand U12676 (N_12676,N_9690,N_6562);
and U12677 (N_12677,N_6387,N_6313);
nand U12678 (N_12678,N_5712,N_6466);
and U12679 (N_12679,N_5863,N_8482);
xor U12680 (N_12680,N_9933,N_5807);
or U12681 (N_12681,N_7075,N_5119);
nor U12682 (N_12682,N_8433,N_9010);
nand U12683 (N_12683,N_9592,N_8633);
nor U12684 (N_12684,N_8597,N_8358);
or U12685 (N_12685,N_8138,N_5549);
or U12686 (N_12686,N_5583,N_9902);
xor U12687 (N_12687,N_8593,N_8969);
nand U12688 (N_12688,N_7468,N_7026);
xor U12689 (N_12689,N_8766,N_6258);
or U12690 (N_12690,N_5423,N_9913);
and U12691 (N_12691,N_6122,N_9316);
or U12692 (N_12692,N_8463,N_5473);
and U12693 (N_12693,N_7544,N_5679);
or U12694 (N_12694,N_7590,N_8604);
nor U12695 (N_12695,N_8795,N_9260);
nand U12696 (N_12696,N_8741,N_5027);
nand U12697 (N_12697,N_7357,N_8324);
or U12698 (N_12698,N_5514,N_9519);
and U12699 (N_12699,N_6579,N_6970);
and U12700 (N_12700,N_9722,N_6875);
or U12701 (N_12701,N_9834,N_8706);
or U12702 (N_12702,N_6637,N_5021);
and U12703 (N_12703,N_6957,N_8493);
nor U12704 (N_12704,N_8560,N_8173);
nor U12705 (N_12705,N_9312,N_6385);
or U12706 (N_12706,N_8563,N_8423);
or U12707 (N_12707,N_7158,N_8419);
nand U12708 (N_12708,N_9437,N_9557);
or U12709 (N_12709,N_6279,N_6684);
xor U12710 (N_12710,N_7546,N_9894);
nand U12711 (N_12711,N_8738,N_6283);
or U12712 (N_12712,N_5297,N_5043);
nand U12713 (N_12713,N_9476,N_5808);
nor U12714 (N_12714,N_7308,N_6599);
and U12715 (N_12715,N_7985,N_6404);
nor U12716 (N_12716,N_5712,N_6197);
nor U12717 (N_12717,N_8871,N_9364);
nand U12718 (N_12718,N_9656,N_8643);
and U12719 (N_12719,N_9594,N_7989);
nor U12720 (N_12720,N_6842,N_5240);
nor U12721 (N_12721,N_6217,N_8152);
or U12722 (N_12722,N_7486,N_6267);
nor U12723 (N_12723,N_9287,N_5711);
nor U12724 (N_12724,N_5674,N_6217);
nor U12725 (N_12725,N_6746,N_5644);
nor U12726 (N_12726,N_6877,N_8144);
nand U12727 (N_12727,N_8284,N_5400);
nand U12728 (N_12728,N_8832,N_7683);
or U12729 (N_12729,N_8140,N_5769);
nor U12730 (N_12730,N_5290,N_5693);
nand U12731 (N_12731,N_9637,N_9951);
nand U12732 (N_12732,N_9345,N_8663);
or U12733 (N_12733,N_9979,N_7566);
nor U12734 (N_12734,N_8847,N_9697);
and U12735 (N_12735,N_7023,N_6314);
nor U12736 (N_12736,N_7760,N_7361);
or U12737 (N_12737,N_6428,N_9016);
nor U12738 (N_12738,N_5925,N_8903);
and U12739 (N_12739,N_8277,N_5004);
or U12740 (N_12740,N_8966,N_8656);
and U12741 (N_12741,N_8640,N_7273);
nand U12742 (N_12742,N_7065,N_6219);
nand U12743 (N_12743,N_9090,N_5209);
nand U12744 (N_12744,N_7921,N_5973);
nand U12745 (N_12745,N_5152,N_8893);
and U12746 (N_12746,N_5371,N_9431);
or U12747 (N_12747,N_7377,N_9189);
and U12748 (N_12748,N_5488,N_7055);
or U12749 (N_12749,N_9700,N_8500);
and U12750 (N_12750,N_9888,N_5338);
nand U12751 (N_12751,N_6261,N_7388);
nor U12752 (N_12752,N_9969,N_6260);
nand U12753 (N_12753,N_5722,N_8054);
and U12754 (N_12754,N_5262,N_8716);
or U12755 (N_12755,N_6134,N_8875);
nor U12756 (N_12756,N_7327,N_7006);
and U12757 (N_12757,N_5870,N_6058);
nand U12758 (N_12758,N_6382,N_6460);
and U12759 (N_12759,N_9604,N_6384);
nor U12760 (N_12760,N_5595,N_8449);
and U12761 (N_12761,N_5007,N_8262);
and U12762 (N_12762,N_8246,N_7276);
nand U12763 (N_12763,N_5392,N_9143);
or U12764 (N_12764,N_8773,N_5434);
nand U12765 (N_12765,N_5651,N_8655);
or U12766 (N_12766,N_5931,N_5033);
or U12767 (N_12767,N_9852,N_6635);
or U12768 (N_12768,N_8173,N_8923);
or U12769 (N_12769,N_7233,N_5049);
nand U12770 (N_12770,N_9800,N_7118);
and U12771 (N_12771,N_8421,N_6351);
nor U12772 (N_12772,N_6467,N_8338);
or U12773 (N_12773,N_7183,N_9353);
and U12774 (N_12774,N_6669,N_9747);
xor U12775 (N_12775,N_9651,N_6241);
or U12776 (N_12776,N_5907,N_9508);
nor U12777 (N_12777,N_5036,N_7487);
xor U12778 (N_12778,N_5227,N_6540);
nor U12779 (N_12779,N_9426,N_6766);
nand U12780 (N_12780,N_6567,N_5679);
and U12781 (N_12781,N_9433,N_7403);
or U12782 (N_12782,N_8858,N_7705);
or U12783 (N_12783,N_7357,N_6375);
nor U12784 (N_12784,N_6196,N_7508);
nor U12785 (N_12785,N_9209,N_6568);
and U12786 (N_12786,N_6345,N_8056);
and U12787 (N_12787,N_5055,N_5081);
or U12788 (N_12788,N_5588,N_8522);
nor U12789 (N_12789,N_7814,N_9601);
or U12790 (N_12790,N_8772,N_7810);
nand U12791 (N_12791,N_5281,N_6258);
or U12792 (N_12792,N_9138,N_8763);
and U12793 (N_12793,N_8589,N_6842);
or U12794 (N_12794,N_9343,N_7855);
and U12795 (N_12795,N_8604,N_7958);
nand U12796 (N_12796,N_6969,N_5451);
nor U12797 (N_12797,N_8153,N_9278);
or U12798 (N_12798,N_8554,N_5635);
nor U12799 (N_12799,N_9109,N_6719);
and U12800 (N_12800,N_9482,N_8483);
and U12801 (N_12801,N_5179,N_7183);
nand U12802 (N_12802,N_8129,N_9748);
nor U12803 (N_12803,N_9561,N_7349);
xor U12804 (N_12804,N_7149,N_9511);
nor U12805 (N_12805,N_5820,N_7101);
nor U12806 (N_12806,N_9528,N_7222);
nor U12807 (N_12807,N_6658,N_8241);
and U12808 (N_12808,N_8967,N_7840);
nand U12809 (N_12809,N_9636,N_9589);
nand U12810 (N_12810,N_9576,N_5392);
nor U12811 (N_12811,N_8497,N_8950);
or U12812 (N_12812,N_5429,N_6662);
or U12813 (N_12813,N_7911,N_6903);
nor U12814 (N_12814,N_7112,N_8601);
and U12815 (N_12815,N_5723,N_7369);
and U12816 (N_12816,N_5387,N_6119);
nor U12817 (N_12817,N_6894,N_9723);
nand U12818 (N_12818,N_9926,N_7049);
and U12819 (N_12819,N_9428,N_6178);
and U12820 (N_12820,N_8479,N_5837);
nand U12821 (N_12821,N_9017,N_9185);
nand U12822 (N_12822,N_7472,N_5749);
nor U12823 (N_12823,N_7514,N_7902);
xor U12824 (N_12824,N_6348,N_7476);
nor U12825 (N_12825,N_5771,N_9807);
nand U12826 (N_12826,N_8080,N_6590);
nand U12827 (N_12827,N_9004,N_6229);
and U12828 (N_12828,N_6076,N_8458);
nand U12829 (N_12829,N_5626,N_5841);
nor U12830 (N_12830,N_8721,N_9800);
nand U12831 (N_12831,N_7025,N_6289);
or U12832 (N_12832,N_6656,N_9254);
and U12833 (N_12833,N_9900,N_8415);
or U12834 (N_12834,N_8513,N_8575);
nand U12835 (N_12835,N_7381,N_5020);
and U12836 (N_12836,N_9440,N_9339);
nor U12837 (N_12837,N_8829,N_6208);
nand U12838 (N_12838,N_7320,N_8895);
and U12839 (N_12839,N_6577,N_6543);
nor U12840 (N_12840,N_5369,N_8541);
and U12841 (N_12841,N_7846,N_6961);
nand U12842 (N_12842,N_9669,N_9918);
nand U12843 (N_12843,N_9476,N_7657);
or U12844 (N_12844,N_9802,N_5700);
xnor U12845 (N_12845,N_8577,N_8580);
or U12846 (N_12846,N_6461,N_6783);
or U12847 (N_12847,N_7144,N_7931);
or U12848 (N_12848,N_5253,N_9233);
or U12849 (N_12849,N_9761,N_9092);
and U12850 (N_12850,N_6474,N_6873);
and U12851 (N_12851,N_6603,N_6060);
or U12852 (N_12852,N_6127,N_7347);
nor U12853 (N_12853,N_7041,N_5347);
xnor U12854 (N_12854,N_7333,N_8378);
or U12855 (N_12855,N_5149,N_6133);
nand U12856 (N_12856,N_5429,N_6550);
and U12857 (N_12857,N_9924,N_5373);
or U12858 (N_12858,N_6630,N_6461);
and U12859 (N_12859,N_5247,N_8281);
or U12860 (N_12860,N_8269,N_6527);
or U12861 (N_12861,N_8151,N_7327);
nand U12862 (N_12862,N_9062,N_9762);
and U12863 (N_12863,N_8961,N_6819);
nand U12864 (N_12864,N_9487,N_5342);
or U12865 (N_12865,N_8555,N_5980);
nand U12866 (N_12866,N_7194,N_7132);
nor U12867 (N_12867,N_8603,N_7167);
nand U12868 (N_12868,N_6310,N_7844);
nand U12869 (N_12869,N_9095,N_9285);
nor U12870 (N_12870,N_9868,N_9755);
nand U12871 (N_12871,N_8598,N_6807);
or U12872 (N_12872,N_9163,N_6502);
nor U12873 (N_12873,N_8665,N_5137);
or U12874 (N_12874,N_8140,N_7697);
nor U12875 (N_12875,N_5449,N_5732);
and U12876 (N_12876,N_8164,N_9754);
or U12877 (N_12877,N_8778,N_9274);
or U12878 (N_12878,N_5129,N_5685);
and U12879 (N_12879,N_9117,N_5029);
or U12880 (N_12880,N_8025,N_9752);
and U12881 (N_12881,N_5615,N_9708);
or U12882 (N_12882,N_6459,N_9358);
nand U12883 (N_12883,N_8327,N_5843);
and U12884 (N_12884,N_6938,N_8108);
and U12885 (N_12885,N_6016,N_9795);
nand U12886 (N_12886,N_7647,N_9524);
nor U12887 (N_12887,N_9530,N_6054);
nand U12888 (N_12888,N_9405,N_9658);
or U12889 (N_12889,N_9839,N_8368);
and U12890 (N_12890,N_9839,N_8159);
nor U12891 (N_12891,N_9262,N_8037);
or U12892 (N_12892,N_5046,N_8747);
nand U12893 (N_12893,N_6381,N_7960);
nor U12894 (N_12894,N_9620,N_6756);
or U12895 (N_12895,N_9139,N_5800);
and U12896 (N_12896,N_6288,N_9423);
or U12897 (N_12897,N_5466,N_6571);
nand U12898 (N_12898,N_5521,N_8769);
or U12899 (N_12899,N_8178,N_6227);
and U12900 (N_12900,N_5435,N_8942);
nor U12901 (N_12901,N_6490,N_7387);
and U12902 (N_12902,N_5553,N_7862);
and U12903 (N_12903,N_6200,N_8683);
nor U12904 (N_12904,N_7623,N_5390);
nor U12905 (N_12905,N_7363,N_8587);
and U12906 (N_12906,N_9067,N_5262);
and U12907 (N_12907,N_5898,N_8057);
or U12908 (N_12908,N_9990,N_7088);
or U12909 (N_12909,N_9264,N_6398);
and U12910 (N_12910,N_9612,N_5912);
or U12911 (N_12911,N_8902,N_9640);
or U12912 (N_12912,N_8259,N_9305);
nand U12913 (N_12913,N_6861,N_7103);
nand U12914 (N_12914,N_8135,N_6543);
nand U12915 (N_12915,N_5835,N_7003);
and U12916 (N_12916,N_7848,N_8524);
or U12917 (N_12917,N_9320,N_6562);
nand U12918 (N_12918,N_7652,N_8788);
nor U12919 (N_12919,N_9651,N_5086);
or U12920 (N_12920,N_5983,N_8883);
nor U12921 (N_12921,N_9442,N_8017);
and U12922 (N_12922,N_6769,N_8921);
and U12923 (N_12923,N_5072,N_8097);
nor U12924 (N_12924,N_8554,N_5434);
nor U12925 (N_12925,N_6429,N_7800);
or U12926 (N_12926,N_7519,N_8782);
nor U12927 (N_12927,N_5912,N_8545);
nand U12928 (N_12928,N_8145,N_7394);
or U12929 (N_12929,N_6208,N_5552);
or U12930 (N_12930,N_8288,N_6988);
or U12931 (N_12931,N_7406,N_8607);
nand U12932 (N_12932,N_7861,N_8686);
and U12933 (N_12933,N_9480,N_8662);
nand U12934 (N_12934,N_5216,N_7269);
and U12935 (N_12935,N_5549,N_6920);
nor U12936 (N_12936,N_5362,N_8316);
and U12937 (N_12937,N_8627,N_5158);
nand U12938 (N_12938,N_9891,N_9698);
nand U12939 (N_12939,N_5543,N_9788);
nor U12940 (N_12940,N_6375,N_9841);
nor U12941 (N_12941,N_6647,N_8364);
nand U12942 (N_12942,N_7854,N_6984);
and U12943 (N_12943,N_5647,N_5609);
or U12944 (N_12944,N_8700,N_5117);
nand U12945 (N_12945,N_8513,N_6568);
nor U12946 (N_12946,N_7609,N_9470);
and U12947 (N_12947,N_6679,N_9393);
or U12948 (N_12948,N_8526,N_5548);
or U12949 (N_12949,N_9722,N_7228);
and U12950 (N_12950,N_6688,N_7240);
nand U12951 (N_12951,N_7657,N_5749);
nor U12952 (N_12952,N_5519,N_9792);
nand U12953 (N_12953,N_7838,N_8937);
and U12954 (N_12954,N_5152,N_8849);
or U12955 (N_12955,N_7018,N_5919);
nor U12956 (N_12956,N_7478,N_8600);
and U12957 (N_12957,N_6504,N_8721);
or U12958 (N_12958,N_5887,N_7970);
nor U12959 (N_12959,N_9758,N_5493);
nand U12960 (N_12960,N_6377,N_9868);
or U12961 (N_12961,N_8075,N_5944);
nand U12962 (N_12962,N_9199,N_5262);
or U12963 (N_12963,N_9797,N_7872);
nand U12964 (N_12964,N_9759,N_9227);
nor U12965 (N_12965,N_6400,N_8612);
or U12966 (N_12966,N_7732,N_6916);
nor U12967 (N_12967,N_5800,N_8792);
or U12968 (N_12968,N_5552,N_8417);
nand U12969 (N_12969,N_5546,N_7072);
nor U12970 (N_12970,N_5557,N_7477);
or U12971 (N_12971,N_7505,N_9226);
nand U12972 (N_12972,N_9711,N_9218);
or U12973 (N_12973,N_6026,N_9701);
nand U12974 (N_12974,N_9702,N_7305);
nand U12975 (N_12975,N_7362,N_6875);
nand U12976 (N_12976,N_8077,N_7927);
nand U12977 (N_12977,N_8936,N_6088);
nand U12978 (N_12978,N_5121,N_5265);
nand U12979 (N_12979,N_9498,N_5380);
and U12980 (N_12980,N_7293,N_8873);
nor U12981 (N_12981,N_6143,N_5226);
or U12982 (N_12982,N_5523,N_5847);
or U12983 (N_12983,N_9022,N_7566);
or U12984 (N_12984,N_9727,N_8875);
nor U12985 (N_12985,N_9173,N_8978);
and U12986 (N_12986,N_5675,N_9071);
and U12987 (N_12987,N_8003,N_5167);
or U12988 (N_12988,N_7359,N_5769);
and U12989 (N_12989,N_5030,N_9353);
nor U12990 (N_12990,N_8671,N_9233);
and U12991 (N_12991,N_5033,N_5437);
and U12992 (N_12992,N_8979,N_7314);
and U12993 (N_12993,N_6449,N_7396);
nor U12994 (N_12994,N_6715,N_8770);
xor U12995 (N_12995,N_6020,N_9073);
nand U12996 (N_12996,N_9330,N_5109);
or U12997 (N_12997,N_8873,N_8022);
nor U12998 (N_12998,N_5403,N_7151);
nor U12999 (N_12999,N_9057,N_9394);
or U13000 (N_13000,N_7104,N_9356);
or U13001 (N_13001,N_8958,N_8725);
nand U13002 (N_13002,N_6378,N_5150);
and U13003 (N_13003,N_9414,N_5203);
nand U13004 (N_13004,N_6861,N_6908);
and U13005 (N_13005,N_5842,N_8155);
nand U13006 (N_13006,N_8722,N_5592);
nor U13007 (N_13007,N_6718,N_7135);
and U13008 (N_13008,N_5375,N_9890);
nand U13009 (N_13009,N_7838,N_9420);
nand U13010 (N_13010,N_9034,N_5800);
and U13011 (N_13011,N_6169,N_8282);
nand U13012 (N_13012,N_9922,N_8011);
nor U13013 (N_13013,N_5821,N_7465);
or U13014 (N_13014,N_8215,N_7061);
nor U13015 (N_13015,N_6183,N_9435);
and U13016 (N_13016,N_5729,N_6151);
or U13017 (N_13017,N_5892,N_5246);
nand U13018 (N_13018,N_9938,N_9273);
or U13019 (N_13019,N_8071,N_8562);
nor U13020 (N_13020,N_9544,N_7623);
nor U13021 (N_13021,N_7427,N_9123);
nor U13022 (N_13022,N_7514,N_7892);
nor U13023 (N_13023,N_5018,N_7978);
nor U13024 (N_13024,N_8299,N_5288);
nand U13025 (N_13025,N_9733,N_6340);
or U13026 (N_13026,N_7136,N_9035);
or U13027 (N_13027,N_9702,N_9764);
nor U13028 (N_13028,N_7442,N_6504);
nand U13029 (N_13029,N_9653,N_6844);
nor U13030 (N_13030,N_8344,N_8916);
and U13031 (N_13031,N_7620,N_8494);
or U13032 (N_13032,N_9789,N_8533);
nor U13033 (N_13033,N_6716,N_8433);
and U13034 (N_13034,N_6550,N_8199);
and U13035 (N_13035,N_8593,N_9844);
or U13036 (N_13036,N_7169,N_8047);
and U13037 (N_13037,N_9316,N_8832);
and U13038 (N_13038,N_8323,N_8763);
or U13039 (N_13039,N_6206,N_8268);
nand U13040 (N_13040,N_6257,N_7725);
nand U13041 (N_13041,N_9146,N_8283);
nand U13042 (N_13042,N_5161,N_5029);
and U13043 (N_13043,N_5624,N_6765);
and U13044 (N_13044,N_5294,N_8389);
nor U13045 (N_13045,N_7807,N_8937);
or U13046 (N_13046,N_5915,N_8176);
nand U13047 (N_13047,N_9961,N_5000);
nor U13048 (N_13048,N_6577,N_9562);
nand U13049 (N_13049,N_7437,N_6223);
xor U13050 (N_13050,N_9377,N_5099);
or U13051 (N_13051,N_7448,N_5882);
nor U13052 (N_13052,N_7671,N_6935);
or U13053 (N_13053,N_5213,N_5852);
and U13054 (N_13054,N_9553,N_8464);
or U13055 (N_13055,N_5227,N_9962);
or U13056 (N_13056,N_7837,N_8491);
and U13057 (N_13057,N_7820,N_5594);
and U13058 (N_13058,N_8485,N_5082);
and U13059 (N_13059,N_8903,N_8521);
nor U13060 (N_13060,N_7661,N_7997);
nor U13061 (N_13061,N_5666,N_8454);
xnor U13062 (N_13062,N_8889,N_6145);
and U13063 (N_13063,N_6382,N_6739);
nand U13064 (N_13064,N_5540,N_8550);
nand U13065 (N_13065,N_9509,N_7618);
or U13066 (N_13066,N_7238,N_5330);
or U13067 (N_13067,N_8681,N_8085);
or U13068 (N_13068,N_9010,N_8407);
and U13069 (N_13069,N_6081,N_6920);
xor U13070 (N_13070,N_7052,N_9388);
and U13071 (N_13071,N_6581,N_5906);
nand U13072 (N_13072,N_8181,N_6956);
or U13073 (N_13073,N_7873,N_8131);
nor U13074 (N_13074,N_7016,N_9557);
xor U13075 (N_13075,N_6710,N_7283);
nand U13076 (N_13076,N_9870,N_5969);
nor U13077 (N_13077,N_5698,N_6586);
or U13078 (N_13078,N_5562,N_6105);
nor U13079 (N_13079,N_6399,N_7571);
nor U13080 (N_13080,N_9518,N_6999);
and U13081 (N_13081,N_5006,N_7588);
nand U13082 (N_13082,N_7860,N_5143);
nand U13083 (N_13083,N_9965,N_7513);
and U13084 (N_13084,N_9130,N_8925);
xor U13085 (N_13085,N_7272,N_9858);
and U13086 (N_13086,N_9325,N_9246);
and U13087 (N_13087,N_5587,N_6627);
nand U13088 (N_13088,N_7149,N_5677);
or U13089 (N_13089,N_6942,N_6535);
or U13090 (N_13090,N_5351,N_7720);
nor U13091 (N_13091,N_9349,N_5603);
nand U13092 (N_13092,N_7788,N_6801);
or U13093 (N_13093,N_7234,N_8028);
and U13094 (N_13094,N_7462,N_5910);
nor U13095 (N_13095,N_6190,N_9084);
or U13096 (N_13096,N_9881,N_7065);
nor U13097 (N_13097,N_9077,N_7089);
nand U13098 (N_13098,N_8501,N_7089);
and U13099 (N_13099,N_8750,N_5720);
nand U13100 (N_13100,N_6559,N_8038);
nor U13101 (N_13101,N_7753,N_7053);
and U13102 (N_13102,N_5887,N_5737);
nor U13103 (N_13103,N_8866,N_5339);
or U13104 (N_13104,N_8064,N_6510);
nor U13105 (N_13105,N_6880,N_7265);
or U13106 (N_13106,N_9299,N_9818);
nand U13107 (N_13107,N_8872,N_7047);
and U13108 (N_13108,N_9264,N_9655);
nand U13109 (N_13109,N_5788,N_7276);
and U13110 (N_13110,N_5764,N_8990);
nand U13111 (N_13111,N_7497,N_6345);
or U13112 (N_13112,N_8458,N_6280);
nand U13113 (N_13113,N_5407,N_7517);
and U13114 (N_13114,N_7937,N_7935);
nor U13115 (N_13115,N_5201,N_9582);
and U13116 (N_13116,N_5389,N_7565);
xnor U13117 (N_13117,N_8927,N_5141);
or U13118 (N_13118,N_9717,N_6252);
and U13119 (N_13119,N_9461,N_8249);
nand U13120 (N_13120,N_9857,N_6249);
nor U13121 (N_13121,N_7555,N_7647);
nand U13122 (N_13122,N_6485,N_5330);
and U13123 (N_13123,N_5269,N_9709);
and U13124 (N_13124,N_7447,N_8448);
nor U13125 (N_13125,N_8717,N_8865);
nor U13126 (N_13126,N_9012,N_8769);
and U13127 (N_13127,N_7235,N_7317);
nand U13128 (N_13128,N_8699,N_5852);
nand U13129 (N_13129,N_8908,N_6084);
nand U13130 (N_13130,N_6247,N_6447);
or U13131 (N_13131,N_8928,N_7110);
nand U13132 (N_13132,N_5462,N_6708);
or U13133 (N_13133,N_9972,N_6878);
nand U13134 (N_13134,N_5302,N_6405);
nor U13135 (N_13135,N_6060,N_9641);
or U13136 (N_13136,N_9594,N_5270);
nor U13137 (N_13137,N_8821,N_7863);
nor U13138 (N_13138,N_9624,N_9799);
and U13139 (N_13139,N_9026,N_5299);
or U13140 (N_13140,N_8830,N_5692);
nand U13141 (N_13141,N_9372,N_8148);
or U13142 (N_13142,N_5378,N_5943);
and U13143 (N_13143,N_7800,N_9613);
or U13144 (N_13144,N_9091,N_7551);
nand U13145 (N_13145,N_9558,N_8684);
nor U13146 (N_13146,N_9417,N_5765);
nand U13147 (N_13147,N_5976,N_6171);
nor U13148 (N_13148,N_5930,N_9544);
and U13149 (N_13149,N_7295,N_6656);
or U13150 (N_13150,N_5268,N_7109);
nor U13151 (N_13151,N_8636,N_8944);
and U13152 (N_13152,N_9785,N_9210);
nor U13153 (N_13153,N_7355,N_5639);
nand U13154 (N_13154,N_9424,N_8277);
nand U13155 (N_13155,N_9210,N_8341);
or U13156 (N_13156,N_7843,N_7093);
nor U13157 (N_13157,N_9938,N_7363);
nand U13158 (N_13158,N_7402,N_7841);
nor U13159 (N_13159,N_8855,N_9016);
nand U13160 (N_13160,N_5016,N_7200);
nand U13161 (N_13161,N_6437,N_7816);
or U13162 (N_13162,N_5007,N_5488);
or U13163 (N_13163,N_5561,N_7865);
nor U13164 (N_13164,N_8067,N_7810);
and U13165 (N_13165,N_9186,N_5202);
nand U13166 (N_13166,N_8762,N_9003);
nand U13167 (N_13167,N_9558,N_9941);
and U13168 (N_13168,N_5640,N_5347);
nand U13169 (N_13169,N_8917,N_6769);
and U13170 (N_13170,N_5355,N_9722);
nor U13171 (N_13171,N_6502,N_7542);
nor U13172 (N_13172,N_6814,N_8005);
nand U13173 (N_13173,N_5566,N_7681);
nor U13174 (N_13174,N_6937,N_5177);
nand U13175 (N_13175,N_7926,N_9031);
nand U13176 (N_13176,N_9598,N_7512);
nor U13177 (N_13177,N_8716,N_8548);
nor U13178 (N_13178,N_5087,N_6433);
nor U13179 (N_13179,N_8756,N_9853);
and U13180 (N_13180,N_6898,N_9839);
nand U13181 (N_13181,N_8225,N_5919);
nor U13182 (N_13182,N_9004,N_7006);
nand U13183 (N_13183,N_5195,N_6722);
or U13184 (N_13184,N_7288,N_5117);
nand U13185 (N_13185,N_5469,N_6675);
or U13186 (N_13186,N_9404,N_5409);
and U13187 (N_13187,N_5366,N_6475);
or U13188 (N_13188,N_6632,N_6937);
or U13189 (N_13189,N_8971,N_6219);
and U13190 (N_13190,N_9126,N_6745);
or U13191 (N_13191,N_5768,N_7390);
or U13192 (N_13192,N_5505,N_7890);
nand U13193 (N_13193,N_6694,N_6658);
nor U13194 (N_13194,N_9680,N_9453);
and U13195 (N_13195,N_6186,N_8712);
xnor U13196 (N_13196,N_6767,N_9762);
or U13197 (N_13197,N_8218,N_8323);
nand U13198 (N_13198,N_6716,N_5417);
nor U13199 (N_13199,N_7389,N_5579);
and U13200 (N_13200,N_5749,N_6700);
nand U13201 (N_13201,N_9545,N_5851);
nand U13202 (N_13202,N_9909,N_9447);
and U13203 (N_13203,N_6147,N_7029);
nand U13204 (N_13204,N_8589,N_8832);
nor U13205 (N_13205,N_7318,N_9170);
nand U13206 (N_13206,N_5747,N_7876);
and U13207 (N_13207,N_7265,N_9140);
nor U13208 (N_13208,N_5825,N_9942);
or U13209 (N_13209,N_8705,N_8725);
and U13210 (N_13210,N_9988,N_7451);
and U13211 (N_13211,N_9819,N_6745);
nor U13212 (N_13212,N_6635,N_6895);
xnor U13213 (N_13213,N_5376,N_6002);
and U13214 (N_13214,N_8752,N_9765);
nand U13215 (N_13215,N_6991,N_8222);
nor U13216 (N_13216,N_6456,N_8223);
and U13217 (N_13217,N_6717,N_7900);
nor U13218 (N_13218,N_7163,N_6271);
xor U13219 (N_13219,N_9233,N_9345);
nand U13220 (N_13220,N_8741,N_8570);
and U13221 (N_13221,N_7970,N_5348);
or U13222 (N_13222,N_9541,N_7691);
nor U13223 (N_13223,N_9621,N_7257);
nor U13224 (N_13224,N_5331,N_9699);
nand U13225 (N_13225,N_5945,N_5180);
nor U13226 (N_13226,N_6963,N_9764);
xor U13227 (N_13227,N_7560,N_6316);
nor U13228 (N_13228,N_6406,N_9019);
or U13229 (N_13229,N_6861,N_9565);
and U13230 (N_13230,N_6899,N_5970);
nand U13231 (N_13231,N_9267,N_6728);
nor U13232 (N_13232,N_9254,N_6883);
or U13233 (N_13233,N_6806,N_6169);
nand U13234 (N_13234,N_8739,N_8534);
nor U13235 (N_13235,N_9692,N_6963);
nand U13236 (N_13236,N_5354,N_6235);
nand U13237 (N_13237,N_7525,N_9911);
or U13238 (N_13238,N_7987,N_8730);
and U13239 (N_13239,N_8536,N_6483);
nand U13240 (N_13240,N_9009,N_7632);
nor U13241 (N_13241,N_7964,N_7017);
and U13242 (N_13242,N_7205,N_8064);
nand U13243 (N_13243,N_8965,N_8258);
or U13244 (N_13244,N_5280,N_9963);
or U13245 (N_13245,N_8922,N_5304);
or U13246 (N_13246,N_9488,N_9674);
or U13247 (N_13247,N_8706,N_9557);
or U13248 (N_13248,N_8366,N_7679);
and U13249 (N_13249,N_5680,N_5750);
nand U13250 (N_13250,N_6374,N_8300);
nor U13251 (N_13251,N_9081,N_7631);
xor U13252 (N_13252,N_9577,N_8763);
nor U13253 (N_13253,N_5634,N_5693);
nor U13254 (N_13254,N_6147,N_9824);
or U13255 (N_13255,N_8327,N_8724);
and U13256 (N_13256,N_5838,N_8364);
nor U13257 (N_13257,N_7249,N_7670);
nand U13258 (N_13258,N_8840,N_7216);
or U13259 (N_13259,N_5778,N_6530);
or U13260 (N_13260,N_5685,N_9217);
or U13261 (N_13261,N_6598,N_9981);
nand U13262 (N_13262,N_5772,N_7578);
and U13263 (N_13263,N_8570,N_5431);
nand U13264 (N_13264,N_6588,N_9001);
nor U13265 (N_13265,N_7715,N_9608);
nand U13266 (N_13266,N_7956,N_7502);
and U13267 (N_13267,N_5342,N_6866);
nor U13268 (N_13268,N_8590,N_6196);
nand U13269 (N_13269,N_7120,N_8700);
nor U13270 (N_13270,N_6317,N_9848);
or U13271 (N_13271,N_7682,N_6152);
or U13272 (N_13272,N_8378,N_6956);
nor U13273 (N_13273,N_6954,N_6302);
nor U13274 (N_13274,N_6888,N_9646);
nor U13275 (N_13275,N_6611,N_5956);
and U13276 (N_13276,N_7099,N_8392);
or U13277 (N_13277,N_9987,N_5100);
nor U13278 (N_13278,N_6844,N_7399);
or U13279 (N_13279,N_6975,N_8276);
and U13280 (N_13280,N_9182,N_6742);
nor U13281 (N_13281,N_5010,N_8810);
nor U13282 (N_13282,N_7853,N_9788);
and U13283 (N_13283,N_6541,N_7972);
nor U13284 (N_13284,N_7490,N_5132);
xnor U13285 (N_13285,N_5225,N_8363);
nor U13286 (N_13286,N_7556,N_7464);
and U13287 (N_13287,N_9157,N_8535);
nand U13288 (N_13288,N_6399,N_9108);
nand U13289 (N_13289,N_8222,N_6634);
and U13290 (N_13290,N_8120,N_9362);
nor U13291 (N_13291,N_6546,N_8188);
nor U13292 (N_13292,N_8141,N_9880);
nand U13293 (N_13293,N_6610,N_8663);
nand U13294 (N_13294,N_9273,N_9034);
and U13295 (N_13295,N_6896,N_9338);
or U13296 (N_13296,N_8615,N_7289);
or U13297 (N_13297,N_5172,N_8556);
nor U13298 (N_13298,N_9209,N_8301);
or U13299 (N_13299,N_6638,N_5271);
nand U13300 (N_13300,N_5066,N_7479);
nand U13301 (N_13301,N_8817,N_9040);
nor U13302 (N_13302,N_6373,N_8045);
nand U13303 (N_13303,N_8734,N_5437);
nor U13304 (N_13304,N_6593,N_5668);
or U13305 (N_13305,N_5112,N_5949);
and U13306 (N_13306,N_7980,N_6205);
nor U13307 (N_13307,N_8224,N_9261);
or U13308 (N_13308,N_7232,N_6157);
nand U13309 (N_13309,N_8838,N_9250);
and U13310 (N_13310,N_7753,N_6520);
nor U13311 (N_13311,N_8142,N_7226);
and U13312 (N_13312,N_8356,N_5703);
or U13313 (N_13313,N_5200,N_9606);
xnor U13314 (N_13314,N_8624,N_7904);
and U13315 (N_13315,N_8920,N_5797);
or U13316 (N_13316,N_6377,N_5049);
nor U13317 (N_13317,N_8347,N_7703);
or U13318 (N_13318,N_6563,N_5157);
nor U13319 (N_13319,N_7213,N_5433);
nand U13320 (N_13320,N_9531,N_7143);
nor U13321 (N_13321,N_6265,N_5843);
nor U13322 (N_13322,N_8456,N_6487);
nor U13323 (N_13323,N_7901,N_8968);
and U13324 (N_13324,N_7333,N_5694);
xnor U13325 (N_13325,N_8728,N_7695);
nor U13326 (N_13326,N_7151,N_9125);
and U13327 (N_13327,N_5086,N_6188);
nand U13328 (N_13328,N_9847,N_5291);
nor U13329 (N_13329,N_7152,N_7274);
nand U13330 (N_13330,N_7624,N_7497);
nand U13331 (N_13331,N_6931,N_8857);
nor U13332 (N_13332,N_8432,N_8981);
nand U13333 (N_13333,N_7971,N_5935);
nand U13334 (N_13334,N_8167,N_7755);
or U13335 (N_13335,N_7656,N_9473);
nand U13336 (N_13336,N_9287,N_7983);
xnor U13337 (N_13337,N_7788,N_8375);
nand U13338 (N_13338,N_8333,N_5087);
or U13339 (N_13339,N_9374,N_5904);
xor U13340 (N_13340,N_6040,N_5357);
or U13341 (N_13341,N_8865,N_6672);
and U13342 (N_13342,N_6780,N_7200);
nor U13343 (N_13343,N_6142,N_8995);
and U13344 (N_13344,N_8506,N_6701);
and U13345 (N_13345,N_5910,N_9660);
and U13346 (N_13346,N_7852,N_5372);
or U13347 (N_13347,N_7619,N_7340);
or U13348 (N_13348,N_8824,N_5066);
and U13349 (N_13349,N_6822,N_6450);
nor U13350 (N_13350,N_6920,N_9495);
nand U13351 (N_13351,N_5298,N_8924);
and U13352 (N_13352,N_9619,N_5416);
and U13353 (N_13353,N_5402,N_9765);
and U13354 (N_13354,N_7851,N_5437);
nor U13355 (N_13355,N_5416,N_7775);
or U13356 (N_13356,N_9204,N_6125);
nand U13357 (N_13357,N_7587,N_7008);
or U13358 (N_13358,N_8645,N_9449);
xor U13359 (N_13359,N_6619,N_8021);
and U13360 (N_13360,N_6594,N_9695);
or U13361 (N_13361,N_5719,N_8214);
or U13362 (N_13362,N_7348,N_8106);
nand U13363 (N_13363,N_8135,N_8261);
or U13364 (N_13364,N_6136,N_5882);
or U13365 (N_13365,N_7147,N_6866);
and U13366 (N_13366,N_6054,N_7863);
and U13367 (N_13367,N_9552,N_6662);
nor U13368 (N_13368,N_7093,N_5092);
xnor U13369 (N_13369,N_8113,N_8028);
nand U13370 (N_13370,N_6490,N_9057);
or U13371 (N_13371,N_9298,N_6107);
nor U13372 (N_13372,N_9986,N_6038);
nor U13373 (N_13373,N_9056,N_5702);
nand U13374 (N_13374,N_6259,N_7633);
nand U13375 (N_13375,N_8372,N_8563);
nor U13376 (N_13376,N_7323,N_9042);
and U13377 (N_13377,N_9659,N_6443);
nor U13378 (N_13378,N_9607,N_7718);
and U13379 (N_13379,N_5839,N_5540);
and U13380 (N_13380,N_5160,N_5505);
nand U13381 (N_13381,N_6725,N_8452);
nor U13382 (N_13382,N_7353,N_7774);
and U13383 (N_13383,N_9615,N_5953);
nand U13384 (N_13384,N_7012,N_5168);
and U13385 (N_13385,N_9148,N_5169);
nor U13386 (N_13386,N_5836,N_6976);
nand U13387 (N_13387,N_7154,N_6950);
or U13388 (N_13388,N_9757,N_6237);
nand U13389 (N_13389,N_7771,N_8711);
nand U13390 (N_13390,N_9620,N_7719);
nand U13391 (N_13391,N_9320,N_9907);
and U13392 (N_13392,N_7483,N_8698);
or U13393 (N_13393,N_7918,N_8234);
and U13394 (N_13394,N_8935,N_5045);
nor U13395 (N_13395,N_5991,N_8740);
nor U13396 (N_13396,N_9058,N_9723);
nand U13397 (N_13397,N_9549,N_6462);
or U13398 (N_13398,N_6474,N_5356);
nand U13399 (N_13399,N_6850,N_7597);
nand U13400 (N_13400,N_8409,N_5380);
or U13401 (N_13401,N_9255,N_8913);
nor U13402 (N_13402,N_7766,N_9075);
nor U13403 (N_13403,N_7902,N_6553);
nand U13404 (N_13404,N_5575,N_5421);
nand U13405 (N_13405,N_6098,N_5003);
nor U13406 (N_13406,N_8694,N_5100);
nand U13407 (N_13407,N_6650,N_6224);
nand U13408 (N_13408,N_5016,N_9622);
and U13409 (N_13409,N_7503,N_6515);
and U13410 (N_13410,N_9197,N_7496);
and U13411 (N_13411,N_8191,N_6623);
nor U13412 (N_13412,N_9026,N_5335);
xor U13413 (N_13413,N_7365,N_7258);
or U13414 (N_13414,N_9857,N_6261);
nand U13415 (N_13415,N_7152,N_6142);
nor U13416 (N_13416,N_9650,N_5143);
xor U13417 (N_13417,N_8073,N_8023);
nand U13418 (N_13418,N_6727,N_6605);
nor U13419 (N_13419,N_6390,N_6883);
or U13420 (N_13420,N_8994,N_7992);
nor U13421 (N_13421,N_8647,N_7348);
or U13422 (N_13422,N_8160,N_7247);
nor U13423 (N_13423,N_7102,N_7387);
nand U13424 (N_13424,N_8715,N_8806);
nor U13425 (N_13425,N_9946,N_7229);
and U13426 (N_13426,N_9177,N_6247);
nor U13427 (N_13427,N_9292,N_5694);
or U13428 (N_13428,N_9808,N_7170);
nor U13429 (N_13429,N_6491,N_9260);
nand U13430 (N_13430,N_6490,N_7896);
nand U13431 (N_13431,N_7101,N_8194);
xor U13432 (N_13432,N_9303,N_6724);
nor U13433 (N_13433,N_8727,N_8649);
nand U13434 (N_13434,N_7361,N_9534);
nand U13435 (N_13435,N_7789,N_7327);
and U13436 (N_13436,N_6500,N_5532);
nor U13437 (N_13437,N_8749,N_5439);
nor U13438 (N_13438,N_6535,N_7490);
or U13439 (N_13439,N_8271,N_5160);
nand U13440 (N_13440,N_8238,N_9887);
nand U13441 (N_13441,N_8975,N_7046);
nand U13442 (N_13442,N_8543,N_8514);
and U13443 (N_13443,N_8890,N_8295);
nor U13444 (N_13444,N_5640,N_9708);
nand U13445 (N_13445,N_6114,N_6197);
nor U13446 (N_13446,N_9476,N_9891);
and U13447 (N_13447,N_9011,N_9614);
or U13448 (N_13448,N_7772,N_6928);
and U13449 (N_13449,N_7438,N_7246);
and U13450 (N_13450,N_7995,N_5116);
nand U13451 (N_13451,N_5231,N_5138);
nor U13452 (N_13452,N_9788,N_6422);
or U13453 (N_13453,N_5713,N_7944);
nor U13454 (N_13454,N_5106,N_8969);
or U13455 (N_13455,N_5653,N_9543);
nand U13456 (N_13456,N_5299,N_9690);
nand U13457 (N_13457,N_9528,N_8342);
and U13458 (N_13458,N_9607,N_9525);
or U13459 (N_13459,N_8873,N_9305);
and U13460 (N_13460,N_9517,N_6360);
nor U13461 (N_13461,N_5935,N_5223);
or U13462 (N_13462,N_7928,N_5833);
nand U13463 (N_13463,N_5171,N_8223);
or U13464 (N_13464,N_7819,N_7869);
nand U13465 (N_13465,N_9149,N_9121);
or U13466 (N_13466,N_5492,N_9316);
and U13467 (N_13467,N_8979,N_6464);
and U13468 (N_13468,N_6829,N_6998);
and U13469 (N_13469,N_8524,N_7425);
nor U13470 (N_13470,N_7531,N_8057);
or U13471 (N_13471,N_8911,N_9142);
nand U13472 (N_13472,N_9356,N_6369);
or U13473 (N_13473,N_8250,N_8203);
or U13474 (N_13474,N_8497,N_5198);
or U13475 (N_13475,N_5621,N_7886);
or U13476 (N_13476,N_7544,N_8363);
and U13477 (N_13477,N_6267,N_7226);
or U13478 (N_13478,N_6285,N_7896);
nor U13479 (N_13479,N_8836,N_8940);
nand U13480 (N_13480,N_9715,N_5720);
or U13481 (N_13481,N_7285,N_9323);
nor U13482 (N_13482,N_7985,N_5279);
nand U13483 (N_13483,N_7255,N_6496);
nor U13484 (N_13484,N_5383,N_7501);
or U13485 (N_13485,N_8168,N_5652);
nand U13486 (N_13486,N_5664,N_9685);
nand U13487 (N_13487,N_5870,N_6908);
nor U13488 (N_13488,N_8505,N_7193);
or U13489 (N_13489,N_5385,N_5615);
nand U13490 (N_13490,N_9234,N_5303);
and U13491 (N_13491,N_5162,N_9361);
nand U13492 (N_13492,N_7894,N_5113);
or U13493 (N_13493,N_7069,N_9492);
or U13494 (N_13494,N_6340,N_5134);
xor U13495 (N_13495,N_8122,N_7226);
nor U13496 (N_13496,N_8498,N_5532);
and U13497 (N_13497,N_5270,N_8773);
nand U13498 (N_13498,N_5129,N_5063);
or U13499 (N_13499,N_5510,N_8059);
nand U13500 (N_13500,N_5604,N_6113);
nand U13501 (N_13501,N_5962,N_5687);
or U13502 (N_13502,N_9059,N_9052);
and U13503 (N_13503,N_5061,N_6348);
nand U13504 (N_13504,N_5592,N_5509);
or U13505 (N_13505,N_6220,N_8409);
nor U13506 (N_13506,N_9191,N_9985);
or U13507 (N_13507,N_6227,N_6410);
nand U13508 (N_13508,N_6872,N_6723);
and U13509 (N_13509,N_5655,N_5085);
and U13510 (N_13510,N_8590,N_5789);
nand U13511 (N_13511,N_9239,N_6748);
or U13512 (N_13512,N_6000,N_7511);
nor U13513 (N_13513,N_6186,N_7389);
or U13514 (N_13514,N_7276,N_8097);
nand U13515 (N_13515,N_5608,N_8624);
or U13516 (N_13516,N_7586,N_8600);
nor U13517 (N_13517,N_9007,N_6020);
nor U13518 (N_13518,N_5168,N_6209);
nor U13519 (N_13519,N_6452,N_7440);
nor U13520 (N_13520,N_6613,N_6982);
and U13521 (N_13521,N_6906,N_7952);
nor U13522 (N_13522,N_6756,N_8989);
nor U13523 (N_13523,N_6961,N_6312);
or U13524 (N_13524,N_9830,N_6537);
nand U13525 (N_13525,N_9604,N_6418);
nor U13526 (N_13526,N_9159,N_9464);
nand U13527 (N_13527,N_7411,N_5142);
or U13528 (N_13528,N_7551,N_5381);
and U13529 (N_13529,N_7902,N_6495);
or U13530 (N_13530,N_8867,N_7848);
xnor U13531 (N_13531,N_6588,N_6443);
or U13532 (N_13532,N_8875,N_8240);
or U13533 (N_13533,N_8727,N_7799);
or U13534 (N_13534,N_5051,N_9251);
and U13535 (N_13535,N_5573,N_5308);
nor U13536 (N_13536,N_9066,N_9118);
or U13537 (N_13537,N_5972,N_6642);
nor U13538 (N_13538,N_9602,N_8774);
and U13539 (N_13539,N_8325,N_8639);
and U13540 (N_13540,N_5515,N_8415);
and U13541 (N_13541,N_6374,N_7243);
or U13542 (N_13542,N_7806,N_7415);
nand U13543 (N_13543,N_9258,N_7503);
nand U13544 (N_13544,N_5357,N_7708);
and U13545 (N_13545,N_6388,N_7240);
nand U13546 (N_13546,N_9487,N_5205);
nor U13547 (N_13547,N_8326,N_6390);
xor U13548 (N_13548,N_7267,N_8034);
and U13549 (N_13549,N_5646,N_9559);
or U13550 (N_13550,N_9121,N_5865);
nor U13551 (N_13551,N_7870,N_5125);
nand U13552 (N_13552,N_8755,N_5939);
nand U13553 (N_13553,N_7453,N_6114);
nand U13554 (N_13554,N_9905,N_7504);
and U13555 (N_13555,N_5595,N_5824);
nor U13556 (N_13556,N_8315,N_8991);
or U13557 (N_13557,N_8270,N_9004);
nand U13558 (N_13558,N_9982,N_8529);
nor U13559 (N_13559,N_8262,N_5175);
or U13560 (N_13560,N_6312,N_8097);
or U13561 (N_13561,N_5752,N_9577);
nor U13562 (N_13562,N_6552,N_8913);
and U13563 (N_13563,N_5384,N_9430);
and U13564 (N_13564,N_8348,N_9758);
nor U13565 (N_13565,N_7302,N_8684);
nor U13566 (N_13566,N_9594,N_8306);
or U13567 (N_13567,N_8876,N_8489);
and U13568 (N_13568,N_9534,N_5341);
nor U13569 (N_13569,N_5215,N_5160);
nand U13570 (N_13570,N_9826,N_5859);
nor U13571 (N_13571,N_7185,N_8872);
nand U13572 (N_13572,N_8652,N_9816);
or U13573 (N_13573,N_7784,N_7016);
nor U13574 (N_13574,N_8877,N_9330);
nand U13575 (N_13575,N_9118,N_7819);
nor U13576 (N_13576,N_5511,N_8713);
and U13577 (N_13577,N_9816,N_8226);
and U13578 (N_13578,N_6505,N_9585);
nor U13579 (N_13579,N_6186,N_6371);
and U13580 (N_13580,N_9778,N_8563);
nor U13581 (N_13581,N_7422,N_7821);
nor U13582 (N_13582,N_5272,N_5343);
or U13583 (N_13583,N_6764,N_5730);
nor U13584 (N_13584,N_6674,N_6214);
nand U13585 (N_13585,N_6490,N_7836);
nor U13586 (N_13586,N_7417,N_5960);
and U13587 (N_13587,N_7287,N_6630);
and U13588 (N_13588,N_6237,N_5635);
nand U13589 (N_13589,N_9757,N_9316);
nor U13590 (N_13590,N_6790,N_8132);
and U13591 (N_13591,N_9044,N_7890);
nand U13592 (N_13592,N_9663,N_9424);
nor U13593 (N_13593,N_8359,N_5595);
or U13594 (N_13594,N_7255,N_9328);
and U13595 (N_13595,N_5945,N_6413);
nor U13596 (N_13596,N_5543,N_6133);
nor U13597 (N_13597,N_8770,N_6239);
nand U13598 (N_13598,N_7463,N_5170);
or U13599 (N_13599,N_7831,N_5929);
nor U13600 (N_13600,N_7185,N_5679);
xnor U13601 (N_13601,N_5903,N_5727);
nor U13602 (N_13602,N_6301,N_7761);
and U13603 (N_13603,N_5029,N_9589);
nand U13604 (N_13604,N_5774,N_7514);
or U13605 (N_13605,N_6423,N_6179);
or U13606 (N_13606,N_7487,N_5087);
and U13607 (N_13607,N_9911,N_6221);
or U13608 (N_13608,N_5847,N_6357);
and U13609 (N_13609,N_6743,N_6251);
nand U13610 (N_13610,N_6899,N_7411);
nor U13611 (N_13611,N_6499,N_7903);
nand U13612 (N_13612,N_8428,N_7729);
nand U13613 (N_13613,N_9924,N_6347);
and U13614 (N_13614,N_7365,N_5901);
and U13615 (N_13615,N_6413,N_8664);
and U13616 (N_13616,N_7710,N_8288);
and U13617 (N_13617,N_6324,N_8786);
nor U13618 (N_13618,N_5441,N_9697);
nor U13619 (N_13619,N_8579,N_5103);
nor U13620 (N_13620,N_8966,N_7800);
nand U13621 (N_13621,N_6229,N_5445);
xnor U13622 (N_13622,N_8034,N_5569);
and U13623 (N_13623,N_9983,N_8612);
xnor U13624 (N_13624,N_8605,N_9456);
and U13625 (N_13625,N_5524,N_6213);
or U13626 (N_13626,N_9503,N_6486);
or U13627 (N_13627,N_7419,N_8835);
and U13628 (N_13628,N_8894,N_8422);
nor U13629 (N_13629,N_5240,N_6309);
nor U13630 (N_13630,N_8109,N_7663);
or U13631 (N_13631,N_5544,N_7285);
or U13632 (N_13632,N_9402,N_9802);
nor U13633 (N_13633,N_5140,N_6617);
nand U13634 (N_13634,N_9594,N_6944);
and U13635 (N_13635,N_8148,N_8043);
or U13636 (N_13636,N_7742,N_6896);
or U13637 (N_13637,N_9279,N_7755);
xnor U13638 (N_13638,N_8206,N_7624);
or U13639 (N_13639,N_7684,N_7625);
nand U13640 (N_13640,N_9348,N_6935);
or U13641 (N_13641,N_9062,N_6087);
and U13642 (N_13642,N_7717,N_6013);
nand U13643 (N_13643,N_5358,N_9448);
nor U13644 (N_13644,N_8864,N_7623);
nand U13645 (N_13645,N_6956,N_9661);
xor U13646 (N_13646,N_6408,N_9565);
nand U13647 (N_13647,N_9426,N_5274);
xor U13648 (N_13648,N_9573,N_8055);
nor U13649 (N_13649,N_8894,N_5451);
or U13650 (N_13650,N_8346,N_9171);
nand U13651 (N_13651,N_9693,N_5509);
nor U13652 (N_13652,N_7313,N_8436);
nand U13653 (N_13653,N_6923,N_8395);
nor U13654 (N_13654,N_7864,N_9295);
or U13655 (N_13655,N_6712,N_9306);
nand U13656 (N_13656,N_5740,N_6178);
nand U13657 (N_13657,N_6118,N_9137);
or U13658 (N_13658,N_6139,N_7744);
or U13659 (N_13659,N_8072,N_7857);
nand U13660 (N_13660,N_5303,N_7438);
nand U13661 (N_13661,N_8416,N_7721);
nor U13662 (N_13662,N_8259,N_7318);
nor U13663 (N_13663,N_6408,N_7742);
or U13664 (N_13664,N_6984,N_9939);
or U13665 (N_13665,N_5397,N_9419);
or U13666 (N_13666,N_8303,N_5036);
or U13667 (N_13667,N_9534,N_8878);
nor U13668 (N_13668,N_9490,N_6611);
or U13669 (N_13669,N_9571,N_9047);
and U13670 (N_13670,N_7597,N_5900);
nand U13671 (N_13671,N_8841,N_9244);
or U13672 (N_13672,N_9608,N_7996);
nand U13673 (N_13673,N_8325,N_7841);
nand U13674 (N_13674,N_9877,N_6942);
or U13675 (N_13675,N_9890,N_9108);
or U13676 (N_13676,N_5891,N_8677);
or U13677 (N_13677,N_6330,N_8196);
or U13678 (N_13678,N_7058,N_5551);
and U13679 (N_13679,N_8170,N_5868);
and U13680 (N_13680,N_9676,N_8217);
nor U13681 (N_13681,N_7773,N_5533);
nand U13682 (N_13682,N_7932,N_6295);
and U13683 (N_13683,N_9217,N_5270);
xnor U13684 (N_13684,N_6283,N_9753);
nand U13685 (N_13685,N_9868,N_6175);
and U13686 (N_13686,N_7953,N_9923);
or U13687 (N_13687,N_9347,N_7771);
nand U13688 (N_13688,N_8169,N_9594);
or U13689 (N_13689,N_5527,N_9564);
nand U13690 (N_13690,N_5736,N_7310);
nor U13691 (N_13691,N_8583,N_9044);
or U13692 (N_13692,N_5494,N_8587);
nor U13693 (N_13693,N_5071,N_6858);
or U13694 (N_13694,N_7004,N_7830);
and U13695 (N_13695,N_6773,N_8466);
nand U13696 (N_13696,N_5060,N_8399);
nor U13697 (N_13697,N_9967,N_9621);
nand U13698 (N_13698,N_5562,N_6687);
and U13699 (N_13699,N_8819,N_8786);
and U13700 (N_13700,N_7075,N_5270);
nor U13701 (N_13701,N_9039,N_7267);
and U13702 (N_13702,N_7610,N_8269);
or U13703 (N_13703,N_6315,N_5057);
nor U13704 (N_13704,N_9257,N_8624);
nor U13705 (N_13705,N_9876,N_8442);
nor U13706 (N_13706,N_5936,N_8443);
xnor U13707 (N_13707,N_8656,N_5881);
or U13708 (N_13708,N_7418,N_9782);
or U13709 (N_13709,N_6689,N_5830);
and U13710 (N_13710,N_5255,N_5536);
or U13711 (N_13711,N_9589,N_6958);
nor U13712 (N_13712,N_6037,N_8762);
or U13713 (N_13713,N_6619,N_7656);
nand U13714 (N_13714,N_6850,N_9423);
or U13715 (N_13715,N_9378,N_7426);
or U13716 (N_13716,N_5124,N_7090);
nand U13717 (N_13717,N_6655,N_6268);
nor U13718 (N_13718,N_8755,N_8919);
and U13719 (N_13719,N_7527,N_7585);
and U13720 (N_13720,N_5567,N_8589);
nor U13721 (N_13721,N_6484,N_8129);
nand U13722 (N_13722,N_6029,N_7790);
nor U13723 (N_13723,N_7276,N_7583);
nor U13724 (N_13724,N_9030,N_5523);
nand U13725 (N_13725,N_5468,N_9749);
and U13726 (N_13726,N_5857,N_6983);
nand U13727 (N_13727,N_8234,N_6071);
nor U13728 (N_13728,N_8512,N_7575);
and U13729 (N_13729,N_6483,N_5016);
xnor U13730 (N_13730,N_5451,N_5442);
or U13731 (N_13731,N_9258,N_7971);
nor U13732 (N_13732,N_5177,N_9511);
or U13733 (N_13733,N_8284,N_6945);
or U13734 (N_13734,N_6740,N_7333);
and U13735 (N_13735,N_7996,N_9273);
nand U13736 (N_13736,N_5082,N_9842);
and U13737 (N_13737,N_9035,N_8782);
and U13738 (N_13738,N_8520,N_9940);
and U13739 (N_13739,N_6893,N_5873);
nor U13740 (N_13740,N_5527,N_7220);
or U13741 (N_13741,N_6695,N_9995);
nand U13742 (N_13742,N_9755,N_8236);
nand U13743 (N_13743,N_8216,N_8297);
and U13744 (N_13744,N_7104,N_9008);
or U13745 (N_13745,N_9221,N_5877);
and U13746 (N_13746,N_5075,N_6986);
and U13747 (N_13747,N_5556,N_5835);
and U13748 (N_13748,N_8176,N_7244);
and U13749 (N_13749,N_5828,N_6406);
nand U13750 (N_13750,N_7868,N_8132);
nand U13751 (N_13751,N_8680,N_6989);
or U13752 (N_13752,N_5130,N_7977);
and U13753 (N_13753,N_6153,N_5019);
nand U13754 (N_13754,N_6084,N_6326);
and U13755 (N_13755,N_8101,N_8004);
nor U13756 (N_13756,N_7085,N_7818);
nand U13757 (N_13757,N_9558,N_6685);
or U13758 (N_13758,N_9135,N_9734);
or U13759 (N_13759,N_8591,N_8127);
and U13760 (N_13760,N_9078,N_6279);
and U13761 (N_13761,N_9572,N_8396);
nand U13762 (N_13762,N_9379,N_7027);
nor U13763 (N_13763,N_5661,N_7781);
and U13764 (N_13764,N_8105,N_6756);
nand U13765 (N_13765,N_6279,N_7759);
nor U13766 (N_13766,N_7886,N_8531);
or U13767 (N_13767,N_7607,N_9899);
nor U13768 (N_13768,N_7370,N_9560);
nor U13769 (N_13769,N_9031,N_8101);
or U13770 (N_13770,N_7442,N_5655);
nand U13771 (N_13771,N_5881,N_9948);
nand U13772 (N_13772,N_6342,N_5225);
nor U13773 (N_13773,N_6003,N_6022);
or U13774 (N_13774,N_7643,N_9757);
nand U13775 (N_13775,N_6824,N_6174);
nand U13776 (N_13776,N_7154,N_9852);
or U13777 (N_13777,N_8558,N_6109);
and U13778 (N_13778,N_5043,N_5057);
nand U13779 (N_13779,N_6666,N_7530);
nor U13780 (N_13780,N_7273,N_9282);
nand U13781 (N_13781,N_5434,N_9754);
nand U13782 (N_13782,N_7822,N_7710);
and U13783 (N_13783,N_5872,N_7065);
nor U13784 (N_13784,N_5745,N_5201);
nor U13785 (N_13785,N_8278,N_7934);
nand U13786 (N_13786,N_5820,N_6581);
nor U13787 (N_13787,N_7294,N_6212);
and U13788 (N_13788,N_6924,N_8227);
xnor U13789 (N_13789,N_8821,N_5155);
or U13790 (N_13790,N_5550,N_5631);
nand U13791 (N_13791,N_7172,N_7755);
or U13792 (N_13792,N_5916,N_7002);
or U13793 (N_13793,N_5747,N_8876);
and U13794 (N_13794,N_6431,N_7781);
and U13795 (N_13795,N_8748,N_8862);
nor U13796 (N_13796,N_7018,N_6751);
or U13797 (N_13797,N_7572,N_5982);
and U13798 (N_13798,N_9054,N_9257);
nand U13799 (N_13799,N_8094,N_8586);
nor U13800 (N_13800,N_7570,N_9514);
nor U13801 (N_13801,N_7039,N_6900);
nand U13802 (N_13802,N_9679,N_9859);
or U13803 (N_13803,N_8097,N_7419);
or U13804 (N_13804,N_7091,N_6019);
nand U13805 (N_13805,N_8015,N_5980);
and U13806 (N_13806,N_7212,N_7994);
and U13807 (N_13807,N_6449,N_5430);
or U13808 (N_13808,N_6699,N_9849);
or U13809 (N_13809,N_7307,N_6652);
nor U13810 (N_13810,N_8434,N_9259);
and U13811 (N_13811,N_9987,N_7231);
and U13812 (N_13812,N_9799,N_9280);
nor U13813 (N_13813,N_6411,N_7023);
xor U13814 (N_13814,N_5241,N_7608);
nand U13815 (N_13815,N_6490,N_8453);
or U13816 (N_13816,N_5064,N_8160);
nor U13817 (N_13817,N_9277,N_6111);
nand U13818 (N_13818,N_7318,N_6616);
or U13819 (N_13819,N_5336,N_8930);
nor U13820 (N_13820,N_7047,N_7771);
nor U13821 (N_13821,N_6797,N_5124);
nor U13822 (N_13822,N_6355,N_8571);
or U13823 (N_13823,N_8807,N_5211);
or U13824 (N_13824,N_5844,N_7013);
nand U13825 (N_13825,N_7417,N_8291);
nand U13826 (N_13826,N_6032,N_8491);
nand U13827 (N_13827,N_8873,N_9953);
or U13828 (N_13828,N_6459,N_5670);
and U13829 (N_13829,N_8950,N_9638);
or U13830 (N_13830,N_5471,N_7799);
and U13831 (N_13831,N_9986,N_5592);
nor U13832 (N_13832,N_8542,N_7887);
or U13833 (N_13833,N_9218,N_7379);
nand U13834 (N_13834,N_8582,N_6682);
and U13835 (N_13835,N_9060,N_8457);
or U13836 (N_13836,N_5472,N_7583);
and U13837 (N_13837,N_7735,N_6495);
or U13838 (N_13838,N_7663,N_9887);
nor U13839 (N_13839,N_9584,N_7573);
and U13840 (N_13840,N_7164,N_5111);
or U13841 (N_13841,N_9341,N_7075);
nand U13842 (N_13842,N_8491,N_9588);
or U13843 (N_13843,N_9848,N_5892);
nor U13844 (N_13844,N_9910,N_6241);
xnor U13845 (N_13845,N_9556,N_7059);
or U13846 (N_13846,N_7226,N_5249);
and U13847 (N_13847,N_9363,N_5756);
nor U13848 (N_13848,N_8177,N_8610);
nor U13849 (N_13849,N_8970,N_9374);
or U13850 (N_13850,N_9604,N_7990);
or U13851 (N_13851,N_9558,N_6886);
or U13852 (N_13852,N_7988,N_6527);
and U13853 (N_13853,N_5120,N_9544);
or U13854 (N_13854,N_6367,N_5927);
nor U13855 (N_13855,N_5273,N_6346);
nor U13856 (N_13856,N_5124,N_7826);
or U13857 (N_13857,N_6841,N_9513);
and U13858 (N_13858,N_9352,N_6086);
and U13859 (N_13859,N_5176,N_5846);
and U13860 (N_13860,N_5852,N_5832);
and U13861 (N_13861,N_5347,N_8091);
and U13862 (N_13862,N_6399,N_7741);
and U13863 (N_13863,N_5586,N_6880);
and U13864 (N_13864,N_8087,N_5678);
or U13865 (N_13865,N_7861,N_9573);
and U13866 (N_13866,N_9695,N_9603);
nor U13867 (N_13867,N_6315,N_9386);
or U13868 (N_13868,N_5882,N_9001);
nand U13869 (N_13869,N_9488,N_9446);
nor U13870 (N_13870,N_9660,N_8851);
nand U13871 (N_13871,N_6619,N_7237);
and U13872 (N_13872,N_5354,N_7367);
and U13873 (N_13873,N_7018,N_6096);
or U13874 (N_13874,N_5036,N_8625);
and U13875 (N_13875,N_6306,N_8023);
nor U13876 (N_13876,N_7856,N_8016);
and U13877 (N_13877,N_8380,N_5519);
and U13878 (N_13878,N_9901,N_7772);
nand U13879 (N_13879,N_5681,N_8709);
xor U13880 (N_13880,N_6729,N_7536);
or U13881 (N_13881,N_7680,N_7594);
and U13882 (N_13882,N_5514,N_8907);
and U13883 (N_13883,N_8730,N_9933);
nand U13884 (N_13884,N_8831,N_5517);
and U13885 (N_13885,N_5477,N_6052);
nand U13886 (N_13886,N_7151,N_6374);
or U13887 (N_13887,N_8530,N_8845);
and U13888 (N_13888,N_6989,N_6852);
or U13889 (N_13889,N_7716,N_6148);
or U13890 (N_13890,N_5303,N_7844);
or U13891 (N_13891,N_6069,N_8932);
nor U13892 (N_13892,N_7001,N_7866);
and U13893 (N_13893,N_6406,N_6249);
nand U13894 (N_13894,N_5652,N_6626);
nor U13895 (N_13895,N_5438,N_8511);
or U13896 (N_13896,N_6951,N_5335);
or U13897 (N_13897,N_9132,N_6425);
nand U13898 (N_13898,N_9203,N_6769);
or U13899 (N_13899,N_8493,N_5785);
or U13900 (N_13900,N_5561,N_6931);
nor U13901 (N_13901,N_8429,N_7874);
nor U13902 (N_13902,N_5207,N_9500);
and U13903 (N_13903,N_7646,N_9294);
nor U13904 (N_13904,N_6171,N_6204);
or U13905 (N_13905,N_7982,N_9628);
and U13906 (N_13906,N_9450,N_5102);
and U13907 (N_13907,N_5874,N_8916);
and U13908 (N_13908,N_9339,N_9780);
nand U13909 (N_13909,N_7865,N_8472);
and U13910 (N_13910,N_9543,N_8704);
nor U13911 (N_13911,N_6414,N_9147);
nor U13912 (N_13912,N_5520,N_8237);
nor U13913 (N_13913,N_8021,N_9609);
and U13914 (N_13914,N_6510,N_6829);
nand U13915 (N_13915,N_5963,N_5431);
or U13916 (N_13916,N_6243,N_9414);
or U13917 (N_13917,N_7510,N_5973);
nand U13918 (N_13918,N_8823,N_7474);
and U13919 (N_13919,N_8307,N_7661);
nor U13920 (N_13920,N_8070,N_9054);
or U13921 (N_13921,N_5418,N_6629);
nand U13922 (N_13922,N_6900,N_8846);
nand U13923 (N_13923,N_7199,N_6517);
and U13924 (N_13924,N_9688,N_9166);
xor U13925 (N_13925,N_5990,N_9257);
nor U13926 (N_13926,N_9357,N_6659);
or U13927 (N_13927,N_7083,N_5783);
nor U13928 (N_13928,N_5406,N_7712);
nand U13929 (N_13929,N_6778,N_5752);
nor U13930 (N_13930,N_7589,N_6518);
or U13931 (N_13931,N_6237,N_5328);
and U13932 (N_13932,N_7519,N_7633);
or U13933 (N_13933,N_7627,N_8719);
nor U13934 (N_13934,N_9752,N_9498);
or U13935 (N_13935,N_5969,N_8638);
and U13936 (N_13936,N_7379,N_7371);
and U13937 (N_13937,N_7948,N_9211);
or U13938 (N_13938,N_6831,N_7199);
nand U13939 (N_13939,N_9983,N_5932);
or U13940 (N_13940,N_7319,N_5548);
or U13941 (N_13941,N_9090,N_9309);
or U13942 (N_13942,N_8865,N_9888);
nand U13943 (N_13943,N_8389,N_9382);
nor U13944 (N_13944,N_7296,N_6727);
nor U13945 (N_13945,N_8474,N_9700);
nor U13946 (N_13946,N_7187,N_8299);
nor U13947 (N_13947,N_7706,N_9833);
or U13948 (N_13948,N_5740,N_8820);
nor U13949 (N_13949,N_9318,N_6385);
or U13950 (N_13950,N_9543,N_6763);
or U13951 (N_13951,N_5685,N_5679);
nand U13952 (N_13952,N_5788,N_9180);
nand U13953 (N_13953,N_5585,N_8112);
nor U13954 (N_13954,N_5233,N_9834);
nor U13955 (N_13955,N_5342,N_9206);
and U13956 (N_13956,N_6957,N_6738);
or U13957 (N_13957,N_8638,N_8959);
and U13958 (N_13958,N_8480,N_5555);
nor U13959 (N_13959,N_8598,N_5161);
xor U13960 (N_13960,N_8096,N_7091);
nor U13961 (N_13961,N_5122,N_5821);
nor U13962 (N_13962,N_7246,N_9518);
nand U13963 (N_13963,N_8662,N_9349);
and U13964 (N_13964,N_9889,N_6087);
and U13965 (N_13965,N_5716,N_5213);
xor U13966 (N_13966,N_8662,N_8689);
nand U13967 (N_13967,N_7596,N_7599);
nand U13968 (N_13968,N_8848,N_6529);
nor U13969 (N_13969,N_9147,N_5879);
or U13970 (N_13970,N_7316,N_5761);
and U13971 (N_13971,N_6229,N_5036);
and U13972 (N_13972,N_7977,N_5429);
or U13973 (N_13973,N_7604,N_7905);
nor U13974 (N_13974,N_5613,N_6787);
nand U13975 (N_13975,N_8554,N_8047);
nand U13976 (N_13976,N_8541,N_8258);
nand U13977 (N_13977,N_8953,N_6671);
and U13978 (N_13978,N_8616,N_9226);
or U13979 (N_13979,N_6143,N_9761);
and U13980 (N_13980,N_9553,N_5545);
nand U13981 (N_13981,N_9157,N_5386);
and U13982 (N_13982,N_9687,N_7999);
and U13983 (N_13983,N_8364,N_5186);
nor U13984 (N_13984,N_5677,N_5048);
nand U13985 (N_13985,N_7676,N_8620);
nor U13986 (N_13986,N_6358,N_9891);
and U13987 (N_13987,N_8149,N_5585);
nor U13988 (N_13988,N_5405,N_7472);
or U13989 (N_13989,N_6646,N_9140);
nor U13990 (N_13990,N_7483,N_8631);
or U13991 (N_13991,N_9334,N_8467);
nand U13992 (N_13992,N_9883,N_7985);
nor U13993 (N_13993,N_9046,N_5759);
nand U13994 (N_13994,N_5363,N_7979);
and U13995 (N_13995,N_5778,N_6105);
nand U13996 (N_13996,N_9646,N_7773);
nand U13997 (N_13997,N_5962,N_5511);
nor U13998 (N_13998,N_7309,N_7401);
and U13999 (N_13999,N_7272,N_7100);
and U14000 (N_14000,N_9370,N_8866);
and U14001 (N_14001,N_9253,N_6413);
nand U14002 (N_14002,N_6330,N_8418);
nor U14003 (N_14003,N_7215,N_5463);
or U14004 (N_14004,N_7978,N_7276);
nand U14005 (N_14005,N_7683,N_6766);
nand U14006 (N_14006,N_6620,N_8880);
or U14007 (N_14007,N_8093,N_9012);
or U14008 (N_14008,N_5040,N_7685);
or U14009 (N_14009,N_6764,N_5379);
or U14010 (N_14010,N_6135,N_7113);
nand U14011 (N_14011,N_8918,N_9147);
nand U14012 (N_14012,N_6123,N_5526);
or U14013 (N_14013,N_9403,N_9522);
or U14014 (N_14014,N_8271,N_8350);
or U14015 (N_14015,N_6728,N_7088);
or U14016 (N_14016,N_8340,N_6698);
and U14017 (N_14017,N_6725,N_7839);
xor U14018 (N_14018,N_7959,N_7403);
nand U14019 (N_14019,N_8334,N_5162);
or U14020 (N_14020,N_5717,N_6067);
nor U14021 (N_14021,N_6726,N_8322);
or U14022 (N_14022,N_5862,N_5363);
nand U14023 (N_14023,N_9674,N_6173);
or U14024 (N_14024,N_9597,N_5623);
nor U14025 (N_14025,N_9333,N_8479);
nor U14026 (N_14026,N_6185,N_8570);
nor U14027 (N_14027,N_7494,N_8270);
and U14028 (N_14028,N_9951,N_8362);
or U14029 (N_14029,N_8290,N_5562);
nor U14030 (N_14030,N_5307,N_9671);
and U14031 (N_14031,N_6681,N_6491);
or U14032 (N_14032,N_9400,N_9121);
and U14033 (N_14033,N_6926,N_5348);
nand U14034 (N_14034,N_8159,N_7700);
nand U14035 (N_14035,N_9457,N_7732);
and U14036 (N_14036,N_8201,N_7730);
and U14037 (N_14037,N_7879,N_9325);
nand U14038 (N_14038,N_9876,N_7870);
or U14039 (N_14039,N_8293,N_8036);
nand U14040 (N_14040,N_8678,N_8883);
or U14041 (N_14041,N_6068,N_6817);
nand U14042 (N_14042,N_9331,N_8180);
or U14043 (N_14043,N_6167,N_7167);
nand U14044 (N_14044,N_5686,N_9804);
and U14045 (N_14045,N_5298,N_8267);
nor U14046 (N_14046,N_8365,N_6243);
and U14047 (N_14047,N_5933,N_9634);
nor U14048 (N_14048,N_5504,N_9477);
or U14049 (N_14049,N_9032,N_8452);
or U14050 (N_14050,N_6375,N_5641);
nand U14051 (N_14051,N_6843,N_8668);
nand U14052 (N_14052,N_5127,N_9049);
and U14053 (N_14053,N_6369,N_9612);
and U14054 (N_14054,N_6448,N_8603);
and U14055 (N_14055,N_6164,N_6592);
nor U14056 (N_14056,N_7694,N_9454);
and U14057 (N_14057,N_5879,N_9628);
nor U14058 (N_14058,N_5860,N_5591);
nand U14059 (N_14059,N_8466,N_7550);
and U14060 (N_14060,N_5684,N_7351);
or U14061 (N_14061,N_7585,N_7784);
or U14062 (N_14062,N_9283,N_6985);
nand U14063 (N_14063,N_6747,N_9210);
and U14064 (N_14064,N_5857,N_8489);
and U14065 (N_14065,N_9679,N_9972);
nor U14066 (N_14066,N_7635,N_8519);
nor U14067 (N_14067,N_5234,N_5225);
or U14068 (N_14068,N_8453,N_6946);
nand U14069 (N_14069,N_5773,N_9407);
nand U14070 (N_14070,N_8319,N_7638);
or U14071 (N_14071,N_9170,N_8929);
nand U14072 (N_14072,N_8613,N_6336);
nor U14073 (N_14073,N_8474,N_6922);
xnor U14074 (N_14074,N_5292,N_6607);
and U14075 (N_14075,N_5981,N_6677);
nand U14076 (N_14076,N_5801,N_9076);
and U14077 (N_14077,N_8797,N_6558);
and U14078 (N_14078,N_9160,N_8830);
and U14079 (N_14079,N_8920,N_7710);
or U14080 (N_14080,N_6419,N_9180);
nor U14081 (N_14081,N_5144,N_7927);
nor U14082 (N_14082,N_6846,N_9215);
nand U14083 (N_14083,N_8768,N_8496);
nor U14084 (N_14084,N_9061,N_5709);
nand U14085 (N_14085,N_9198,N_7191);
nand U14086 (N_14086,N_7948,N_8286);
nor U14087 (N_14087,N_7880,N_6982);
nand U14088 (N_14088,N_7833,N_9184);
nand U14089 (N_14089,N_8928,N_6199);
nand U14090 (N_14090,N_6094,N_5427);
nand U14091 (N_14091,N_7621,N_9730);
nand U14092 (N_14092,N_9810,N_8780);
and U14093 (N_14093,N_5779,N_7493);
nand U14094 (N_14094,N_7530,N_7358);
and U14095 (N_14095,N_8923,N_9774);
nor U14096 (N_14096,N_7639,N_9767);
nand U14097 (N_14097,N_9166,N_9460);
and U14098 (N_14098,N_8486,N_5924);
nand U14099 (N_14099,N_6022,N_7810);
nor U14100 (N_14100,N_8020,N_8900);
nand U14101 (N_14101,N_5537,N_9420);
nand U14102 (N_14102,N_8528,N_7065);
nor U14103 (N_14103,N_6306,N_9631);
nor U14104 (N_14104,N_5298,N_9382);
nor U14105 (N_14105,N_5984,N_8072);
nand U14106 (N_14106,N_8296,N_5506);
nor U14107 (N_14107,N_5093,N_6932);
nand U14108 (N_14108,N_7771,N_7284);
nand U14109 (N_14109,N_7130,N_6484);
and U14110 (N_14110,N_6710,N_8014);
nand U14111 (N_14111,N_5407,N_7503);
nand U14112 (N_14112,N_9095,N_8285);
xor U14113 (N_14113,N_6449,N_8942);
nor U14114 (N_14114,N_7593,N_8826);
nand U14115 (N_14115,N_8170,N_8684);
nor U14116 (N_14116,N_7681,N_9045);
or U14117 (N_14117,N_7882,N_8752);
and U14118 (N_14118,N_5390,N_9686);
or U14119 (N_14119,N_9579,N_9364);
and U14120 (N_14120,N_5366,N_7237);
nand U14121 (N_14121,N_8896,N_5745);
and U14122 (N_14122,N_7065,N_5805);
nor U14123 (N_14123,N_5080,N_9231);
or U14124 (N_14124,N_6098,N_8422);
nand U14125 (N_14125,N_8886,N_7686);
nor U14126 (N_14126,N_6976,N_9944);
or U14127 (N_14127,N_8554,N_7802);
nor U14128 (N_14128,N_7262,N_5494);
and U14129 (N_14129,N_6119,N_5535);
nor U14130 (N_14130,N_9454,N_7420);
or U14131 (N_14131,N_8165,N_7585);
nor U14132 (N_14132,N_8650,N_5213);
or U14133 (N_14133,N_8089,N_6131);
and U14134 (N_14134,N_7159,N_6788);
or U14135 (N_14135,N_8062,N_5687);
nand U14136 (N_14136,N_7442,N_5642);
nand U14137 (N_14137,N_9471,N_9531);
nor U14138 (N_14138,N_5502,N_7286);
nor U14139 (N_14139,N_6051,N_6118);
or U14140 (N_14140,N_8241,N_9281);
or U14141 (N_14141,N_5311,N_8426);
nand U14142 (N_14142,N_6935,N_8337);
or U14143 (N_14143,N_9415,N_9110);
or U14144 (N_14144,N_7604,N_6798);
and U14145 (N_14145,N_6754,N_5728);
and U14146 (N_14146,N_7086,N_5589);
or U14147 (N_14147,N_8294,N_7018);
or U14148 (N_14148,N_7139,N_5576);
and U14149 (N_14149,N_6939,N_8746);
nor U14150 (N_14150,N_7904,N_7125);
nand U14151 (N_14151,N_6643,N_8978);
nand U14152 (N_14152,N_7009,N_5832);
or U14153 (N_14153,N_9494,N_5239);
nand U14154 (N_14154,N_7957,N_9199);
nor U14155 (N_14155,N_6265,N_7581);
and U14156 (N_14156,N_5058,N_5829);
or U14157 (N_14157,N_6944,N_5189);
and U14158 (N_14158,N_6883,N_9994);
nand U14159 (N_14159,N_5816,N_9606);
xor U14160 (N_14160,N_9019,N_9822);
nand U14161 (N_14161,N_9304,N_5429);
or U14162 (N_14162,N_8250,N_7733);
nor U14163 (N_14163,N_8764,N_9155);
nand U14164 (N_14164,N_6065,N_8115);
and U14165 (N_14165,N_9087,N_9702);
and U14166 (N_14166,N_9257,N_7808);
nor U14167 (N_14167,N_5719,N_9531);
nor U14168 (N_14168,N_9365,N_5124);
or U14169 (N_14169,N_8776,N_9618);
or U14170 (N_14170,N_7140,N_6047);
or U14171 (N_14171,N_9450,N_8720);
nor U14172 (N_14172,N_8691,N_7655);
nand U14173 (N_14173,N_9696,N_9516);
or U14174 (N_14174,N_6156,N_9298);
or U14175 (N_14175,N_9519,N_9656);
or U14176 (N_14176,N_7534,N_7476);
and U14177 (N_14177,N_9982,N_8403);
or U14178 (N_14178,N_8803,N_9272);
and U14179 (N_14179,N_7050,N_7331);
nor U14180 (N_14180,N_5543,N_5650);
and U14181 (N_14181,N_9154,N_9011);
nor U14182 (N_14182,N_8591,N_9934);
and U14183 (N_14183,N_5578,N_6502);
xnor U14184 (N_14184,N_8053,N_7052);
nor U14185 (N_14185,N_7602,N_7745);
or U14186 (N_14186,N_8302,N_7518);
and U14187 (N_14187,N_9232,N_9305);
nor U14188 (N_14188,N_6830,N_7430);
nand U14189 (N_14189,N_9485,N_7177);
nor U14190 (N_14190,N_9266,N_6174);
or U14191 (N_14191,N_5132,N_5162);
nand U14192 (N_14192,N_6629,N_6680);
nand U14193 (N_14193,N_5527,N_7632);
and U14194 (N_14194,N_6536,N_5595);
or U14195 (N_14195,N_9137,N_9563);
nand U14196 (N_14196,N_9864,N_5563);
nor U14197 (N_14197,N_6801,N_7131);
nor U14198 (N_14198,N_7621,N_6203);
nand U14199 (N_14199,N_7682,N_8334);
nor U14200 (N_14200,N_7347,N_9534);
nor U14201 (N_14201,N_6241,N_5428);
or U14202 (N_14202,N_5886,N_8365);
or U14203 (N_14203,N_6846,N_7159);
or U14204 (N_14204,N_6230,N_5000);
and U14205 (N_14205,N_8461,N_7687);
or U14206 (N_14206,N_9466,N_6450);
nand U14207 (N_14207,N_5376,N_6698);
xnor U14208 (N_14208,N_8070,N_6771);
nand U14209 (N_14209,N_8781,N_7352);
nor U14210 (N_14210,N_7702,N_7850);
nor U14211 (N_14211,N_7593,N_6988);
and U14212 (N_14212,N_5163,N_6288);
and U14213 (N_14213,N_6422,N_7344);
nand U14214 (N_14214,N_7915,N_5438);
and U14215 (N_14215,N_5211,N_9965);
or U14216 (N_14216,N_9096,N_8028);
and U14217 (N_14217,N_5737,N_8668);
nand U14218 (N_14218,N_6438,N_8317);
nand U14219 (N_14219,N_5050,N_6953);
nand U14220 (N_14220,N_7591,N_7530);
nand U14221 (N_14221,N_9511,N_5704);
and U14222 (N_14222,N_9194,N_5057);
nand U14223 (N_14223,N_7876,N_6927);
or U14224 (N_14224,N_6817,N_6775);
nand U14225 (N_14225,N_9124,N_7994);
nor U14226 (N_14226,N_9812,N_5784);
nand U14227 (N_14227,N_5751,N_6960);
or U14228 (N_14228,N_9066,N_8701);
and U14229 (N_14229,N_8789,N_6203);
or U14230 (N_14230,N_5779,N_6354);
nor U14231 (N_14231,N_5952,N_6696);
or U14232 (N_14232,N_5916,N_7186);
nor U14233 (N_14233,N_6082,N_8824);
and U14234 (N_14234,N_8119,N_5259);
or U14235 (N_14235,N_8489,N_9659);
nor U14236 (N_14236,N_6598,N_9946);
and U14237 (N_14237,N_8662,N_9337);
and U14238 (N_14238,N_5702,N_7703);
or U14239 (N_14239,N_8376,N_7112);
and U14240 (N_14240,N_5464,N_8648);
nor U14241 (N_14241,N_8971,N_7017);
nor U14242 (N_14242,N_9571,N_8686);
and U14243 (N_14243,N_7817,N_9683);
and U14244 (N_14244,N_8084,N_6854);
nor U14245 (N_14245,N_9142,N_8063);
nor U14246 (N_14246,N_7117,N_9728);
and U14247 (N_14247,N_8454,N_5091);
nor U14248 (N_14248,N_5979,N_7713);
nand U14249 (N_14249,N_6596,N_8963);
nor U14250 (N_14250,N_6438,N_7621);
or U14251 (N_14251,N_7148,N_8928);
nor U14252 (N_14252,N_8010,N_9793);
and U14253 (N_14253,N_9989,N_7868);
nand U14254 (N_14254,N_5077,N_9524);
nor U14255 (N_14255,N_7754,N_6291);
or U14256 (N_14256,N_5498,N_9571);
nor U14257 (N_14257,N_5553,N_9918);
and U14258 (N_14258,N_8534,N_6950);
and U14259 (N_14259,N_5346,N_7262);
nand U14260 (N_14260,N_8174,N_9654);
or U14261 (N_14261,N_7595,N_8135);
or U14262 (N_14262,N_9840,N_9348);
nor U14263 (N_14263,N_8405,N_5289);
nand U14264 (N_14264,N_5904,N_8560);
and U14265 (N_14265,N_5726,N_9891);
nor U14266 (N_14266,N_9869,N_8409);
and U14267 (N_14267,N_7316,N_9546);
and U14268 (N_14268,N_8518,N_8752);
and U14269 (N_14269,N_7330,N_5843);
nand U14270 (N_14270,N_7165,N_8839);
nor U14271 (N_14271,N_8174,N_7210);
nor U14272 (N_14272,N_8590,N_9210);
and U14273 (N_14273,N_7275,N_9858);
nand U14274 (N_14274,N_9730,N_6207);
or U14275 (N_14275,N_9581,N_8362);
nand U14276 (N_14276,N_8451,N_5065);
and U14277 (N_14277,N_6179,N_9096);
and U14278 (N_14278,N_9972,N_7054);
nor U14279 (N_14279,N_5512,N_7994);
nand U14280 (N_14280,N_6935,N_5591);
nor U14281 (N_14281,N_6737,N_5454);
nor U14282 (N_14282,N_6478,N_6702);
nor U14283 (N_14283,N_9289,N_9620);
nor U14284 (N_14284,N_5100,N_6369);
nand U14285 (N_14285,N_9864,N_5038);
nor U14286 (N_14286,N_9980,N_8145);
nor U14287 (N_14287,N_8765,N_5469);
nor U14288 (N_14288,N_9666,N_6648);
and U14289 (N_14289,N_6787,N_5545);
nor U14290 (N_14290,N_8087,N_9465);
and U14291 (N_14291,N_7829,N_7467);
and U14292 (N_14292,N_9659,N_6124);
nand U14293 (N_14293,N_7887,N_6679);
nor U14294 (N_14294,N_9847,N_8676);
xnor U14295 (N_14295,N_8166,N_5118);
or U14296 (N_14296,N_9571,N_8687);
nand U14297 (N_14297,N_9768,N_9674);
nand U14298 (N_14298,N_5338,N_7030);
or U14299 (N_14299,N_5308,N_7677);
and U14300 (N_14300,N_6610,N_9757);
nand U14301 (N_14301,N_8854,N_6443);
nor U14302 (N_14302,N_8029,N_8670);
or U14303 (N_14303,N_6738,N_6376);
nand U14304 (N_14304,N_6748,N_5466);
nand U14305 (N_14305,N_8335,N_6030);
and U14306 (N_14306,N_5393,N_5218);
or U14307 (N_14307,N_8280,N_5282);
or U14308 (N_14308,N_9247,N_7600);
nand U14309 (N_14309,N_6293,N_8265);
or U14310 (N_14310,N_5650,N_6656);
and U14311 (N_14311,N_7813,N_8042);
or U14312 (N_14312,N_9349,N_5069);
xor U14313 (N_14313,N_7189,N_9798);
nor U14314 (N_14314,N_9968,N_8893);
or U14315 (N_14315,N_8738,N_5834);
and U14316 (N_14316,N_7414,N_9864);
and U14317 (N_14317,N_7764,N_5215);
or U14318 (N_14318,N_6709,N_9272);
and U14319 (N_14319,N_6793,N_6125);
or U14320 (N_14320,N_8730,N_9246);
and U14321 (N_14321,N_9951,N_6443);
and U14322 (N_14322,N_8140,N_8874);
nor U14323 (N_14323,N_6795,N_5717);
nor U14324 (N_14324,N_8046,N_8165);
and U14325 (N_14325,N_7138,N_7671);
or U14326 (N_14326,N_8125,N_8351);
nor U14327 (N_14327,N_6415,N_7991);
xnor U14328 (N_14328,N_9204,N_9959);
nand U14329 (N_14329,N_8605,N_8598);
xor U14330 (N_14330,N_5364,N_6800);
nand U14331 (N_14331,N_6282,N_5788);
and U14332 (N_14332,N_8357,N_8941);
or U14333 (N_14333,N_6508,N_7966);
nor U14334 (N_14334,N_9510,N_9570);
nor U14335 (N_14335,N_9209,N_5182);
nand U14336 (N_14336,N_8123,N_8897);
or U14337 (N_14337,N_8157,N_7182);
or U14338 (N_14338,N_7497,N_8313);
nor U14339 (N_14339,N_5931,N_6947);
or U14340 (N_14340,N_9357,N_9382);
nor U14341 (N_14341,N_7394,N_8486);
nand U14342 (N_14342,N_8006,N_5755);
nor U14343 (N_14343,N_5719,N_6686);
nand U14344 (N_14344,N_7817,N_9678);
nand U14345 (N_14345,N_9256,N_9933);
nor U14346 (N_14346,N_8558,N_8258);
nor U14347 (N_14347,N_9321,N_8609);
nor U14348 (N_14348,N_6332,N_9111);
nor U14349 (N_14349,N_8494,N_7273);
nand U14350 (N_14350,N_6935,N_9547);
nor U14351 (N_14351,N_9211,N_8610);
and U14352 (N_14352,N_5471,N_6732);
or U14353 (N_14353,N_6765,N_6439);
nor U14354 (N_14354,N_6916,N_8243);
and U14355 (N_14355,N_7097,N_8691);
nand U14356 (N_14356,N_8411,N_8449);
nor U14357 (N_14357,N_9256,N_7085);
nor U14358 (N_14358,N_9541,N_7696);
nor U14359 (N_14359,N_9287,N_6332);
nand U14360 (N_14360,N_5398,N_8956);
nor U14361 (N_14361,N_8575,N_6808);
or U14362 (N_14362,N_9955,N_5676);
nor U14363 (N_14363,N_8281,N_9902);
or U14364 (N_14364,N_5965,N_7707);
or U14365 (N_14365,N_7407,N_6087);
nor U14366 (N_14366,N_5630,N_9568);
nand U14367 (N_14367,N_7860,N_8813);
nor U14368 (N_14368,N_5668,N_6018);
and U14369 (N_14369,N_6088,N_8624);
and U14370 (N_14370,N_8926,N_9883);
nor U14371 (N_14371,N_6375,N_5593);
or U14372 (N_14372,N_7542,N_7126);
or U14373 (N_14373,N_9260,N_5871);
and U14374 (N_14374,N_6418,N_5559);
and U14375 (N_14375,N_5548,N_8265);
nor U14376 (N_14376,N_5805,N_9663);
or U14377 (N_14377,N_6777,N_7060);
nor U14378 (N_14378,N_6500,N_9880);
or U14379 (N_14379,N_6030,N_5962);
nand U14380 (N_14380,N_5955,N_7718);
and U14381 (N_14381,N_7227,N_6910);
and U14382 (N_14382,N_7743,N_9868);
or U14383 (N_14383,N_9981,N_7370);
or U14384 (N_14384,N_9046,N_7516);
nand U14385 (N_14385,N_8652,N_8201);
or U14386 (N_14386,N_9043,N_7467);
and U14387 (N_14387,N_5470,N_8242);
nand U14388 (N_14388,N_5519,N_7389);
or U14389 (N_14389,N_7099,N_8101);
nor U14390 (N_14390,N_5065,N_6086);
or U14391 (N_14391,N_8786,N_8245);
or U14392 (N_14392,N_8993,N_7878);
or U14393 (N_14393,N_9870,N_8137);
nor U14394 (N_14394,N_9172,N_9351);
nand U14395 (N_14395,N_7740,N_5204);
nand U14396 (N_14396,N_8205,N_8790);
nor U14397 (N_14397,N_5768,N_5940);
nand U14398 (N_14398,N_6060,N_5406);
and U14399 (N_14399,N_7103,N_7085);
xnor U14400 (N_14400,N_7733,N_9572);
nor U14401 (N_14401,N_7692,N_9957);
nor U14402 (N_14402,N_8562,N_9561);
and U14403 (N_14403,N_5345,N_8070);
and U14404 (N_14404,N_7936,N_9368);
or U14405 (N_14405,N_7597,N_6780);
nand U14406 (N_14406,N_9501,N_8968);
or U14407 (N_14407,N_5854,N_5206);
nand U14408 (N_14408,N_7586,N_8315);
or U14409 (N_14409,N_9442,N_8976);
nor U14410 (N_14410,N_6912,N_5402);
nor U14411 (N_14411,N_6732,N_6412);
and U14412 (N_14412,N_6128,N_8231);
or U14413 (N_14413,N_5761,N_6572);
nand U14414 (N_14414,N_7950,N_8348);
or U14415 (N_14415,N_6857,N_9643);
nor U14416 (N_14416,N_9968,N_6734);
and U14417 (N_14417,N_8694,N_7435);
and U14418 (N_14418,N_9119,N_9115);
or U14419 (N_14419,N_9820,N_7779);
nor U14420 (N_14420,N_6853,N_9739);
or U14421 (N_14421,N_6675,N_8166);
nor U14422 (N_14422,N_7719,N_5207);
or U14423 (N_14423,N_8819,N_7786);
nor U14424 (N_14424,N_8715,N_9299);
and U14425 (N_14425,N_8520,N_8767);
xnor U14426 (N_14426,N_6087,N_9608);
nor U14427 (N_14427,N_6423,N_8132);
and U14428 (N_14428,N_6337,N_8291);
and U14429 (N_14429,N_9429,N_8367);
or U14430 (N_14430,N_7731,N_5957);
and U14431 (N_14431,N_8628,N_5049);
nor U14432 (N_14432,N_7539,N_7029);
or U14433 (N_14433,N_7194,N_5534);
nor U14434 (N_14434,N_9743,N_6810);
nand U14435 (N_14435,N_7641,N_9520);
and U14436 (N_14436,N_7021,N_8207);
or U14437 (N_14437,N_7969,N_9630);
or U14438 (N_14438,N_8264,N_6863);
nor U14439 (N_14439,N_5636,N_6596);
and U14440 (N_14440,N_6852,N_8318);
or U14441 (N_14441,N_8604,N_5429);
nand U14442 (N_14442,N_8101,N_7102);
nor U14443 (N_14443,N_9417,N_8570);
nand U14444 (N_14444,N_7068,N_5938);
or U14445 (N_14445,N_8999,N_9805);
nor U14446 (N_14446,N_6814,N_9475);
or U14447 (N_14447,N_9588,N_8346);
and U14448 (N_14448,N_9200,N_8793);
and U14449 (N_14449,N_7705,N_5856);
nand U14450 (N_14450,N_7011,N_9014);
or U14451 (N_14451,N_8091,N_8074);
or U14452 (N_14452,N_7501,N_7188);
nor U14453 (N_14453,N_6844,N_5527);
and U14454 (N_14454,N_8701,N_6632);
or U14455 (N_14455,N_8079,N_6996);
or U14456 (N_14456,N_9003,N_7168);
and U14457 (N_14457,N_9487,N_5893);
nor U14458 (N_14458,N_6266,N_8452);
or U14459 (N_14459,N_5400,N_6149);
xnor U14460 (N_14460,N_7413,N_6303);
nor U14461 (N_14461,N_8276,N_7247);
nor U14462 (N_14462,N_9009,N_8084);
or U14463 (N_14463,N_7800,N_7959);
and U14464 (N_14464,N_7668,N_8243);
or U14465 (N_14465,N_7911,N_9902);
and U14466 (N_14466,N_5788,N_8242);
nand U14467 (N_14467,N_5861,N_5905);
nor U14468 (N_14468,N_6067,N_5520);
nor U14469 (N_14469,N_6726,N_6082);
nor U14470 (N_14470,N_8333,N_8745);
or U14471 (N_14471,N_5953,N_9304);
or U14472 (N_14472,N_9787,N_6755);
nand U14473 (N_14473,N_6531,N_6984);
nor U14474 (N_14474,N_7781,N_9903);
nand U14475 (N_14475,N_6095,N_9565);
and U14476 (N_14476,N_9402,N_6403);
or U14477 (N_14477,N_9345,N_9275);
nor U14478 (N_14478,N_8688,N_7240);
and U14479 (N_14479,N_5215,N_9552);
nor U14480 (N_14480,N_8975,N_6802);
nand U14481 (N_14481,N_8855,N_5139);
or U14482 (N_14482,N_8177,N_6875);
xor U14483 (N_14483,N_8243,N_8917);
nor U14484 (N_14484,N_9749,N_5348);
nand U14485 (N_14485,N_5014,N_7949);
nor U14486 (N_14486,N_9021,N_5163);
and U14487 (N_14487,N_8362,N_6016);
nor U14488 (N_14488,N_6973,N_5946);
nand U14489 (N_14489,N_5801,N_7871);
and U14490 (N_14490,N_6536,N_8765);
or U14491 (N_14491,N_6145,N_8316);
nand U14492 (N_14492,N_5031,N_5864);
or U14493 (N_14493,N_8304,N_5732);
nand U14494 (N_14494,N_6546,N_7187);
nor U14495 (N_14495,N_5266,N_6343);
nor U14496 (N_14496,N_5737,N_9100);
and U14497 (N_14497,N_8990,N_8031);
or U14498 (N_14498,N_6827,N_9377);
or U14499 (N_14499,N_5626,N_9461);
or U14500 (N_14500,N_6894,N_5559);
or U14501 (N_14501,N_8458,N_9891);
nor U14502 (N_14502,N_9513,N_7904);
nor U14503 (N_14503,N_8752,N_7141);
or U14504 (N_14504,N_7718,N_9622);
nor U14505 (N_14505,N_5950,N_6609);
or U14506 (N_14506,N_6955,N_5602);
and U14507 (N_14507,N_7314,N_5967);
nand U14508 (N_14508,N_5816,N_7802);
nor U14509 (N_14509,N_9307,N_7424);
and U14510 (N_14510,N_8369,N_7491);
and U14511 (N_14511,N_6753,N_8559);
and U14512 (N_14512,N_8118,N_7751);
or U14513 (N_14513,N_7183,N_5963);
nand U14514 (N_14514,N_8529,N_6057);
and U14515 (N_14515,N_9654,N_8510);
and U14516 (N_14516,N_5881,N_5789);
nor U14517 (N_14517,N_5342,N_9338);
nor U14518 (N_14518,N_8650,N_6536);
and U14519 (N_14519,N_8156,N_9160);
nor U14520 (N_14520,N_5278,N_8829);
nand U14521 (N_14521,N_7232,N_5786);
nand U14522 (N_14522,N_7342,N_5099);
or U14523 (N_14523,N_9580,N_6745);
xnor U14524 (N_14524,N_5990,N_5221);
nand U14525 (N_14525,N_9788,N_8209);
nand U14526 (N_14526,N_5394,N_8217);
nand U14527 (N_14527,N_6708,N_6106);
nand U14528 (N_14528,N_5016,N_5392);
nand U14529 (N_14529,N_7313,N_9934);
and U14530 (N_14530,N_9905,N_8590);
or U14531 (N_14531,N_7547,N_7020);
and U14532 (N_14532,N_6891,N_5400);
or U14533 (N_14533,N_9440,N_5163);
xor U14534 (N_14534,N_6124,N_8630);
and U14535 (N_14535,N_9571,N_6314);
nor U14536 (N_14536,N_5324,N_6390);
or U14537 (N_14537,N_9720,N_5394);
or U14538 (N_14538,N_6321,N_9639);
nor U14539 (N_14539,N_6721,N_5722);
or U14540 (N_14540,N_8837,N_8337);
nand U14541 (N_14541,N_5411,N_8367);
and U14542 (N_14542,N_6029,N_8141);
or U14543 (N_14543,N_6480,N_9720);
nor U14544 (N_14544,N_6546,N_9606);
or U14545 (N_14545,N_9839,N_7116);
and U14546 (N_14546,N_5711,N_5485);
and U14547 (N_14547,N_5711,N_9355);
or U14548 (N_14548,N_5529,N_5632);
and U14549 (N_14549,N_7184,N_9915);
or U14550 (N_14550,N_8199,N_8102);
nor U14551 (N_14551,N_9309,N_6328);
or U14552 (N_14552,N_9817,N_6247);
nand U14553 (N_14553,N_9526,N_7766);
or U14554 (N_14554,N_7947,N_5687);
nand U14555 (N_14555,N_5924,N_5795);
or U14556 (N_14556,N_6078,N_5674);
nand U14557 (N_14557,N_8428,N_6770);
and U14558 (N_14558,N_6930,N_6782);
and U14559 (N_14559,N_8624,N_7224);
nor U14560 (N_14560,N_6205,N_6911);
nor U14561 (N_14561,N_8470,N_9600);
nand U14562 (N_14562,N_8704,N_8636);
or U14563 (N_14563,N_5710,N_8401);
xnor U14564 (N_14564,N_8392,N_7564);
nor U14565 (N_14565,N_7574,N_5930);
nor U14566 (N_14566,N_9419,N_6842);
and U14567 (N_14567,N_8898,N_7146);
and U14568 (N_14568,N_9289,N_6996);
xnor U14569 (N_14569,N_9747,N_5556);
or U14570 (N_14570,N_8589,N_8000);
nor U14571 (N_14571,N_8512,N_6264);
and U14572 (N_14572,N_8544,N_5926);
nand U14573 (N_14573,N_5858,N_9091);
nor U14574 (N_14574,N_5568,N_9572);
nand U14575 (N_14575,N_6191,N_8171);
nor U14576 (N_14576,N_9152,N_5911);
nand U14577 (N_14577,N_6440,N_9720);
or U14578 (N_14578,N_6210,N_9620);
or U14579 (N_14579,N_6626,N_6116);
or U14580 (N_14580,N_6398,N_6870);
nand U14581 (N_14581,N_9134,N_7557);
or U14582 (N_14582,N_9616,N_7290);
nor U14583 (N_14583,N_5426,N_5268);
nor U14584 (N_14584,N_9058,N_8674);
nor U14585 (N_14585,N_8545,N_7111);
or U14586 (N_14586,N_7561,N_6570);
or U14587 (N_14587,N_5201,N_7632);
and U14588 (N_14588,N_6200,N_6066);
xnor U14589 (N_14589,N_9120,N_8306);
nor U14590 (N_14590,N_5607,N_7951);
nor U14591 (N_14591,N_9973,N_9381);
or U14592 (N_14592,N_7534,N_7860);
and U14593 (N_14593,N_7232,N_6179);
and U14594 (N_14594,N_6940,N_5693);
and U14595 (N_14595,N_8253,N_5411);
and U14596 (N_14596,N_7864,N_5772);
nor U14597 (N_14597,N_8700,N_6746);
nor U14598 (N_14598,N_8277,N_9599);
and U14599 (N_14599,N_9913,N_9364);
or U14600 (N_14600,N_6425,N_9275);
and U14601 (N_14601,N_8889,N_9565);
or U14602 (N_14602,N_8912,N_9711);
nand U14603 (N_14603,N_9741,N_6195);
and U14604 (N_14604,N_9745,N_5621);
nand U14605 (N_14605,N_8171,N_6196);
nand U14606 (N_14606,N_8476,N_8255);
or U14607 (N_14607,N_9518,N_9123);
or U14608 (N_14608,N_8081,N_5309);
and U14609 (N_14609,N_8802,N_6052);
and U14610 (N_14610,N_5967,N_5495);
xor U14611 (N_14611,N_9562,N_9677);
nor U14612 (N_14612,N_5779,N_5404);
or U14613 (N_14613,N_8143,N_8645);
xnor U14614 (N_14614,N_8310,N_7470);
nand U14615 (N_14615,N_7940,N_7306);
nor U14616 (N_14616,N_6708,N_7794);
or U14617 (N_14617,N_9898,N_9392);
and U14618 (N_14618,N_7471,N_9750);
nor U14619 (N_14619,N_6960,N_6083);
nor U14620 (N_14620,N_8350,N_5583);
or U14621 (N_14621,N_9481,N_8583);
or U14622 (N_14622,N_5417,N_6202);
and U14623 (N_14623,N_7749,N_5535);
xnor U14624 (N_14624,N_7083,N_9220);
nor U14625 (N_14625,N_8922,N_6905);
nand U14626 (N_14626,N_8679,N_8479);
or U14627 (N_14627,N_5025,N_6291);
nand U14628 (N_14628,N_7698,N_7786);
and U14629 (N_14629,N_9990,N_8517);
and U14630 (N_14630,N_6953,N_7399);
nor U14631 (N_14631,N_6283,N_6077);
or U14632 (N_14632,N_5862,N_5315);
and U14633 (N_14633,N_5116,N_6285);
and U14634 (N_14634,N_8072,N_7774);
and U14635 (N_14635,N_5196,N_8169);
nand U14636 (N_14636,N_6515,N_7768);
nor U14637 (N_14637,N_9498,N_7365);
nand U14638 (N_14638,N_5781,N_5912);
nand U14639 (N_14639,N_5994,N_6453);
or U14640 (N_14640,N_6570,N_6059);
or U14641 (N_14641,N_5971,N_7934);
nor U14642 (N_14642,N_9031,N_9525);
and U14643 (N_14643,N_8746,N_9724);
and U14644 (N_14644,N_7458,N_5161);
nand U14645 (N_14645,N_6488,N_7824);
and U14646 (N_14646,N_5576,N_9488);
nor U14647 (N_14647,N_8745,N_6430);
nor U14648 (N_14648,N_7064,N_9375);
and U14649 (N_14649,N_6234,N_6181);
and U14650 (N_14650,N_9330,N_9012);
nand U14651 (N_14651,N_8579,N_9318);
or U14652 (N_14652,N_8138,N_9451);
nor U14653 (N_14653,N_5469,N_8433);
and U14654 (N_14654,N_7219,N_6272);
nand U14655 (N_14655,N_8245,N_5644);
xnor U14656 (N_14656,N_9010,N_6849);
and U14657 (N_14657,N_5045,N_8734);
nand U14658 (N_14658,N_8859,N_8767);
and U14659 (N_14659,N_5155,N_6210);
and U14660 (N_14660,N_7832,N_8414);
nand U14661 (N_14661,N_5875,N_6867);
or U14662 (N_14662,N_7456,N_8626);
nor U14663 (N_14663,N_6052,N_5131);
nand U14664 (N_14664,N_6379,N_6047);
nand U14665 (N_14665,N_8417,N_7356);
nor U14666 (N_14666,N_7329,N_9338);
nand U14667 (N_14667,N_7278,N_9395);
or U14668 (N_14668,N_8319,N_8427);
or U14669 (N_14669,N_5020,N_8664);
and U14670 (N_14670,N_6597,N_6933);
xor U14671 (N_14671,N_9529,N_8549);
nor U14672 (N_14672,N_5470,N_7918);
and U14673 (N_14673,N_9535,N_6195);
and U14674 (N_14674,N_8647,N_7526);
nand U14675 (N_14675,N_5156,N_8385);
or U14676 (N_14676,N_9344,N_5741);
nand U14677 (N_14677,N_6183,N_5136);
or U14678 (N_14678,N_9578,N_7955);
or U14679 (N_14679,N_8158,N_6175);
and U14680 (N_14680,N_6884,N_6513);
nor U14681 (N_14681,N_6461,N_7982);
nor U14682 (N_14682,N_5270,N_7628);
and U14683 (N_14683,N_5272,N_7873);
nor U14684 (N_14684,N_5965,N_9583);
and U14685 (N_14685,N_9619,N_5377);
or U14686 (N_14686,N_6707,N_5268);
nor U14687 (N_14687,N_8769,N_8070);
nand U14688 (N_14688,N_6921,N_7759);
nand U14689 (N_14689,N_5960,N_6965);
nor U14690 (N_14690,N_8731,N_5197);
or U14691 (N_14691,N_5683,N_8332);
and U14692 (N_14692,N_7483,N_7865);
nand U14693 (N_14693,N_9569,N_7965);
nand U14694 (N_14694,N_5514,N_5890);
nor U14695 (N_14695,N_9429,N_6260);
or U14696 (N_14696,N_5676,N_6220);
and U14697 (N_14697,N_7797,N_8076);
xor U14698 (N_14698,N_6318,N_9235);
xor U14699 (N_14699,N_6419,N_9064);
and U14700 (N_14700,N_5869,N_6010);
or U14701 (N_14701,N_8591,N_5177);
nand U14702 (N_14702,N_6919,N_5949);
nand U14703 (N_14703,N_8213,N_8784);
nand U14704 (N_14704,N_8247,N_8341);
or U14705 (N_14705,N_5196,N_8364);
or U14706 (N_14706,N_8413,N_6729);
or U14707 (N_14707,N_5234,N_6005);
and U14708 (N_14708,N_8939,N_6631);
or U14709 (N_14709,N_7299,N_5793);
nand U14710 (N_14710,N_6262,N_5759);
nand U14711 (N_14711,N_9408,N_5013);
or U14712 (N_14712,N_9790,N_8334);
and U14713 (N_14713,N_6639,N_7134);
nand U14714 (N_14714,N_7608,N_9678);
or U14715 (N_14715,N_9845,N_7130);
nand U14716 (N_14716,N_9218,N_7562);
nand U14717 (N_14717,N_7448,N_9357);
nand U14718 (N_14718,N_7866,N_5549);
nand U14719 (N_14719,N_7478,N_5050);
nor U14720 (N_14720,N_5361,N_6057);
nand U14721 (N_14721,N_7687,N_5764);
or U14722 (N_14722,N_7474,N_9363);
and U14723 (N_14723,N_9871,N_7562);
and U14724 (N_14724,N_9311,N_5925);
or U14725 (N_14725,N_8340,N_5785);
xnor U14726 (N_14726,N_8285,N_5918);
and U14727 (N_14727,N_8080,N_6883);
nor U14728 (N_14728,N_9045,N_9651);
or U14729 (N_14729,N_8789,N_9476);
and U14730 (N_14730,N_6302,N_6393);
or U14731 (N_14731,N_7167,N_7393);
nand U14732 (N_14732,N_7740,N_7691);
and U14733 (N_14733,N_6943,N_6287);
and U14734 (N_14734,N_7679,N_6724);
nor U14735 (N_14735,N_8364,N_6887);
or U14736 (N_14736,N_5805,N_9153);
or U14737 (N_14737,N_6046,N_5853);
and U14738 (N_14738,N_7641,N_6826);
or U14739 (N_14739,N_8618,N_5179);
nand U14740 (N_14740,N_8888,N_8741);
nor U14741 (N_14741,N_8089,N_6726);
nor U14742 (N_14742,N_9529,N_8067);
nor U14743 (N_14743,N_9179,N_8358);
nor U14744 (N_14744,N_6409,N_7086);
nor U14745 (N_14745,N_8714,N_7850);
nor U14746 (N_14746,N_8014,N_9551);
and U14747 (N_14747,N_7097,N_7589);
nand U14748 (N_14748,N_8249,N_7062);
nor U14749 (N_14749,N_7426,N_6362);
nor U14750 (N_14750,N_5681,N_6911);
or U14751 (N_14751,N_8703,N_5109);
and U14752 (N_14752,N_7063,N_5887);
nor U14753 (N_14753,N_5477,N_9022);
xor U14754 (N_14754,N_6956,N_9289);
or U14755 (N_14755,N_7116,N_6537);
nand U14756 (N_14756,N_8612,N_9354);
or U14757 (N_14757,N_5129,N_5508);
nand U14758 (N_14758,N_9974,N_8301);
xnor U14759 (N_14759,N_5295,N_6848);
nand U14760 (N_14760,N_7899,N_7757);
nor U14761 (N_14761,N_6629,N_7286);
or U14762 (N_14762,N_5361,N_5433);
and U14763 (N_14763,N_8437,N_9877);
and U14764 (N_14764,N_9975,N_6301);
and U14765 (N_14765,N_5906,N_5184);
nor U14766 (N_14766,N_6646,N_8813);
or U14767 (N_14767,N_7005,N_7623);
nand U14768 (N_14768,N_9318,N_6332);
and U14769 (N_14769,N_8910,N_7285);
and U14770 (N_14770,N_6622,N_9390);
and U14771 (N_14771,N_8430,N_8543);
and U14772 (N_14772,N_5466,N_5085);
nand U14773 (N_14773,N_7132,N_9918);
nor U14774 (N_14774,N_5311,N_6151);
and U14775 (N_14775,N_8611,N_9068);
and U14776 (N_14776,N_7906,N_9197);
and U14777 (N_14777,N_6985,N_5135);
and U14778 (N_14778,N_7908,N_9987);
nor U14779 (N_14779,N_5462,N_6780);
nor U14780 (N_14780,N_5104,N_9547);
and U14781 (N_14781,N_9245,N_6817);
and U14782 (N_14782,N_8478,N_9009);
xor U14783 (N_14783,N_8033,N_7115);
nor U14784 (N_14784,N_8895,N_9247);
and U14785 (N_14785,N_9383,N_6417);
nor U14786 (N_14786,N_5420,N_7245);
nand U14787 (N_14787,N_7832,N_7338);
nor U14788 (N_14788,N_9435,N_7351);
nand U14789 (N_14789,N_9273,N_7924);
and U14790 (N_14790,N_7787,N_7083);
and U14791 (N_14791,N_7411,N_6896);
nor U14792 (N_14792,N_9965,N_9946);
or U14793 (N_14793,N_6492,N_8873);
nor U14794 (N_14794,N_9641,N_5075);
nand U14795 (N_14795,N_5902,N_6569);
nand U14796 (N_14796,N_8107,N_9115);
and U14797 (N_14797,N_6149,N_5903);
nor U14798 (N_14798,N_8456,N_6304);
nor U14799 (N_14799,N_7844,N_9756);
and U14800 (N_14800,N_8383,N_6203);
nand U14801 (N_14801,N_9295,N_7649);
or U14802 (N_14802,N_5645,N_6179);
or U14803 (N_14803,N_9345,N_8448);
nand U14804 (N_14804,N_8311,N_8686);
nand U14805 (N_14805,N_9601,N_9091);
nand U14806 (N_14806,N_6823,N_6714);
nor U14807 (N_14807,N_8517,N_7136);
and U14808 (N_14808,N_9765,N_7481);
nor U14809 (N_14809,N_6670,N_5332);
and U14810 (N_14810,N_7262,N_6138);
nand U14811 (N_14811,N_7411,N_6937);
nand U14812 (N_14812,N_9879,N_7634);
nor U14813 (N_14813,N_9140,N_6237);
nor U14814 (N_14814,N_7917,N_9352);
and U14815 (N_14815,N_6295,N_6837);
or U14816 (N_14816,N_5265,N_5867);
nor U14817 (N_14817,N_8209,N_6019);
nor U14818 (N_14818,N_7984,N_7332);
or U14819 (N_14819,N_6597,N_9143);
nand U14820 (N_14820,N_8925,N_8936);
nor U14821 (N_14821,N_9508,N_5377);
and U14822 (N_14822,N_6589,N_9778);
nor U14823 (N_14823,N_8518,N_5127);
xor U14824 (N_14824,N_7013,N_7557);
and U14825 (N_14825,N_7789,N_6700);
xor U14826 (N_14826,N_9518,N_5883);
and U14827 (N_14827,N_8758,N_6076);
nand U14828 (N_14828,N_8905,N_9825);
nand U14829 (N_14829,N_9352,N_6459);
nor U14830 (N_14830,N_6826,N_6843);
nor U14831 (N_14831,N_9977,N_9457);
nor U14832 (N_14832,N_8002,N_8302);
nand U14833 (N_14833,N_9042,N_7211);
or U14834 (N_14834,N_7901,N_7380);
and U14835 (N_14835,N_8290,N_9781);
nor U14836 (N_14836,N_5884,N_6877);
nor U14837 (N_14837,N_7799,N_9034);
and U14838 (N_14838,N_9514,N_7359);
nand U14839 (N_14839,N_5551,N_6663);
or U14840 (N_14840,N_6506,N_6005);
nand U14841 (N_14841,N_8288,N_6036);
or U14842 (N_14842,N_6454,N_8518);
and U14843 (N_14843,N_9149,N_5417);
and U14844 (N_14844,N_8788,N_9508);
or U14845 (N_14845,N_6824,N_8754);
nand U14846 (N_14846,N_9835,N_5405);
and U14847 (N_14847,N_8213,N_5704);
or U14848 (N_14848,N_7493,N_6018);
nor U14849 (N_14849,N_8316,N_7878);
nor U14850 (N_14850,N_5739,N_9663);
nand U14851 (N_14851,N_5763,N_6069);
or U14852 (N_14852,N_7073,N_7474);
or U14853 (N_14853,N_6308,N_7755);
and U14854 (N_14854,N_6751,N_9626);
and U14855 (N_14855,N_9996,N_6864);
and U14856 (N_14856,N_5971,N_5999);
nand U14857 (N_14857,N_7870,N_7416);
nor U14858 (N_14858,N_8339,N_8129);
nor U14859 (N_14859,N_5705,N_6015);
nand U14860 (N_14860,N_9865,N_8940);
nand U14861 (N_14861,N_8749,N_7567);
nor U14862 (N_14862,N_5163,N_9578);
nand U14863 (N_14863,N_6741,N_7673);
or U14864 (N_14864,N_6488,N_6066);
and U14865 (N_14865,N_8822,N_5930);
nand U14866 (N_14866,N_7122,N_8969);
nor U14867 (N_14867,N_8308,N_7952);
or U14868 (N_14868,N_8533,N_8197);
nor U14869 (N_14869,N_6963,N_6453);
xor U14870 (N_14870,N_6971,N_6084);
nand U14871 (N_14871,N_9850,N_6014);
or U14872 (N_14872,N_9739,N_5861);
or U14873 (N_14873,N_6084,N_7929);
nor U14874 (N_14874,N_5940,N_9829);
nand U14875 (N_14875,N_5342,N_9909);
and U14876 (N_14876,N_6293,N_8557);
or U14877 (N_14877,N_7353,N_8046);
or U14878 (N_14878,N_6464,N_6202);
and U14879 (N_14879,N_5663,N_7753);
nor U14880 (N_14880,N_8315,N_6596);
nor U14881 (N_14881,N_5143,N_7464);
nor U14882 (N_14882,N_9176,N_6873);
nor U14883 (N_14883,N_8237,N_5060);
or U14884 (N_14884,N_8069,N_8614);
and U14885 (N_14885,N_8910,N_9482);
nor U14886 (N_14886,N_9483,N_5779);
or U14887 (N_14887,N_5476,N_9674);
nor U14888 (N_14888,N_6851,N_6472);
or U14889 (N_14889,N_9175,N_9605);
or U14890 (N_14890,N_7606,N_8129);
nor U14891 (N_14891,N_5502,N_5560);
or U14892 (N_14892,N_7969,N_5464);
nand U14893 (N_14893,N_9090,N_7352);
nor U14894 (N_14894,N_7090,N_6290);
or U14895 (N_14895,N_8503,N_8180);
and U14896 (N_14896,N_5694,N_5665);
or U14897 (N_14897,N_8341,N_5702);
nor U14898 (N_14898,N_8918,N_9369);
nor U14899 (N_14899,N_8971,N_8306);
xor U14900 (N_14900,N_6754,N_6628);
nand U14901 (N_14901,N_9129,N_5456);
nand U14902 (N_14902,N_8318,N_8618);
or U14903 (N_14903,N_7375,N_5444);
nand U14904 (N_14904,N_7310,N_6664);
nor U14905 (N_14905,N_5529,N_7724);
nor U14906 (N_14906,N_6803,N_5674);
or U14907 (N_14907,N_7978,N_8714);
and U14908 (N_14908,N_9749,N_6839);
nand U14909 (N_14909,N_5820,N_7535);
nor U14910 (N_14910,N_6009,N_5033);
nor U14911 (N_14911,N_8055,N_6228);
or U14912 (N_14912,N_9901,N_8795);
and U14913 (N_14913,N_5175,N_6131);
and U14914 (N_14914,N_8761,N_7733);
nand U14915 (N_14915,N_9961,N_9909);
or U14916 (N_14916,N_7885,N_5485);
nand U14917 (N_14917,N_8349,N_5430);
and U14918 (N_14918,N_5525,N_6451);
and U14919 (N_14919,N_8296,N_7414);
nor U14920 (N_14920,N_8109,N_7265);
or U14921 (N_14921,N_5861,N_9055);
nand U14922 (N_14922,N_6481,N_9243);
and U14923 (N_14923,N_6148,N_7884);
nor U14924 (N_14924,N_8594,N_7551);
nand U14925 (N_14925,N_5233,N_6375);
nor U14926 (N_14926,N_9758,N_6032);
nand U14927 (N_14927,N_5695,N_9430);
xnor U14928 (N_14928,N_8698,N_9038);
or U14929 (N_14929,N_8817,N_7509);
and U14930 (N_14930,N_8186,N_8719);
and U14931 (N_14931,N_7454,N_5566);
nor U14932 (N_14932,N_7015,N_7173);
nor U14933 (N_14933,N_9145,N_5165);
nand U14934 (N_14934,N_7743,N_8733);
or U14935 (N_14935,N_7034,N_7406);
nor U14936 (N_14936,N_6075,N_6468);
or U14937 (N_14937,N_9998,N_5064);
nor U14938 (N_14938,N_5324,N_7740);
and U14939 (N_14939,N_7304,N_7594);
and U14940 (N_14940,N_5020,N_8999);
or U14941 (N_14941,N_9822,N_6774);
nor U14942 (N_14942,N_8158,N_8247);
nand U14943 (N_14943,N_6182,N_8321);
nor U14944 (N_14944,N_6433,N_6928);
nand U14945 (N_14945,N_7151,N_5590);
or U14946 (N_14946,N_9168,N_5490);
and U14947 (N_14947,N_7050,N_8557);
or U14948 (N_14948,N_6247,N_9033);
nor U14949 (N_14949,N_7541,N_5415);
nand U14950 (N_14950,N_6860,N_9585);
and U14951 (N_14951,N_6010,N_6769);
nor U14952 (N_14952,N_8959,N_6329);
and U14953 (N_14953,N_9877,N_8641);
or U14954 (N_14954,N_6302,N_5603);
and U14955 (N_14955,N_7924,N_6391);
and U14956 (N_14956,N_6392,N_6079);
nor U14957 (N_14957,N_5433,N_5990);
and U14958 (N_14958,N_5287,N_6742);
and U14959 (N_14959,N_9753,N_7940);
nand U14960 (N_14960,N_6784,N_5247);
nor U14961 (N_14961,N_9068,N_7056);
nor U14962 (N_14962,N_8595,N_8808);
nor U14963 (N_14963,N_5903,N_9018);
nand U14964 (N_14964,N_8838,N_9570);
nand U14965 (N_14965,N_7916,N_9958);
nand U14966 (N_14966,N_9309,N_5040);
nor U14967 (N_14967,N_5138,N_9018);
xnor U14968 (N_14968,N_6758,N_7494);
nand U14969 (N_14969,N_9841,N_6130);
nand U14970 (N_14970,N_6877,N_9244);
nand U14971 (N_14971,N_5227,N_5307);
or U14972 (N_14972,N_5270,N_9715);
nor U14973 (N_14973,N_8286,N_8653);
or U14974 (N_14974,N_8446,N_6962);
nand U14975 (N_14975,N_6962,N_7724);
and U14976 (N_14976,N_6673,N_8390);
and U14977 (N_14977,N_7813,N_9974);
or U14978 (N_14978,N_8983,N_7399);
or U14979 (N_14979,N_8331,N_6575);
or U14980 (N_14980,N_6613,N_6935);
or U14981 (N_14981,N_9127,N_6309);
xnor U14982 (N_14982,N_9385,N_5208);
or U14983 (N_14983,N_8438,N_8309);
nand U14984 (N_14984,N_6126,N_5663);
and U14985 (N_14985,N_6890,N_7795);
or U14986 (N_14986,N_9952,N_8412);
nor U14987 (N_14987,N_9484,N_8182);
and U14988 (N_14988,N_9137,N_7737);
nand U14989 (N_14989,N_9897,N_8976);
nor U14990 (N_14990,N_7501,N_9667);
or U14991 (N_14991,N_8311,N_8725);
or U14992 (N_14992,N_6104,N_5914);
nand U14993 (N_14993,N_7475,N_7898);
or U14994 (N_14994,N_9097,N_9828);
or U14995 (N_14995,N_7369,N_5868);
or U14996 (N_14996,N_7679,N_8839);
and U14997 (N_14997,N_8539,N_7008);
nand U14998 (N_14998,N_7221,N_8438);
xnor U14999 (N_14999,N_6667,N_5251);
or U15000 (N_15000,N_11963,N_12766);
or U15001 (N_15001,N_12185,N_12095);
and U15002 (N_15002,N_10432,N_13778);
and U15003 (N_15003,N_11496,N_13094);
xor U15004 (N_15004,N_13903,N_10901);
or U15005 (N_15005,N_10188,N_12067);
or U15006 (N_15006,N_10455,N_14040);
or U15007 (N_15007,N_10521,N_14257);
nand U15008 (N_15008,N_14229,N_10912);
and U15009 (N_15009,N_11951,N_11944);
or U15010 (N_15010,N_14647,N_14846);
or U15011 (N_15011,N_11250,N_12254);
or U15012 (N_15012,N_12860,N_10866);
nor U15013 (N_15013,N_14592,N_14021);
nand U15014 (N_15014,N_12042,N_14476);
and U15015 (N_15015,N_12794,N_13686);
and U15016 (N_15016,N_10559,N_10066);
nor U15017 (N_15017,N_12942,N_11643);
nor U15018 (N_15018,N_13419,N_13490);
or U15019 (N_15019,N_14253,N_11238);
xor U15020 (N_15020,N_13418,N_11519);
nand U15021 (N_15021,N_11403,N_10451);
nand U15022 (N_15022,N_10771,N_12366);
or U15023 (N_15023,N_13374,N_13351);
and U15024 (N_15024,N_12946,N_14435);
or U15025 (N_15025,N_14239,N_14748);
nor U15026 (N_15026,N_14161,N_13481);
or U15027 (N_15027,N_10716,N_14404);
and U15028 (N_15028,N_10080,N_11919);
nand U15029 (N_15029,N_14783,N_11443);
nor U15030 (N_15030,N_10693,N_13372);
or U15031 (N_15031,N_14993,N_13296);
xnor U15032 (N_15032,N_11954,N_11381);
nand U15033 (N_15033,N_10916,N_14262);
and U15034 (N_15034,N_13067,N_14817);
nand U15035 (N_15035,N_11349,N_12813);
and U15036 (N_15036,N_12575,N_12260);
or U15037 (N_15037,N_14156,N_12983);
or U15038 (N_15038,N_11716,N_13550);
and U15039 (N_15039,N_12805,N_13926);
nor U15040 (N_15040,N_10187,N_11074);
nor U15041 (N_15041,N_13641,N_13097);
and U15042 (N_15042,N_13442,N_12989);
nor U15043 (N_15043,N_12675,N_11147);
nand U15044 (N_15044,N_11423,N_14552);
nand U15045 (N_15045,N_11794,N_13913);
xnor U15046 (N_15046,N_13895,N_10090);
nor U15047 (N_15047,N_13518,N_12775);
nand U15048 (N_15048,N_12714,N_10851);
or U15049 (N_15049,N_10904,N_10788);
and U15050 (N_15050,N_14584,N_12374);
and U15051 (N_15051,N_14589,N_12189);
or U15052 (N_15052,N_10454,N_10342);
nand U15053 (N_15053,N_10838,N_12331);
nand U15054 (N_15054,N_13478,N_14216);
and U15055 (N_15055,N_11180,N_13405);
or U15056 (N_15056,N_10573,N_11620);
nor U15057 (N_15057,N_13533,N_12330);
and U15058 (N_15058,N_11137,N_10965);
or U15059 (N_15059,N_10744,N_12174);
nand U15060 (N_15060,N_11214,N_14692);
nand U15061 (N_15061,N_12621,N_10151);
or U15062 (N_15062,N_14325,N_12886);
and U15063 (N_15063,N_13431,N_11715);
nor U15064 (N_15064,N_10329,N_10500);
nand U15065 (N_15065,N_12633,N_11828);
and U15066 (N_15066,N_10355,N_14917);
nand U15067 (N_15067,N_10483,N_10259);
nor U15068 (N_15068,N_10294,N_12285);
nand U15069 (N_15069,N_13615,N_14649);
and U15070 (N_15070,N_14116,N_14859);
or U15071 (N_15071,N_12949,N_12565);
nor U15072 (N_15072,N_14000,N_11192);
or U15073 (N_15073,N_10150,N_10540);
nand U15074 (N_15074,N_13654,N_11590);
nand U15075 (N_15075,N_13681,N_11523);
nor U15076 (N_15076,N_14258,N_14309);
or U15077 (N_15077,N_10801,N_13127);
nand U15078 (N_15078,N_10073,N_10597);
nor U15079 (N_15079,N_14541,N_10932);
nand U15080 (N_15080,N_12716,N_10939);
nand U15081 (N_15081,N_14833,N_12554);
or U15082 (N_15082,N_11538,N_13295);
or U15083 (N_15083,N_11277,N_13639);
and U15084 (N_15084,N_13629,N_14891);
or U15085 (N_15085,N_13173,N_14168);
and U15086 (N_15086,N_11497,N_10522);
or U15087 (N_15087,N_12743,N_12239);
nand U15088 (N_15088,N_13217,N_10183);
and U15089 (N_15089,N_13355,N_10344);
or U15090 (N_15090,N_12881,N_14805);
and U15091 (N_15091,N_14678,N_13437);
or U15092 (N_15092,N_12078,N_13682);
and U15093 (N_15093,N_11167,N_12514);
or U15094 (N_15094,N_14458,N_10244);
or U15095 (N_15095,N_12157,N_11021);
and U15096 (N_15096,N_12650,N_10730);
or U15097 (N_15097,N_13027,N_10269);
and U15098 (N_15098,N_12995,N_11219);
and U15099 (N_15099,N_11713,N_13080);
xor U15100 (N_15100,N_10872,N_11553);
nor U15101 (N_15101,N_10669,N_12273);
or U15102 (N_15102,N_13354,N_10858);
nor U15103 (N_15103,N_13253,N_13875);
nor U15104 (N_15104,N_12441,N_14276);
nand U15105 (N_15105,N_13964,N_14611);
and U15106 (N_15106,N_10917,N_10778);
nand U15107 (N_15107,N_11097,N_14208);
nor U15108 (N_15108,N_11187,N_13118);
nand U15109 (N_15109,N_12102,N_10331);
nand U15110 (N_15110,N_14271,N_10144);
or U15111 (N_15111,N_14585,N_11695);
nand U15112 (N_15112,N_13218,N_11357);
and U15113 (N_15113,N_14619,N_13501);
nor U15114 (N_15114,N_14065,N_11048);
or U15115 (N_15115,N_13312,N_13940);
or U15116 (N_15116,N_11071,N_13346);
or U15117 (N_15117,N_14511,N_10889);
or U15118 (N_15118,N_13908,N_14631);
and U15119 (N_15119,N_13404,N_14010);
nand U15120 (N_15120,N_12215,N_11194);
and U15121 (N_15121,N_14071,N_14219);
nand U15122 (N_15122,N_13553,N_12403);
xnor U15123 (N_15123,N_11863,N_12390);
and U15124 (N_15124,N_11790,N_12868);
nand U15125 (N_15125,N_10781,N_14462);
nand U15126 (N_15126,N_12652,N_12092);
or U15127 (N_15127,N_14890,N_12883);
or U15128 (N_15128,N_10935,N_12384);
and U15129 (N_15129,N_10678,N_11022);
or U15130 (N_15130,N_11193,N_13901);
nor U15131 (N_15131,N_14154,N_14326);
nor U15132 (N_15132,N_14043,N_13017);
and U15133 (N_15133,N_14111,N_11545);
and U15134 (N_15134,N_14428,N_11310);
nand U15135 (N_15135,N_13379,N_14495);
nand U15136 (N_15136,N_12933,N_11366);
nand U15137 (N_15137,N_14132,N_12188);
nand U15138 (N_15138,N_13558,N_10464);
or U15139 (N_15139,N_10941,N_13304);
and U15140 (N_15140,N_14122,N_11121);
nor U15141 (N_15141,N_14670,N_14164);
or U15142 (N_15142,N_12319,N_12404);
nand U15143 (N_15143,N_14743,N_10083);
and U15144 (N_15144,N_14714,N_10079);
and U15145 (N_15145,N_13590,N_12753);
nor U15146 (N_15146,N_11678,N_12300);
nor U15147 (N_15147,N_14725,N_12550);
nand U15148 (N_15148,N_10088,N_13666);
or U15149 (N_15149,N_13849,N_12664);
or U15150 (N_15150,N_11294,N_14110);
and U15151 (N_15151,N_14041,N_11639);
and U15152 (N_15152,N_10829,N_10366);
nor U15153 (N_15153,N_11400,N_13636);
nor U15154 (N_15154,N_11166,N_14706);
nor U15155 (N_15155,N_12169,N_11049);
nor U15156 (N_15156,N_13147,N_12894);
nand U15157 (N_15157,N_14615,N_12286);
and U15158 (N_15158,N_11897,N_10425);
and U15159 (N_15159,N_11099,N_14583);
or U15160 (N_15160,N_14144,N_12712);
nand U15161 (N_15161,N_11059,N_11693);
nor U15162 (N_15162,N_14823,N_12064);
and U15163 (N_15163,N_14701,N_13890);
and U15164 (N_15164,N_10395,N_13795);
nand U15165 (N_15165,N_10056,N_12419);
nor U15166 (N_15166,N_10240,N_13115);
nand U15167 (N_15167,N_11637,N_10074);
nand U15168 (N_15168,N_12569,N_10779);
nand U15169 (N_15169,N_10867,N_12443);
nor U15170 (N_15170,N_10427,N_11182);
or U15171 (N_15171,N_11664,N_14259);
and U15172 (N_15172,N_12503,N_11632);
and U15173 (N_15173,N_12896,N_12435);
nor U15174 (N_15174,N_14475,N_14245);
or U15175 (N_15175,N_14512,N_14183);
and U15176 (N_15176,N_10591,N_13240);
or U15177 (N_15177,N_10270,N_14313);
nand U15178 (N_15178,N_10969,N_11125);
nor U15179 (N_15179,N_12468,N_11660);
and U15180 (N_15180,N_10845,N_12681);
nand U15181 (N_15181,N_13283,N_10286);
nand U15182 (N_15182,N_14365,N_10566);
and U15183 (N_15183,N_11265,N_12504);
nand U15184 (N_15184,N_13063,N_14738);
and U15185 (N_15185,N_14553,N_12402);
and U15186 (N_15186,N_11718,N_11318);
and U15187 (N_15187,N_13341,N_12464);
nor U15188 (N_15188,N_11183,N_11613);
or U15189 (N_15189,N_13994,N_11737);
nor U15190 (N_15190,N_12969,N_11405);
nor U15191 (N_15191,N_14436,N_13934);
or U15192 (N_15192,N_10707,N_13579);
and U15193 (N_15193,N_14503,N_10646);
nor U15194 (N_15194,N_13664,N_10158);
and U15195 (N_15195,N_14836,N_14414);
and U15196 (N_15196,N_12201,N_11406);
and U15197 (N_15197,N_12352,N_11110);
nor U15198 (N_15198,N_11775,N_12270);
or U15199 (N_15199,N_12000,N_11898);
and U15200 (N_15200,N_11766,N_12426);
and U15201 (N_15201,N_13053,N_12884);
nand U15202 (N_15202,N_12072,N_12658);
or U15203 (N_15203,N_12710,N_10061);
and U15204 (N_15204,N_10319,N_14078);
or U15205 (N_15205,N_12872,N_11745);
and U15206 (N_15206,N_13648,N_13715);
or U15207 (N_15207,N_14928,N_10039);
and U15208 (N_15208,N_10385,N_10775);
or U15209 (N_15209,N_14662,N_13110);
and U15210 (N_15210,N_11453,N_12740);
nand U15211 (N_15211,N_12774,N_14347);
nand U15212 (N_15212,N_10304,N_13035);
nor U15213 (N_15213,N_14375,N_13894);
nand U15214 (N_15214,N_12773,N_12516);
or U15215 (N_15215,N_10834,N_12857);
xnor U15216 (N_15216,N_13560,N_14599);
nor U15217 (N_15217,N_12945,N_10589);
nand U15218 (N_15218,N_10992,N_12928);
and U15219 (N_15219,N_12120,N_10252);
nand U15220 (N_15220,N_11699,N_11033);
or U15221 (N_15221,N_11704,N_14205);
and U15222 (N_15222,N_13669,N_10810);
or U15223 (N_15223,N_12071,N_10870);
nand U15224 (N_15224,N_13181,N_10453);
or U15225 (N_15225,N_11055,N_11656);
and U15226 (N_15226,N_11384,N_11966);
or U15227 (N_15227,N_10795,N_13897);
nor U15228 (N_15228,N_14453,N_10792);
and U15229 (N_15229,N_14389,N_12321);
or U15230 (N_15230,N_11311,N_13876);
nor U15231 (N_15231,N_10293,N_13852);
nand U15232 (N_15232,N_12485,N_14731);
and U15233 (N_15233,N_12738,N_10207);
nor U15234 (N_15234,N_10607,N_10980);
nor U15235 (N_15235,N_10816,N_13893);
nand U15236 (N_15236,N_14422,N_14286);
and U15237 (N_15237,N_14001,N_11540);
nor U15238 (N_15238,N_10112,N_12973);
nor U15239 (N_15239,N_11007,N_14391);
and U15240 (N_15240,N_13251,N_10025);
nand U15241 (N_15241,N_11968,N_11600);
or U15242 (N_15242,N_11874,N_13220);
nand U15243 (N_15243,N_13289,N_12373);
xor U15244 (N_15244,N_10605,N_11563);
or U15245 (N_15245,N_11139,N_11090);
and U15246 (N_15246,N_12132,N_14782);
nor U15247 (N_15247,N_14038,N_14763);
nor U15248 (N_15248,N_11953,N_14328);
or U15249 (N_15249,N_14430,N_11106);
nand U15250 (N_15250,N_13366,N_10362);
nand U15251 (N_15251,N_13642,N_11128);
or U15252 (N_15252,N_12627,N_10557);
nor U15253 (N_15253,N_11950,N_14268);
nand U15254 (N_15254,N_13935,N_12493);
or U15255 (N_15255,N_12326,N_12608);
nand U15256 (N_15256,N_10403,N_14096);
or U15257 (N_15257,N_10755,N_10960);
or U15258 (N_15258,N_10302,N_12168);
and U15259 (N_15259,N_11235,N_10296);
nor U15260 (N_15260,N_14489,N_14514);
nand U15261 (N_15261,N_11358,N_10449);
nor U15262 (N_15262,N_14753,N_14023);
nor U15263 (N_15263,N_10840,N_11293);
nand U15264 (N_15264,N_13002,N_13523);
or U15265 (N_15265,N_11959,N_10919);
or U15266 (N_15266,N_14955,N_10223);
and U15267 (N_15267,N_10414,N_12180);
or U15268 (N_15268,N_11998,N_14883);
xor U15269 (N_15269,N_14233,N_10898);
xnor U15270 (N_15270,N_13505,N_10624);
or U15271 (N_15271,N_11515,N_10632);
nand U15272 (N_15272,N_13272,N_10814);
or U15273 (N_15273,N_14146,N_12291);
nand U15274 (N_15274,N_13618,N_12039);
or U15275 (N_15275,N_10488,N_12127);
xnor U15276 (N_15276,N_12899,N_14620);
nor U15277 (N_15277,N_13631,N_10094);
and U15278 (N_15278,N_10283,N_12372);
nand U15279 (N_15279,N_14267,N_11645);
or U15280 (N_15280,N_11368,N_14314);
and U15281 (N_15281,N_12557,N_12737);
and U15282 (N_15282,N_10552,N_13252);
and U15283 (N_15283,N_13224,N_12361);
or U15284 (N_15284,N_14440,N_10794);
or U15285 (N_15285,N_13765,N_10239);
nor U15286 (N_15286,N_13064,N_13473);
nand U15287 (N_15287,N_13772,N_14897);
and U15288 (N_15288,N_11113,N_10208);
nor U15289 (N_15289,N_14801,N_12564);
or U15290 (N_15290,N_13136,N_13983);
nand U15291 (N_15291,N_14171,N_12453);
nand U15292 (N_15292,N_13273,N_12387);
nand U15293 (N_15293,N_14965,N_13278);
nor U15294 (N_15294,N_12205,N_13541);
nand U15295 (N_15295,N_13241,N_11041);
or U15296 (N_15296,N_12267,N_11323);
xnor U15297 (N_15297,N_13925,N_12531);
or U15298 (N_15298,N_13454,N_13160);
nand U15299 (N_15299,N_12505,N_13867);
or U15300 (N_15300,N_13122,N_10837);
and U15301 (N_15301,N_13172,N_14998);
and U15302 (N_15302,N_11741,N_11485);
or U15303 (N_15303,N_12880,N_10620);
xnor U15304 (N_15304,N_10175,N_13169);
and U15305 (N_15305,N_11578,N_12873);
nor U15306 (N_15306,N_11031,N_14691);
nand U15307 (N_15307,N_10790,N_13259);
nand U15308 (N_15308,N_11539,N_12948);
and U15309 (N_15309,N_13754,N_10234);
nor U15310 (N_15310,N_13905,N_11252);
nor U15311 (N_15311,N_14720,N_10878);
xor U15312 (N_15312,N_10146,N_10527);
nor U15313 (N_15313,N_11602,N_10676);
or U15314 (N_15314,N_13076,N_12467);
nor U15315 (N_15315,N_11160,N_11258);
or U15316 (N_15316,N_10653,N_10558);
nor U15317 (N_15317,N_11224,N_13318);
and U15318 (N_15318,N_10871,N_14047);
nand U15319 (N_15319,N_13095,N_14169);
and U15320 (N_15320,N_13347,N_12047);
nand U15321 (N_15321,N_13081,N_13577);
and U15322 (N_15322,N_14613,N_12902);
and U15323 (N_15323,N_13958,N_13892);
or U15324 (N_15324,N_13924,N_11978);
nor U15325 (N_15325,N_10312,N_12457);
nor U15326 (N_15326,N_14341,N_11216);
xor U15327 (N_15327,N_12228,N_11326);
and U15328 (N_15328,N_13663,N_12034);
or U15329 (N_15329,N_11475,N_13909);
and U15330 (N_15330,N_14996,N_13422);
nand U15331 (N_15331,N_12898,N_10906);
nor U15332 (N_15332,N_14186,N_10346);
nor U15333 (N_15333,N_10567,N_14492);
and U15334 (N_15334,N_12206,N_13254);
nor U15335 (N_15335,N_13691,N_13000);
and U15336 (N_15336,N_10382,N_14627);
or U15337 (N_15337,N_13495,N_10934);
nand U15338 (N_15338,N_12576,N_14191);
nand U15339 (N_15339,N_11478,N_14634);
or U15340 (N_15340,N_11824,N_13256);
and U15341 (N_15341,N_13712,N_12281);
xnor U15342 (N_15342,N_10347,N_10574);
nand U15343 (N_15343,N_12012,N_13670);
and U15344 (N_15344,N_14401,N_12250);
nor U15345 (N_15345,N_11548,N_11474);
or U15346 (N_15346,N_11616,N_10937);
nand U15347 (N_15347,N_11859,N_14166);
nor U15348 (N_15348,N_11719,N_10373);
and U15349 (N_15349,N_11787,N_13689);
and U15350 (N_15350,N_14415,N_11179);
nor U15351 (N_15351,N_11499,N_14768);
nor U15352 (N_15352,N_14074,N_14352);
or U15353 (N_15353,N_13697,N_14354);
nand U15354 (N_15354,N_11388,N_14056);
or U15355 (N_15355,N_14222,N_11208);
and U15356 (N_15356,N_10446,N_10374);
or U15357 (N_15357,N_11864,N_11518);
or U15358 (N_15358,N_14560,N_13604);
and U15359 (N_15359,N_12213,N_13554);
nand U15360 (N_15360,N_11512,N_11914);
nor U15361 (N_15361,N_14604,N_13015);
and U15362 (N_15362,N_10272,N_11972);
nor U15363 (N_15363,N_11995,N_14220);
xor U15364 (N_15364,N_11758,N_12887);
nor U15365 (N_15365,N_11034,N_11291);
or U15366 (N_15366,N_14903,N_10448);
and U15367 (N_15367,N_12466,N_14451);
or U15368 (N_15368,N_13592,N_10593);
or U15369 (N_15369,N_14162,N_12110);
and U15370 (N_15370,N_13919,N_10823);
nand U15371 (N_15371,N_10193,N_14598);
nand U15372 (N_15372,N_12397,N_14247);
nor U15373 (N_15373,N_14690,N_10751);
and U15374 (N_15374,N_12770,N_14573);
or U15375 (N_15375,N_13622,N_11267);
and U15376 (N_15376,N_11196,N_12121);
or U15377 (N_15377,N_11671,N_12629);
nand U15378 (N_15378,N_11749,N_10128);
and U15379 (N_15379,N_10824,N_13555);
or U15380 (N_15380,N_11687,N_12323);
xor U15381 (N_15381,N_14134,N_12606);
and U15382 (N_15382,N_11594,N_12107);
nor U15383 (N_15383,N_10804,N_13507);
nor U15384 (N_15384,N_10267,N_10445);
nor U15385 (N_15385,N_11390,N_13825);
nor U15386 (N_15386,N_13003,N_11644);
or U15387 (N_15387,N_12670,N_12549);
and U15388 (N_15388,N_14024,N_14515);
nor U15389 (N_15389,N_14656,N_13265);
nor U15390 (N_15390,N_14697,N_10245);
nand U15391 (N_15391,N_13588,N_14209);
nand U15392 (N_15392,N_13263,N_14042);
and U15393 (N_15393,N_14032,N_11047);
and U15394 (N_15394,N_11136,N_12358);
nand U15395 (N_15395,N_14105,N_14048);
and U15396 (N_15396,N_10159,N_11469);
nand U15397 (N_15397,N_13415,N_11338);
nand U15398 (N_15398,N_13452,N_10876);
nor U15399 (N_15399,N_14084,N_11501);
or U15400 (N_15400,N_12878,N_12261);
and U15401 (N_15401,N_10882,N_11852);
nor U15402 (N_15402,N_10990,N_14360);
nand U15403 (N_15403,N_10058,N_12046);
nand U15404 (N_15404,N_10981,N_14223);
or U15405 (N_15405,N_12226,N_12312);
nand U15406 (N_15406,N_11391,N_10152);
nor U15407 (N_15407,N_10623,N_14735);
and U15408 (N_15408,N_11920,N_11712);
nand U15409 (N_15409,N_12561,N_10043);
nand U15410 (N_15410,N_10023,N_10135);
nor U15411 (N_15411,N_13717,N_11989);
nand U15412 (N_15412,N_13491,N_14848);
and U15413 (N_15413,N_14128,N_10137);
nand U15414 (N_15414,N_10466,N_13159);
or U15415 (N_15415,N_14063,N_10408);
and U15416 (N_15416,N_10098,N_13634);
nand U15417 (N_15417,N_10952,N_10474);
nor U15418 (N_15418,N_13839,N_10450);
nand U15419 (N_15419,N_12314,N_10631);
nand U15420 (N_15420,N_14305,N_11581);
and U15421 (N_15421,N_11230,N_12771);
nor U15422 (N_15422,N_12377,N_12746);
nand U15423 (N_15423,N_11408,N_12028);
or U15424 (N_15424,N_14264,N_13292);
and U15425 (N_15425,N_13793,N_14590);
and U15426 (N_15426,N_12170,N_11268);
nand U15427 (N_15427,N_11170,N_10011);
and U15428 (N_15428,N_12761,N_10734);
and U15429 (N_15429,N_11426,N_12547);
and U15430 (N_15430,N_13291,N_13863);
nor U15431 (N_15431,N_10599,N_12425);
nand U15432 (N_15432,N_13727,N_14982);
and U15433 (N_15433,N_12368,N_10726);
and U15434 (N_15434,N_13988,N_11000);
nor U15435 (N_15435,N_11754,N_10407);
nand U15436 (N_15436,N_13930,N_10160);
or U15437 (N_15437,N_11974,N_12742);
nor U15438 (N_15438,N_12255,N_10622);
and U15439 (N_15439,N_11820,N_10070);
nand U15440 (N_15440,N_13843,N_13310);
and U15441 (N_15441,N_12673,N_13862);
and U15442 (N_15442,N_14083,N_12200);
nand U15443 (N_15443,N_14101,N_12543);
and U15444 (N_15444,N_11781,N_10496);
nor U15445 (N_15445,N_10603,N_10478);
nand U15446 (N_15446,N_12479,N_13223);
and U15447 (N_15447,N_13834,N_10401);
or U15448 (N_15448,N_11883,N_12066);
and U15449 (N_15449,N_10026,N_13128);
or U15450 (N_15450,N_13174,N_14398);
nor U15451 (N_15451,N_13284,N_12927);
or U15452 (N_15452,N_11274,N_11472);
and U15453 (N_15453,N_12982,N_14505);
nor U15454 (N_15454,N_14922,N_11517);
nor U15455 (N_15455,N_12007,N_11172);
and U15456 (N_15456,N_14987,N_12055);
nor U15457 (N_15457,N_10576,N_14509);
and U15458 (N_15458,N_14501,N_10752);
nand U15459 (N_15459,N_12423,N_12919);
and U15460 (N_15460,N_13877,N_10807);
nor U15461 (N_15461,N_14878,N_13358);
nor U15462 (N_15462,N_14909,N_12651);
nor U15463 (N_15463,N_10295,N_12932);
or U15464 (N_15464,N_10554,N_11276);
or U15465 (N_15465,N_11459,N_12334);
or U15466 (N_15466,N_12636,N_11836);
nor U15467 (N_15467,N_11801,N_12665);
and U15468 (N_15468,N_11077,N_13477);
nand U15469 (N_15469,N_12903,N_10007);
and U15470 (N_15470,N_13707,N_11269);
or U15471 (N_15471,N_13480,N_13954);
and U15472 (N_15472,N_13539,N_12490);
and U15473 (N_15473,N_11881,N_11661);
nand U15474 (N_15474,N_10060,N_10133);
or U15475 (N_15475,N_13120,N_11329);
and U15476 (N_15476,N_11120,N_11451);
nand U15477 (N_15477,N_11526,N_14676);
and U15478 (N_15478,N_14332,N_12449);
nor U15479 (N_15479,N_13808,N_12257);
or U15480 (N_15480,N_12768,N_11087);
nor U15481 (N_15481,N_11360,N_13783);
and U15482 (N_15482,N_13829,N_12142);
or U15483 (N_15483,N_11566,N_11514);
nand U15484 (N_15484,N_14761,N_10409);
nor U15485 (N_15485,N_14170,N_13536);
nand U15486 (N_15486,N_11642,N_11455);
and U15487 (N_15487,N_10767,N_13466);
nand U15488 (N_15488,N_13640,N_10423);
and U15489 (N_15489,N_14901,N_10630);
and U15490 (N_15490,N_10699,N_12780);
nor U15491 (N_15491,N_10940,N_14815);
nor U15492 (N_15492,N_10668,N_12371);
nor U15493 (N_15493,N_11407,N_14853);
nor U15494 (N_15494,N_14976,N_14716);
or U15495 (N_15495,N_12063,N_13219);
nor U15496 (N_15496,N_13149,N_12527);
nor U15497 (N_15497,N_11690,N_10594);
nor U15498 (N_15498,N_10104,N_11906);
nand U15499 (N_15499,N_12835,N_14793);
nor U15500 (N_15500,N_10274,N_10719);
nand U15501 (N_15501,N_14323,N_10570);
or U15502 (N_15502,N_14315,N_14832);
and U15503 (N_15503,N_13900,N_12182);
or U15504 (N_15504,N_12099,N_14945);
or U15505 (N_15505,N_12691,N_10063);
nor U15506 (N_15506,N_12274,N_14185);
and U15507 (N_15507,N_10708,N_10264);
nor U15508 (N_15508,N_10830,N_13785);
and U15509 (N_15509,N_13912,N_10683);
or U15510 (N_15510,N_10809,N_14977);
and U15511 (N_15511,N_13661,N_13319);
nand U15512 (N_15512,N_13428,N_12461);
and U15513 (N_15513,N_10379,N_11673);
nand U15514 (N_15514,N_11502,N_11783);
or U15515 (N_15515,N_13710,N_12191);
or U15516 (N_15516,N_12867,N_13525);
nand U15517 (N_15517,N_12644,N_11527);
or U15518 (N_15518,N_12506,N_11707);
nor U15519 (N_15519,N_12240,N_10565);
xnor U15520 (N_15520,N_11228,N_10818);
and U15521 (N_15521,N_13457,N_10880);
nor U15522 (N_15522,N_10943,N_10741);
and U15523 (N_15523,N_13907,N_11397);
nand U15524 (N_15524,N_11511,N_10459);
nand U15525 (N_15525,N_11143,N_12106);
or U15526 (N_15526,N_14317,N_10325);
nor U15527 (N_15527,N_11321,N_13221);
nand U15528 (N_15528,N_12661,N_14037);
or U15529 (N_15529,N_14461,N_11355);
nor U15530 (N_15530,N_14073,N_12214);
or U15531 (N_15531,N_12444,N_12486);
or U15532 (N_15532,N_13566,N_14246);
nor U15533 (N_15533,N_10333,N_12613);
nor U15534 (N_15534,N_10463,N_10213);
nor U15535 (N_15535,N_12941,N_14696);
nor U15536 (N_15536,N_13809,N_13183);
and U15537 (N_15537,N_13784,N_10749);
or U15538 (N_15538,N_13782,N_14668);
or U15539 (N_15539,N_12723,N_12552);
nand U15540 (N_15540,N_10041,N_12408);
and U15541 (N_15541,N_14644,N_12147);
nand U15542 (N_15542,N_13594,N_14582);
nand U15543 (N_15543,N_14641,N_11155);
nor U15544 (N_15544,N_14607,N_11763);
nor U15545 (N_15545,N_14275,N_11188);
nand U15546 (N_15546,N_12588,N_12765);
and U15547 (N_15547,N_11061,N_12530);
nor U15548 (N_15548,N_14973,N_12784);
nor U15549 (N_15549,N_14985,N_14674);
or U15550 (N_15550,N_12440,N_11727);
or U15551 (N_15551,N_13407,N_14726);
and U15552 (N_15552,N_12581,N_12525);
nor U15553 (N_15553,N_10196,N_12161);
or U15554 (N_15554,N_12802,N_13879);
or U15555 (N_15555,N_13156,N_13343);
xnor U15556 (N_15556,N_13943,N_10614);
and U15557 (N_15557,N_12744,N_11484);
or U15558 (N_15558,N_10485,N_13673);
and U15559 (N_15559,N_12568,N_11279);
nand U15560 (N_15560,N_10950,N_12615);
or U15561 (N_15561,N_10857,N_10909);
and U15562 (N_15562,N_10106,N_11516);
nand U15563 (N_15563,N_11887,N_13416);
nor U15564 (N_15564,N_14740,N_14609);
and U15565 (N_15565,N_14938,N_10307);
nor U15566 (N_15566,N_14009,N_11768);
nor U15567 (N_15567,N_14951,N_12823);
or U15568 (N_15568,N_10968,N_11722);
and U15569 (N_15569,N_12858,N_11879);
nand U15570 (N_15570,N_11948,N_11975);
or U15571 (N_15571,N_14302,N_10174);
and U15572 (N_15572,N_11410,N_13230);
nand U15573 (N_15573,N_13856,N_14485);
and U15574 (N_15574,N_12961,N_14137);
xnor U15575 (N_15575,N_11721,N_10335);
nand U15576 (N_15576,N_14773,N_14337);
nor U15577 (N_15577,N_12296,N_12030);
nor U15578 (N_15578,N_13544,N_11858);
nor U15579 (N_15579,N_12841,N_11510);
nor U15580 (N_15580,N_10995,N_10220);
nand U15581 (N_15581,N_13260,N_13906);
or U15582 (N_15582,N_13492,N_13233);
nand U15583 (N_15583,N_12010,N_10883);
and U15584 (N_15584,N_12912,N_14921);
nor U15585 (N_15585,N_10209,N_11565);
or U15586 (N_15586,N_11889,N_12448);
xnor U15587 (N_15587,N_11977,N_10194);
and U15588 (N_15588,N_13889,N_12962);
xnor U15589 (N_15589,N_10938,N_13129);
nor U15590 (N_15590,N_10813,N_14139);
and U15591 (N_15591,N_14577,N_10211);
nor U15592 (N_15592,N_13424,N_10243);
nand U15593 (N_15593,N_14650,N_10036);
nor U15594 (N_15594,N_11709,N_12176);
nor U15595 (N_15595,N_11035,N_12879);
nand U15596 (N_15596,N_13917,N_13476);
xor U15597 (N_15597,N_11465,N_13973);
or U15598 (N_15598,N_13770,N_12223);
or U15599 (N_15599,N_14638,N_14454);
nor U15600 (N_15600,N_11454,N_12041);
nand U15601 (N_15601,N_10231,N_14752);
or U15602 (N_15602,N_11913,N_12114);
and U15603 (N_15603,N_11039,N_13228);
nand U15604 (N_15604,N_13249,N_12692);
or U15605 (N_15605,N_12827,N_12602);
nor U15606 (N_15606,N_11934,N_11873);
nand U15607 (N_15607,N_14316,N_12657);
nand U15608 (N_15608,N_12626,N_12264);
and U15609 (N_15609,N_10419,N_12265);
or U15610 (N_15610,N_13048,N_12079);
nand U15611 (N_15611,N_12639,N_10024);
or U15612 (N_15612,N_10684,N_11473);
nand U15613 (N_15613,N_13551,N_14478);
and U15614 (N_15614,N_11651,N_10092);
nand U15615 (N_15615,N_14082,N_13870);
and U15616 (N_15616,N_12367,N_12175);
or U15617 (N_15617,N_14682,N_12342);
nor U15618 (N_15618,N_13132,N_10686);
xor U15619 (N_15619,N_14114,N_12382);
nand U15620 (N_15620,N_13660,N_14292);
nor U15621 (N_15621,N_11375,N_10290);
nand U15622 (N_15622,N_10203,N_14500);
or U15623 (N_15623,N_13538,N_13699);
nor U15624 (N_15624,N_14044,N_13920);
or U15625 (N_15625,N_13649,N_10121);
and U15626 (N_15626,N_13196,N_11409);
nor U15627 (N_15627,N_10487,N_12134);
nand U15628 (N_15628,N_10439,N_13929);
nor U15629 (N_15629,N_14713,N_10279);
nor U15630 (N_15630,N_10462,N_12566);
or U15631 (N_15631,N_10704,N_11767);
nor U15632 (N_15632,N_13397,N_11532);
and U15633 (N_15633,N_13506,N_13276);
nor U15634 (N_15634,N_10030,N_13377);
or U15635 (N_15635,N_10173,N_14855);
nand U15636 (N_15636,N_10132,N_13166);
nand U15637 (N_15637,N_13497,N_11838);
nand U15638 (N_15638,N_13915,N_14799);
or U15639 (N_15639,N_14811,N_12810);
or U15640 (N_15640,N_13087,N_11271);
or U15641 (N_15641,N_10215,N_14758);
nand U15642 (N_15642,N_12004,N_14545);
nand U15643 (N_15643,N_14914,N_11597);
or U15644 (N_15644,N_12393,N_14942);
nand U15645 (N_15645,N_13148,N_12293);
nor U15646 (N_15646,N_14762,N_13059);
nor U15647 (N_15647,N_11990,N_13987);
nor U15648 (N_15648,N_13298,N_11088);
and U15649 (N_15649,N_12332,N_12497);
or U15650 (N_15650,N_14721,N_10885);
nor U15651 (N_15651,N_10037,N_10982);
nand U15652 (N_15652,N_10651,N_14646);
or U15653 (N_15653,N_11657,N_14665);
and U15654 (N_15654,N_11544,N_14510);
nand U15655 (N_15655,N_11788,N_11072);
and U15656 (N_15656,N_11826,N_10345);
xor U15657 (N_15657,N_13864,N_11026);
nand U15658 (N_15658,N_13184,N_10948);
and U15659 (N_15659,N_11348,N_11122);
or U15660 (N_15660,N_10071,N_12341);
nor U15661 (N_15661,N_10310,N_13731);
or U15662 (N_15662,N_12577,N_10954);
or U15663 (N_15663,N_10093,N_12571);
and U15664 (N_15664,N_10629,N_13222);
nand U15665 (N_15665,N_11916,N_12991);
nor U15666 (N_15666,N_14707,N_14984);
and U15667 (N_15667,N_11822,N_12739);
nor U15668 (N_15668,N_12400,N_12659);
nor U15669 (N_15669,N_11330,N_13979);
and U15670 (N_15670,N_14370,N_12966);
and U15671 (N_15671,N_13367,N_10797);
nor U15672 (N_15672,N_11280,N_12960);
or U15673 (N_15673,N_14015,N_10583);
nand U15674 (N_15674,N_13317,N_13730);
nand U15675 (N_15675,N_14029,N_11605);
nand U15676 (N_15676,N_13373,N_14614);
nand U15677 (N_15677,N_10327,N_13561);
or U15678 (N_15678,N_14351,N_13033);
or U15679 (N_15679,N_14539,N_12792);
and U15680 (N_15680,N_13807,N_14464);
and U15681 (N_15681,N_14603,N_11301);
nand U15682 (N_15682,N_10431,N_13902);
and U15683 (N_15683,N_12796,N_14491);
and U15684 (N_15684,N_14684,N_10354);
nand U15685 (N_15685,N_12167,N_11751);
and U15686 (N_15686,N_10210,N_11461);
nor U15687 (N_15687,N_12668,N_13823);
or U15688 (N_15688,N_13177,N_10349);
and U15689 (N_15689,N_11851,N_10214);
nor U15690 (N_15690,N_13364,N_11247);
nand U15691 (N_15691,N_10200,N_13309);
nand U15692 (N_15692,N_12646,N_11666);
nand U15693 (N_15693,N_10162,N_13383);
or U15694 (N_15694,N_10914,N_14588);
nand U15695 (N_15695,N_14792,N_11922);
xnor U15696 (N_15696,N_12696,N_10006);
and U15697 (N_15697,N_10616,N_12537);
and U15698 (N_15698,N_11316,N_10731);
and U15699 (N_15699,N_10052,N_12600);
nand U15700 (N_15700,N_14311,N_14357);
and U15701 (N_15701,N_13880,N_13657);
and U15702 (N_15702,N_13565,N_14648);
nand U15703 (N_15703,N_10510,N_14586);
nand U15704 (N_15704,N_13899,N_10662);
nand U15705 (N_15705,N_14936,N_14858);
and U15706 (N_15706,N_11008,N_12230);
or U15707 (N_15707,N_13022,N_13108);
nand U15708 (N_15708,N_12166,N_10514);
nor U15709 (N_15709,N_12855,N_13887);
or U15710 (N_15710,N_10314,N_12755);
nor U15711 (N_15711,N_10947,N_10854);
xnor U15712 (N_15712,N_14460,N_11986);
nand U15713 (N_15713,N_11377,N_14473);
and U15714 (N_15714,N_12298,N_12011);
xnor U15715 (N_15715,N_10156,N_14946);
or U15716 (N_15716,N_13847,N_13044);
xnor U15717 (N_15717,N_13333,N_12287);
and U15718 (N_15718,N_11629,N_11830);
nor U15719 (N_15719,N_13855,N_14457);
and U15720 (N_15720,N_10802,N_10126);
and U15721 (N_15721,N_10352,N_10185);
xnor U15722 (N_15722,N_13171,N_12986);
nand U15723 (N_15723,N_11069,N_13306);
nand U15724 (N_15724,N_14273,N_11757);
and U15725 (N_15725,N_13187,N_14265);
and U15726 (N_15726,N_13564,N_10096);
nor U15727 (N_15727,N_12747,N_14283);
or U15728 (N_15728,N_10397,N_10787);
nor U15729 (N_15729,N_10361,N_11242);
nor U15730 (N_15730,N_14808,N_14596);
and U15731 (N_15731,N_10167,N_11201);
nand U15732 (N_15732,N_11085,N_12062);
and U15733 (N_15733,N_11591,N_12623);
and U15734 (N_15734,N_14948,N_14287);
nor U15735 (N_15735,N_10777,N_12465);
nor U15736 (N_15736,N_12578,N_10625);
and U15737 (N_15737,N_10280,N_14088);
or U15738 (N_15738,N_10886,N_13342);
or U15739 (N_15739,N_13078,N_13720);
or U15740 (N_15740,N_14941,N_10698);
nor U15741 (N_15741,N_10641,N_10059);
nor U15742 (N_15742,N_10291,N_12522);
or U15743 (N_15743,N_13100,N_11356);
xor U15744 (N_15744,N_12278,N_12178);
nor U15745 (N_15745,N_13653,N_11756);
nand U15746 (N_15746,N_12216,N_13910);
nand U15747 (N_15747,N_13685,N_13747);
and U15748 (N_15748,N_14953,N_13293);
xnor U15749 (N_15749,N_10523,N_13213);
nor U15750 (N_15750,N_11038,N_11880);
nand U15751 (N_15751,N_11100,N_13804);
nor U15752 (N_15752,N_12520,N_11435);
nand U15753 (N_15753,N_14397,N_13395);
nor U15754 (N_15754,N_13739,N_10311);
xor U15755 (N_15755,N_14474,N_11001);
and U15756 (N_15756,N_12049,N_11431);
nor U15757 (N_15757,N_10004,N_14809);
xor U15758 (N_15758,N_13039,N_14441);
nor U15759 (N_15759,N_12849,N_10581);
or U15760 (N_15760,N_12463,N_12515);
or U15761 (N_15761,N_11197,N_13779);
nor U15762 (N_15762,N_14845,N_14962);
or U15763 (N_15763,N_10911,N_13953);
and U15764 (N_15764,N_11601,N_11134);
and U15765 (N_15765,N_14699,N_12288);
or U15766 (N_15766,N_14971,N_12061);
or U15767 (N_15767,N_10222,N_10657);
or U15768 (N_15768,N_12192,N_14263);
nor U15769 (N_15769,N_13993,N_13647);
nand U15770 (N_15770,N_11254,N_14595);
nand U15771 (N_15771,N_12844,N_13813);
or U15772 (N_15772,N_13737,N_14378);
nor U15773 (N_15773,N_14954,N_13266);
or U15774 (N_15774,N_13514,N_10105);
and U15775 (N_15775,N_14757,N_13736);
nand U15776 (N_15776,N_14636,N_10642);
and U15777 (N_15777,N_12413,N_14338);
and U15778 (N_15778,N_14959,N_11521);
and U15779 (N_15779,N_10402,N_12271);
nor U15780 (N_15780,N_11175,N_13959);
or U15781 (N_15781,N_10002,N_12380);
or U15782 (N_15782,N_11670,N_11023);
and U15783 (N_15783,N_10706,N_11753);
or U15784 (N_15784,N_11307,N_11846);
or U15785 (N_15785,N_11229,N_11957);
and U15786 (N_15786,N_10165,N_14046);
nor U15787 (N_15787,N_13949,N_13280);
nor U15788 (N_15788,N_10747,N_10481);
nand U15789 (N_15789,N_13024,N_10853);
or U15790 (N_15790,N_12698,N_13299);
nor U15791 (N_15791,N_11466,N_11032);
nand U15792 (N_15792,N_13467,N_13975);
nand U15793 (N_15793,N_11505,N_12173);
or U15794 (N_15794,N_12507,N_13257);
nor U15795 (N_15795,N_10770,N_11547);
or U15796 (N_15796,N_11283,N_14304);
nand U15797 (N_15797,N_14194,N_10793);
and U15798 (N_15798,N_11150,N_10931);
and U15799 (N_15799,N_11985,N_12357);
or U15800 (N_15800,N_14459,N_14215);
and U15801 (N_15801,N_13655,N_10050);
or U15802 (N_15802,N_10471,N_14356);
and U15803 (N_15803,N_12779,N_10966);
nand U15804 (N_15804,N_12153,N_10645);
or U15805 (N_15805,N_11354,N_10820);
xor U15806 (N_15806,N_12786,N_11380);
xnor U15807 (N_15807,N_12437,N_13746);
and U15808 (N_15808,N_11612,N_13537);
nor U15809 (N_15809,N_14479,N_12597);
nor U15810 (N_15810,N_10328,N_11792);
and U15811 (N_15811,N_11815,N_13386);
or U15812 (N_15812,N_13684,N_13874);
and U15813 (N_15813,N_14580,N_13458);
or U15814 (N_15814,N_14051,N_14810);
nand U15815 (N_15815,N_14028,N_11619);
nor U15816 (N_15816,N_13186,N_11302);
and U15817 (N_15817,N_14957,N_12731);
nor U15818 (N_15818,N_11002,N_14175);
nand U15819 (N_15819,N_12889,N_13288);
nor U15820 (N_15820,N_13714,N_13562);
and U15821 (N_15821,N_12977,N_10650);
and U15822 (N_15822,N_12125,N_14786);
nand U15823 (N_15823,N_14140,N_13742);
nor U15824 (N_15824,N_12526,N_14373);
nor U15825 (N_15825,N_13029,N_13179);
nor U15826 (N_15826,N_13938,N_12370);
nor U15827 (N_15827,N_14002,N_14003);
nand U15828 (N_15828,N_13144,N_10494);
nand U15829 (N_15829,N_12491,N_12724);
nor U15830 (N_15830,N_11776,N_12052);
and U15831 (N_15831,N_10649,N_11654);
and U15832 (N_15832,N_11270,N_11037);
or U15833 (N_15833,N_14306,N_11575);
and U15834 (N_15834,N_13854,N_13061);
or U15835 (N_15835,N_14095,N_11181);
and U15836 (N_15836,N_13195,N_10561);
or U15837 (N_15837,N_10596,N_11129);
or U15838 (N_15838,N_12864,N_14155);
and U15839 (N_15839,N_11655,N_11123);
or U15840 (N_15840,N_10796,N_11872);
and U15841 (N_15841,N_11198,N_12082);
or U15842 (N_15842,N_13921,N_11839);
and U15843 (N_15843,N_11111,N_12632);
or U15844 (N_15844,N_14498,N_13700);
and U15845 (N_15845,N_12450,N_13494);
nand U15846 (N_15846,N_14899,N_12251);
nor U15847 (N_15847,N_14250,N_12767);
nand U15848 (N_15848,N_12655,N_12975);
and U15849 (N_15849,N_11845,N_14730);
xnor U15850 (N_15850,N_13471,N_14016);
and U15851 (N_15851,N_12707,N_14226);
nand U15852 (N_15852,N_13521,N_10045);
nor U15853 (N_15853,N_11130,N_14147);
nand U15854 (N_15854,N_11823,N_10737);
and U15855 (N_15855,N_12567,N_14533);
xnor U15856 (N_15856,N_13142,N_13331);
nor U15857 (N_15857,N_11045,N_14570);
or U15858 (N_15858,N_14849,N_12700);
nand U15859 (N_15859,N_13549,N_13595);
nand U15860 (N_15860,N_10309,N_11503);
nand U15861 (N_15861,N_13517,N_14390);
nand U15862 (N_15862,N_13117,N_14026);
and U15863 (N_15863,N_12607,N_14983);
nor U15864 (N_15864,N_10976,N_14324);
and U15865 (N_15865,N_10181,N_14834);
nand U15866 (N_15866,N_10170,N_11012);
nand U15867 (N_15867,N_12411,N_13332);
and U15868 (N_15868,N_10501,N_12918);
or U15869 (N_15869,N_11324,N_13677);
nor U15870 (N_15870,N_10863,N_14550);
or U15871 (N_15871,N_14874,N_11650);
or U15872 (N_15872,N_14744,N_11158);
nor U15873 (N_15873,N_14445,N_12050);
or U15874 (N_15874,N_12190,N_14666);
nand U15875 (N_15875,N_13605,N_10022);
and U15876 (N_15876,N_12430,N_13303);
and U15877 (N_15877,N_14318,N_12140);
nand U15878 (N_15878,N_13945,N_12421);
nand U15879 (N_15879,N_11156,N_13005);
nand U15880 (N_15880,N_13608,N_11531);
nand U15881 (N_15881,N_12356,N_14235);
nand U15882 (N_15882,N_11631,N_14523);
nand U15883 (N_15883,N_12398,N_13821);
and U15884 (N_15884,N_14158,N_10069);
and U15885 (N_15885,N_11108,N_10404);
nor U15886 (N_15886,N_11915,N_12704);
and U15887 (N_15887,N_10723,N_11585);
nand U15888 (N_15888,N_10984,N_13583);
or U15889 (N_15889,N_12538,N_11477);
nand U15890 (N_15890,N_11350,N_13083);
and U15891 (N_15891,N_14712,N_14837);
nand U15892 (N_15892,N_12979,N_12489);
nor U15893 (N_15893,N_10748,N_12981);
nand U15894 (N_15894,N_13315,N_11325);
and U15895 (N_15895,N_13151,N_12388);
nor U15896 (N_15896,N_14297,N_12163);
and U15897 (N_15897,N_12728,N_13130);
or U15898 (N_15898,N_11019,N_14568);
nand U15899 (N_15899,N_10111,N_14054);
nand U15900 (N_15900,N_13401,N_12294);
nand U15901 (N_15901,N_11683,N_10680);
nand U15902 (N_15902,N_13226,N_12111);
or U15903 (N_15903,N_14559,N_12137);
and U15904 (N_15904,N_14939,N_14967);
nor U15905 (N_15905,N_14488,N_12446);
nand U15906 (N_15906,N_13216,N_12938);
nor U15907 (N_15907,N_10469,N_14868);
and U15908 (N_15908,N_11347,N_13425);
and U15909 (N_15909,N_11681,N_14880);
or U15910 (N_15910,N_10671,N_10677);
nor U15911 (N_15911,N_11396,N_13045);
or U15912 (N_15912,N_13827,N_13750);
and U15913 (N_15913,N_12350,N_13427);
or U15914 (N_15914,N_12343,N_13390);
nand U15915 (N_15915,N_14165,N_11028);
nand U15916 (N_15916,N_10915,N_12616);
and U15917 (N_15917,N_13327,N_14723);
nor U15918 (N_15918,N_13300,N_13482);
nor U15919 (N_15919,N_11171,N_13556);
or U15920 (N_15920,N_13623,N_13690);
nand U15921 (N_15921,N_10841,N_12434);
or U15922 (N_15922,N_14866,N_12130);
nand U15923 (N_15923,N_11411,N_11557);
xnor U15924 (N_15924,N_11641,N_12160);
or U15925 (N_15925,N_13314,N_14270);
or U15926 (N_15926,N_13972,N_12913);
and U15927 (N_15927,N_13322,N_11385);
nor U15928 (N_15928,N_12611,N_12346);
nand U15929 (N_15929,N_12247,N_10562);
and U15930 (N_15930,N_10913,N_13270);
and U15931 (N_15931,N_14182,N_11996);
nor U15932 (N_15932,N_13567,N_13628);
or U15933 (N_15933,N_10964,N_12196);
or U15934 (N_15934,N_13014,N_10003);
nand U15935 (N_15935,N_10848,N_11064);
and U15936 (N_15936,N_10972,N_14289);
xor U15937 (N_15937,N_10391,N_13865);
or U15938 (N_15938,N_11394,N_11762);
nand U15939 (N_15939,N_13426,N_14385);
nand U15940 (N_15940,N_11440,N_13456);
and U15941 (N_15941,N_13502,N_11339);
xnor U15942 (N_15942,N_14795,N_11369);
and U15943 (N_15943,N_14399,N_14819);
and U15944 (N_15944,N_14469,N_10051);
nand U15945 (N_15945,N_10769,N_14143);
nor U15946 (N_15946,N_12840,N_10721);
nand U15947 (N_15947,N_10654,N_14377);
nor U15948 (N_15948,N_12729,N_10441);
or U15949 (N_15949,N_10191,N_12139);
and U15950 (N_15950,N_12301,N_12469);
and U15951 (N_15951,N_13950,N_13701);
nand U15952 (N_15952,N_14230,N_13512);
or U15953 (N_15953,N_11593,N_13868);
and U15954 (N_15954,N_10542,N_10568);
or U15955 (N_15955,N_11105,N_14380);
nand U15956 (N_15956,N_12202,N_10868);
and U15957 (N_15957,N_14529,N_13557);
nand U15958 (N_15958,N_14518,N_13066);
nor U15959 (N_15959,N_12422,N_11983);
or U15960 (N_15960,N_14902,N_13450);
or U15961 (N_15961,N_14862,N_13350);
nand U15962 (N_15962,N_14617,N_11212);
nand U15963 (N_15963,N_13410,N_10918);
or U15964 (N_15964,N_10532,N_12473);
or U15965 (N_15965,N_11614,N_14802);
nand U15966 (N_15966,N_14212,N_13713);
nand U15967 (N_15967,N_11569,N_12401);
nand U15968 (N_15968,N_12777,N_14109);
nor U15969 (N_15969,N_10492,N_12475);
or U15970 (N_15970,N_12002,N_11608);
xnor U15971 (N_15971,N_11213,N_10229);
or U15972 (N_15972,N_14645,N_12900);
or U15973 (N_15973,N_12501,N_13429);
or U15974 (N_15974,N_11142,N_14221);
xnor U15975 (N_15975,N_10718,N_10553);
and U15976 (N_15976,N_11273,N_12256);
or U15977 (N_15977,N_13703,N_10120);
or U15978 (N_15978,N_12534,N_11961);
and U15979 (N_15979,N_14978,N_14734);
or U15980 (N_15980,N_13493,N_12573);
nor U15981 (N_15981,N_13520,N_12998);
nor U15982 (N_15982,N_10235,N_11726);
and U15983 (N_15983,N_12500,N_13070);
and U15984 (N_15984,N_11686,N_14499);
nor U15985 (N_15985,N_11684,N_14371);
or U15986 (N_15986,N_13609,N_14900);
or U15987 (N_15987,N_14172,N_13370);
nor U15988 (N_15988,N_11480,N_13399);
and U15989 (N_15989,N_14269,N_13610);
and U15990 (N_15990,N_12194,N_14432);
and U15991 (N_15991,N_12797,N_13250);
nor U15992 (N_15992,N_13098,N_13459);
and U15993 (N_15993,N_13584,N_14869);
nor U15994 (N_15994,N_10910,N_10587);
and U15995 (N_15995,N_14949,N_14569);
and U15996 (N_15996,N_12016,N_13627);
nor U15997 (N_15997,N_12183,N_10665);
and U15998 (N_15998,N_14387,N_14574);
xnor U15999 (N_15999,N_13388,N_12593);
xnor U16000 (N_16000,N_10772,N_13728);
nand U16001 (N_16001,N_10690,N_11592);
nor U16002 (N_16002,N_10638,N_14363);
and U16003 (N_16003,N_14966,N_14919);
and U16004 (N_16004,N_14771,N_10298);
nor U16005 (N_16005,N_11596,N_11263);
or U16006 (N_16006,N_12798,N_13353);
or U16007 (N_16007,N_13469,N_13574);
xor U16008 (N_16008,N_11813,N_13898);
nor U16009 (N_16009,N_11926,N_11004);
nor U16010 (N_16010,N_14530,N_14346);
nor U16011 (N_16011,N_12009,N_10292);
nand U16012 (N_16012,N_12663,N_13914);
or U16013 (N_16013,N_13812,N_13247);
and U16014 (N_16014,N_14411,N_13625);
nand U16015 (N_16015,N_11648,N_11589);
nor U16016 (N_16016,N_10555,N_13786);
nand U16017 (N_16017,N_13028,N_11840);
and U16018 (N_16018,N_10493,N_14076);
or U16019 (N_16019,N_14256,N_13816);
nor U16020 (N_16020,N_11742,N_10843);
nand U16021 (N_16021,N_12410,N_14827);
nor U16022 (N_16022,N_11821,N_14754);
nor U16023 (N_16023,N_10697,N_13810);
and U16024 (N_16024,N_13091,N_13421);
nand U16025 (N_16025,N_12906,N_13391);
nor U16026 (N_16026,N_13056,N_11067);
nand U16027 (N_16027,N_12259,N_13305);
nor U16028 (N_16028,N_10484,N_12513);
nand U16029 (N_16029,N_12244,N_12151);
and U16030 (N_16030,N_12131,N_12972);
and U16031 (N_16031,N_14663,N_13872);
and U16032 (N_16032,N_11649,N_12854);
nor U16033 (N_16033,N_12123,N_12645);
and U16034 (N_16034,N_11225,N_11127);
nand U16035 (N_16035,N_12922,N_11970);
or U16036 (N_16036,N_12128,N_10860);
and U16037 (N_16037,N_11809,N_11272);
nand U16038 (N_16038,N_14248,N_12705);
nand U16039 (N_16039,N_13841,N_13019);
and U16040 (N_16040,N_10661,N_11806);
or U16041 (N_16041,N_13942,N_13239);
and U16042 (N_16042,N_14093,N_11588);
nand U16043 (N_16043,N_12329,N_10065);
or U16044 (N_16044,N_11932,N_14367);
nand U16045 (N_16045,N_13844,N_13741);
or U16046 (N_16046,N_10097,N_14379);
nor U16047 (N_16047,N_11980,N_11093);
and U16048 (N_16048,N_13057,N_11364);
nand U16049 (N_16049,N_14452,N_11189);
nor U16050 (N_16050,N_14189,N_10811);
or U16051 (N_16051,N_12711,N_10881);
nor U16052 (N_16052,N_10664,N_10526);
nor U16053 (N_16053,N_14751,N_10343);
or U16054 (N_16054,N_14112,N_13974);
nand U16055 (N_16055,N_14555,N_12680);
xnor U16056 (N_16056,N_11869,N_14687);
nand U16057 (N_16057,N_13965,N_11264);
nand U16058 (N_16058,N_11089,N_14572);
and U16059 (N_16059,N_13733,N_13324);
nor U16060 (N_16060,N_14766,N_12819);
or U16061 (N_16061,N_14228,N_12848);
nand U16062 (N_16062,N_14203,N_12481);
nor U16063 (N_16063,N_11892,N_11116);
or U16064 (N_16064,N_12378,N_11290);
nand U16065 (N_16065,N_14211,N_14525);
nand U16066 (N_16066,N_12562,N_13274);
nor U16067 (N_16067,N_14947,N_14594);
or U16068 (N_16068,N_10666,N_13192);
nand U16069 (N_16069,N_10221,N_14626);
nand U16070 (N_16070,N_11560,N_14520);
and U16071 (N_16071,N_10759,N_10430);
and U16072 (N_16072,N_10341,N_14640);
and U16073 (N_16073,N_10873,N_10864);
nand U16074 (N_16074,N_12582,N_14655);
xnor U16075 (N_16075,N_13271,N_10115);
or U16076 (N_16076,N_14675,N_12038);
and U16077 (N_16077,N_13519,N_12791);
or U16078 (N_16078,N_11795,N_12210);
or U16079 (N_16079,N_12392,N_13820);
and U16080 (N_16080,N_13662,N_13861);
nor U16081 (N_16081,N_11236,N_13916);
and U16082 (N_16082,N_10438,N_12037);
and U16083 (N_16083,N_12462,N_11576);
nor U16084 (N_16084,N_11555,N_10305);
nand U16085 (N_16085,N_14343,N_10299);
nand U16086 (N_16086,N_13886,N_10503);
and U16087 (N_16087,N_13202,N_11925);
or U16088 (N_16088,N_14201,N_13788);
nand U16089 (N_16089,N_11210,N_10001);
nor U16090 (N_16090,N_10029,N_12838);
nor U16091 (N_16091,N_11833,N_12069);
nand U16092 (N_16092,N_14437,N_11389);
nand U16093 (N_16093,N_11877,N_13123);
nor U16094 (N_16094,N_13485,N_13931);
and U16095 (N_16095,N_13402,N_14642);
nand U16096 (N_16096,N_11058,N_12220);
or U16097 (N_16097,N_13326,N_10444);
nand U16098 (N_16098,N_12888,N_12517);
nand U16099 (N_16099,N_10504,N_12836);
nor U16100 (N_16100,N_10258,N_10618);
nand U16101 (N_16101,N_13578,N_14673);
nand U16102 (N_16102,N_10612,N_10991);
nand U16103 (N_16103,N_10786,N_14658);
nand U16104 (N_16104,N_11154,N_10710);
nand U16105 (N_16105,N_12143,N_11382);
or U16106 (N_16106,N_12592,N_12234);
and U16107 (N_16107,N_11227,N_12752);
xor U16108 (N_16108,N_13702,N_11421);
nor U16109 (N_16109,N_11797,N_14911);
nor U16110 (N_16110,N_12231,N_12806);
nand U16111 (N_16111,N_14920,N_13290);
and U16112 (N_16112,N_10892,N_10324);
or U16113 (N_16113,N_12818,N_10016);
and U16114 (N_16114,N_11253,N_12246);
and U16115 (N_16115,N_11705,N_12685);
and U16116 (N_16116,N_10053,N_14031);
or U16117 (N_16117,N_10608,N_10903);
xnor U16118 (N_16118,N_13819,N_14180);
nand U16119 (N_16119,N_12085,N_11736);
nor U16120 (N_16120,N_12897,N_11735);
nand U16121 (N_16121,N_12086,N_12893);
and U16122 (N_16122,N_14895,N_13328);
nor U16123 (N_16123,N_13191,N_11580);
or U16124 (N_16124,N_12145,N_13764);
nand U16125 (N_16125,N_13320,N_11468);
nor U16126 (N_16126,N_13601,N_12625);
nor U16127 (N_16127,N_10908,N_11470);
or U16128 (N_16128,N_11126,N_11761);
or U16129 (N_16129,N_14011,N_13037);
nor U16130 (N_16130,N_11739,N_12734);
and U16131 (N_16131,N_12068,N_14532);
nor U16132 (N_16132,N_10852,N_12262);
and U16133 (N_16133,N_11131,N_12096);
nor U16134 (N_16134,N_12832,N_12495);
nor U16135 (N_16135,N_10833,N_11832);
nand U16136 (N_16136,N_12524,N_13952);
and U16137 (N_16137,N_13814,N_14145);
nand U16138 (N_16138,N_10524,N_11094);
nor U16139 (N_16139,N_10370,N_13345);
nand U16140 (N_16140,N_13038,N_11239);
nand U16141 (N_16141,N_12105,N_12115);
nor U16142 (N_16142,N_14299,N_11365);
or U16143 (N_16143,N_11119,N_12783);
and U16144 (N_16144,N_14188,N_10420);
nand U16145 (N_16145,N_10129,N_13944);
nand U16146 (N_16146,N_14423,N_14234);
nand U16147 (N_16147,N_10846,N_12222);
and U16148 (N_16148,N_11988,N_14516);
nand U16149 (N_16149,N_12053,N_12572);
or U16150 (N_16150,N_10862,N_14824);
nand U16151 (N_16151,N_10812,N_12951);
or U16152 (N_16152,N_10728,N_10284);
or U16153 (N_16153,N_13971,N_12866);
and U16154 (N_16154,N_11628,N_14605);
or U16155 (N_16155,N_13792,N_13946);
nand U16156 (N_16156,N_13141,N_13393);
and U16157 (N_16157,N_10736,N_11476);
and U16158 (N_16158,N_14528,N_12129);
or U16159 (N_16159,N_14564,N_14893);
or U16160 (N_16160,N_10376,N_11303);
nor U16161 (N_16161,N_13937,N_14438);
nand U16162 (N_16162,N_14425,N_10507);
and U16163 (N_16163,N_12340,N_12328);
nor U16164 (N_16164,N_12335,N_12845);
xor U16165 (N_16165,N_14100,N_12874);
and U16166 (N_16166,N_13683,N_14526);
nor U16167 (N_16167,N_13706,N_13546);
and U16168 (N_16168,N_12025,N_10386);
or U16169 (N_16169,N_13708,N_11899);
and U16170 (N_16170,N_12292,N_12097);
and U16171 (N_16171,N_14217,N_10323);
nor U16172 (N_16172,N_14127,N_13569);
nand U16173 (N_16173,N_12327,N_12032);
nand U16174 (N_16174,N_14160,N_11102);
nor U16175 (N_16175,N_12622,N_11924);
nor U16176 (N_16176,N_12800,N_14240);
or U16177 (N_16177,N_11647,N_10033);
nand U16178 (N_16178,N_10348,N_11595);
and U16179 (N_16179,N_10357,N_13385);
nor U16180 (N_16180,N_10250,N_11159);
and U16181 (N_16181,N_10390,N_11215);
xnor U16182 (N_16182,N_12703,N_14374);
nand U16183 (N_16183,N_13099,N_10962);
or U16184 (N_16184,N_11178,N_13599);
xnor U16185 (N_16185,N_10571,N_10467);
nor U16186 (N_16186,N_10682,N_12221);
nand U16187 (N_16187,N_13760,N_14992);
and U16188 (N_16188,N_11163,N_11513);
nand U16189 (N_16189,N_13297,N_12237);
nor U16190 (N_16190,N_14892,N_11495);
and U16191 (N_16191,N_14694,N_11955);
and U16192 (N_16192,N_12118,N_10547);
and U16193 (N_16193,N_14197,N_11507);
or U16194 (N_16194,N_14022,N_11278);
nand U16195 (N_16195,N_10316,N_11371);
and U16196 (N_16196,N_13650,N_14014);
nand U16197 (N_16197,N_14200,N_12708);
nand U16198 (N_16198,N_12492,N_11133);
nand U16199 (N_16199,N_14336,N_14077);
xor U16200 (N_16200,N_11458,N_12459);
nor U16201 (N_16201,N_13992,N_14405);
nor U16202 (N_16202,N_10595,N_13771);
and U16203 (N_16203,N_10089,N_12144);
nand U16204 (N_16204,N_14120,N_11750);
or U16205 (N_16205,N_14266,N_14784);
or U16206 (N_16206,N_10893,N_10363);
nor U16207 (N_16207,N_14227,N_11298);
or U16208 (N_16208,N_10177,N_10338);
nor U16209 (N_16209,N_14635,N_12787);
or U16210 (N_16210,N_13600,N_11482);
or U16211 (N_16211,N_11488,N_10997);
and U16212 (N_16212,N_13050,N_11870);
and U16213 (N_16213,N_13170,N_14546);
and U16214 (N_16214,N_12232,N_10768);
and U16215 (N_16215,N_11910,N_14236);
nor U16216 (N_16216,N_14791,N_11850);
or U16217 (N_16217,N_13759,N_13238);
nand U16218 (N_16218,N_10255,N_10044);
and U16219 (N_16219,N_12677,N_11734);
and U16220 (N_16220,N_13797,N_11169);
nor U16221 (N_16221,N_13051,N_11351);
and U16222 (N_16222,N_12587,N_13818);
or U16223 (N_16223,N_14727,N_10199);
nand U16224 (N_16224,N_14693,N_11297);
and U16225 (N_16225,N_11743,N_14481);
nand U16226 (N_16226,N_12036,N_13777);
nand U16227 (N_16227,N_12474,N_13463);
nor U16228 (N_16228,N_14794,N_12233);
and U16229 (N_16229,N_14249,N_11427);
or U16230 (N_16230,N_13435,N_12604);
nand U16231 (N_16231,N_12245,N_14549);
or U16232 (N_16232,N_10888,N_12360);
nor U16233 (N_16233,N_11938,N_11804);
or U16234 (N_16234,N_13308,N_12926);
and U16235 (N_16235,N_14571,N_10776);
nand U16236 (N_16236,N_10924,N_13277);
and U16237 (N_16237,N_10054,N_13484);
and U16238 (N_16238,N_11528,N_12325);
and U16239 (N_16239,N_11240,N_14865);
and U16240 (N_16240,N_14710,N_10495);
and U16241 (N_16241,N_11905,N_12480);
nor U16242 (N_16242,N_11626,N_14524);
nand U16243 (N_16243,N_14747,N_11144);
and U16244 (N_16244,N_14308,N_12598);
nor U16245 (N_16245,N_12512,N_14830);
and U16246 (N_16246,N_11314,N_12885);
nor U16247 (N_16247,N_13763,N_14497);
or U16248 (N_16248,N_14484,N_13444);
or U16249 (N_16249,N_12386,N_10815);
or U16250 (N_16250,N_14456,N_14099);
or U16251 (N_16251,N_13977,N_10278);
nor U16252 (N_16252,N_13723,N_13178);
nand U16253 (N_16253,N_11894,N_11630);
nor U16254 (N_16254,N_13075,N_10865);
and U16255 (N_16255,N_14660,N_13201);
nor U16256 (N_16256,N_11506,N_13542);
and U16257 (N_16257,N_12060,N_14722);
nand U16258 (N_16258,N_11896,N_13596);
nor U16259 (N_16259,N_10956,N_10145);
or U16260 (N_16260,N_12809,N_10447);
and U16261 (N_16261,N_11051,N_13922);
or U16262 (N_16262,N_10602,N_13400);
or U16263 (N_16263,N_12353,N_14418);
nor U16264 (N_16264,N_14542,N_10384);
xnor U16265 (N_16265,N_14652,N_12580);
and U16266 (N_16266,N_13652,N_10700);
nor U16267 (N_16267,N_13264,N_11733);
nor U16268 (N_16268,N_10582,N_10989);
or U16269 (N_16269,N_13243,N_12563);
or U16270 (N_16270,N_12289,N_13524);
and U16271 (N_16271,N_14392,N_11936);
and U16272 (N_16272,N_13498,N_10276);
nor U16273 (N_16273,N_11256,N_11882);
or U16274 (N_16274,N_14622,N_10891);
nand U16275 (N_16275,N_11731,N_13790);
nand U16276 (N_16276,N_14322,N_11777);
nor U16277 (N_16277,N_12788,N_10856);
and U16278 (N_16278,N_12856,N_10907);
and U16279 (N_16279,N_14281,N_11782);
nor U16280 (N_16280,N_11025,N_14179);
nand U16281 (N_16281,N_12158,N_12965);
nand U16282 (N_16282,N_11888,N_11967);
nand U16283 (N_16283,N_14661,N_12307);
and U16284 (N_16284,N_10505,N_12101);
or U16285 (N_16285,N_13211,N_11207);
or U16286 (N_16286,N_12309,N_11574);
and U16287 (N_16287,N_14125,N_10660);
nor U16288 (N_16288,N_14718,N_13236);
or U16289 (N_16289,N_13696,N_10010);
and U16290 (N_16290,N_11063,N_10472);
or U16291 (N_16291,N_10247,N_10225);
xnor U16292 (N_16292,N_14925,N_12135);
nor U16293 (N_16293,N_14664,N_12094);
nand U16294 (N_16294,N_12472,N_10248);
or U16295 (N_16295,N_14904,N_12594);
and U16296 (N_16296,N_13244,N_14547);
nor U16297 (N_16297,N_13302,N_14013);
or U16298 (N_16298,N_12133,N_10271);
nor U16299 (N_16299,N_11266,N_11844);
or U16300 (N_16300,N_14471,N_13633);
and U16301 (N_16301,N_10202,N_14335);
and U16302 (N_16302,N_13644,N_11680);
nor U16303 (N_16303,N_14348,N_13175);
or U16304 (N_16304,N_13363,N_12669);
or U16305 (N_16305,N_14470,N_14106);
nor U16306 (N_16306,N_13540,N_13133);
and U16307 (N_16307,N_14192,N_14157);
and U16308 (N_16308,N_13073,N_12684);
and U16309 (N_16309,N_10819,N_14839);
nand U16310 (N_16310,N_11571,N_13552);
xnor U16311 (N_16311,N_10091,N_12758);
or U16312 (N_16312,N_10988,N_13235);
or U16313 (N_16313,N_11943,N_11457);
and U16314 (N_16314,N_10739,N_10897);
and U16315 (N_16315,N_14407,N_10611);
nand U16316 (N_16316,N_10879,N_14840);
nor U16317 (N_16317,N_13824,N_11186);
nand U16318 (N_16318,N_13121,N_13103);
nand U16319 (N_16319,N_13225,N_13695);
and U16320 (N_16320,N_12804,N_13088);
nand U16321 (N_16321,N_14382,N_14831);
or U16322 (N_16322,N_13282,N_10201);
and U16323 (N_16323,N_11449,N_12795);
or U16324 (N_16324,N_14433,N_10442);
and U16325 (N_16325,N_12824,N_13748);
nor U16326 (N_16326,N_12455,N_13190);
nor U16327 (N_16327,N_10164,N_11177);
nand U16328 (N_16328,N_10332,N_12364);
or U16329 (N_16329,N_14797,N_12116);
and U16330 (N_16330,N_14755,N_14950);
or U16331 (N_16331,N_10068,N_11598);
nor U16332 (N_16332,N_12428,N_10163);
nor U16333 (N_16333,N_13008,N_14821);
xor U16334 (N_16334,N_12925,N_11114);
nor U16335 (N_16335,N_12937,N_14991);
nor U16336 (N_16336,N_11800,N_12308);
and U16337 (N_16337,N_10633,N_12749);
or U16338 (N_16338,N_13145,N_11060);
nor U16339 (N_16339,N_14280,N_12718);
and U16340 (N_16340,N_11190,N_11609);
or U16341 (N_16341,N_13470,N_12138);
nor U16342 (N_16342,N_13384,N_11050);
and U16343 (N_16343,N_13152,N_14218);
nand U16344 (N_16344,N_14455,N_13671);
and U16345 (N_16345,N_14069,N_10149);
and U16346 (N_16346,N_12953,N_12040);
nand U16347 (N_16347,N_13032,N_11424);
nor U16348 (N_16348,N_10986,N_14294);
and U16349 (N_16349,N_11940,N_14927);
or U16350 (N_16350,N_10356,N_10738);
xnor U16351 (N_16351,N_11191,N_12821);
nand U16352 (N_16352,N_12154,N_10334);
nor U16353 (N_16353,N_14540,N_12057);
nand U16354 (N_16354,N_10610,N_10015);
xnor U16355 (N_16355,N_11446,N_12585);
nand U16356 (N_16356,N_11933,N_14121);
nand U16357 (N_16357,N_10936,N_14534);
or U16358 (N_16358,N_12620,N_10530);
or U16359 (N_16359,N_10921,N_11778);
nand U16360 (N_16360,N_13740,N_12058);
or U16361 (N_16361,N_12141,N_11981);
or U16362 (N_16362,N_10087,N_11275);
xor U16363 (N_16363,N_13617,N_10040);
or U16364 (N_16364,N_13483,N_11676);
xnor U16365 (N_16365,N_10859,N_12345);
and U16366 (N_16366,N_10513,N_14075);
or U16367 (N_16367,N_14008,N_14715);
and U16368 (N_16368,N_14703,N_14486);
or U16369 (N_16369,N_13991,N_14142);
nand U16370 (N_16370,N_13980,N_10821);
nand U16371 (N_16371,N_12641,N_12776);
nand U16372 (N_16372,N_13687,N_11640);
or U16373 (N_16373,N_13751,N_10758);
nand U16374 (N_16374,N_12302,N_10268);
nand U16375 (N_16375,N_13423,N_11568);
nand U16376 (N_16376,N_14163,N_13069);
nor U16377 (N_16377,N_13009,N_12649);
nor U16378 (N_16378,N_11587,N_12427);
and U16379 (N_16379,N_10537,N_11313);
and U16380 (N_16380,N_12610,N_14421);
and U16381 (N_16381,N_14719,N_14633);
or U16382 (N_16382,N_10979,N_14729);
nand U16383 (N_16383,N_11027,N_11098);
or U16384 (N_16384,N_13316,N_10475);
or U16385 (N_16385,N_11209,N_12235);
or U16386 (N_16386,N_12283,N_12996);
xor U16387 (N_16387,N_10392,N_14575);
nand U16388 (N_16388,N_10154,N_14884);
nor U16389 (N_16389,N_12243,N_10372);
or U16390 (N_16390,N_13180,N_11415);
and U16391 (N_16391,N_13010,N_11491);
and U16392 (N_16392,N_14173,N_11818);
nor U16393 (N_16393,N_14686,N_11875);
nand U16394 (N_16394,N_14403,N_13439);
nand U16395 (N_16395,N_11359,N_12418);
or U16396 (N_16396,N_12337,N_12065);
and U16397 (N_16397,N_13023,N_14689);
or U16398 (N_16398,N_10711,N_11153);
nand U16399 (N_16399,N_13193,N_10095);
and U16400 (N_16400,N_14704,N_12266);
or U16401 (N_16401,N_14080,N_12355);
nand U16402 (N_16402,N_14926,N_13698);
or U16403 (N_16403,N_11206,N_14591);
xor U16404 (N_16404,N_10502,N_11095);
nor U16405 (N_16405,N_14732,N_13735);
or U16406 (N_16406,N_10754,N_14362);
or U16407 (N_16407,N_10339,N_11336);
nor U16408 (N_16408,N_10477,N_11665);
or U16409 (N_16409,N_11941,N_13488);
nor U16410 (N_16410,N_11164,N_11245);
nor U16411 (N_16411,N_11634,N_13357);
or U16412 (N_16412,N_12630,N_10486);
nand U16413 (N_16413,N_11723,N_14654);
xor U16414 (N_16414,N_10353,N_11621);
or U16415 (N_16415,N_12075,N_14210);
or U16416 (N_16416,N_14413,N_13643);
and U16417 (N_16417,N_12306,N_12967);
or U16418 (N_16418,N_14870,N_12124);
nand U16419 (N_16419,N_10377,N_14548);
nor U16420 (N_16420,N_13607,N_14447);
nand U16421 (N_16421,N_13828,N_12529);
or U16422 (N_16422,N_10452,N_11861);
nor U16423 (N_16423,N_13767,N_11030);
nand U16424 (N_16424,N_10828,N_14295);
nor U16425 (N_16425,N_10617,N_11556);
nand U16426 (N_16426,N_10985,N_12596);
or U16427 (N_16427,N_14214,N_14477);
nand U16428 (N_16428,N_14494,N_12591);
nor U16429 (N_16429,N_10933,N_10109);
nor U16430 (N_16430,N_12447,N_12686);
and U16431 (N_16431,N_10009,N_13205);
nand U16432 (N_16432,N_14685,N_14813);
nor U16433 (N_16433,N_11416,N_12056);
xor U16434 (N_16434,N_10689,N_11819);
nand U16435 (N_16435,N_10987,N_14034);
or U16436 (N_16436,N_10123,N_11237);
and U16437 (N_16437,N_14778,N_13489);
or U16438 (N_16438,N_14178,N_12023);
nor U16439 (N_16439,N_11691,N_13046);
nand U16440 (N_16440,N_12544,N_13446);
nand U16441 (N_16441,N_14123,N_14968);
or U16442 (N_16442,N_13104,N_14052);
nand U16443 (N_16443,N_14728,N_14049);
nand U16444 (N_16444,N_14007,N_12315);
and U16445 (N_16445,N_12310,N_14621);
or U16446 (N_16446,N_14537,N_14986);
and U16447 (N_16447,N_13866,N_10826);
nor U16448 (N_16448,N_10434,N_10180);
and U16449 (N_16449,N_11420,N_11810);
nor U16450 (N_16450,N_10887,N_13768);
and U16451 (N_16451,N_12077,N_10688);
nand U16452 (N_16452,N_14860,N_10929);
or U16453 (N_16453,N_10288,N_13116);
and U16454 (N_16454,N_12605,N_14442);
or U16455 (N_16455,N_14408,N_10647);
and U16456 (N_16456,N_10005,N_10640);
and U16457 (N_16457,N_14225,N_13189);
and U16458 (N_16458,N_10764,N_10656);
and U16459 (N_16459,N_13694,N_13799);
and U16460 (N_16460,N_13016,N_11232);
and U16461 (N_16461,N_11462,N_11483);
nand U16462 (N_16462,N_10062,N_14567);
or U16463 (N_16463,N_14321,N_11636);
nor U16464 (N_16464,N_12431,N_11903);
nand U16465 (N_16465,N_14881,N_14285);
and U16466 (N_16466,N_11018,N_10367);
or U16467 (N_16467,N_13668,N_10393);
or U16468 (N_16468,N_11011,N_13998);
or U16469 (N_16469,N_13451,N_13692);
nor U16470 (N_16470,N_14910,N_13999);
and U16471 (N_16471,N_12451,N_10539);
nand U16472 (N_16472,N_14995,N_14742);
nor U16473 (N_16473,N_10416,N_11295);
and U16474 (N_16474,N_13062,N_11714);
nor U16475 (N_16475,N_13464,N_10153);
and U16476 (N_16476,N_11773,N_12923);
or U16477 (N_16477,N_13074,N_12035);
nor U16478 (N_16478,N_11398,N_11176);
nand U16479 (N_16479,N_10303,N_12993);
and U16480 (N_16480,N_14108,N_13939);
and U16481 (N_16481,N_14841,N_11079);
nand U16482 (N_16482,N_14937,N_13711);
or U16483 (N_16483,N_12642,N_14769);
and U16484 (N_16484,N_12162,N_11317);
nor U16485 (N_16485,N_14610,N_14756);
nand U16486 (N_16486,N_14581,N_10760);
nand U16487 (N_16487,N_11583,N_10437);
and U16488 (N_16488,N_11379,N_10099);
nand U16489 (N_16489,N_12690,N_14057);
nand U16490 (N_16490,N_13858,N_12059);
or U16491 (N_16491,N_12171,N_12842);
and U16492 (N_16492,N_10701,N_11492);
xnor U16493 (N_16493,N_11604,N_13575);
nand U16494 (N_16494,N_10637,N_11417);
and U16495 (N_16495,N_11148,N_10116);
or U16496 (N_16496,N_10627,N_11885);
or U16497 (N_16497,N_13448,N_10460);
or U16498 (N_16498,N_12901,N_14006);
nor U16499 (N_16499,N_13406,N_13646);
or U16500 (N_16500,N_14717,N_13504);
nand U16501 (N_16501,N_11149,N_14152);
nand U16502 (N_16502,N_10691,N_13207);
nand U16503 (N_16503,N_12679,N_13749);
nor U16504 (N_16504,N_14138,N_12971);
or U16505 (N_16505,N_14632,N_10136);
nand U16506 (N_16506,N_13339,N_11827);
and U16507 (N_16507,N_12882,N_12236);
and U16508 (N_16508,N_11841,N_14174);
nand U16509 (N_16509,N_13111,N_11765);
nor U16510 (N_16510,N_13842,N_12676);
nand U16511 (N_16511,N_14482,N_13680);
and U16512 (N_16512,N_12483,N_10461);
and U16513 (N_16513,N_13840,N_14329);
or U16514 (N_16514,N_14788,N_12268);
or U16515 (N_16515,N_11522,N_10034);
nand U16516 (N_16516,N_11627,N_14683);
and U16517 (N_16517,N_10927,N_11689);
and U16518 (N_16518,N_10763,N_10695);
nand U16519 (N_16519,N_11141,N_14050);
nand U16520 (N_16520,N_13313,N_13150);
and U16521 (N_16521,N_13651,N_14342);
nor U16522 (N_16522,N_11068,N_11319);
or U16523 (N_16523,N_14466,N_12406);
nor U16524 (N_16524,N_12954,N_12599);
nor U16525 (N_16525,N_11053,N_14521);
nand U16526 (N_16526,N_13624,N_14536);
nand U16527 (N_16527,N_10114,N_10110);
or U16528 (N_16528,N_10113,N_11062);
or U16529 (N_16529,N_14940,N_10216);
nor U16530 (N_16530,N_11976,N_13732);
nand U16531 (N_16531,N_12399,N_11577);
nand U16532 (N_16532,N_10717,N_10388);
and U16533 (N_16533,N_13658,N_10681);
and U16534 (N_16534,N_12721,N_10470);
nor U16535 (N_16535,N_12333,N_13096);
nor U16536 (N_16536,N_14284,N_12999);
nor U16537 (N_16537,N_11928,N_12741);
nor U16538 (N_16538,N_13242,N_13203);
nor U16539 (N_16539,N_13445,N_12808);
xor U16540 (N_16540,N_12282,N_12763);
nor U16541 (N_16541,N_14629,N_14333);
nand U16542 (N_16542,N_13928,N_13408);
and U16543 (N_16543,N_10019,N_10424);
or U16544 (N_16544,N_11890,N_11617);
xnor U16545 (N_16545,N_13962,N_13486);
or U16546 (N_16546,N_10655,N_12305);
and U16547 (N_16547,N_13286,N_12959);
and U16548 (N_16548,N_12027,N_14130);
nor U16549 (N_16549,N_13675,N_10973);
nand U16550 (N_16550,N_10218,N_12764);
nor U16551 (N_16551,N_14339,N_12811);
and U16552 (N_16552,N_13645,N_13348);
or U16553 (N_16553,N_10961,N_13597);
nand U16554 (N_16554,N_14843,N_14680);
nand U16555 (N_16555,N_12136,N_14745);
nand U16556 (N_16556,N_11659,N_11345);
or U16557 (N_16557,N_12336,N_11871);
or U16558 (N_16558,N_12720,N_11993);
nand U16559 (N_16559,N_13107,N_13375);
nand U16560 (N_16560,N_13510,N_14393);
and U16561 (N_16561,N_14906,N_12968);
or U16562 (N_16562,N_13801,N_10412);
nor U16563 (N_16563,N_11353,N_14237);
and U16564 (N_16564,N_11490,N_14814);
nand U16565 (N_16565,N_12656,N_11205);
nand U16566 (N_16566,N_13417,N_14376);
and U16567 (N_16567,N_11161,N_10727);
and U16568 (N_16568,N_12322,N_10396);
nor U16569 (N_16569,N_10381,N_11537);
nand U16570 (N_16570,N_13837,N_13789);
nor U16571 (N_16571,N_11559,N_11376);
nor U16572 (N_16572,N_14677,N_11808);
nor U16573 (N_16573,N_10141,N_12814);
or U16574 (N_16574,N_11942,N_10993);
nor U16575 (N_16575,N_12249,N_13321);
nor U16576 (N_16576,N_10190,N_10405);
nor U16577 (N_16577,N_12748,N_12476);
nand U16578 (N_16578,N_11701,N_11487);
and U16579 (N_16579,N_12556,N_11029);
or U16580 (N_16580,N_11015,N_11493);
nor U16581 (N_16581,N_14657,N_11402);
nand U16582 (N_16582,N_10257,N_13817);
nand U16583 (N_16583,N_14724,N_13092);
or U16584 (N_16584,N_11662,N_11997);
nor U16585 (N_16585,N_14988,N_11322);
and U16586 (N_16586,N_12429,N_12532);
or U16587 (N_16587,N_13124,N_14759);
nand U16588 (N_16588,N_10743,N_13359);
nor U16589 (N_16589,N_11076,N_10756);
or U16590 (N_16590,N_13527,N_10850);
and U16591 (N_16591,N_10369,N_11445);
and U16592 (N_16592,N_12417,N_12553);
nor U16593 (N_16593,N_12369,N_12790);
nand U16594 (N_16594,N_10055,N_13055);
or U16595 (N_16595,N_11014,N_13381);
xnor U16596 (N_16596,N_11929,N_12955);
nor U16597 (N_16597,N_14119,N_13534);
and U16598 (N_16598,N_12054,N_11173);
and U16599 (N_16599,N_12816,N_10326);
and U16600 (N_16600,N_11829,N_12412);
and U16601 (N_16601,N_12984,N_13743);
nand U16602 (N_16602,N_13472,N_12688);
or U16603 (N_16603,N_12916,N_13352);
nand U16604 (N_16604,N_12217,N_13976);
nor U16605 (N_16605,N_14089,N_12699);
or U16606 (N_16606,N_11202,N_14700);
nor U16607 (N_16607,N_10516,N_12952);
nor U16608 (N_16608,N_13378,N_14254);
and U16609 (N_16609,N_12853,N_13034);
or U16610 (N_16610,N_12985,N_12560);
or U16611 (N_16611,N_14272,N_10923);
nand U16612 (N_16612,N_13745,N_10592);
or U16613 (N_16613,N_13362,N_14746);
or U16614 (N_16614,N_10529,N_11387);
and U16615 (N_16615,N_14064,N_10822);
or U16616 (N_16616,N_14774,N_11702);
nor U16617 (N_16617,N_11233,N_14039);
and U16618 (N_16618,N_14608,N_12482);
nand U16619 (N_16619,N_14618,N_14961);
or U16620 (N_16620,N_14290,N_13461);
nor U16621 (N_16621,N_10192,N_11494);
and U16622 (N_16622,N_13369,N_13474);
and U16623 (N_16623,N_11285,N_12089);
nor U16624 (N_16624,N_14907,N_12199);
and U16625 (N_16625,N_14504,N_10413);
nor U16626 (N_16626,N_12347,N_13606);
or U16627 (N_16627,N_14085,N_14625);
nand U16628 (N_16628,N_10509,N_11533);
nand U16629 (N_16629,N_14750,N_10117);
and U16630 (N_16630,N_10765,N_10619);
nor U16631 (N_16631,N_12164,N_10946);
and U16632 (N_16632,N_12439,N_10544);
nor U16633 (N_16633,N_13957,N_11346);
and U16634 (N_16634,N_14923,N_12033);
and U16635 (N_16635,N_11682,N_10480);
nand U16636 (N_16636,N_11909,N_13020);
nand U16637 (N_16637,N_12001,N_14030);
nor U16638 (N_16638,N_12772,N_11586);
nor U16639 (N_16639,N_13165,N_10546);
and U16640 (N_16640,N_12875,N_13398);
and U16641 (N_16641,N_10491,N_13582);
or U16642 (N_16642,N_13734,N_13800);
and U16643 (N_16643,N_14058,N_11973);
xor U16644 (N_16644,N_12934,N_11927);
and U16645 (N_16645,N_14005,N_12276);
or U16646 (N_16646,N_14033,N_10417);
or U16647 (N_16647,N_10713,N_10839);
or U16648 (N_16648,N_11261,N_13871);
or U16649 (N_16649,N_14736,N_12803);
nor U16650 (N_16650,N_10241,N_13997);
xor U16651 (N_16651,N_14772,N_12365);
or U16652 (N_16652,N_11374,N_12022);
or U16653 (N_16653,N_10735,N_10435);
or U16654 (N_16654,N_10297,N_10928);
or U16655 (N_16655,N_12865,N_13440);
xor U16656 (N_16656,N_11811,N_11341);
or U16657 (N_16657,N_12910,N_13725);
nand U16658 (N_16658,N_13227,N_11006);
and U16659 (N_16659,N_13716,N_11774);
and U16660 (N_16660,N_12117,N_11607);
or U16661 (N_16661,N_10142,N_13462);
or U16662 (N_16662,N_12181,N_12339);
nand U16663 (N_16663,N_11361,N_10499);
and U16664 (N_16664,N_13503,N_14770);
or U16665 (N_16665,N_11760,N_11399);
nand U16666 (N_16666,N_14331,N_12311);
and U16667 (N_16667,N_13465,N_13775);
or U16668 (N_16668,N_12994,N_13932);
nor U16669 (N_16669,N_11288,N_12719);
and U16670 (N_16670,N_12950,N_13496);
or U16671 (N_16671,N_14176,N_12904);
and U16672 (N_16672,N_14487,N_13878);
or U16673 (N_16673,N_10101,N_12424);
and U16674 (N_16674,N_13602,N_14852);
nor U16675 (N_16675,N_12997,N_11337);
or U16676 (N_16676,N_10600,N_12119);
nor U16677 (N_16677,N_11434,N_11546);
nand U16678 (N_16678,N_11785,N_12093);
nor U16679 (N_16679,N_11174,N_10217);
nor U16680 (N_16680,N_14468,N_12511);
nor U16681 (N_16681,N_10077,N_10212);
nor U16682 (N_16682,N_10598,N_11070);
nor U16683 (N_16683,N_11992,N_11848);
or U16684 (N_16684,N_12197,N_11260);
or U16685 (N_16685,N_10028,N_14406);
and U16686 (N_16686,N_10131,N_10543);
nand U16687 (N_16687,N_14764,N_11044);
xnor U16688 (N_16688,N_11991,N_12458);
nand U16689 (N_16689,N_10675,N_12165);
and U16690 (N_16690,N_14876,N_13667);
nor U16691 (N_16691,N_11622,N_10032);
nor U16692 (N_16692,N_13571,N_10251);
and U16693 (N_16693,N_11138,N_14231);
nor U16694 (N_16694,N_11211,N_12713);
nor U16695 (N_16695,N_11724,N_11082);
and U16696 (N_16696,N_14045,N_10782);
or U16697 (N_16697,N_12496,N_12363);
or U16698 (N_16698,N_13065,N_12487);
and U16699 (N_16699,N_10399,N_13530);
nand U16700 (N_16700,N_14301,N_11442);
and U16701 (N_16701,N_12006,N_11103);
or U16702 (N_16702,N_11524,N_14777);
nand U16703 (N_16703,N_12395,N_10536);
nor U16704 (N_16704,N_13619,N_14115);
or U16705 (N_16705,N_14812,N_14522);
nor U16706 (N_16706,N_11151,N_14070);
nor U16707 (N_16707,N_14300,N_13869);
and U16708 (N_16708,N_12375,N_12076);
and U16709 (N_16709,N_10613,N_12847);
or U16710 (N_16710,N_12113,N_12407);
nor U16711 (N_16711,N_13576,N_12584);
and U16712 (N_16712,N_13436,N_14918);
or U16713 (N_16713,N_10301,N_10421);
and U16714 (N_16714,N_12624,N_10808);
nand U16715 (N_16715,N_12409,N_13006);
nand U16716 (N_16716,N_10832,N_13721);
or U16717 (N_16717,N_14563,N_14999);
nor U16718 (N_16718,N_14244,N_11092);
nand U16719 (N_16719,N_10609,N_13138);
xor U16720 (N_16720,N_11748,N_13985);
or U16721 (N_16721,N_10171,N_11679);
nor U16722 (N_16722,N_14519,N_14915);
and U16723 (N_16723,N_12193,N_14449);
or U16724 (N_16724,N_12026,N_12736);
and U16725 (N_16725,N_13433,N_12242);
and U16726 (N_16726,N_10715,N_13547);
and U16727 (N_16727,N_11124,N_13086);
nor U16728 (N_16728,N_12958,N_14361);
nor U16729 (N_16729,N_12706,N_10443);
nand U16730 (N_16730,N_11162,N_12207);
and U16731 (N_16731,N_10047,N_13559);
nand U16732 (N_16732,N_10306,N_10256);
and U16733 (N_16733,N_10896,N_13511);
nand U16734 (N_16734,N_12640,N_14600);
nor U16735 (N_16735,N_14061,N_11947);
or U16736 (N_16736,N_14296,N_14079);
nand U16737 (N_16737,N_13989,N_13275);
and U16738 (N_16738,N_14017,N_12921);
nor U16739 (N_16739,N_10317,N_12988);
or U16740 (N_16740,N_11327,N_11343);
and U16741 (N_16741,N_13509,N_10560);
and U16742 (N_16742,N_11222,N_11525);
or U16743 (N_16743,N_10254,N_10422);
nor U16744 (N_16744,N_12509,N_12674);
nand U16745 (N_16745,N_10746,N_12963);
and U16746 (N_16746,N_13389,N_13773);
nor U16747 (N_16747,N_14467,N_13229);
nor U16748 (N_16748,N_14204,N_13387);
nand U16749 (N_16749,N_10994,N_10712);
or U16750 (N_16750,N_12103,N_11091);
nand U16751 (N_16751,N_12391,N_10525);
nor U16752 (N_16752,N_10578,N_11779);
nand U16753 (N_16753,N_10575,N_13204);
or U16754 (N_16754,N_11855,N_11075);
nor U16755 (N_16755,N_14344,N_13620);
nor U16756 (N_16756,N_13585,N_10884);
and U16757 (N_16757,N_14932,N_12502);
nand U16758 (N_16758,N_10702,N_11046);
and U16759 (N_16759,N_10983,N_13161);
or U16760 (N_16760,N_13787,N_11287);
or U16761 (N_16761,N_13572,N_11857);
and U16762 (N_16762,N_10556,N_13287);
or U16763 (N_16763,N_14463,N_12195);
or U16764 (N_16764,N_11834,N_14825);
nor U16765 (N_16765,N_12637,N_12224);
nand U16766 (N_16766,N_11878,N_12048);
nand U16767 (N_16767,N_10761,N_14055);
nand U16768 (N_16768,N_10371,N_11140);
and U16769 (N_16769,N_10184,N_11429);
nor U16770 (N_16770,N_11334,N_10588);
nor U16771 (N_16771,N_11500,N_14103);
nand U16772 (N_16772,N_10182,N_14975);
or U16773 (N_16773,N_12519,N_11717);
nand U16774 (N_16774,N_14087,N_14334);
and U16775 (N_16775,N_11118,N_10729);
xnor U16776 (N_16776,N_11835,N_11923);
nand U16777 (N_16777,N_13054,N_12508);
or U16778 (N_16778,N_12290,N_11688);
and U16779 (N_16779,N_12184,N_11217);
nand U16780 (N_16780,N_11436,N_13356);
or U16781 (N_16781,N_10584,N_12031);
and U16782 (N_16782,N_11248,N_12717);
or U16783 (N_16783,N_10433,N_11558);
and U16784 (N_16784,N_13269,N_12452);
nor U16785 (N_16785,N_14427,N_13531);
or U16786 (N_16786,N_11930,N_14450);
or U16787 (N_16787,N_11729,N_13058);
nand U16788 (N_16788,N_10076,N_12781);
and U16789 (N_16789,N_13665,N_13153);
nor U16790 (N_16790,N_13535,N_13155);
nand U16791 (N_16791,N_12297,N_12542);
nand U16792 (N_16792,N_14576,N_10538);
or U16793 (N_16793,N_13329,N_13036);
nand U16794 (N_16794,N_11668,N_12976);
or U16795 (N_16795,N_11711,N_12272);
nand U16796 (N_16796,N_12929,N_13368);
and U16797 (N_16797,N_12317,N_13301);
nand U16798 (N_16798,N_12829,N_12238);
nor U16799 (N_16799,N_10020,N_13826);
nor U16800 (N_16800,N_13927,N_14887);
and U16801 (N_16801,N_11286,N_12990);
and U16802 (N_16802,N_12709,N_13268);
or U16803 (N_16803,N_10945,N_13970);
nand U16804 (N_16804,N_14779,N_14136);
or U16805 (N_16805,N_12956,N_13382);
or U16806 (N_16806,N_11969,N_11669);
nand U16807 (N_16807,N_10228,N_13679);
nand U16808 (N_16808,N_12280,N_14882);
or U16809 (N_16809,N_10703,N_14431);
or U16810 (N_16810,N_11255,N_11418);
nor U16811 (N_16811,N_11908,N_11949);
or U16812 (N_16812,N_13744,N_11653);
nor U16813 (N_16813,N_13468,N_13139);
and U16814 (N_16814,N_12846,N_12715);
nand U16815 (N_16815,N_11570,N_10108);
nor U16816 (N_16816,N_10648,N_13761);
or U16817 (N_16817,N_14924,N_11081);
nor U16818 (N_16818,N_12631,N_11812);
nor U16819 (N_16819,N_11703,N_10899);
nand U16820 (N_16820,N_13755,N_12785);
and U16821 (N_16821,N_10197,N_11096);
nand U16822 (N_16822,N_12488,N_10008);
or U16823 (N_16823,N_13360,N_13403);
or U16824 (N_16824,N_10226,N_11732);
and U16825 (N_16825,N_12789,N_12080);
nand U16826 (N_16826,N_11979,N_13344);
and U16827 (N_16827,N_13432,N_10955);
and U16828 (N_16828,N_12204,N_10189);
and U16829 (N_16829,N_10157,N_12782);
and U16830 (N_16830,N_10102,N_13105);
nand U16831 (N_16831,N_10012,N_12666);
nor U16832 (N_16832,N_13803,N_12702);
or U16833 (N_16833,N_10140,N_13248);
and U16834 (N_16834,N_12647,N_13013);
and U16835 (N_16835,N_12044,N_13836);
or U16836 (N_16836,N_14195,N_11907);
and U16837 (N_16837,N_10798,N_11441);
nor U16838 (N_16838,N_14974,N_12351);
nand U16839 (N_16839,N_13261,N_14384);
and U16840 (N_16840,N_12545,N_11562);
and U16841 (N_16841,N_12258,N_12697);
nor U16842 (N_16842,N_10275,N_12146);
and U16843 (N_16843,N_13157,N_13093);
nor U16844 (N_16844,N_10206,N_11333);
and U16845 (N_16845,N_14952,N_12660);
nand U16846 (N_16846,N_13231,N_10398);
nand U16847 (N_16847,N_13413,N_14252);
xnor U16848 (N_16848,N_13068,N_13850);
nor U16849 (N_16849,N_10740,N_10253);
nand U16850 (N_16850,N_14020,N_12098);
nand U16851 (N_16851,N_11438,N_12420);
or U16852 (N_16852,N_13131,N_14086);
or U16853 (N_16853,N_13757,N_13499);
and U16854 (N_16854,N_13090,N_10757);
or U16855 (N_16855,N_12396,N_10687);
or U16856 (N_16856,N_14282,N_12614);
nor U16857 (N_16857,N_13025,N_11769);
and U16858 (N_16858,N_10415,N_12843);
and U16859 (N_16859,N_12769,N_11498);
nand U16860 (N_16860,N_13031,N_12851);
nand U16861 (N_16861,N_11672,N_11530);
and U16862 (N_16862,N_14807,N_13941);
and U16863 (N_16863,N_11911,N_13140);
or U16864 (N_16864,N_13762,N_11633);
nand U16865 (N_16865,N_14789,N_13573);
nand U16866 (N_16866,N_14118,N_13960);
nor U16867 (N_16867,N_12253,N_14135);
and U16868 (N_16868,N_14551,N_14651);
or U16869 (N_16869,N_14420,N_10195);
and U16870 (N_16870,N_14129,N_10549);
and U16871 (N_16871,N_11946,N_14278);
and U16872 (N_16872,N_14349,N_11856);
or U16873 (N_16873,N_12471,N_12088);
nand U16874 (N_16874,N_14531,N_12359);
or U16875 (N_16875,N_14963,N_10580);
nand U16876 (N_16876,N_11168,N_11535);
nor U16877 (N_16877,N_14081,N_11960);
and U16878 (N_16878,N_11658,N_14602);
or U16879 (N_16879,N_13904,N_10262);
and U16880 (N_16880,N_13529,N_14737);
nand U16881 (N_16881,N_14969,N_14243);
and U16882 (N_16882,N_11289,N_10178);
nor U16883 (N_16883,N_12152,N_11904);
nor U16884 (N_16884,N_12218,N_13845);
and U16885 (N_16885,N_10468,N_11825);
nand U16886 (N_16886,N_10340,N_10615);
or U16887 (N_16887,N_13279,N_13851);
nand U16888 (N_16888,N_14358,N_12546);
nand U16889 (N_16889,N_11677,N_10977);
and U16890 (N_16890,N_10805,N_13182);
and U16891 (N_16891,N_11414,N_10057);
and U16892 (N_16892,N_12909,N_13545);
or U16893 (N_16893,N_13246,N_13859);
nor U16894 (N_16894,N_14193,N_12432);
or U16895 (N_16895,N_11618,N_11223);
nor U16896 (N_16896,N_13262,N_13198);
nor U16897 (N_16897,N_10550,N_12227);
nor U16898 (N_16898,N_11685,N_11220);
nand U16899 (N_16899,N_11865,N_13612);
and U16900 (N_16900,N_11606,N_12318);
or U16901 (N_16901,N_11803,N_14775);
nor U16902 (N_16902,N_14059,N_10635);
or U16903 (N_16903,N_12727,N_14372);
nand U16904 (N_16904,N_11893,N_14419);
nand U16905 (N_16905,N_14153,N_13676);
nand U16906 (N_16906,N_14765,N_12730);
and U16907 (N_16907,N_11430,N_10130);
nand U16908 (N_16908,N_14241,N_10320);
nor U16909 (N_16909,N_10081,N_13593);
nand U16910 (N_16910,N_13508,N_11257);
and U16911 (N_16911,N_13726,N_11615);
nand U16912 (N_16912,N_10204,N_10122);
or U16913 (N_16913,N_10360,N_12091);
or U16914 (N_16914,N_11444,N_11016);
nor U16915 (N_16915,N_14557,N_14767);
nor U16916 (N_16916,N_12295,N_10490);
nand U16917 (N_16917,N_14395,N_10266);
nand U16918 (N_16918,N_14053,N_11866);
xnor U16919 (N_16919,N_14698,N_14578);
nor U16920 (N_16920,N_10249,N_14238);
nand U16921 (N_16921,N_13281,N_10579);
and U16922 (N_16922,N_10072,N_11481);
or U16923 (N_16923,N_11362,N_13990);
nand U16924 (N_16924,N_13883,N_10086);
nor U16925 (N_16925,N_11392,N_13041);
nand U16926 (N_16926,N_11816,N_14543);
or U16927 (N_16927,N_11935,N_14446);
or U16928 (N_16928,N_13532,N_14623);
nor U16929 (N_16929,N_13380,N_13077);
and U16930 (N_16930,N_14733,N_11509);
xor U16931 (N_16931,N_14705,N_10400);
or U16932 (N_16932,N_14989,N_10874);
and U16933 (N_16933,N_13026,N_10639);
nor U16934 (N_16934,N_11921,N_12617);
nand U16935 (N_16935,N_11300,N_13568);
nor U16936 (N_16936,N_10784,N_13678);
nor U16937 (N_16937,N_13042,N_10380);
and U16938 (N_16938,N_14260,N_12915);
or U16939 (N_16939,N_14066,N_13781);
nand U16940 (N_16940,N_12541,N_14804);
nand U16941 (N_16941,N_10027,N_13756);
or U16942 (N_16942,N_10512,N_11554);
or U16943 (N_16943,N_11195,N_10817);
nor U16944 (N_16944,N_13948,N_10855);
nor U16945 (N_16945,N_14426,N_13752);
nand U16946 (N_16946,N_11010,N_10541);
nor U16947 (N_16947,N_10508,N_11747);
nor U16948 (N_16948,N_10440,N_10018);
xnor U16949 (N_16949,N_12830,N_12612);
or U16950 (N_16950,N_11352,N_13882);
and U16951 (N_16951,N_12820,N_11728);
nor U16952 (N_16952,N_12911,N_10998);
or U16953 (N_16953,N_11520,N_13012);
nand U16954 (N_16954,N_14098,N_11796);
and U16955 (N_16955,N_14929,N_14126);
nand U16956 (N_16956,N_11312,N_14785);
and U16957 (N_16957,N_11043,N_11802);
or U16958 (N_16958,N_11203,N_14854);
and U16959 (N_16959,N_13040,N_10042);
nand U16960 (N_16960,N_10375,N_12324);
or U16961 (N_16961,N_12045,N_12931);
and U16962 (N_16962,N_14561,N_11798);
or U16963 (N_16963,N_10411,N_11412);
or U16964 (N_16964,N_12320,N_11218);
nand U16965 (N_16965,N_10169,N_13134);
nor U16966 (N_16966,N_13630,N_14094);
or U16967 (N_16967,N_14261,N_11738);
xor U16968 (N_16968,N_13791,N_10265);
and U16969 (N_16969,N_13089,N_10161);
or U16970 (N_16970,N_10313,N_12478);
or U16971 (N_16971,N_13255,N_14847);
or U16972 (N_16972,N_10569,N_14202);
or U16973 (N_16973,N_12754,N_10732);
nor U16974 (N_16974,N_11958,N_14293);
nor U16975 (N_16975,N_13011,N_11931);
nor U16976 (N_16976,N_10067,N_14672);
nand U16977 (N_16977,N_14781,N_11552);
and U16978 (N_16978,N_12590,N_11770);
nor U16979 (N_16979,N_14319,N_11342);
and U16980 (N_16980,N_13933,N_14097);
or U16981 (N_16981,N_14368,N_14800);
xor U16982 (N_16982,N_14232,N_12751);
and U16983 (N_16983,N_11582,N_12725);
nor U16984 (N_16984,N_14330,N_14803);
nor U16985 (N_16985,N_14630,N_14829);
and U16986 (N_16986,N_14141,N_11529);
nor U16987 (N_16987,N_10281,N_10260);
or U16988 (N_16988,N_14196,N_13365);
or U16989 (N_16989,N_11066,N_10869);
nand U16990 (N_16990,N_10720,N_13891);
nor U16991 (N_16991,N_14935,N_14429);
and U16992 (N_16992,N_12081,N_11786);
nand U16993 (N_16993,N_10679,N_14027);
or U16994 (N_16994,N_11912,N_11799);
nand U16995 (N_16995,N_12583,N_13071);
nor U16996 (N_16996,N_11467,N_13361);
nand U16997 (N_16997,N_12877,N_12263);
and U16998 (N_16998,N_13434,N_13753);
or U16999 (N_16999,N_13515,N_13614);
nor U17000 (N_17000,N_13449,N_10944);
nor U17001 (N_17001,N_11962,N_10014);
or U17002 (N_17002,N_11744,N_11489);
and U17003 (N_17003,N_12203,N_13896);
nor U17004 (N_17004,N_12839,N_11204);
and U17005 (N_17005,N_12654,N_11401);
nand U17006 (N_17006,N_10999,N_10789);
nor U17007 (N_17007,N_11635,N_12678);
nor U17008 (N_17008,N_13307,N_10545);
and U17009 (N_17009,N_13982,N_13969);
nor U17010 (N_17010,N_10978,N_10895);
and U17011 (N_17011,N_12362,N_10692);
nor U17012 (N_17012,N_12284,N_14062);
nor U17013 (N_17013,N_14980,N_12732);
nand U17014 (N_17014,N_11895,N_12433);
nand U17015 (N_17015,N_11306,N_10563);
nand U17016 (N_17016,N_11793,N_12376);
nand U17017 (N_17017,N_12470,N_10844);
nor U17018 (N_17018,N_10890,N_14667);
nand U17019 (N_17019,N_12914,N_10387);
nor U17020 (N_17020,N_10318,N_10875);
or U17021 (N_17021,N_10745,N_10902);
nand U17022 (N_17022,N_14790,N_14224);
nand U17023 (N_17023,N_12416,N_11534);
and U17024 (N_17024,N_14597,N_13336);
or U17025 (N_17025,N_13185,N_12499);
or U17026 (N_17026,N_13412,N_11536);
nor U17027 (N_17027,N_12579,N_13967);
and U17028 (N_17028,N_14472,N_11603);
or U17029 (N_17029,N_12757,N_13780);
nor U17030 (N_17030,N_13659,N_12943);
and U17031 (N_17031,N_11504,N_11817);
and U17032 (N_17032,N_12394,N_10368);
nand U17033 (N_17033,N_12694,N_11764);
nand U17034 (N_17034,N_10282,N_14864);
or U17035 (N_17035,N_12876,N_11036);
nor U17036 (N_17036,N_11891,N_13570);
nor U17037 (N_17037,N_11309,N_10643);
and U17038 (N_17038,N_10389,N_11564);
or U17039 (N_17039,N_12084,N_12155);
and U17040 (N_17040,N_13888,N_13101);
xnor U17041 (N_17041,N_10604,N_10900);
nor U17042 (N_17042,N_10564,N_11674);
or U17043 (N_17043,N_13693,N_10709);
and U17044 (N_17044,N_13911,N_10783);
and U17045 (N_17045,N_11837,N_11109);
nand U17046 (N_17046,N_11831,N_10365);
or U17047 (N_17047,N_12523,N_10035);
nand U17048 (N_17048,N_11054,N_14708);
and U17049 (N_17049,N_13961,N_14538);
and U17050 (N_17050,N_11246,N_11999);
nor U17051 (N_17051,N_10227,N_11393);
and U17052 (N_17052,N_13392,N_14739);
or U17053 (N_17053,N_14434,N_12683);
nor U17054 (N_17054,N_11432,N_11902);
and U17055 (N_17055,N_13126,N_10078);
nand U17056 (N_17056,N_14151,N_14312);
nor U17057 (N_17057,N_12024,N_14213);
nor U17058 (N_17058,N_10013,N_13637);
and U17059 (N_17059,N_14838,N_11335);
or U17060 (N_17060,N_14894,N_11772);
or U17061 (N_17061,N_12186,N_14255);
nand U17062 (N_17062,N_10242,N_14181);
xor U17063 (N_17063,N_13563,N_14150);
and U17064 (N_17064,N_12643,N_13591);
nor U17065 (N_17065,N_12891,N_14366);
xor U17066 (N_17066,N_14886,N_13587);
nor U17067 (N_17067,N_14350,N_12693);
xor U17068 (N_17068,N_14749,N_13955);
and U17069 (N_17069,N_13267,N_10418);
or U17070 (N_17070,N_13334,N_11464);
and U17071 (N_17071,N_14102,N_14198);
or U17072 (N_17072,N_13885,N_12344);
nand U17073 (N_17073,N_13340,N_11282);
nand U17074 (N_17074,N_10825,N_10456);
and U17075 (N_17075,N_14544,N_11363);
nor U17076 (N_17076,N_13109,N_10148);
nor U17077 (N_17077,N_13674,N_11937);
or U17078 (N_17078,N_10186,N_13981);
nor U17079 (N_17079,N_13146,N_14355);
nand U17080 (N_17080,N_10705,N_10925);
nor U17081 (N_17081,N_12385,N_13688);
and U17082 (N_17082,N_11437,N_11107);
nor U17083 (N_17083,N_13396,N_14579);
and U17084 (N_17084,N_12087,N_13830);
or U17085 (N_17085,N_13200,N_13164);
or U17086 (N_17086,N_14439,N_12083);
or U17087 (N_17087,N_14444,N_14369);
and U17088 (N_17088,N_10049,N_14688);
or U17089 (N_17089,N_14517,N_13210);
or U17090 (N_17090,N_10233,N_14659);
nand U17091 (N_17091,N_10791,N_11234);
and U17092 (N_17092,N_11221,N_10673);
and U17093 (N_17093,N_13021,N_13873);
nand U17094 (N_17094,N_11331,N_13776);
or U17095 (N_17095,N_12349,N_13513);
nor U17096 (N_17096,N_10773,N_13632);
or U17097 (N_17097,N_14381,N_12219);
or U17098 (N_17098,N_10230,N_10064);
nand U17099 (N_17099,N_10762,N_12348);
and U17100 (N_17100,N_13528,N_10658);
xnor U17101 (N_17101,N_11460,N_14386);
and U17102 (N_17102,N_12618,N_12559);
or U17103 (N_17103,N_11567,N_12947);
or U17104 (N_17104,N_14851,N_14303);
or U17105 (N_17105,N_13918,N_12438);
and U17106 (N_17106,N_12574,N_12156);
nand U17107 (N_17107,N_10958,N_14898);
or U17108 (N_17108,N_12148,N_13049);
or U17109 (N_17109,N_13984,N_10273);
nor U17110 (N_17110,N_10261,N_14068);
nand U17111 (N_17111,N_10300,N_11413);
or U17112 (N_17112,N_12980,N_11638);
xor U17113 (N_17113,N_11710,N_11675);
or U17114 (N_17114,N_10198,N_12695);
nor U17115 (N_17115,N_14877,N_14593);
nor U17116 (N_17116,N_13176,N_11854);
nor U17117 (N_17117,N_10084,N_13487);
and U17118 (N_17118,N_12014,N_14711);
or U17119 (N_17119,N_14067,N_12628);
and U17120 (N_17120,N_13209,N_14251);
or U17121 (N_17121,N_12277,N_12112);
nor U17122 (N_17122,N_14653,N_12279);
nor U17123 (N_17123,N_13805,N_12074);
or U17124 (N_17124,N_10219,N_10383);
nor U17125 (N_17125,N_10277,N_10236);
and U17126 (N_17126,N_13769,N_11994);
nand U17127 (N_17127,N_12405,N_10520);
or U17128 (N_17128,N_13163,N_11971);
and U17129 (N_17129,N_12619,N_10155);
xnor U17130 (N_17130,N_11450,N_11165);
nand U17131 (N_17131,N_11231,N_14508);
or U17132 (N_17132,N_10548,N_13371);
and U17133 (N_17133,N_11471,N_13831);
nor U17134 (N_17134,N_13323,N_14842);
and U17135 (N_17135,N_12018,N_13853);
nand U17136 (N_17136,N_10166,N_14206);
nor U17137 (N_17137,N_12974,N_12733);
nor U17138 (N_17138,N_10048,N_10498);
and U17139 (N_17139,N_10975,N_13455);
or U17140 (N_17140,N_14913,N_13986);
and U17141 (N_17141,N_14353,N_11901);
nand U17142 (N_17142,N_12555,N_14396);
nand U17143 (N_17143,N_13079,N_14483);
nor U17144 (N_17144,N_11956,N_11784);
nand U17145 (N_17145,N_14669,N_12108);
and U17146 (N_17146,N_11952,N_11479);
or U17147 (N_17147,N_14760,N_11009);
and U17148 (N_17148,N_13621,N_11452);
nor U17149 (N_17149,N_14091,N_10351);
or U17150 (N_17150,N_10714,N_14857);
or U17151 (N_17151,N_11244,N_13718);
or U17152 (N_17152,N_12414,N_11117);
nand U17153 (N_17153,N_14796,N_10733);
and U17154 (N_17154,N_10358,N_13815);
and U17155 (N_17155,N_13335,N_12863);
and U17156 (N_17156,N_11965,N_10533);
or U17157 (N_17157,N_10534,N_12812);
or U17158 (N_17158,N_11020,N_12379);
nor U17159 (N_17159,N_11439,N_11771);
nor U17160 (N_17160,N_10831,N_14124);
nand U17161 (N_17161,N_11448,N_13857);
nand U17162 (N_17162,N_13611,N_13589);
and U17163 (N_17163,N_12778,N_12662);
or U17164 (N_17164,N_14190,N_14997);
nor U17165 (N_17165,N_14554,N_12269);
or U17166 (N_17166,N_10685,N_12570);
xor U17167 (N_17167,N_14875,N_12442);
or U17168 (N_17168,N_12536,N_14702);
and U17169 (N_17169,N_11652,N_12852);
and U17170 (N_17170,N_14288,N_13167);
xor U17171 (N_17171,N_12924,N_12017);
nor U17172 (N_17172,N_14184,N_11624);
or U17173 (N_17173,N_14340,N_14956);
or U17174 (N_17174,N_10951,N_11843);
nand U17175 (N_17175,N_10350,N_13212);
nand U17176 (N_17176,N_13586,N_12454);
nor U17177 (N_17177,N_11086,N_10742);
or U17178 (N_17178,N_12149,N_12211);
xnor U17179 (N_17179,N_13616,N_12638);
nand U17180 (N_17180,N_14943,N_12667);
and U17181 (N_17181,N_12892,N_11780);
and U17182 (N_17182,N_13835,N_11984);
nor U17183 (N_17183,N_13626,N_12436);
and U17184 (N_17184,N_13113,N_14409);
and U17185 (N_17185,N_12029,N_10285);
nor U17186 (N_17186,N_12817,N_10847);
or U17187 (N_17187,N_12745,N_10515);
xnor U17188 (N_17188,N_11370,N_14527);
nor U17189 (N_17189,N_12241,N_11463);
xnor U17190 (N_17190,N_12648,N_14850);
nand U17191 (N_17191,N_13199,N_12944);
nor U17192 (N_17192,N_10205,N_11862);
nand U17193 (N_17193,N_10287,N_12498);
and U17194 (N_17194,N_13443,N_14443);
nor U17195 (N_17195,N_11057,N_12609);
or U17196 (N_17196,N_14835,N_12043);
nor U17197 (N_17197,N_11610,N_13447);
and U17198 (N_17198,N_14587,N_10038);
or U17199 (N_17199,N_13143,N_13338);
and U17200 (N_17200,N_12871,N_14199);
or U17201 (N_17201,N_10519,N_11791);
or U17202 (N_17202,N_12862,N_13951);
nand U17203 (N_17203,N_12551,N_14931);
and U17204 (N_17204,N_10971,N_13325);
nor U17205 (N_17205,N_10172,N_12936);
and U17206 (N_17206,N_12905,N_11549);
nand U17207 (N_17207,N_11886,N_13438);
or U17208 (N_17208,N_11551,N_14639);
nand U17209 (N_17209,N_13311,N_12940);
nand U17210 (N_17210,N_12090,N_12540);
and U17211 (N_17211,N_12109,N_10021);
nand U17212 (N_17212,N_10953,N_13598);
nand U17213 (N_17213,N_12510,N_10315);
and U17214 (N_17214,N_11611,N_11814);
or U17215 (N_17215,N_14981,N_10119);
or U17216 (N_17216,N_10118,N_10722);
nor U17217 (N_17217,N_10949,N_12682);
nand U17218 (N_17218,N_12907,N_11372);
and U17219 (N_17219,N_13112,N_10694);
or U17220 (N_17220,N_14908,N_11572);
nor U17221 (N_17221,N_13724,N_13052);
nand U17222 (N_17222,N_12187,N_14400);
xnor U17223 (N_17223,N_13705,N_14606);
or U17224 (N_17224,N_11696,N_13704);
or U17225 (N_17225,N_12870,N_12801);
nor U17226 (N_17226,N_14159,N_12383);
nor U17227 (N_17227,N_14424,N_12828);
and U17228 (N_17228,N_14496,N_13963);
nor U17229 (N_17229,N_12760,N_11157);
nor U17230 (N_17230,N_11386,N_10577);
nor U17231 (N_17231,N_11805,N_11200);
nor U17232 (N_17232,N_14933,N_13936);
or U17233 (N_17233,N_12389,N_10849);
or U17234 (N_17234,N_12019,N_10621);
or U17235 (N_17235,N_12225,N_14113);
nor U17236 (N_17236,N_14872,N_13860);
and U17237 (N_17237,N_11259,N_10667);
and U17238 (N_17238,N_14912,N_10103);
nand U17239 (N_17239,N_11184,N_14879);
nand U17240 (N_17240,N_10406,N_12687);
xor U17241 (N_17241,N_11299,N_13802);
and U17242 (N_17242,N_13258,N_10774);
nand U17243 (N_17243,N_10750,N_14310);
and U17244 (N_17244,N_11073,N_14905);
or U17245 (N_17245,N_11013,N_10497);
xnor U17246 (N_17246,N_10659,N_14970);
and U17247 (N_17247,N_12833,N_14104);
nor U17248 (N_17248,N_11508,N_11332);
nor U17249 (N_17249,N_14964,N_12861);
or U17250 (N_17250,N_11104,N_10803);
nand U17251 (N_17251,N_13001,N_10489);
and U17252 (N_17252,N_13330,N_11900);
or U17253 (N_17253,N_14004,N_13237);
or U17254 (N_17254,N_12825,N_14388);
nand U17255 (N_17255,N_14934,N_13603);
and U17256 (N_17256,N_11853,N_12837);
nor U17257 (N_17257,N_11024,N_13638);
and U17258 (N_17258,N_12229,N_11304);
xor U17259 (N_17259,N_10147,N_13838);
nand U17260 (N_17260,N_13500,N_11152);
or U17261 (N_17261,N_10518,N_10724);
and U17262 (N_17262,N_10877,N_12073);
or U17263 (N_17263,N_11561,N_11789);
nor U17264 (N_17264,N_11550,N_13811);
nand U17265 (N_17265,N_10330,N_14018);
nand U17266 (N_17266,N_12126,N_14207);
or U17267 (N_17267,N_10075,N_13774);
nor U17268 (N_17268,N_10800,N_11112);
and U17269 (N_17269,N_12935,N_11663);
or U17270 (N_17270,N_10082,N_12198);
or U17271 (N_17271,N_13580,N_12589);
nand U17272 (N_17272,N_14873,N_10674);
or U17273 (N_17273,N_11251,N_13234);
and U17274 (N_17274,N_12456,N_13047);
and U17275 (N_17275,N_14818,N_13232);
nand U17276 (N_17276,N_10143,N_10138);
or U17277 (N_17277,N_13441,N_14798);
nand U17278 (N_17278,N_13833,N_13548);
or U17279 (N_17279,N_11425,N_13137);
and U17280 (N_17280,N_14826,N_12381);
and U17281 (N_17281,N_14624,N_10957);
nand U17282 (N_17282,N_14490,N_10601);
nand U17283 (N_17283,N_14019,N_12859);
or U17284 (N_17284,N_14359,N_10959);
or U17285 (N_17285,N_13516,N_10046);
nor U17286 (N_17286,N_14327,N_13154);
and U17287 (N_17287,N_12815,N_13215);
nor U17288 (N_17288,N_11706,N_10806);
nand U17289 (N_17289,N_10238,N_14916);
nand U17290 (N_17290,N_14616,N_13978);
and U17291 (N_17291,N_13135,N_13722);
nand U17292 (N_17292,N_11241,N_12672);
nor U17293 (N_17293,N_14601,N_10289);
and U17294 (N_17294,N_11447,N_11328);
nor U17295 (N_17295,N_10535,N_10842);
and U17296 (N_17296,N_14867,N_12750);
and U17297 (N_17297,N_13084,N_12104);
and U17298 (N_17298,N_10436,N_11698);
nand U17299 (N_17299,N_12172,N_14480);
xor U17300 (N_17300,N_14888,N_11700);
or U17301 (N_17301,N_14274,N_13656);
nor U17302 (N_17302,N_12807,N_10364);
nand U17303 (N_17303,N_11395,N_10920);
or U17304 (N_17304,N_10224,N_12338);
or U17305 (N_17305,N_11945,N_12150);
and U17306 (N_17306,N_14025,N_11939);
or U17307 (N_17307,N_13479,N_10780);
nor U17308 (N_17308,N_13729,N_10107);
nor U17309 (N_17309,N_13376,N_10246);
and U17310 (N_17310,N_13832,N_11052);
and U17311 (N_17311,N_10457,N_12939);
nand U17312 (N_17312,N_10232,N_10134);
or U17313 (N_17313,N_10799,N_10482);
nand U17314 (N_17314,N_12756,N_12122);
and U17315 (N_17315,N_13738,N_11080);
and U17316 (N_17316,N_13060,N_13522);
or U17317 (N_17317,N_13923,N_14187);
nand U17318 (N_17318,N_12159,N_11541);
nor U17319 (N_17319,N_10586,N_12890);
nand U17320 (N_17320,N_14863,N_14402);
and U17321 (N_17321,N_13004,N_12964);
or U17322 (N_17322,N_14416,N_11226);
and U17323 (N_17323,N_13162,N_10652);
nor U17324 (N_17324,N_14092,N_10479);
nand U17325 (N_17325,N_11486,N_13420);
and U17326 (N_17326,N_12484,N_10785);
nand U17327 (N_17327,N_10905,N_14820);
nand U17328 (N_17328,N_14090,N_10974);
nand U17329 (N_17329,N_10085,N_10585);
nand U17330 (N_17330,N_13294,N_12477);
nand U17331 (N_17331,N_10590,N_14972);
nor U17332 (N_17332,N_12548,N_11320);
nor U17333 (N_17333,N_14558,N_13796);
nand U17334 (N_17334,N_13794,N_14871);
and U17335 (N_17335,N_11042,N_12021);
and U17336 (N_17336,N_13102,N_13995);
nor U17337 (N_17337,N_14896,N_13453);
nor U17338 (N_17338,N_10308,N_12248);
nor U17339 (N_17339,N_13409,N_14417);
nor U17340 (N_17340,N_14958,N_14816);
or U17341 (N_17341,N_11249,N_12415);
or U17342 (N_17342,N_11543,N_11987);
or U17343 (N_17343,N_10394,N_10100);
and U17344 (N_17344,N_12558,N_14806);
or U17345 (N_17345,N_10963,N_10176);
or U17346 (N_17346,N_14513,N_12015);
or U17347 (N_17347,N_13543,N_14012);
or U17348 (N_17348,N_11884,N_14979);
nand U17349 (N_17349,N_13966,N_11740);
or U17350 (N_17350,N_10663,N_10996);
or U17351 (N_17351,N_11305,N_13119);
nand U17352 (N_17352,N_14822,N_13411);
nor U17353 (N_17353,N_10970,N_13881);
and U17354 (N_17354,N_12518,N_14133);
or U17355 (N_17355,N_10237,N_11419);
xor U17356 (N_17356,N_12303,N_12895);
or U17357 (N_17357,N_10458,N_14131);
and U17358 (N_17358,N_13285,N_11573);
nand U17359 (N_17359,N_13475,N_13581);
and U17360 (N_17360,N_11292,N_13349);
nor U17361 (N_17361,N_11725,N_14562);
nand U17362 (N_17362,N_10426,N_12208);
nand U17363 (N_17363,N_11867,N_12100);
nand U17364 (N_17364,N_14383,N_14787);
or U17365 (N_17365,N_14291,N_11185);
or U17366 (N_17366,N_11692,N_14412);
or U17367 (N_17367,N_14279,N_14990);
or U17368 (N_17368,N_14307,N_11145);
or U17369 (N_17369,N_11344,N_11422);
or U17370 (N_17370,N_12252,N_11542);
and U17371 (N_17371,N_12051,N_14776);
nor U17372 (N_17372,N_12653,N_10827);
or U17373 (N_17373,N_10626,N_12535);
nor U17374 (N_17374,N_11433,N_10942);
nand U17375 (N_17375,N_11296,N_11694);
nor U17376 (N_17376,N_11964,N_12869);
and U17377 (N_17377,N_14507,N_10725);
or U17378 (N_17378,N_11623,N_12275);
or U17379 (N_17379,N_13206,N_14780);
or U17380 (N_17380,N_12992,N_11625);
or U17381 (N_17381,N_11040,N_11646);
and U17382 (N_17382,N_14844,N_14889);
or U17383 (N_17383,N_12978,N_10429);
nand U17384 (N_17384,N_12304,N_13043);
nand U17385 (N_17385,N_13822,N_11262);
nand U17386 (N_17386,N_11146,N_13460);
nor U17387 (N_17387,N_10336,N_10861);
and U17388 (N_17388,N_13214,N_13758);
nand U17389 (N_17389,N_10517,N_11428);
nand U17390 (N_17390,N_14167,N_12930);
nor U17391 (N_17391,N_14493,N_11842);
or U17392 (N_17392,N_13208,N_12799);
and U17393 (N_17393,N_12354,N_11720);
or U17394 (N_17394,N_13245,N_11315);
nand U17395 (N_17395,N_11367,N_14320);
nand U17396 (N_17396,N_10930,N_14148);
and U17397 (N_17397,N_12826,N_11284);
nand U17398 (N_17398,N_10410,N_14944);
nand U17399 (N_17399,N_14177,N_10168);
or U17400 (N_17400,N_10476,N_12595);
and U17401 (N_17401,N_10634,N_11065);
or U17402 (N_17402,N_13168,N_12601);
xnor U17403 (N_17403,N_10465,N_10672);
or U17404 (N_17404,N_14506,N_11730);
nor U17405 (N_17405,N_13613,N_11876);
or U17406 (N_17406,N_13947,N_14117);
and U17407 (N_17407,N_11847,N_12460);
and U17408 (N_17408,N_13158,N_11667);
nor U17409 (N_17409,N_14681,N_12539);
nor U17410 (N_17410,N_13106,N_11746);
or U17411 (N_17411,N_11579,N_14242);
nor U17412 (N_17412,N_14448,N_13072);
nor U17413 (N_17413,N_10031,N_11083);
or U17414 (N_17414,N_14535,N_13672);
nor U17415 (N_17415,N_14741,N_10670);
nand U17416 (N_17416,N_13956,N_12209);
nor U17417 (N_17417,N_12831,N_11378);
and U17418 (N_17418,N_12212,N_14637);
and U17419 (N_17419,N_12299,N_11868);
nand U17420 (N_17420,N_14671,N_10572);
nor U17421 (N_17421,N_12735,N_13766);
nor U17422 (N_17422,N_10337,N_12528);
nor U17423 (N_17423,N_12005,N_11849);
nand U17424 (N_17424,N_13884,N_14298);
and U17425 (N_17425,N_10766,N_13996);
nor U17426 (N_17426,N_13018,N_12834);
nor U17427 (N_17427,N_14502,N_12762);
and U17428 (N_17428,N_10606,N_13394);
nor U17429 (N_17429,N_14566,N_10428);
and U17430 (N_17430,N_10124,N_11599);
nor U17431 (N_17431,N_10125,N_10506);
nor U17432 (N_17432,N_13709,N_11982);
or U17433 (N_17433,N_10696,N_14960);
nand U17434 (N_17434,N_14643,N_11135);
nor U17435 (N_17435,N_11243,N_11697);
nand U17436 (N_17436,N_14060,N_12759);
nand U17437 (N_17437,N_10321,N_13798);
nor U17438 (N_17438,N_14465,N_12070);
nand U17439 (N_17439,N_12917,N_10753);
nand U17440 (N_17440,N_12722,N_14565);
nor U17441 (N_17441,N_13414,N_11584);
or U17442 (N_17442,N_14556,N_14107);
nor U17443 (N_17443,N_13114,N_10017);
nor U17444 (N_17444,N_11860,N_10359);
or U17445 (N_17445,N_13337,N_12970);
and U17446 (N_17446,N_11917,N_12013);
or U17447 (N_17447,N_10179,N_14856);
nand U17448 (N_17448,N_10967,N_12822);
and U17449 (N_17449,N_11708,N_13719);
and U17450 (N_17450,N_13197,N_13806);
or U17451 (N_17451,N_14994,N_12445);
xnor U17452 (N_17452,N_11003,N_12908);
and U17453 (N_17453,N_11101,N_12020);
or U17454 (N_17454,N_11404,N_11383);
and U17455 (N_17455,N_10531,N_11752);
nand U17456 (N_17456,N_13082,N_11199);
nand U17457 (N_17457,N_14394,N_10322);
and U17458 (N_17458,N_10511,N_11078);
or U17459 (N_17459,N_14072,N_12634);
and U17460 (N_17460,N_11759,N_12957);
and U17461 (N_17461,N_10836,N_14885);
nor U17462 (N_17462,N_13085,N_13848);
nand U17463 (N_17463,N_10127,N_14410);
or U17464 (N_17464,N_10835,N_13125);
nor U17465 (N_17465,N_14679,N_11373);
nor U17466 (N_17466,N_11281,N_12701);
nor U17467 (N_17467,N_10378,N_10551);
nand U17468 (N_17468,N_13430,N_10636);
nand U17469 (N_17469,N_10139,N_11056);
and U17470 (N_17470,N_11340,N_14149);
and U17471 (N_17471,N_14930,N_11017);
nor U17472 (N_17472,N_11918,N_12177);
nor U17473 (N_17473,N_12003,N_12603);
xnor U17474 (N_17474,N_12671,N_14695);
nand U17475 (N_17475,N_12726,N_14035);
nand U17476 (N_17476,N_13194,N_12494);
xnor U17477 (N_17477,N_10473,N_12313);
nor U17478 (N_17478,N_13635,N_10926);
and U17479 (N_17479,N_12689,N_12008);
nor U17480 (N_17480,N_12793,N_12586);
nand U17481 (N_17481,N_12316,N_10628);
xor U17482 (N_17482,N_12533,N_10922);
nor U17483 (N_17483,N_14709,N_10000);
or U17484 (N_17484,N_10263,N_10644);
or U17485 (N_17485,N_12179,N_12635);
or U17486 (N_17486,N_11456,N_14364);
nor U17487 (N_17487,N_11755,N_10528);
or U17488 (N_17488,N_12987,N_12521);
and U17489 (N_17489,N_13526,N_14628);
or U17490 (N_17490,N_11308,N_13846);
or U17491 (N_17491,N_11807,N_14861);
nand U17492 (N_17492,N_10894,N_14036);
nand U17493 (N_17493,N_13188,N_13030);
or U17494 (N_17494,N_14612,N_13968);
and U17495 (N_17495,N_11005,N_11115);
and U17496 (N_17496,N_12920,N_11084);
nand U17497 (N_17497,N_12850,N_14345);
and U17498 (N_17498,N_13007,N_11132);
or U17499 (N_17499,N_14277,N_14828);
and U17500 (N_17500,N_13537,N_11456);
or U17501 (N_17501,N_14339,N_10982);
nor U17502 (N_17502,N_10186,N_14670);
nor U17503 (N_17503,N_10743,N_10614);
and U17504 (N_17504,N_10334,N_12380);
or U17505 (N_17505,N_12456,N_10583);
nand U17506 (N_17506,N_14703,N_12099);
nor U17507 (N_17507,N_10539,N_11748);
and U17508 (N_17508,N_14797,N_14627);
nand U17509 (N_17509,N_12104,N_14676);
and U17510 (N_17510,N_13594,N_14917);
nand U17511 (N_17511,N_12461,N_14904);
or U17512 (N_17512,N_11183,N_12506);
or U17513 (N_17513,N_13893,N_14035);
nor U17514 (N_17514,N_11945,N_10671);
or U17515 (N_17515,N_14618,N_10159);
nand U17516 (N_17516,N_10033,N_14948);
nor U17517 (N_17517,N_12412,N_13957);
nand U17518 (N_17518,N_13928,N_14434);
nor U17519 (N_17519,N_12133,N_13268);
or U17520 (N_17520,N_12225,N_14041);
nor U17521 (N_17521,N_10336,N_12593);
nand U17522 (N_17522,N_11250,N_11456);
and U17523 (N_17523,N_13993,N_11187);
nand U17524 (N_17524,N_10151,N_10396);
nand U17525 (N_17525,N_10004,N_14758);
nor U17526 (N_17526,N_11781,N_13990);
and U17527 (N_17527,N_11988,N_12535);
nand U17528 (N_17528,N_11293,N_13283);
and U17529 (N_17529,N_10505,N_12457);
nor U17530 (N_17530,N_14496,N_13181);
or U17531 (N_17531,N_13370,N_10018);
nor U17532 (N_17532,N_11123,N_12687);
nor U17533 (N_17533,N_11096,N_10514);
nand U17534 (N_17534,N_12606,N_13082);
or U17535 (N_17535,N_14574,N_14712);
or U17536 (N_17536,N_10382,N_14413);
nor U17537 (N_17537,N_11253,N_12205);
and U17538 (N_17538,N_10037,N_12382);
xor U17539 (N_17539,N_14946,N_13915);
nand U17540 (N_17540,N_14435,N_10989);
nor U17541 (N_17541,N_11865,N_12759);
and U17542 (N_17542,N_13967,N_12417);
or U17543 (N_17543,N_13824,N_12672);
or U17544 (N_17544,N_10440,N_12854);
or U17545 (N_17545,N_12197,N_12093);
nand U17546 (N_17546,N_13622,N_11732);
or U17547 (N_17547,N_11428,N_10360);
nor U17548 (N_17548,N_12895,N_13271);
or U17549 (N_17549,N_11742,N_11834);
nand U17550 (N_17550,N_14927,N_13271);
nor U17551 (N_17551,N_11500,N_13098);
or U17552 (N_17552,N_10590,N_11675);
nor U17553 (N_17553,N_13709,N_10650);
nand U17554 (N_17554,N_12680,N_12147);
and U17555 (N_17555,N_13950,N_10520);
or U17556 (N_17556,N_14024,N_13512);
nand U17557 (N_17557,N_11314,N_14225);
nand U17558 (N_17558,N_14898,N_13086);
nand U17559 (N_17559,N_13570,N_12959);
nand U17560 (N_17560,N_12198,N_10889);
and U17561 (N_17561,N_10831,N_12373);
or U17562 (N_17562,N_14544,N_12369);
nand U17563 (N_17563,N_11172,N_14145);
nor U17564 (N_17564,N_13044,N_14987);
nor U17565 (N_17565,N_12828,N_14796);
nand U17566 (N_17566,N_13232,N_11484);
or U17567 (N_17567,N_10320,N_12116);
or U17568 (N_17568,N_14810,N_11369);
or U17569 (N_17569,N_14684,N_11501);
or U17570 (N_17570,N_12336,N_14782);
or U17571 (N_17571,N_12475,N_12403);
and U17572 (N_17572,N_12928,N_10525);
or U17573 (N_17573,N_12583,N_13348);
and U17574 (N_17574,N_10657,N_12319);
or U17575 (N_17575,N_11665,N_13628);
or U17576 (N_17576,N_13622,N_11297);
or U17577 (N_17577,N_12311,N_11606);
nor U17578 (N_17578,N_13881,N_14202);
nand U17579 (N_17579,N_12998,N_10129);
nor U17580 (N_17580,N_14334,N_13516);
and U17581 (N_17581,N_12894,N_12178);
nor U17582 (N_17582,N_12790,N_10318);
nor U17583 (N_17583,N_11605,N_12772);
or U17584 (N_17584,N_10206,N_13927);
or U17585 (N_17585,N_14151,N_11167);
nand U17586 (N_17586,N_13191,N_11058);
and U17587 (N_17587,N_12940,N_13648);
or U17588 (N_17588,N_14333,N_14989);
xnor U17589 (N_17589,N_14679,N_11510);
nand U17590 (N_17590,N_11604,N_12117);
nand U17591 (N_17591,N_12443,N_10591);
nor U17592 (N_17592,N_12325,N_12402);
nor U17593 (N_17593,N_14157,N_12849);
nand U17594 (N_17594,N_12180,N_10974);
and U17595 (N_17595,N_14480,N_11186);
nor U17596 (N_17596,N_14428,N_10107);
nand U17597 (N_17597,N_10508,N_11995);
nand U17598 (N_17598,N_11521,N_10961);
and U17599 (N_17599,N_14921,N_10854);
nand U17600 (N_17600,N_12414,N_11480);
and U17601 (N_17601,N_12783,N_12029);
or U17602 (N_17602,N_14929,N_11929);
nand U17603 (N_17603,N_14893,N_12642);
and U17604 (N_17604,N_14751,N_10003);
and U17605 (N_17605,N_11991,N_14179);
nand U17606 (N_17606,N_14616,N_10452);
nor U17607 (N_17607,N_11993,N_13493);
nor U17608 (N_17608,N_10306,N_14963);
or U17609 (N_17609,N_11477,N_11536);
and U17610 (N_17610,N_10357,N_14026);
or U17611 (N_17611,N_13027,N_10829);
nand U17612 (N_17612,N_11973,N_14318);
or U17613 (N_17613,N_10456,N_11913);
and U17614 (N_17614,N_11370,N_11771);
and U17615 (N_17615,N_14583,N_11102);
and U17616 (N_17616,N_14998,N_12329);
nand U17617 (N_17617,N_14500,N_14358);
nand U17618 (N_17618,N_13752,N_10363);
nand U17619 (N_17619,N_10465,N_12081);
or U17620 (N_17620,N_12187,N_14386);
or U17621 (N_17621,N_12014,N_10888);
nor U17622 (N_17622,N_11921,N_10042);
nand U17623 (N_17623,N_10741,N_12100);
and U17624 (N_17624,N_12910,N_10841);
or U17625 (N_17625,N_14071,N_12712);
nand U17626 (N_17626,N_14050,N_14099);
nand U17627 (N_17627,N_10566,N_10713);
and U17628 (N_17628,N_12439,N_13458);
nor U17629 (N_17629,N_10436,N_11061);
nor U17630 (N_17630,N_10488,N_11581);
or U17631 (N_17631,N_14350,N_13019);
and U17632 (N_17632,N_10657,N_13555);
or U17633 (N_17633,N_12868,N_13754);
nor U17634 (N_17634,N_10477,N_12762);
nor U17635 (N_17635,N_14407,N_10034);
nor U17636 (N_17636,N_13310,N_14491);
or U17637 (N_17637,N_12174,N_11295);
nor U17638 (N_17638,N_12363,N_11387);
and U17639 (N_17639,N_13862,N_14088);
and U17640 (N_17640,N_13091,N_11965);
or U17641 (N_17641,N_10078,N_10215);
and U17642 (N_17642,N_10156,N_14518);
or U17643 (N_17643,N_12618,N_14795);
and U17644 (N_17644,N_12603,N_11518);
nand U17645 (N_17645,N_12986,N_10383);
nor U17646 (N_17646,N_10898,N_12733);
nand U17647 (N_17647,N_12498,N_10925);
or U17648 (N_17648,N_11027,N_11367);
xor U17649 (N_17649,N_11034,N_14604);
and U17650 (N_17650,N_14551,N_10677);
xnor U17651 (N_17651,N_13827,N_11581);
nand U17652 (N_17652,N_14610,N_11598);
nor U17653 (N_17653,N_13542,N_12006);
and U17654 (N_17654,N_12874,N_14176);
or U17655 (N_17655,N_13052,N_12604);
nand U17656 (N_17656,N_13333,N_12542);
nor U17657 (N_17657,N_13902,N_11930);
and U17658 (N_17658,N_10066,N_14105);
nor U17659 (N_17659,N_13559,N_10827);
nand U17660 (N_17660,N_12899,N_10179);
nor U17661 (N_17661,N_13655,N_12872);
or U17662 (N_17662,N_10505,N_10495);
and U17663 (N_17663,N_10936,N_14334);
or U17664 (N_17664,N_10831,N_13417);
nor U17665 (N_17665,N_10458,N_13177);
and U17666 (N_17666,N_10996,N_11418);
or U17667 (N_17667,N_10319,N_10976);
and U17668 (N_17668,N_10023,N_10842);
nor U17669 (N_17669,N_10607,N_11985);
nand U17670 (N_17670,N_14595,N_11987);
and U17671 (N_17671,N_14326,N_14437);
nand U17672 (N_17672,N_10009,N_10572);
or U17673 (N_17673,N_12558,N_12660);
nor U17674 (N_17674,N_14399,N_12200);
nand U17675 (N_17675,N_14011,N_12210);
and U17676 (N_17676,N_13526,N_11674);
or U17677 (N_17677,N_12903,N_13874);
or U17678 (N_17678,N_10594,N_14423);
nor U17679 (N_17679,N_10455,N_13739);
or U17680 (N_17680,N_13352,N_12289);
or U17681 (N_17681,N_14004,N_12261);
and U17682 (N_17682,N_10117,N_14518);
and U17683 (N_17683,N_14899,N_14529);
or U17684 (N_17684,N_12836,N_10183);
or U17685 (N_17685,N_14299,N_12069);
and U17686 (N_17686,N_13923,N_12627);
and U17687 (N_17687,N_13070,N_14593);
and U17688 (N_17688,N_10288,N_10949);
or U17689 (N_17689,N_10417,N_11777);
nor U17690 (N_17690,N_12724,N_13989);
and U17691 (N_17691,N_11135,N_13346);
or U17692 (N_17692,N_10930,N_12209);
or U17693 (N_17693,N_14656,N_10760);
or U17694 (N_17694,N_10722,N_12531);
or U17695 (N_17695,N_14156,N_10407);
nand U17696 (N_17696,N_14015,N_11595);
nand U17697 (N_17697,N_14094,N_11561);
nand U17698 (N_17698,N_11136,N_10311);
and U17699 (N_17699,N_14112,N_10952);
nor U17700 (N_17700,N_10437,N_11472);
or U17701 (N_17701,N_13484,N_14628);
nand U17702 (N_17702,N_10822,N_13876);
and U17703 (N_17703,N_12069,N_10196);
nor U17704 (N_17704,N_10359,N_14628);
or U17705 (N_17705,N_11456,N_12737);
nor U17706 (N_17706,N_10281,N_11507);
and U17707 (N_17707,N_12971,N_13695);
nor U17708 (N_17708,N_14044,N_14122);
nand U17709 (N_17709,N_12718,N_11591);
or U17710 (N_17710,N_12407,N_14495);
and U17711 (N_17711,N_13989,N_13568);
or U17712 (N_17712,N_13248,N_14849);
nor U17713 (N_17713,N_12110,N_13664);
or U17714 (N_17714,N_11128,N_12721);
nor U17715 (N_17715,N_11286,N_11986);
or U17716 (N_17716,N_10962,N_11468);
or U17717 (N_17717,N_14630,N_14980);
and U17718 (N_17718,N_13161,N_13831);
or U17719 (N_17719,N_10676,N_11165);
or U17720 (N_17720,N_10362,N_12028);
or U17721 (N_17721,N_12085,N_13001);
or U17722 (N_17722,N_11296,N_11023);
xor U17723 (N_17723,N_13368,N_12722);
nand U17724 (N_17724,N_13455,N_13786);
nor U17725 (N_17725,N_13004,N_11071);
nand U17726 (N_17726,N_11492,N_14141);
xor U17727 (N_17727,N_13375,N_11366);
nor U17728 (N_17728,N_11196,N_10845);
and U17729 (N_17729,N_11345,N_13863);
nand U17730 (N_17730,N_10090,N_13791);
and U17731 (N_17731,N_10675,N_13645);
or U17732 (N_17732,N_13015,N_13729);
and U17733 (N_17733,N_10198,N_14695);
or U17734 (N_17734,N_14764,N_10198);
and U17735 (N_17735,N_14612,N_13766);
or U17736 (N_17736,N_13927,N_12179);
nor U17737 (N_17737,N_11652,N_14605);
and U17738 (N_17738,N_11884,N_11719);
nand U17739 (N_17739,N_14437,N_14581);
nand U17740 (N_17740,N_11772,N_12447);
nor U17741 (N_17741,N_10252,N_11663);
and U17742 (N_17742,N_12718,N_14017);
and U17743 (N_17743,N_12503,N_14490);
or U17744 (N_17744,N_12167,N_14319);
xor U17745 (N_17745,N_10396,N_10139);
or U17746 (N_17746,N_11281,N_14577);
nor U17747 (N_17747,N_11474,N_13190);
or U17748 (N_17748,N_11897,N_14027);
and U17749 (N_17749,N_10448,N_11687);
nor U17750 (N_17750,N_12865,N_10000);
nand U17751 (N_17751,N_14527,N_10216);
or U17752 (N_17752,N_12480,N_14711);
nor U17753 (N_17753,N_12705,N_13885);
and U17754 (N_17754,N_10457,N_14675);
or U17755 (N_17755,N_14351,N_10169);
or U17756 (N_17756,N_13285,N_13713);
nand U17757 (N_17757,N_10722,N_10008);
nand U17758 (N_17758,N_13497,N_14125);
or U17759 (N_17759,N_10042,N_13146);
nand U17760 (N_17760,N_14245,N_10972);
or U17761 (N_17761,N_10231,N_11683);
nor U17762 (N_17762,N_12314,N_14738);
and U17763 (N_17763,N_11404,N_11876);
nand U17764 (N_17764,N_13623,N_11754);
nor U17765 (N_17765,N_10482,N_12972);
nor U17766 (N_17766,N_11067,N_14901);
or U17767 (N_17767,N_14100,N_10608);
nand U17768 (N_17768,N_10108,N_12017);
and U17769 (N_17769,N_11175,N_10907);
or U17770 (N_17770,N_10160,N_12496);
or U17771 (N_17771,N_13238,N_10043);
or U17772 (N_17772,N_10287,N_12687);
nor U17773 (N_17773,N_14411,N_13729);
xor U17774 (N_17774,N_14888,N_10210);
or U17775 (N_17775,N_12466,N_11196);
nand U17776 (N_17776,N_11159,N_14971);
or U17777 (N_17777,N_10427,N_10570);
or U17778 (N_17778,N_12589,N_13801);
or U17779 (N_17779,N_12945,N_10610);
or U17780 (N_17780,N_11449,N_12054);
or U17781 (N_17781,N_13756,N_12695);
and U17782 (N_17782,N_14497,N_10655);
nand U17783 (N_17783,N_13774,N_14512);
nand U17784 (N_17784,N_10166,N_10920);
nor U17785 (N_17785,N_12595,N_12395);
nor U17786 (N_17786,N_14174,N_14683);
or U17787 (N_17787,N_13128,N_10453);
nor U17788 (N_17788,N_13482,N_13431);
and U17789 (N_17789,N_14350,N_14043);
nand U17790 (N_17790,N_11129,N_11437);
or U17791 (N_17791,N_14366,N_14396);
or U17792 (N_17792,N_11614,N_13217);
nor U17793 (N_17793,N_14792,N_13613);
and U17794 (N_17794,N_10724,N_11335);
nor U17795 (N_17795,N_14158,N_14781);
nor U17796 (N_17796,N_12780,N_10576);
or U17797 (N_17797,N_10637,N_14171);
nor U17798 (N_17798,N_14364,N_10852);
and U17799 (N_17799,N_14737,N_10410);
xor U17800 (N_17800,N_11143,N_10770);
nand U17801 (N_17801,N_14240,N_14586);
nor U17802 (N_17802,N_10597,N_13476);
or U17803 (N_17803,N_12652,N_13470);
and U17804 (N_17804,N_13194,N_11006);
or U17805 (N_17805,N_12854,N_11057);
or U17806 (N_17806,N_14444,N_10097);
nor U17807 (N_17807,N_10826,N_11441);
nand U17808 (N_17808,N_11478,N_14704);
and U17809 (N_17809,N_14129,N_14138);
xor U17810 (N_17810,N_14230,N_14715);
nor U17811 (N_17811,N_10169,N_12697);
and U17812 (N_17812,N_11930,N_11984);
and U17813 (N_17813,N_13396,N_12678);
nand U17814 (N_17814,N_13159,N_13323);
and U17815 (N_17815,N_14021,N_12704);
nand U17816 (N_17816,N_11680,N_12673);
nand U17817 (N_17817,N_11726,N_10667);
or U17818 (N_17818,N_11605,N_12654);
or U17819 (N_17819,N_11434,N_13858);
and U17820 (N_17820,N_11806,N_14116);
nor U17821 (N_17821,N_11874,N_14302);
and U17822 (N_17822,N_11476,N_12599);
nor U17823 (N_17823,N_13939,N_13870);
or U17824 (N_17824,N_12015,N_13757);
nand U17825 (N_17825,N_13187,N_11025);
and U17826 (N_17826,N_11324,N_13434);
nor U17827 (N_17827,N_10261,N_10926);
and U17828 (N_17828,N_12582,N_10209);
and U17829 (N_17829,N_14383,N_12680);
or U17830 (N_17830,N_13788,N_11938);
and U17831 (N_17831,N_10512,N_12243);
and U17832 (N_17832,N_10510,N_11935);
nor U17833 (N_17833,N_13153,N_10134);
or U17834 (N_17834,N_13946,N_10848);
nor U17835 (N_17835,N_11552,N_14168);
nand U17836 (N_17836,N_14643,N_12210);
and U17837 (N_17837,N_14296,N_10942);
nand U17838 (N_17838,N_10875,N_13500);
nand U17839 (N_17839,N_14672,N_14384);
or U17840 (N_17840,N_13768,N_11829);
nor U17841 (N_17841,N_10214,N_10571);
nor U17842 (N_17842,N_14439,N_14349);
and U17843 (N_17843,N_13618,N_10045);
and U17844 (N_17844,N_12092,N_13409);
nand U17845 (N_17845,N_12648,N_11422);
nand U17846 (N_17846,N_12657,N_12022);
and U17847 (N_17847,N_11635,N_13449);
and U17848 (N_17848,N_10737,N_10655);
nor U17849 (N_17849,N_14207,N_14072);
nand U17850 (N_17850,N_14465,N_14514);
nor U17851 (N_17851,N_13255,N_11252);
or U17852 (N_17852,N_12992,N_14872);
nand U17853 (N_17853,N_11629,N_11621);
nand U17854 (N_17854,N_12259,N_14527);
nand U17855 (N_17855,N_12141,N_10332);
or U17856 (N_17856,N_12670,N_11688);
nand U17857 (N_17857,N_13754,N_14569);
or U17858 (N_17858,N_12922,N_13573);
and U17859 (N_17859,N_12738,N_11817);
and U17860 (N_17860,N_12992,N_14250);
and U17861 (N_17861,N_11290,N_14725);
nand U17862 (N_17862,N_11128,N_10207);
nor U17863 (N_17863,N_11503,N_12523);
nand U17864 (N_17864,N_13705,N_13105);
nor U17865 (N_17865,N_12463,N_14855);
nor U17866 (N_17866,N_13196,N_13419);
nor U17867 (N_17867,N_12710,N_14434);
nor U17868 (N_17868,N_14463,N_10540);
or U17869 (N_17869,N_12567,N_14123);
or U17870 (N_17870,N_14508,N_13106);
nand U17871 (N_17871,N_11894,N_14450);
nor U17872 (N_17872,N_12575,N_12989);
nand U17873 (N_17873,N_14512,N_12640);
and U17874 (N_17874,N_12521,N_14846);
and U17875 (N_17875,N_10540,N_12386);
nand U17876 (N_17876,N_14979,N_11845);
nand U17877 (N_17877,N_13735,N_14300);
nand U17878 (N_17878,N_11232,N_13112);
nand U17879 (N_17879,N_13116,N_11746);
xor U17880 (N_17880,N_14359,N_12816);
or U17881 (N_17881,N_11573,N_10604);
or U17882 (N_17882,N_10239,N_13892);
nand U17883 (N_17883,N_14750,N_10330);
nand U17884 (N_17884,N_14918,N_11225);
or U17885 (N_17885,N_12830,N_11298);
and U17886 (N_17886,N_13869,N_10960);
xor U17887 (N_17887,N_13649,N_13290);
nand U17888 (N_17888,N_12594,N_12253);
nand U17889 (N_17889,N_12760,N_10121);
or U17890 (N_17890,N_14767,N_14030);
and U17891 (N_17891,N_14785,N_11354);
or U17892 (N_17892,N_11457,N_12676);
or U17893 (N_17893,N_11441,N_14690);
nand U17894 (N_17894,N_11464,N_11283);
nor U17895 (N_17895,N_10168,N_14988);
nand U17896 (N_17896,N_12764,N_13747);
nand U17897 (N_17897,N_10866,N_12932);
or U17898 (N_17898,N_14377,N_13784);
and U17899 (N_17899,N_11481,N_10819);
nor U17900 (N_17900,N_10255,N_12533);
nor U17901 (N_17901,N_13309,N_12901);
xnor U17902 (N_17902,N_11484,N_12681);
nand U17903 (N_17903,N_11548,N_14091);
and U17904 (N_17904,N_11826,N_13709);
nand U17905 (N_17905,N_14028,N_13486);
or U17906 (N_17906,N_11373,N_11355);
or U17907 (N_17907,N_12811,N_13930);
or U17908 (N_17908,N_10248,N_12646);
nand U17909 (N_17909,N_14715,N_14114);
nor U17910 (N_17910,N_14856,N_10211);
xor U17911 (N_17911,N_11846,N_11694);
or U17912 (N_17912,N_12196,N_11914);
and U17913 (N_17913,N_11988,N_11665);
nand U17914 (N_17914,N_14683,N_10607);
nor U17915 (N_17915,N_13379,N_11248);
and U17916 (N_17916,N_14196,N_13161);
or U17917 (N_17917,N_12324,N_10494);
nand U17918 (N_17918,N_14485,N_12058);
nor U17919 (N_17919,N_14437,N_10216);
nand U17920 (N_17920,N_14988,N_10184);
nor U17921 (N_17921,N_10929,N_12008);
or U17922 (N_17922,N_10130,N_12163);
nor U17923 (N_17923,N_14833,N_11115);
nand U17924 (N_17924,N_11859,N_12396);
nor U17925 (N_17925,N_10189,N_13444);
nand U17926 (N_17926,N_12038,N_14613);
or U17927 (N_17927,N_11887,N_12613);
nand U17928 (N_17928,N_14032,N_10584);
or U17929 (N_17929,N_10014,N_14023);
and U17930 (N_17930,N_13908,N_14278);
and U17931 (N_17931,N_11301,N_11184);
nor U17932 (N_17932,N_10537,N_10339);
or U17933 (N_17933,N_10216,N_12922);
and U17934 (N_17934,N_12140,N_11020);
nand U17935 (N_17935,N_11634,N_10425);
and U17936 (N_17936,N_10915,N_11712);
nor U17937 (N_17937,N_10545,N_14173);
nor U17938 (N_17938,N_14312,N_13366);
or U17939 (N_17939,N_11245,N_14323);
nor U17940 (N_17940,N_11487,N_13833);
nand U17941 (N_17941,N_12580,N_11448);
nor U17942 (N_17942,N_10807,N_12788);
and U17943 (N_17943,N_12595,N_10401);
nor U17944 (N_17944,N_10582,N_11597);
or U17945 (N_17945,N_14353,N_11608);
or U17946 (N_17946,N_10715,N_10967);
nand U17947 (N_17947,N_12084,N_10074);
nor U17948 (N_17948,N_13181,N_14748);
nor U17949 (N_17949,N_11436,N_14312);
and U17950 (N_17950,N_14799,N_10592);
nor U17951 (N_17951,N_10055,N_14034);
or U17952 (N_17952,N_13700,N_13908);
nand U17953 (N_17953,N_11945,N_10533);
and U17954 (N_17954,N_11223,N_10558);
nand U17955 (N_17955,N_11533,N_10735);
and U17956 (N_17956,N_14520,N_13802);
and U17957 (N_17957,N_11889,N_11628);
or U17958 (N_17958,N_11697,N_13515);
and U17959 (N_17959,N_12650,N_10815);
and U17960 (N_17960,N_14965,N_13021);
nand U17961 (N_17961,N_13714,N_11904);
nand U17962 (N_17962,N_14879,N_14317);
and U17963 (N_17963,N_14759,N_13243);
or U17964 (N_17964,N_13661,N_12649);
and U17965 (N_17965,N_11230,N_12735);
and U17966 (N_17966,N_11565,N_12576);
and U17967 (N_17967,N_14032,N_13246);
nand U17968 (N_17968,N_12859,N_12335);
nand U17969 (N_17969,N_14831,N_12827);
and U17970 (N_17970,N_14706,N_11977);
nand U17971 (N_17971,N_13818,N_11274);
nand U17972 (N_17972,N_13309,N_11578);
or U17973 (N_17973,N_11751,N_14812);
nor U17974 (N_17974,N_11840,N_11462);
and U17975 (N_17975,N_10557,N_14342);
and U17976 (N_17976,N_10042,N_11585);
nor U17977 (N_17977,N_13058,N_14678);
nor U17978 (N_17978,N_13045,N_14691);
and U17979 (N_17979,N_12811,N_10432);
or U17980 (N_17980,N_11690,N_12117);
nor U17981 (N_17981,N_14868,N_12250);
nor U17982 (N_17982,N_13450,N_11642);
nand U17983 (N_17983,N_12308,N_14246);
nor U17984 (N_17984,N_14384,N_13605);
or U17985 (N_17985,N_11982,N_11005);
and U17986 (N_17986,N_13875,N_14228);
nor U17987 (N_17987,N_10462,N_14490);
nand U17988 (N_17988,N_11571,N_13043);
or U17989 (N_17989,N_12584,N_13848);
nand U17990 (N_17990,N_12337,N_12255);
or U17991 (N_17991,N_14297,N_10231);
nand U17992 (N_17992,N_12096,N_14105);
nor U17993 (N_17993,N_14374,N_13828);
nor U17994 (N_17994,N_14871,N_14679);
or U17995 (N_17995,N_14193,N_12221);
and U17996 (N_17996,N_11422,N_10673);
and U17997 (N_17997,N_14641,N_11004);
or U17998 (N_17998,N_12474,N_13988);
or U17999 (N_17999,N_10132,N_14174);
and U18000 (N_18000,N_11113,N_11326);
and U18001 (N_18001,N_13639,N_13372);
nand U18002 (N_18002,N_14924,N_13931);
nand U18003 (N_18003,N_14825,N_12640);
xnor U18004 (N_18004,N_10903,N_12006);
nor U18005 (N_18005,N_10779,N_12625);
nor U18006 (N_18006,N_14164,N_14625);
or U18007 (N_18007,N_14567,N_13863);
nor U18008 (N_18008,N_13618,N_11168);
or U18009 (N_18009,N_14954,N_10740);
or U18010 (N_18010,N_12852,N_12911);
and U18011 (N_18011,N_11273,N_13515);
nor U18012 (N_18012,N_10342,N_10101);
nand U18013 (N_18013,N_12922,N_11726);
nand U18014 (N_18014,N_13625,N_11966);
or U18015 (N_18015,N_10844,N_14633);
or U18016 (N_18016,N_10170,N_10823);
and U18017 (N_18017,N_14998,N_14797);
nor U18018 (N_18018,N_13657,N_12349);
nor U18019 (N_18019,N_12273,N_11634);
nand U18020 (N_18020,N_13419,N_12156);
or U18021 (N_18021,N_11028,N_10537);
nor U18022 (N_18022,N_10791,N_10778);
and U18023 (N_18023,N_10295,N_12480);
nor U18024 (N_18024,N_10757,N_14871);
or U18025 (N_18025,N_10749,N_10095);
nor U18026 (N_18026,N_12263,N_11612);
xnor U18027 (N_18027,N_12346,N_11102);
nand U18028 (N_18028,N_10028,N_12106);
nand U18029 (N_18029,N_12190,N_10916);
and U18030 (N_18030,N_14182,N_12027);
or U18031 (N_18031,N_12423,N_12714);
or U18032 (N_18032,N_14059,N_13949);
nor U18033 (N_18033,N_14072,N_14071);
nor U18034 (N_18034,N_10528,N_13793);
or U18035 (N_18035,N_13081,N_10329);
xnor U18036 (N_18036,N_14970,N_14975);
nor U18037 (N_18037,N_12601,N_14369);
nand U18038 (N_18038,N_14566,N_11804);
or U18039 (N_18039,N_13601,N_14489);
and U18040 (N_18040,N_11860,N_12103);
nand U18041 (N_18041,N_14905,N_12084);
or U18042 (N_18042,N_14919,N_13674);
or U18043 (N_18043,N_11469,N_12242);
nand U18044 (N_18044,N_14155,N_13887);
nand U18045 (N_18045,N_14453,N_11567);
nand U18046 (N_18046,N_12287,N_10342);
nor U18047 (N_18047,N_12877,N_10936);
or U18048 (N_18048,N_14271,N_10802);
and U18049 (N_18049,N_10281,N_11021);
and U18050 (N_18050,N_14513,N_13832);
nand U18051 (N_18051,N_14469,N_12802);
nor U18052 (N_18052,N_13687,N_12793);
and U18053 (N_18053,N_14877,N_12060);
or U18054 (N_18054,N_12084,N_10333);
nor U18055 (N_18055,N_12273,N_13243);
nor U18056 (N_18056,N_13853,N_10541);
nor U18057 (N_18057,N_14619,N_11604);
nand U18058 (N_18058,N_13197,N_11308);
and U18059 (N_18059,N_10997,N_13865);
and U18060 (N_18060,N_14948,N_13643);
nand U18061 (N_18061,N_11015,N_11968);
and U18062 (N_18062,N_14816,N_14115);
and U18063 (N_18063,N_13470,N_14764);
or U18064 (N_18064,N_13665,N_14048);
nand U18065 (N_18065,N_14046,N_10696);
nand U18066 (N_18066,N_14012,N_11036);
and U18067 (N_18067,N_10949,N_14724);
nor U18068 (N_18068,N_13529,N_11784);
nor U18069 (N_18069,N_13114,N_12767);
nand U18070 (N_18070,N_14508,N_10416);
and U18071 (N_18071,N_11694,N_12874);
nor U18072 (N_18072,N_14319,N_12841);
and U18073 (N_18073,N_14766,N_13380);
nor U18074 (N_18074,N_10978,N_12974);
or U18075 (N_18075,N_13395,N_12422);
nor U18076 (N_18076,N_14601,N_12105);
and U18077 (N_18077,N_12241,N_14988);
nor U18078 (N_18078,N_10777,N_14738);
or U18079 (N_18079,N_12833,N_12226);
nor U18080 (N_18080,N_12808,N_12095);
and U18081 (N_18081,N_12237,N_14322);
or U18082 (N_18082,N_13876,N_12849);
or U18083 (N_18083,N_12171,N_12479);
nor U18084 (N_18084,N_12096,N_11980);
xnor U18085 (N_18085,N_12453,N_10708);
and U18086 (N_18086,N_10481,N_10605);
nor U18087 (N_18087,N_12141,N_11413);
and U18088 (N_18088,N_12295,N_10554);
and U18089 (N_18089,N_13885,N_13216);
nand U18090 (N_18090,N_11965,N_14822);
nor U18091 (N_18091,N_14317,N_10155);
xor U18092 (N_18092,N_10630,N_13120);
or U18093 (N_18093,N_12423,N_13682);
nand U18094 (N_18094,N_12512,N_10517);
nand U18095 (N_18095,N_10219,N_11678);
and U18096 (N_18096,N_10054,N_11493);
nand U18097 (N_18097,N_10854,N_14609);
xnor U18098 (N_18098,N_10451,N_12908);
nand U18099 (N_18099,N_10054,N_13510);
nor U18100 (N_18100,N_13859,N_13706);
and U18101 (N_18101,N_12499,N_14522);
nand U18102 (N_18102,N_13920,N_12456);
nor U18103 (N_18103,N_11148,N_12705);
or U18104 (N_18104,N_13139,N_12672);
and U18105 (N_18105,N_10171,N_10926);
nor U18106 (N_18106,N_12282,N_10958);
nand U18107 (N_18107,N_12927,N_14191);
or U18108 (N_18108,N_10607,N_10981);
or U18109 (N_18109,N_13940,N_14230);
and U18110 (N_18110,N_12552,N_11089);
and U18111 (N_18111,N_11303,N_12895);
or U18112 (N_18112,N_11819,N_11274);
or U18113 (N_18113,N_13082,N_13027);
nand U18114 (N_18114,N_13938,N_12545);
and U18115 (N_18115,N_13894,N_12656);
or U18116 (N_18116,N_14170,N_11430);
or U18117 (N_18117,N_12907,N_14286);
or U18118 (N_18118,N_13790,N_10203);
or U18119 (N_18119,N_14126,N_14770);
nor U18120 (N_18120,N_12751,N_13920);
and U18121 (N_18121,N_12780,N_12693);
nand U18122 (N_18122,N_11832,N_12483);
and U18123 (N_18123,N_12512,N_10052);
nand U18124 (N_18124,N_13956,N_10666);
or U18125 (N_18125,N_13819,N_11911);
nor U18126 (N_18126,N_10400,N_14434);
or U18127 (N_18127,N_12857,N_13653);
nand U18128 (N_18128,N_14352,N_11141);
nor U18129 (N_18129,N_12724,N_10698);
nor U18130 (N_18130,N_10879,N_14036);
nand U18131 (N_18131,N_13259,N_12648);
nor U18132 (N_18132,N_10107,N_10914);
and U18133 (N_18133,N_13111,N_14085);
nand U18134 (N_18134,N_12328,N_11542);
and U18135 (N_18135,N_14074,N_11466);
nor U18136 (N_18136,N_14864,N_12505);
or U18137 (N_18137,N_13842,N_13967);
nor U18138 (N_18138,N_14369,N_12699);
and U18139 (N_18139,N_10549,N_11580);
nand U18140 (N_18140,N_10016,N_10562);
and U18141 (N_18141,N_14383,N_13494);
nand U18142 (N_18142,N_13214,N_12217);
nand U18143 (N_18143,N_10533,N_11505);
or U18144 (N_18144,N_13078,N_12790);
nor U18145 (N_18145,N_13275,N_12292);
or U18146 (N_18146,N_14660,N_11237);
or U18147 (N_18147,N_11235,N_14657);
and U18148 (N_18148,N_12903,N_12764);
and U18149 (N_18149,N_14462,N_12662);
nand U18150 (N_18150,N_11031,N_11229);
nor U18151 (N_18151,N_14954,N_10035);
nor U18152 (N_18152,N_13454,N_12715);
nand U18153 (N_18153,N_12101,N_14475);
nor U18154 (N_18154,N_10050,N_14369);
and U18155 (N_18155,N_14882,N_11822);
or U18156 (N_18156,N_12689,N_11918);
nor U18157 (N_18157,N_14760,N_14892);
nand U18158 (N_18158,N_11386,N_13752);
nand U18159 (N_18159,N_13626,N_12299);
or U18160 (N_18160,N_12897,N_12070);
and U18161 (N_18161,N_13354,N_13160);
or U18162 (N_18162,N_13973,N_10609);
nand U18163 (N_18163,N_14081,N_14794);
and U18164 (N_18164,N_12115,N_13582);
nor U18165 (N_18165,N_10914,N_13090);
xnor U18166 (N_18166,N_11771,N_12417);
and U18167 (N_18167,N_11581,N_13516);
nor U18168 (N_18168,N_14727,N_11038);
nor U18169 (N_18169,N_10954,N_11548);
and U18170 (N_18170,N_14212,N_10185);
nand U18171 (N_18171,N_11066,N_14767);
and U18172 (N_18172,N_11768,N_14714);
nand U18173 (N_18173,N_13246,N_10981);
nor U18174 (N_18174,N_11934,N_11793);
nand U18175 (N_18175,N_14316,N_10672);
nor U18176 (N_18176,N_12282,N_11257);
nand U18177 (N_18177,N_14279,N_10858);
nor U18178 (N_18178,N_14392,N_14252);
and U18179 (N_18179,N_12503,N_10541);
and U18180 (N_18180,N_13751,N_13709);
and U18181 (N_18181,N_10640,N_14222);
nand U18182 (N_18182,N_14276,N_13746);
nand U18183 (N_18183,N_14866,N_13541);
nor U18184 (N_18184,N_10549,N_14652);
and U18185 (N_18185,N_10201,N_13517);
nor U18186 (N_18186,N_11427,N_11337);
nor U18187 (N_18187,N_11971,N_10605);
nor U18188 (N_18188,N_12810,N_14430);
nor U18189 (N_18189,N_14353,N_13362);
nand U18190 (N_18190,N_10311,N_12019);
or U18191 (N_18191,N_10423,N_10620);
xor U18192 (N_18192,N_14215,N_12535);
nand U18193 (N_18193,N_11082,N_14305);
nor U18194 (N_18194,N_10375,N_10097);
or U18195 (N_18195,N_11378,N_13932);
nand U18196 (N_18196,N_12742,N_12905);
or U18197 (N_18197,N_10663,N_10553);
and U18198 (N_18198,N_11516,N_13629);
or U18199 (N_18199,N_12463,N_12364);
nor U18200 (N_18200,N_11293,N_13840);
or U18201 (N_18201,N_11315,N_13156);
nand U18202 (N_18202,N_10581,N_12791);
nand U18203 (N_18203,N_11348,N_12271);
nor U18204 (N_18204,N_10444,N_14959);
nand U18205 (N_18205,N_13697,N_14288);
and U18206 (N_18206,N_14764,N_14669);
and U18207 (N_18207,N_14574,N_12147);
nor U18208 (N_18208,N_10200,N_14346);
and U18209 (N_18209,N_13169,N_14620);
or U18210 (N_18210,N_14564,N_13053);
and U18211 (N_18211,N_10772,N_12352);
and U18212 (N_18212,N_14676,N_11195);
or U18213 (N_18213,N_13441,N_14676);
or U18214 (N_18214,N_10367,N_13690);
nand U18215 (N_18215,N_14089,N_14703);
nand U18216 (N_18216,N_11316,N_10748);
and U18217 (N_18217,N_10274,N_12069);
and U18218 (N_18218,N_12716,N_11896);
and U18219 (N_18219,N_14324,N_14425);
nor U18220 (N_18220,N_11350,N_13271);
nor U18221 (N_18221,N_10797,N_10876);
nand U18222 (N_18222,N_14915,N_10756);
xor U18223 (N_18223,N_14001,N_13030);
or U18224 (N_18224,N_13593,N_13450);
and U18225 (N_18225,N_12124,N_12379);
or U18226 (N_18226,N_10459,N_13035);
or U18227 (N_18227,N_12319,N_11096);
nand U18228 (N_18228,N_12862,N_14253);
nor U18229 (N_18229,N_11556,N_11393);
and U18230 (N_18230,N_13030,N_10400);
nand U18231 (N_18231,N_13266,N_13365);
nor U18232 (N_18232,N_11303,N_14076);
and U18233 (N_18233,N_13448,N_14297);
or U18234 (N_18234,N_12356,N_14651);
nand U18235 (N_18235,N_14328,N_10372);
nand U18236 (N_18236,N_11981,N_13493);
or U18237 (N_18237,N_14170,N_12678);
or U18238 (N_18238,N_11718,N_12312);
and U18239 (N_18239,N_14947,N_10093);
or U18240 (N_18240,N_11597,N_12553);
nand U18241 (N_18241,N_14026,N_10128);
and U18242 (N_18242,N_12881,N_12434);
nand U18243 (N_18243,N_13131,N_13773);
nand U18244 (N_18244,N_14605,N_12155);
or U18245 (N_18245,N_13686,N_13828);
nand U18246 (N_18246,N_13726,N_12369);
nand U18247 (N_18247,N_12839,N_11449);
and U18248 (N_18248,N_11178,N_14223);
or U18249 (N_18249,N_14990,N_10218);
and U18250 (N_18250,N_13837,N_13459);
nand U18251 (N_18251,N_13820,N_14600);
nand U18252 (N_18252,N_11459,N_13238);
or U18253 (N_18253,N_13927,N_14756);
nor U18254 (N_18254,N_14555,N_14681);
and U18255 (N_18255,N_14813,N_14053);
nor U18256 (N_18256,N_10449,N_13842);
nand U18257 (N_18257,N_12480,N_10401);
or U18258 (N_18258,N_11142,N_10842);
and U18259 (N_18259,N_12157,N_10160);
nor U18260 (N_18260,N_11538,N_12156);
nor U18261 (N_18261,N_11178,N_11228);
and U18262 (N_18262,N_10944,N_11792);
and U18263 (N_18263,N_11911,N_11841);
nor U18264 (N_18264,N_12521,N_11205);
nor U18265 (N_18265,N_12817,N_10980);
and U18266 (N_18266,N_10982,N_10774);
and U18267 (N_18267,N_13874,N_12155);
and U18268 (N_18268,N_10239,N_13456);
nor U18269 (N_18269,N_14296,N_10605);
nand U18270 (N_18270,N_14313,N_14993);
and U18271 (N_18271,N_13517,N_14369);
nand U18272 (N_18272,N_13614,N_12431);
or U18273 (N_18273,N_12268,N_10354);
nand U18274 (N_18274,N_14372,N_11735);
nand U18275 (N_18275,N_13870,N_10509);
or U18276 (N_18276,N_10083,N_11951);
or U18277 (N_18277,N_10564,N_11292);
nand U18278 (N_18278,N_13633,N_10679);
or U18279 (N_18279,N_13178,N_12740);
nand U18280 (N_18280,N_13409,N_12699);
nand U18281 (N_18281,N_12159,N_13234);
and U18282 (N_18282,N_13569,N_14458);
and U18283 (N_18283,N_12596,N_14935);
nand U18284 (N_18284,N_12947,N_13658);
nor U18285 (N_18285,N_14688,N_14396);
xnor U18286 (N_18286,N_13414,N_12363);
nor U18287 (N_18287,N_11010,N_10967);
and U18288 (N_18288,N_14074,N_11076);
and U18289 (N_18289,N_11342,N_12242);
nand U18290 (N_18290,N_14567,N_11192);
and U18291 (N_18291,N_12064,N_14780);
nand U18292 (N_18292,N_14108,N_10824);
or U18293 (N_18293,N_12488,N_13221);
or U18294 (N_18294,N_13891,N_10966);
or U18295 (N_18295,N_13944,N_13982);
nor U18296 (N_18296,N_13826,N_13663);
or U18297 (N_18297,N_11967,N_13341);
nor U18298 (N_18298,N_13312,N_14853);
or U18299 (N_18299,N_11670,N_11018);
or U18300 (N_18300,N_10555,N_13041);
nand U18301 (N_18301,N_10684,N_13437);
and U18302 (N_18302,N_14244,N_11256);
nor U18303 (N_18303,N_13177,N_10195);
or U18304 (N_18304,N_13395,N_11155);
or U18305 (N_18305,N_14602,N_12730);
and U18306 (N_18306,N_14924,N_13044);
or U18307 (N_18307,N_11777,N_14353);
nand U18308 (N_18308,N_13181,N_14874);
nor U18309 (N_18309,N_10932,N_14296);
nor U18310 (N_18310,N_10175,N_14159);
nand U18311 (N_18311,N_13792,N_12723);
nor U18312 (N_18312,N_11197,N_12428);
or U18313 (N_18313,N_14141,N_12905);
nor U18314 (N_18314,N_13122,N_11372);
nor U18315 (N_18315,N_11216,N_11510);
or U18316 (N_18316,N_13759,N_12137);
and U18317 (N_18317,N_11242,N_13007);
and U18318 (N_18318,N_10108,N_14050);
nor U18319 (N_18319,N_10132,N_11924);
and U18320 (N_18320,N_12082,N_14593);
nand U18321 (N_18321,N_14691,N_13911);
nand U18322 (N_18322,N_12066,N_10729);
and U18323 (N_18323,N_10309,N_13597);
nor U18324 (N_18324,N_10876,N_14095);
or U18325 (N_18325,N_12434,N_13323);
nand U18326 (N_18326,N_11342,N_12730);
and U18327 (N_18327,N_12540,N_12506);
and U18328 (N_18328,N_12218,N_12504);
nand U18329 (N_18329,N_11282,N_10176);
and U18330 (N_18330,N_14579,N_12996);
or U18331 (N_18331,N_13695,N_11393);
or U18332 (N_18332,N_10264,N_13076);
and U18333 (N_18333,N_10196,N_10838);
and U18334 (N_18334,N_11856,N_14288);
nor U18335 (N_18335,N_11387,N_13540);
nand U18336 (N_18336,N_12680,N_10188);
and U18337 (N_18337,N_14432,N_14422);
nor U18338 (N_18338,N_11472,N_11072);
nand U18339 (N_18339,N_12912,N_14242);
xnor U18340 (N_18340,N_12729,N_13246);
and U18341 (N_18341,N_14312,N_12126);
nor U18342 (N_18342,N_12767,N_10325);
nor U18343 (N_18343,N_11617,N_13943);
and U18344 (N_18344,N_12823,N_13637);
nand U18345 (N_18345,N_10578,N_11625);
and U18346 (N_18346,N_12540,N_10325);
and U18347 (N_18347,N_11138,N_11687);
nor U18348 (N_18348,N_10812,N_10381);
xor U18349 (N_18349,N_13969,N_12264);
and U18350 (N_18350,N_11607,N_14683);
nor U18351 (N_18351,N_11914,N_12790);
nand U18352 (N_18352,N_11123,N_14456);
nor U18353 (N_18353,N_11135,N_12412);
and U18354 (N_18354,N_13154,N_14406);
and U18355 (N_18355,N_13783,N_12014);
nand U18356 (N_18356,N_10167,N_13796);
nor U18357 (N_18357,N_11216,N_13132);
and U18358 (N_18358,N_12090,N_13188);
nand U18359 (N_18359,N_11148,N_11068);
xor U18360 (N_18360,N_11111,N_10863);
nor U18361 (N_18361,N_12986,N_13845);
and U18362 (N_18362,N_10692,N_12828);
or U18363 (N_18363,N_14489,N_12600);
nor U18364 (N_18364,N_11771,N_10871);
nand U18365 (N_18365,N_12589,N_14327);
xor U18366 (N_18366,N_11838,N_14467);
nand U18367 (N_18367,N_10372,N_10957);
nand U18368 (N_18368,N_14192,N_11873);
nor U18369 (N_18369,N_10709,N_10879);
or U18370 (N_18370,N_13252,N_10045);
and U18371 (N_18371,N_14351,N_14263);
nand U18372 (N_18372,N_11410,N_11230);
and U18373 (N_18373,N_11886,N_14915);
or U18374 (N_18374,N_14777,N_13631);
nand U18375 (N_18375,N_12067,N_11333);
nand U18376 (N_18376,N_10915,N_14429);
and U18377 (N_18377,N_13070,N_13151);
xor U18378 (N_18378,N_14551,N_14003);
nand U18379 (N_18379,N_14410,N_12039);
or U18380 (N_18380,N_13412,N_10973);
nor U18381 (N_18381,N_13600,N_12882);
or U18382 (N_18382,N_14093,N_13901);
and U18383 (N_18383,N_13977,N_10932);
nor U18384 (N_18384,N_11657,N_10071);
nand U18385 (N_18385,N_14185,N_13895);
nand U18386 (N_18386,N_11786,N_13800);
or U18387 (N_18387,N_11915,N_10465);
or U18388 (N_18388,N_11347,N_13867);
nor U18389 (N_18389,N_14708,N_12749);
nor U18390 (N_18390,N_13597,N_11676);
and U18391 (N_18391,N_11232,N_10766);
nor U18392 (N_18392,N_14678,N_14918);
and U18393 (N_18393,N_13637,N_14570);
or U18394 (N_18394,N_11869,N_14789);
or U18395 (N_18395,N_14538,N_13431);
and U18396 (N_18396,N_11254,N_14126);
and U18397 (N_18397,N_11392,N_12585);
or U18398 (N_18398,N_11149,N_12444);
nor U18399 (N_18399,N_12376,N_14036);
or U18400 (N_18400,N_11664,N_13480);
nor U18401 (N_18401,N_11851,N_13137);
nor U18402 (N_18402,N_10296,N_13426);
and U18403 (N_18403,N_12143,N_11003);
or U18404 (N_18404,N_10624,N_10094);
nand U18405 (N_18405,N_11400,N_12070);
nand U18406 (N_18406,N_12873,N_10537);
nor U18407 (N_18407,N_13509,N_11688);
and U18408 (N_18408,N_10242,N_10306);
nor U18409 (N_18409,N_13935,N_11481);
or U18410 (N_18410,N_12933,N_12429);
or U18411 (N_18411,N_10068,N_10568);
nand U18412 (N_18412,N_12717,N_14107);
and U18413 (N_18413,N_10702,N_14927);
and U18414 (N_18414,N_11165,N_10579);
nor U18415 (N_18415,N_14562,N_14023);
and U18416 (N_18416,N_11370,N_13032);
or U18417 (N_18417,N_10659,N_14084);
or U18418 (N_18418,N_10500,N_12034);
and U18419 (N_18419,N_13169,N_11883);
and U18420 (N_18420,N_12330,N_10570);
or U18421 (N_18421,N_11276,N_10561);
nand U18422 (N_18422,N_10994,N_13308);
nand U18423 (N_18423,N_14216,N_11779);
xor U18424 (N_18424,N_13303,N_14858);
or U18425 (N_18425,N_12197,N_14560);
nand U18426 (N_18426,N_14069,N_12194);
or U18427 (N_18427,N_13080,N_14151);
xnor U18428 (N_18428,N_10132,N_11102);
or U18429 (N_18429,N_12637,N_14564);
and U18430 (N_18430,N_13786,N_14463);
nand U18431 (N_18431,N_10466,N_13812);
and U18432 (N_18432,N_10295,N_14576);
nor U18433 (N_18433,N_13378,N_14920);
nor U18434 (N_18434,N_14199,N_14231);
nor U18435 (N_18435,N_14850,N_12816);
nor U18436 (N_18436,N_13926,N_12130);
and U18437 (N_18437,N_12080,N_11889);
nand U18438 (N_18438,N_14027,N_10562);
nand U18439 (N_18439,N_12811,N_14200);
nand U18440 (N_18440,N_11401,N_11375);
nand U18441 (N_18441,N_10173,N_13455);
and U18442 (N_18442,N_12440,N_12606);
nor U18443 (N_18443,N_10700,N_13179);
nor U18444 (N_18444,N_12207,N_14746);
nor U18445 (N_18445,N_13354,N_11911);
or U18446 (N_18446,N_14269,N_11443);
nand U18447 (N_18447,N_12422,N_10253);
nand U18448 (N_18448,N_13185,N_12641);
nor U18449 (N_18449,N_12188,N_13315);
nor U18450 (N_18450,N_10768,N_11150);
or U18451 (N_18451,N_10940,N_11763);
nand U18452 (N_18452,N_11732,N_12617);
nand U18453 (N_18453,N_14952,N_14767);
or U18454 (N_18454,N_11481,N_14891);
nor U18455 (N_18455,N_10849,N_14608);
nor U18456 (N_18456,N_11995,N_12308);
and U18457 (N_18457,N_14173,N_13177);
nor U18458 (N_18458,N_12242,N_13101);
or U18459 (N_18459,N_14063,N_10754);
or U18460 (N_18460,N_10907,N_13043);
nand U18461 (N_18461,N_11837,N_13268);
nor U18462 (N_18462,N_13500,N_14097);
and U18463 (N_18463,N_12178,N_10471);
or U18464 (N_18464,N_12237,N_13391);
nor U18465 (N_18465,N_14163,N_12353);
nor U18466 (N_18466,N_10774,N_13060);
nand U18467 (N_18467,N_13999,N_14997);
and U18468 (N_18468,N_12925,N_10312);
nor U18469 (N_18469,N_13249,N_13094);
nand U18470 (N_18470,N_12024,N_11734);
nor U18471 (N_18471,N_13576,N_10198);
xor U18472 (N_18472,N_10430,N_11247);
nand U18473 (N_18473,N_12357,N_14614);
nand U18474 (N_18474,N_10408,N_13030);
nand U18475 (N_18475,N_12618,N_11248);
nand U18476 (N_18476,N_10687,N_10371);
nand U18477 (N_18477,N_12038,N_13961);
or U18478 (N_18478,N_11761,N_12380);
nand U18479 (N_18479,N_11379,N_13058);
nand U18480 (N_18480,N_10969,N_12330);
nand U18481 (N_18481,N_10318,N_14121);
and U18482 (N_18482,N_11011,N_12519);
and U18483 (N_18483,N_13813,N_10473);
or U18484 (N_18484,N_13184,N_12695);
or U18485 (N_18485,N_13742,N_14561);
and U18486 (N_18486,N_10471,N_11947);
or U18487 (N_18487,N_10075,N_13787);
nand U18488 (N_18488,N_14577,N_12607);
or U18489 (N_18489,N_13819,N_11210);
nand U18490 (N_18490,N_12436,N_10742);
or U18491 (N_18491,N_12032,N_12565);
nor U18492 (N_18492,N_13543,N_12012);
or U18493 (N_18493,N_14434,N_13474);
and U18494 (N_18494,N_10579,N_14036);
and U18495 (N_18495,N_14305,N_14833);
or U18496 (N_18496,N_13533,N_11401);
nor U18497 (N_18497,N_12250,N_13812);
nor U18498 (N_18498,N_10480,N_14016);
and U18499 (N_18499,N_11111,N_12530);
or U18500 (N_18500,N_13208,N_10651);
nor U18501 (N_18501,N_14090,N_10327);
nand U18502 (N_18502,N_12964,N_12879);
and U18503 (N_18503,N_13131,N_14658);
or U18504 (N_18504,N_11202,N_10578);
or U18505 (N_18505,N_13399,N_14365);
nor U18506 (N_18506,N_10539,N_11914);
xor U18507 (N_18507,N_12785,N_11599);
nor U18508 (N_18508,N_11296,N_13065);
nand U18509 (N_18509,N_13467,N_14853);
and U18510 (N_18510,N_11628,N_13107);
nor U18511 (N_18511,N_11573,N_13877);
nand U18512 (N_18512,N_13378,N_12851);
nand U18513 (N_18513,N_13203,N_11189);
or U18514 (N_18514,N_12242,N_14890);
nand U18515 (N_18515,N_10591,N_14351);
or U18516 (N_18516,N_12377,N_13157);
or U18517 (N_18517,N_12758,N_10525);
nand U18518 (N_18518,N_12775,N_12546);
nand U18519 (N_18519,N_11774,N_10730);
nor U18520 (N_18520,N_11641,N_11640);
nor U18521 (N_18521,N_11567,N_10868);
nand U18522 (N_18522,N_13214,N_13960);
nor U18523 (N_18523,N_12373,N_12099);
or U18524 (N_18524,N_13857,N_12326);
or U18525 (N_18525,N_13836,N_14178);
and U18526 (N_18526,N_10701,N_11064);
nor U18527 (N_18527,N_14362,N_14949);
nor U18528 (N_18528,N_13159,N_12642);
nand U18529 (N_18529,N_14227,N_10926);
and U18530 (N_18530,N_14865,N_14175);
nand U18531 (N_18531,N_12845,N_11510);
nand U18532 (N_18532,N_11687,N_10935);
or U18533 (N_18533,N_14726,N_14964);
or U18534 (N_18534,N_11900,N_11907);
nand U18535 (N_18535,N_12436,N_14222);
and U18536 (N_18536,N_13598,N_11770);
and U18537 (N_18537,N_12404,N_14835);
nand U18538 (N_18538,N_14969,N_11056);
or U18539 (N_18539,N_10927,N_10435);
or U18540 (N_18540,N_11856,N_10816);
nand U18541 (N_18541,N_11920,N_12254);
nor U18542 (N_18542,N_10383,N_11376);
nor U18543 (N_18543,N_10538,N_13003);
or U18544 (N_18544,N_13397,N_11880);
nand U18545 (N_18545,N_10378,N_12990);
or U18546 (N_18546,N_12336,N_13138);
nand U18547 (N_18547,N_14558,N_13680);
and U18548 (N_18548,N_11818,N_10168);
nor U18549 (N_18549,N_12953,N_11558);
nand U18550 (N_18550,N_14528,N_10359);
and U18551 (N_18551,N_14305,N_11250);
and U18552 (N_18552,N_14164,N_10250);
xnor U18553 (N_18553,N_11511,N_13365);
nor U18554 (N_18554,N_10803,N_14474);
nand U18555 (N_18555,N_11355,N_12777);
nand U18556 (N_18556,N_10304,N_14970);
xnor U18557 (N_18557,N_12108,N_12528);
nand U18558 (N_18558,N_11792,N_11855);
nand U18559 (N_18559,N_13325,N_14053);
nor U18560 (N_18560,N_10877,N_13043);
and U18561 (N_18561,N_14566,N_14590);
or U18562 (N_18562,N_11373,N_10440);
and U18563 (N_18563,N_14213,N_13871);
or U18564 (N_18564,N_12496,N_13414);
nand U18565 (N_18565,N_11591,N_10107);
nor U18566 (N_18566,N_12819,N_12337);
nor U18567 (N_18567,N_14113,N_10157);
nor U18568 (N_18568,N_11425,N_13459);
nand U18569 (N_18569,N_14635,N_13197);
nand U18570 (N_18570,N_14189,N_12946);
nand U18571 (N_18571,N_14509,N_14937);
nand U18572 (N_18572,N_14100,N_13345);
nand U18573 (N_18573,N_13772,N_13747);
and U18574 (N_18574,N_13356,N_10954);
nor U18575 (N_18575,N_12778,N_12136);
and U18576 (N_18576,N_14538,N_10955);
and U18577 (N_18577,N_13797,N_13065);
nor U18578 (N_18578,N_12025,N_13183);
nor U18579 (N_18579,N_14973,N_10119);
nor U18580 (N_18580,N_10808,N_13153);
nor U18581 (N_18581,N_11447,N_13845);
nand U18582 (N_18582,N_11455,N_12751);
nand U18583 (N_18583,N_11843,N_11369);
or U18584 (N_18584,N_14244,N_12619);
and U18585 (N_18585,N_12143,N_14480);
and U18586 (N_18586,N_13979,N_10711);
nor U18587 (N_18587,N_12822,N_14781);
or U18588 (N_18588,N_10408,N_10130);
and U18589 (N_18589,N_10292,N_12758);
nor U18590 (N_18590,N_11128,N_12272);
nand U18591 (N_18591,N_13828,N_11918);
nand U18592 (N_18592,N_10573,N_14270);
and U18593 (N_18593,N_14023,N_13819);
nor U18594 (N_18594,N_13253,N_10922);
nand U18595 (N_18595,N_14917,N_11926);
and U18596 (N_18596,N_11502,N_13221);
nor U18597 (N_18597,N_11177,N_12491);
and U18598 (N_18598,N_11789,N_12638);
nor U18599 (N_18599,N_10127,N_14620);
nand U18600 (N_18600,N_11130,N_12834);
nand U18601 (N_18601,N_10714,N_11660);
and U18602 (N_18602,N_11141,N_10924);
or U18603 (N_18603,N_14968,N_12551);
nand U18604 (N_18604,N_14205,N_14925);
and U18605 (N_18605,N_11914,N_14532);
nand U18606 (N_18606,N_13975,N_11042);
nor U18607 (N_18607,N_13033,N_11657);
or U18608 (N_18608,N_11811,N_13110);
nand U18609 (N_18609,N_11387,N_12991);
or U18610 (N_18610,N_11284,N_13706);
nand U18611 (N_18611,N_13557,N_14367);
nor U18612 (N_18612,N_12795,N_14131);
nor U18613 (N_18613,N_11705,N_11677);
or U18614 (N_18614,N_11378,N_11211);
or U18615 (N_18615,N_13092,N_14863);
or U18616 (N_18616,N_12205,N_13688);
nor U18617 (N_18617,N_12579,N_12382);
nor U18618 (N_18618,N_13238,N_13909);
or U18619 (N_18619,N_13374,N_12872);
and U18620 (N_18620,N_11211,N_10748);
nor U18621 (N_18621,N_12369,N_13610);
nand U18622 (N_18622,N_14902,N_12477);
nor U18623 (N_18623,N_10627,N_11411);
nand U18624 (N_18624,N_12846,N_14244);
nand U18625 (N_18625,N_11789,N_14816);
nand U18626 (N_18626,N_11116,N_12516);
or U18627 (N_18627,N_10138,N_11094);
nor U18628 (N_18628,N_12098,N_14957);
nand U18629 (N_18629,N_12180,N_14421);
nand U18630 (N_18630,N_14552,N_10039);
nand U18631 (N_18631,N_14845,N_12816);
nor U18632 (N_18632,N_10965,N_13357);
nand U18633 (N_18633,N_13942,N_10837);
and U18634 (N_18634,N_10583,N_11380);
nor U18635 (N_18635,N_14290,N_13920);
nand U18636 (N_18636,N_10375,N_14230);
or U18637 (N_18637,N_10415,N_12628);
nor U18638 (N_18638,N_10818,N_10367);
nor U18639 (N_18639,N_11792,N_11093);
nor U18640 (N_18640,N_14386,N_11518);
or U18641 (N_18641,N_13103,N_14843);
or U18642 (N_18642,N_10253,N_11332);
nand U18643 (N_18643,N_10075,N_14763);
xor U18644 (N_18644,N_11156,N_12118);
nor U18645 (N_18645,N_13185,N_10555);
or U18646 (N_18646,N_12496,N_11782);
and U18647 (N_18647,N_13098,N_13923);
and U18648 (N_18648,N_13232,N_13284);
nand U18649 (N_18649,N_14042,N_10160);
or U18650 (N_18650,N_14104,N_14673);
and U18651 (N_18651,N_14914,N_11572);
or U18652 (N_18652,N_13791,N_11902);
nor U18653 (N_18653,N_10893,N_10854);
nor U18654 (N_18654,N_10686,N_14976);
nand U18655 (N_18655,N_11722,N_13248);
nor U18656 (N_18656,N_13577,N_11721);
nor U18657 (N_18657,N_12936,N_10127);
nor U18658 (N_18658,N_12232,N_13640);
or U18659 (N_18659,N_11355,N_10686);
or U18660 (N_18660,N_13829,N_14249);
nand U18661 (N_18661,N_14102,N_11882);
nor U18662 (N_18662,N_13259,N_11476);
xnor U18663 (N_18663,N_12326,N_11563);
nand U18664 (N_18664,N_12703,N_10345);
nor U18665 (N_18665,N_13578,N_14652);
xor U18666 (N_18666,N_11221,N_10405);
and U18667 (N_18667,N_14615,N_11564);
and U18668 (N_18668,N_12476,N_11964);
nand U18669 (N_18669,N_14053,N_14998);
or U18670 (N_18670,N_11364,N_10407);
or U18671 (N_18671,N_14438,N_14564);
nor U18672 (N_18672,N_11057,N_14376);
and U18673 (N_18673,N_11189,N_13216);
and U18674 (N_18674,N_10205,N_10913);
nand U18675 (N_18675,N_13243,N_12993);
and U18676 (N_18676,N_14534,N_11230);
or U18677 (N_18677,N_14988,N_11883);
or U18678 (N_18678,N_13323,N_11485);
nor U18679 (N_18679,N_11074,N_14268);
or U18680 (N_18680,N_10354,N_13760);
nand U18681 (N_18681,N_12191,N_14161);
or U18682 (N_18682,N_12927,N_11309);
or U18683 (N_18683,N_12679,N_11160);
nand U18684 (N_18684,N_14889,N_11391);
nor U18685 (N_18685,N_14405,N_13995);
and U18686 (N_18686,N_10139,N_11068);
nor U18687 (N_18687,N_11317,N_11022);
and U18688 (N_18688,N_12903,N_12296);
nand U18689 (N_18689,N_12934,N_13033);
nor U18690 (N_18690,N_14251,N_10087);
or U18691 (N_18691,N_13460,N_10404);
or U18692 (N_18692,N_10075,N_12008);
nand U18693 (N_18693,N_12646,N_12486);
or U18694 (N_18694,N_14801,N_12866);
xor U18695 (N_18695,N_10259,N_11984);
and U18696 (N_18696,N_12285,N_12659);
nand U18697 (N_18697,N_10565,N_12914);
nor U18698 (N_18698,N_10211,N_13184);
nor U18699 (N_18699,N_11163,N_14454);
nor U18700 (N_18700,N_14534,N_14349);
nand U18701 (N_18701,N_14233,N_14478);
xnor U18702 (N_18702,N_13991,N_14995);
and U18703 (N_18703,N_11158,N_14926);
nand U18704 (N_18704,N_13821,N_13987);
and U18705 (N_18705,N_10075,N_11276);
and U18706 (N_18706,N_13090,N_11791);
and U18707 (N_18707,N_10322,N_13659);
and U18708 (N_18708,N_11672,N_10663);
nor U18709 (N_18709,N_11728,N_13176);
and U18710 (N_18710,N_11173,N_11983);
nand U18711 (N_18711,N_12326,N_10523);
or U18712 (N_18712,N_11602,N_14414);
or U18713 (N_18713,N_10014,N_11197);
nand U18714 (N_18714,N_13896,N_10238);
nand U18715 (N_18715,N_12070,N_12201);
nand U18716 (N_18716,N_12987,N_12824);
and U18717 (N_18717,N_10921,N_13645);
nor U18718 (N_18718,N_13273,N_14216);
or U18719 (N_18719,N_14835,N_14479);
and U18720 (N_18720,N_13877,N_11510);
or U18721 (N_18721,N_11722,N_11187);
or U18722 (N_18722,N_13654,N_12065);
nand U18723 (N_18723,N_14833,N_13779);
nand U18724 (N_18724,N_12914,N_14642);
nor U18725 (N_18725,N_14699,N_10375);
nand U18726 (N_18726,N_14246,N_10359);
nor U18727 (N_18727,N_13897,N_10719);
nor U18728 (N_18728,N_10281,N_11253);
and U18729 (N_18729,N_10644,N_12982);
and U18730 (N_18730,N_14605,N_11205);
and U18731 (N_18731,N_12844,N_11763);
nor U18732 (N_18732,N_14408,N_12619);
xnor U18733 (N_18733,N_13933,N_11769);
and U18734 (N_18734,N_14269,N_14211);
and U18735 (N_18735,N_14914,N_12387);
nor U18736 (N_18736,N_10886,N_13106);
nor U18737 (N_18737,N_11495,N_13367);
or U18738 (N_18738,N_10588,N_14887);
and U18739 (N_18739,N_13062,N_10990);
nor U18740 (N_18740,N_12140,N_12185);
and U18741 (N_18741,N_14653,N_14148);
nand U18742 (N_18742,N_10706,N_12719);
nor U18743 (N_18743,N_14032,N_14136);
nand U18744 (N_18744,N_14224,N_14098);
or U18745 (N_18745,N_12539,N_10678);
nand U18746 (N_18746,N_14789,N_12316);
or U18747 (N_18747,N_12614,N_14318);
nand U18748 (N_18748,N_10455,N_13804);
nand U18749 (N_18749,N_12211,N_10584);
xor U18750 (N_18750,N_11732,N_14618);
or U18751 (N_18751,N_11497,N_12346);
or U18752 (N_18752,N_13238,N_14098);
and U18753 (N_18753,N_12397,N_10814);
and U18754 (N_18754,N_10306,N_11987);
or U18755 (N_18755,N_12404,N_10545);
and U18756 (N_18756,N_10580,N_12416);
or U18757 (N_18757,N_12250,N_13843);
and U18758 (N_18758,N_14567,N_14040);
nand U18759 (N_18759,N_14165,N_10405);
and U18760 (N_18760,N_13422,N_11070);
nand U18761 (N_18761,N_10798,N_14514);
or U18762 (N_18762,N_12007,N_10775);
nand U18763 (N_18763,N_10609,N_14766);
and U18764 (N_18764,N_10610,N_13211);
nor U18765 (N_18765,N_13468,N_14184);
and U18766 (N_18766,N_11552,N_10102);
and U18767 (N_18767,N_14895,N_10567);
nand U18768 (N_18768,N_14172,N_11163);
and U18769 (N_18769,N_12697,N_10677);
xnor U18770 (N_18770,N_14592,N_11546);
nand U18771 (N_18771,N_11351,N_14571);
nor U18772 (N_18772,N_11539,N_11486);
nor U18773 (N_18773,N_14026,N_12506);
and U18774 (N_18774,N_11111,N_14420);
or U18775 (N_18775,N_12409,N_14748);
nor U18776 (N_18776,N_10131,N_12848);
nand U18777 (N_18777,N_10631,N_14920);
nand U18778 (N_18778,N_10451,N_10057);
nor U18779 (N_18779,N_10346,N_10896);
nor U18780 (N_18780,N_13020,N_14401);
or U18781 (N_18781,N_12087,N_10118);
nand U18782 (N_18782,N_14447,N_14107);
or U18783 (N_18783,N_10118,N_11822);
and U18784 (N_18784,N_10273,N_10111);
nor U18785 (N_18785,N_10992,N_13188);
nor U18786 (N_18786,N_12087,N_12041);
and U18787 (N_18787,N_11196,N_13496);
nand U18788 (N_18788,N_11644,N_12610);
nor U18789 (N_18789,N_13556,N_11639);
nor U18790 (N_18790,N_10086,N_11654);
nand U18791 (N_18791,N_13237,N_14315);
nand U18792 (N_18792,N_12347,N_12019);
nand U18793 (N_18793,N_11029,N_14460);
nand U18794 (N_18794,N_10187,N_14924);
and U18795 (N_18795,N_13454,N_11235);
nand U18796 (N_18796,N_12532,N_13516);
or U18797 (N_18797,N_11520,N_14437);
or U18798 (N_18798,N_14488,N_14487);
nor U18799 (N_18799,N_11293,N_14838);
and U18800 (N_18800,N_10491,N_14017);
or U18801 (N_18801,N_10430,N_14401);
or U18802 (N_18802,N_11015,N_11746);
and U18803 (N_18803,N_13376,N_12927);
nor U18804 (N_18804,N_11735,N_11400);
xnor U18805 (N_18805,N_10010,N_12417);
xnor U18806 (N_18806,N_12633,N_14182);
nor U18807 (N_18807,N_13696,N_13560);
nand U18808 (N_18808,N_11038,N_11973);
nor U18809 (N_18809,N_11391,N_14700);
nor U18810 (N_18810,N_10024,N_14476);
nor U18811 (N_18811,N_14503,N_10121);
and U18812 (N_18812,N_14748,N_14707);
nand U18813 (N_18813,N_11834,N_10575);
and U18814 (N_18814,N_10599,N_12478);
nand U18815 (N_18815,N_11281,N_14680);
or U18816 (N_18816,N_11140,N_14088);
nor U18817 (N_18817,N_10659,N_10051);
nor U18818 (N_18818,N_12037,N_14294);
nor U18819 (N_18819,N_13251,N_11587);
and U18820 (N_18820,N_10721,N_14953);
and U18821 (N_18821,N_10938,N_14114);
or U18822 (N_18822,N_11354,N_11242);
or U18823 (N_18823,N_10922,N_11153);
nor U18824 (N_18824,N_10691,N_10233);
nor U18825 (N_18825,N_13295,N_11131);
nor U18826 (N_18826,N_14513,N_11875);
nor U18827 (N_18827,N_12952,N_13473);
or U18828 (N_18828,N_13909,N_13411);
nand U18829 (N_18829,N_12657,N_13377);
and U18830 (N_18830,N_10099,N_14367);
and U18831 (N_18831,N_12160,N_14227);
or U18832 (N_18832,N_11713,N_14181);
nand U18833 (N_18833,N_14422,N_14876);
or U18834 (N_18834,N_13087,N_13783);
nand U18835 (N_18835,N_14761,N_13331);
and U18836 (N_18836,N_11113,N_14241);
nand U18837 (N_18837,N_12929,N_14284);
and U18838 (N_18838,N_14596,N_13507);
or U18839 (N_18839,N_13154,N_12321);
or U18840 (N_18840,N_11427,N_10878);
and U18841 (N_18841,N_14916,N_13886);
nor U18842 (N_18842,N_14326,N_11886);
nor U18843 (N_18843,N_10459,N_12220);
or U18844 (N_18844,N_10990,N_11535);
or U18845 (N_18845,N_13845,N_14072);
or U18846 (N_18846,N_11594,N_14438);
or U18847 (N_18847,N_14753,N_12684);
and U18848 (N_18848,N_10772,N_11924);
or U18849 (N_18849,N_11291,N_10211);
nand U18850 (N_18850,N_10493,N_10721);
and U18851 (N_18851,N_13047,N_10929);
or U18852 (N_18852,N_11119,N_11869);
nand U18853 (N_18853,N_13459,N_10029);
and U18854 (N_18854,N_13241,N_10123);
nand U18855 (N_18855,N_10612,N_10083);
or U18856 (N_18856,N_10981,N_14371);
or U18857 (N_18857,N_12460,N_10083);
xor U18858 (N_18858,N_12714,N_14334);
nor U18859 (N_18859,N_14726,N_13549);
or U18860 (N_18860,N_12309,N_12445);
nor U18861 (N_18861,N_12118,N_11673);
nand U18862 (N_18862,N_14938,N_13682);
xor U18863 (N_18863,N_12175,N_13422);
or U18864 (N_18864,N_13225,N_13096);
nor U18865 (N_18865,N_11951,N_12540);
nor U18866 (N_18866,N_13344,N_12322);
or U18867 (N_18867,N_11038,N_12642);
and U18868 (N_18868,N_11860,N_12279);
or U18869 (N_18869,N_14251,N_13139);
nor U18870 (N_18870,N_10304,N_12310);
nand U18871 (N_18871,N_11860,N_12793);
nor U18872 (N_18872,N_13322,N_10939);
or U18873 (N_18873,N_12425,N_13157);
or U18874 (N_18874,N_12536,N_10202);
nor U18875 (N_18875,N_10151,N_10926);
nor U18876 (N_18876,N_14996,N_12600);
xor U18877 (N_18877,N_12917,N_10302);
nand U18878 (N_18878,N_13691,N_12531);
or U18879 (N_18879,N_10377,N_12950);
xnor U18880 (N_18880,N_10254,N_10300);
and U18881 (N_18881,N_10139,N_11142);
and U18882 (N_18882,N_11737,N_14440);
or U18883 (N_18883,N_12571,N_12794);
nand U18884 (N_18884,N_10936,N_12093);
or U18885 (N_18885,N_12840,N_12578);
or U18886 (N_18886,N_13704,N_11015);
and U18887 (N_18887,N_14862,N_14404);
or U18888 (N_18888,N_10762,N_12696);
nand U18889 (N_18889,N_14778,N_12600);
and U18890 (N_18890,N_12121,N_11781);
nand U18891 (N_18891,N_13414,N_13772);
nand U18892 (N_18892,N_12275,N_11343);
and U18893 (N_18893,N_10063,N_11873);
or U18894 (N_18894,N_13339,N_14489);
nor U18895 (N_18895,N_10093,N_11595);
nor U18896 (N_18896,N_12164,N_14300);
and U18897 (N_18897,N_14102,N_13152);
nor U18898 (N_18898,N_13213,N_13570);
and U18899 (N_18899,N_11197,N_11056);
nand U18900 (N_18900,N_14794,N_10383);
or U18901 (N_18901,N_10879,N_11169);
xor U18902 (N_18902,N_14300,N_13229);
or U18903 (N_18903,N_14463,N_14500);
or U18904 (N_18904,N_12723,N_14034);
and U18905 (N_18905,N_10312,N_11203);
nor U18906 (N_18906,N_12594,N_11658);
nor U18907 (N_18907,N_11437,N_12035);
nor U18908 (N_18908,N_11606,N_10319);
nand U18909 (N_18909,N_12221,N_13317);
nand U18910 (N_18910,N_10318,N_14015);
nor U18911 (N_18911,N_11921,N_13349);
or U18912 (N_18912,N_12755,N_13189);
nand U18913 (N_18913,N_12889,N_13178);
xor U18914 (N_18914,N_10931,N_12902);
or U18915 (N_18915,N_14624,N_10782);
and U18916 (N_18916,N_12966,N_14531);
nand U18917 (N_18917,N_14948,N_10612);
nand U18918 (N_18918,N_10473,N_13242);
nand U18919 (N_18919,N_14023,N_13653);
nand U18920 (N_18920,N_13700,N_10848);
nand U18921 (N_18921,N_14170,N_12583);
and U18922 (N_18922,N_12304,N_11198);
nor U18923 (N_18923,N_13778,N_12791);
nor U18924 (N_18924,N_10286,N_12944);
nand U18925 (N_18925,N_10678,N_11034);
and U18926 (N_18926,N_13999,N_12171);
and U18927 (N_18927,N_11423,N_14239);
or U18928 (N_18928,N_10386,N_14095);
or U18929 (N_18929,N_10854,N_10379);
and U18930 (N_18930,N_14689,N_11145);
and U18931 (N_18931,N_11672,N_10946);
and U18932 (N_18932,N_14292,N_10347);
or U18933 (N_18933,N_12257,N_10589);
or U18934 (N_18934,N_14082,N_13490);
or U18935 (N_18935,N_14424,N_13476);
or U18936 (N_18936,N_11068,N_11946);
or U18937 (N_18937,N_10206,N_13461);
nor U18938 (N_18938,N_13749,N_10767);
nand U18939 (N_18939,N_12113,N_11890);
or U18940 (N_18940,N_10573,N_10075);
or U18941 (N_18941,N_11407,N_13843);
or U18942 (N_18942,N_10310,N_12605);
nand U18943 (N_18943,N_14061,N_14082);
nand U18944 (N_18944,N_12752,N_14123);
nor U18945 (N_18945,N_12144,N_14304);
or U18946 (N_18946,N_13439,N_11407);
nand U18947 (N_18947,N_11775,N_10756);
nand U18948 (N_18948,N_11805,N_14317);
or U18949 (N_18949,N_11003,N_10332);
and U18950 (N_18950,N_14186,N_13539);
or U18951 (N_18951,N_12674,N_13883);
and U18952 (N_18952,N_13879,N_10977);
and U18953 (N_18953,N_11552,N_14859);
and U18954 (N_18954,N_14615,N_13001);
or U18955 (N_18955,N_13881,N_14599);
nand U18956 (N_18956,N_10386,N_11046);
nand U18957 (N_18957,N_13560,N_11745);
nand U18958 (N_18958,N_13038,N_10270);
nand U18959 (N_18959,N_14734,N_12044);
and U18960 (N_18960,N_10813,N_10785);
nand U18961 (N_18961,N_13960,N_10760);
and U18962 (N_18962,N_10150,N_12893);
nor U18963 (N_18963,N_11163,N_10436);
or U18964 (N_18964,N_13066,N_11750);
xor U18965 (N_18965,N_11312,N_10419);
or U18966 (N_18966,N_14484,N_14441);
or U18967 (N_18967,N_14878,N_11587);
nand U18968 (N_18968,N_13038,N_11075);
or U18969 (N_18969,N_12966,N_10184);
nor U18970 (N_18970,N_13061,N_11943);
nand U18971 (N_18971,N_13906,N_14815);
xor U18972 (N_18972,N_10699,N_10784);
nor U18973 (N_18973,N_14669,N_11091);
and U18974 (N_18974,N_11011,N_11975);
or U18975 (N_18975,N_11484,N_14582);
nand U18976 (N_18976,N_10799,N_12970);
xnor U18977 (N_18977,N_13785,N_11972);
and U18978 (N_18978,N_11184,N_13556);
nand U18979 (N_18979,N_14618,N_13852);
and U18980 (N_18980,N_13199,N_14524);
nand U18981 (N_18981,N_12939,N_14738);
or U18982 (N_18982,N_13951,N_14569);
nand U18983 (N_18983,N_14117,N_11906);
nand U18984 (N_18984,N_10778,N_12447);
nor U18985 (N_18985,N_11213,N_14067);
nor U18986 (N_18986,N_10907,N_14945);
or U18987 (N_18987,N_14235,N_14987);
xor U18988 (N_18988,N_13136,N_12336);
nand U18989 (N_18989,N_14271,N_14120);
and U18990 (N_18990,N_11534,N_13126);
nor U18991 (N_18991,N_11423,N_11872);
nand U18992 (N_18992,N_14299,N_10884);
and U18993 (N_18993,N_14363,N_11778);
or U18994 (N_18994,N_11537,N_10435);
nor U18995 (N_18995,N_12945,N_10776);
or U18996 (N_18996,N_11002,N_14418);
or U18997 (N_18997,N_14748,N_11023);
and U18998 (N_18998,N_14451,N_10570);
nand U18999 (N_18999,N_14263,N_13052);
nand U19000 (N_19000,N_11309,N_13833);
nor U19001 (N_19001,N_11173,N_11170);
or U19002 (N_19002,N_10070,N_11123);
or U19003 (N_19003,N_13256,N_10470);
or U19004 (N_19004,N_14612,N_13724);
or U19005 (N_19005,N_10166,N_12946);
or U19006 (N_19006,N_10252,N_10978);
and U19007 (N_19007,N_12898,N_10182);
nand U19008 (N_19008,N_12657,N_12029);
or U19009 (N_19009,N_12691,N_10742);
and U19010 (N_19010,N_12645,N_11374);
and U19011 (N_19011,N_14676,N_14719);
and U19012 (N_19012,N_10659,N_11859);
and U19013 (N_19013,N_14209,N_12850);
and U19014 (N_19014,N_11449,N_12423);
nor U19015 (N_19015,N_12092,N_10768);
and U19016 (N_19016,N_13539,N_13589);
and U19017 (N_19017,N_10270,N_14738);
nand U19018 (N_19018,N_12940,N_13845);
nand U19019 (N_19019,N_12696,N_12090);
or U19020 (N_19020,N_14452,N_10014);
nor U19021 (N_19021,N_14258,N_13079);
nor U19022 (N_19022,N_13703,N_12340);
nand U19023 (N_19023,N_12942,N_10495);
nor U19024 (N_19024,N_12100,N_12698);
and U19025 (N_19025,N_11105,N_11038);
and U19026 (N_19026,N_11164,N_12923);
or U19027 (N_19027,N_10958,N_13589);
nor U19028 (N_19028,N_10333,N_12996);
nor U19029 (N_19029,N_10067,N_11748);
nor U19030 (N_19030,N_10478,N_12618);
or U19031 (N_19031,N_13499,N_11834);
nand U19032 (N_19032,N_11273,N_12204);
nand U19033 (N_19033,N_13256,N_13134);
nor U19034 (N_19034,N_10272,N_13633);
and U19035 (N_19035,N_14472,N_11819);
or U19036 (N_19036,N_13675,N_10915);
or U19037 (N_19037,N_14543,N_13248);
nand U19038 (N_19038,N_14937,N_11402);
nand U19039 (N_19039,N_14183,N_14607);
nor U19040 (N_19040,N_12707,N_13412);
or U19041 (N_19041,N_14863,N_12304);
nand U19042 (N_19042,N_14835,N_13568);
nor U19043 (N_19043,N_11668,N_11018);
nand U19044 (N_19044,N_10227,N_11126);
nor U19045 (N_19045,N_12577,N_10133);
or U19046 (N_19046,N_11324,N_10720);
nor U19047 (N_19047,N_14777,N_14539);
or U19048 (N_19048,N_13452,N_14272);
nor U19049 (N_19049,N_12282,N_10947);
nor U19050 (N_19050,N_11345,N_13543);
and U19051 (N_19051,N_14417,N_10482);
nand U19052 (N_19052,N_10896,N_11921);
nand U19053 (N_19053,N_11547,N_11077);
or U19054 (N_19054,N_12296,N_12491);
or U19055 (N_19055,N_10920,N_10904);
nor U19056 (N_19056,N_10802,N_14771);
nor U19057 (N_19057,N_12625,N_11733);
nand U19058 (N_19058,N_12250,N_14988);
or U19059 (N_19059,N_12093,N_11293);
and U19060 (N_19060,N_10391,N_11419);
nor U19061 (N_19061,N_14837,N_11700);
and U19062 (N_19062,N_14183,N_14281);
nand U19063 (N_19063,N_13275,N_10403);
nand U19064 (N_19064,N_11080,N_12082);
or U19065 (N_19065,N_11946,N_13165);
nand U19066 (N_19066,N_12240,N_13599);
and U19067 (N_19067,N_10344,N_12964);
or U19068 (N_19068,N_12793,N_14216);
nand U19069 (N_19069,N_10053,N_11879);
nand U19070 (N_19070,N_14973,N_12388);
nand U19071 (N_19071,N_12487,N_13241);
nand U19072 (N_19072,N_11606,N_12697);
and U19073 (N_19073,N_13050,N_14295);
or U19074 (N_19074,N_14995,N_14796);
nand U19075 (N_19075,N_11721,N_14234);
or U19076 (N_19076,N_11868,N_13331);
nor U19077 (N_19077,N_12686,N_12831);
nand U19078 (N_19078,N_14185,N_11457);
nand U19079 (N_19079,N_11587,N_11578);
nor U19080 (N_19080,N_12990,N_12361);
or U19081 (N_19081,N_13360,N_10329);
xnor U19082 (N_19082,N_10196,N_12581);
nor U19083 (N_19083,N_14105,N_12219);
nor U19084 (N_19084,N_12137,N_14314);
and U19085 (N_19085,N_14237,N_11355);
and U19086 (N_19086,N_11068,N_12939);
nand U19087 (N_19087,N_12466,N_10527);
nand U19088 (N_19088,N_11157,N_10086);
nand U19089 (N_19089,N_14592,N_14942);
or U19090 (N_19090,N_14214,N_12735);
and U19091 (N_19091,N_11912,N_14797);
or U19092 (N_19092,N_10199,N_10838);
nand U19093 (N_19093,N_11645,N_10145);
nor U19094 (N_19094,N_10824,N_10111);
xor U19095 (N_19095,N_11185,N_14255);
nand U19096 (N_19096,N_10320,N_14938);
nand U19097 (N_19097,N_12012,N_14519);
nand U19098 (N_19098,N_10245,N_11286);
xnor U19099 (N_19099,N_13468,N_14858);
and U19100 (N_19100,N_11769,N_14232);
and U19101 (N_19101,N_13943,N_14890);
and U19102 (N_19102,N_11479,N_12908);
nand U19103 (N_19103,N_14745,N_10197);
nand U19104 (N_19104,N_13503,N_10965);
nand U19105 (N_19105,N_10400,N_11088);
and U19106 (N_19106,N_13922,N_10485);
or U19107 (N_19107,N_10417,N_13300);
or U19108 (N_19108,N_12502,N_14253);
nand U19109 (N_19109,N_12242,N_14195);
nand U19110 (N_19110,N_11200,N_14760);
nand U19111 (N_19111,N_13490,N_13220);
or U19112 (N_19112,N_14572,N_13611);
and U19113 (N_19113,N_13784,N_10615);
or U19114 (N_19114,N_10066,N_12929);
nor U19115 (N_19115,N_14490,N_13046);
or U19116 (N_19116,N_13743,N_12600);
nor U19117 (N_19117,N_11157,N_10390);
nand U19118 (N_19118,N_11682,N_10851);
nand U19119 (N_19119,N_11694,N_14179);
nor U19120 (N_19120,N_14817,N_12489);
and U19121 (N_19121,N_12400,N_11447);
nand U19122 (N_19122,N_13480,N_14664);
or U19123 (N_19123,N_10439,N_10238);
nor U19124 (N_19124,N_14514,N_14747);
or U19125 (N_19125,N_12070,N_10992);
xnor U19126 (N_19126,N_11159,N_14566);
or U19127 (N_19127,N_11629,N_14348);
or U19128 (N_19128,N_12864,N_12901);
or U19129 (N_19129,N_11064,N_14438);
nand U19130 (N_19130,N_11540,N_13807);
and U19131 (N_19131,N_14563,N_12427);
or U19132 (N_19132,N_12039,N_10128);
nand U19133 (N_19133,N_12572,N_12198);
nor U19134 (N_19134,N_11000,N_14773);
nand U19135 (N_19135,N_12772,N_12131);
nor U19136 (N_19136,N_11988,N_14314);
nor U19137 (N_19137,N_14394,N_13018);
or U19138 (N_19138,N_14049,N_10724);
and U19139 (N_19139,N_14416,N_12872);
and U19140 (N_19140,N_14698,N_10721);
nand U19141 (N_19141,N_11822,N_14405);
or U19142 (N_19142,N_11178,N_14669);
nand U19143 (N_19143,N_14560,N_10951);
or U19144 (N_19144,N_13744,N_10647);
nor U19145 (N_19145,N_13649,N_12401);
and U19146 (N_19146,N_14979,N_12873);
and U19147 (N_19147,N_14359,N_14599);
or U19148 (N_19148,N_10506,N_11016);
and U19149 (N_19149,N_14479,N_11866);
nor U19150 (N_19150,N_10304,N_13848);
nor U19151 (N_19151,N_10097,N_11172);
or U19152 (N_19152,N_12367,N_10808);
or U19153 (N_19153,N_12909,N_14955);
or U19154 (N_19154,N_12824,N_13277);
or U19155 (N_19155,N_13809,N_10332);
or U19156 (N_19156,N_14475,N_13908);
nor U19157 (N_19157,N_12055,N_12718);
nor U19158 (N_19158,N_12628,N_11367);
or U19159 (N_19159,N_13878,N_12068);
nand U19160 (N_19160,N_13763,N_14848);
or U19161 (N_19161,N_13260,N_10082);
nand U19162 (N_19162,N_10488,N_10664);
nand U19163 (N_19163,N_10378,N_12420);
or U19164 (N_19164,N_11825,N_11855);
and U19165 (N_19165,N_14797,N_14037);
nand U19166 (N_19166,N_13076,N_13848);
or U19167 (N_19167,N_14255,N_13661);
nor U19168 (N_19168,N_14286,N_11662);
nor U19169 (N_19169,N_13658,N_11539);
or U19170 (N_19170,N_13104,N_11179);
nor U19171 (N_19171,N_10994,N_11507);
nor U19172 (N_19172,N_12322,N_10219);
or U19173 (N_19173,N_11194,N_12814);
nor U19174 (N_19174,N_14331,N_11931);
or U19175 (N_19175,N_13259,N_12580);
and U19176 (N_19176,N_12932,N_10868);
nor U19177 (N_19177,N_10597,N_14761);
and U19178 (N_19178,N_12635,N_10629);
nor U19179 (N_19179,N_10077,N_14195);
nand U19180 (N_19180,N_14106,N_14780);
xor U19181 (N_19181,N_14728,N_14604);
and U19182 (N_19182,N_11446,N_14517);
xnor U19183 (N_19183,N_14115,N_11660);
and U19184 (N_19184,N_11408,N_12231);
and U19185 (N_19185,N_13053,N_13510);
nand U19186 (N_19186,N_11056,N_12462);
or U19187 (N_19187,N_13819,N_14587);
or U19188 (N_19188,N_10564,N_10828);
or U19189 (N_19189,N_12692,N_13737);
nor U19190 (N_19190,N_12948,N_10307);
or U19191 (N_19191,N_14403,N_14538);
nor U19192 (N_19192,N_10882,N_12834);
nor U19193 (N_19193,N_10900,N_10324);
nor U19194 (N_19194,N_13860,N_14907);
or U19195 (N_19195,N_11111,N_12535);
nor U19196 (N_19196,N_10060,N_13169);
and U19197 (N_19197,N_13216,N_13150);
nand U19198 (N_19198,N_12214,N_10968);
and U19199 (N_19199,N_13675,N_14746);
nor U19200 (N_19200,N_11492,N_12347);
and U19201 (N_19201,N_13709,N_13889);
nand U19202 (N_19202,N_14420,N_10017);
or U19203 (N_19203,N_11889,N_12388);
nor U19204 (N_19204,N_11518,N_11350);
nand U19205 (N_19205,N_10114,N_10852);
and U19206 (N_19206,N_10165,N_13636);
nor U19207 (N_19207,N_13912,N_10518);
or U19208 (N_19208,N_12791,N_11113);
nand U19209 (N_19209,N_13218,N_10471);
and U19210 (N_19210,N_12749,N_14698);
and U19211 (N_19211,N_11984,N_10242);
or U19212 (N_19212,N_11381,N_14962);
or U19213 (N_19213,N_14656,N_12385);
nor U19214 (N_19214,N_12512,N_10573);
nor U19215 (N_19215,N_13843,N_10202);
nor U19216 (N_19216,N_11913,N_14284);
nand U19217 (N_19217,N_14672,N_12835);
nor U19218 (N_19218,N_13431,N_14068);
and U19219 (N_19219,N_11594,N_12485);
or U19220 (N_19220,N_10076,N_11218);
or U19221 (N_19221,N_11886,N_13463);
and U19222 (N_19222,N_12380,N_11344);
nand U19223 (N_19223,N_12516,N_13441);
nor U19224 (N_19224,N_11725,N_10921);
and U19225 (N_19225,N_11254,N_11873);
nor U19226 (N_19226,N_14930,N_10604);
or U19227 (N_19227,N_12088,N_14165);
nor U19228 (N_19228,N_14109,N_11061);
nand U19229 (N_19229,N_11980,N_11303);
nor U19230 (N_19230,N_10593,N_12971);
or U19231 (N_19231,N_10226,N_10055);
nand U19232 (N_19232,N_13328,N_13077);
nand U19233 (N_19233,N_12106,N_13270);
and U19234 (N_19234,N_13792,N_13677);
nor U19235 (N_19235,N_11380,N_12984);
and U19236 (N_19236,N_11095,N_14619);
nand U19237 (N_19237,N_14536,N_13429);
nand U19238 (N_19238,N_10406,N_14735);
nor U19239 (N_19239,N_13793,N_10040);
or U19240 (N_19240,N_10749,N_14333);
and U19241 (N_19241,N_11719,N_13355);
nand U19242 (N_19242,N_10426,N_11519);
or U19243 (N_19243,N_10382,N_10476);
nor U19244 (N_19244,N_14728,N_10347);
and U19245 (N_19245,N_10591,N_10407);
or U19246 (N_19246,N_10467,N_12177);
nor U19247 (N_19247,N_13479,N_12147);
nor U19248 (N_19248,N_13084,N_13223);
and U19249 (N_19249,N_13030,N_14077);
nor U19250 (N_19250,N_10030,N_13791);
nand U19251 (N_19251,N_10450,N_12164);
xor U19252 (N_19252,N_11319,N_10360);
nand U19253 (N_19253,N_12396,N_12429);
nor U19254 (N_19254,N_11647,N_14366);
and U19255 (N_19255,N_11199,N_12772);
nor U19256 (N_19256,N_14227,N_13293);
nor U19257 (N_19257,N_13898,N_14534);
nand U19258 (N_19258,N_14618,N_14163);
or U19259 (N_19259,N_10429,N_12927);
nand U19260 (N_19260,N_12543,N_13776);
or U19261 (N_19261,N_11336,N_10395);
nand U19262 (N_19262,N_12097,N_10761);
xor U19263 (N_19263,N_12784,N_14857);
or U19264 (N_19264,N_10200,N_10569);
or U19265 (N_19265,N_13922,N_12478);
xnor U19266 (N_19266,N_10953,N_11391);
nor U19267 (N_19267,N_11836,N_11118);
or U19268 (N_19268,N_14669,N_14504);
or U19269 (N_19269,N_13586,N_12780);
nand U19270 (N_19270,N_13828,N_12141);
and U19271 (N_19271,N_10127,N_11859);
nor U19272 (N_19272,N_14570,N_14356);
nand U19273 (N_19273,N_14145,N_14752);
and U19274 (N_19274,N_10659,N_11028);
or U19275 (N_19275,N_10423,N_12163);
and U19276 (N_19276,N_11107,N_14219);
or U19277 (N_19277,N_11803,N_13940);
and U19278 (N_19278,N_14980,N_10396);
nand U19279 (N_19279,N_13218,N_10743);
nand U19280 (N_19280,N_14779,N_12324);
or U19281 (N_19281,N_14130,N_12270);
nor U19282 (N_19282,N_14273,N_12722);
xnor U19283 (N_19283,N_14001,N_13425);
and U19284 (N_19284,N_11650,N_14803);
or U19285 (N_19285,N_12403,N_14110);
and U19286 (N_19286,N_13034,N_11017);
nand U19287 (N_19287,N_11471,N_12350);
or U19288 (N_19288,N_14696,N_13070);
nor U19289 (N_19289,N_11997,N_12783);
nand U19290 (N_19290,N_11913,N_14304);
and U19291 (N_19291,N_11442,N_11471);
nand U19292 (N_19292,N_14254,N_11209);
nand U19293 (N_19293,N_11510,N_13569);
or U19294 (N_19294,N_12971,N_14704);
and U19295 (N_19295,N_10748,N_12835);
or U19296 (N_19296,N_14478,N_14056);
nand U19297 (N_19297,N_14535,N_10416);
or U19298 (N_19298,N_12790,N_13380);
and U19299 (N_19299,N_13477,N_11793);
xnor U19300 (N_19300,N_10561,N_11816);
nand U19301 (N_19301,N_10790,N_12248);
nor U19302 (N_19302,N_14621,N_12936);
and U19303 (N_19303,N_11866,N_11407);
nor U19304 (N_19304,N_13414,N_11986);
nor U19305 (N_19305,N_11914,N_12820);
nor U19306 (N_19306,N_13302,N_13312);
nand U19307 (N_19307,N_11566,N_11438);
nand U19308 (N_19308,N_14709,N_13462);
and U19309 (N_19309,N_12358,N_11212);
nand U19310 (N_19310,N_14604,N_12282);
or U19311 (N_19311,N_11596,N_14512);
and U19312 (N_19312,N_10705,N_11801);
nand U19313 (N_19313,N_10503,N_13098);
and U19314 (N_19314,N_10237,N_10443);
nor U19315 (N_19315,N_14059,N_12777);
nand U19316 (N_19316,N_10923,N_14231);
nand U19317 (N_19317,N_10438,N_14918);
nor U19318 (N_19318,N_13406,N_11787);
nor U19319 (N_19319,N_12183,N_12108);
nor U19320 (N_19320,N_10755,N_14581);
and U19321 (N_19321,N_12721,N_13308);
and U19322 (N_19322,N_11180,N_13393);
nor U19323 (N_19323,N_14445,N_14749);
or U19324 (N_19324,N_12221,N_12441);
or U19325 (N_19325,N_10508,N_13207);
and U19326 (N_19326,N_14491,N_14424);
nand U19327 (N_19327,N_13202,N_12656);
nand U19328 (N_19328,N_11448,N_14928);
nand U19329 (N_19329,N_13504,N_11425);
or U19330 (N_19330,N_10532,N_13587);
nor U19331 (N_19331,N_11521,N_14149);
nor U19332 (N_19332,N_11643,N_14308);
or U19333 (N_19333,N_13257,N_11605);
and U19334 (N_19334,N_13479,N_13170);
nand U19335 (N_19335,N_12211,N_13693);
xor U19336 (N_19336,N_10498,N_14848);
xnor U19337 (N_19337,N_12868,N_11726);
nand U19338 (N_19338,N_14784,N_12024);
and U19339 (N_19339,N_10342,N_13328);
nand U19340 (N_19340,N_10849,N_10740);
and U19341 (N_19341,N_11340,N_10940);
and U19342 (N_19342,N_12814,N_12759);
nand U19343 (N_19343,N_12156,N_12971);
xnor U19344 (N_19344,N_13404,N_10169);
or U19345 (N_19345,N_11801,N_13158);
or U19346 (N_19346,N_11027,N_10611);
nand U19347 (N_19347,N_12941,N_12128);
or U19348 (N_19348,N_10020,N_13218);
nor U19349 (N_19349,N_10211,N_11683);
or U19350 (N_19350,N_14818,N_13783);
and U19351 (N_19351,N_13231,N_14288);
nor U19352 (N_19352,N_14582,N_14792);
nor U19353 (N_19353,N_10648,N_13354);
nand U19354 (N_19354,N_13963,N_14226);
or U19355 (N_19355,N_14893,N_13525);
or U19356 (N_19356,N_14206,N_11123);
or U19357 (N_19357,N_12075,N_13273);
or U19358 (N_19358,N_14111,N_11781);
nor U19359 (N_19359,N_10042,N_12653);
nand U19360 (N_19360,N_11005,N_14559);
nand U19361 (N_19361,N_13217,N_11792);
or U19362 (N_19362,N_12330,N_14970);
nand U19363 (N_19363,N_13700,N_10854);
nor U19364 (N_19364,N_14184,N_14653);
nand U19365 (N_19365,N_12924,N_12071);
nand U19366 (N_19366,N_11351,N_12264);
or U19367 (N_19367,N_14739,N_13742);
and U19368 (N_19368,N_10764,N_11787);
nand U19369 (N_19369,N_10943,N_12546);
nor U19370 (N_19370,N_11529,N_12593);
nor U19371 (N_19371,N_12129,N_12970);
nand U19372 (N_19372,N_10351,N_10937);
nor U19373 (N_19373,N_13527,N_12296);
nand U19374 (N_19374,N_13148,N_13568);
nand U19375 (N_19375,N_11957,N_10814);
and U19376 (N_19376,N_11237,N_13256);
nand U19377 (N_19377,N_10131,N_12167);
or U19378 (N_19378,N_14383,N_12745);
or U19379 (N_19379,N_13972,N_13281);
or U19380 (N_19380,N_11236,N_14164);
nand U19381 (N_19381,N_13243,N_14196);
nor U19382 (N_19382,N_12341,N_12278);
or U19383 (N_19383,N_11043,N_13283);
or U19384 (N_19384,N_14657,N_14332);
or U19385 (N_19385,N_12022,N_14340);
nand U19386 (N_19386,N_14006,N_12232);
or U19387 (N_19387,N_13313,N_10525);
nand U19388 (N_19388,N_13731,N_12508);
nand U19389 (N_19389,N_12642,N_14684);
and U19390 (N_19390,N_14420,N_10361);
and U19391 (N_19391,N_14536,N_13564);
xnor U19392 (N_19392,N_12061,N_12041);
and U19393 (N_19393,N_11253,N_11419);
nand U19394 (N_19394,N_12425,N_13568);
nor U19395 (N_19395,N_12591,N_13687);
nor U19396 (N_19396,N_11819,N_14097);
xor U19397 (N_19397,N_14343,N_10959);
nor U19398 (N_19398,N_13585,N_13875);
nor U19399 (N_19399,N_12558,N_10333);
or U19400 (N_19400,N_11838,N_10805);
and U19401 (N_19401,N_10710,N_12671);
and U19402 (N_19402,N_13907,N_12711);
nor U19403 (N_19403,N_13125,N_10894);
nor U19404 (N_19404,N_14318,N_11470);
and U19405 (N_19405,N_14057,N_10409);
or U19406 (N_19406,N_13894,N_13413);
and U19407 (N_19407,N_11419,N_13438);
nor U19408 (N_19408,N_12139,N_13101);
nor U19409 (N_19409,N_10209,N_14184);
and U19410 (N_19410,N_14246,N_10379);
nor U19411 (N_19411,N_14986,N_14059);
and U19412 (N_19412,N_12718,N_10150);
or U19413 (N_19413,N_10550,N_10479);
and U19414 (N_19414,N_13598,N_12732);
or U19415 (N_19415,N_12005,N_11536);
or U19416 (N_19416,N_14232,N_13975);
and U19417 (N_19417,N_11099,N_10745);
and U19418 (N_19418,N_12645,N_12408);
nand U19419 (N_19419,N_13782,N_14241);
nand U19420 (N_19420,N_11682,N_12553);
nand U19421 (N_19421,N_10346,N_11292);
or U19422 (N_19422,N_12147,N_14302);
or U19423 (N_19423,N_10127,N_11194);
and U19424 (N_19424,N_14526,N_14363);
nand U19425 (N_19425,N_11882,N_10425);
nand U19426 (N_19426,N_10080,N_14180);
or U19427 (N_19427,N_12673,N_14051);
nand U19428 (N_19428,N_10917,N_13140);
or U19429 (N_19429,N_11156,N_13788);
nand U19430 (N_19430,N_12119,N_10376);
nor U19431 (N_19431,N_12529,N_12932);
or U19432 (N_19432,N_11734,N_14493);
nor U19433 (N_19433,N_11322,N_14217);
and U19434 (N_19434,N_14600,N_12518);
and U19435 (N_19435,N_13324,N_10895);
nor U19436 (N_19436,N_11736,N_12547);
or U19437 (N_19437,N_13535,N_11979);
nand U19438 (N_19438,N_14927,N_13183);
and U19439 (N_19439,N_14240,N_12883);
nor U19440 (N_19440,N_11415,N_14135);
and U19441 (N_19441,N_14946,N_13538);
and U19442 (N_19442,N_14022,N_11936);
and U19443 (N_19443,N_11350,N_10155);
nand U19444 (N_19444,N_11590,N_12331);
nor U19445 (N_19445,N_14038,N_14507);
and U19446 (N_19446,N_14594,N_14651);
or U19447 (N_19447,N_11773,N_12472);
nand U19448 (N_19448,N_11992,N_11362);
nand U19449 (N_19449,N_14858,N_14675);
nand U19450 (N_19450,N_13047,N_11463);
nand U19451 (N_19451,N_10070,N_14638);
and U19452 (N_19452,N_11523,N_12174);
nand U19453 (N_19453,N_11945,N_10024);
and U19454 (N_19454,N_14531,N_14051);
nand U19455 (N_19455,N_12583,N_12145);
and U19456 (N_19456,N_13535,N_11414);
nand U19457 (N_19457,N_11882,N_14039);
nor U19458 (N_19458,N_11102,N_11431);
nor U19459 (N_19459,N_14552,N_14914);
or U19460 (N_19460,N_11180,N_14934);
nand U19461 (N_19461,N_10661,N_10521);
nand U19462 (N_19462,N_14170,N_12886);
or U19463 (N_19463,N_12462,N_14881);
and U19464 (N_19464,N_11397,N_11761);
nand U19465 (N_19465,N_12897,N_14336);
nand U19466 (N_19466,N_12326,N_12149);
or U19467 (N_19467,N_10166,N_13330);
and U19468 (N_19468,N_12553,N_10081);
nand U19469 (N_19469,N_14469,N_14915);
nor U19470 (N_19470,N_13644,N_12740);
and U19471 (N_19471,N_11124,N_11767);
nor U19472 (N_19472,N_11541,N_13734);
nor U19473 (N_19473,N_11619,N_13081);
nand U19474 (N_19474,N_12987,N_11519);
and U19475 (N_19475,N_12610,N_14279);
nand U19476 (N_19476,N_12914,N_11317);
and U19477 (N_19477,N_14128,N_10212);
nor U19478 (N_19478,N_14390,N_10993);
and U19479 (N_19479,N_13743,N_14285);
nor U19480 (N_19480,N_12855,N_11994);
nand U19481 (N_19481,N_13560,N_14278);
or U19482 (N_19482,N_12422,N_10389);
nand U19483 (N_19483,N_11905,N_10524);
nand U19484 (N_19484,N_12994,N_11995);
nand U19485 (N_19485,N_10245,N_11580);
nor U19486 (N_19486,N_14824,N_12442);
nor U19487 (N_19487,N_10119,N_11797);
or U19488 (N_19488,N_10331,N_13358);
and U19489 (N_19489,N_13697,N_11369);
xor U19490 (N_19490,N_10027,N_14864);
and U19491 (N_19491,N_14992,N_12232);
nor U19492 (N_19492,N_12889,N_10865);
and U19493 (N_19493,N_14338,N_14155);
nand U19494 (N_19494,N_14849,N_12942);
or U19495 (N_19495,N_11869,N_10417);
or U19496 (N_19496,N_11696,N_13644);
and U19497 (N_19497,N_10571,N_13198);
or U19498 (N_19498,N_13999,N_10696);
xor U19499 (N_19499,N_12422,N_10009);
nand U19500 (N_19500,N_10983,N_11915);
and U19501 (N_19501,N_11016,N_11988);
or U19502 (N_19502,N_11722,N_11082);
nor U19503 (N_19503,N_10074,N_13782);
nand U19504 (N_19504,N_11956,N_10423);
or U19505 (N_19505,N_13993,N_11510);
xor U19506 (N_19506,N_11647,N_14608);
and U19507 (N_19507,N_10372,N_10725);
nand U19508 (N_19508,N_14522,N_13808);
nor U19509 (N_19509,N_11803,N_12654);
nor U19510 (N_19510,N_14831,N_12744);
nand U19511 (N_19511,N_11947,N_14225);
or U19512 (N_19512,N_10189,N_14567);
nor U19513 (N_19513,N_14394,N_13221);
nor U19514 (N_19514,N_13402,N_12233);
nor U19515 (N_19515,N_11479,N_11427);
or U19516 (N_19516,N_10817,N_10885);
or U19517 (N_19517,N_10350,N_14924);
nor U19518 (N_19518,N_12473,N_11443);
xnor U19519 (N_19519,N_13860,N_12724);
or U19520 (N_19520,N_11055,N_10842);
nor U19521 (N_19521,N_14648,N_14431);
and U19522 (N_19522,N_11647,N_11053);
nand U19523 (N_19523,N_11877,N_11739);
nand U19524 (N_19524,N_11703,N_13801);
or U19525 (N_19525,N_12552,N_12132);
nand U19526 (N_19526,N_13121,N_12300);
or U19527 (N_19527,N_14885,N_13218);
nor U19528 (N_19528,N_14295,N_13575);
nand U19529 (N_19529,N_10322,N_13093);
and U19530 (N_19530,N_10477,N_13217);
nor U19531 (N_19531,N_10153,N_12977);
or U19532 (N_19532,N_14275,N_13212);
or U19533 (N_19533,N_11509,N_12880);
and U19534 (N_19534,N_12807,N_13965);
or U19535 (N_19535,N_13732,N_10649);
nand U19536 (N_19536,N_14206,N_10112);
nand U19537 (N_19537,N_11728,N_13606);
nand U19538 (N_19538,N_13754,N_12268);
nand U19539 (N_19539,N_14907,N_14400);
nand U19540 (N_19540,N_13067,N_10993);
nor U19541 (N_19541,N_10862,N_11634);
and U19542 (N_19542,N_10954,N_10816);
nand U19543 (N_19543,N_11191,N_12889);
nor U19544 (N_19544,N_13534,N_13924);
nor U19545 (N_19545,N_11390,N_14577);
nand U19546 (N_19546,N_13812,N_13167);
or U19547 (N_19547,N_11111,N_11567);
or U19548 (N_19548,N_13766,N_11325);
or U19549 (N_19549,N_14693,N_13420);
or U19550 (N_19550,N_13044,N_12381);
and U19551 (N_19551,N_10289,N_14522);
nor U19552 (N_19552,N_11108,N_10120);
nand U19553 (N_19553,N_13548,N_14581);
and U19554 (N_19554,N_14139,N_11007);
and U19555 (N_19555,N_13150,N_10555);
nor U19556 (N_19556,N_12239,N_10726);
or U19557 (N_19557,N_11977,N_10409);
and U19558 (N_19558,N_10428,N_12065);
nand U19559 (N_19559,N_12260,N_10975);
or U19560 (N_19560,N_10941,N_12204);
nand U19561 (N_19561,N_14715,N_12033);
nor U19562 (N_19562,N_12620,N_11233);
or U19563 (N_19563,N_14107,N_13183);
nand U19564 (N_19564,N_10501,N_10745);
and U19565 (N_19565,N_14679,N_14699);
nand U19566 (N_19566,N_14879,N_10373);
nor U19567 (N_19567,N_10287,N_14033);
or U19568 (N_19568,N_11819,N_13202);
nor U19569 (N_19569,N_11631,N_14655);
and U19570 (N_19570,N_11940,N_10210);
and U19571 (N_19571,N_12748,N_12876);
nor U19572 (N_19572,N_13743,N_12938);
nor U19573 (N_19573,N_13635,N_10595);
nor U19574 (N_19574,N_14256,N_11815);
nor U19575 (N_19575,N_13803,N_10795);
and U19576 (N_19576,N_12616,N_14203);
or U19577 (N_19577,N_11024,N_11261);
and U19578 (N_19578,N_13745,N_14273);
nand U19579 (N_19579,N_10250,N_12032);
or U19580 (N_19580,N_14271,N_10698);
or U19581 (N_19581,N_12636,N_10860);
nor U19582 (N_19582,N_11754,N_12835);
nand U19583 (N_19583,N_11939,N_12630);
or U19584 (N_19584,N_13927,N_13591);
and U19585 (N_19585,N_10870,N_12651);
nand U19586 (N_19586,N_11934,N_13468);
or U19587 (N_19587,N_11281,N_13164);
and U19588 (N_19588,N_14934,N_11603);
nor U19589 (N_19589,N_13618,N_13093);
or U19590 (N_19590,N_10800,N_10802);
and U19591 (N_19591,N_12654,N_10727);
nand U19592 (N_19592,N_10321,N_13835);
and U19593 (N_19593,N_13495,N_12689);
nor U19594 (N_19594,N_13177,N_12650);
nor U19595 (N_19595,N_11670,N_10064);
and U19596 (N_19596,N_11628,N_10494);
nor U19597 (N_19597,N_12393,N_12637);
and U19598 (N_19598,N_10637,N_10655);
and U19599 (N_19599,N_14667,N_12779);
nand U19600 (N_19600,N_10738,N_14174);
or U19601 (N_19601,N_13960,N_14714);
and U19602 (N_19602,N_11601,N_10134);
or U19603 (N_19603,N_10406,N_13279);
and U19604 (N_19604,N_11364,N_10060);
nor U19605 (N_19605,N_13551,N_13404);
nand U19606 (N_19606,N_13504,N_11286);
and U19607 (N_19607,N_11522,N_13491);
nand U19608 (N_19608,N_11198,N_12785);
nor U19609 (N_19609,N_14777,N_13045);
and U19610 (N_19610,N_13248,N_12120);
or U19611 (N_19611,N_11582,N_13850);
nand U19612 (N_19612,N_13507,N_13157);
nor U19613 (N_19613,N_10719,N_14925);
and U19614 (N_19614,N_13736,N_14422);
xnor U19615 (N_19615,N_13758,N_13493);
or U19616 (N_19616,N_12593,N_11841);
or U19617 (N_19617,N_14737,N_10144);
nand U19618 (N_19618,N_12453,N_12264);
and U19619 (N_19619,N_14740,N_11614);
or U19620 (N_19620,N_13662,N_13297);
and U19621 (N_19621,N_10344,N_10220);
and U19622 (N_19622,N_11279,N_14418);
nand U19623 (N_19623,N_10184,N_11268);
nand U19624 (N_19624,N_13788,N_12257);
or U19625 (N_19625,N_10888,N_14773);
nand U19626 (N_19626,N_14143,N_14390);
nor U19627 (N_19627,N_10402,N_12184);
nor U19628 (N_19628,N_14563,N_14887);
nand U19629 (N_19629,N_13860,N_10031);
nand U19630 (N_19630,N_11610,N_10022);
nor U19631 (N_19631,N_10935,N_13313);
and U19632 (N_19632,N_12278,N_12143);
nor U19633 (N_19633,N_14989,N_12879);
nand U19634 (N_19634,N_12095,N_11216);
or U19635 (N_19635,N_10734,N_10370);
or U19636 (N_19636,N_14927,N_14477);
nand U19637 (N_19637,N_12627,N_13194);
or U19638 (N_19638,N_14049,N_10088);
nor U19639 (N_19639,N_11723,N_14562);
or U19640 (N_19640,N_14840,N_13898);
or U19641 (N_19641,N_11550,N_11357);
or U19642 (N_19642,N_11354,N_14269);
nand U19643 (N_19643,N_14898,N_12443);
nand U19644 (N_19644,N_10933,N_10291);
nand U19645 (N_19645,N_12650,N_13784);
nand U19646 (N_19646,N_12822,N_14895);
nor U19647 (N_19647,N_10101,N_12418);
nand U19648 (N_19648,N_10052,N_10004);
nor U19649 (N_19649,N_14347,N_10794);
and U19650 (N_19650,N_14931,N_14783);
nand U19651 (N_19651,N_12618,N_11015);
nor U19652 (N_19652,N_11813,N_14376);
or U19653 (N_19653,N_13041,N_11940);
nor U19654 (N_19654,N_11777,N_14739);
nand U19655 (N_19655,N_12692,N_10633);
nor U19656 (N_19656,N_12079,N_10664);
and U19657 (N_19657,N_12467,N_11736);
or U19658 (N_19658,N_10155,N_13849);
nand U19659 (N_19659,N_12422,N_13992);
and U19660 (N_19660,N_13087,N_10849);
nor U19661 (N_19661,N_11662,N_11623);
nand U19662 (N_19662,N_10213,N_13136);
or U19663 (N_19663,N_13017,N_11909);
or U19664 (N_19664,N_14446,N_12934);
or U19665 (N_19665,N_13636,N_13859);
nor U19666 (N_19666,N_10156,N_13361);
or U19667 (N_19667,N_14031,N_14766);
nand U19668 (N_19668,N_10302,N_14321);
nor U19669 (N_19669,N_10708,N_11181);
nor U19670 (N_19670,N_10839,N_10062);
or U19671 (N_19671,N_14097,N_12570);
nor U19672 (N_19672,N_11977,N_11258);
or U19673 (N_19673,N_10370,N_11452);
nand U19674 (N_19674,N_11247,N_11144);
or U19675 (N_19675,N_11804,N_14168);
nand U19676 (N_19676,N_14773,N_13912);
nand U19677 (N_19677,N_10875,N_13259);
and U19678 (N_19678,N_12181,N_12868);
nand U19679 (N_19679,N_12446,N_10680);
nor U19680 (N_19680,N_14750,N_10997);
nand U19681 (N_19681,N_12238,N_10548);
nor U19682 (N_19682,N_11319,N_10173);
and U19683 (N_19683,N_11698,N_13765);
nor U19684 (N_19684,N_14367,N_12565);
or U19685 (N_19685,N_10491,N_11709);
and U19686 (N_19686,N_14667,N_14477);
nand U19687 (N_19687,N_13763,N_13969);
nor U19688 (N_19688,N_10926,N_11777);
or U19689 (N_19689,N_10622,N_11590);
and U19690 (N_19690,N_10713,N_11960);
and U19691 (N_19691,N_11464,N_10612);
nor U19692 (N_19692,N_10495,N_11339);
and U19693 (N_19693,N_10573,N_14146);
or U19694 (N_19694,N_13659,N_13435);
nand U19695 (N_19695,N_13949,N_13573);
or U19696 (N_19696,N_14970,N_12431);
nor U19697 (N_19697,N_12883,N_13816);
nor U19698 (N_19698,N_11296,N_12994);
and U19699 (N_19699,N_13389,N_13262);
or U19700 (N_19700,N_11243,N_12845);
nand U19701 (N_19701,N_10918,N_13572);
xnor U19702 (N_19702,N_10140,N_12999);
and U19703 (N_19703,N_12063,N_12727);
or U19704 (N_19704,N_10224,N_12152);
nor U19705 (N_19705,N_11428,N_14802);
and U19706 (N_19706,N_13907,N_12897);
and U19707 (N_19707,N_13289,N_14769);
nor U19708 (N_19708,N_14657,N_10489);
and U19709 (N_19709,N_11104,N_11681);
and U19710 (N_19710,N_10706,N_14612);
nand U19711 (N_19711,N_11239,N_12834);
nor U19712 (N_19712,N_10946,N_10911);
xor U19713 (N_19713,N_14628,N_11513);
nor U19714 (N_19714,N_11421,N_11885);
nor U19715 (N_19715,N_11208,N_13065);
nor U19716 (N_19716,N_12181,N_10179);
or U19717 (N_19717,N_13215,N_14621);
and U19718 (N_19718,N_12512,N_14683);
nand U19719 (N_19719,N_10485,N_10640);
and U19720 (N_19720,N_12473,N_13132);
nor U19721 (N_19721,N_14008,N_11878);
nor U19722 (N_19722,N_13188,N_12910);
and U19723 (N_19723,N_11660,N_13259);
or U19724 (N_19724,N_14819,N_13656);
nand U19725 (N_19725,N_10238,N_11191);
nand U19726 (N_19726,N_12539,N_14593);
or U19727 (N_19727,N_13426,N_10099);
xor U19728 (N_19728,N_11231,N_10821);
or U19729 (N_19729,N_13115,N_14726);
or U19730 (N_19730,N_14773,N_13609);
nor U19731 (N_19731,N_13410,N_10881);
and U19732 (N_19732,N_11736,N_13297);
and U19733 (N_19733,N_12433,N_12520);
and U19734 (N_19734,N_10279,N_14546);
xor U19735 (N_19735,N_11595,N_13005);
or U19736 (N_19736,N_12878,N_14801);
xor U19737 (N_19737,N_11405,N_10493);
nor U19738 (N_19738,N_10311,N_10505);
nor U19739 (N_19739,N_14623,N_10968);
and U19740 (N_19740,N_10188,N_10982);
nor U19741 (N_19741,N_14960,N_12358);
nor U19742 (N_19742,N_13186,N_10755);
nand U19743 (N_19743,N_14009,N_12655);
nand U19744 (N_19744,N_11073,N_10662);
and U19745 (N_19745,N_11881,N_12688);
and U19746 (N_19746,N_13684,N_12969);
nand U19747 (N_19747,N_12420,N_10751);
nor U19748 (N_19748,N_11276,N_11520);
xor U19749 (N_19749,N_13552,N_10909);
and U19750 (N_19750,N_11047,N_12351);
xnor U19751 (N_19751,N_11754,N_14829);
or U19752 (N_19752,N_12893,N_13731);
nand U19753 (N_19753,N_11351,N_12342);
nand U19754 (N_19754,N_13605,N_14420);
nand U19755 (N_19755,N_11708,N_10018);
or U19756 (N_19756,N_14166,N_11062);
nand U19757 (N_19757,N_12953,N_14042);
and U19758 (N_19758,N_13258,N_11879);
or U19759 (N_19759,N_12144,N_10733);
nand U19760 (N_19760,N_13032,N_12752);
nand U19761 (N_19761,N_14450,N_13870);
nor U19762 (N_19762,N_14765,N_14982);
xnor U19763 (N_19763,N_13740,N_13714);
nor U19764 (N_19764,N_13919,N_14442);
or U19765 (N_19765,N_10385,N_13857);
nor U19766 (N_19766,N_14319,N_11501);
nand U19767 (N_19767,N_12554,N_11661);
and U19768 (N_19768,N_11614,N_10271);
and U19769 (N_19769,N_11970,N_13214);
and U19770 (N_19770,N_10917,N_11664);
nor U19771 (N_19771,N_12726,N_13356);
nor U19772 (N_19772,N_11495,N_13814);
nor U19773 (N_19773,N_11035,N_12116);
and U19774 (N_19774,N_13198,N_13420);
and U19775 (N_19775,N_10715,N_14448);
or U19776 (N_19776,N_13525,N_13922);
nand U19777 (N_19777,N_10106,N_11081);
and U19778 (N_19778,N_10551,N_11283);
xnor U19779 (N_19779,N_12244,N_10644);
nor U19780 (N_19780,N_14352,N_13777);
nor U19781 (N_19781,N_14936,N_14961);
nand U19782 (N_19782,N_10552,N_11128);
or U19783 (N_19783,N_11675,N_13572);
nor U19784 (N_19784,N_10461,N_14979);
and U19785 (N_19785,N_11751,N_14711);
nor U19786 (N_19786,N_11806,N_10264);
nand U19787 (N_19787,N_12689,N_13372);
nor U19788 (N_19788,N_11170,N_10731);
nor U19789 (N_19789,N_11485,N_12415);
or U19790 (N_19790,N_13200,N_14283);
nor U19791 (N_19791,N_10723,N_13262);
or U19792 (N_19792,N_14820,N_12703);
nor U19793 (N_19793,N_11882,N_14392);
nor U19794 (N_19794,N_13607,N_13385);
or U19795 (N_19795,N_13431,N_13583);
and U19796 (N_19796,N_10892,N_11952);
nor U19797 (N_19797,N_11311,N_13323);
or U19798 (N_19798,N_12731,N_14095);
nor U19799 (N_19799,N_13240,N_12375);
nand U19800 (N_19800,N_11819,N_10775);
nor U19801 (N_19801,N_12914,N_10886);
nor U19802 (N_19802,N_14638,N_11770);
nor U19803 (N_19803,N_12824,N_14598);
xnor U19804 (N_19804,N_10910,N_12150);
or U19805 (N_19805,N_13584,N_13881);
nand U19806 (N_19806,N_13100,N_13014);
nand U19807 (N_19807,N_12768,N_10855);
and U19808 (N_19808,N_11759,N_11435);
nand U19809 (N_19809,N_12313,N_10275);
or U19810 (N_19810,N_10473,N_13655);
nand U19811 (N_19811,N_11292,N_11119);
nand U19812 (N_19812,N_14950,N_14220);
nor U19813 (N_19813,N_11315,N_14144);
or U19814 (N_19814,N_13469,N_12633);
and U19815 (N_19815,N_13058,N_10261);
or U19816 (N_19816,N_11021,N_14782);
xnor U19817 (N_19817,N_10059,N_12672);
and U19818 (N_19818,N_10276,N_11063);
or U19819 (N_19819,N_11426,N_11676);
nor U19820 (N_19820,N_12931,N_13866);
or U19821 (N_19821,N_10085,N_11713);
nor U19822 (N_19822,N_11747,N_11164);
xor U19823 (N_19823,N_11886,N_14916);
nor U19824 (N_19824,N_11030,N_10389);
and U19825 (N_19825,N_10756,N_10328);
nand U19826 (N_19826,N_12557,N_13913);
or U19827 (N_19827,N_11723,N_14684);
nand U19828 (N_19828,N_13759,N_10517);
nand U19829 (N_19829,N_12020,N_12796);
or U19830 (N_19830,N_12385,N_13988);
or U19831 (N_19831,N_12933,N_11722);
nor U19832 (N_19832,N_13002,N_11315);
and U19833 (N_19833,N_13588,N_14000);
nor U19834 (N_19834,N_12299,N_11238);
and U19835 (N_19835,N_10880,N_10871);
or U19836 (N_19836,N_11860,N_10846);
and U19837 (N_19837,N_14163,N_10318);
or U19838 (N_19838,N_14036,N_11593);
and U19839 (N_19839,N_12006,N_13358);
nand U19840 (N_19840,N_11407,N_14024);
and U19841 (N_19841,N_10710,N_12817);
nor U19842 (N_19842,N_11566,N_10249);
and U19843 (N_19843,N_14506,N_10795);
nand U19844 (N_19844,N_10231,N_12155);
and U19845 (N_19845,N_13493,N_11856);
nand U19846 (N_19846,N_10809,N_14000);
nor U19847 (N_19847,N_11172,N_14672);
or U19848 (N_19848,N_13715,N_12001);
or U19849 (N_19849,N_14866,N_13153);
or U19850 (N_19850,N_10194,N_11675);
or U19851 (N_19851,N_11902,N_13335);
and U19852 (N_19852,N_12840,N_13771);
and U19853 (N_19853,N_13344,N_12750);
or U19854 (N_19854,N_11379,N_11068);
or U19855 (N_19855,N_14460,N_11241);
nor U19856 (N_19856,N_11616,N_11855);
and U19857 (N_19857,N_12762,N_12289);
and U19858 (N_19858,N_13012,N_10132);
nand U19859 (N_19859,N_13365,N_11096);
and U19860 (N_19860,N_13333,N_12905);
and U19861 (N_19861,N_13794,N_12495);
and U19862 (N_19862,N_13848,N_14322);
or U19863 (N_19863,N_12163,N_10103);
nor U19864 (N_19864,N_11942,N_14344);
or U19865 (N_19865,N_10748,N_13917);
or U19866 (N_19866,N_13484,N_13799);
nand U19867 (N_19867,N_13602,N_10736);
or U19868 (N_19868,N_11869,N_13119);
and U19869 (N_19869,N_14454,N_14811);
nand U19870 (N_19870,N_11364,N_12886);
or U19871 (N_19871,N_12511,N_12694);
or U19872 (N_19872,N_14933,N_11904);
nand U19873 (N_19873,N_14635,N_11768);
or U19874 (N_19874,N_10300,N_10742);
nor U19875 (N_19875,N_12044,N_12114);
and U19876 (N_19876,N_13708,N_11833);
nor U19877 (N_19877,N_10748,N_14882);
and U19878 (N_19878,N_12650,N_10627);
and U19879 (N_19879,N_12697,N_14597);
nand U19880 (N_19880,N_13197,N_11575);
nor U19881 (N_19881,N_13248,N_13113);
nor U19882 (N_19882,N_13063,N_12405);
and U19883 (N_19883,N_13463,N_14213);
or U19884 (N_19884,N_11076,N_11133);
or U19885 (N_19885,N_13271,N_12499);
nor U19886 (N_19886,N_13993,N_10601);
or U19887 (N_19887,N_10620,N_10475);
nand U19888 (N_19888,N_10888,N_14730);
nor U19889 (N_19889,N_11404,N_11326);
or U19890 (N_19890,N_11811,N_14154);
xnor U19891 (N_19891,N_13102,N_14550);
and U19892 (N_19892,N_12391,N_11265);
or U19893 (N_19893,N_14106,N_12128);
nor U19894 (N_19894,N_11040,N_10146);
nand U19895 (N_19895,N_13957,N_14742);
and U19896 (N_19896,N_10592,N_11960);
and U19897 (N_19897,N_14052,N_11660);
or U19898 (N_19898,N_12038,N_14828);
nand U19899 (N_19899,N_14291,N_11566);
or U19900 (N_19900,N_10789,N_10254);
and U19901 (N_19901,N_11339,N_13461);
nand U19902 (N_19902,N_13039,N_10555);
nor U19903 (N_19903,N_10807,N_11455);
and U19904 (N_19904,N_14756,N_14401);
and U19905 (N_19905,N_14057,N_10377);
nand U19906 (N_19906,N_14579,N_12398);
nand U19907 (N_19907,N_12708,N_12641);
and U19908 (N_19908,N_11006,N_14289);
and U19909 (N_19909,N_12955,N_10287);
or U19910 (N_19910,N_10652,N_14954);
nor U19911 (N_19911,N_11216,N_10554);
or U19912 (N_19912,N_11654,N_14637);
and U19913 (N_19913,N_13343,N_13563);
or U19914 (N_19914,N_10509,N_13756);
and U19915 (N_19915,N_11860,N_14586);
and U19916 (N_19916,N_13008,N_10187);
nand U19917 (N_19917,N_11608,N_14349);
nor U19918 (N_19918,N_11852,N_13397);
nand U19919 (N_19919,N_14327,N_13097);
xnor U19920 (N_19920,N_13198,N_13201);
and U19921 (N_19921,N_10182,N_12076);
nand U19922 (N_19922,N_13697,N_13135);
and U19923 (N_19923,N_10514,N_11538);
and U19924 (N_19924,N_11377,N_13989);
nand U19925 (N_19925,N_10096,N_12449);
nand U19926 (N_19926,N_14648,N_12060);
or U19927 (N_19927,N_12021,N_10533);
and U19928 (N_19928,N_13401,N_11116);
nand U19929 (N_19929,N_13111,N_12515);
nor U19930 (N_19930,N_13562,N_13097);
nand U19931 (N_19931,N_10615,N_11932);
nand U19932 (N_19932,N_14751,N_13768);
and U19933 (N_19933,N_12774,N_11776);
and U19934 (N_19934,N_10856,N_10557);
nand U19935 (N_19935,N_14408,N_11566);
nand U19936 (N_19936,N_14998,N_11754);
and U19937 (N_19937,N_11293,N_12753);
nand U19938 (N_19938,N_13937,N_13089);
and U19939 (N_19939,N_10111,N_10636);
nand U19940 (N_19940,N_14222,N_11686);
or U19941 (N_19941,N_11724,N_13008);
and U19942 (N_19942,N_12802,N_13792);
nand U19943 (N_19943,N_14360,N_14765);
nor U19944 (N_19944,N_10009,N_13189);
or U19945 (N_19945,N_10939,N_12336);
or U19946 (N_19946,N_12524,N_13615);
nand U19947 (N_19947,N_11140,N_14056);
and U19948 (N_19948,N_14010,N_12384);
nand U19949 (N_19949,N_10606,N_11901);
nor U19950 (N_19950,N_10154,N_14634);
nand U19951 (N_19951,N_10479,N_12290);
and U19952 (N_19952,N_13425,N_10820);
nand U19953 (N_19953,N_14192,N_13141);
or U19954 (N_19954,N_11226,N_10197);
nor U19955 (N_19955,N_11645,N_10123);
or U19956 (N_19956,N_10704,N_11882);
and U19957 (N_19957,N_11084,N_14872);
and U19958 (N_19958,N_10264,N_10739);
nand U19959 (N_19959,N_11244,N_10521);
nand U19960 (N_19960,N_14305,N_13030);
nor U19961 (N_19961,N_10253,N_13438);
or U19962 (N_19962,N_10647,N_13913);
nand U19963 (N_19963,N_14606,N_12756);
nor U19964 (N_19964,N_11451,N_13410);
nor U19965 (N_19965,N_10275,N_12535);
or U19966 (N_19966,N_12374,N_12497);
or U19967 (N_19967,N_13946,N_13970);
nor U19968 (N_19968,N_10034,N_11501);
nor U19969 (N_19969,N_14338,N_14069);
and U19970 (N_19970,N_10162,N_13190);
nand U19971 (N_19971,N_11029,N_14845);
nand U19972 (N_19972,N_13082,N_11950);
and U19973 (N_19973,N_12299,N_13692);
nand U19974 (N_19974,N_10705,N_13436);
and U19975 (N_19975,N_10861,N_12476);
nand U19976 (N_19976,N_14957,N_13538);
or U19977 (N_19977,N_11118,N_10726);
nand U19978 (N_19978,N_14657,N_10348);
and U19979 (N_19979,N_14096,N_10088);
nor U19980 (N_19980,N_12416,N_10232);
nor U19981 (N_19981,N_13394,N_12133);
and U19982 (N_19982,N_14109,N_10468);
or U19983 (N_19983,N_11876,N_12520);
and U19984 (N_19984,N_13968,N_10830);
or U19985 (N_19985,N_11412,N_11729);
or U19986 (N_19986,N_10263,N_11458);
nand U19987 (N_19987,N_14271,N_13502);
nor U19988 (N_19988,N_10281,N_12643);
xor U19989 (N_19989,N_13870,N_10754);
and U19990 (N_19990,N_14030,N_13054);
nor U19991 (N_19991,N_13798,N_12802);
nand U19992 (N_19992,N_11784,N_10326);
nand U19993 (N_19993,N_14432,N_11541);
or U19994 (N_19994,N_14889,N_10520);
or U19995 (N_19995,N_14186,N_11819);
nor U19996 (N_19996,N_11700,N_10753);
or U19997 (N_19997,N_13503,N_12174);
and U19998 (N_19998,N_10005,N_14515);
nand U19999 (N_19999,N_10504,N_14088);
nand U20000 (N_20000,N_15007,N_17423);
nand U20001 (N_20001,N_15544,N_16754);
xor U20002 (N_20002,N_19995,N_18018);
or U20003 (N_20003,N_19207,N_16158);
and U20004 (N_20004,N_19453,N_18916);
nor U20005 (N_20005,N_15966,N_15304);
nand U20006 (N_20006,N_19872,N_19214);
nand U20007 (N_20007,N_15367,N_18017);
nor U20008 (N_20008,N_15332,N_19085);
nor U20009 (N_20009,N_15254,N_16163);
or U20010 (N_20010,N_15798,N_17433);
nand U20011 (N_20011,N_18592,N_15112);
and U20012 (N_20012,N_16977,N_19646);
nor U20013 (N_20013,N_19736,N_15842);
nor U20014 (N_20014,N_19640,N_17513);
nand U20015 (N_20015,N_16644,N_17012);
and U20016 (N_20016,N_16277,N_16054);
nor U20017 (N_20017,N_16190,N_15527);
xor U20018 (N_20018,N_18545,N_18232);
or U20019 (N_20019,N_15503,N_17021);
and U20020 (N_20020,N_17326,N_15376);
nor U20021 (N_20021,N_16021,N_15105);
nor U20022 (N_20022,N_18346,N_18779);
nand U20023 (N_20023,N_18289,N_19755);
or U20024 (N_20024,N_15999,N_17372);
nor U20025 (N_20025,N_16883,N_16155);
and U20026 (N_20026,N_17610,N_18104);
or U20027 (N_20027,N_15433,N_19092);
and U20028 (N_20028,N_17307,N_17358);
or U20029 (N_20029,N_18848,N_16249);
or U20030 (N_20030,N_17774,N_18627);
nor U20031 (N_20031,N_17560,N_15997);
and U20032 (N_20032,N_15971,N_18874);
nor U20033 (N_20033,N_16999,N_15557);
nand U20034 (N_20034,N_16445,N_18756);
and U20035 (N_20035,N_18934,N_18682);
and U20036 (N_20036,N_17547,N_16306);
or U20037 (N_20037,N_15745,N_18641);
and U20038 (N_20038,N_19395,N_16814);
and U20039 (N_20039,N_17179,N_19933);
nand U20040 (N_20040,N_18768,N_16447);
nor U20041 (N_20041,N_16459,N_18458);
nor U20042 (N_20042,N_16211,N_17244);
nand U20043 (N_20043,N_15601,N_19303);
nand U20044 (N_20044,N_15813,N_15988);
nand U20045 (N_20045,N_17435,N_16386);
nand U20046 (N_20046,N_19376,N_19131);
and U20047 (N_20047,N_19823,N_15872);
nand U20048 (N_20048,N_16052,N_15531);
xnor U20049 (N_20049,N_19289,N_16144);
or U20050 (N_20050,N_16038,N_16889);
or U20051 (N_20051,N_17988,N_17576);
and U20052 (N_20052,N_17355,N_16597);
nor U20053 (N_20053,N_15055,N_15486);
or U20054 (N_20054,N_17837,N_18199);
or U20055 (N_20055,N_16598,N_15054);
or U20056 (N_20056,N_17336,N_19913);
nand U20057 (N_20057,N_19259,N_16474);
nor U20058 (N_20058,N_16684,N_15663);
nand U20059 (N_20059,N_19546,N_15672);
or U20060 (N_20060,N_15518,N_16851);
nor U20061 (N_20061,N_16116,N_18800);
and U20062 (N_20062,N_19048,N_18067);
and U20063 (N_20063,N_15692,N_19989);
nand U20064 (N_20064,N_18659,N_17063);
and U20065 (N_20065,N_19330,N_15668);
and U20066 (N_20066,N_17084,N_16040);
nand U20067 (N_20067,N_18028,N_18580);
nor U20068 (N_20068,N_16000,N_17432);
nor U20069 (N_20069,N_19648,N_15599);
or U20070 (N_20070,N_15019,N_17263);
nor U20071 (N_20071,N_16241,N_16724);
nor U20072 (N_20072,N_19469,N_15691);
nor U20073 (N_20073,N_16162,N_16132);
nand U20074 (N_20074,N_15270,N_18147);
nor U20075 (N_20075,N_17691,N_16149);
and U20076 (N_20076,N_16252,N_18698);
or U20077 (N_20077,N_17896,N_16645);
and U20078 (N_20078,N_18224,N_18843);
nor U20079 (N_20079,N_15982,N_16524);
nand U20080 (N_20080,N_19084,N_19237);
and U20081 (N_20081,N_18142,N_17217);
or U20082 (N_20082,N_17274,N_18498);
nand U20083 (N_20083,N_15409,N_17945);
nand U20084 (N_20084,N_15155,N_19815);
nand U20085 (N_20085,N_19532,N_17071);
nand U20086 (N_20086,N_17738,N_17474);
and U20087 (N_20087,N_17016,N_17471);
nor U20088 (N_20088,N_18574,N_19548);
and U20089 (N_20089,N_17374,N_17710);
nand U20090 (N_20090,N_17283,N_18528);
and U20091 (N_20091,N_18382,N_18593);
nand U20092 (N_20092,N_15983,N_18890);
nand U20093 (N_20093,N_19619,N_16228);
nand U20094 (N_20094,N_15522,N_16746);
nor U20095 (N_20095,N_15126,N_19592);
nor U20096 (N_20096,N_19809,N_18949);
or U20097 (N_20097,N_19526,N_17612);
nand U20098 (N_20098,N_16551,N_17462);
nor U20099 (N_20099,N_16657,N_17754);
nor U20100 (N_20100,N_15578,N_16946);
or U20101 (N_20101,N_17431,N_19580);
nand U20102 (N_20102,N_17556,N_19360);
or U20103 (N_20103,N_19263,N_19482);
nand U20104 (N_20104,N_17644,N_15925);
nand U20105 (N_20105,N_18968,N_17871);
and U20106 (N_20106,N_16152,N_16947);
or U20107 (N_20107,N_15725,N_16579);
or U20108 (N_20108,N_15284,N_15477);
and U20109 (N_20109,N_15080,N_16559);
or U20110 (N_20110,N_16067,N_15896);
and U20111 (N_20111,N_18096,N_17128);
and U20112 (N_20112,N_17598,N_18970);
nand U20113 (N_20113,N_19002,N_16505);
and U20114 (N_20114,N_15905,N_16010);
nor U20115 (N_20115,N_15754,N_17378);
or U20116 (N_20116,N_17704,N_19921);
and U20117 (N_20117,N_18564,N_19910);
xnor U20118 (N_20118,N_15528,N_19795);
and U20119 (N_20119,N_17543,N_15504);
nor U20120 (N_20120,N_17282,N_19404);
nand U20121 (N_20121,N_19448,N_15891);
or U20122 (N_20122,N_17999,N_16079);
xor U20123 (N_20123,N_19027,N_17497);
nor U20124 (N_20124,N_19599,N_19598);
xor U20125 (N_20125,N_17745,N_15078);
nor U20126 (N_20126,N_18470,N_15776);
nand U20127 (N_20127,N_19649,N_19043);
and U20128 (N_20128,N_16929,N_16206);
nor U20129 (N_20129,N_15481,N_19536);
or U20130 (N_20130,N_18584,N_16385);
nor U20131 (N_20131,N_18771,N_16357);
nor U20132 (N_20132,N_17522,N_16689);
nand U20133 (N_20133,N_17763,N_18048);
and U20134 (N_20134,N_15136,N_16775);
or U20135 (N_20135,N_19262,N_18110);
nor U20136 (N_20136,N_18332,N_15073);
or U20137 (N_20137,N_18190,N_16519);
and U20138 (N_20138,N_15196,N_15303);
nor U20139 (N_20139,N_17105,N_19265);
nor U20140 (N_20140,N_16265,N_17510);
nand U20141 (N_20141,N_15897,N_18141);
and U20142 (N_20142,N_18500,N_15742);
or U20143 (N_20143,N_18654,N_18098);
and U20144 (N_20144,N_17491,N_15764);
or U20145 (N_20145,N_19126,N_15492);
nor U20146 (N_20146,N_15717,N_17359);
nor U20147 (N_20147,N_15931,N_19747);
and U20148 (N_20148,N_19839,N_15084);
or U20149 (N_20149,N_17487,N_19614);
and U20150 (N_20150,N_16708,N_16203);
nor U20151 (N_20151,N_15551,N_19275);
or U20152 (N_20152,N_19993,N_16778);
and U20153 (N_20153,N_17311,N_18724);
and U20154 (N_20154,N_17696,N_18219);
nor U20155 (N_20155,N_16840,N_16284);
nand U20156 (N_20156,N_17042,N_16870);
nand U20157 (N_20157,N_17113,N_15107);
or U20158 (N_20158,N_19515,N_18857);
nor U20159 (N_20159,N_15350,N_18745);
and U20160 (N_20160,N_19877,N_17571);
or U20161 (N_20161,N_18414,N_18058);
nor U20162 (N_20162,N_19684,N_18272);
or U20163 (N_20163,N_16272,N_18230);
and U20164 (N_20164,N_15986,N_18073);
nor U20165 (N_20165,N_17175,N_17818);
nand U20166 (N_20166,N_19762,N_16658);
nand U20167 (N_20167,N_16329,N_15859);
and U20168 (N_20168,N_18364,N_17149);
or U20169 (N_20169,N_15626,N_16570);
nand U20170 (N_20170,N_16630,N_17390);
nand U20171 (N_20171,N_16457,N_18555);
and U20172 (N_20172,N_18841,N_16412);
nor U20173 (N_20173,N_16012,N_18533);
nor U20174 (N_20174,N_15427,N_18467);
and U20175 (N_20175,N_15684,N_15398);
and U20176 (N_20176,N_18097,N_18312);
nand U20177 (N_20177,N_15563,N_18475);
nor U20178 (N_20178,N_18892,N_17756);
or U20179 (N_20179,N_17044,N_16450);
or U20180 (N_20180,N_17317,N_17156);
nand U20181 (N_20181,N_17421,N_16339);
nand U20182 (N_20182,N_18180,N_15980);
and U20183 (N_20183,N_15787,N_15086);
and U20184 (N_20184,N_19600,N_15840);
and U20185 (N_20185,N_18981,N_15232);
nand U20186 (N_20186,N_18819,N_17451);
or U20187 (N_20187,N_19887,N_17511);
nand U20188 (N_20188,N_19590,N_19644);
or U20189 (N_20189,N_17564,N_19885);
or U20190 (N_20190,N_15043,N_15830);
nand U20191 (N_20191,N_18342,N_15794);
nor U20192 (N_20192,N_19555,N_17979);
or U20193 (N_20193,N_15883,N_17797);
nand U20194 (N_20194,N_18294,N_19777);
or U20195 (N_20195,N_16654,N_19452);
nand U20196 (N_20196,N_16709,N_16777);
nor U20197 (N_20197,N_16632,N_16990);
nor U20198 (N_20198,N_17893,N_17253);
nand U20199 (N_20199,N_15489,N_16673);
nor U20200 (N_20200,N_19786,N_19561);
and U20201 (N_20201,N_17873,N_18055);
and U20202 (N_20202,N_17989,N_18443);
or U20203 (N_20203,N_18568,N_15027);
nand U20204 (N_20204,N_15822,N_15092);
or U20205 (N_20205,N_18491,N_16750);
and U20206 (N_20206,N_15795,N_16944);
and U20207 (N_20207,N_17791,N_16415);
and U20208 (N_20208,N_19868,N_16702);
and U20209 (N_20209,N_19204,N_18728);
nand U20210 (N_20210,N_17736,N_15166);
nand U20211 (N_20211,N_15289,N_16390);
nor U20212 (N_20212,N_15103,N_17948);
nand U20213 (N_20213,N_17847,N_19512);
nor U20214 (N_20214,N_16343,N_16358);
nor U20215 (N_20215,N_16454,N_18661);
or U20216 (N_20216,N_19003,N_15603);
nor U20217 (N_20217,N_16989,N_19165);
nor U20218 (N_20218,N_15538,N_16594);
nand U20219 (N_20219,N_19090,N_17897);
nand U20220 (N_20220,N_19685,N_18281);
nand U20221 (N_20221,N_17565,N_15115);
nand U20222 (N_20222,N_16431,N_18709);
or U20223 (N_20223,N_15446,N_19593);
nor U20224 (N_20224,N_18559,N_15298);
and U20225 (N_20225,N_16695,N_19146);
nand U20226 (N_20226,N_16651,N_17383);
nor U20227 (N_20227,N_17561,N_18982);
nand U20228 (N_20228,N_16810,N_18197);
xnor U20229 (N_20229,N_17722,N_19865);
nor U20230 (N_20230,N_17220,N_17213);
and U20231 (N_20231,N_17324,N_17536);
nand U20232 (N_20232,N_16568,N_17650);
nand U20233 (N_20233,N_19752,N_15900);
xnor U20234 (N_20234,N_19970,N_19254);
and U20235 (N_20235,N_19336,N_15970);
nand U20236 (N_20236,N_17699,N_17203);
or U20237 (N_20237,N_19082,N_17864);
nand U20238 (N_20238,N_18239,N_19225);
and U20239 (N_20239,N_18166,N_16636);
nor U20240 (N_20240,N_18674,N_15960);
nor U20241 (N_20241,N_18328,N_16212);
nor U20242 (N_20242,N_15256,N_19790);
or U20243 (N_20243,N_18653,N_15632);
or U20244 (N_20244,N_17687,N_19270);
and U20245 (N_20245,N_18207,N_18815);
and U20246 (N_20246,N_17657,N_15331);
and U20247 (N_20247,N_16569,N_18024);
or U20248 (N_20248,N_15362,N_19929);
or U20249 (N_20249,N_18179,N_18705);
and U20250 (N_20250,N_17166,N_16541);
nor U20251 (N_20251,N_19034,N_16895);
and U20252 (N_20252,N_15629,N_18325);
or U20253 (N_20253,N_18373,N_18181);
nand U20254 (N_20254,N_15734,N_19629);
nand U20255 (N_20255,N_15193,N_16083);
or U20256 (N_20256,N_19630,N_16194);
nor U20257 (N_20257,N_15349,N_19334);
or U20258 (N_20258,N_18652,N_19927);
or U20259 (N_20259,N_17257,N_15886);
nor U20260 (N_20260,N_16100,N_19906);
nor U20261 (N_20261,N_17360,N_18769);
or U20262 (N_20262,N_19153,N_15517);
nor U20263 (N_20263,N_16987,N_16732);
and U20264 (N_20264,N_19185,N_17539);
nand U20265 (N_20265,N_18943,N_16548);
nand U20266 (N_20266,N_16910,N_18339);
and U20267 (N_20267,N_17859,N_16314);
and U20268 (N_20268,N_15442,N_19797);
and U20269 (N_20269,N_15954,N_16026);
nor U20270 (N_20270,N_18957,N_19415);
nand U20271 (N_20271,N_17005,N_15228);
nand U20272 (N_20272,N_17039,N_19350);
nor U20273 (N_20273,N_16302,N_16951);
nor U20274 (N_20274,N_17357,N_17122);
xor U20275 (N_20275,N_19535,N_19645);
nand U20276 (N_20276,N_19953,N_15849);
and U20277 (N_20277,N_16036,N_18433);
and U20278 (N_20278,N_17240,N_15004);
or U20279 (N_20279,N_19145,N_19198);
and U20280 (N_20280,N_18523,N_15001);
nand U20281 (N_20281,N_15688,N_19641);
or U20282 (N_20282,N_17537,N_15952);
and U20283 (N_20283,N_16124,N_19819);
and U20284 (N_20284,N_16716,N_19338);
or U20285 (N_20285,N_18174,N_19321);
or U20286 (N_20286,N_15565,N_15185);
or U20287 (N_20287,N_17027,N_17698);
nor U20288 (N_20288,N_17860,N_19991);
nor U20289 (N_20289,N_16995,N_17173);
nand U20290 (N_20290,N_18838,N_18374);
nor U20291 (N_20291,N_17183,N_17377);
or U20292 (N_20292,N_18863,N_17425);
nand U20293 (N_20293,N_15485,N_17599);
and U20294 (N_20294,N_15633,N_16239);
nand U20295 (N_20295,N_18948,N_17373);
nor U20296 (N_20296,N_17690,N_19331);
nand U20297 (N_20297,N_18835,N_18877);
and U20298 (N_20298,N_17572,N_16982);
or U20299 (N_20299,N_16070,N_15833);
nand U20300 (N_20300,N_16525,N_16837);
nand U20301 (N_20301,N_19860,N_19783);
or U20302 (N_20302,N_18214,N_19770);
nand U20303 (N_20303,N_18327,N_19669);
or U20304 (N_20304,N_18810,N_17463);
nand U20305 (N_20305,N_17822,N_18353);
nand U20306 (N_20306,N_17507,N_15440);
and U20307 (N_20307,N_19665,N_17557);
nor U20308 (N_20308,N_16515,N_19516);
nand U20309 (N_20309,N_17768,N_17008);
and U20310 (N_20310,N_17652,N_15324);
nor U20311 (N_20311,N_18717,N_17215);
or U20312 (N_20312,N_19772,N_15595);
nand U20313 (N_20313,N_19503,N_15455);
nor U20314 (N_20314,N_19743,N_15790);
nor U20315 (N_20315,N_19227,N_18681);
nand U20316 (N_20316,N_16690,N_18340);
nand U20317 (N_20317,N_16127,N_19086);
and U20318 (N_20318,N_17582,N_17700);
nand U20319 (N_20319,N_19681,N_16309);
nand U20320 (N_20320,N_18990,N_19308);
nand U20321 (N_20321,N_19831,N_16146);
and U20322 (N_20322,N_17050,N_18090);
nor U20323 (N_20323,N_17025,N_17277);
nor U20324 (N_20324,N_16172,N_17194);
nand U20325 (N_20325,N_18394,N_18971);
nor U20326 (N_20326,N_15188,N_16405);
or U20327 (N_20327,N_16563,N_17226);
or U20328 (N_20328,N_17920,N_15307);
nor U20329 (N_20329,N_19682,N_16109);
nor U20330 (N_20330,N_19720,N_17888);
nor U20331 (N_20331,N_17943,N_15806);
nand U20332 (N_20332,N_15260,N_16262);
nor U20333 (N_20333,N_16134,N_18308);
and U20334 (N_20334,N_15809,N_19015);
nor U20335 (N_20335,N_16011,N_16136);
nor U20336 (N_20336,N_16751,N_16108);
or U20337 (N_20337,N_17713,N_18927);
xor U20338 (N_20338,N_19359,N_18463);
nor U20339 (N_20339,N_17007,N_18495);
nand U20340 (N_20340,N_19344,N_15829);
and U20341 (N_20341,N_16983,N_19464);
or U20342 (N_20342,N_15868,N_18131);
or U20343 (N_20343,N_16041,N_19813);
or U20344 (N_20344,N_16811,N_15501);
nor U20345 (N_20345,N_18758,N_18019);
nand U20346 (N_20346,N_15106,N_16813);
nand U20347 (N_20347,N_15958,N_16609);
and U20348 (N_20348,N_18626,N_19725);
or U20349 (N_20349,N_15206,N_16841);
nor U20350 (N_20350,N_18229,N_18573);
nand U20351 (N_20351,N_18608,N_17239);
nand U20352 (N_20352,N_16659,N_16089);
nor U20353 (N_20353,N_17829,N_18752);
xor U20354 (N_20354,N_17589,N_17028);
nand U20355 (N_20355,N_18792,N_17424);
nor U20356 (N_20356,N_15977,N_19459);
nor U20357 (N_20357,N_15010,N_15549);
nand U20358 (N_20358,N_15119,N_15100);
nor U20359 (N_20359,N_17692,N_19194);
and U20360 (N_20360,N_18985,N_19834);
and U20361 (N_20361,N_17827,N_15290);
or U20362 (N_20362,N_15909,N_18689);
and U20363 (N_20363,N_17825,N_15101);
or U20364 (N_20364,N_16122,N_15340);
or U20365 (N_20365,N_18749,N_15377);
or U20366 (N_20366,N_18284,N_16739);
and U20367 (N_20367,N_15799,N_19647);
and U20368 (N_20368,N_16062,N_16937);
or U20369 (N_20369,N_15898,N_16063);
or U20370 (N_20370,N_15940,N_18226);
xnor U20371 (N_20371,N_16802,N_18338);
nand U20372 (N_20372,N_19867,N_18140);
nand U20373 (N_20373,N_17255,N_18032);
nor U20374 (N_20374,N_19243,N_15575);
nand U20375 (N_20375,N_17444,N_18020);
and U20376 (N_20376,N_16963,N_16035);
or U20377 (N_20377,N_18014,N_16890);
and U20378 (N_20378,N_15144,N_17428);
and U20379 (N_20379,N_18788,N_17558);
and U20380 (N_20380,N_16111,N_17461);
or U20381 (N_20381,N_18896,N_15018);
and U20382 (N_20382,N_16534,N_15189);
and U20383 (N_20383,N_19693,N_16591);
nand U20384 (N_20384,N_17342,N_18793);
and U20385 (N_20385,N_16219,N_15525);
and U20386 (N_20386,N_18726,N_18718);
and U20387 (N_20387,N_16726,N_16599);
nor U20388 (N_20388,N_17081,N_15917);
xor U20389 (N_20389,N_15863,N_16589);
xnor U20390 (N_20390,N_16336,N_15475);
nand U20391 (N_20391,N_16285,N_18802);
nand U20392 (N_20392,N_17490,N_18127);
nor U20393 (N_20393,N_17985,N_16113);
nand U20394 (N_20394,N_16528,N_17750);
or U20395 (N_20395,N_15152,N_17514);
nor U20396 (N_20396,N_15893,N_17010);
and U20397 (N_20397,N_17889,N_17781);
nor U20398 (N_20398,N_19127,N_15327);
and U20399 (N_20399,N_17190,N_16740);
and U20400 (N_20400,N_19656,N_17370);
nand U20401 (N_20401,N_18737,N_19607);
and U20402 (N_20402,N_16847,N_15716);
or U20403 (N_20403,N_19825,N_19829);
xor U20404 (N_20404,N_16117,N_19869);
or U20405 (N_20405,N_19317,N_16959);
nand U20406 (N_20406,N_16560,N_17879);
nand U20407 (N_20407,N_18212,N_19862);
and U20408 (N_20408,N_17392,N_17919);
nand U20409 (N_20409,N_16527,N_18829);
nor U20410 (N_20410,N_19827,N_17794);
or U20411 (N_20411,N_18952,N_18506);
nand U20412 (N_20412,N_17052,N_17637);
and U20413 (N_20413,N_19922,N_19689);
or U20414 (N_20414,N_19022,N_17209);
nor U20415 (N_20415,N_18822,N_18736);
or U20416 (N_20416,N_19703,N_16015);
or U20417 (N_20417,N_17445,N_16872);
or U20418 (N_20418,N_15523,N_17562);
nor U20419 (N_20419,N_18108,N_19242);
nor U20420 (N_20420,N_19140,N_18796);
nand U20421 (N_20421,N_16857,N_17400);
nor U20422 (N_20422,N_16341,N_15636);
nand U20423 (N_20423,N_15939,N_15096);
nand U20424 (N_20424,N_16271,N_17110);
nand U20425 (N_20425,N_15212,N_15546);
nor U20426 (N_20426,N_16796,N_17676);
and U20427 (N_20427,N_17295,N_19983);
or U20428 (N_20428,N_18424,N_18638);
nor U20429 (N_20429,N_19282,N_16342);
nor U20430 (N_20430,N_18008,N_18917);
or U20431 (N_20431,N_15582,N_15561);
nor U20432 (N_20432,N_16578,N_15192);
nor U20433 (N_20433,N_16940,N_19800);
nor U20434 (N_20434,N_15461,N_16631);
nand U20435 (N_20435,N_15956,N_19302);
nor U20436 (N_20436,N_18449,N_16417);
nor U20437 (N_20437,N_16974,N_19591);
or U20438 (N_20438,N_15593,N_19496);
and U20439 (N_20439,N_18201,N_19558);
and U20440 (N_20440,N_17312,N_16622);
and U20441 (N_20441,N_17026,N_15877);
or U20442 (N_20442,N_19602,N_15443);
or U20443 (N_20443,N_15610,N_19695);
nand U20444 (N_20444,N_17662,N_17484);
nand U20445 (N_20445,N_17218,N_18692);
and U20446 (N_20446,N_16295,N_19622);
and U20447 (N_20447,N_16808,N_16312);
or U20448 (N_20448,N_19139,N_17581);
and U20449 (N_20449,N_16626,N_18902);
or U20450 (N_20450,N_17647,N_18235);
or U20451 (N_20451,N_19491,N_18748);
or U20452 (N_20452,N_16091,N_16220);
nand U20453 (N_20453,N_16546,N_17862);
nor U20454 (N_20454,N_15836,N_17129);
or U20455 (N_20455,N_18852,N_19858);
nor U20456 (N_20456,N_17866,N_18196);
and U20457 (N_20457,N_17199,N_19540);
nand U20458 (N_20458,N_15341,N_17502);
and U20459 (N_20459,N_18731,N_17249);
xnor U20460 (N_20460,N_17578,N_15639);
and U20461 (N_20461,N_19509,N_17877);
or U20462 (N_20462,N_19979,N_16481);
and U20463 (N_20463,N_18036,N_15354);
nand U20464 (N_20464,N_19796,N_17865);
or U20465 (N_20465,N_16706,N_19332);
nand U20466 (N_20466,N_18377,N_17752);
or U20467 (N_20467,N_15305,N_17627);
nor U20468 (N_20468,N_19735,N_15360);
and U20469 (N_20469,N_16086,N_16676);
and U20470 (N_20470,N_17251,N_18352);
or U20471 (N_20471,N_15365,N_17212);
nor U20472 (N_20472,N_17732,N_15195);
nand U20473 (N_20473,N_15457,N_15889);
and U20474 (N_20474,N_15286,N_17088);
nor U20475 (N_20475,N_16416,N_17348);
nand U20476 (N_20476,N_19610,N_17819);
nand U20477 (N_20477,N_15227,N_18539);
xnor U20478 (N_20478,N_17334,N_19613);
or U20479 (N_20479,N_19477,N_16171);
nor U20480 (N_20480,N_15899,N_18972);
and U20481 (N_20481,N_16905,N_15385);
or U20482 (N_20482,N_17418,N_19731);
nor U20483 (N_20483,N_16887,N_15170);
and U20484 (N_20484,N_18801,N_16962);
and U20485 (N_20485,N_19000,N_15056);
and U20486 (N_20486,N_17869,N_15214);
and U20487 (N_20487,N_18384,N_15731);
or U20488 (N_20488,N_18043,N_19776);
or U20489 (N_20489,N_18926,N_18202);
nand U20490 (N_20490,N_16024,N_15448);
or U20491 (N_20491,N_17172,N_19577);
or U20492 (N_20492,N_19779,N_19741);
nand U20493 (N_20493,N_16251,N_18040);
or U20494 (N_20494,N_18345,N_19506);
and U20495 (N_20495,N_19470,N_16120);
or U20496 (N_20496,N_15548,N_19171);
nand U20497 (N_20497,N_16282,N_18033);
nor U20498 (N_20498,N_17741,N_18037);
nand U20499 (N_20499,N_18025,N_19866);
and U20500 (N_20500,N_15817,N_16587);
and U20501 (N_20501,N_18157,N_18651);
or U20502 (N_20502,N_18408,N_15515);
nor U20503 (N_20503,N_18265,N_19801);
nor U20504 (N_20504,N_19864,N_19908);
and U20505 (N_20505,N_19963,N_15049);
or U20506 (N_20506,N_18160,N_16820);
nand U20507 (N_20507,N_19356,N_18407);
nand U20508 (N_20508,N_17272,N_18082);
or U20509 (N_20509,N_17623,N_16006);
and U20510 (N_20510,N_18326,N_18649);
nor U20511 (N_20511,N_15099,N_16540);
or U20512 (N_20512,N_17024,N_15707);
nand U20513 (N_20513,N_19926,N_19769);
or U20514 (N_20514,N_15678,N_19534);
and U20515 (N_20515,N_18818,N_15468);
or U20516 (N_20516,N_19420,N_17622);
and U20517 (N_20517,N_19634,N_19729);
nand U20518 (N_20518,N_19007,N_16865);
nor U20519 (N_20519,N_18359,N_17624);
nor U20520 (N_20520,N_19038,N_16939);
and U20521 (N_20521,N_17772,N_17712);
nand U20522 (N_20522,N_19472,N_17509);
or U20523 (N_20523,N_18825,N_15416);
nand U20524 (N_20524,N_17064,N_15723);
nand U20525 (N_20525,N_16861,N_16033);
and U20526 (N_20526,N_16866,N_16529);
and U20527 (N_20527,N_19394,N_15769);
or U20528 (N_20528,N_17689,N_18178);
or U20529 (N_20529,N_19016,N_17930);
or U20530 (N_20530,N_19316,N_18453);
nand U20531 (N_20531,N_15791,N_15357);
nor U20532 (N_20532,N_18931,N_19440);
or U20533 (N_20533,N_19627,N_18172);
nor U20534 (N_20534,N_15567,N_15081);
nand U20535 (N_20535,N_15064,N_18150);
nor U20536 (N_20536,N_19942,N_15431);
nand U20537 (N_20537,N_16147,N_18089);
nand U20538 (N_20538,N_19271,N_18669);
and U20539 (N_20539,N_16526,N_16180);
and U20540 (N_20540,N_17760,N_18283);
and U20541 (N_20541,N_19545,N_17685);
and U20542 (N_20542,N_19652,N_15987);
or U20543 (N_20543,N_18060,N_19672);
nor U20544 (N_20544,N_18906,N_17832);
and U20545 (N_20545,N_19474,N_15540);
nor U20546 (N_20546,N_15111,N_18534);
and U20547 (N_20547,N_16463,N_16005);
or U20548 (N_20548,N_15320,N_18850);
nor U20549 (N_20549,N_17036,N_15529);
xnor U20550 (N_20550,N_18349,N_16602);
nor U20551 (N_20551,N_19278,N_17160);
and U20552 (N_20552,N_18124,N_15858);
or U20553 (N_20553,N_15646,N_18770);
and U20554 (N_20554,N_17116,N_16722);
nor U20555 (N_20555,N_19728,N_19386);
and U20556 (N_20556,N_18541,N_16835);
and U20557 (N_20557,N_17403,N_16886);
nor U20558 (N_20558,N_16363,N_16649);
nand U20559 (N_20559,N_19907,N_19818);
and U20560 (N_20560,N_16647,N_16742);
nor U20561 (N_20561,N_17932,N_17803);
and U20562 (N_20562,N_18233,N_17293);
and U20563 (N_20563,N_15374,N_15429);
and U20564 (N_20564,N_17167,N_18930);
nand U20565 (N_20565,N_15653,N_19190);
nand U20566 (N_20566,N_15138,N_15222);
nand U20567 (N_20567,N_15647,N_16513);
nor U20568 (N_20568,N_17531,N_19552);
or U20569 (N_20569,N_16613,N_17946);
nand U20570 (N_20570,N_17069,N_18388);
or U20571 (N_20571,N_18113,N_16776);
and U20572 (N_20572,N_15623,N_15181);
or U20573 (N_20573,N_19151,N_19025);
or U20574 (N_20574,N_18266,N_16806);
or U20575 (N_20575,N_17135,N_15867);
or U20576 (N_20576,N_18248,N_18455);
or U20577 (N_20577,N_18962,N_15651);
xor U20578 (N_20578,N_15389,N_18220);
nor U20579 (N_20579,N_18960,N_16489);
and U20580 (N_20580,N_16173,N_19195);
or U20581 (N_20581,N_17330,N_17955);
and U20582 (N_20582,N_18395,N_19863);
and U20583 (N_20583,N_19258,N_16704);
nand U20584 (N_20584,N_18954,N_15165);
nand U20585 (N_20585,N_16797,N_18511);
nor U20586 (N_20586,N_17905,N_17248);
or U20587 (N_20587,N_19596,N_16214);
nor U20588 (N_20588,N_17242,N_17775);
nand U20589 (N_20589,N_18288,N_19110);
or U20590 (N_20590,N_18767,N_19696);
and U20591 (N_20591,N_16842,N_17538);
or U20592 (N_20592,N_19917,N_18079);
and U20593 (N_20593,N_16004,N_15265);
nand U20594 (N_20594,N_19851,N_18938);
and U20595 (N_20595,N_19285,N_19586);
nor U20596 (N_20596,N_19919,N_15024);
or U20597 (N_20597,N_16465,N_15381);
and U20598 (N_20598,N_19216,N_17563);
nor U20599 (N_20599,N_17308,N_15770);
nor U20600 (N_20600,N_16919,N_19612);
nor U20601 (N_20601,N_19298,N_19678);
and U20602 (N_20602,N_15419,N_16762);
nor U20603 (N_20603,N_16656,N_15611);
and U20604 (N_20604,N_18347,N_16097);
or U20605 (N_20605,N_17450,N_16174);
or U20606 (N_20606,N_18120,N_16681);
nand U20607 (N_20607,N_19401,N_15146);
and U20608 (N_20608,N_17523,N_15919);
or U20609 (N_20609,N_17123,N_15441);
nand U20610 (N_20610,N_18757,N_19840);
nand U20611 (N_20611,N_18389,N_17385);
and U20612 (N_20612,N_17082,N_17727);
nor U20613 (N_20613,N_17653,N_17328);
or U20614 (N_20614,N_17494,N_16733);
nor U20615 (N_20615,N_16682,N_19276);
nor U20616 (N_20616,N_18189,N_18459);
or U20617 (N_20617,N_17058,N_17535);
and U20618 (N_20618,N_16891,N_17566);
and U20619 (N_20619,N_19980,N_18794);
nand U20620 (N_20620,N_19020,N_18367);
and U20621 (N_20621,N_18194,N_15275);
nor U20622 (N_20622,N_17405,N_18677);
nor U20623 (N_20623,N_17788,N_19410);
xnor U20624 (N_20624,N_18085,N_16586);
nor U20625 (N_20625,N_18601,N_16965);
and U20626 (N_20626,N_15733,N_19319);
and U20627 (N_20627,N_17735,N_17352);
or U20628 (N_20628,N_18891,N_18121);
xor U20629 (N_20629,N_15091,N_16616);
nand U20630 (N_20630,N_19396,N_18099);
or U20631 (N_20631,N_16590,N_16210);
nand U20632 (N_20632,N_16169,N_17458);
or U20633 (N_20633,N_15800,N_15712);
or U20634 (N_20634,N_16839,N_17144);
and U20635 (N_20635,N_18276,N_15771);
nor U20636 (N_20636,N_18341,N_18291);
and U20637 (N_20637,N_18610,N_15729);
xor U20638 (N_20638,N_15255,N_17040);
or U20639 (N_20639,N_19969,N_18117);
nand U20640 (N_20640,N_16380,N_18831);
nand U20641 (N_20641,N_19423,N_16475);
nand U20642 (N_20642,N_18513,N_19894);
or U20643 (N_20643,N_19550,N_16060);
and U20644 (N_20644,N_15277,N_18278);
nand U20645 (N_20645,N_18440,N_16068);
nand U20646 (N_20646,N_18029,N_17613);
nor U20647 (N_20647,N_17184,N_19408);
nand U20648 (N_20648,N_17753,N_18222);
nand U20649 (N_20649,N_15343,N_17776);
xor U20650 (N_20650,N_17369,N_18507);
nor U20651 (N_20651,N_18645,N_18816);
xnor U20652 (N_20652,N_16713,N_19076);
nor U20653 (N_20653,N_17035,N_16348);
nand U20654 (N_20654,N_18668,N_17294);
nand U20655 (N_20655,N_16670,N_17952);
xor U20656 (N_20656,N_17815,N_18888);
nor U20657 (N_20657,N_15157,N_17926);
nand U20658 (N_20658,N_19362,N_15701);
nor U20659 (N_20659,N_17228,N_19322);
or U20660 (N_20660,N_19643,N_18897);
or U20661 (N_20661,N_18518,N_15355);
or U20662 (N_20662,N_19058,N_18116);
nand U20663 (N_20663,N_18561,N_17660);
nor U20664 (N_20664,N_18072,N_16803);
and U20665 (N_20665,N_19019,N_17959);
nor U20666 (N_20666,N_19104,N_17634);
nor U20667 (N_20667,N_19531,N_19281);
and U20668 (N_20668,N_19373,N_18723);
or U20669 (N_20669,N_17271,N_17663);
and U20670 (N_20670,N_19901,N_19390);
nand U20671 (N_20671,N_15116,N_16918);
nand U20672 (N_20672,N_19467,N_18773);
nand U20673 (N_20673,N_16728,N_15197);
nor U20674 (N_20674,N_17874,N_15346);
and U20675 (N_20675,N_15180,N_17060);
and U20676 (N_20676,N_18362,N_16687);
nor U20677 (N_20677,N_19603,N_17137);
or U20678 (N_20678,N_18720,N_15009);
nand U20679 (N_20679,N_16507,N_17922);
and U20680 (N_20680,N_17824,N_19782);
nor U20681 (N_20681,N_17666,N_18218);
and U20682 (N_20682,N_19481,N_16485);
and U20683 (N_20683,N_15801,N_19845);
or U20684 (N_20684,N_16338,N_16972);
or U20685 (N_20685,N_17890,N_15759);
nand U20686 (N_20686,N_15159,N_17520);
xnor U20687 (N_20687,N_17820,N_18746);
or U20688 (N_20688,N_19071,N_18319);
nor U20689 (N_20689,N_18824,N_19269);
and U20690 (N_20690,N_15676,N_17929);
or U20691 (N_20691,N_16648,N_17414);
nand U20692 (N_20692,N_15129,N_15747);
nand U20693 (N_20693,N_18155,N_19008);
nor U20694 (N_20694,N_16663,N_18400);
or U20695 (N_20695,N_15741,N_19924);
nand U20696 (N_20696,N_16868,N_18602);
or U20697 (N_20697,N_16167,N_17619);
or U20698 (N_20698,N_15474,N_17857);
xnor U20699 (N_20699,N_17047,N_15174);
or U20700 (N_20700,N_15005,N_19049);
or U20701 (N_20701,N_19737,N_19802);
nand U20702 (N_20702,N_15746,N_15781);
nand U20703 (N_20703,N_19519,N_15990);
xor U20704 (N_20704,N_19609,N_18062);
or U20705 (N_20705,N_18684,N_19997);
nand U20706 (N_20706,N_19878,N_18725);
nor U20707 (N_20707,N_18630,N_17579);
and U20708 (N_20708,N_17051,N_19734);
and U20709 (N_20709,N_19808,N_16730);
nand U20710 (N_20710,N_15606,N_19523);
or U20711 (N_20711,N_16934,N_18109);
nor U20712 (N_20712,N_15395,N_19686);
nand U20713 (N_20713,N_16611,N_19758);
and U20714 (N_20714,N_16471,N_17602);
nand U20715 (N_20715,N_19117,N_15464);
nor U20716 (N_20716,N_19182,N_19325);
and U20717 (N_20717,N_18612,N_15089);
or U20718 (N_20718,N_16201,N_16661);
nand U20719 (N_20719,N_15432,N_17971);
nor U20720 (N_20720,N_16023,N_15450);
nor U20721 (N_20721,N_17814,N_15083);
or U20722 (N_20722,N_16215,N_16830);
and U20723 (N_20723,N_17921,N_15766);
or U20724 (N_20724,N_18297,N_15579);
and U20725 (N_20725,N_16854,N_19520);
nor U20726 (N_20726,N_19073,N_17821);
and U20727 (N_20727,N_15887,N_19632);
nand U20728 (N_20728,N_17632,N_15364);
nor U20729 (N_20729,N_17269,N_19041);
and U20730 (N_20730,N_18567,N_15151);
and U20731 (N_20731,N_15521,N_17705);
and U20732 (N_20732,N_19508,N_18893);
or U20733 (N_20733,N_16396,N_19974);
and U20734 (N_20734,N_16002,N_18582);
nor U20735 (N_20735,N_18290,N_19446);
nand U20736 (N_20736,N_19952,N_15607);
nand U20737 (N_20737,N_17133,N_16877);
nor U20738 (N_20738,N_16221,N_16580);
xnor U20739 (N_20739,N_17473,N_16297);
nor U20740 (N_20740,N_17196,N_15727);
nor U20741 (N_20741,N_17725,N_17104);
or U20742 (N_20742,N_19653,N_18441);
nand U20743 (N_20743,N_17384,N_16931);
or U20744 (N_20744,N_18144,N_19637);
nand U20745 (N_20745,N_15309,N_17998);
or U20746 (N_20746,N_15248,N_18678);
xor U20747 (N_20747,N_17020,N_17394);
nor U20748 (N_20748,N_16638,N_15621);
and U20749 (N_20749,N_17376,N_18809);
nor U20750 (N_20750,N_18743,N_15753);
nand U20751 (N_20751,N_17454,N_18393);
nor U20752 (N_20752,N_15386,N_16286);
or U20753 (N_20753,N_18078,N_15554);
nand U20754 (N_20754,N_19197,N_17671);
nor U20755 (N_20755,N_15124,N_18137);
nor U20756 (N_20756,N_16948,N_15117);
nor U20757 (N_20757,N_16533,N_19132);
and U20758 (N_20758,N_15259,N_17074);
or U20759 (N_20759,N_16355,N_15231);
or U20760 (N_20760,N_16885,N_18125);
nor U20761 (N_20761,N_17031,N_19147);
and U20762 (N_20762,N_17789,N_19437);
nand U20763 (N_20763,N_18343,N_18331);
or U20764 (N_20764,N_17102,N_18210);
and U20765 (N_20765,N_18295,N_19854);
or U20766 (N_20766,N_19100,N_15696);
or U20767 (N_20767,N_15533,N_18517);
or U20768 (N_20768,N_19438,N_19700);
and U20769 (N_20769,N_16430,N_15453);
and U20770 (N_20770,N_17004,N_19215);
nor U20771 (N_20771,N_19832,N_15452);
or U20772 (N_20772,N_19284,N_15618);
nand U20773 (N_20773,N_15969,N_15943);
nor U20774 (N_20774,N_16170,N_19575);
and U20775 (N_20775,N_15574,N_19419);
nand U20776 (N_20776,N_18867,N_18485);
nand U20777 (N_20777,N_16392,N_17111);
and U20778 (N_20778,N_16498,N_15585);
nand U20779 (N_20779,N_19340,N_17983);
or U20780 (N_20780,N_18995,N_19938);
or U20781 (N_20781,N_17397,N_15536);
nand U20782 (N_20782,N_15519,N_19017);
nor U20783 (N_20783,N_16607,N_19358);
nor U20784 (N_20784,N_17427,N_17583);
and U20785 (N_20785,N_19756,N_15657);
nor U20786 (N_20786,N_15823,N_18522);
nand U20787 (N_20787,N_18363,N_16980);
or U20788 (N_20788,N_19177,N_15445);
and U20789 (N_20789,N_16466,N_18997);
or U20790 (N_20790,N_19642,N_17097);
xnor U20791 (N_20791,N_19256,N_16275);
xnor U20792 (N_20792,N_18504,N_17211);
or U20793 (N_20793,N_18253,N_18263);
xor U20794 (N_20794,N_19366,N_19130);
and U20795 (N_20795,N_19722,N_19943);
and U20796 (N_20796,N_17960,N_18279);
or U20797 (N_20797,N_16008,N_16186);
or U20798 (N_20798,N_16952,N_16514);
nor U20799 (N_20799,N_19674,N_19150);
or U20800 (N_20800,N_18169,N_19846);
nand U20801 (N_20801,N_17073,N_18051);
nor U20802 (N_20802,N_15237,N_17780);
and U20803 (N_20803,N_17095,N_16434);
and U20804 (N_20804,N_18899,N_15656);
nand U20805 (N_20805,N_18759,N_17157);
nor U20806 (N_20806,N_19057,N_18337);
and U20807 (N_20807,N_19538,N_16490);
or U20808 (N_20808,N_17399,N_15029);
or U20809 (N_20809,N_19021,N_17214);
nand U20810 (N_20810,N_15074,N_18679);
nor U20811 (N_20811,N_17546,N_19502);
nor U20812 (N_20812,N_16182,N_17206);
nor U20813 (N_20813,N_18243,N_15921);
xnor U20814 (N_20814,N_17972,N_19426);
nand U20815 (N_20815,N_16317,N_16853);
nor U20816 (N_20816,N_15037,N_15478);
or U20817 (N_20817,N_19903,N_15665);
nor U20818 (N_20818,N_18175,N_16672);
or U20819 (N_20819,N_19333,N_17440);
and U20820 (N_20820,N_18929,N_15927);
or U20821 (N_20821,N_16102,N_17965);
and U20822 (N_20822,N_19711,N_15470);
nand U20823 (N_20823,N_19412,N_17270);
or U20824 (N_20824,N_17717,N_18225);
nor U20825 (N_20825,N_17011,N_19954);
nand U20826 (N_20826,N_19588,N_17590);
or U20827 (N_20827,N_16539,N_16095);
and U20828 (N_20828,N_16044,N_18501);
xnor U20829 (N_20829,N_16826,N_18396);
nor U20830 (N_20830,N_17446,N_16639);
xnor U20831 (N_20831,N_16749,N_15907);
or U20832 (N_20832,N_18685,N_15721);
nor U20833 (N_20833,N_19389,N_19180);
and U20834 (N_20834,N_17739,N_17260);
nor U20835 (N_20835,N_15796,N_16482);
nand U20836 (N_20836,N_17828,N_17664);
and U20837 (N_20837,N_19764,N_16969);
nor U20838 (N_20838,N_16581,N_17029);
and U20839 (N_20839,N_19814,N_18429);
nand U20840 (N_20840,N_17986,N_17387);
nand U20841 (N_20841,N_16273,N_18646);
nand U20842 (N_20842,N_18417,N_18741);
nor U20843 (N_20843,N_18286,N_18676);
nor U20844 (N_20844,N_18105,N_17608);
and U20845 (N_20845,N_18618,N_18722);
nand U20846 (N_20846,N_16763,N_19381);
nand U20847 (N_20847,N_16502,N_18171);
nor U20848 (N_20848,N_18719,N_17907);
nand U20849 (N_20849,N_17769,N_15098);
or U20850 (N_20850,N_17568,N_19768);
and U20851 (N_20851,N_19848,N_19203);
and U20852 (N_20852,N_15666,N_15156);
xnor U20853 (N_20853,N_19835,N_16432);
nand U20854 (N_20854,N_16858,N_17350);
and U20855 (N_20855,N_15178,N_19047);
or U20856 (N_20856,N_16073,N_18492);
or U20857 (N_20857,N_15961,N_18311);
nand U20858 (N_20858,N_17009,N_15989);
and U20859 (N_20859,N_19393,N_16468);
nand U20860 (N_20860,N_16992,N_17994);
nor U20861 (N_20861,N_18548,N_18324);
nor U20862 (N_20862,N_18693,N_19012);
nand U20863 (N_20863,N_16495,N_17908);
nand U20864 (N_20864,N_19088,N_19717);
nand U20865 (N_20865,N_19075,N_19222);
nand U20866 (N_20866,N_16032,N_19014);
and U20867 (N_20867,N_15079,N_17549);
and U20868 (N_20868,N_17938,N_19988);
and U20869 (N_20869,N_18271,N_16072);
nand U20870 (N_20870,N_18524,N_15944);
or U20871 (N_20871,N_15493,N_18039);
nor U20872 (N_20872,N_18292,N_15406);
nand U20873 (N_20873,N_16408,N_18161);
or U20874 (N_20874,N_17527,N_17455);
nor U20875 (N_20875,N_18551,N_16909);
or U20876 (N_20876,N_17759,N_17661);
and U20877 (N_20877,N_15797,N_19740);
or U20878 (N_20878,N_15015,N_16101);
or U20879 (N_20879,N_15161,N_16753);
nor U20880 (N_20880,N_19201,N_18560);
and U20881 (N_20881,N_15953,N_19931);
or U20882 (N_20882,N_15689,N_16958);
nor U20883 (N_20883,N_16494,N_17168);
nor U20884 (N_20884,N_17724,N_16442);
nand U20885 (N_20885,N_15458,N_17106);
and U20886 (N_20886,N_17100,N_17422);
and U20887 (N_20887,N_17015,N_17525);
nand U20888 (N_20888,N_19836,N_19673);
nand U20889 (N_20889,N_18476,N_16664);
nor U20890 (N_20890,N_17191,N_18708);
nor U20891 (N_20891,N_19441,N_18603);
and U20892 (N_20892,N_18094,N_18826);
nand U20893 (N_20893,N_16583,N_15071);
nor U20894 (N_20894,N_15946,N_15634);
or U20895 (N_20895,N_17164,N_17614);
xnor U20896 (N_20896,N_19918,N_18740);
nand U20897 (N_20897,N_19094,N_17259);
nor U20898 (N_20898,N_16293,N_15642);
nand U20899 (N_20899,N_15358,N_15860);
or U20900 (N_20900,N_16917,N_19746);
nor U20901 (N_20901,N_15649,N_17287);
nand U20902 (N_20902,N_17718,N_15383);
and U20903 (N_20903,N_15818,N_19698);
nand U20904 (N_20904,N_15506,N_15526);
nand U20905 (N_20905,N_16970,N_18101);
nor U20906 (N_20906,N_18223,N_16027);
or U20907 (N_20907,N_17630,N_15985);
nand U20908 (N_20908,N_19578,N_15694);
nand U20909 (N_20909,N_18031,N_19402);
or U20910 (N_20910,N_18922,N_17766);
nand U20911 (N_20911,N_17701,N_18460);
nor U20912 (N_20912,N_17476,N_19347);
nand U20913 (N_20913,N_15811,N_19288);
or U20914 (N_20914,N_17306,N_16259);
and U20915 (N_20915,N_16880,N_17187);
and U20916 (N_20916,N_16255,N_18215);
nor U20917 (N_20917,N_16371,N_18209);
nor U20918 (N_20918,N_16470,N_17210);
and U20919 (N_20919,N_18010,N_17247);
nand U20920 (N_20920,N_18571,N_15109);
nor U20921 (N_20921,N_16118,N_17439);
nor U20922 (N_20922,N_18493,N_17301);
and U20923 (N_20923,N_19902,N_15930);
nor U20924 (N_20924,N_17262,N_15315);
and U20925 (N_20925,N_15876,N_18366);
and U20926 (N_20926,N_19941,N_16818);
nor U20927 (N_20927,N_19937,N_19950);
nor U20928 (N_20928,N_16772,N_19709);
and U20929 (N_20929,N_16264,N_17408);
nor U20930 (N_20930,N_19625,N_17256);
nand U20931 (N_20931,N_19246,N_19473);
and U20932 (N_20932,N_18375,N_19101);
or U20933 (N_20933,N_17616,N_17407);
nor U20934 (N_20934,N_19702,N_18041);
and U20935 (N_20935,N_19045,N_18071);
or U20936 (N_20936,N_15590,N_18213);
nand U20937 (N_20937,N_18047,N_16743);
nand U20938 (N_20938,N_16543,N_18228);
or U20939 (N_20939,N_17798,N_16752);
and U20940 (N_20940,N_15239,N_17053);
or U20941 (N_20941,N_18992,N_15447);
nand U20942 (N_20942,N_17067,N_18154);
or U20943 (N_20943,N_15072,N_18832);
and U20944 (N_20944,N_15683,N_18845);
or U20945 (N_20945,N_16792,N_19042);
nor U20946 (N_20946,N_19727,N_19361);
or U20947 (N_20947,N_16398,N_15730);
nand U20948 (N_20948,N_19228,N_16267);
nor U20949 (N_20949,N_16584,N_18456);
or U20950 (N_20950,N_17674,N_19326);
nand U20951 (N_20951,N_17807,N_17038);
and U20952 (N_20952,N_15920,N_16410);
nor U20953 (N_20953,N_15285,N_16247);
and U20954 (N_20954,N_19122,N_17366);
or U20955 (N_20955,N_18776,N_16815);
and U20956 (N_20956,N_15856,N_17415);
nand U20957 (N_20957,N_18680,N_15810);
or U20958 (N_20958,N_15224,N_19187);
nand U20959 (N_20959,N_17396,N_18066);
and U20960 (N_20960,N_17675,N_17098);
and U20961 (N_20961,N_17349,N_19120);
nand U20962 (N_20962,N_18937,N_15933);
nand U20963 (N_20963,N_16053,N_16666);
and U20964 (N_20964,N_15133,N_18333);
nor U20965 (N_20965,N_17516,N_15573);
nand U20966 (N_20966,N_17083,N_15890);
nand U20967 (N_20967,N_16473,N_19606);
or U20968 (N_20968,N_15208,N_16085);
and U20969 (N_20969,N_19337,N_17288);
and U20970 (N_20970,N_15951,N_15276);
nor U20971 (N_20971,N_15855,N_16446);
and U20972 (N_20972,N_19972,N_18817);
or U20973 (N_20973,N_19184,N_18820);
or U20974 (N_20974,N_15635,N_17804);
or U20975 (N_20975,N_18296,N_17059);
nand U20976 (N_20976,N_15615,N_16107);
nand U20977 (N_20977,N_17169,N_19915);
nor U20978 (N_20978,N_19923,N_19456);
and U20979 (N_20979,N_19909,N_18195);
nor U20980 (N_20980,N_19152,N_17551);
and U20981 (N_20981,N_17289,N_16104);
nor U20982 (N_20982,N_18001,N_19428);
xnor U20983 (N_20983,N_16084,N_15862);
and U20984 (N_20984,N_17816,N_16403);
or U20985 (N_20985,N_19701,N_15749);
or U20986 (N_20986,N_15700,N_16202);
or U20987 (N_20987,N_18951,N_15060);
and U20988 (N_20988,N_16973,N_18624);
and U20989 (N_20989,N_17673,N_15901);
or U20990 (N_20990,N_15269,N_17969);
and U20991 (N_20991,N_18915,N_17709);
nor U20992 (N_20992,N_18486,N_17902);
and U20993 (N_20993,N_19290,N_18361);
nor U20994 (N_20994,N_15213,N_18376);
nand U20995 (N_20995,N_18191,N_18293);
and U20996 (N_20996,N_16372,N_15513);
nand U20997 (N_20997,N_16619,N_15462);
or U20998 (N_20998,N_17830,N_16968);
nor U20999 (N_20999,N_16574,N_18544);
or U21000 (N_21000,N_16192,N_18625);
nand U21001 (N_21001,N_16444,N_15583);
nor U21002 (N_21002,N_17529,N_18164);
xnor U21003 (N_21003,N_18368,N_18526);
and U21004 (N_21004,N_15592,N_18383);
or U21005 (N_21005,N_17987,N_15281);
nor U21006 (N_21006,N_16126,N_15627);
nor U21007 (N_21007,N_18575,N_18823);
or U21008 (N_21008,N_16025,N_15844);
nand U21009 (N_21009,N_19461,N_19987);
nor U21010 (N_21010,N_17291,N_17316);
nor U21011 (N_21011,N_15272,N_16869);
or U21012 (N_21012,N_19312,N_19378);
nand U21013 (N_21013,N_15233,N_18106);
nor U21014 (N_21014,N_16137,N_19500);
nor U21015 (N_21015,N_18437,N_18027);
or U21016 (N_21016,N_19061,N_17597);
and U21017 (N_21017,N_16767,N_19385);
nand U21018 (N_21018,N_19671,N_19060);
and U21019 (N_21019,N_17504,N_17409);
or U21020 (N_21020,N_19160,N_18193);
nor U21021 (N_21021,N_17101,N_15496);
nor U21022 (N_21022,N_18895,N_15761);
and U21023 (N_21023,N_16235,N_16020);
nand U21024 (N_21024,N_18490,N_19044);
nor U21025 (N_21025,N_16771,N_19462);
nor U21026 (N_21026,N_17846,N_18984);
and U21027 (N_21027,N_19168,N_18656);
and U21028 (N_21028,N_16635,N_17799);
or U21029 (N_21029,N_15775,N_19095);
and U21030 (N_21030,N_19973,N_18477);
and U21031 (N_21031,N_17438,N_16836);
or U21032 (N_21032,N_17812,N_19369);
nand U21033 (N_21033,N_18302,N_15038);
and U21034 (N_21034,N_18980,N_19141);
nand U21035 (N_21035,N_16925,N_15782);
nand U21036 (N_21036,N_17749,N_17351);
nand U21037 (N_21037,N_18790,N_17693);
or U21038 (N_21038,N_16351,N_17851);
or U21039 (N_21039,N_17204,N_18760);
nand U21040 (N_21040,N_18570,N_15735);
nor U21041 (N_21041,N_18146,N_17266);
nand U21042 (N_21042,N_16226,N_17364);
and U21043 (N_21043,N_15922,N_17065);
xnor U21044 (N_21044,N_15311,N_18785);
nor U21045 (N_21045,N_16279,N_18013);
nor U21046 (N_21046,N_19413,N_17268);
nand U21047 (N_21047,N_16409,N_18688);
nor U21048 (N_21048,N_16500,N_17596);
nor U21049 (N_21049,N_15299,N_15916);
nor U21050 (N_21050,N_17216,N_16093);
and U21051 (N_21051,N_18907,N_15832);
nand U21052 (N_21052,N_19098,N_16867);
nand U21053 (N_21053,N_16058,N_17974);
or U21054 (N_21054,N_16313,N_15690);
nand U21055 (N_21055,N_19219,N_19403);
nand U21056 (N_21056,N_15042,N_15915);
and U21057 (N_21057,N_17231,N_18259);
nand U21058 (N_21058,N_17237,N_15542);
nand U21059 (N_21059,N_16458,N_16773);
nor U21060 (N_21060,N_19582,N_15267);
nand U21061 (N_21061,N_19335,N_18670);
nor U21062 (N_21062,N_16734,N_18122);
nor U21063 (N_21063,N_17436,N_16356);
nand U21064 (N_21064,N_15292,N_17706);
xor U21065 (N_21065,N_16151,N_19876);
nand U21066 (N_21066,N_18701,N_19478);
or U21067 (N_21067,N_18482,N_19749);
xnor U21068 (N_21068,N_19169,N_19398);
nor U21069 (N_21069,N_15210,N_16055);
nand U21070 (N_21070,N_15708,N_17174);
or U21071 (N_21071,N_16585,N_19490);
nand U21072 (N_21072,N_15912,N_15421);
and U21073 (N_21073,N_15067,N_19217);
or U21074 (N_21074,N_16737,N_16596);
or U21075 (N_21075,N_19579,N_18786);
nor U21076 (N_21076,N_18742,N_16345);
or U21077 (N_21077,N_15728,N_16013);
and U21078 (N_21078,N_17426,N_15654);
nor U21079 (N_21079,N_17770,N_16860);
or U21080 (N_21080,N_18474,N_19765);
nand U21081 (N_21081,N_18583,N_16047);
and U21082 (N_21082,N_19348,N_19934);
or U21083 (N_21083,N_16523,N_18941);
nor U21084 (N_21084,N_16007,N_17876);
nand U21085 (N_21085,N_15031,N_17670);
or U21086 (N_21086,N_15560,N_19511);
or U21087 (N_21087,N_17962,N_15564);
or U21088 (N_21088,N_17155,N_16864);
nor U21089 (N_21089,N_15737,N_15740);
nand U21090 (N_21090,N_15068,N_17202);
nand U21091 (N_21091,N_16367,N_16469);
nor U21092 (N_21092,N_18691,N_17737);
or U21093 (N_21093,N_16437,N_19300);
and U21094 (N_21094,N_15302,N_17621);
or U21095 (N_21095,N_18185,N_18132);
nor U21096 (N_21096,N_19881,N_19664);
xnor U21097 (N_21097,N_18321,N_17861);
nor U21098 (N_21098,N_19179,N_18502);
or U21099 (N_21099,N_18011,N_16197);
and U21100 (N_21100,N_15882,N_19706);
xor U21101 (N_21101,N_19113,N_16300);
nand U21102 (N_21102,N_17119,N_18023);
and U21103 (N_21103,N_16135,N_15685);
or U21104 (N_21104,N_15967,N_17134);
or U21105 (N_21105,N_16571,N_16653);
nor U21106 (N_21106,N_15187,N_16049);
nor U21107 (N_21107,N_19422,N_15387);
and U21108 (N_21108,N_15711,N_18833);
nand U21109 (N_21109,N_19107,N_16449);
and U21110 (N_21110,N_17620,N_19091);
nand U21111 (N_21111,N_17688,N_17524);
nand U21112 (N_21112,N_16790,N_16164);
and U21113 (N_21113,N_17891,N_17371);
or U21114 (N_21114,N_15628,N_17625);
nor U21115 (N_21115,N_18619,N_15175);
xor U21116 (N_21116,N_15164,N_16399);
nor U21117 (N_21117,N_19387,N_19850);
nand U21118 (N_21118,N_15190,N_17254);
xor U21119 (N_21119,N_15288,N_18986);
and U21120 (N_21120,N_16274,N_16183);
xor U21121 (N_21121,N_18489,N_18432);
or U21122 (N_21122,N_19365,N_18317);
and U21123 (N_21123,N_16037,N_18650);
or U21124 (N_21124,N_18955,N_15347);
nand U21125 (N_21125,N_17154,N_15238);
xnor U21126 (N_21126,N_19384,N_19707);
nor U21127 (N_21127,N_18764,N_18430);
nor U21128 (N_21128,N_15757,N_19460);
and U21129 (N_21129,N_15816,N_19488);
or U21130 (N_21130,N_18639,N_17580);
or U21131 (N_21131,N_15661,N_16161);
nand U21132 (N_21132,N_18529,N_18596);
nand U21133 (N_21133,N_19904,N_18076);
and U21134 (N_21134,N_18320,N_16650);
nor U21135 (N_21135,N_19784,N_16855);
or U21136 (N_21136,N_17570,N_18176);
nor U21137 (N_21137,N_18973,N_15234);
nand U21138 (N_21138,N_15390,N_19439);
nand U21139 (N_21139,N_18974,N_16090);
nor U21140 (N_21140,N_18270,N_19957);
or U21141 (N_21141,N_19726,N_19080);
and U21142 (N_21142,N_15444,N_15738);
and U21143 (N_21143,N_16059,N_19886);
and U21144 (N_21144,N_17465,N_18847);
or U21145 (N_21145,N_16996,N_18846);
nor U21146 (N_21146,N_18134,N_16957);
or U21147 (N_21147,N_15439,N_18979);
and U21148 (N_21148,N_19137,N_16364);
nand U21149 (N_21149,N_19031,N_19174);
and U21150 (N_21150,N_18478,N_15604);
and U21151 (N_21151,N_18026,N_19998);
and U21152 (N_21152,N_16427,N_19286);
or U21153 (N_21153,N_15507,N_19791);
nor U21154 (N_21154,N_15132,N_16985);
nor U21155 (N_21155,N_17606,N_18667);
nand U21156 (N_21156,N_16334,N_16896);
nand U21157 (N_21157,N_18939,N_15077);
nand U21158 (N_21158,N_16674,N_17904);
nand U21159 (N_21159,N_15558,N_17333);
and U21160 (N_21160,N_18369,N_16031);
nand U21161 (N_21161,N_15039,N_17305);
xor U21162 (N_21162,N_15134,N_16467);
nor U21163 (N_21163,N_18021,N_15087);
and U21164 (N_21164,N_16142,N_15878);
nor U21165 (N_21165,N_17924,N_18969);
nor U21166 (N_21166,N_18431,N_16926);
nand U21167 (N_21167,N_18221,N_15147);
nand U21168 (N_21168,N_16736,N_19046);
nor U21169 (N_21169,N_17013,N_16422);
nor U21170 (N_21170,N_16310,N_17521);
or U21171 (N_21171,N_18961,N_18690);
and U21172 (N_21172,N_18446,N_15182);
or U21173 (N_21173,N_19164,N_15342);
and U21174 (N_21174,N_17980,N_18686);
or U21175 (N_21175,N_16139,N_15614);
or U21176 (N_21176,N_18102,N_17410);
nor U21177 (N_21177,N_19837,N_16927);
nor U21178 (N_21178,N_15758,N_17903);
nor U21179 (N_21179,N_19949,N_18256);
and U21180 (N_21180,N_16244,N_16222);
nand U21181 (N_21181,N_19780,N_18015);
or U21182 (N_21182,N_16693,N_18585);
or U21183 (N_21183,N_16205,N_17894);
nor U21184 (N_21184,N_15736,N_18156);
or U21185 (N_21185,N_15580,N_19280);
nand U21186 (N_21186,N_16299,N_17850);
nor U21187 (N_21187,N_15050,N_19399);
or U21188 (N_21188,N_19556,N_15392);
or U21189 (N_21189,N_16921,N_15821);
nand U21190 (N_21190,N_15359,N_17982);
nor U21191 (N_21191,N_19212,N_16801);
nor U21192 (N_21192,N_19463,N_19449);
nand U21193 (N_21193,N_19134,N_18406);
or U21194 (N_21194,N_17077,N_16646);
or U21195 (N_21195,N_15682,N_16287);
nor U21196 (N_21196,N_18244,N_17234);
nor U21197 (N_21197,N_17353,N_18426);
nor U21198 (N_21198,N_16712,N_19148);
nand U21199 (N_21199,N_15778,N_17322);
and U21200 (N_21200,N_17515,N_19220);
nand U21201 (N_21201,N_16141,N_17898);
nor U21202 (N_21202,N_17875,N_16506);
and U21203 (N_21203,N_16115,N_16069);
and U21204 (N_21204,N_19191,N_19411);
and U21205 (N_21205,N_19856,N_15502);
nand U21206 (N_21206,N_18655,N_18704);
nand U21207 (N_21207,N_19965,N_16154);
nand U21208 (N_21208,N_18360,N_16483);
nor U21209 (N_21209,N_16593,N_18153);
and U21210 (N_21210,N_16915,N_17103);
nor U21211 (N_21211,N_16850,N_18473);
and U21212 (N_21212,N_18287,N_19544);
or U21213 (N_21213,N_18797,N_18152);
nor U21214 (N_21214,N_17142,N_17771);
and U21215 (N_21215,N_18238,N_18273);
or U21216 (N_21216,N_16844,N_15287);
and U21217 (N_21217,N_19662,N_19097);
and U21218 (N_21218,N_16976,N_18372);
and U21219 (N_21219,N_15814,N_16871);
or U21220 (N_21220,N_19033,N_19986);
xor U21221 (N_21221,N_16140,N_18274);
nor U21222 (N_21222,N_18738,N_18647);
nor U21223 (N_21223,N_19353,N_18996);
nor U21224 (N_21224,N_18520,N_16240);
nand U21225 (N_21225,N_18866,N_16876);
xor U21226 (N_21226,N_17182,N_16143);
or U21227 (N_21227,N_17141,N_16787);
nor U21228 (N_21228,N_16455,N_17045);
and U21229 (N_21229,N_15602,N_19173);
nand U21230 (N_21230,N_17201,N_17882);
or U21231 (N_21231,N_17367,N_19816);
and U21232 (N_21232,N_18988,N_19793);
and U21233 (N_21233,N_18351,N_19616);
nand U21234 (N_21234,N_15718,N_17153);
or U21235 (N_21235,N_15576,N_17443);
and U21236 (N_21236,N_15568,N_19855);
and U21237 (N_21237,N_18795,N_18261);
nand U21238 (N_21238,N_16066,N_17734);
nand U21239 (N_21239,N_17790,N_17467);
nand U21240 (N_21240,N_15363,N_15932);
or U21241 (N_21241,N_17868,N_19154);
nand U21242 (N_21242,N_18648,N_18525);
nor U21243 (N_21243,N_18615,N_19925);
nor U21244 (N_21244,N_16092,N_15023);
nor U21245 (N_21245,N_16894,N_16805);
nor U21246 (N_21246,N_16019,N_18159);
or U21247 (N_21247,N_15936,N_18119);
or U21248 (N_21248,N_19301,N_17925);
nand U21249 (N_21249,N_17585,N_18634);
nor U21250 (N_21250,N_15118,N_18578);
nor U21251 (N_21251,N_16231,N_15559);
nor U21252 (N_21252,N_16368,N_15994);
nand U21253 (N_21253,N_17838,N_16326);
nor U21254 (N_21254,N_15824,N_17279);
nor U21255 (N_21255,N_15514,N_18703);
nand U21256 (N_21256,N_18487,N_18403);
or U21257 (N_21257,N_19721,N_18236);
or U21258 (N_21258,N_18086,N_18882);
and U21259 (N_21259,N_19186,N_17548);
nand U21260 (N_21260,N_17495,N_19547);
or U21261 (N_21261,N_17937,N_18355);
xor U21262 (N_21262,N_19486,N_16694);
nor U21263 (N_21263,N_16378,N_18632);
nand U21264 (N_21264,N_17092,N_18538);
nand U21265 (N_21265,N_18439,N_16330);
or U21266 (N_21266,N_18145,N_19880);
nor U21267 (N_21267,N_19803,N_16491);
or U21268 (N_21268,N_17225,N_19896);
nor U21269 (N_21269,N_15006,N_15911);
nor U21270 (N_21270,N_15947,N_17362);
and U21271 (N_21271,N_16208,N_17747);
and U21272 (N_21272,N_16881,N_18942);
nand U21273 (N_21273,N_19843,N_19458);
and U21274 (N_21274,N_15317,N_15871);
and U21275 (N_21275,N_18700,N_15594);
or U21276 (N_21276,N_17361,N_18410);
xor U21277 (N_21277,N_15020,N_19601);
or U21278 (N_21278,N_15002,N_16414);
nor U21279 (N_21279,N_19224,N_15945);
or U21280 (N_21280,N_19847,N_16045);
nor U21281 (N_21281,N_15283,N_19875);
xor U21282 (N_21282,N_16319,N_18399);
nor U21283 (N_21283,N_16688,N_17459);
nand U21284 (N_21284,N_17464,N_18315);
nand U21285 (N_21285,N_16375,N_16785);
nand U21286 (N_21286,N_19231,N_15839);
nor U21287 (N_21287,N_16346,N_19208);
or U21288 (N_21288,N_16246,N_19341);
or U21289 (N_21289,N_16625,N_18249);
nor U21290 (N_21290,N_15041,N_15053);
nor U21291 (N_21291,N_16050,N_16099);
and U21292 (N_21292,N_17870,N_15714);
and U21293 (N_21293,N_19261,N_19176);
nor U21294 (N_21294,N_15013,N_17037);
nand U21295 (N_21295,N_17075,N_18313);
xnor U21296 (N_21296,N_18543,N_16179);
or U21297 (N_21297,N_18516,N_15848);
or U21298 (N_21298,N_15410,N_16863);
or U21299 (N_21299,N_17264,N_15211);
nor U21300 (N_21300,N_19183,N_18398);
nor U21301 (N_21301,N_17604,N_17854);
and U21302 (N_21302,N_15014,N_17730);
nor U21303 (N_21303,N_16710,N_17329);
and U21304 (N_21304,N_19388,N_16377);
nand U21305 (N_21305,N_17642,N_15913);
nor U21306 (N_21306,N_15826,N_16472);
xor U21307 (N_21307,N_16731,N_17638);
and U21308 (N_21308,N_15929,N_16479);
nor U21309 (N_21309,N_16997,N_18420);
nor U21310 (N_21310,N_15581,N_16407);
nand U21311 (N_21311,N_19936,N_15906);
or U21312 (N_21312,N_15724,N_19879);
or U21313 (N_21313,N_19539,N_17057);
and U21314 (N_21314,N_19745,N_15918);
nor U21315 (N_21315,N_17453,N_19971);
nand U21316 (N_21316,N_18644,N_19798);
nor U21317 (N_21317,N_16029,N_19118);
nand U21318 (N_21318,N_15879,N_16234);
nor U21319 (N_21319,N_17834,N_15903);
nor U21320 (N_21320,N_18056,N_17339);
or U21321 (N_21321,N_16845,N_18350);
and U21322 (N_21322,N_19367,N_18285);
and U21323 (N_21323,N_16933,N_15588);
nand U21324 (N_21324,N_19787,N_19391);
or U21325 (N_21325,N_17501,N_19433);
nand U21326 (N_21326,N_19379,N_17331);
nand U21327 (N_21327,N_17872,N_16770);
or U21328 (N_21328,N_16250,N_17779);
xor U21329 (N_21329,N_19615,N_19157);
nor U21330 (N_21330,N_15160,N_16610);
nand U21331 (N_21331,N_19994,N_16315);
or U21332 (N_21332,N_18812,N_17066);
and U21333 (N_21333,N_19585,N_16998);
or U21334 (N_21334,N_19155,N_15030);
nand U21335 (N_21335,N_16233,N_15344);
nand U21336 (N_21336,N_18837,N_15631);
and U21337 (N_21337,N_16438,N_17721);
xnor U21338 (N_21338,N_17014,N_17276);
and U21339 (N_21339,N_15995,N_16902);
nand U21340 (N_21340,N_16979,N_17588);
nand U21341 (N_21341,N_17574,N_18778);
nand U21342 (N_21342,N_18588,N_17354);
nor U21343 (N_21343,N_17796,N_15179);
xnor U21344 (N_21344,N_19267,N_18488);
nand U21345 (N_21345,N_17398,N_18933);
nor U21346 (N_21346,N_15388,N_17441);
nor U21347 (N_21347,N_18177,N_17915);
nor U21348 (N_21348,N_19328,N_19967);
nand U21349 (N_21349,N_18546,N_16668);
and U21350 (N_21350,N_19051,N_17146);
or U21351 (N_21351,N_19677,N_17654);
xor U21352 (N_21352,N_18950,N_16757);
and U21353 (N_21353,N_17899,N_16402);
nor U21354 (N_21354,N_17076,N_17420);
nor U21355 (N_21355,N_16374,N_17180);
or U21356 (N_21356,N_15282,N_19457);
nand U21357 (N_21357,N_19723,N_19099);
or U21358 (N_21358,N_19680,N_16882);
and U21359 (N_21359,N_19368,N_15622);
nand U21360 (N_21360,N_19343,N_19525);
and U21361 (N_21361,N_15278,N_15273);
and U21362 (N_21362,N_18254,N_18227);
or U21363 (N_21363,N_15391,N_17680);
and U21364 (N_21364,N_19572,N_18211);
and U21365 (N_21365,N_17555,N_19781);
and U21366 (N_21366,N_17878,N_17388);
nor U21367 (N_21367,N_16828,N_18251);
or U21368 (N_21368,N_15131,N_15011);
and U21369 (N_21369,N_15772,N_18563);
and U21370 (N_21370,N_17679,N_17554);
and U21371 (N_21371,N_19557,N_18702);
nand U21372 (N_21372,N_17341,N_16238);
nand U21373 (N_21373,N_17286,N_18840);
and U21374 (N_21374,N_15973,N_19382);
or U21375 (N_21375,N_16875,N_19499);
or U21376 (N_21376,N_16456,N_15271);
and U21377 (N_21377,N_19266,N_17430);
nor U21378 (N_21378,N_16366,N_18966);
nand U21379 (N_21379,N_17048,N_17235);
and U21380 (N_21380,N_17858,N_19069);
nor U21381 (N_21381,N_18264,N_15697);
and U21382 (N_21382,N_15645,N_19255);
nand U21383 (N_21383,N_19279,N_17826);
nor U21384 (N_21384,N_17836,N_19958);
xor U21385 (N_21385,N_18744,N_18204);
nor U21386 (N_21386,N_17881,N_16846);
xor U21387 (N_21387,N_17258,N_17990);
nor U21388 (N_21388,N_15263,N_18510);
nor U21389 (N_21389,N_19895,N_18814);
nor U21390 (N_21390,N_15016,N_17412);
nor U21391 (N_21391,N_18139,N_19392);
nand U21392 (N_21392,N_18206,N_15979);
nand U21393 (N_21393,N_18878,N_18908);
and U21394 (N_21394,N_17070,N_17281);
nand U21395 (N_21395,N_16781,N_15650);
and U21396 (N_21396,N_15490,N_15619);
nand U21397 (N_21397,N_16094,N_17236);
and U21398 (N_21398,N_16936,N_19029);
and U21399 (N_21399,N_16791,N_15135);
nand U21400 (N_21400,N_17517,N_18107);
nand U21401 (N_21401,N_16960,N_15057);
nor U21402 (N_21402,N_18964,N_18834);
nor U21403 (N_21403,N_17043,N_15261);
and U21404 (N_21404,N_19618,N_16303);
or U21405 (N_21405,N_17429,N_19635);
nand U21406 (N_21406,N_15652,N_16671);
nor U21407 (N_21407,N_18936,N_19870);
or U21408 (N_21408,N_16928,N_18378);
nor U21409 (N_21409,N_19077,N_16504);
and U21410 (N_21410,N_18064,N_15003);
nor U21411 (N_21411,N_18853,N_19166);
and U21412 (N_21412,N_17170,N_15372);
nor U21413 (N_21413,N_19295,N_16492);
nand U21414 (N_21414,N_19418,N_19771);
and U21415 (N_21415,N_16956,N_18879);
nand U21416 (N_21416,N_19005,N_19529);
xnor U21417 (N_21417,N_16662,N_17956);
and U21418 (N_21418,N_15494,N_18255);
xor U21419 (N_21419,N_16725,N_17448);
and U21420 (N_21420,N_18123,N_17575);
nor U21421 (N_21421,N_19450,N_17643);
or U21422 (N_21422,N_19633,N_18549);
nor U21423 (N_21423,N_16323,N_19424);
xor U21424 (N_21424,N_18442,N_16320);
or U21425 (N_21425,N_16360,N_18621);
and U21426 (N_21426,N_15706,N_18851);
nand U21427 (N_21427,N_19260,N_19961);
xnor U21428 (N_21428,N_19946,N_15539);
or U21429 (N_21429,N_15598,N_19708);
and U21430 (N_21430,N_15148,N_16633);
and U21431 (N_21431,N_17835,N_15434);
or U21432 (N_21432,N_15638,N_19024);
or U21433 (N_21433,N_16420,N_19898);
or U21434 (N_21434,N_17677,N_18300);
nand U21435 (N_21435,N_15659,N_15827);
and U21436 (N_21436,N_18084,N_18422);
nor U21437 (N_21437,N_15408,N_18712);
nor U21438 (N_21438,N_17761,N_17018);
or U21439 (N_21439,N_15853,N_17176);
and U21440 (N_21440,N_15767,N_15895);
nor U21441 (N_21441,N_15719,N_17842);
or U21442 (N_21442,N_16542,N_16332);
or U21443 (N_21443,N_15655,N_19939);
and U21444 (N_21444,N_16641,N_18186);
xor U21445 (N_21445,N_16130,N_16592);
or U21446 (N_21446,N_17611,N_18531);
and U21447 (N_21447,N_18989,N_16532);
and U21448 (N_21448,N_18133,N_15914);
nand U21449 (N_21449,N_17460,N_15804);
or U21450 (N_21450,N_16795,N_19767);
and U21451 (N_21451,N_19920,N_16518);
nand U21452 (N_21452,N_15338,N_19766);
or U21453 (N_21453,N_19497,N_15552);
or U21454 (N_21454,N_15715,N_18754);
nand U21455 (N_21455,N_19018,N_17740);
or U21456 (N_21456,N_17617,N_18068);
nor U21457 (N_21457,N_17227,N_17126);
nor U21458 (N_21458,N_17480,N_18633);
nand U21459 (N_21459,N_18087,N_15000);
or U21460 (N_21460,N_16862,N_18241);
or U21461 (N_21461,N_16148,N_17640);
or U21462 (N_21462,N_15550,N_15861);
or U21463 (N_21463,N_16361,N_15036);
nand U21464 (N_21464,N_18304,N_15783);
nor U21465 (N_21465,N_18257,N_16193);
or U21466 (N_21466,N_19882,N_18766);
nand U21467 (N_21467,N_16852,N_17032);
xor U21468 (N_21468,N_19314,N_16331);
nor U21469 (N_21469,N_15061,N_19483);
or U21470 (N_21470,N_16337,N_16176);
or U21471 (N_21471,N_18309,N_18953);
nor U21472 (N_21472,N_18128,N_18721);
nand U21473 (N_21473,N_15570,N_18565);
or U21474 (N_21474,N_16916,N_17914);
and U21475 (N_21475,N_18262,N_17086);
and U21476 (N_21476,N_15793,N_15524);
nand U21477 (N_21477,N_16383,N_16493);
nor U21478 (N_21478,N_15972,N_19323);
or U21479 (N_21479,N_19476,N_17635);
or U21480 (N_21480,N_15625,N_18042);
nand U21481 (N_21481,N_15545,N_16893);
nand U21482 (N_21482,N_18397,N_18126);
nor U21483 (N_21483,N_17577,N_16018);
nand U21484 (N_21484,N_17626,N_18165);
nand U21485 (N_21485,N_18521,N_17278);
nor U21486 (N_21486,N_15870,N_16679);
nor U21487 (N_21487,N_16153,N_19188);
nand U21488 (N_21488,N_16448,N_15589);
or U21489 (N_21489,N_17290,N_19666);
and U21490 (N_21490,N_18401,N_19884);
and U21491 (N_21491,N_16779,N_16961);
nor U21492 (N_21492,N_17125,N_18411);
or U21493 (N_21493,N_19406,N_15726);
and U21494 (N_21494,N_16879,N_19468);
and U21495 (N_21495,N_17382,N_16705);
nand U21496 (N_21496,N_17449,N_19889);
nand U21497 (N_21497,N_16098,N_19240);
and U21498 (N_21498,N_15251,N_17792);
and U21499 (N_21499,N_16223,N_17844);
nor U21500 (N_21500,N_19063,N_16608);
nor U21501 (N_21501,N_16950,N_15201);
and U21502 (N_21502,N_18598,N_19239);
or U21503 (N_21503,N_15323,N_19806);
nand U21504 (N_21504,N_18844,N_18091);
nor U21505 (N_21505,N_16156,N_15236);
nor U21506 (N_21506,N_17853,N_16967);
or U21507 (N_21507,N_16892,N_15819);
and U21508 (N_21508,N_15417,N_18242);
nor U21509 (N_21509,N_18924,N_17886);
or U21510 (N_21510,N_18587,N_16760);
or U21511 (N_21511,N_16833,N_19571);
and U21512 (N_21512,N_15673,N_17913);
or U21513 (N_21513,N_17041,N_17910);
nand U21514 (N_21514,N_19638,N_17393);
nor U21515 (N_21515,N_15250,N_19710);
or U21516 (N_21516,N_19495,N_17944);
and U21517 (N_21517,N_17152,N_15828);
or U21518 (N_21518,N_19223,N_15679);
and U21519 (N_21519,N_19053,N_15491);
and U21520 (N_21520,N_15667,N_18444);
nand U21521 (N_21521,N_16800,N_19893);
or U21522 (N_21522,N_18519,N_19654);
nor U21523 (N_21523,N_15572,N_15296);
or U21524 (N_21524,N_17417,N_19631);
and U21525 (N_21525,N_19416,N_18898);
nand U21526 (N_21526,N_16793,N_16943);
and U21527 (N_21527,N_17631,N_15114);
nor U21528 (N_21528,N_19471,N_19313);
or U21529 (N_21529,N_15221,N_16376);
nand U21530 (N_21530,N_17061,N_18138);
nand U21531 (N_21531,N_18716,N_15257);
nand U21532 (N_21532,N_17600,N_16898);
nand U21533 (N_21533,N_17681,N_17957);
or U21534 (N_21534,N_15396,N_18946);
and U21535 (N_21535,N_15894,N_15785);
and U21536 (N_21536,N_16269,N_18316);
nand U21537 (N_21537,N_18747,N_16133);
or U21538 (N_21538,N_15658,N_19143);
nor U21539 (N_21539,N_18909,N_15596);
and U21540 (N_21540,N_17686,N_19380);
and U21541 (N_21541,N_17482,N_19775);
nand U21542 (N_21542,N_16565,N_19573);
nor U21543 (N_21543,N_15090,N_17831);
nand U21544 (N_21544,N_18438,N_17181);
or U21545 (N_21545,N_16369,N_18889);
nor U21546 (N_21546,N_15070,N_16229);
nor U21547 (N_21547,N_16401,N_15145);
or U21548 (N_21548,N_16516,N_17532);
and U21549 (N_21549,N_16322,N_16419);
xnor U21550 (N_21550,N_15864,N_18103);
xnor U21551 (N_21551,N_19560,N_18515);
and U21552 (N_21552,N_17840,N_15569);
xor U21553 (N_21553,N_17726,N_16552);
nor U21554 (N_21554,N_16439,N_17198);
and U21555 (N_21555,N_17800,N_17177);
nor U21556 (N_21556,N_19247,N_15566);
and U21557 (N_21557,N_17413,N_15415);
or U21558 (N_21558,N_15928,N_19050);
or U21559 (N_21559,N_18216,N_19299);
and U21560 (N_21560,N_15012,N_19985);
nor U21561 (N_21561,N_17499,N_18836);
nand U21562 (N_21562,N_17519,N_16196);
nor U21563 (N_21563,N_16227,N_19897);
or U21564 (N_21564,N_17707,N_15926);
nor U21565 (N_21565,N_18699,N_18755);
nor U21566 (N_21566,N_16678,N_15942);
nand U21567 (N_21567,N_18804,N_16503);
and U21568 (N_21568,N_18589,N_16225);
nor U21569 (N_21569,N_18115,N_18558);
nand U21570 (N_21570,N_19951,N_19799);
nor U21571 (N_21571,N_16822,N_17651);
and U21572 (N_21572,N_15088,N_15229);
nand U21573 (N_21573,N_18059,N_18100);
nor U21574 (N_21574,N_16614,N_15644);
nand U21575 (N_21575,N_16129,N_18660);
and U21576 (N_21576,N_17936,N_19608);
or U21577 (N_21577,N_18448,N_15418);
or U21578 (N_21578,N_15348,N_18237);
and U21579 (N_21579,N_17299,N_15243);
and U21580 (N_21580,N_18784,N_18976);
or U21581 (N_21581,N_15680,N_19562);
nor U21582 (N_21582,N_15875,N_17130);
nand U21583 (N_21583,N_17646,N_17981);
nand U21584 (N_21584,N_19687,N_19001);
nand U21585 (N_21585,N_16558,N_16922);
or U21586 (N_21586,N_19447,N_18535);
and U21587 (N_21587,N_16087,N_17542);
or U21588 (N_21588,N_16224,N_15851);
nor U21589 (N_21589,N_16305,N_19309);
or U21590 (N_21590,N_15356,N_16510);
nand U21591 (N_21591,N_16081,N_16522);
or U21592 (N_21592,N_17136,N_18616);
or U21593 (N_21593,N_15739,N_17933);
or U21594 (N_21594,N_19158,N_17841);
and U21595 (N_21595,N_16741,N_17711);
or U21596 (N_21596,N_16292,N_15293);
or U21597 (N_21597,N_17300,N_18967);
nand U21598 (N_21598,N_19914,N_18465);
or U21599 (N_21599,N_17813,N_18881);
nand U21600 (N_21600,N_16859,N_16765);
or U21601 (N_21601,N_19209,N_16030);
and U21602 (N_21602,N_15541,N_16266);
or U21603 (N_21603,N_15153,N_19899);
nor U21604 (N_21604,N_18464,N_17996);
or U21605 (N_21605,N_17503,N_17633);
and U21606 (N_21606,N_15695,N_19444);
or U21607 (N_21607,N_17942,N_17823);
nand U21608 (N_21608,N_16843,N_16243);
or U21609 (N_21609,N_17017,N_18617);
or U21610 (N_21610,N_17208,N_19501);
or U21611 (N_21611,N_19339,N_15750);
nand U21612 (N_21612,N_17786,N_18299);
and U21613 (N_21613,N_15121,N_18038);
nor U21614 (N_21614,N_17658,N_15399);
nand U21615 (N_21615,N_19537,N_18977);
nor U21616 (N_21616,N_19824,N_16564);
and U21617 (N_21617,N_15154,N_18070);
or U21618 (N_21618,N_18335,N_18246);
nor U21619 (N_21619,N_15760,N_17793);
nor U21620 (N_21620,N_16276,N_19036);
nand U21621 (N_21621,N_16604,N_17559);
nand U21622 (N_21622,N_19487,N_15773);
and U21623 (N_21623,N_18007,N_18170);
and U21624 (N_21624,N_17139,N_19812);
nand U21625 (N_21625,N_18392,N_16121);
or U21626 (N_21626,N_17801,N_18045);
and U21627 (N_21627,N_18469,N_15669);
nor U21628 (N_21628,N_18586,N_16642);
nor U21629 (N_21629,N_16213,N_17285);
nand U21630 (N_21630,N_15516,N_19283);
nand U21631 (N_21631,N_17534,N_19694);
nor U21632 (N_21632,N_16537,N_18483);
and U21633 (N_21633,N_16637,N_16218);
or U21634 (N_21634,N_19202,N_19089);
and U21635 (N_21635,N_19329,N_18462);
and U21636 (N_21636,N_19873,N_17275);
nor U21637 (N_21637,N_16291,N_19070);
nand U21638 (N_21638,N_15219,N_15902);
or U21639 (N_21639,N_18913,N_16145);
and U21640 (N_21640,N_15722,N_15150);
nor U21641 (N_21641,N_18666,N_19170);
and U21642 (N_21642,N_17992,N_15469);
and U21643 (N_21643,N_17309,N_19479);
and U21644 (N_21644,N_18112,N_16435);
xor U21645 (N_21645,N_15451,N_19037);
and U21646 (N_21646,N_15866,N_16615);
nand U21647 (N_21647,N_18314,N_16577);
nand U21648 (N_21648,N_19109,N_18547);
or U21649 (N_21649,N_17022,N_19232);
nand U21650 (N_21650,N_16088,N_19105);
nand U21651 (N_21651,N_15449,N_15686);
nand U21652 (N_21652,N_16461,N_15280);
or U21653 (N_21653,N_18808,N_19119);
or U21654 (N_21654,N_17708,N_19838);
or U21655 (N_21655,N_17892,N_17863);
or U21656 (N_21656,N_19697,N_15959);
nand U21657 (N_21657,N_18550,N_18069);
nor U21658 (N_21658,N_18074,N_19211);
nand U21659 (N_21659,N_16697,N_15122);
and U21660 (N_21660,N_15329,N_18370);
and U21661 (N_21661,N_19968,N_15173);
nand U21662 (N_21662,N_18065,N_18734);
nand U21663 (N_21663,N_17138,N_18000);
nand U21664 (N_21664,N_18622,N_18998);
nor U21665 (N_21665,N_16907,N_17492);
and U21666 (N_21666,N_15397,N_17158);
nor U21667 (N_21667,N_19565,N_19115);
or U21668 (N_21668,N_15353,N_17783);
and U21669 (N_21669,N_19443,N_17470);
nand U21670 (N_21670,N_18557,N_16349);
nand U21671 (N_21671,N_15094,N_16908);
nor U21672 (N_21672,N_17200,N_17941);
and U21673 (N_21673,N_19200,N_15025);
nand U21674 (N_21674,N_15373,N_19108);
and U21675 (N_21675,N_16554,N_15235);
nand U21676 (N_21676,N_15319,N_18805);
or U21677 (N_21677,N_18694,N_17855);
nor U21678 (N_21678,N_16187,N_17762);
or U21679 (N_21679,N_19445,N_17928);
and U21680 (N_21680,N_15670,N_16288);
nand U21681 (N_21681,N_17221,N_19992);
or U21682 (N_21682,N_19257,N_18143);
or U21683 (N_21683,N_16103,N_18912);
or U21684 (N_21684,N_18348,N_17587);
or U21685 (N_21685,N_19417,N_17880);
nor U21686 (N_21686,N_17550,N_17694);
and U21687 (N_21687,N_15616,N_17280);
nand U21688 (N_21688,N_16175,N_17486);
nand U21689 (N_21689,N_15483,N_18975);
and U21690 (N_21690,N_16849,N_16298);
or U21691 (N_21691,N_19944,N_16707);
nor U21692 (N_21692,N_18732,N_17808);
or U21693 (N_21693,N_19724,N_15108);
nand U21694 (N_21694,N_16575,N_16606);
and U21695 (N_21695,N_16436,N_16966);
and U21696 (N_21696,N_16311,N_19052);
and U21697 (N_21697,N_16181,N_19712);
nor U21698 (N_21698,N_15139,N_18664);
and U21699 (N_21699,N_19492,N_18569);
nand U21700 (N_21700,N_15984,N_15393);
or U21701 (N_21701,N_15505,N_15047);
nor U21702 (N_21702,N_16237,N_17261);
and U21703 (N_21703,N_19794,N_19149);
nand U21704 (N_21704,N_19959,N_15370);
nand U21705 (N_21705,N_17594,N_19714);
nand U21706 (N_21706,N_18358,N_15314);
and U21707 (N_21707,N_18629,N_16764);
and U21708 (N_21708,N_19650,N_15702);
and U21709 (N_21709,N_19306,N_18675);
xnor U21710 (N_21710,N_15498,N_18864);
nand U21711 (N_21711,N_17145,N_15687);
or U21712 (N_21712,N_17901,N_15008);
or U21713 (N_21713,N_17954,N_17667);
or U21714 (N_21714,N_16780,N_15321);
nand U21715 (N_21715,N_16074,N_19205);
and U21716 (N_21716,N_16384,N_19748);
and U21717 (N_21717,N_19235,N_18269);
or U21718 (N_21718,N_15834,N_19960);
nand U21719 (N_21719,N_16333,N_15034);
nor U21720 (N_21720,N_15597,N_16421);
and U21721 (N_21721,N_19732,N_17498);
or U21722 (N_21722,N_17733,N_15537);
or U21723 (N_21723,N_16804,N_17601);
and U21724 (N_21724,N_15225,N_15904);
or U21725 (N_21725,N_19124,N_16703);
nand U21726 (N_21726,N_16114,N_16391);
and U21727 (N_21727,N_16603,N_17115);
and U21728 (N_21728,N_15846,N_17108);
or U21729 (N_21729,N_19442,N_19305);
nor U21730 (N_21730,N_16057,N_19400);
nand U21731 (N_21731,N_16794,N_19810);
nor U21732 (N_21732,N_18739,N_19570);
and U21733 (N_21733,N_17682,N_17406);
and U21734 (N_21734,N_17743,N_16204);
or U21735 (N_21735,N_15709,N_18919);
and U21736 (N_21736,N_17716,N_17469);
or U21737 (N_21737,N_16623,N_16945);
nor U21738 (N_21738,N_18762,N_17795);
nand U21739 (N_21739,N_15765,N_16878);
nand U21740 (N_21740,N_19844,N_15617);
nor U21741 (N_21741,N_18200,N_17883);
or U21742 (N_21742,N_17884,N_19670);
and U21743 (N_21743,N_19081,N_18581);
and U21744 (N_21744,N_18925,N_19349);
or U21745 (N_21745,N_18030,N_15209);
nand U21746 (N_21746,N_15964,N_16511);
or U21747 (N_21747,N_18499,N_15934);
and U21748 (N_21748,N_19990,N_16207);
or U21749 (N_21749,N_17978,N_19133);
and U21750 (N_21750,N_15463,N_15847);
nor U21751 (N_21751,N_18484,N_18658);
nor U21752 (N_21752,N_16400,N_17478);
or U21753 (N_21753,N_19013,N_18613);
nand U21754 (N_21754,N_18855,N_18234);
or U21755 (N_21755,N_16411,N_19676);
nand U21756 (N_21756,N_15368,N_18665);
nor U21757 (N_21757,N_15093,N_17178);
xor U21758 (N_21758,N_19667,N_17296);
or U21759 (N_21759,N_16316,N_18963);
nand U21760 (N_21760,N_18923,N_15720);
or U21761 (N_21761,N_17265,N_18532);
or U21762 (N_21762,N_15382,N_18054);
or U21763 (N_21763,N_16281,N_19125);
nor U21764 (N_21764,N_16711,N_15756);
and U21765 (N_21765,N_15199,N_15394);
xnor U21766 (N_21766,N_15535,N_19975);
nor U21767 (N_21767,N_18454,N_17584);
nor U21768 (N_21768,N_17297,N_19241);
nor U21769 (N_21769,N_15768,N_18640);
or U21770 (N_21770,N_15130,N_19751);
or U21771 (N_21771,N_19374,N_16425);
nand U21772 (N_21772,N_17968,N_19792);
nand U21773 (N_21773,N_18994,N_18553);
or U21774 (N_21774,N_15467,N_19742);
xor U21775 (N_21775,N_15142,N_17118);
nor U21776 (N_21776,N_18003,N_15127);
nor U21777 (N_21777,N_19234,N_19763);
nand U21778 (N_21778,N_17489,N_15748);
or U21779 (N_21779,N_15191,N_15937);
nand U21780 (N_21780,N_15674,N_19023);
or U21781 (N_21781,N_19817,N_19683);
nand U21782 (N_21782,N_15266,N_18380);
or U21783 (N_21783,N_19221,N_17655);
and U21784 (N_21784,N_15202,N_17939);
nand U21785 (N_21785,N_15699,N_17062);
and U21786 (N_21786,N_17238,N_19252);
nor U21787 (N_21787,N_15476,N_18280);
or U21788 (N_21788,N_16195,N_17787);
or U21789 (N_21789,N_19436,N_16718);
xor U21790 (N_21790,N_16799,N_17318);
and U21791 (N_21791,N_15258,N_16046);
nor U21792 (N_21792,N_15744,N_18282);
and U21793 (N_21793,N_18605,N_19977);
nor U21794 (N_21794,N_15751,N_15245);
or U21795 (N_21795,N_15097,N_19821);
nand U21796 (N_21796,N_16691,N_16774);
or U21797 (N_21797,N_19510,N_18885);
and U21798 (N_21798,N_19659,N_18849);
and U21799 (N_21799,N_19524,N_15587);
or U21800 (N_21800,N_15743,N_17485);
nor U21801 (N_21801,N_17346,N_18807);
or U21802 (N_21802,N_17618,N_19930);
and U21803 (N_21803,N_17806,N_17940);
and U21804 (N_21804,N_17748,N_17171);
and U21805 (N_21805,N_17810,N_19604);
and U21806 (N_21806,N_19274,N_19493);
nand U21807 (N_21807,N_16784,N_17391);
nand U21808 (N_21808,N_17553,N_15454);
or U21809 (N_21809,N_17303,N_15168);
nor U21810 (N_21810,N_15379,N_18905);
nor U21811 (N_21811,N_15641,N_15949);
or U21812 (N_21812,N_19691,N_18163);
xnor U21813 (N_21813,N_18554,N_15935);
and U21814 (N_21814,N_17001,N_15420);
or U21815 (N_21815,N_16555,N_19569);
and U21816 (N_21816,N_17165,N_18450);
and U21817 (N_21817,N_17958,N_16549);
nor U21818 (N_21818,N_19624,N_19744);
nand U21819 (N_21819,N_17319,N_15500);
or U21820 (N_21820,N_19996,N_15609);
nor U21821 (N_21821,N_15424,N_15792);
nor U21822 (N_21822,N_15774,N_16462);
and U21823 (N_21823,N_18075,N_18611);
or U21824 (N_21824,N_16014,N_18217);
and U21825 (N_21825,N_15562,N_19828);
nor U21826 (N_21826,N_16189,N_19056);
nand U21827 (N_21827,N_16755,N_19514);
and U21828 (N_21828,N_17605,N_18903);
nor U21829 (N_21829,N_16165,N_17481);
nor U21830 (N_21830,N_16535,N_18250);
nor U21831 (N_21831,N_15066,N_19272);
nand U21832 (N_21832,N_15955,N_18606);
and U21833 (N_21833,N_18231,N_17540);
and U21834 (N_21834,N_16488,N_15295);
or U21835 (N_21835,N_18623,N_15241);
nor U21836 (N_21836,N_17951,N_16832);
and U21837 (N_21837,N_18130,N_16388);
or U21838 (N_21838,N_19346,N_16075);
and U21839 (N_21839,N_16901,N_15509);
or U21840 (N_21840,N_19370,N_18514);
or U21841 (N_21841,N_16738,N_15624);
nor U21842 (N_21842,N_16257,N_18168);
nor U21843 (N_21843,N_18599,N_16394);
and U21844 (N_21844,N_19040,N_19663);
nand U21845 (N_21845,N_19945,N_15369);
nand U21846 (N_21846,N_17541,N_16698);
or U21847 (N_21847,N_16717,N_16125);
or U21848 (N_21848,N_15313,N_17091);
nand U21849 (N_21849,N_15435,N_19981);
and U21850 (N_21850,N_19162,N_15892);
or U21851 (N_21851,N_19507,N_15378);
or U21852 (N_21852,N_19068,N_16735);
nor U21853 (N_21853,N_18080,N_15040);
and U21854 (N_21854,N_17006,N_17267);
or U21855 (N_21855,N_19826,N_16536);
or U21856 (N_21856,N_16248,N_16496);
nand U21857 (N_21857,N_18821,N_18480);
nor U21858 (N_21858,N_18880,N_16721);
and U21859 (N_21859,N_16106,N_15026);
nand U21860 (N_21860,N_19760,N_16168);
xor U21861 (N_21861,N_17072,N_16756);
nand U21862 (N_21862,N_19628,N_15484);
nor U21863 (N_21863,N_15048,N_18987);
or U21864 (N_21864,N_19911,N_15465);
and U21865 (N_21865,N_16256,N_16572);
and U21866 (N_21866,N_15143,N_18149);
nand U21867 (N_21867,N_17345,N_17112);
and U21868 (N_21868,N_16198,N_19517);
nor U21869 (N_21869,N_19956,N_18956);
nand U21870 (N_21870,N_15336,N_16941);
and U21871 (N_21871,N_17395,N_19842);
nand U21872 (N_21872,N_16562,N_18798);
and U21873 (N_21873,N_19905,N_17337);
or U21874 (N_21874,N_15755,N_15125);
or U21875 (N_21875,N_19861,N_15613);
nor U21876 (N_21876,N_17649,N_16395);
nor U21877 (N_21877,N_15637,N_19574);
and U21878 (N_21878,N_18192,N_19425);
nand U21879 (N_21879,N_19189,N_18859);
or U21880 (N_21880,N_16200,N_17984);
and U21881 (N_21881,N_18330,N_15128);
nor U21882 (N_21882,N_15046,N_17483);
nand U21883 (N_21883,N_17784,N_16620);
or U21884 (N_21884,N_15884,N_19718);
or U21885 (N_21885,N_16077,N_19074);
nand U21886 (N_21886,N_16912,N_15520);
or U21887 (N_21887,N_19192,N_17090);
nor U21888 (N_21888,N_19172,N_19087);
and U21889 (N_21889,N_17246,N_16017);
nand U21890 (N_21890,N_19430,N_16042);
or U21891 (N_21891,N_18323,N_17586);
nor U21892 (N_21892,N_19553,N_16769);
nand U21893 (N_21893,N_19504,N_16484);
nor U21894 (N_21894,N_18435,N_19704);
nand U21895 (N_21895,N_18750,N_15203);
or U21896 (N_21896,N_15437,N_16270);
nand U21897 (N_21897,N_16942,N_16253);
or U21898 (N_21898,N_18503,N_15835);
or U21899 (N_21899,N_18258,N_18993);
nand U21900 (N_21900,N_19822,N_15534);
and U21901 (N_21901,N_19789,N_17668);
and U21902 (N_21902,N_19657,N_17757);
nor U21903 (N_21903,N_16652,N_17054);
nor U21904 (N_21904,N_15962,N_18730);
and U21905 (N_21905,N_15186,N_17250);
nor U21906 (N_21906,N_17327,N_19206);
nor U21907 (N_21907,N_15035,N_19688);
nand U21908 (N_21908,N_19010,N_16834);
and U21909 (N_21909,N_16199,N_17927);
nor U21910 (N_21910,N_19679,N_18710);
or U21911 (N_21911,N_17591,N_18151);
nand U21912 (N_21912,N_15556,N_16624);
nand U21913 (N_21913,N_18415,N_19976);
or U21914 (N_21914,N_16230,N_16440);
nand U21915 (N_21915,N_17636,N_17080);
or U21916 (N_21916,N_18904,N_15841);
nor U21917 (N_21917,N_17304,N_16185);
and U21918 (N_21918,N_16324,N_17375);
and U21919 (N_21919,N_17950,N_19096);
or U21920 (N_21920,N_17219,N_15167);
or U21921 (N_21921,N_18053,N_18607);
nor U21922 (N_21922,N_15643,N_15366);
and U21923 (N_21923,N_18591,N_19297);
nor U21924 (N_21924,N_16848,N_19465);
nor U21925 (N_21925,N_17315,N_15547);
or U21926 (N_21926,N_18959,N_15605);
nor U21927 (N_21927,N_19397,N_16381);
xnor U21928 (N_21928,N_15021,N_17107);
and U21929 (N_21929,N_15423,N_19805);
and U21930 (N_21930,N_17731,N_17000);
and U21931 (N_21931,N_15996,N_18208);
xor U21932 (N_21932,N_19639,N_15176);
and U21933 (N_21933,N_19318,N_19962);
and U21934 (N_21934,N_16819,N_17607);
nor U21935 (N_21935,N_19530,N_19841);
nor U21936 (N_21936,N_17923,N_16119);
or U21937 (N_21937,N_18620,N_17703);
nor U21938 (N_21938,N_18129,N_18451);
and U21939 (N_21939,N_15456,N_17310);
and U21940 (N_21940,N_15218,N_16096);
nor U21941 (N_21941,N_19883,N_19940);
nand U21942 (N_21942,N_19114,N_15069);
nand U21943 (N_21943,N_18252,N_18628);
nor U21944 (N_21944,N_16530,N_18114);
nand U21945 (N_21945,N_18576,N_15762);
nand U21946 (N_21946,N_17659,N_18556);
or U21947 (N_21947,N_16354,N_16280);
and U21948 (N_21948,N_16655,N_19138);
or U21949 (N_21949,N_16150,N_19383);
and U21950 (N_21950,N_15948,N_17773);
nor U21951 (N_21951,N_15123,N_18542);
nand U21952 (N_21952,N_16112,N_16955);
nor U21953 (N_21953,N_17127,N_18050);
and U21954 (N_21954,N_19754,N_19455);
and U21955 (N_21955,N_16547,N_16994);
nor U21956 (N_21956,N_18385,N_15401);
nor U21957 (N_21957,N_17321,N_18861);
or U21958 (N_21958,N_18409,N_17019);
and U21959 (N_21959,N_15045,N_17778);
nor U21960 (N_21960,N_16362,N_16719);
and U21961 (N_21961,N_16508,N_18537);
nor U21962 (N_21962,N_16812,N_18035);
or U21963 (N_21963,N_15335,N_15978);
nor U21964 (N_21964,N_18876,N_16914);
and U21965 (N_21965,N_16476,N_19236);
and U21966 (N_21966,N_16906,N_16160);
nand U21967 (N_21967,N_16643,N_17802);
nand U21968 (N_21968,N_18873,N_19984);
and U21969 (N_21969,N_15612,N_15553);
and U21970 (N_21970,N_15226,N_16954);
and U21971 (N_21971,N_17755,N_19773);
nand U21972 (N_21972,N_16379,N_18479);
and U21973 (N_21973,N_15063,N_17079);
or U21974 (N_21974,N_18944,N_18777);
xor U21975 (N_21975,N_19611,N_16071);
nor U21976 (N_21976,N_15268,N_19857);
or U21977 (N_21977,N_19597,N_17434);
or U21978 (N_21978,N_17785,N_15677);
nor U21979 (N_21979,N_15274,N_19175);
xnor U21980 (N_21980,N_15850,N_15865);
and U21981 (N_21981,N_15620,N_17456);
nor U21982 (N_21982,N_17518,N_17386);
and U21983 (N_21983,N_15571,N_19739);
nand U21984 (N_21984,N_19932,N_19811);
and U21985 (N_21985,N_15110,N_18301);
and U21986 (N_21986,N_18643,N_15974);
and U21987 (N_21987,N_19230,N_18136);
nor U21988 (N_21988,N_16634,N_15252);
and U21989 (N_21989,N_15880,N_18095);
nor U21990 (N_21990,N_17845,N_15831);
nor U21991 (N_21991,N_18447,N_18828);
nor U21992 (N_21992,N_15414,N_16043);
nand U21993 (N_21993,N_19435,N_15495);
nand U21994 (N_21994,N_15460,N_19489);
or U21995 (N_21995,N_19485,N_15140);
nand U21996 (N_21996,N_15993,N_17758);
and U21997 (N_21997,N_16443,N_16258);
nor U21998 (N_21998,N_17411,N_15808);
nor U21999 (N_21999,N_15820,N_16499);
or U22000 (N_22000,N_19244,N_18277);
and U22001 (N_22001,N_17909,N_16701);
or U22002 (N_22002,N_16627,N_18009);
and U22003 (N_22003,N_19564,N_17447);
and U22004 (N_22004,N_16745,N_18865);
and U22005 (N_22005,N_16605,N_17452);
and U22006 (N_22006,N_19675,N_18683);
nor U22007 (N_22007,N_17545,N_19123);
nor U22008 (N_22008,N_17809,N_19498);
nand U22009 (N_22009,N_19352,N_16123);
nor U22010 (N_22010,N_17068,N_17131);
or U22011 (N_22011,N_17437,N_18421);
and U22012 (N_22012,N_17273,N_19311);
and U22013 (N_22013,N_15240,N_15698);
nor U22014 (N_22014,N_19658,N_17592);
and U22015 (N_22015,N_15923,N_17684);
nor U22016 (N_22016,N_15428,N_16426);
or U22017 (N_22017,N_18914,N_18310);
or U22018 (N_22018,N_17049,N_16993);
nor U22019 (N_22019,N_19121,N_17715);
and U22020 (N_22020,N_18344,N_16807);
or U22021 (N_22021,N_17120,N_16509);
nor U22022 (N_22022,N_15407,N_18631);
or U22023 (N_22023,N_15788,N_19128);
and U22024 (N_22024,N_19761,N_15384);
or U22025 (N_22025,N_18900,N_16245);
nor U22026 (N_22026,N_15869,N_16128);
nand U22027 (N_22027,N_19135,N_17506);
nor U22028 (N_22028,N_19163,N_19966);
nand U22029 (N_22029,N_17975,N_15981);
or U22030 (N_22030,N_18600,N_18921);
or U22031 (N_22031,N_16184,N_16723);
nor U22032 (N_22032,N_16667,N_17885);
and U22033 (N_22033,N_16714,N_16873);
nor U22034 (N_22034,N_17895,N_16278);
and U22035 (N_22035,N_18092,N_19661);
nor U22036 (N_22036,N_16350,N_17848);
and U22037 (N_22037,N_15881,N_18413);
and U22038 (N_22038,N_19617,N_17245);
or U22039 (N_22039,N_15120,N_19891);
or U22040 (N_22040,N_17419,N_18356);
nand U22041 (N_22041,N_19999,N_19563);
or U22042 (N_22042,N_16216,N_19451);
and U22043 (N_22043,N_16932,N_17232);
nand U22044 (N_22044,N_16759,N_18267);
nor U22045 (N_22045,N_16904,N_18419);
and U22046 (N_22046,N_16913,N_18842);
nand U22047 (N_22047,N_15963,N_18562);
and U22048 (N_22048,N_15297,N_15482);
and U22049 (N_22049,N_16034,N_16824);
nand U22050 (N_22050,N_16829,N_19948);
and U22051 (N_22051,N_17030,N_19226);
nor U22052 (N_22052,N_16531,N_17380);
and U22053 (N_22053,N_18566,N_15950);
xor U22054 (N_22054,N_18405,N_17723);
and U22055 (N_22055,N_15310,N_18428);
nor U22056 (N_22056,N_19527,N_17702);
nand U22057 (N_22057,N_19888,N_19788);
or U22058 (N_22058,N_17140,N_17093);
and U22059 (N_22059,N_19551,N_15158);
or U22060 (N_22060,N_17401,N_16460);
nor U22061 (N_22061,N_15968,N_16261);
or U22062 (N_22062,N_19405,N_19009);
nor U22063 (N_22063,N_17114,N_18595);
nor U22064 (N_22064,N_16387,N_15752);
nand U22065 (N_22065,N_19541,N_19660);
or U22066 (N_22066,N_19595,N_19955);
nor U22067 (N_22067,N_19371,N_15065);
nand U22068 (N_22068,N_16308,N_15062);
nor U22069 (N_22069,N_19026,N_16453);
or U22070 (N_22070,N_15308,N_18004);
nor U22071 (N_22071,N_16157,N_16048);
and U22072 (N_22072,N_19528,N_16911);
nand U22073 (N_22073,N_16039,N_19414);
nand U22074 (N_22074,N_17320,N_16727);
nand U22075 (N_22075,N_16178,N_16981);
nand U22076 (N_22076,N_17056,N_17976);
nor U22077 (N_22077,N_15425,N_18240);
xor U22078 (N_22078,N_19715,N_16669);
nor U22079 (N_22079,N_18452,N_18088);
nor U22080 (N_22080,N_16545,N_15436);
and U22081 (N_22081,N_19759,N_17526);
nand U22082 (N_22082,N_17343,N_18614);
nor U22083 (N_22083,N_16501,N_18813);
and U22084 (N_22084,N_15405,N_19605);
nor U22085 (N_22085,N_18910,N_17973);
or U22086 (N_22086,N_18496,N_18390);
nand U22087 (N_22087,N_16975,N_18901);
or U22088 (N_22088,N_16628,N_15780);
nor U22089 (N_22089,N_15085,N_18713);
and U22090 (N_22090,N_17918,N_18425);
xor U22091 (N_22091,N_19668,N_15488);
and U22092 (N_22092,N_19364,N_15805);
nor U22093 (N_22093,N_15318,N_17970);
and U22094 (N_22094,N_19136,N_15246);
nand U22095 (N_22095,N_17645,N_16825);
or U22096 (N_22096,N_17094,N_16561);
nand U22097 (N_22097,N_17782,N_16816);
nor U22098 (N_22098,N_17192,N_16595);
and U22099 (N_22099,N_18188,N_18687);
and U22100 (N_22100,N_18275,N_18461);
and U22101 (N_22101,N_17096,N_19916);
nor U22102 (N_22102,N_18775,N_18772);
nor U22103 (N_22103,N_19249,N_17124);
and U22104 (N_22104,N_18167,N_15411);
or U22105 (N_22105,N_18245,N_15852);
and U22106 (N_22106,N_17089,N_15184);
nor U22107 (N_22107,N_15215,N_19363);
xnor U22108 (N_22108,N_16352,N_19004);
nor U22109 (N_22109,N_17953,N_15220);
nor U22110 (N_22110,N_17243,N_17678);
and U22111 (N_22111,N_19566,N_15075);
nor U22112 (N_22112,N_15786,N_19310);
nand U22113 (N_22113,N_19859,N_16016);
and U22114 (N_22114,N_15854,N_16768);
nor U22115 (N_22115,N_15924,N_17335);
nand U22116 (N_22116,N_16660,N_18005);
and U22117 (N_22117,N_19833,N_17193);
and U22118 (N_22118,N_19078,N_15471);
nor U22119 (N_22119,N_15975,N_18671);
and U22120 (N_22120,N_18868,N_17949);
or U22121 (N_22121,N_16692,N_18594);
nor U22122 (N_22122,N_17991,N_18799);
nand U22123 (N_22123,N_17087,N_19719);
or U22124 (N_22124,N_18579,N_15230);
or U22125 (N_22125,N_15141,N_19377);
and U22126 (N_22126,N_15802,N_15630);
and U22127 (N_22127,N_19250,N_15681);
nor U22128 (N_22128,N_18706,N_19636);
nand U22129 (N_22129,N_15998,N_17817);
nor U22130 (N_22130,N_15807,N_15177);
nor U22131 (N_22131,N_15763,N_17843);
or U22132 (N_22132,N_16788,N_17839);
nor U22133 (N_22133,N_19620,N_18497);
and U22134 (N_22134,N_19233,N_18870);
nor U22135 (N_22135,N_18883,N_18662);
or U22136 (N_22136,N_18577,N_17314);
nor U22137 (N_22137,N_17615,N_18298);
nand U22138 (N_22138,N_17767,N_17230);
nor U22139 (N_22139,N_15885,N_16335);
or U22140 (N_22140,N_16382,N_15438);
or U22141 (N_22141,N_18044,N_19287);
or U22142 (N_22142,N_16617,N_19427);
nor U22143 (N_22143,N_19757,N_16984);
and U22144 (N_22144,N_16217,N_16477);
nand U22145 (N_22145,N_19296,N_18135);
or U22146 (N_22146,N_16188,N_18002);
nor U22147 (N_22147,N_16680,N_15803);
nand U22148 (N_22148,N_19589,N_15244);
or U22149 (N_22149,N_17977,N_19978);
nand U22150 (N_22150,N_15857,N_17197);
nand U22151 (N_22151,N_15380,N_19699);
nor U22152 (N_22152,N_19292,N_16675);
xor U22153 (N_22153,N_17764,N_15403);
or U22154 (N_22154,N_19277,N_16344);
nor U22155 (N_22155,N_17292,N_19892);
and U22156 (N_22156,N_18247,N_15102);
nand U22157 (N_22157,N_16538,N_15294);
or U22158 (N_22158,N_15703,N_17344);
or U22159 (N_22159,N_16191,N_18862);
and U22160 (N_22160,N_15198,N_16340);
and U22161 (N_22161,N_18781,N_16159);
nand U22162 (N_22162,N_17205,N_18657);
or U22163 (N_22163,N_16677,N_19626);
nor U22164 (N_22164,N_16557,N_17906);
and U22165 (N_22165,N_18081,N_19533);
and U22166 (N_22166,N_17917,N_17533);
nor U22167 (N_22167,N_16418,N_18012);
or U22168 (N_22168,N_19705,N_17323);
nand U22169 (N_22169,N_15608,N_18457);
and U22170 (N_22170,N_19062,N_18552);
and U22171 (N_22171,N_17023,N_17233);
nor U22172 (N_22172,N_17356,N_17751);
nand U22173 (N_22173,N_17313,N_17856);
and U22174 (N_22174,N_16290,N_19568);
or U22175 (N_22175,N_17603,N_17189);
and U22176 (N_22176,N_18416,N_16260);
nand U22177 (N_22177,N_16618,N_15591);
or U22178 (N_22178,N_19055,N_18022);
or U22179 (N_22179,N_18733,N_15247);
nand U22180 (N_22180,N_19621,N_17229);
and U22181 (N_22181,N_19454,N_18763);
and U22182 (N_22182,N_16328,N_16971);
and U22183 (N_22183,N_19264,N_15204);
nor U22184 (N_22184,N_16321,N_19011);
and U22185 (N_22185,N_15479,N_19549);
and U22186 (N_22186,N_15710,N_17967);
nor U22187 (N_22187,N_17947,N_16242);
nand U22188 (N_22188,N_15466,N_19079);
and U22189 (N_22189,N_15361,N_17099);
nor U22190 (N_22190,N_15345,N_19431);
nor U22191 (N_22191,N_15555,N_19804);
or U22192 (N_22192,N_18509,N_17252);
xnor U22193 (N_22193,N_17222,N_19351);
and U22194 (N_22194,N_15032,N_16888);
xnor U22195 (N_22195,N_17284,N_16821);
or U22196 (N_22196,N_15938,N_19475);
xor U22197 (N_22197,N_17472,N_18077);
nand U22198 (N_22198,N_18418,N_19407);
nand U22199 (N_22199,N_18427,N_18148);
and U22200 (N_22200,N_16553,N_15253);
nor U22201 (N_22201,N_18978,N_16301);
nand U22202 (N_22202,N_19738,N_18791);
xnor U22203 (N_22203,N_19713,N_18111);
nor U22204 (N_22204,N_19103,N_18787);
or U22205 (N_22205,N_18391,N_19357);
and U22206 (N_22206,N_18049,N_16938);
and U22207 (N_22207,N_18322,N_15137);
nor U22208 (N_22208,N_16897,N_18371);
nor U22209 (N_22209,N_19083,N_17389);
nor U22210 (N_22210,N_18063,N_16003);
or U22211 (N_22211,N_15705,N_16105);
nor U22212 (N_22212,N_16404,N_18735);
nor U22213 (N_22213,N_17997,N_15473);
nor U22214 (N_22214,N_15662,N_16700);
or U22215 (N_22215,N_18727,N_17159);
and U22216 (N_22216,N_19054,N_16289);
nand U22217 (N_22217,N_18672,N_17609);
and U22218 (N_22218,N_15205,N_18886);
or U22219 (N_22219,N_15413,N_17744);
nor U22220 (N_22220,N_15510,N_15162);
or U22221 (N_22221,N_17224,N_19106);
nand U22222 (N_22222,N_16930,N_16487);
and U22223 (N_22223,N_17728,N_17714);
nand U22224 (N_22224,N_15459,N_16783);
and U22225 (N_22225,N_15838,N_19315);
and U22226 (N_22226,N_15577,N_15217);
nor U22227 (N_22227,N_16683,N_17151);
nand U22228 (N_22228,N_18198,N_17003);
nand U22229 (N_22229,N_18387,N_18260);
nand U22230 (N_22230,N_18061,N_18839);
nor U22231 (N_22231,N_17628,N_16304);
nand U22232 (N_22232,N_18635,N_19028);
nor U22233 (N_22233,N_19576,N_18609);
nor U22234 (N_22234,N_18006,N_15586);
or U22235 (N_22235,N_16550,N_19355);
or U22236 (N_22236,N_19193,N_19324);
nor U22237 (N_22237,N_19181,N_19421);
nand U22238 (N_22238,N_17147,N_16556);
or U22239 (N_22239,N_19030,N_17935);
or U22240 (N_22240,N_18572,N_15337);
nor U22241 (N_22241,N_16521,N_19006);
and U22242 (N_22242,N_17852,N_17223);
and U22243 (N_22243,N_17573,N_19327);
nor U22244 (N_22244,N_17639,N_18958);
and U22245 (N_22245,N_17629,N_18714);
nor U22246 (N_22246,N_15328,N_16353);
and U22247 (N_22247,N_17085,N_16720);
nand U22248 (N_22248,N_19581,N_16782);
nor U22249 (N_22249,N_15784,N_16640);
nand U22250 (N_22250,N_15033,N_15223);
or U22251 (N_22251,N_15163,N_16582);
nor U22252 (N_22252,N_15584,N_17993);
nor U22253 (N_22253,N_15530,N_15242);
nand U22254 (N_22254,N_18530,N_15976);
nor U22255 (N_22255,N_17402,N_19273);
or U22256 (N_22256,N_17742,N_16424);
and U22257 (N_22257,N_19554,N_15306);
nand U22258 (N_22258,N_17805,N_18856);
or U22259 (N_22259,N_16138,N_18162);
and U22260 (N_22260,N_19251,N_17150);
nor U22261 (N_22261,N_17595,N_15965);
and U22262 (N_22262,N_18947,N_19293);
or U22263 (N_22263,N_16001,N_19982);
or U22264 (N_22264,N_19059,N_18381);
nor U22265 (N_22265,N_19750,N_18642);
and U22266 (N_22266,N_17185,N_19690);
or U22267 (N_22267,N_15194,N_16022);
and U22268 (N_22268,N_15543,N_17849);
nand U22269 (N_22269,N_16874,N_16573);
and U22270 (N_22270,N_17931,N_15837);
nand U22271 (N_22271,N_16748,N_15845);
nand U22272 (N_22272,N_18884,N_19196);
nand U22273 (N_22273,N_15044,N_17963);
and U22274 (N_22274,N_18512,N_18918);
nand U22275 (N_22275,N_17163,N_18182);
nor U22276 (N_22276,N_19035,N_18057);
and U22277 (N_22277,N_18696,N_19567);
and U22278 (N_22278,N_18663,N_17363);
nand U22279 (N_22279,N_16798,N_19623);
and U22280 (N_22280,N_17900,N_19039);
or U22281 (N_22281,N_15497,N_18811);
nor U22282 (N_22282,N_18354,N_16209);
nand U22283 (N_22283,N_18827,N_16566);
nand U22284 (N_22284,N_19559,N_16978);
nand U22285 (N_22285,N_19429,N_16078);
nor U22286 (N_22286,N_19853,N_17078);
and U22287 (N_22287,N_19730,N_19871);
or U22288 (N_22288,N_15664,N_15511);
and U22289 (N_22289,N_16236,N_17567);
or U22290 (N_22290,N_16953,N_19116);
or U22291 (N_22291,N_19199,N_19375);
or U22292 (N_22292,N_16761,N_18318);
and U22293 (N_22293,N_17505,N_17477);
nand U22294 (N_22294,N_17496,N_15322);
nand U22295 (N_22295,N_16747,N_17528);
nor U22296 (N_22296,N_16082,N_18830);
nor U22297 (N_22297,N_18965,N_17298);
and U22298 (N_22298,N_15316,N_19518);
or U22299 (N_22299,N_16428,N_17404);
and U22300 (N_22300,N_18412,N_16923);
and U22301 (N_22301,N_16177,N_15671);
or U22302 (N_22302,N_18540,N_15339);
nor U22303 (N_22303,N_15400,N_15815);
nor U22304 (N_22304,N_19245,N_16373);
nand U22305 (N_22305,N_18379,N_16567);
or U22306 (N_22306,N_17544,N_15171);
nor U22307 (N_22307,N_15874,N_15330);
nor U22308 (N_22308,N_16307,N_16406);
nor U22309 (N_22309,N_15017,N_16283);
nor U22310 (N_22310,N_19432,N_17161);
nor U22311 (N_22311,N_18305,N_18920);
nand U22312 (N_22312,N_15022,N_16900);
or U22313 (N_22313,N_19505,N_17479);
or U22314 (N_22314,N_18183,N_16166);
nor U22315 (N_22315,N_17648,N_19785);
nand U22316 (N_22316,N_15058,N_15169);
or U22317 (N_22317,N_17530,N_15325);
and U22318 (N_22318,N_16520,N_17729);
nand U22319 (N_22319,N_17195,N_15941);
nand U22320 (N_22320,N_16080,N_15825);
nor U22321 (N_22321,N_15326,N_19830);
or U22322 (N_22322,N_16452,N_17241);
and U22323 (N_22323,N_17697,N_18780);
nand U22324 (N_22324,N_17912,N_15908);
nand U22325 (N_22325,N_15430,N_15051);
or U22326 (N_22326,N_15333,N_19912);
nand U22327 (N_22327,N_17162,N_15640);
nand U22328 (N_22328,N_16920,N_17046);
or U22329 (N_22329,N_18494,N_16451);
or U22330 (N_22330,N_18673,N_19947);
nand U22331 (N_22331,N_17033,N_19144);
and U22332 (N_22332,N_19129,N_16823);
nand U22333 (N_22333,N_16715,N_19852);
or U22334 (N_22334,N_15422,N_17325);
nand U22335 (N_22335,N_16480,N_17966);
or U22336 (N_22336,N_18753,N_15279);
and U22337 (N_22337,N_17034,N_15301);
and U22338 (N_22338,N_15843,N_16397);
and U22339 (N_22339,N_18173,N_17777);
nor U22340 (N_22340,N_19542,N_19521);
or U22341 (N_22341,N_18887,N_19345);
and U22342 (N_22342,N_17867,N_15371);
or U22343 (N_22343,N_18871,N_16056);
or U22344 (N_22344,N_16789,N_19716);
nand U22345 (N_22345,N_19159,N_15512);
and U22346 (N_22346,N_18402,N_19354);
or U22347 (N_22347,N_16268,N_16685);
nor U22348 (N_22348,N_19229,N_18928);
or U22349 (N_22349,N_17719,N_16464);
and U22350 (N_22350,N_16370,N_16512);
and U22351 (N_22351,N_17332,N_18858);
or U22352 (N_22352,N_18466,N_18505);
nor U22353 (N_22353,N_19307,N_15480);
nor U22354 (N_22354,N_16413,N_18034);
or U22355 (N_22355,N_18046,N_15426);
or U22356 (N_22356,N_17379,N_16009);
and U22357 (N_22357,N_19874,N_16766);
or U22358 (N_22358,N_16696,N_18774);
and U22359 (N_22359,N_17493,N_16924);
and U22360 (N_22360,N_17669,N_17833);
and U22361 (N_22361,N_17186,N_16686);
nand U22362 (N_22362,N_15351,N_15172);
xor U22363 (N_22363,N_17207,N_19692);
or U22364 (N_22364,N_19733,N_18118);
and U22365 (N_22365,N_18707,N_18445);
nand U22366 (N_22366,N_15693,N_19584);
nand U22367 (N_22367,N_17109,N_19178);
and U22368 (N_22368,N_19093,N_17593);
nand U22369 (N_22369,N_17500,N_19072);
nand U22370 (N_22370,N_16497,N_18695);
nor U22371 (N_22371,N_18365,N_18789);
nand U22372 (N_22372,N_19480,N_18386);
nand U22373 (N_22373,N_15992,N_19142);
or U22374 (N_22374,N_16365,N_17148);
or U22375 (N_22375,N_15104,N_15789);
nor U22376 (N_22376,N_15076,N_19210);
and U22377 (N_22377,N_19434,N_16544);
nand U22378 (N_22378,N_16232,N_15264);
or U22379 (N_22379,N_19513,N_16612);
and U22380 (N_22380,N_18597,N_18894);
nor U22381 (N_22381,N_18481,N_17765);
or U22382 (N_22382,N_17695,N_18336);
and U22383 (N_22383,N_19807,N_18307);
or U22384 (N_22384,N_18158,N_15812);
nor U22385 (N_22385,N_16517,N_15660);
nand U22386 (N_22386,N_17641,N_18761);
and U22387 (N_22387,N_16817,N_18468);
and U22388 (N_22388,N_17887,N_15779);
nor U22389 (N_22389,N_18471,N_16478);
and U22390 (N_22390,N_15052,N_18527);
and U22391 (N_22391,N_15508,N_17656);
and U22392 (N_22392,N_16131,N_16347);
or U22393 (N_22393,N_18536,N_17468);
or U22394 (N_22394,N_17365,N_19167);
nand U22395 (N_22395,N_17340,N_16359);
nand U22396 (N_22396,N_17132,N_16051);
and U22397 (N_22397,N_17347,N_17995);
or U22398 (N_22398,N_15312,N_17381);
or U22399 (N_22399,N_16991,N_19066);
nor U22400 (N_22400,N_18508,N_19372);
nand U22401 (N_22401,N_19102,N_15600);
or U22402 (N_22402,N_15300,N_15149);
and U22403 (N_22403,N_16601,N_19820);
nor U22404 (N_22404,N_19900,N_16831);
nand U22405 (N_22405,N_18052,N_18306);
nand U22406 (N_22406,N_16600,N_16986);
nand U22407 (N_22407,N_16899,N_18636);
and U22408 (N_22408,N_18806,N_17552);
or U22409 (N_22409,N_17488,N_19964);
nor U22410 (N_22410,N_18932,N_15059);
or U22411 (N_22411,N_18205,N_16576);
xor U22412 (N_22412,N_16621,N_16325);
and U22413 (N_22413,N_18983,N_17143);
nand U22414 (N_22414,N_16076,N_15777);
and U22415 (N_22415,N_15472,N_16389);
or U22416 (N_22416,N_18751,N_15675);
or U22417 (N_22417,N_19583,N_18765);
or U22418 (N_22418,N_19064,N_19543);
nand U22419 (N_22419,N_19065,N_15648);
or U22420 (N_22420,N_16318,N_16827);
nor U22421 (N_22421,N_16629,N_15113);
nor U22422 (N_22422,N_17302,N_17512);
nor U22423 (N_22423,N_19753,N_15487);
or U22424 (N_22424,N_15028,N_19161);
nand U22425 (N_22425,N_17811,N_16061);
nor U22426 (N_22426,N_16988,N_15713);
or U22427 (N_22427,N_16884,N_18872);
nor U22428 (N_22428,N_18940,N_16327);
and U22429 (N_22429,N_16441,N_18472);
nor U22430 (N_22430,N_19111,N_15095);
or U22431 (N_22431,N_15352,N_16809);
and U22432 (N_22432,N_18783,N_15183);
nand U22433 (N_22433,N_17475,N_16423);
or U22434 (N_22434,N_19156,N_18911);
nor U22435 (N_22435,N_17911,N_19268);
nand U22436 (N_22436,N_19067,N_16064);
nor U22437 (N_22437,N_18991,N_18999);
and U22438 (N_22438,N_18268,N_15262);
nor U22439 (N_22439,N_16296,N_18935);
nor U22440 (N_22440,N_18711,N_19494);
nand U22441 (N_22441,N_19213,N_19320);
nand U22442 (N_22442,N_15704,N_18697);
nor U22443 (N_22443,N_16949,N_18016);
nor U22444 (N_22444,N_18329,N_17442);
nand U22445 (N_22445,N_19849,N_17117);
and U22446 (N_22446,N_15532,N_18203);
nand U22447 (N_22447,N_15375,N_19248);
nand U22448 (N_22448,N_19655,N_16429);
or U22449 (N_22449,N_18637,N_17055);
nand U22450 (N_22450,N_18854,N_16903);
and U22451 (N_22451,N_17338,N_17466);
and U22452 (N_22452,N_15334,N_15499);
nor U22453 (N_22453,N_19466,N_18404);
nor U22454 (N_22454,N_17665,N_19238);
or U22455 (N_22455,N_18423,N_19587);
or U22456 (N_22456,N_17368,N_19218);
nand U22457 (N_22457,N_17683,N_18604);
nand U22458 (N_22458,N_15291,N_19409);
nor U22459 (N_22459,N_15402,N_15404);
nand U22460 (N_22460,N_18093,N_16254);
and U22461 (N_22461,N_18875,N_16758);
and U22462 (N_22462,N_15873,N_16028);
nor U22463 (N_22463,N_16699,N_18945);
nor U22464 (N_22464,N_19112,N_17720);
nor U22465 (N_22465,N_19032,N_17121);
and U22466 (N_22466,N_15957,N_16744);
or U22467 (N_22467,N_18187,N_15200);
nor U22468 (N_22468,N_18303,N_16263);
nor U22469 (N_22469,N_17672,N_19484);
nor U22470 (N_22470,N_15991,N_15082);
or U22471 (N_22471,N_19522,N_19304);
nor U22472 (N_22472,N_18436,N_18083);
xnor U22473 (N_22473,N_15216,N_18869);
and U22474 (N_22474,N_15249,N_19774);
nand U22475 (N_22475,N_16729,N_18860);
or U22476 (N_22476,N_17746,N_16433);
nor U22477 (N_22477,N_16486,N_18729);
or U22478 (N_22478,N_16935,N_18715);
nand U22479 (N_22479,N_17416,N_16786);
nand U22480 (N_22480,N_19778,N_16393);
nor U22481 (N_22481,N_19935,N_17508);
nor U22482 (N_22482,N_19342,N_17457);
nor U22483 (N_22483,N_16838,N_16065);
nor U22484 (N_22484,N_15910,N_17964);
and U22485 (N_22485,N_18334,N_17934);
and U22486 (N_22486,N_15888,N_18782);
or U22487 (N_22487,N_18357,N_16856);
and U22488 (N_22488,N_15207,N_19294);
nand U22489 (N_22489,N_17916,N_16588);
or U22490 (N_22490,N_19651,N_18590);
nor U22491 (N_22491,N_15412,N_17569);
or U22492 (N_22492,N_16665,N_16964);
nor U22493 (N_22493,N_19928,N_19594);
or U22494 (N_22494,N_18184,N_16294);
nand U22495 (N_22495,N_15732,N_17188);
nand U22496 (N_22496,N_17002,N_19253);
nor U22497 (N_22497,N_18803,N_16110);
nand U22498 (N_22498,N_18434,N_17961);
nand U22499 (N_22499,N_19291,N_19890);
nand U22500 (N_22500,N_19220,N_18450);
and U22501 (N_22501,N_15894,N_19268);
nor U22502 (N_22502,N_16185,N_16686);
or U22503 (N_22503,N_18537,N_16335);
xnor U22504 (N_22504,N_17522,N_17597);
or U22505 (N_22505,N_17948,N_19311);
nand U22506 (N_22506,N_16033,N_16838);
xnor U22507 (N_22507,N_19892,N_18936);
or U22508 (N_22508,N_15412,N_19870);
nand U22509 (N_22509,N_15376,N_17283);
nor U22510 (N_22510,N_19598,N_16398);
nor U22511 (N_22511,N_18661,N_15493);
and U22512 (N_22512,N_16735,N_15216);
nor U22513 (N_22513,N_18722,N_19572);
nor U22514 (N_22514,N_16622,N_19374);
and U22515 (N_22515,N_18115,N_15165);
or U22516 (N_22516,N_19612,N_16636);
and U22517 (N_22517,N_19008,N_16746);
and U22518 (N_22518,N_15692,N_15708);
or U22519 (N_22519,N_19555,N_15157);
nand U22520 (N_22520,N_19088,N_16992);
and U22521 (N_22521,N_15888,N_18093);
or U22522 (N_22522,N_17050,N_19074);
and U22523 (N_22523,N_19189,N_17943);
and U22524 (N_22524,N_15540,N_15393);
and U22525 (N_22525,N_16548,N_16186);
nand U22526 (N_22526,N_15983,N_15245);
nand U22527 (N_22527,N_19505,N_16828);
or U22528 (N_22528,N_18588,N_17268);
nor U22529 (N_22529,N_18505,N_15784);
or U22530 (N_22530,N_16208,N_17826);
and U22531 (N_22531,N_18594,N_16385);
nor U22532 (N_22532,N_18220,N_19751);
nor U22533 (N_22533,N_18161,N_17961);
nor U22534 (N_22534,N_18073,N_18889);
nor U22535 (N_22535,N_18384,N_19934);
nor U22536 (N_22536,N_15614,N_15298);
or U22537 (N_22537,N_16154,N_16761);
nor U22538 (N_22538,N_17437,N_19024);
and U22539 (N_22539,N_15549,N_17268);
or U22540 (N_22540,N_15073,N_15225);
nand U22541 (N_22541,N_16187,N_18949);
nand U22542 (N_22542,N_18949,N_16362);
nand U22543 (N_22543,N_15888,N_18256);
or U22544 (N_22544,N_19415,N_16584);
nor U22545 (N_22545,N_15931,N_16408);
and U22546 (N_22546,N_17870,N_19904);
and U22547 (N_22547,N_16855,N_16362);
nand U22548 (N_22548,N_18149,N_19148);
nand U22549 (N_22549,N_15844,N_15823);
and U22550 (N_22550,N_17789,N_18261);
and U22551 (N_22551,N_15666,N_18673);
and U22552 (N_22552,N_16958,N_19106);
or U22553 (N_22553,N_18007,N_15157);
nor U22554 (N_22554,N_19807,N_19211);
or U22555 (N_22555,N_19590,N_19130);
xor U22556 (N_22556,N_19687,N_18083);
xnor U22557 (N_22557,N_16412,N_18792);
and U22558 (N_22558,N_18559,N_16738);
nor U22559 (N_22559,N_16567,N_18997);
and U22560 (N_22560,N_18926,N_15188);
nor U22561 (N_22561,N_17727,N_15788);
or U22562 (N_22562,N_17809,N_15936);
or U22563 (N_22563,N_16820,N_16913);
nor U22564 (N_22564,N_17150,N_19117);
or U22565 (N_22565,N_17839,N_19150);
and U22566 (N_22566,N_16131,N_15530);
nor U22567 (N_22567,N_18069,N_17575);
and U22568 (N_22568,N_18940,N_16803);
nand U22569 (N_22569,N_15455,N_15992);
and U22570 (N_22570,N_17310,N_17725);
or U22571 (N_22571,N_17093,N_18718);
or U22572 (N_22572,N_17704,N_18203);
nand U22573 (N_22573,N_18444,N_19186);
or U22574 (N_22574,N_19357,N_16763);
and U22575 (N_22575,N_15961,N_18549);
or U22576 (N_22576,N_19073,N_16745);
or U22577 (N_22577,N_15987,N_19122);
nand U22578 (N_22578,N_15227,N_16168);
or U22579 (N_22579,N_16103,N_18891);
nor U22580 (N_22580,N_17877,N_19711);
and U22581 (N_22581,N_16211,N_16743);
or U22582 (N_22582,N_15456,N_15609);
nor U22583 (N_22583,N_17767,N_15877);
nand U22584 (N_22584,N_17991,N_19341);
nand U22585 (N_22585,N_18427,N_17176);
nor U22586 (N_22586,N_19877,N_17799);
nor U22587 (N_22587,N_17423,N_16037);
and U22588 (N_22588,N_17568,N_18848);
nor U22589 (N_22589,N_16353,N_17892);
nor U22590 (N_22590,N_15603,N_17696);
and U22591 (N_22591,N_19273,N_16379);
or U22592 (N_22592,N_19986,N_18302);
nand U22593 (N_22593,N_19915,N_18198);
or U22594 (N_22594,N_16160,N_18015);
nand U22595 (N_22595,N_19332,N_18525);
xor U22596 (N_22596,N_17541,N_17722);
and U22597 (N_22597,N_16081,N_16068);
or U22598 (N_22598,N_15974,N_16881);
nand U22599 (N_22599,N_17255,N_17389);
and U22600 (N_22600,N_16965,N_17329);
xor U22601 (N_22601,N_16501,N_17349);
nand U22602 (N_22602,N_17813,N_16103);
or U22603 (N_22603,N_19004,N_16378);
or U22604 (N_22604,N_18459,N_15046);
nand U22605 (N_22605,N_19349,N_17312);
or U22606 (N_22606,N_17390,N_15433);
and U22607 (N_22607,N_16956,N_19490);
nand U22608 (N_22608,N_17478,N_19715);
nand U22609 (N_22609,N_17867,N_16503);
and U22610 (N_22610,N_18086,N_17393);
or U22611 (N_22611,N_16224,N_16323);
nor U22612 (N_22612,N_19607,N_18079);
or U22613 (N_22613,N_19129,N_15677);
nand U22614 (N_22614,N_19899,N_18370);
xor U22615 (N_22615,N_18836,N_16749);
and U22616 (N_22616,N_19556,N_18994);
and U22617 (N_22617,N_15866,N_19123);
or U22618 (N_22618,N_15490,N_15476);
or U22619 (N_22619,N_19701,N_17395);
and U22620 (N_22620,N_17104,N_16760);
and U22621 (N_22621,N_16139,N_17272);
nor U22622 (N_22622,N_15952,N_17179);
nand U22623 (N_22623,N_16510,N_15882);
nor U22624 (N_22624,N_19652,N_15964);
and U22625 (N_22625,N_15395,N_19618);
and U22626 (N_22626,N_17014,N_17617);
nor U22627 (N_22627,N_18406,N_19858);
nor U22628 (N_22628,N_16119,N_17620);
nor U22629 (N_22629,N_19149,N_16538);
or U22630 (N_22630,N_19006,N_15724);
nand U22631 (N_22631,N_19804,N_16402);
nor U22632 (N_22632,N_16929,N_15324);
nor U22633 (N_22633,N_18367,N_19538);
or U22634 (N_22634,N_18211,N_17191);
nand U22635 (N_22635,N_15396,N_18085);
and U22636 (N_22636,N_18296,N_16852);
xor U22637 (N_22637,N_17926,N_18265);
and U22638 (N_22638,N_16200,N_17273);
or U22639 (N_22639,N_18437,N_18680);
or U22640 (N_22640,N_18366,N_18439);
nand U22641 (N_22641,N_15395,N_16391);
nand U22642 (N_22642,N_17508,N_16835);
nor U22643 (N_22643,N_19399,N_19359);
nand U22644 (N_22644,N_17921,N_15551);
xor U22645 (N_22645,N_16757,N_16314);
or U22646 (N_22646,N_17129,N_17081);
nand U22647 (N_22647,N_16208,N_19243);
or U22648 (N_22648,N_16989,N_17092);
or U22649 (N_22649,N_18762,N_18558);
or U22650 (N_22650,N_15159,N_16722);
or U22651 (N_22651,N_18189,N_15236);
or U22652 (N_22652,N_16825,N_15632);
nand U22653 (N_22653,N_16162,N_19170);
nand U22654 (N_22654,N_17932,N_18964);
or U22655 (N_22655,N_16341,N_16291);
nor U22656 (N_22656,N_18235,N_15624);
or U22657 (N_22657,N_19058,N_19917);
and U22658 (N_22658,N_16702,N_15939);
nor U22659 (N_22659,N_19175,N_18638);
xnor U22660 (N_22660,N_19709,N_16065);
nand U22661 (N_22661,N_19423,N_16748);
nand U22662 (N_22662,N_18415,N_18824);
and U22663 (N_22663,N_17689,N_16044);
nand U22664 (N_22664,N_17896,N_16878);
and U22665 (N_22665,N_19398,N_18034);
and U22666 (N_22666,N_17876,N_18373);
and U22667 (N_22667,N_16712,N_17211);
nor U22668 (N_22668,N_15449,N_19510);
nand U22669 (N_22669,N_18145,N_17810);
nor U22670 (N_22670,N_18860,N_19913);
nor U22671 (N_22671,N_16979,N_19434);
nor U22672 (N_22672,N_16401,N_17122);
or U22673 (N_22673,N_17203,N_17578);
and U22674 (N_22674,N_16701,N_16998);
or U22675 (N_22675,N_19783,N_15621);
and U22676 (N_22676,N_19836,N_17894);
and U22677 (N_22677,N_17350,N_19246);
and U22678 (N_22678,N_15881,N_17781);
nor U22679 (N_22679,N_16749,N_18103);
nand U22680 (N_22680,N_15067,N_17642);
or U22681 (N_22681,N_19826,N_17324);
or U22682 (N_22682,N_19865,N_18746);
nor U22683 (N_22683,N_18593,N_15501);
and U22684 (N_22684,N_19952,N_16203);
and U22685 (N_22685,N_18814,N_17211);
nand U22686 (N_22686,N_16884,N_16517);
nor U22687 (N_22687,N_17725,N_15076);
or U22688 (N_22688,N_19340,N_19835);
and U22689 (N_22689,N_18264,N_16589);
nand U22690 (N_22690,N_18405,N_17740);
nor U22691 (N_22691,N_19395,N_16834);
and U22692 (N_22692,N_16263,N_16043);
nor U22693 (N_22693,N_19739,N_15918);
nand U22694 (N_22694,N_18185,N_15127);
nand U22695 (N_22695,N_18552,N_15816);
nor U22696 (N_22696,N_17602,N_19557);
and U22697 (N_22697,N_16689,N_18051);
and U22698 (N_22698,N_17387,N_16743);
or U22699 (N_22699,N_18606,N_15026);
and U22700 (N_22700,N_15228,N_16313);
or U22701 (N_22701,N_16200,N_18093);
nand U22702 (N_22702,N_19536,N_19518);
nor U22703 (N_22703,N_15383,N_19303);
nand U22704 (N_22704,N_15653,N_18256);
or U22705 (N_22705,N_18185,N_18626);
and U22706 (N_22706,N_15230,N_16565);
and U22707 (N_22707,N_17315,N_19606);
nand U22708 (N_22708,N_18985,N_16236);
nand U22709 (N_22709,N_16413,N_15990);
or U22710 (N_22710,N_15778,N_16077);
nor U22711 (N_22711,N_16473,N_18095);
or U22712 (N_22712,N_19528,N_18861);
and U22713 (N_22713,N_16636,N_19517);
nand U22714 (N_22714,N_17863,N_15031);
nor U22715 (N_22715,N_17323,N_16352);
nor U22716 (N_22716,N_15902,N_16314);
nand U22717 (N_22717,N_18065,N_19091);
nor U22718 (N_22718,N_16064,N_19591);
or U22719 (N_22719,N_17079,N_19635);
nor U22720 (N_22720,N_15830,N_15371);
nor U22721 (N_22721,N_16214,N_16353);
or U22722 (N_22722,N_15821,N_18362);
nor U22723 (N_22723,N_18962,N_15758);
nand U22724 (N_22724,N_16563,N_19995);
and U22725 (N_22725,N_18786,N_19082);
or U22726 (N_22726,N_15397,N_17839);
nand U22727 (N_22727,N_17235,N_17749);
xor U22728 (N_22728,N_15668,N_19743);
nand U22729 (N_22729,N_15848,N_15167);
or U22730 (N_22730,N_17614,N_15647);
and U22731 (N_22731,N_15852,N_18635);
and U22732 (N_22732,N_19999,N_16731);
or U22733 (N_22733,N_18940,N_16181);
and U22734 (N_22734,N_15028,N_15722);
or U22735 (N_22735,N_15581,N_19107);
or U22736 (N_22736,N_19889,N_16156);
or U22737 (N_22737,N_17703,N_15311);
and U22738 (N_22738,N_18030,N_17476);
or U22739 (N_22739,N_19710,N_18230);
and U22740 (N_22740,N_16907,N_19798);
and U22741 (N_22741,N_16063,N_19241);
xnor U22742 (N_22742,N_17160,N_17287);
nand U22743 (N_22743,N_16112,N_19363);
or U22744 (N_22744,N_17534,N_15560);
nand U22745 (N_22745,N_15429,N_19020);
nor U22746 (N_22746,N_15599,N_16197);
and U22747 (N_22747,N_17399,N_17031);
nand U22748 (N_22748,N_16147,N_16527);
and U22749 (N_22749,N_16762,N_18538);
nand U22750 (N_22750,N_16505,N_17938);
nor U22751 (N_22751,N_17618,N_19499);
and U22752 (N_22752,N_17249,N_15236);
nand U22753 (N_22753,N_17507,N_19376);
and U22754 (N_22754,N_16419,N_15842);
or U22755 (N_22755,N_19583,N_17228);
or U22756 (N_22756,N_19872,N_15233);
and U22757 (N_22757,N_18023,N_18152);
nor U22758 (N_22758,N_16969,N_15255);
or U22759 (N_22759,N_16031,N_17135);
nand U22760 (N_22760,N_15036,N_15824);
or U22761 (N_22761,N_16325,N_17438);
and U22762 (N_22762,N_19075,N_16854);
and U22763 (N_22763,N_15479,N_16445);
nand U22764 (N_22764,N_19047,N_18499);
nand U22765 (N_22765,N_16054,N_15970);
nor U22766 (N_22766,N_18286,N_16609);
and U22767 (N_22767,N_16588,N_18329);
or U22768 (N_22768,N_15053,N_19842);
nor U22769 (N_22769,N_15212,N_17886);
nor U22770 (N_22770,N_16507,N_19178);
or U22771 (N_22771,N_16224,N_18291);
nand U22772 (N_22772,N_17704,N_19296);
nor U22773 (N_22773,N_16902,N_18185);
nand U22774 (N_22774,N_15272,N_16874);
nand U22775 (N_22775,N_16594,N_16908);
and U22776 (N_22776,N_16353,N_16873);
or U22777 (N_22777,N_15038,N_18869);
nand U22778 (N_22778,N_17809,N_17332);
nor U22779 (N_22779,N_16089,N_17186);
nor U22780 (N_22780,N_16792,N_15058);
nand U22781 (N_22781,N_19477,N_16652);
and U22782 (N_22782,N_16924,N_19875);
nor U22783 (N_22783,N_17925,N_16940);
nand U22784 (N_22784,N_19902,N_18201);
xor U22785 (N_22785,N_17584,N_17439);
and U22786 (N_22786,N_18490,N_17497);
nand U22787 (N_22787,N_17687,N_16448);
nand U22788 (N_22788,N_17048,N_15165);
or U22789 (N_22789,N_15074,N_16869);
or U22790 (N_22790,N_17101,N_19393);
and U22791 (N_22791,N_18568,N_18678);
nand U22792 (N_22792,N_17068,N_17959);
xor U22793 (N_22793,N_18871,N_16110);
nand U22794 (N_22794,N_16928,N_18530);
nor U22795 (N_22795,N_17080,N_17818);
or U22796 (N_22796,N_18707,N_18406);
nand U22797 (N_22797,N_16604,N_18180);
nor U22798 (N_22798,N_17893,N_16028);
nor U22799 (N_22799,N_16802,N_18023);
nand U22800 (N_22800,N_15817,N_16412);
nor U22801 (N_22801,N_19429,N_19696);
or U22802 (N_22802,N_17860,N_19227);
and U22803 (N_22803,N_18771,N_17010);
nand U22804 (N_22804,N_17028,N_18404);
nor U22805 (N_22805,N_16383,N_18862);
nand U22806 (N_22806,N_19034,N_17898);
or U22807 (N_22807,N_17213,N_16787);
nand U22808 (N_22808,N_19646,N_16350);
or U22809 (N_22809,N_19862,N_18323);
or U22810 (N_22810,N_19051,N_16899);
or U22811 (N_22811,N_18556,N_17553);
or U22812 (N_22812,N_18472,N_16961);
nand U22813 (N_22813,N_18861,N_18352);
nand U22814 (N_22814,N_15980,N_19869);
nand U22815 (N_22815,N_16196,N_15765);
nand U22816 (N_22816,N_18728,N_19118);
or U22817 (N_22817,N_19180,N_17386);
or U22818 (N_22818,N_15516,N_15673);
and U22819 (N_22819,N_15643,N_17511);
or U22820 (N_22820,N_17717,N_18410);
or U22821 (N_22821,N_16029,N_18159);
xor U22822 (N_22822,N_18352,N_15735);
or U22823 (N_22823,N_15195,N_16870);
nand U22824 (N_22824,N_16624,N_16385);
or U22825 (N_22825,N_16836,N_15531);
and U22826 (N_22826,N_19831,N_15098);
nand U22827 (N_22827,N_17372,N_15741);
or U22828 (N_22828,N_19164,N_15997);
or U22829 (N_22829,N_19245,N_19000);
nand U22830 (N_22830,N_18674,N_15235);
and U22831 (N_22831,N_17993,N_19843);
and U22832 (N_22832,N_18224,N_18098);
or U22833 (N_22833,N_16855,N_16148);
nor U22834 (N_22834,N_17214,N_16757);
nor U22835 (N_22835,N_15982,N_15598);
nor U22836 (N_22836,N_18611,N_17365);
nor U22837 (N_22837,N_18021,N_19246);
and U22838 (N_22838,N_15901,N_18632);
and U22839 (N_22839,N_19165,N_17952);
or U22840 (N_22840,N_18647,N_15081);
and U22841 (N_22841,N_15144,N_16875);
nor U22842 (N_22842,N_18755,N_18131);
nand U22843 (N_22843,N_15485,N_19180);
nand U22844 (N_22844,N_17666,N_19850);
nand U22845 (N_22845,N_16853,N_15058);
nor U22846 (N_22846,N_15370,N_18275);
nand U22847 (N_22847,N_16043,N_16703);
nand U22848 (N_22848,N_19764,N_19543);
nand U22849 (N_22849,N_17739,N_19278);
nor U22850 (N_22850,N_19303,N_19740);
and U22851 (N_22851,N_16198,N_18473);
or U22852 (N_22852,N_15533,N_16293);
or U22853 (N_22853,N_16016,N_18130);
and U22854 (N_22854,N_17136,N_17515);
nor U22855 (N_22855,N_15917,N_17770);
and U22856 (N_22856,N_19722,N_15313);
or U22857 (N_22857,N_19251,N_18749);
nor U22858 (N_22858,N_17950,N_15242);
nor U22859 (N_22859,N_19962,N_18600);
nor U22860 (N_22860,N_17571,N_19074);
nor U22861 (N_22861,N_16243,N_19728);
nor U22862 (N_22862,N_17026,N_19849);
and U22863 (N_22863,N_18659,N_15515);
nor U22864 (N_22864,N_19767,N_18453);
or U22865 (N_22865,N_19232,N_18136);
nor U22866 (N_22866,N_17469,N_18086);
or U22867 (N_22867,N_15780,N_17393);
and U22868 (N_22868,N_18076,N_18872);
and U22869 (N_22869,N_18519,N_16140);
and U22870 (N_22870,N_18642,N_18746);
or U22871 (N_22871,N_15179,N_18374);
or U22872 (N_22872,N_17239,N_18399);
and U22873 (N_22873,N_15107,N_15820);
and U22874 (N_22874,N_16686,N_15947);
and U22875 (N_22875,N_16405,N_19947);
or U22876 (N_22876,N_18471,N_16228);
nor U22877 (N_22877,N_18476,N_19890);
nand U22878 (N_22878,N_19007,N_15499);
or U22879 (N_22879,N_18406,N_18928);
nor U22880 (N_22880,N_17491,N_16385);
nand U22881 (N_22881,N_16918,N_19561);
or U22882 (N_22882,N_15251,N_15983);
or U22883 (N_22883,N_16629,N_15499);
nand U22884 (N_22884,N_15318,N_18526);
or U22885 (N_22885,N_16145,N_17410);
nor U22886 (N_22886,N_19100,N_17044);
nor U22887 (N_22887,N_15514,N_18521);
and U22888 (N_22888,N_15284,N_15233);
nor U22889 (N_22889,N_15131,N_18886);
and U22890 (N_22890,N_18125,N_19087);
nand U22891 (N_22891,N_17085,N_19463);
nand U22892 (N_22892,N_16648,N_17693);
or U22893 (N_22893,N_15242,N_16203);
and U22894 (N_22894,N_18695,N_16706);
nor U22895 (N_22895,N_16741,N_16048);
and U22896 (N_22896,N_18586,N_16390);
nor U22897 (N_22897,N_17212,N_18026);
or U22898 (N_22898,N_18073,N_17617);
nor U22899 (N_22899,N_16082,N_17635);
nor U22900 (N_22900,N_19759,N_19387);
nor U22901 (N_22901,N_19530,N_16581);
nor U22902 (N_22902,N_15204,N_15709);
nand U22903 (N_22903,N_18595,N_18049);
nand U22904 (N_22904,N_16924,N_15614);
nor U22905 (N_22905,N_19433,N_15477);
nor U22906 (N_22906,N_16419,N_16230);
nand U22907 (N_22907,N_16906,N_18943);
xnor U22908 (N_22908,N_15519,N_17530);
nor U22909 (N_22909,N_16513,N_15253);
or U22910 (N_22910,N_17566,N_15341);
or U22911 (N_22911,N_17760,N_17294);
nand U22912 (N_22912,N_19499,N_17774);
nor U22913 (N_22913,N_17725,N_18789);
and U22914 (N_22914,N_18892,N_15686);
nor U22915 (N_22915,N_17398,N_18019);
nor U22916 (N_22916,N_18163,N_16172);
or U22917 (N_22917,N_15567,N_19347);
or U22918 (N_22918,N_16389,N_15116);
or U22919 (N_22919,N_16910,N_19134);
and U22920 (N_22920,N_15348,N_18143);
xnor U22921 (N_22921,N_19326,N_19718);
nand U22922 (N_22922,N_17504,N_18212);
nor U22923 (N_22923,N_15844,N_19789);
nor U22924 (N_22924,N_17843,N_16016);
or U22925 (N_22925,N_18046,N_18529);
and U22926 (N_22926,N_15321,N_15283);
nor U22927 (N_22927,N_19055,N_17234);
or U22928 (N_22928,N_17393,N_18720);
nor U22929 (N_22929,N_19456,N_17092);
and U22930 (N_22930,N_18062,N_17986);
or U22931 (N_22931,N_16315,N_18830);
nor U22932 (N_22932,N_18627,N_19444);
nand U22933 (N_22933,N_16832,N_16578);
nand U22934 (N_22934,N_18490,N_16424);
nor U22935 (N_22935,N_16380,N_18432);
or U22936 (N_22936,N_15991,N_19863);
and U22937 (N_22937,N_15165,N_15763);
and U22938 (N_22938,N_17644,N_18862);
or U22939 (N_22939,N_19437,N_19897);
or U22940 (N_22940,N_15991,N_19143);
nor U22941 (N_22941,N_17041,N_16291);
or U22942 (N_22942,N_17920,N_18431);
and U22943 (N_22943,N_19051,N_15969);
nand U22944 (N_22944,N_16959,N_17823);
or U22945 (N_22945,N_17350,N_15640);
nand U22946 (N_22946,N_16781,N_15056);
or U22947 (N_22947,N_19364,N_19135);
nand U22948 (N_22948,N_15825,N_15962);
nor U22949 (N_22949,N_19527,N_16414);
or U22950 (N_22950,N_19432,N_16659);
or U22951 (N_22951,N_16609,N_19726);
or U22952 (N_22952,N_18355,N_15110);
or U22953 (N_22953,N_16252,N_15390);
nand U22954 (N_22954,N_17883,N_16475);
or U22955 (N_22955,N_17967,N_19916);
and U22956 (N_22956,N_16235,N_19591);
nor U22957 (N_22957,N_17701,N_15674);
or U22958 (N_22958,N_19585,N_18177);
and U22959 (N_22959,N_16306,N_15548);
nand U22960 (N_22960,N_15767,N_19202);
nand U22961 (N_22961,N_18177,N_18649);
or U22962 (N_22962,N_17760,N_18065);
nand U22963 (N_22963,N_15576,N_16644);
and U22964 (N_22964,N_15282,N_15000);
and U22965 (N_22965,N_18798,N_19825);
and U22966 (N_22966,N_18463,N_19201);
nand U22967 (N_22967,N_15590,N_16157);
or U22968 (N_22968,N_17992,N_19216);
nand U22969 (N_22969,N_16639,N_18738);
nand U22970 (N_22970,N_16050,N_18340);
xnor U22971 (N_22971,N_19183,N_16616);
or U22972 (N_22972,N_16800,N_16160);
and U22973 (N_22973,N_16648,N_18623);
nand U22974 (N_22974,N_18709,N_15792);
nor U22975 (N_22975,N_16302,N_15648);
and U22976 (N_22976,N_15777,N_16262);
and U22977 (N_22977,N_19481,N_17356);
or U22978 (N_22978,N_18010,N_15964);
and U22979 (N_22979,N_17084,N_16660);
or U22980 (N_22980,N_19669,N_19122);
nand U22981 (N_22981,N_16086,N_19208);
or U22982 (N_22982,N_15950,N_18085);
nor U22983 (N_22983,N_15214,N_18167);
or U22984 (N_22984,N_17662,N_16876);
nand U22985 (N_22985,N_16906,N_19650);
or U22986 (N_22986,N_17566,N_17639);
or U22987 (N_22987,N_16179,N_19744);
and U22988 (N_22988,N_16261,N_15610);
or U22989 (N_22989,N_16420,N_17678);
nor U22990 (N_22990,N_18510,N_15726);
and U22991 (N_22991,N_17575,N_15602);
nand U22992 (N_22992,N_16035,N_17494);
nor U22993 (N_22993,N_17348,N_19583);
nand U22994 (N_22994,N_19981,N_15651);
or U22995 (N_22995,N_18807,N_18542);
nand U22996 (N_22996,N_16685,N_16026);
and U22997 (N_22997,N_15654,N_19126);
nor U22998 (N_22998,N_16996,N_19636);
and U22999 (N_22999,N_16906,N_15473);
or U23000 (N_23000,N_19695,N_15646);
nor U23001 (N_23001,N_15454,N_19456);
and U23002 (N_23002,N_17663,N_19351);
or U23003 (N_23003,N_15351,N_15536);
nand U23004 (N_23004,N_15956,N_18365);
or U23005 (N_23005,N_16511,N_19570);
or U23006 (N_23006,N_15827,N_16653);
nor U23007 (N_23007,N_17519,N_17559);
and U23008 (N_23008,N_16464,N_17083);
nand U23009 (N_23009,N_17596,N_15767);
nor U23010 (N_23010,N_17245,N_18141);
xor U23011 (N_23011,N_15046,N_19480);
nor U23012 (N_23012,N_16867,N_19639);
nand U23013 (N_23013,N_17585,N_16479);
nand U23014 (N_23014,N_19066,N_19638);
or U23015 (N_23015,N_18232,N_15896);
nand U23016 (N_23016,N_15672,N_19166);
nor U23017 (N_23017,N_17508,N_15484);
nand U23018 (N_23018,N_19786,N_16926);
or U23019 (N_23019,N_17432,N_17891);
and U23020 (N_23020,N_16752,N_15867);
or U23021 (N_23021,N_17043,N_15835);
nand U23022 (N_23022,N_15292,N_16752);
and U23023 (N_23023,N_18880,N_18217);
or U23024 (N_23024,N_18994,N_16818);
and U23025 (N_23025,N_15638,N_15460);
nand U23026 (N_23026,N_15491,N_16939);
or U23027 (N_23027,N_19760,N_15052);
and U23028 (N_23028,N_17363,N_17441);
and U23029 (N_23029,N_15462,N_16272);
and U23030 (N_23030,N_18685,N_17531);
or U23031 (N_23031,N_15941,N_15130);
or U23032 (N_23032,N_15438,N_15573);
or U23033 (N_23033,N_18217,N_17057);
nor U23034 (N_23034,N_17096,N_17841);
nor U23035 (N_23035,N_17144,N_19224);
or U23036 (N_23036,N_15834,N_15809);
nor U23037 (N_23037,N_19438,N_15825);
nor U23038 (N_23038,N_19358,N_16046);
nand U23039 (N_23039,N_15685,N_15715);
or U23040 (N_23040,N_15974,N_15800);
nor U23041 (N_23041,N_16299,N_19666);
nand U23042 (N_23042,N_16472,N_15298);
or U23043 (N_23043,N_15984,N_19770);
nor U23044 (N_23044,N_18916,N_16539);
nand U23045 (N_23045,N_18139,N_17952);
nor U23046 (N_23046,N_17138,N_15248);
or U23047 (N_23047,N_15415,N_18140);
nand U23048 (N_23048,N_15290,N_16400);
nand U23049 (N_23049,N_19244,N_15375);
nor U23050 (N_23050,N_17229,N_15045);
or U23051 (N_23051,N_19591,N_17238);
nand U23052 (N_23052,N_16696,N_19077);
xor U23053 (N_23053,N_17651,N_16349);
or U23054 (N_23054,N_18559,N_16827);
nor U23055 (N_23055,N_17550,N_18818);
nand U23056 (N_23056,N_18716,N_15924);
and U23057 (N_23057,N_15294,N_17967);
nor U23058 (N_23058,N_17688,N_18858);
and U23059 (N_23059,N_16364,N_17589);
nor U23060 (N_23060,N_15647,N_16161);
nor U23061 (N_23061,N_15413,N_18723);
and U23062 (N_23062,N_18009,N_18762);
or U23063 (N_23063,N_17269,N_15381);
and U23064 (N_23064,N_17318,N_17040);
nand U23065 (N_23065,N_19447,N_17031);
nor U23066 (N_23066,N_19794,N_19520);
and U23067 (N_23067,N_18376,N_15631);
and U23068 (N_23068,N_19917,N_19550);
or U23069 (N_23069,N_17666,N_18528);
nor U23070 (N_23070,N_15747,N_17175);
or U23071 (N_23071,N_15478,N_15168);
nor U23072 (N_23072,N_19949,N_17940);
or U23073 (N_23073,N_15977,N_17455);
or U23074 (N_23074,N_16123,N_19446);
or U23075 (N_23075,N_19930,N_18874);
and U23076 (N_23076,N_18564,N_19005);
nand U23077 (N_23077,N_17071,N_15603);
nand U23078 (N_23078,N_15128,N_18170);
nor U23079 (N_23079,N_16144,N_17907);
and U23080 (N_23080,N_15443,N_18567);
nor U23081 (N_23081,N_16222,N_18683);
nor U23082 (N_23082,N_15502,N_17869);
nand U23083 (N_23083,N_18006,N_16316);
nand U23084 (N_23084,N_16772,N_17307);
nand U23085 (N_23085,N_15468,N_18513);
and U23086 (N_23086,N_18297,N_18976);
nand U23087 (N_23087,N_17003,N_18689);
nor U23088 (N_23088,N_16071,N_18567);
or U23089 (N_23089,N_19353,N_16542);
nand U23090 (N_23090,N_18793,N_17050);
and U23091 (N_23091,N_15250,N_17031);
or U23092 (N_23092,N_17416,N_19112);
or U23093 (N_23093,N_17591,N_17628);
nor U23094 (N_23094,N_16831,N_18439);
and U23095 (N_23095,N_17531,N_19639);
nor U23096 (N_23096,N_19944,N_15366);
nor U23097 (N_23097,N_15409,N_17844);
or U23098 (N_23098,N_16786,N_19685);
nor U23099 (N_23099,N_16592,N_17386);
or U23100 (N_23100,N_19903,N_16124);
nand U23101 (N_23101,N_16590,N_19940);
or U23102 (N_23102,N_16137,N_19436);
and U23103 (N_23103,N_19313,N_19955);
and U23104 (N_23104,N_16659,N_18652);
or U23105 (N_23105,N_19585,N_18364);
and U23106 (N_23106,N_15017,N_15190);
and U23107 (N_23107,N_18120,N_19689);
nor U23108 (N_23108,N_16794,N_15310);
nor U23109 (N_23109,N_17614,N_18375);
and U23110 (N_23110,N_15843,N_17765);
or U23111 (N_23111,N_16422,N_19502);
and U23112 (N_23112,N_15933,N_16926);
and U23113 (N_23113,N_18935,N_15030);
or U23114 (N_23114,N_16850,N_16742);
nor U23115 (N_23115,N_16462,N_15964);
or U23116 (N_23116,N_17501,N_19514);
xor U23117 (N_23117,N_19047,N_18655);
nor U23118 (N_23118,N_15602,N_16430);
or U23119 (N_23119,N_18384,N_17005);
nand U23120 (N_23120,N_15590,N_17968);
nand U23121 (N_23121,N_19174,N_16548);
nand U23122 (N_23122,N_15882,N_19968);
or U23123 (N_23123,N_18511,N_16125);
xor U23124 (N_23124,N_15595,N_19252);
or U23125 (N_23125,N_18677,N_17808);
or U23126 (N_23126,N_17970,N_15725);
nand U23127 (N_23127,N_17727,N_18498);
or U23128 (N_23128,N_16036,N_18059);
or U23129 (N_23129,N_17782,N_16835);
and U23130 (N_23130,N_19101,N_17063);
nor U23131 (N_23131,N_16852,N_15803);
or U23132 (N_23132,N_17761,N_16382);
nand U23133 (N_23133,N_18766,N_15089);
nand U23134 (N_23134,N_17755,N_15191);
nand U23135 (N_23135,N_18399,N_19247);
nand U23136 (N_23136,N_17632,N_19690);
nor U23137 (N_23137,N_18541,N_15875);
or U23138 (N_23138,N_18393,N_17316);
nor U23139 (N_23139,N_15509,N_19826);
or U23140 (N_23140,N_18313,N_15553);
and U23141 (N_23141,N_17105,N_18433);
nand U23142 (N_23142,N_18250,N_19252);
and U23143 (N_23143,N_18404,N_15028);
nand U23144 (N_23144,N_19224,N_17838);
or U23145 (N_23145,N_18666,N_18033);
and U23146 (N_23146,N_15007,N_19542);
nor U23147 (N_23147,N_16899,N_15784);
xnor U23148 (N_23148,N_18555,N_15420);
nor U23149 (N_23149,N_17841,N_15961);
or U23150 (N_23150,N_16549,N_19014);
or U23151 (N_23151,N_17183,N_17682);
nand U23152 (N_23152,N_19218,N_18481);
xor U23153 (N_23153,N_17208,N_17236);
and U23154 (N_23154,N_16540,N_17099);
and U23155 (N_23155,N_19769,N_19563);
nand U23156 (N_23156,N_17332,N_15457);
or U23157 (N_23157,N_15927,N_19150);
nand U23158 (N_23158,N_18383,N_19101);
or U23159 (N_23159,N_15597,N_16470);
or U23160 (N_23160,N_18549,N_17690);
nand U23161 (N_23161,N_16510,N_19497);
nand U23162 (N_23162,N_15494,N_18005);
nor U23163 (N_23163,N_17265,N_17313);
nand U23164 (N_23164,N_19970,N_18115);
nand U23165 (N_23165,N_17342,N_15040);
nand U23166 (N_23166,N_18513,N_17501);
and U23167 (N_23167,N_19683,N_16182);
nand U23168 (N_23168,N_18174,N_15692);
and U23169 (N_23169,N_18423,N_17248);
or U23170 (N_23170,N_15772,N_19287);
or U23171 (N_23171,N_15153,N_15208);
or U23172 (N_23172,N_17822,N_19751);
and U23173 (N_23173,N_17389,N_17560);
or U23174 (N_23174,N_18110,N_19683);
nor U23175 (N_23175,N_16746,N_16334);
and U23176 (N_23176,N_15722,N_16010);
and U23177 (N_23177,N_17589,N_19846);
and U23178 (N_23178,N_18024,N_16778);
or U23179 (N_23179,N_19687,N_17885);
or U23180 (N_23180,N_19445,N_19162);
nor U23181 (N_23181,N_17829,N_16832);
and U23182 (N_23182,N_16775,N_18505);
nor U23183 (N_23183,N_15998,N_18960);
or U23184 (N_23184,N_16737,N_15893);
nor U23185 (N_23185,N_17029,N_15234);
nor U23186 (N_23186,N_17206,N_19400);
and U23187 (N_23187,N_17126,N_16303);
nand U23188 (N_23188,N_17754,N_17616);
or U23189 (N_23189,N_17897,N_15751);
nor U23190 (N_23190,N_16869,N_18068);
xor U23191 (N_23191,N_16213,N_15581);
nor U23192 (N_23192,N_16681,N_17613);
and U23193 (N_23193,N_19434,N_16044);
or U23194 (N_23194,N_16253,N_15532);
and U23195 (N_23195,N_16348,N_15408);
nand U23196 (N_23196,N_17701,N_17097);
and U23197 (N_23197,N_15770,N_15840);
nand U23198 (N_23198,N_17049,N_16879);
nand U23199 (N_23199,N_19496,N_16409);
nand U23200 (N_23200,N_19054,N_16894);
and U23201 (N_23201,N_15616,N_18704);
xnor U23202 (N_23202,N_16992,N_16145);
or U23203 (N_23203,N_16352,N_17020);
or U23204 (N_23204,N_16367,N_15810);
nor U23205 (N_23205,N_19633,N_16642);
or U23206 (N_23206,N_15666,N_18111);
nand U23207 (N_23207,N_16781,N_15090);
nand U23208 (N_23208,N_16209,N_19147);
and U23209 (N_23209,N_19013,N_16411);
nand U23210 (N_23210,N_18288,N_15892);
and U23211 (N_23211,N_16242,N_15942);
or U23212 (N_23212,N_17593,N_16821);
nand U23213 (N_23213,N_15547,N_18981);
nor U23214 (N_23214,N_19758,N_15462);
nand U23215 (N_23215,N_17973,N_19695);
and U23216 (N_23216,N_17266,N_17105);
and U23217 (N_23217,N_17629,N_15043);
nor U23218 (N_23218,N_19951,N_17367);
nor U23219 (N_23219,N_16147,N_19721);
or U23220 (N_23220,N_19191,N_19580);
or U23221 (N_23221,N_16974,N_18539);
xnor U23222 (N_23222,N_17206,N_18183);
nand U23223 (N_23223,N_16652,N_15956);
or U23224 (N_23224,N_17079,N_16880);
nand U23225 (N_23225,N_15531,N_17192);
nor U23226 (N_23226,N_16618,N_17845);
nand U23227 (N_23227,N_19783,N_17950);
nand U23228 (N_23228,N_16448,N_16006);
nor U23229 (N_23229,N_15066,N_16130);
nor U23230 (N_23230,N_15238,N_18585);
or U23231 (N_23231,N_19868,N_19829);
or U23232 (N_23232,N_15651,N_16312);
nand U23233 (N_23233,N_17818,N_19232);
and U23234 (N_23234,N_17448,N_15762);
or U23235 (N_23235,N_16808,N_17866);
and U23236 (N_23236,N_16767,N_15787);
nor U23237 (N_23237,N_16307,N_16079);
nand U23238 (N_23238,N_18445,N_17186);
nor U23239 (N_23239,N_15317,N_19931);
nand U23240 (N_23240,N_19866,N_15812);
and U23241 (N_23241,N_17418,N_18177);
nand U23242 (N_23242,N_16300,N_16651);
nor U23243 (N_23243,N_18602,N_15234);
or U23244 (N_23244,N_19216,N_16503);
or U23245 (N_23245,N_18237,N_18097);
nor U23246 (N_23246,N_16613,N_18645);
nand U23247 (N_23247,N_17956,N_17516);
nand U23248 (N_23248,N_18211,N_18129);
and U23249 (N_23249,N_16937,N_16978);
or U23250 (N_23250,N_19739,N_16720);
nor U23251 (N_23251,N_15367,N_19110);
nor U23252 (N_23252,N_19165,N_17292);
nand U23253 (N_23253,N_19551,N_15018);
or U23254 (N_23254,N_16949,N_17902);
and U23255 (N_23255,N_19333,N_16580);
nand U23256 (N_23256,N_17930,N_18467);
nor U23257 (N_23257,N_17300,N_19461);
nand U23258 (N_23258,N_17134,N_17441);
or U23259 (N_23259,N_15361,N_17284);
or U23260 (N_23260,N_15638,N_18753);
and U23261 (N_23261,N_16044,N_16983);
or U23262 (N_23262,N_17863,N_16307);
or U23263 (N_23263,N_15824,N_16278);
nand U23264 (N_23264,N_19418,N_18652);
xor U23265 (N_23265,N_15018,N_19346);
nor U23266 (N_23266,N_15966,N_18980);
or U23267 (N_23267,N_17967,N_16892);
or U23268 (N_23268,N_18512,N_17948);
nand U23269 (N_23269,N_17453,N_15099);
or U23270 (N_23270,N_16106,N_19948);
and U23271 (N_23271,N_16424,N_15506);
or U23272 (N_23272,N_17223,N_19901);
and U23273 (N_23273,N_15747,N_15508);
nor U23274 (N_23274,N_17188,N_15391);
or U23275 (N_23275,N_17537,N_16105);
or U23276 (N_23276,N_18505,N_15123);
or U23277 (N_23277,N_15417,N_16589);
nand U23278 (N_23278,N_17865,N_18237);
nor U23279 (N_23279,N_19908,N_15354);
xor U23280 (N_23280,N_19016,N_18310);
nand U23281 (N_23281,N_17390,N_16509);
nor U23282 (N_23282,N_17072,N_17621);
or U23283 (N_23283,N_15210,N_15966);
or U23284 (N_23284,N_16170,N_17164);
or U23285 (N_23285,N_16854,N_18009);
nor U23286 (N_23286,N_15798,N_17704);
nor U23287 (N_23287,N_15236,N_15957);
nand U23288 (N_23288,N_17090,N_17956);
nor U23289 (N_23289,N_19395,N_15528);
or U23290 (N_23290,N_19233,N_19759);
nor U23291 (N_23291,N_15056,N_18291);
nor U23292 (N_23292,N_16875,N_17897);
nand U23293 (N_23293,N_15384,N_19099);
and U23294 (N_23294,N_15457,N_15456);
and U23295 (N_23295,N_19127,N_15649);
and U23296 (N_23296,N_16404,N_16091);
nor U23297 (N_23297,N_19831,N_18914);
or U23298 (N_23298,N_15879,N_17417);
nand U23299 (N_23299,N_18867,N_17351);
nand U23300 (N_23300,N_16780,N_15874);
or U23301 (N_23301,N_19857,N_16774);
nor U23302 (N_23302,N_16260,N_17353);
and U23303 (N_23303,N_15860,N_15446);
or U23304 (N_23304,N_19731,N_17000);
nand U23305 (N_23305,N_19453,N_18368);
and U23306 (N_23306,N_16844,N_19564);
nand U23307 (N_23307,N_16713,N_15552);
or U23308 (N_23308,N_18010,N_19078);
nand U23309 (N_23309,N_19613,N_18582);
and U23310 (N_23310,N_15211,N_17837);
or U23311 (N_23311,N_15291,N_17334);
and U23312 (N_23312,N_15770,N_15353);
nor U23313 (N_23313,N_18225,N_15856);
or U23314 (N_23314,N_19439,N_16690);
nand U23315 (N_23315,N_16733,N_16000);
or U23316 (N_23316,N_15774,N_16228);
nor U23317 (N_23317,N_16235,N_18808);
nor U23318 (N_23318,N_15553,N_19431);
nand U23319 (N_23319,N_16298,N_17143);
nor U23320 (N_23320,N_18866,N_15088);
or U23321 (N_23321,N_17459,N_17952);
or U23322 (N_23322,N_15485,N_17463);
and U23323 (N_23323,N_17465,N_17108);
nor U23324 (N_23324,N_15402,N_19751);
or U23325 (N_23325,N_17609,N_19230);
or U23326 (N_23326,N_15093,N_15128);
nor U23327 (N_23327,N_17725,N_16409);
nand U23328 (N_23328,N_16886,N_18714);
or U23329 (N_23329,N_17978,N_19508);
nand U23330 (N_23330,N_15674,N_17993);
xnor U23331 (N_23331,N_16821,N_17425);
or U23332 (N_23332,N_19019,N_17369);
or U23333 (N_23333,N_17331,N_16618);
and U23334 (N_23334,N_15171,N_18878);
and U23335 (N_23335,N_15388,N_18413);
xnor U23336 (N_23336,N_15256,N_17563);
nand U23337 (N_23337,N_16991,N_19931);
nor U23338 (N_23338,N_18078,N_18999);
or U23339 (N_23339,N_18592,N_19713);
or U23340 (N_23340,N_18358,N_19285);
and U23341 (N_23341,N_19756,N_19712);
or U23342 (N_23342,N_15548,N_16492);
xnor U23343 (N_23343,N_19849,N_17743);
or U23344 (N_23344,N_15416,N_19037);
and U23345 (N_23345,N_19115,N_16272);
nor U23346 (N_23346,N_17567,N_17411);
nand U23347 (N_23347,N_18271,N_16555);
or U23348 (N_23348,N_16345,N_19622);
nor U23349 (N_23349,N_17427,N_19148);
nor U23350 (N_23350,N_19694,N_15757);
and U23351 (N_23351,N_18900,N_18599);
and U23352 (N_23352,N_15112,N_17118);
nor U23353 (N_23353,N_15760,N_16785);
and U23354 (N_23354,N_19770,N_16207);
nor U23355 (N_23355,N_15890,N_18352);
and U23356 (N_23356,N_19505,N_15849);
xor U23357 (N_23357,N_18035,N_15709);
nor U23358 (N_23358,N_16997,N_18250);
xnor U23359 (N_23359,N_16397,N_18742);
and U23360 (N_23360,N_19851,N_16259);
nand U23361 (N_23361,N_19034,N_16929);
or U23362 (N_23362,N_16640,N_19047);
and U23363 (N_23363,N_17003,N_16122);
and U23364 (N_23364,N_19155,N_19332);
or U23365 (N_23365,N_18483,N_18414);
nand U23366 (N_23366,N_16545,N_17378);
or U23367 (N_23367,N_16656,N_15410);
nand U23368 (N_23368,N_16877,N_15434);
and U23369 (N_23369,N_16744,N_19975);
or U23370 (N_23370,N_19604,N_19349);
xnor U23371 (N_23371,N_17945,N_16982);
or U23372 (N_23372,N_19401,N_19702);
and U23373 (N_23373,N_16781,N_16886);
or U23374 (N_23374,N_17579,N_18961);
and U23375 (N_23375,N_16881,N_16000);
and U23376 (N_23376,N_19793,N_18868);
nor U23377 (N_23377,N_16149,N_15041);
nand U23378 (N_23378,N_17699,N_19858);
nand U23379 (N_23379,N_15003,N_17667);
and U23380 (N_23380,N_19377,N_17272);
and U23381 (N_23381,N_15293,N_17579);
and U23382 (N_23382,N_19327,N_19862);
nor U23383 (N_23383,N_17934,N_18109);
nand U23384 (N_23384,N_15809,N_17815);
nand U23385 (N_23385,N_17685,N_18302);
xnor U23386 (N_23386,N_16434,N_17271);
nor U23387 (N_23387,N_19762,N_15487);
and U23388 (N_23388,N_15270,N_16078);
nand U23389 (N_23389,N_15733,N_17119);
nor U23390 (N_23390,N_17354,N_18142);
nor U23391 (N_23391,N_16795,N_15707);
and U23392 (N_23392,N_19377,N_19042);
or U23393 (N_23393,N_18423,N_18081);
or U23394 (N_23394,N_19221,N_17986);
nand U23395 (N_23395,N_16064,N_15863);
xnor U23396 (N_23396,N_15674,N_15770);
nor U23397 (N_23397,N_16001,N_17504);
xor U23398 (N_23398,N_19460,N_15796);
nor U23399 (N_23399,N_19879,N_19040);
nand U23400 (N_23400,N_18205,N_17126);
nor U23401 (N_23401,N_18489,N_17478);
nand U23402 (N_23402,N_16538,N_15420);
and U23403 (N_23403,N_17438,N_16386);
nor U23404 (N_23404,N_15776,N_19487);
nand U23405 (N_23405,N_16341,N_17268);
or U23406 (N_23406,N_15459,N_15227);
and U23407 (N_23407,N_16523,N_15435);
nand U23408 (N_23408,N_15322,N_16884);
nand U23409 (N_23409,N_19838,N_18597);
nand U23410 (N_23410,N_15340,N_16422);
or U23411 (N_23411,N_16785,N_17553);
or U23412 (N_23412,N_16606,N_15652);
xor U23413 (N_23413,N_16151,N_15979);
and U23414 (N_23414,N_19335,N_17530);
nor U23415 (N_23415,N_19462,N_19005);
nor U23416 (N_23416,N_17945,N_15557);
and U23417 (N_23417,N_17970,N_18748);
and U23418 (N_23418,N_17697,N_19686);
nand U23419 (N_23419,N_18687,N_17607);
nor U23420 (N_23420,N_15107,N_17997);
or U23421 (N_23421,N_19485,N_19606);
nand U23422 (N_23422,N_18261,N_16252);
and U23423 (N_23423,N_19173,N_16266);
xor U23424 (N_23424,N_17335,N_19546);
nand U23425 (N_23425,N_18078,N_17952);
and U23426 (N_23426,N_19759,N_16527);
nand U23427 (N_23427,N_16048,N_18755);
nand U23428 (N_23428,N_16161,N_15138);
or U23429 (N_23429,N_18749,N_19387);
and U23430 (N_23430,N_15815,N_18916);
nor U23431 (N_23431,N_19146,N_15177);
nor U23432 (N_23432,N_17100,N_17277);
or U23433 (N_23433,N_17466,N_17874);
and U23434 (N_23434,N_19093,N_15776);
nor U23435 (N_23435,N_19294,N_18712);
and U23436 (N_23436,N_18236,N_19381);
nor U23437 (N_23437,N_15381,N_15770);
and U23438 (N_23438,N_16490,N_16743);
xnor U23439 (N_23439,N_19488,N_15992);
nand U23440 (N_23440,N_19449,N_16502);
nand U23441 (N_23441,N_19628,N_16124);
and U23442 (N_23442,N_15414,N_17686);
nor U23443 (N_23443,N_17682,N_17118);
and U23444 (N_23444,N_16678,N_17562);
nand U23445 (N_23445,N_17779,N_19770);
and U23446 (N_23446,N_16016,N_16523);
nand U23447 (N_23447,N_15515,N_17822);
nand U23448 (N_23448,N_15024,N_18037);
nand U23449 (N_23449,N_19185,N_18353);
and U23450 (N_23450,N_18259,N_19503);
or U23451 (N_23451,N_15503,N_15771);
nand U23452 (N_23452,N_16806,N_19250);
or U23453 (N_23453,N_16970,N_15941);
and U23454 (N_23454,N_15191,N_19862);
nor U23455 (N_23455,N_15202,N_19151);
nor U23456 (N_23456,N_15623,N_16289);
or U23457 (N_23457,N_17101,N_18626);
or U23458 (N_23458,N_16984,N_17733);
and U23459 (N_23459,N_18396,N_18535);
or U23460 (N_23460,N_17237,N_18272);
and U23461 (N_23461,N_16372,N_16129);
nor U23462 (N_23462,N_17139,N_17743);
nor U23463 (N_23463,N_15374,N_17437);
nor U23464 (N_23464,N_15314,N_15362);
or U23465 (N_23465,N_18814,N_17420);
nand U23466 (N_23466,N_16925,N_16617);
nand U23467 (N_23467,N_19342,N_17668);
nor U23468 (N_23468,N_18846,N_16731);
nand U23469 (N_23469,N_15190,N_16905);
or U23470 (N_23470,N_16827,N_17631);
and U23471 (N_23471,N_19862,N_16401);
nand U23472 (N_23472,N_17023,N_19896);
nor U23473 (N_23473,N_16024,N_16881);
and U23474 (N_23474,N_17149,N_18819);
nand U23475 (N_23475,N_16034,N_18596);
nor U23476 (N_23476,N_16894,N_15526);
xor U23477 (N_23477,N_16270,N_16214);
nand U23478 (N_23478,N_19484,N_18504);
nand U23479 (N_23479,N_18611,N_19151);
xor U23480 (N_23480,N_16885,N_16309);
or U23481 (N_23481,N_19878,N_15136);
nand U23482 (N_23482,N_17242,N_15179);
nand U23483 (N_23483,N_18223,N_16748);
or U23484 (N_23484,N_19995,N_16841);
and U23485 (N_23485,N_18049,N_17353);
and U23486 (N_23486,N_15166,N_19249);
nor U23487 (N_23487,N_15374,N_18550);
nor U23488 (N_23488,N_19425,N_19981);
or U23489 (N_23489,N_17015,N_19521);
and U23490 (N_23490,N_16960,N_18485);
and U23491 (N_23491,N_15243,N_15896);
and U23492 (N_23492,N_15810,N_19741);
or U23493 (N_23493,N_17337,N_18438);
nand U23494 (N_23494,N_19662,N_17069);
nand U23495 (N_23495,N_18877,N_15127);
and U23496 (N_23496,N_15436,N_18225);
or U23497 (N_23497,N_16871,N_18369);
nor U23498 (N_23498,N_16215,N_18629);
or U23499 (N_23499,N_19085,N_17394);
nor U23500 (N_23500,N_18236,N_17573);
or U23501 (N_23501,N_19286,N_17566);
nor U23502 (N_23502,N_17063,N_17030);
nand U23503 (N_23503,N_16213,N_15077);
nor U23504 (N_23504,N_16154,N_16203);
nand U23505 (N_23505,N_15669,N_18778);
and U23506 (N_23506,N_19389,N_16248);
nor U23507 (N_23507,N_16833,N_17909);
and U23508 (N_23508,N_18661,N_19886);
and U23509 (N_23509,N_16169,N_15579);
xnor U23510 (N_23510,N_18414,N_18964);
nand U23511 (N_23511,N_15533,N_18819);
or U23512 (N_23512,N_19114,N_19720);
nand U23513 (N_23513,N_17313,N_18772);
and U23514 (N_23514,N_16118,N_18775);
nand U23515 (N_23515,N_18525,N_17417);
and U23516 (N_23516,N_15875,N_18776);
or U23517 (N_23517,N_16075,N_19823);
or U23518 (N_23518,N_18448,N_18401);
or U23519 (N_23519,N_17595,N_16233);
nor U23520 (N_23520,N_19435,N_17476);
or U23521 (N_23521,N_16839,N_15620);
or U23522 (N_23522,N_17152,N_18372);
and U23523 (N_23523,N_19219,N_19275);
nor U23524 (N_23524,N_16970,N_17848);
nand U23525 (N_23525,N_17537,N_17151);
nor U23526 (N_23526,N_15059,N_19901);
or U23527 (N_23527,N_15348,N_18980);
and U23528 (N_23528,N_19694,N_17800);
nor U23529 (N_23529,N_17908,N_15058);
or U23530 (N_23530,N_16545,N_18771);
and U23531 (N_23531,N_16054,N_16712);
nor U23532 (N_23532,N_19670,N_19671);
and U23533 (N_23533,N_18091,N_19572);
and U23534 (N_23534,N_15737,N_17165);
nor U23535 (N_23535,N_15121,N_18186);
and U23536 (N_23536,N_17669,N_17223);
or U23537 (N_23537,N_16067,N_16733);
nand U23538 (N_23538,N_18096,N_16863);
nand U23539 (N_23539,N_19768,N_19561);
and U23540 (N_23540,N_18574,N_15754);
xor U23541 (N_23541,N_18177,N_17420);
nor U23542 (N_23542,N_15235,N_17025);
nand U23543 (N_23543,N_17902,N_15909);
or U23544 (N_23544,N_19782,N_15454);
nand U23545 (N_23545,N_15937,N_16625);
nand U23546 (N_23546,N_18063,N_17180);
nand U23547 (N_23547,N_16144,N_17774);
nor U23548 (N_23548,N_17442,N_17993);
and U23549 (N_23549,N_16930,N_19502);
and U23550 (N_23550,N_16372,N_17367);
and U23551 (N_23551,N_17770,N_19498);
nor U23552 (N_23552,N_19560,N_19581);
nand U23553 (N_23553,N_16705,N_18925);
or U23554 (N_23554,N_18389,N_19429);
nor U23555 (N_23555,N_18034,N_17633);
and U23556 (N_23556,N_18932,N_16354);
nand U23557 (N_23557,N_19121,N_17413);
and U23558 (N_23558,N_17570,N_17665);
and U23559 (N_23559,N_17612,N_17223);
nand U23560 (N_23560,N_18036,N_19965);
and U23561 (N_23561,N_16628,N_18116);
and U23562 (N_23562,N_15327,N_17327);
or U23563 (N_23563,N_15430,N_18791);
nand U23564 (N_23564,N_17443,N_16050);
nor U23565 (N_23565,N_17760,N_18437);
nor U23566 (N_23566,N_16732,N_15180);
nor U23567 (N_23567,N_17013,N_16387);
xnor U23568 (N_23568,N_17140,N_18972);
and U23569 (N_23569,N_18180,N_15683);
nand U23570 (N_23570,N_15528,N_17879);
and U23571 (N_23571,N_16363,N_15006);
or U23572 (N_23572,N_16512,N_19549);
or U23573 (N_23573,N_15146,N_17515);
nor U23574 (N_23574,N_17896,N_16991);
nand U23575 (N_23575,N_16889,N_16611);
and U23576 (N_23576,N_16034,N_19424);
nor U23577 (N_23577,N_18382,N_18167);
xor U23578 (N_23578,N_16422,N_18591);
xor U23579 (N_23579,N_18852,N_19795);
and U23580 (N_23580,N_19997,N_18920);
and U23581 (N_23581,N_19224,N_16952);
or U23582 (N_23582,N_15243,N_19716);
and U23583 (N_23583,N_17594,N_19095);
or U23584 (N_23584,N_16318,N_18334);
xor U23585 (N_23585,N_16618,N_19196);
nand U23586 (N_23586,N_17926,N_17547);
nand U23587 (N_23587,N_17414,N_19137);
or U23588 (N_23588,N_16786,N_18030);
or U23589 (N_23589,N_17957,N_16203);
nand U23590 (N_23590,N_15639,N_16066);
nor U23591 (N_23591,N_15901,N_15419);
nor U23592 (N_23592,N_15608,N_15204);
or U23593 (N_23593,N_17864,N_19715);
and U23594 (N_23594,N_16725,N_16078);
or U23595 (N_23595,N_18179,N_18241);
and U23596 (N_23596,N_19310,N_16592);
or U23597 (N_23597,N_17463,N_18792);
nor U23598 (N_23598,N_19838,N_15982);
or U23599 (N_23599,N_18472,N_19601);
and U23600 (N_23600,N_17625,N_16567);
nor U23601 (N_23601,N_19679,N_19808);
or U23602 (N_23602,N_19332,N_19006);
nand U23603 (N_23603,N_15847,N_19963);
and U23604 (N_23604,N_18234,N_19308);
or U23605 (N_23605,N_16438,N_16494);
or U23606 (N_23606,N_16771,N_16656);
and U23607 (N_23607,N_16165,N_17663);
or U23608 (N_23608,N_16140,N_18175);
or U23609 (N_23609,N_16227,N_18785);
nor U23610 (N_23610,N_17061,N_19144);
or U23611 (N_23611,N_19852,N_17669);
nor U23612 (N_23612,N_18452,N_17117);
or U23613 (N_23613,N_19269,N_18127);
or U23614 (N_23614,N_18627,N_15050);
nor U23615 (N_23615,N_16011,N_19625);
and U23616 (N_23616,N_17789,N_16134);
or U23617 (N_23617,N_16091,N_15098);
nand U23618 (N_23618,N_16280,N_19468);
or U23619 (N_23619,N_16293,N_18489);
nor U23620 (N_23620,N_19052,N_16488);
or U23621 (N_23621,N_17413,N_17556);
nand U23622 (N_23622,N_16180,N_17991);
and U23623 (N_23623,N_16055,N_17996);
and U23624 (N_23624,N_15978,N_15398);
nor U23625 (N_23625,N_16035,N_19356);
or U23626 (N_23626,N_15542,N_19067);
nor U23627 (N_23627,N_19171,N_19925);
nor U23628 (N_23628,N_18111,N_18694);
nor U23629 (N_23629,N_17441,N_17606);
and U23630 (N_23630,N_16926,N_18729);
or U23631 (N_23631,N_17790,N_16481);
nand U23632 (N_23632,N_19733,N_15193);
nor U23633 (N_23633,N_18008,N_16268);
or U23634 (N_23634,N_16395,N_17811);
nor U23635 (N_23635,N_16516,N_19214);
and U23636 (N_23636,N_17803,N_15589);
and U23637 (N_23637,N_19985,N_17298);
and U23638 (N_23638,N_16637,N_17219);
nand U23639 (N_23639,N_18430,N_17636);
nand U23640 (N_23640,N_18214,N_16913);
or U23641 (N_23641,N_15464,N_17700);
or U23642 (N_23642,N_19813,N_17587);
nor U23643 (N_23643,N_18208,N_19614);
and U23644 (N_23644,N_17733,N_19133);
nand U23645 (N_23645,N_19577,N_17388);
and U23646 (N_23646,N_15578,N_18483);
nand U23647 (N_23647,N_18036,N_19749);
or U23648 (N_23648,N_18697,N_18305);
nand U23649 (N_23649,N_15276,N_15089);
nor U23650 (N_23650,N_16010,N_16556);
or U23651 (N_23651,N_18635,N_19232);
nor U23652 (N_23652,N_15077,N_18923);
or U23653 (N_23653,N_18201,N_19226);
or U23654 (N_23654,N_16264,N_18624);
nor U23655 (N_23655,N_19237,N_18981);
nor U23656 (N_23656,N_19619,N_19538);
nand U23657 (N_23657,N_15049,N_19245);
nand U23658 (N_23658,N_17628,N_15222);
and U23659 (N_23659,N_16748,N_15459);
nor U23660 (N_23660,N_19615,N_18027);
or U23661 (N_23661,N_15111,N_17300);
and U23662 (N_23662,N_16461,N_17309);
or U23663 (N_23663,N_18343,N_17822);
nor U23664 (N_23664,N_19241,N_18214);
or U23665 (N_23665,N_19918,N_18975);
and U23666 (N_23666,N_15495,N_17349);
and U23667 (N_23667,N_19757,N_19271);
or U23668 (N_23668,N_16433,N_17417);
nand U23669 (N_23669,N_15371,N_15908);
nand U23670 (N_23670,N_16563,N_16286);
nand U23671 (N_23671,N_15008,N_16659);
or U23672 (N_23672,N_15384,N_19399);
nand U23673 (N_23673,N_16451,N_16599);
nand U23674 (N_23674,N_17536,N_15336);
or U23675 (N_23675,N_16210,N_17163);
nand U23676 (N_23676,N_15759,N_16879);
or U23677 (N_23677,N_19354,N_15580);
nor U23678 (N_23678,N_18564,N_17700);
nand U23679 (N_23679,N_16018,N_16548);
or U23680 (N_23680,N_16241,N_17486);
nand U23681 (N_23681,N_18536,N_17116);
nand U23682 (N_23682,N_16335,N_16654);
and U23683 (N_23683,N_15401,N_18094);
or U23684 (N_23684,N_18193,N_19074);
nand U23685 (N_23685,N_15416,N_16377);
or U23686 (N_23686,N_15979,N_18668);
and U23687 (N_23687,N_17646,N_17545);
nand U23688 (N_23688,N_18640,N_16353);
nand U23689 (N_23689,N_16575,N_18173);
or U23690 (N_23690,N_16285,N_19295);
and U23691 (N_23691,N_17673,N_15111);
nor U23692 (N_23692,N_17458,N_17423);
nand U23693 (N_23693,N_19500,N_19408);
nand U23694 (N_23694,N_16011,N_19212);
and U23695 (N_23695,N_19978,N_19038);
nand U23696 (N_23696,N_16421,N_15704);
xnor U23697 (N_23697,N_19046,N_16764);
and U23698 (N_23698,N_16450,N_18939);
and U23699 (N_23699,N_16356,N_17564);
nand U23700 (N_23700,N_18671,N_15982);
nand U23701 (N_23701,N_18221,N_15131);
nor U23702 (N_23702,N_18191,N_19884);
nor U23703 (N_23703,N_16443,N_17362);
nor U23704 (N_23704,N_19299,N_17520);
or U23705 (N_23705,N_19537,N_16385);
and U23706 (N_23706,N_17162,N_17501);
and U23707 (N_23707,N_18656,N_17454);
or U23708 (N_23708,N_15588,N_15291);
or U23709 (N_23709,N_15373,N_18740);
nor U23710 (N_23710,N_16320,N_16538);
nor U23711 (N_23711,N_17583,N_16060);
and U23712 (N_23712,N_19605,N_17491);
nor U23713 (N_23713,N_15530,N_15504);
nand U23714 (N_23714,N_19589,N_15351);
xnor U23715 (N_23715,N_17856,N_15283);
nor U23716 (N_23716,N_16208,N_17582);
nand U23717 (N_23717,N_18542,N_17224);
or U23718 (N_23718,N_19063,N_15489);
nor U23719 (N_23719,N_18935,N_17179);
or U23720 (N_23720,N_15623,N_17908);
or U23721 (N_23721,N_18918,N_18253);
nor U23722 (N_23722,N_18618,N_18914);
nor U23723 (N_23723,N_16067,N_18375);
and U23724 (N_23724,N_17237,N_19726);
or U23725 (N_23725,N_15969,N_15779);
nor U23726 (N_23726,N_18551,N_19055);
nand U23727 (N_23727,N_19171,N_19768);
and U23728 (N_23728,N_17739,N_17847);
xor U23729 (N_23729,N_16406,N_15022);
and U23730 (N_23730,N_17296,N_15121);
nand U23731 (N_23731,N_18220,N_17835);
nor U23732 (N_23732,N_18755,N_15572);
nand U23733 (N_23733,N_15055,N_17753);
nand U23734 (N_23734,N_16291,N_19829);
xor U23735 (N_23735,N_19695,N_16748);
nor U23736 (N_23736,N_18447,N_16330);
or U23737 (N_23737,N_16325,N_17244);
nor U23738 (N_23738,N_18577,N_19094);
nor U23739 (N_23739,N_17732,N_15197);
or U23740 (N_23740,N_17424,N_15738);
nor U23741 (N_23741,N_18120,N_18649);
and U23742 (N_23742,N_18746,N_18720);
xor U23743 (N_23743,N_18599,N_18551);
or U23744 (N_23744,N_19712,N_16763);
xor U23745 (N_23745,N_16619,N_17818);
nand U23746 (N_23746,N_19820,N_17218);
and U23747 (N_23747,N_19359,N_19467);
or U23748 (N_23748,N_18912,N_15020);
and U23749 (N_23749,N_15993,N_19166);
xnor U23750 (N_23750,N_19345,N_19812);
or U23751 (N_23751,N_19376,N_17864);
nand U23752 (N_23752,N_16897,N_15861);
and U23753 (N_23753,N_16241,N_15894);
or U23754 (N_23754,N_19379,N_18927);
or U23755 (N_23755,N_19605,N_19199);
and U23756 (N_23756,N_17895,N_18205);
and U23757 (N_23757,N_19938,N_18145);
or U23758 (N_23758,N_19582,N_18986);
nand U23759 (N_23759,N_15409,N_17174);
nand U23760 (N_23760,N_19546,N_16370);
and U23761 (N_23761,N_15807,N_15097);
nand U23762 (N_23762,N_18433,N_16061);
or U23763 (N_23763,N_16624,N_17363);
or U23764 (N_23764,N_15958,N_17890);
and U23765 (N_23765,N_15465,N_17562);
nor U23766 (N_23766,N_15159,N_15483);
nor U23767 (N_23767,N_19947,N_16947);
and U23768 (N_23768,N_15124,N_15120);
nand U23769 (N_23769,N_17313,N_18865);
nor U23770 (N_23770,N_18100,N_17651);
nand U23771 (N_23771,N_15683,N_15087);
nand U23772 (N_23772,N_16875,N_18325);
nand U23773 (N_23773,N_17110,N_18470);
nor U23774 (N_23774,N_15636,N_16118);
and U23775 (N_23775,N_19110,N_19436);
xnor U23776 (N_23776,N_15198,N_15683);
or U23777 (N_23777,N_18766,N_16471);
and U23778 (N_23778,N_17412,N_19611);
nand U23779 (N_23779,N_16359,N_19898);
nand U23780 (N_23780,N_18060,N_18451);
nor U23781 (N_23781,N_16814,N_15155);
and U23782 (N_23782,N_19912,N_19234);
and U23783 (N_23783,N_17696,N_16877);
and U23784 (N_23784,N_15004,N_17114);
or U23785 (N_23785,N_17227,N_18454);
and U23786 (N_23786,N_18829,N_16058);
nor U23787 (N_23787,N_15198,N_17900);
nand U23788 (N_23788,N_16691,N_18669);
or U23789 (N_23789,N_16609,N_15068);
nor U23790 (N_23790,N_16725,N_16095);
or U23791 (N_23791,N_18646,N_17857);
nand U23792 (N_23792,N_16220,N_16029);
and U23793 (N_23793,N_17065,N_15547);
nand U23794 (N_23794,N_16376,N_17260);
nand U23795 (N_23795,N_17356,N_16052);
nor U23796 (N_23796,N_16969,N_19856);
xnor U23797 (N_23797,N_19297,N_17759);
and U23798 (N_23798,N_17822,N_15748);
nor U23799 (N_23799,N_17008,N_19103);
nor U23800 (N_23800,N_15547,N_18262);
or U23801 (N_23801,N_19759,N_16502);
nand U23802 (N_23802,N_15668,N_17242);
nand U23803 (N_23803,N_16571,N_17049);
nand U23804 (N_23804,N_19121,N_19154);
and U23805 (N_23805,N_15275,N_17215);
xor U23806 (N_23806,N_18565,N_17509);
nor U23807 (N_23807,N_16541,N_16899);
and U23808 (N_23808,N_18577,N_17395);
nor U23809 (N_23809,N_19509,N_17523);
nand U23810 (N_23810,N_18370,N_16984);
nor U23811 (N_23811,N_18840,N_17489);
xnor U23812 (N_23812,N_19562,N_15003);
nand U23813 (N_23813,N_19755,N_16955);
and U23814 (N_23814,N_18683,N_19934);
nor U23815 (N_23815,N_19435,N_19919);
and U23816 (N_23816,N_19646,N_18164);
nor U23817 (N_23817,N_15480,N_18746);
or U23818 (N_23818,N_18273,N_17700);
or U23819 (N_23819,N_16257,N_15661);
and U23820 (N_23820,N_18373,N_17769);
nor U23821 (N_23821,N_18261,N_18074);
or U23822 (N_23822,N_19280,N_15067);
or U23823 (N_23823,N_17910,N_16999);
or U23824 (N_23824,N_17988,N_17231);
nor U23825 (N_23825,N_15306,N_18830);
and U23826 (N_23826,N_16303,N_15676);
or U23827 (N_23827,N_19155,N_19660);
and U23828 (N_23828,N_16763,N_17773);
nand U23829 (N_23829,N_16274,N_17246);
and U23830 (N_23830,N_17303,N_17149);
and U23831 (N_23831,N_15250,N_17325);
nand U23832 (N_23832,N_16483,N_19276);
or U23833 (N_23833,N_18387,N_17027);
or U23834 (N_23834,N_15569,N_15343);
and U23835 (N_23835,N_19474,N_17241);
nand U23836 (N_23836,N_16308,N_15779);
nor U23837 (N_23837,N_19296,N_16585);
nand U23838 (N_23838,N_16067,N_19810);
and U23839 (N_23839,N_19446,N_16496);
nand U23840 (N_23840,N_17887,N_18311);
nand U23841 (N_23841,N_19313,N_16157);
nor U23842 (N_23842,N_17593,N_17050);
or U23843 (N_23843,N_17578,N_15177);
nand U23844 (N_23844,N_17321,N_17411);
nand U23845 (N_23845,N_15613,N_19001);
nor U23846 (N_23846,N_17962,N_18453);
xor U23847 (N_23847,N_15503,N_18944);
nand U23848 (N_23848,N_15627,N_15950);
xor U23849 (N_23849,N_17354,N_18154);
or U23850 (N_23850,N_17878,N_15915);
nor U23851 (N_23851,N_18207,N_15549);
or U23852 (N_23852,N_15905,N_19517);
or U23853 (N_23853,N_17742,N_15256);
nor U23854 (N_23854,N_15832,N_17993);
or U23855 (N_23855,N_18861,N_17345);
and U23856 (N_23856,N_15181,N_19112);
nand U23857 (N_23857,N_16046,N_16466);
nand U23858 (N_23858,N_17581,N_17358);
or U23859 (N_23859,N_15596,N_15823);
nand U23860 (N_23860,N_18288,N_17393);
or U23861 (N_23861,N_18051,N_16387);
nand U23862 (N_23862,N_17981,N_16632);
nor U23863 (N_23863,N_15098,N_17975);
nor U23864 (N_23864,N_16083,N_17277);
nand U23865 (N_23865,N_16720,N_16251);
nor U23866 (N_23866,N_18357,N_18852);
and U23867 (N_23867,N_15242,N_19806);
or U23868 (N_23868,N_18494,N_16023);
nor U23869 (N_23869,N_17349,N_17199);
nand U23870 (N_23870,N_17285,N_16745);
nor U23871 (N_23871,N_18826,N_15781);
and U23872 (N_23872,N_15002,N_17965);
or U23873 (N_23873,N_15684,N_19215);
and U23874 (N_23874,N_15495,N_18525);
and U23875 (N_23875,N_15395,N_16047);
or U23876 (N_23876,N_19881,N_17147);
nand U23877 (N_23877,N_18819,N_15813);
nor U23878 (N_23878,N_19181,N_18305);
or U23879 (N_23879,N_15240,N_17189);
nor U23880 (N_23880,N_18150,N_15965);
nor U23881 (N_23881,N_16236,N_18541);
nor U23882 (N_23882,N_17095,N_19808);
and U23883 (N_23883,N_15228,N_16243);
nor U23884 (N_23884,N_15612,N_15147);
and U23885 (N_23885,N_17181,N_16658);
nand U23886 (N_23886,N_18700,N_19982);
nor U23887 (N_23887,N_17981,N_17450);
nor U23888 (N_23888,N_16227,N_18380);
nor U23889 (N_23889,N_17122,N_15268);
nand U23890 (N_23890,N_19863,N_17521);
and U23891 (N_23891,N_19086,N_18784);
nand U23892 (N_23892,N_17856,N_18375);
and U23893 (N_23893,N_15349,N_15227);
and U23894 (N_23894,N_16425,N_15035);
nor U23895 (N_23895,N_18940,N_16080);
nor U23896 (N_23896,N_15454,N_16061);
and U23897 (N_23897,N_16964,N_16564);
nor U23898 (N_23898,N_16763,N_17316);
nand U23899 (N_23899,N_17719,N_18234);
and U23900 (N_23900,N_18413,N_15700);
nand U23901 (N_23901,N_15642,N_16311);
nand U23902 (N_23902,N_16477,N_18776);
nor U23903 (N_23903,N_15770,N_17537);
nand U23904 (N_23904,N_15792,N_17658);
or U23905 (N_23905,N_18488,N_18707);
xor U23906 (N_23906,N_17975,N_19227);
and U23907 (N_23907,N_19342,N_19361);
nand U23908 (N_23908,N_18181,N_16556);
xnor U23909 (N_23909,N_19030,N_19020);
and U23910 (N_23910,N_16154,N_16544);
nand U23911 (N_23911,N_17354,N_18271);
nor U23912 (N_23912,N_16103,N_18082);
nor U23913 (N_23913,N_15683,N_18946);
xnor U23914 (N_23914,N_15157,N_16645);
nand U23915 (N_23915,N_18613,N_17387);
nor U23916 (N_23916,N_17459,N_16747);
nand U23917 (N_23917,N_15909,N_19827);
nor U23918 (N_23918,N_18876,N_19750);
or U23919 (N_23919,N_17766,N_15269);
nand U23920 (N_23920,N_18025,N_15327);
and U23921 (N_23921,N_18373,N_16247);
or U23922 (N_23922,N_16994,N_19721);
nand U23923 (N_23923,N_18922,N_15918);
nand U23924 (N_23924,N_15735,N_18502);
and U23925 (N_23925,N_18701,N_18067);
nor U23926 (N_23926,N_16667,N_18277);
nor U23927 (N_23927,N_15344,N_15238);
nand U23928 (N_23928,N_15211,N_15976);
nand U23929 (N_23929,N_16977,N_15380);
and U23930 (N_23930,N_19843,N_19402);
or U23931 (N_23931,N_16602,N_19848);
and U23932 (N_23932,N_18965,N_15907);
and U23933 (N_23933,N_16240,N_19011);
nor U23934 (N_23934,N_15781,N_15606);
and U23935 (N_23935,N_18999,N_18666);
nor U23936 (N_23936,N_18837,N_18158);
or U23937 (N_23937,N_17211,N_15189);
and U23938 (N_23938,N_17747,N_19882);
and U23939 (N_23939,N_17968,N_17054);
and U23940 (N_23940,N_19871,N_19177);
or U23941 (N_23941,N_16005,N_15689);
or U23942 (N_23942,N_15591,N_19688);
nor U23943 (N_23943,N_17246,N_16841);
and U23944 (N_23944,N_15178,N_19059);
and U23945 (N_23945,N_19654,N_19627);
and U23946 (N_23946,N_15324,N_19832);
and U23947 (N_23947,N_18880,N_16287);
or U23948 (N_23948,N_16366,N_19622);
nor U23949 (N_23949,N_18733,N_16156);
xnor U23950 (N_23950,N_18416,N_18912);
nor U23951 (N_23951,N_16257,N_18475);
xor U23952 (N_23952,N_18761,N_16384);
or U23953 (N_23953,N_18752,N_17253);
nor U23954 (N_23954,N_18370,N_16114);
or U23955 (N_23955,N_18237,N_17996);
nand U23956 (N_23956,N_16436,N_15933);
nor U23957 (N_23957,N_17183,N_15012);
nand U23958 (N_23958,N_18270,N_19638);
or U23959 (N_23959,N_18538,N_18746);
nor U23960 (N_23960,N_19045,N_18768);
xor U23961 (N_23961,N_19687,N_18080);
and U23962 (N_23962,N_19553,N_18814);
or U23963 (N_23963,N_17319,N_18671);
nor U23964 (N_23964,N_17602,N_17999);
and U23965 (N_23965,N_16159,N_19532);
nor U23966 (N_23966,N_19998,N_15416);
nor U23967 (N_23967,N_18305,N_16707);
and U23968 (N_23968,N_17357,N_18652);
nor U23969 (N_23969,N_15452,N_18640);
nand U23970 (N_23970,N_17079,N_19437);
nor U23971 (N_23971,N_18828,N_15087);
xnor U23972 (N_23972,N_15562,N_16703);
nand U23973 (N_23973,N_17923,N_17695);
nor U23974 (N_23974,N_16156,N_15869);
and U23975 (N_23975,N_16954,N_16865);
and U23976 (N_23976,N_19648,N_15930);
nand U23977 (N_23977,N_15273,N_19835);
nand U23978 (N_23978,N_19350,N_18803);
nand U23979 (N_23979,N_19835,N_15181);
nand U23980 (N_23980,N_19616,N_17629);
and U23981 (N_23981,N_18348,N_16134);
nor U23982 (N_23982,N_16737,N_15519);
or U23983 (N_23983,N_16700,N_18961);
nand U23984 (N_23984,N_17315,N_17952);
and U23985 (N_23985,N_19946,N_17250);
nor U23986 (N_23986,N_16858,N_18231);
xor U23987 (N_23987,N_15137,N_17778);
nand U23988 (N_23988,N_18188,N_15016);
nand U23989 (N_23989,N_16498,N_16817);
nand U23990 (N_23990,N_16704,N_17870);
or U23991 (N_23991,N_15150,N_15642);
nand U23992 (N_23992,N_15225,N_19153);
nor U23993 (N_23993,N_18548,N_18011);
and U23994 (N_23994,N_17709,N_15423);
nand U23995 (N_23995,N_17592,N_16267);
nand U23996 (N_23996,N_16519,N_18580);
nor U23997 (N_23997,N_17813,N_17498);
or U23998 (N_23998,N_15473,N_15537);
nand U23999 (N_23999,N_16045,N_16686);
or U24000 (N_24000,N_16883,N_15535);
or U24001 (N_24001,N_15463,N_15459);
nand U24002 (N_24002,N_17322,N_17033);
nor U24003 (N_24003,N_18052,N_19137);
and U24004 (N_24004,N_19216,N_17086);
nand U24005 (N_24005,N_18795,N_15603);
or U24006 (N_24006,N_18173,N_15062);
nand U24007 (N_24007,N_16903,N_19769);
nand U24008 (N_24008,N_19940,N_19998);
nor U24009 (N_24009,N_19924,N_18880);
nand U24010 (N_24010,N_16034,N_15467);
nand U24011 (N_24011,N_18207,N_17844);
nand U24012 (N_24012,N_18944,N_16795);
nor U24013 (N_24013,N_18574,N_17374);
and U24014 (N_24014,N_16374,N_15463);
and U24015 (N_24015,N_16430,N_18815);
nand U24016 (N_24016,N_19450,N_17060);
or U24017 (N_24017,N_16699,N_16165);
or U24018 (N_24018,N_16338,N_17300);
nor U24019 (N_24019,N_17291,N_19106);
and U24020 (N_24020,N_16362,N_17735);
xor U24021 (N_24021,N_16670,N_16113);
nor U24022 (N_24022,N_18910,N_15788);
nand U24023 (N_24023,N_17461,N_19084);
nand U24024 (N_24024,N_17807,N_15325);
nor U24025 (N_24025,N_19679,N_18897);
and U24026 (N_24026,N_18331,N_19958);
or U24027 (N_24027,N_17702,N_19012);
nor U24028 (N_24028,N_19088,N_18479);
nand U24029 (N_24029,N_17464,N_18858);
xor U24030 (N_24030,N_19456,N_18254);
or U24031 (N_24031,N_16574,N_19292);
nand U24032 (N_24032,N_18503,N_17345);
or U24033 (N_24033,N_16562,N_18210);
or U24034 (N_24034,N_17216,N_16889);
and U24035 (N_24035,N_19438,N_19107);
nand U24036 (N_24036,N_17990,N_17982);
and U24037 (N_24037,N_17217,N_16860);
or U24038 (N_24038,N_17683,N_15710);
or U24039 (N_24039,N_16151,N_16538);
nor U24040 (N_24040,N_16402,N_18011);
or U24041 (N_24041,N_17096,N_19770);
and U24042 (N_24042,N_19760,N_16176);
nand U24043 (N_24043,N_16721,N_16295);
nor U24044 (N_24044,N_18568,N_18854);
or U24045 (N_24045,N_15276,N_15135);
nand U24046 (N_24046,N_15134,N_16091);
and U24047 (N_24047,N_15970,N_16289);
nand U24048 (N_24048,N_18742,N_19280);
nor U24049 (N_24049,N_15456,N_16584);
nand U24050 (N_24050,N_16729,N_16768);
nand U24051 (N_24051,N_19116,N_17564);
or U24052 (N_24052,N_17289,N_16489);
nor U24053 (N_24053,N_16589,N_15711);
and U24054 (N_24054,N_17603,N_16668);
and U24055 (N_24055,N_19284,N_17241);
nor U24056 (N_24056,N_15861,N_19635);
or U24057 (N_24057,N_17155,N_18403);
nand U24058 (N_24058,N_17459,N_19491);
and U24059 (N_24059,N_17180,N_15006);
nand U24060 (N_24060,N_15306,N_16921);
and U24061 (N_24061,N_17579,N_19147);
nand U24062 (N_24062,N_17986,N_17190);
or U24063 (N_24063,N_17278,N_16522);
and U24064 (N_24064,N_15389,N_16375);
nand U24065 (N_24065,N_15733,N_16026);
or U24066 (N_24066,N_18562,N_17974);
and U24067 (N_24067,N_18920,N_17800);
and U24068 (N_24068,N_18292,N_15753);
nand U24069 (N_24069,N_16155,N_19673);
nand U24070 (N_24070,N_16588,N_17403);
nand U24071 (N_24071,N_15591,N_17363);
or U24072 (N_24072,N_16588,N_15458);
or U24073 (N_24073,N_18518,N_19028);
and U24074 (N_24074,N_15165,N_19532);
nor U24075 (N_24075,N_19823,N_16060);
nor U24076 (N_24076,N_18693,N_15329);
or U24077 (N_24077,N_16720,N_15463);
and U24078 (N_24078,N_17038,N_17697);
nor U24079 (N_24079,N_19338,N_18665);
nor U24080 (N_24080,N_15102,N_17895);
or U24081 (N_24081,N_17069,N_18562);
nor U24082 (N_24082,N_15590,N_16903);
nand U24083 (N_24083,N_15869,N_17230);
and U24084 (N_24084,N_19674,N_18286);
and U24085 (N_24085,N_19180,N_17784);
nand U24086 (N_24086,N_16109,N_15155);
nand U24087 (N_24087,N_16712,N_16161);
nand U24088 (N_24088,N_16752,N_15693);
nand U24089 (N_24089,N_17296,N_19040);
nand U24090 (N_24090,N_15546,N_19487);
nand U24091 (N_24091,N_16149,N_15893);
or U24092 (N_24092,N_16670,N_19450);
nand U24093 (N_24093,N_15848,N_15738);
nand U24094 (N_24094,N_15205,N_17883);
nand U24095 (N_24095,N_19958,N_17282);
nand U24096 (N_24096,N_17506,N_17122);
and U24097 (N_24097,N_17271,N_15355);
and U24098 (N_24098,N_17941,N_16039);
or U24099 (N_24099,N_19139,N_17754);
nor U24100 (N_24100,N_19653,N_15413);
nand U24101 (N_24101,N_16018,N_16495);
nor U24102 (N_24102,N_18707,N_17156);
and U24103 (N_24103,N_15355,N_19989);
or U24104 (N_24104,N_17654,N_16459);
nor U24105 (N_24105,N_18038,N_16252);
nand U24106 (N_24106,N_18527,N_16182);
nor U24107 (N_24107,N_16381,N_16664);
nand U24108 (N_24108,N_16339,N_15934);
or U24109 (N_24109,N_18959,N_16192);
nand U24110 (N_24110,N_16016,N_18378);
and U24111 (N_24111,N_16826,N_17710);
or U24112 (N_24112,N_15222,N_19954);
xor U24113 (N_24113,N_18468,N_16853);
nand U24114 (N_24114,N_19545,N_16610);
nand U24115 (N_24115,N_16059,N_18236);
and U24116 (N_24116,N_15171,N_18234);
nand U24117 (N_24117,N_19687,N_18671);
or U24118 (N_24118,N_17190,N_16421);
and U24119 (N_24119,N_16113,N_16249);
nor U24120 (N_24120,N_19509,N_16812);
or U24121 (N_24121,N_15713,N_17885);
or U24122 (N_24122,N_18538,N_18416);
nand U24123 (N_24123,N_17313,N_16607);
nand U24124 (N_24124,N_16795,N_16444);
and U24125 (N_24125,N_16357,N_18894);
or U24126 (N_24126,N_18591,N_15704);
and U24127 (N_24127,N_15709,N_18110);
nand U24128 (N_24128,N_18116,N_18552);
or U24129 (N_24129,N_18901,N_15464);
and U24130 (N_24130,N_15328,N_15182);
nand U24131 (N_24131,N_18469,N_16325);
nand U24132 (N_24132,N_16120,N_17799);
and U24133 (N_24133,N_15855,N_18762);
or U24134 (N_24134,N_19047,N_16568);
nor U24135 (N_24135,N_16705,N_19758);
nand U24136 (N_24136,N_15837,N_17943);
nor U24137 (N_24137,N_19726,N_17056);
or U24138 (N_24138,N_16506,N_16326);
or U24139 (N_24139,N_15859,N_15584);
nor U24140 (N_24140,N_16950,N_18965);
or U24141 (N_24141,N_16980,N_19662);
nand U24142 (N_24142,N_17525,N_18374);
nor U24143 (N_24143,N_15672,N_19075);
nand U24144 (N_24144,N_18567,N_15153);
nor U24145 (N_24145,N_17482,N_17314);
or U24146 (N_24146,N_15701,N_16564);
and U24147 (N_24147,N_16901,N_19999);
nor U24148 (N_24148,N_19549,N_18857);
and U24149 (N_24149,N_17244,N_18120);
nand U24150 (N_24150,N_18769,N_18850);
or U24151 (N_24151,N_17831,N_17047);
and U24152 (N_24152,N_17818,N_18265);
or U24153 (N_24153,N_19067,N_16415);
or U24154 (N_24154,N_15616,N_18846);
nand U24155 (N_24155,N_16192,N_18921);
and U24156 (N_24156,N_17669,N_16713);
and U24157 (N_24157,N_15220,N_16410);
or U24158 (N_24158,N_17278,N_17161);
or U24159 (N_24159,N_19196,N_16644);
nor U24160 (N_24160,N_15085,N_18002);
nor U24161 (N_24161,N_19868,N_17537);
nand U24162 (N_24162,N_17520,N_19576);
or U24163 (N_24163,N_16500,N_15366);
and U24164 (N_24164,N_16474,N_15943);
xor U24165 (N_24165,N_16867,N_19587);
nand U24166 (N_24166,N_17565,N_15807);
or U24167 (N_24167,N_15913,N_19838);
nor U24168 (N_24168,N_16515,N_15969);
nor U24169 (N_24169,N_15282,N_16260);
nand U24170 (N_24170,N_18974,N_18615);
or U24171 (N_24171,N_16943,N_19059);
or U24172 (N_24172,N_17367,N_19466);
nand U24173 (N_24173,N_18021,N_19049);
and U24174 (N_24174,N_19361,N_18968);
and U24175 (N_24175,N_18956,N_15449);
and U24176 (N_24176,N_15031,N_16588);
nor U24177 (N_24177,N_18218,N_17691);
or U24178 (N_24178,N_19817,N_17854);
and U24179 (N_24179,N_18933,N_17078);
or U24180 (N_24180,N_19819,N_16684);
and U24181 (N_24181,N_18370,N_15879);
or U24182 (N_24182,N_16465,N_15450);
or U24183 (N_24183,N_15585,N_15251);
or U24184 (N_24184,N_19179,N_18114);
nor U24185 (N_24185,N_17473,N_15471);
or U24186 (N_24186,N_19173,N_17152);
nand U24187 (N_24187,N_15823,N_17991);
or U24188 (N_24188,N_19921,N_18667);
nor U24189 (N_24189,N_18301,N_16965);
nor U24190 (N_24190,N_18537,N_16941);
or U24191 (N_24191,N_17895,N_17492);
nand U24192 (N_24192,N_15161,N_18353);
nand U24193 (N_24193,N_15502,N_18656);
or U24194 (N_24194,N_16276,N_19640);
nand U24195 (N_24195,N_18449,N_16536);
nor U24196 (N_24196,N_18180,N_19569);
nor U24197 (N_24197,N_16130,N_15658);
nor U24198 (N_24198,N_17949,N_18417);
and U24199 (N_24199,N_17860,N_16986);
nand U24200 (N_24200,N_19253,N_15539);
and U24201 (N_24201,N_19945,N_16918);
nand U24202 (N_24202,N_16557,N_17951);
and U24203 (N_24203,N_19038,N_18897);
and U24204 (N_24204,N_16278,N_18421);
or U24205 (N_24205,N_19867,N_16420);
or U24206 (N_24206,N_17929,N_16790);
and U24207 (N_24207,N_17458,N_18299);
or U24208 (N_24208,N_18018,N_18823);
and U24209 (N_24209,N_17758,N_17533);
or U24210 (N_24210,N_15617,N_16767);
and U24211 (N_24211,N_19519,N_17915);
nor U24212 (N_24212,N_18719,N_15236);
nand U24213 (N_24213,N_17868,N_16699);
nand U24214 (N_24214,N_18257,N_19876);
nand U24215 (N_24215,N_19342,N_16254);
and U24216 (N_24216,N_19076,N_17901);
nand U24217 (N_24217,N_16471,N_17788);
nor U24218 (N_24218,N_18814,N_17113);
nand U24219 (N_24219,N_15746,N_19970);
and U24220 (N_24220,N_15949,N_19929);
nand U24221 (N_24221,N_17843,N_18076);
or U24222 (N_24222,N_17925,N_18126);
or U24223 (N_24223,N_17866,N_17329);
or U24224 (N_24224,N_16667,N_16677);
and U24225 (N_24225,N_17417,N_15208);
nand U24226 (N_24226,N_15209,N_17369);
and U24227 (N_24227,N_19320,N_19014);
and U24228 (N_24228,N_19043,N_16781);
and U24229 (N_24229,N_19637,N_16041);
nand U24230 (N_24230,N_16121,N_18361);
or U24231 (N_24231,N_17180,N_16900);
nor U24232 (N_24232,N_15737,N_18908);
or U24233 (N_24233,N_15131,N_19229);
and U24234 (N_24234,N_15378,N_18382);
nand U24235 (N_24235,N_19235,N_15448);
nor U24236 (N_24236,N_18673,N_15596);
nand U24237 (N_24237,N_19497,N_15171);
and U24238 (N_24238,N_15404,N_17478);
nand U24239 (N_24239,N_17981,N_19886);
and U24240 (N_24240,N_17618,N_18221);
nand U24241 (N_24241,N_19954,N_15364);
and U24242 (N_24242,N_15226,N_19690);
or U24243 (N_24243,N_19272,N_19960);
nand U24244 (N_24244,N_18669,N_18340);
nand U24245 (N_24245,N_15224,N_18982);
xor U24246 (N_24246,N_16353,N_17467);
or U24247 (N_24247,N_15523,N_17726);
and U24248 (N_24248,N_18408,N_18265);
or U24249 (N_24249,N_17729,N_15218);
and U24250 (N_24250,N_18290,N_18711);
nor U24251 (N_24251,N_19969,N_15532);
and U24252 (N_24252,N_18924,N_17062);
nand U24253 (N_24253,N_19444,N_17440);
nand U24254 (N_24254,N_15061,N_16186);
nand U24255 (N_24255,N_17561,N_19612);
and U24256 (N_24256,N_18454,N_17820);
nand U24257 (N_24257,N_16949,N_17750);
xnor U24258 (N_24258,N_15496,N_18431);
nand U24259 (N_24259,N_19398,N_17866);
and U24260 (N_24260,N_19018,N_16267);
or U24261 (N_24261,N_17652,N_15196);
nor U24262 (N_24262,N_16289,N_19999);
nand U24263 (N_24263,N_19958,N_15930);
nand U24264 (N_24264,N_15508,N_17225);
nand U24265 (N_24265,N_16184,N_17887);
nand U24266 (N_24266,N_16016,N_19021);
or U24267 (N_24267,N_18708,N_18035);
nor U24268 (N_24268,N_15761,N_15126);
nand U24269 (N_24269,N_15225,N_17210);
nor U24270 (N_24270,N_15797,N_18242);
nor U24271 (N_24271,N_15351,N_17780);
nand U24272 (N_24272,N_16879,N_18288);
nand U24273 (N_24273,N_17597,N_19459);
nand U24274 (N_24274,N_16387,N_18189);
or U24275 (N_24275,N_15925,N_17689);
nor U24276 (N_24276,N_17957,N_17543);
and U24277 (N_24277,N_18458,N_17890);
nor U24278 (N_24278,N_18896,N_18987);
and U24279 (N_24279,N_15051,N_15461);
nor U24280 (N_24280,N_16494,N_18951);
nor U24281 (N_24281,N_19697,N_18311);
or U24282 (N_24282,N_18569,N_19572);
nand U24283 (N_24283,N_19436,N_15741);
nor U24284 (N_24284,N_16524,N_16920);
and U24285 (N_24285,N_18041,N_19262);
nand U24286 (N_24286,N_15585,N_15311);
or U24287 (N_24287,N_18530,N_19834);
and U24288 (N_24288,N_17487,N_19076);
nand U24289 (N_24289,N_19265,N_17344);
and U24290 (N_24290,N_15212,N_16211);
nor U24291 (N_24291,N_18913,N_16998);
nor U24292 (N_24292,N_16885,N_18639);
nor U24293 (N_24293,N_18247,N_19243);
nor U24294 (N_24294,N_17659,N_15958);
or U24295 (N_24295,N_16741,N_17183);
or U24296 (N_24296,N_18827,N_19895);
nor U24297 (N_24297,N_18902,N_16336);
nand U24298 (N_24298,N_18317,N_16408);
or U24299 (N_24299,N_15534,N_19896);
or U24300 (N_24300,N_18417,N_19301);
or U24301 (N_24301,N_15745,N_18265);
nor U24302 (N_24302,N_17568,N_15811);
or U24303 (N_24303,N_15646,N_18120);
nand U24304 (N_24304,N_16456,N_15942);
nand U24305 (N_24305,N_17773,N_16479);
and U24306 (N_24306,N_15906,N_17883);
nor U24307 (N_24307,N_17607,N_19500);
nand U24308 (N_24308,N_16906,N_15850);
nand U24309 (N_24309,N_19780,N_19124);
or U24310 (N_24310,N_18901,N_15531);
or U24311 (N_24311,N_17021,N_19873);
and U24312 (N_24312,N_17581,N_16076);
or U24313 (N_24313,N_19818,N_17984);
nand U24314 (N_24314,N_15248,N_15044);
nor U24315 (N_24315,N_19541,N_16265);
nor U24316 (N_24316,N_18437,N_17659);
nor U24317 (N_24317,N_19448,N_19222);
or U24318 (N_24318,N_16490,N_19766);
nor U24319 (N_24319,N_16630,N_15435);
nor U24320 (N_24320,N_17667,N_15557);
or U24321 (N_24321,N_16204,N_18334);
nor U24322 (N_24322,N_19999,N_16922);
and U24323 (N_24323,N_18820,N_17428);
or U24324 (N_24324,N_16831,N_17335);
and U24325 (N_24325,N_17561,N_17813);
nand U24326 (N_24326,N_19638,N_17493);
and U24327 (N_24327,N_16764,N_16405);
nor U24328 (N_24328,N_15930,N_17204);
or U24329 (N_24329,N_18791,N_18067);
nand U24330 (N_24330,N_16237,N_18320);
and U24331 (N_24331,N_16377,N_18464);
nand U24332 (N_24332,N_17246,N_19129);
and U24333 (N_24333,N_19728,N_19455);
nor U24334 (N_24334,N_17331,N_16779);
nand U24335 (N_24335,N_19311,N_15085);
and U24336 (N_24336,N_15094,N_16625);
or U24337 (N_24337,N_17900,N_18774);
and U24338 (N_24338,N_15241,N_18081);
nand U24339 (N_24339,N_15189,N_17589);
nand U24340 (N_24340,N_15782,N_15656);
and U24341 (N_24341,N_16061,N_18516);
nor U24342 (N_24342,N_18844,N_16785);
or U24343 (N_24343,N_15046,N_19745);
nand U24344 (N_24344,N_19786,N_17609);
nand U24345 (N_24345,N_16560,N_16489);
nand U24346 (N_24346,N_19094,N_19462);
or U24347 (N_24347,N_18544,N_15457);
and U24348 (N_24348,N_16397,N_15953);
and U24349 (N_24349,N_18763,N_19960);
nand U24350 (N_24350,N_18819,N_16761);
nand U24351 (N_24351,N_16015,N_17025);
nand U24352 (N_24352,N_17039,N_16549);
or U24353 (N_24353,N_18090,N_19177);
nand U24354 (N_24354,N_16339,N_19953);
or U24355 (N_24355,N_19776,N_17905);
or U24356 (N_24356,N_18048,N_18645);
nor U24357 (N_24357,N_18422,N_17838);
and U24358 (N_24358,N_16132,N_15725);
or U24359 (N_24359,N_17998,N_18000);
or U24360 (N_24360,N_16484,N_16091);
or U24361 (N_24361,N_16080,N_17144);
nand U24362 (N_24362,N_19914,N_16654);
and U24363 (N_24363,N_19100,N_18618);
xnor U24364 (N_24364,N_19631,N_16884);
or U24365 (N_24365,N_19863,N_18045);
nor U24366 (N_24366,N_17922,N_16989);
nand U24367 (N_24367,N_16380,N_16524);
nor U24368 (N_24368,N_19201,N_17175);
and U24369 (N_24369,N_16696,N_18479);
nand U24370 (N_24370,N_17951,N_17576);
nand U24371 (N_24371,N_17197,N_18254);
nand U24372 (N_24372,N_15981,N_16008);
nor U24373 (N_24373,N_18293,N_15812);
and U24374 (N_24374,N_18170,N_18028);
and U24375 (N_24375,N_15168,N_19442);
nand U24376 (N_24376,N_15645,N_16497);
nor U24377 (N_24377,N_18281,N_16351);
nand U24378 (N_24378,N_17914,N_17519);
nor U24379 (N_24379,N_16686,N_19131);
nor U24380 (N_24380,N_15015,N_15476);
nand U24381 (N_24381,N_19955,N_16143);
or U24382 (N_24382,N_15183,N_16467);
and U24383 (N_24383,N_15668,N_16420);
or U24384 (N_24384,N_16958,N_15226);
or U24385 (N_24385,N_15277,N_15702);
nor U24386 (N_24386,N_18977,N_15948);
or U24387 (N_24387,N_16101,N_15832);
and U24388 (N_24388,N_18577,N_16027);
or U24389 (N_24389,N_17126,N_17148);
nor U24390 (N_24390,N_16147,N_16135);
and U24391 (N_24391,N_15650,N_16678);
nor U24392 (N_24392,N_15476,N_15884);
and U24393 (N_24393,N_17604,N_15141);
or U24394 (N_24394,N_15346,N_15148);
or U24395 (N_24395,N_19320,N_19451);
and U24396 (N_24396,N_18618,N_17236);
or U24397 (N_24397,N_16952,N_19636);
and U24398 (N_24398,N_17696,N_18828);
or U24399 (N_24399,N_17332,N_18908);
nand U24400 (N_24400,N_17525,N_18471);
nor U24401 (N_24401,N_15929,N_17172);
nor U24402 (N_24402,N_18629,N_18498);
nand U24403 (N_24403,N_15637,N_19507);
or U24404 (N_24404,N_18178,N_18419);
or U24405 (N_24405,N_15529,N_17774);
nor U24406 (N_24406,N_19470,N_19473);
and U24407 (N_24407,N_19863,N_18141);
xor U24408 (N_24408,N_19675,N_17637);
nand U24409 (N_24409,N_18400,N_19361);
nor U24410 (N_24410,N_16337,N_15841);
and U24411 (N_24411,N_16376,N_15352);
or U24412 (N_24412,N_18154,N_16348);
or U24413 (N_24413,N_19071,N_15796);
nand U24414 (N_24414,N_19137,N_17663);
nor U24415 (N_24415,N_16561,N_16896);
and U24416 (N_24416,N_16491,N_16558);
and U24417 (N_24417,N_19329,N_16651);
nand U24418 (N_24418,N_19226,N_16691);
nor U24419 (N_24419,N_19196,N_16269);
and U24420 (N_24420,N_16662,N_19516);
xnor U24421 (N_24421,N_17487,N_17471);
or U24422 (N_24422,N_18479,N_16992);
nor U24423 (N_24423,N_19927,N_17824);
or U24424 (N_24424,N_15493,N_16081);
nand U24425 (N_24425,N_18529,N_19430);
nand U24426 (N_24426,N_15535,N_16923);
or U24427 (N_24427,N_15564,N_16926);
nand U24428 (N_24428,N_18190,N_15661);
nor U24429 (N_24429,N_18633,N_16671);
or U24430 (N_24430,N_18536,N_18764);
nand U24431 (N_24431,N_18079,N_15641);
nand U24432 (N_24432,N_16280,N_16074);
nand U24433 (N_24433,N_16742,N_16777);
or U24434 (N_24434,N_15781,N_19684);
nor U24435 (N_24435,N_15437,N_16218);
and U24436 (N_24436,N_15201,N_17909);
nand U24437 (N_24437,N_15711,N_15612);
nand U24438 (N_24438,N_17539,N_16757);
and U24439 (N_24439,N_16377,N_16757);
or U24440 (N_24440,N_18838,N_18532);
and U24441 (N_24441,N_16266,N_19643);
and U24442 (N_24442,N_19146,N_17240);
nor U24443 (N_24443,N_18719,N_17699);
or U24444 (N_24444,N_16480,N_16623);
nor U24445 (N_24445,N_18530,N_19482);
nor U24446 (N_24446,N_15639,N_17926);
or U24447 (N_24447,N_17962,N_15858);
and U24448 (N_24448,N_17384,N_17151);
or U24449 (N_24449,N_18243,N_16861);
or U24450 (N_24450,N_16081,N_16506);
or U24451 (N_24451,N_17619,N_15484);
and U24452 (N_24452,N_18684,N_17038);
nor U24453 (N_24453,N_18834,N_15230);
nor U24454 (N_24454,N_17452,N_17654);
or U24455 (N_24455,N_15005,N_15947);
and U24456 (N_24456,N_17192,N_17424);
or U24457 (N_24457,N_18785,N_17975);
nand U24458 (N_24458,N_17298,N_17978);
nor U24459 (N_24459,N_19668,N_17143);
nor U24460 (N_24460,N_18826,N_16014);
and U24461 (N_24461,N_19243,N_19594);
or U24462 (N_24462,N_18091,N_17449);
xnor U24463 (N_24463,N_16908,N_16681);
nand U24464 (N_24464,N_15632,N_15143);
nand U24465 (N_24465,N_15896,N_17126);
and U24466 (N_24466,N_16781,N_19607);
nand U24467 (N_24467,N_17445,N_18867);
or U24468 (N_24468,N_15296,N_17460);
or U24469 (N_24469,N_18532,N_17363);
and U24470 (N_24470,N_17864,N_19128);
and U24471 (N_24471,N_18718,N_15783);
nor U24472 (N_24472,N_19000,N_18118);
or U24473 (N_24473,N_16187,N_15517);
nor U24474 (N_24474,N_17297,N_18784);
nor U24475 (N_24475,N_17538,N_19082);
nand U24476 (N_24476,N_16349,N_17638);
nand U24477 (N_24477,N_18026,N_19873);
and U24478 (N_24478,N_15307,N_15159);
nor U24479 (N_24479,N_17180,N_15871);
or U24480 (N_24480,N_19550,N_16588);
nor U24481 (N_24481,N_17606,N_16530);
nor U24482 (N_24482,N_19104,N_16140);
or U24483 (N_24483,N_18824,N_15876);
and U24484 (N_24484,N_19878,N_18135);
nand U24485 (N_24485,N_19922,N_16310);
nand U24486 (N_24486,N_19150,N_18230);
or U24487 (N_24487,N_18712,N_17582);
nand U24488 (N_24488,N_19869,N_15987);
nor U24489 (N_24489,N_19589,N_15612);
nor U24490 (N_24490,N_17033,N_15835);
nor U24491 (N_24491,N_19293,N_16854);
and U24492 (N_24492,N_18100,N_17910);
nand U24493 (N_24493,N_16736,N_16920);
and U24494 (N_24494,N_15483,N_16656);
or U24495 (N_24495,N_19611,N_18168);
or U24496 (N_24496,N_15867,N_16036);
xnor U24497 (N_24497,N_17997,N_19577);
nor U24498 (N_24498,N_15690,N_16320);
and U24499 (N_24499,N_15980,N_17503);
nand U24500 (N_24500,N_18668,N_19853);
and U24501 (N_24501,N_19565,N_15908);
nand U24502 (N_24502,N_15634,N_18698);
or U24503 (N_24503,N_15076,N_18753);
or U24504 (N_24504,N_18597,N_15688);
and U24505 (N_24505,N_17109,N_17712);
nand U24506 (N_24506,N_18182,N_16963);
or U24507 (N_24507,N_18099,N_18173);
nor U24508 (N_24508,N_16065,N_19409);
and U24509 (N_24509,N_18985,N_17725);
nand U24510 (N_24510,N_18895,N_18150);
nand U24511 (N_24511,N_15451,N_17471);
nand U24512 (N_24512,N_16757,N_19806);
nor U24513 (N_24513,N_17284,N_18618);
or U24514 (N_24514,N_15904,N_17199);
or U24515 (N_24515,N_17672,N_16132);
and U24516 (N_24516,N_19435,N_17589);
nor U24517 (N_24517,N_15494,N_18919);
or U24518 (N_24518,N_18518,N_19113);
nand U24519 (N_24519,N_19682,N_19550);
or U24520 (N_24520,N_18977,N_16509);
or U24521 (N_24521,N_17183,N_19361);
nor U24522 (N_24522,N_19003,N_19859);
nor U24523 (N_24523,N_17870,N_15666);
or U24524 (N_24524,N_15792,N_17257);
and U24525 (N_24525,N_15979,N_17206);
xor U24526 (N_24526,N_17034,N_16344);
nand U24527 (N_24527,N_18192,N_18542);
or U24528 (N_24528,N_15239,N_17474);
nand U24529 (N_24529,N_19905,N_18243);
nand U24530 (N_24530,N_16584,N_16493);
nand U24531 (N_24531,N_17304,N_15102);
and U24532 (N_24532,N_16702,N_15668);
or U24533 (N_24533,N_18820,N_16744);
or U24534 (N_24534,N_18715,N_17094);
nand U24535 (N_24535,N_15765,N_16234);
nand U24536 (N_24536,N_15019,N_18269);
nor U24537 (N_24537,N_17527,N_17221);
nor U24538 (N_24538,N_19425,N_19956);
nor U24539 (N_24539,N_17664,N_15813);
nand U24540 (N_24540,N_19892,N_18058);
or U24541 (N_24541,N_17938,N_15617);
nand U24542 (N_24542,N_19494,N_18128);
or U24543 (N_24543,N_17995,N_15511);
nand U24544 (N_24544,N_15781,N_15681);
nor U24545 (N_24545,N_19499,N_17683);
nor U24546 (N_24546,N_17958,N_15282);
nand U24547 (N_24547,N_15242,N_18194);
nor U24548 (N_24548,N_16752,N_19725);
nor U24549 (N_24549,N_18864,N_18414);
xor U24550 (N_24550,N_15115,N_18915);
nor U24551 (N_24551,N_17185,N_15892);
nor U24552 (N_24552,N_19811,N_19990);
nand U24553 (N_24553,N_17106,N_16037);
and U24554 (N_24554,N_18362,N_15264);
and U24555 (N_24555,N_15626,N_16963);
nor U24556 (N_24556,N_17465,N_19993);
or U24557 (N_24557,N_19867,N_17068);
and U24558 (N_24558,N_19100,N_18145);
or U24559 (N_24559,N_16667,N_17446);
nor U24560 (N_24560,N_15342,N_19535);
xnor U24561 (N_24561,N_17587,N_17974);
nand U24562 (N_24562,N_15027,N_17369);
or U24563 (N_24563,N_15791,N_15508);
and U24564 (N_24564,N_18484,N_17379);
or U24565 (N_24565,N_17984,N_16490);
and U24566 (N_24566,N_18701,N_18828);
or U24567 (N_24567,N_17035,N_15206);
nand U24568 (N_24568,N_19598,N_15838);
nor U24569 (N_24569,N_18447,N_19701);
nand U24570 (N_24570,N_18387,N_18909);
or U24571 (N_24571,N_16827,N_19228);
xnor U24572 (N_24572,N_17433,N_17113);
or U24573 (N_24573,N_15951,N_18326);
nand U24574 (N_24574,N_18733,N_19827);
or U24575 (N_24575,N_16952,N_15620);
nand U24576 (N_24576,N_15211,N_18768);
xnor U24577 (N_24577,N_17656,N_16207);
and U24578 (N_24578,N_15506,N_18319);
xnor U24579 (N_24579,N_15034,N_18537);
or U24580 (N_24580,N_19244,N_19824);
nand U24581 (N_24581,N_17016,N_15765);
and U24582 (N_24582,N_19127,N_19919);
and U24583 (N_24583,N_18844,N_15985);
nand U24584 (N_24584,N_18878,N_19360);
nor U24585 (N_24585,N_15772,N_19184);
and U24586 (N_24586,N_18696,N_18353);
and U24587 (N_24587,N_19887,N_18813);
nand U24588 (N_24588,N_19032,N_19564);
or U24589 (N_24589,N_18453,N_15665);
nor U24590 (N_24590,N_18367,N_19222);
nand U24591 (N_24591,N_16441,N_16366);
nor U24592 (N_24592,N_15351,N_16769);
or U24593 (N_24593,N_15598,N_16342);
or U24594 (N_24594,N_15178,N_17945);
and U24595 (N_24595,N_19250,N_18700);
and U24596 (N_24596,N_16547,N_17246);
nor U24597 (N_24597,N_19857,N_17120);
nand U24598 (N_24598,N_15659,N_17451);
xor U24599 (N_24599,N_16077,N_19163);
nor U24600 (N_24600,N_18117,N_17418);
or U24601 (N_24601,N_15677,N_15141);
xnor U24602 (N_24602,N_18345,N_17181);
or U24603 (N_24603,N_18464,N_19815);
or U24604 (N_24604,N_16042,N_19649);
nand U24605 (N_24605,N_16230,N_19473);
nor U24606 (N_24606,N_16348,N_19388);
and U24607 (N_24607,N_18723,N_16986);
or U24608 (N_24608,N_15198,N_17664);
xor U24609 (N_24609,N_19885,N_15154);
nor U24610 (N_24610,N_16447,N_17566);
xnor U24611 (N_24611,N_18909,N_19259);
nand U24612 (N_24612,N_16867,N_16316);
nand U24613 (N_24613,N_18470,N_15037);
and U24614 (N_24614,N_15302,N_15434);
nand U24615 (N_24615,N_17993,N_15223);
nand U24616 (N_24616,N_19758,N_19805);
nor U24617 (N_24617,N_15581,N_19283);
nand U24618 (N_24618,N_18262,N_18365);
nor U24619 (N_24619,N_18873,N_19282);
or U24620 (N_24620,N_18962,N_18624);
and U24621 (N_24621,N_16424,N_16151);
and U24622 (N_24622,N_19944,N_15268);
nand U24623 (N_24623,N_15610,N_16826);
and U24624 (N_24624,N_15593,N_16476);
xnor U24625 (N_24625,N_18423,N_18054);
or U24626 (N_24626,N_19785,N_19051);
or U24627 (N_24627,N_18159,N_16997);
nand U24628 (N_24628,N_18555,N_17388);
nor U24629 (N_24629,N_18774,N_15078);
xnor U24630 (N_24630,N_16707,N_17220);
nor U24631 (N_24631,N_17769,N_18543);
nand U24632 (N_24632,N_19457,N_17830);
nand U24633 (N_24633,N_15613,N_19770);
nand U24634 (N_24634,N_17595,N_18165);
and U24635 (N_24635,N_16956,N_19558);
and U24636 (N_24636,N_18823,N_19811);
nand U24637 (N_24637,N_16061,N_16323);
nand U24638 (N_24638,N_16880,N_16413);
nand U24639 (N_24639,N_19575,N_17561);
or U24640 (N_24640,N_19349,N_18005);
or U24641 (N_24641,N_18743,N_18553);
xor U24642 (N_24642,N_16135,N_15976);
nor U24643 (N_24643,N_15589,N_18508);
and U24644 (N_24644,N_15013,N_19585);
nand U24645 (N_24645,N_17328,N_19141);
or U24646 (N_24646,N_15920,N_15995);
or U24647 (N_24647,N_16000,N_18249);
or U24648 (N_24648,N_16358,N_16928);
and U24649 (N_24649,N_16255,N_17658);
nor U24650 (N_24650,N_15228,N_19062);
and U24651 (N_24651,N_15418,N_17430);
xnor U24652 (N_24652,N_16813,N_19567);
and U24653 (N_24653,N_17310,N_19338);
and U24654 (N_24654,N_16961,N_17761);
and U24655 (N_24655,N_16146,N_19393);
or U24656 (N_24656,N_16616,N_16710);
nor U24657 (N_24657,N_17014,N_16745);
nor U24658 (N_24658,N_17140,N_15459);
nor U24659 (N_24659,N_15200,N_18052);
or U24660 (N_24660,N_19859,N_19279);
and U24661 (N_24661,N_17139,N_16785);
nor U24662 (N_24662,N_15003,N_16164);
nand U24663 (N_24663,N_17089,N_15156);
or U24664 (N_24664,N_18305,N_16015);
nand U24665 (N_24665,N_18587,N_19627);
nor U24666 (N_24666,N_19001,N_19035);
or U24667 (N_24667,N_17731,N_19043);
nor U24668 (N_24668,N_15007,N_15575);
nand U24669 (N_24669,N_19664,N_19361);
and U24670 (N_24670,N_16200,N_18569);
nor U24671 (N_24671,N_19491,N_19323);
or U24672 (N_24672,N_15468,N_17231);
or U24673 (N_24673,N_17941,N_19255);
or U24674 (N_24674,N_15929,N_17963);
nand U24675 (N_24675,N_15999,N_19903);
and U24676 (N_24676,N_18905,N_15656);
and U24677 (N_24677,N_19105,N_15364);
nor U24678 (N_24678,N_18492,N_16600);
nand U24679 (N_24679,N_16470,N_16545);
nor U24680 (N_24680,N_17368,N_17554);
nand U24681 (N_24681,N_18747,N_17108);
and U24682 (N_24682,N_15031,N_17420);
or U24683 (N_24683,N_19792,N_18688);
or U24684 (N_24684,N_16282,N_15944);
or U24685 (N_24685,N_15580,N_18115);
nand U24686 (N_24686,N_17526,N_18849);
and U24687 (N_24687,N_16143,N_18114);
nand U24688 (N_24688,N_18132,N_19948);
or U24689 (N_24689,N_17967,N_18260);
nand U24690 (N_24690,N_15522,N_15714);
and U24691 (N_24691,N_16015,N_16861);
nor U24692 (N_24692,N_19380,N_17823);
and U24693 (N_24693,N_18188,N_19925);
or U24694 (N_24694,N_18732,N_19733);
nor U24695 (N_24695,N_19342,N_15368);
nor U24696 (N_24696,N_17601,N_16374);
or U24697 (N_24697,N_18023,N_17351);
nor U24698 (N_24698,N_18912,N_15304);
nor U24699 (N_24699,N_19550,N_15177);
nor U24700 (N_24700,N_17461,N_15594);
or U24701 (N_24701,N_18180,N_17509);
and U24702 (N_24702,N_18891,N_19316);
and U24703 (N_24703,N_17127,N_17485);
and U24704 (N_24704,N_16142,N_16104);
nor U24705 (N_24705,N_16666,N_15499);
or U24706 (N_24706,N_15076,N_16707);
nand U24707 (N_24707,N_17661,N_19127);
nor U24708 (N_24708,N_18143,N_19842);
nor U24709 (N_24709,N_16518,N_15509);
and U24710 (N_24710,N_15577,N_17751);
or U24711 (N_24711,N_15636,N_15624);
or U24712 (N_24712,N_19885,N_19835);
nor U24713 (N_24713,N_16923,N_17342);
nor U24714 (N_24714,N_17861,N_15880);
or U24715 (N_24715,N_19273,N_15618);
and U24716 (N_24716,N_17375,N_18569);
or U24717 (N_24717,N_15487,N_18270);
or U24718 (N_24718,N_16930,N_15126);
nand U24719 (N_24719,N_16500,N_19318);
and U24720 (N_24720,N_16349,N_19889);
or U24721 (N_24721,N_17117,N_15183);
nor U24722 (N_24722,N_19367,N_15314);
or U24723 (N_24723,N_17293,N_18764);
xor U24724 (N_24724,N_17307,N_19733);
or U24725 (N_24725,N_15865,N_16497);
or U24726 (N_24726,N_17182,N_18721);
nor U24727 (N_24727,N_18574,N_17647);
or U24728 (N_24728,N_19055,N_16979);
nand U24729 (N_24729,N_18712,N_16065);
or U24730 (N_24730,N_16121,N_16518);
nand U24731 (N_24731,N_17058,N_19947);
or U24732 (N_24732,N_18665,N_16908);
nand U24733 (N_24733,N_19918,N_18814);
xnor U24734 (N_24734,N_16448,N_19832);
nand U24735 (N_24735,N_16794,N_16126);
and U24736 (N_24736,N_15988,N_16741);
nor U24737 (N_24737,N_17213,N_18547);
or U24738 (N_24738,N_17607,N_17265);
nand U24739 (N_24739,N_16654,N_19310);
or U24740 (N_24740,N_16593,N_16830);
nand U24741 (N_24741,N_15389,N_18076);
nor U24742 (N_24742,N_18563,N_19007);
nand U24743 (N_24743,N_17033,N_15136);
xor U24744 (N_24744,N_19174,N_17350);
nand U24745 (N_24745,N_16474,N_15576);
and U24746 (N_24746,N_18679,N_19563);
nor U24747 (N_24747,N_19912,N_16932);
or U24748 (N_24748,N_16904,N_16705);
or U24749 (N_24749,N_15167,N_15927);
and U24750 (N_24750,N_19953,N_19590);
or U24751 (N_24751,N_15397,N_15882);
nor U24752 (N_24752,N_17076,N_18367);
or U24753 (N_24753,N_15028,N_17835);
nand U24754 (N_24754,N_18474,N_19443);
nor U24755 (N_24755,N_17812,N_18098);
nand U24756 (N_24756,N_16722,N_15939);
or U24757 (N_24757,N_15383,N_15171);
nor U24758 (N_24758,N_19802,N_19355);
and U24759 (N_24759,N_15851,N_17772);
or U24760 (N_24760,N_15567,N_16941);
nor U24761 (N_24761,N_17556,N_19656);
nand U24762 (N_24762,N_18362,N_17370);
and U24763 (N_24763,N_17930,N_18931);
nor U24764 (N_24764,N_18430,N_15598);
or U24765 (N_24765,N_16692,N_16005);
nand U24766 (N_24766,N_15506,N_18114);
nand U24767 (N_24767,N_19531,N_18694);
nand U24768 (N_24768,N_16227,N_16519);
and U24769 (N_24769,N_18983,N_15631);
nor U24770 (N_24770,N_17837,N_15960);
or U24771 (N_24771,N_16516,N_17992);
or U24772 (N_24772,N_18156,N_17498);
or U24773 (N_24773,N_19533,N_18798);
nor U24774 (N_24774,N_17687,N_15853);
and U24775 (N_24775,N_18838,N_18046);
and U24776 (N_24776,N_17275,N_19464);
and U24777 (N_24777,N_19748,N_17132);
xor U24778 (N_24778,N_17103,N_19134);
and U24779 (N_24779,N_18580,N_16185);
and U24780 (N_24780,N_18962,N_18088);
nand U24781 (N_24781,N_15000,N_19170);
or U24782 (N_24782,N_17950,N_17686);
or U24783 (N_24783,N_19040,N_18166);
or U24784 (N_24784,N_15440,N_19712);
nand U24785 (N_24785,N_18958,N_18239);
and U24786 (N_24786,N_15050,N_18515);
and U24787 (N_24787,N_17090,N_18781);
nor U24788 (N_24788,N_15755,N_15112);
and U24789 (N_24789,N_17854,N_18120);
and U24790 (N_24790,N_16328,N_17421);
nand U24791 (N_24791,N_19268,N_15546);
or U24792 (N_24792,N_18178,N_17326);
nor U24793 (N_24793,N_18381,N_15011);
nand U24794 (N_24794,N_18303,N_17212);
and U24795 (N_24795,N_16446,N_18656);
or U24796 (N_24796,N_15238,N_17872);
xor U24797 (N_24797,N_17522,N_19277);
nand U24798 (N_24798,N_17076,N_15145);
nor U24799 (N_24799,N_18771,N_15617);
nor U24800 (N_24800,N_16270,N_15737);
and U24801 (N_24801,N_18366,N_16563);
or U24802 (N_24802,N_17311,N_17732);
and U24803 (N_24803,N_16089,N_17615);
nand U24804 (N_24804,N_18975,N_15474);
nor U24805 (N_24805,N_16089,N_19033);
and U24806 (N_24806,N_17706,N_17290);
or U24807 (N_24807,N_15093,N_19718);
and U24808 (N_24808,N_19744,N_19751);
xor U24809 (N_24809,N_19973,N_18998);
nand U24810 (N_24810,N_16497,N_17729);
nand U24811 (N_24811,N_17703,N_16185);
and U24812 (N_24812,N_15825,N_19695);
and U24813 (N_24813,N_15033,N_18075);
nor U24814 (N_24814,N_18924,N_16274);
nor U24815 (N_24815,N_17904,N_17937);
nand U24816 (N_24816,N_16549,N_19736);
and U24817 (N_24817,N_15559,N_15621);
nor U24818 (N_24818,N_18759,N_17469);
and U24819 (N_24819,N_18103,N_18127);
nand U24820 (N_24820,N_17384,N_16995);
or U24821 (N_24821,N_19262,N_18411);
nand U24822 (N_24822,N_19801,N_18096);
nand U24823 (N_24823,N_18997,N_18853);
nand U24824 (N_24824,N_19124,N_16114);
nor U24825 (N_24825,N_19651,N_16495);
or U24826 (N_24826,N_19570,N_16881);
or U24827 (N_24827,N_18479,N_15455);
nor U24828 (N_24828,N_16915,N_15738);
nand U24829 (N_24829,N_18858,N_17912);
nor U24830 (N_24830,N_19087,N_15326);
nand U24831 (N_24831,N_17404,N_15663);
and U24832 (N_24832,N_15195,N_19063);
nand U24833 (N_24833,N_19667,N_16991);
or U24834 (N_24834,N_17824,N_17951);
and U24835 (N_24835,N_18171,N_18229);
or U24836 (N_24836,N_17583,N_18068);
and U24837 (N_24837,N_15602,N_15645);
and U24838 (N_24838,N_16354,N_16020);
nor U24839 (N_24839,N_19037,N_17014);
or U24840 (N_24840,N_17251,N_19139);
nand U24841 (N_24841,N_18569,N_16545);
nor U24842 (N_24842,N_18386,N_16366);
nor U24843 (N_24843,N_19093,N_19882);
or U24844 (N_24844,N_15987,N_15222);
nand U24845 (N_24845,N_17273,N_18306);
and U24846 (N_24846,N_18004,N_18425);
or U24847 (N_24847,N_19777,N_16349);
or U24848 (N_24848,N_19693,N_19947);
and U24849 (N_24849,N_18115,N_18911);
xor U24850 (N_24850,N_16219,N_17815);
nor U24851 (N_24851,N_18057,N_15917);
or U24852 (N_24852,N_15290,N_18858);
nand U24853 (N_24853,N_18398,N_19504);
or U24854 (N_24854,N_19316,N_17610);
xnor U24855 (N_24855,N_17301,N_16729);
nand U24856 (N_24856,N_17281,N_18756);
nand U24857 (N_24857,N_16554,N_15262);
or U24858 (N_24858,N_19724,N_15852);
nand U24859 (N_24859,N_15460,N_18379);
nand U24860 (N_24860,N_17217,N_15653);
nor U24861 (N_24861,N_19685,N_18793);
xnor U24862 (N_24862,N_19341,N_16027);
nor U24863 (N_24863,N_17481,N_17472);
or U24864 (N_24864,N_16931,N_16949);
nand U24865 (N_24865,N_19592,N_15940);
nand U24866 (N_24866,N_16356,N_16308);
or U24867 (N_24867,N_15190,N_17693);
and U24868 (N_24868,N_17386,N_18873);
nor U24869 (N_24869,N_19264,N_16578);
nand U24870 (N_24870,N_18156,N_19569);
and U24871 (N_24871,N_15415,N_17629);
nor U24872 (N_24872,N_17407,N_18221);
nor U24873 (N_24873,N_19552,N_18707);
nand U24874 (N_24874,N_18308,N_18157);
and U24875 (N_24875,N_17137,N_18872);
nor U24876 (N_24876,N_16511,N_17225);
or U24877 (N_24877,N_15385,N_17566);
nor U24878 (N_24878,N_16659,N_18370);
nor U24879 (N_24879,N_19379,N_16892);
and U24880 (N_24880,N_19285,N_19928);
nor U24881 (N_24881,N_19817,N_19270);
and U24882 (N_24882,N_18733,N_18826);
and U24883 (N_24883,N_17912,N_15429);
and U24884 (N_24884,N_17575,N_15913);
and U24885 (N_24885,N_19373,N_17856);
and U24886 (N_24886,N_16043,N_15559);
or U24887 (N_24887,N_19612,N_16565);
nand U24888 (N_24888,N_17401,N_19610);
nor U24889 (N_24889,N_19893,N_18421);
nor U24890 (N_24890,N_18309,N_18813);
and U24891 (N_24891,N_15334,N_18735);
and U24892 (N_24892,N_15359,N_15931);
or U24893 (N_24893,N_16688,N_19065);
nand U24894 (N_24894,N_18447,N_19774);
or U24895 (N_24895,N_16453,N_15079);
nand U24896 (N_24896,N_15188,N_19676);
and U24897 (N_24897,N_17530,N_15358);
and U24898 (N_24898,N_18786,N_16802);
and U24899 (N_24899,N_19192,N_18480);
nand U24900 (N_24900,N_19121,N_16445);
or U24901 (N_24901,N_19477,N_16394);
and U24902 (N_24902,N_17298,N_19082);
and U24903 (N_24903,N_15273,N_15948);
nor U24904 (N_24904,N_16473,N_15394);
or U24905 (N_24905,N_19505,N_16120);
or U24906 (N_24906,N_15987,N_17528);
or U24907 (N_24907,N_18305,N_15606);
nor U24908 (N_24908,N_19603,N_18528);
nor U24909 (N_24909,N_19297,N_18832);
and U24910 (N_24910,N_19941,N_15992);
and U24911 (N_24911,N_15287,N_19893);
and U24912 (N_24912,N_19068,N_17551);
and U24913 (N_24913,N_18080,N_17306);
nand U24914 (N_24914,N_16778,N_17056);
nor U24915 (N_24915,N_15863,N_17133);
or U24916 (N_24916,N_19441,N_18984);
and U24917 (N_24917,N_16689,N_17293);
xor U24918 (N_24918,N_16840,N_19258);
nor U24919 (N_24919,N_16527,N_18075);
nor U24920 (N_24920,N_19440,N_17666);
or U24921 (N_24921,N_19617,N_15558);
nand U24922 (N_24922,N_16559,N_16662);
nand U24923 (N_24923,N_17637,N_18834);
or U24924 (N_24924,N_17410,N_17474);
nand U24925 (N_24925,N_19030,N_18144);
nand U24926 (N_24926,N_17911,N_17899);
or U24927 (N_24927,N_15107,N_16403);
nor U24928 (N_24928,N_19085,N_15918);
nor U24929 (N_24929,N_17699,N_19646);
and U24930 (N_24930,N_15543,N_19246);
or U24931 (N_24931,N_18820,N_19450);
and U24932 (N_24932,N_17854,N_18343);
and U24933 (N_24933,N_19466,N_18008);
nand U24934 (N_24934,N_19867,N_17940);
or U24935 (N_24935,N_19784,N_15731);
and U24936 (N_24936,N_17688,N_19394);
and U24937 (N_24937,N_16859,N_18175);
and U24938 (N_24938,N_19909,N_18877);
nand U24939 (N_24939,N_19271,N_19566);
or U24940 (N_24940,N_16747,N_18504);
nor U24941 (N_24941,N_18988,N_16977);
nand U24942 (N_24942,N_15225,N_15049);
or U24943 (N_24943,N_17826,N_15953);
and U24944 (N_24944,N_15911,N_16369);
nor U24945 (N_24945,N_15587,N_18723);
nand U24946 (N_24946,N_15781,N_15596);
or U24947 (N_24947,N_19315,N_15804);
nand U24948 (N_24948,N_16125,N_15286);
nor U24949 (N_24949,N_17732,N_15781);
and U24950 (N_24950,N_18697,N_18060);
xor U24951 (N_24951,N_17564,N_16693);
nor U24952 (N_24952,N_15270,N_16097);
xor U24953 (N_24953,N_16718,N_15014);
and U24954 (N_24954,N_18635,N_18629);
and U24955 (N_24955,N_18358,N_18687);
nor U24956 (N_24956,N_15388,N_19768);
and U24957 (N_24957,N_16599,N_18505);
or U24958 (N_24958,N_16075,N_16111);
or U24959 (N_24959,N_19687,N_19080);
or U24960 (N_24960,N_18449,N_18498);
nand U24961 (N_24961,N_19990,N_16550);
nand U24962 (N_24962,N_19073,N_18729);
and U24963 (N_24963,N_19046,N_18811);
and U24964 (N_24964,N_18340,N_19244);
nor U24965 (N_24965,N_17123,N_16427);
and U24966 (N_24966,N_18868,N_17463);
nand U24967 (N_24967,N_15421,N_17630);
or U24968 (N_24968,N_15115,N_15356);
and U24969 (N_24969,N_16966,N_17060);
or U24970 (N_24970,N_17041,N_15938);
and U24971 (N_24971,N_18776,N_16763);
and U24972 (N_24972,N_17561,N_18492);
and U24973 (N_24973,N_15268,N_15802);
and U24974 (N_24974,N_15638,N_15858);
and U24975 (N_24975,N_19998,N_17113);
nor U24976 (N_24976,N_19366,N_19371);
nand U24977 (N_24977,N_18040,N_19485);
nor U24978 (N_24978,N_17100,N_19243);
and U24979 (N_24979,N_16579,N_19518);
or U24980 (N_24980,N_15141,N_16486);
xor U24981 (N_24981,N_15568,N_16704);
xnor U24982 (N_24982,N_16817,N_17670);
nor U24983 (N_24983,N_16891,N_19054);
or U24984 (N_24984,N_18736,N_16864);
and U24985 (N_24985,N_19167,N_17476);
nor U24986 (N_24986,N_19380,N_19573);
nor U24987 (N_24987,N_18011,N_17640);
or U24988 (N_24988,N_19178,N_17299);
nand U24989 (N_24989,N_15115,N_15853);
and U24990 (N_24990,N_19382,N_15675);
and U24991 (N_24991,N_16335,N_15361);
nor U24992 (N_24992,N_15901,N_19206);
or U24993 (N_24993,N_16139,N_15781);
nand U24994 (N_24994,N_15775,N_19714);
nor U24995 (N_24995,N_15802,N_16983);
nor U24996 (N_24996,N_17008,N_17375);
nand U24997 (N_24997,N_19554,N_16135);
and U24998 (N_24998,N_16645,N_17045);
or U24999 (N_24999,N_15434,N_16081);
nand UO_0 (O_0,N_22306,N_23799);
nand UO_1 (O_1,N_20495,N_23899);
and UO_2 (O_2,N_21576,N_24710);
and UO_3 (O_3,N_22428,N_22049);
nor UO_4 (O_4,N_21169,N_24320);
nand UO_5 (O_5,N_23444,N_24963);
and UO_6 (O_6,N_24134,N_22632);
nand UO_7 (O_7,N_20752,N_24382);
nor UO_8 (O_8,N_21573,N_21622);
nor UO_9 (O_9,N_22562,N_23587);
xor UO_10 (O_10,N_21700,N_20455);
or UO_11 (O_11,N_23892,N_21451);
nand UO_12 (O_12,N_20473,N_22100);
nand UO_13 (O_13,N_21218,N_20984);
nor UO_14 (O_14,N_23699,N_23545);
nor UO_15 (O_15,N_20881,N_21671);
nor UO_16 (O_16,N_24144,N_21315);
and UO_17 (O_17,N_21806,N_22659);
xor UO_18 (O_18,N_22370,N_23188);
nand UO_19 (O_19,N_23311,N_21212);
nor UO_20 (O_20,N_22010,N_22001);
and UO_21 (O_21,N_24688,N_23915);
nor UO_22 (O_22,N_24489,N_22845);
nand UO_23 (O_23,N_24695,N_23912);
nand UO_24 (O_24,N_20899,N_20522);
nor UO_25 (O_25,N_22817,N_22162);
nand UO_26 (O_26,N_22902,N_22666);
nand UO_27 (O_27,N_21987,N_20663);
nand UO_28 (O_28,N_21481,N_21931);
nand UO_29 (O_29,N_21246,N_22851);
nand UO_30 (O_30,N_24509,N_23931);
or UO_31 (O_31,N_24267,N_21697);
nor UO_32 (O_32,N_21929,N_24241);
and UO_33 (O_33,N_21647,N_20976);
and UO_34 (O_34,N_21122,N_22354);
and UO_35 (O_35,N_22805,N_24731);
nand UO_36 (O_36,N_24767,N_22501);
and UO_37 (O_37,N_22264,N_22122);
and UO_38 (O_38,N_21057,N_24886);
nand UO_39 (O_39,N_22292,N_21969);
and UO_40 (O_40,N_24655,N_24178);
nand UO_41 (O_41,N_23150,N_21843);
or UO_42 (O_42,N_22631,N_23178);
nand UO_43 (O_43,N_22947,N_23576);
and UO_44 (O_44,N_20820,N_23564);
nor UO_45 (O_45,N_23754,N_22475);
nor UO_46 (O_46,N_23448,N_20231);
nor UO_47 (O_47,N_23628,N_21019);
nand UO_48 (O_48,N_22432,N_21603);
or UO_49 (O_49,N_22257,N_22516);
xnor UO_50 (O_50,N_20642,N_22300);
and UO_51 (O_51,N_21805,N_21800);
or UO_52 (O_52,N_20694,N_20888);
and UO_53 (O_53,N_23850,N_23003);
or UO_54 (O_54,N_23352,N_24183);
and UO_55 (O_55,N_20062,N_22117);
nor UO_56 (O_56,N_23245,N_23740);
and UO_57 (O_57,N_24833,N_22484);
nand UO_58 (O_58,N_23820,N_24424);
nand UO_59 (O_59,N_20515,N_20192);
and UO_60 (O_60,N_23039,N_20475);
nand UO_61 (O_61,N_20423,N_22070);
nand UO_62 (O_62,N_21660,N_22905);
or UO_63 (O_63,N_22534,N_24974);
or UO_64 (O_64,N_24494,N_23652);
nand UO_65 (O_65,N_21699,N_23404);
nand UO_66 (O_66,N_23745,N_23728);
and UO_67 (O_67,N_24621,N_22310);
nor UO_68 (O_68,N_24238,N_23646);
nor UO_69 (O_69,N_23540,N_21183);
nand UO_70 (O_70,N_22421,N_20632);
or UO_71 (O_71,N_23043,N_20216);
and UO_72 (O_72,N_22706,N_21965);
nand UO_73 (O_73,N_24372,N_24784);
nand UO_74 (O_74,N_24079,N_23796);
and UO_75 (O_75,N_20327,N_24374);
or UO_76 (O_76,N_21126,N_22532);
or UO_77 (O_77,N_22227,N_23447);
nor UO_78 (O_78,N_20341,N_21383);
nand UO_79 (O_79,N_22728,N_20429);
and UO_80 (O_80,N_21932,N_23940);
and UO_81 (O_81,N_21986,N_20595);
nor UO_82 (O_82,N_23443,N_21261);
nor UO_83 (O_83,N_21897,N_20900);
nand UO_84 (O_84,N_23233,N_22163);
and UO_85 (O_85,N_20063,N_22338);
xnor UO_86 (O_86,N_23131,N_24746);
nor UO_87 (O_87,N_20956,N_22127);
and UO_88 (O_88,N_24403,N_23702);
and UO_89 (O_89,N_23044,N_24456);
nor UO_90 (O_90,N_24734,N_24354);
nor UO_91 (O_91,N_24256,N_24818);
and UO_92 (O_92,N_22486,N_22741);
and UO_93 (O_93,N_24443,N_24304);
and UO_94 (O_94,N_24052,N_22963);
and UO_95 (O_95,N_21113,N_24195);
and UO_96 (O_96,N_22431,N_23714);
nand UO_97 (O_97,N_21078,N_20847);
or UO_98 (O_98,N_20271,N_22349);
or UO_99 (O_99,N_22509,N_21559);
nor UO_100 (O_100,N_22298,N_23974);
or UO_101 (O_101,N_22201,N_21295);
nand UO_102 (O_102,N_21884,N_23549);
or UO_103 (O_103,N_21159,N_22858);
nor UO_104 (O_104,N_22525,N_23893);
nor UO_105 (O_105,N_23595,N_24305);
nor UO_106 (O_106,N_23432,N_24425);
nand UO_107 (O_107,N_20343,N_22991);
or UO_108 (O_108,N_24745,N_22857);
xor UO_109 (O_109,N_23857,N_21114);
nand UO_110 (O_110,N_24151,N_21109);
and UO_111 (O_111,N_22740,N_24008);
xor UO_112 (O_112,N_22319,N_23900);
nor UO_113 (O_113,N_20932,N_24798);
nand UO_114 (O_114,N_21031,N_22223);
nor UO_115 (O_115,N_24989,N_23424);
nor UO_116 (O_116,N_21294,N_21182);
nor UO_117 (O_117,N_22941,N_23355);
nand UO_118 (O_118,N_24216,N_20447);
nor UO_119 (O_119,N_22880,N_23826);
and UO_120 (O_120,N_24790,N_22585);
or UO_121 (O_121,N_21721,N_21646);
and UO_122 (O_122,N_21370,N_21421);
nor UO_123 (O_123,N_22553,N_24364);
nor UO_124 (O_124,N_21385,N_21549);
and UO_125 (O_125,N_23774,N_22161);
nand UO_126 (O_126,N_24907,N_21420);
or UO_127 (O_127,N_24359,N_22436);
and UO_128 (O_128,N_23257,N_22850);
and UO_129 (O_129,N_20489,N_22352);
or UO_130 (O_130,N_23722,N_24671);
and UO_131 (O_131,N_23453,N_23956);
and UO_132 (O_132,N_24854,N_23706);
or UO_133 (O_133,N_21045,N_23897);
nand UO_134 (O_134,N_20702,N_20123);
nor UO_135 (O_135,N_23422,N_21896);
and UO_136 (O_136,N_24205,N_22593);
and UO_137 (O_137,N_23149,N_20068);
and UO_138 (O_138,N_24765,N_24128);
nor UO_139 (O_139,N_23005,N_23869);
or UO_140 (O_140,N_20894,N_21832);
nor UO_141 (O_141,N_22521,N_20654);
nand UO_142 (O_142,N_24576,N_23483);
and UO_143 (O_143,N_21708,N_22482);
or UO_144 (O_144,N_23572,N_22255);
nor UO_145 (O_145,N_21855,N_21568);
and UO_146 (O_146,N_21020,N_21709);
and UO_147 (O_147,N_23944,N_21591);
nor UO_148 (O_148,N_23623,N_20529);
nor UO_149 (O_149,N_24788,N_24901);
or UO_150 (O_150,N_21015,N_21203);
nand UO_151 (O_151,N_23504,N_24561);
nand UO_152 (O_152,N_21268,N_23705);
and UO_153 (O_153,N_20322,N_20799);
or UO_154 (O_154,N_23436,N_21042);
and UO_155 (O_155,N_23109,N_24125);
xnor UO_156 (O_156,N_22997,N_21670);
and UO_157 (O_157,N_23023,N_20870);
nor UO_158 (O_158,N_22603,N_24999);
nand UO_159 (O_159,N_23856,N_22897);
nor UO_160 (O_160,N_20664,N_24325);
nor UO_161 (O_161,N_22104,N_20449);
or UO_162 (O_162,N_24712,N_23018);
and UO_163 (O_163,N_20085,N_22158);
or UO_164 (O_164,N_20012,N_22136);
and UO_165 (O_165,N_24067,N_20787);
nor UO_166 (O_166,N_22343,N_23758);
nand UO_167 (O_167,N_23506,N_20046);
nor UO_168 (O_168,N_23086,N_21657);
nand UO_169 (O_169,N_23469,N_20741);
and UO_170 (O_170,N_23530,N_22166);
xor UO_171 (O_171,N_24737,N_22032);
or UO_172 (O_172,N_21144,N_20777);
or UO_173 (O_173,N_22387,N_24020);
and UO_174 (O_174,N_23773,N_22650);
and UO_175 (O_175,N_21167,N_20175);
nor UO_176 (O_176,N_22874,N_24559);
and UO_177 (O_177,N_20933,N_23246);
and UO_178 (O_178,N_20955,N_23708);
and UO_179 (O_179,N_23769,N_24294);
and UO_180 (O_180,N_20259,N_21134);
nor UO_181 (O_181,N_20433,N_22871);
nor UO_182 (O_182,N_24188,N_20811);
and UO_183 (O_183,N_23724,N_22742);
nor UO_184 (O_184,N_23544,N_21796);
nor UO_185 (O_185,N_22124,N_23295);
and UO_186 (O_186,N_23712,N_23379);
and UO_187 (O_187,N_24190,N_22555);
or UO_188 (O_188,N_23327,N_23517);
or UO_189 (O_189,N_21840,N_23201);
nand UO_190 (O_190,N_24293,N_23130);
nand UO_191 (O_191,N_23972,N_22119);
or UO_192 (O_192,N_21077,N_24606);
and UO_193 (O_193,N_24660,N_21394);
nand UO_194 (O_194,N_22846,N_20628);
nand UO_195 (O_195,N_21098,N_22043);
nand UO_196 (O_196,N_21883,N_21522);
nor UO_197 (O_197,N_22508,N_20461);
and UO_198 (O_198,N_20665,N_22220);
or UO_199 (O_199,N_22552,N_23817);
nand UO_200 (O_200,N_21357,N_22138);
or UO_201 (O_201,N_23033,N_23430);
nor UO_202 (O_202,N_23250,N_23846);
nor UO_203 (O_203,N_23841,N_22196);
nor UO_204 (O_204,N_22108,N_22587);
and UO_205 (O_205,N_20960,N_23479);
and UO_206 (O_206,N_22824,N_24402);
xor UO_207 (O_207,N_23965,N_20266);
nor UO_208 (O_208,N_22212,N_22364);
or UO_209 (O_209,N_23613,N_21785);
or UO_210 (O_210,N_21977,N_20531);
nand UO_211 (O_211,N_23942,N_23741);
xnor UO_212 (O_212,N_22887,N_22191);
nor UO_213 (O_213,N_21867,N_21301);
and UO_214 (O_214,N_24613,N_23060);
nor UO_215 (O_215,N_20826,N_24912);
or UO_216 (O_216,N_22397,N_21598);
nor UO_217 (O_217,N_24068,N_23847);
nor UO_218 (O_218,N_21392,N_24251);
nand UO_219 (O_219,N_23076,N_24246);
nand UO_220 (O_220,N_20759,N_24644);
and UO_221 (O_221,N_23375,N_22716);
nor UO_222 (O_222,N_24687,N_21658);
and UO_223 (O_223,N_20188,N_23786);
or UO_224 (O_224,N_20966,N_21736);
nand UO_225 (O_225,N_20672,N_23210);
nand UO_226 (O_226,N_21508,N_24659);
or UO_227 (O_227,N_23871,N_22499);
nor UO_228 (O_228,N_23397,N_23137);
and UO_229 (O_229,N_22356,N_20860);
nor UO_230 (O_230,N_23127,N_22967);
nor UO_231 (O_231,N_23618,N_22937);
nand UO_232 (O_232,N_24626,N_23414);
or UO_233 (O_233,N_20873,N_23451);
nand UO_234 (O_234,N_21360,N_20027);
nor UO_235 (O_235,N_24300,N_20593);
nor UO_236 (O_236,N_21216,N_20073);
and UO_237 (O_237,N_20233,N_20815);
nand UO_238 (O_238,N_22835,N_23600);
or UO_239 (O_239,N_21569,N_22505);
and UO_240 (O_240,N_22760,N_21074);
nand UO_241 (O_241,N_23055,N_20297);
nand UO_242 (O_242,N_23015,N_24579);
nor UO_243 (O_243,N_24445,N_24360);
and UO_244 (O_244,N_22673,N_20993);
and UO_245 (O_245,N_20778,N_20189);
nand UO_246 (O_246,N_24233,N_20358);
nor UO_247 (O_247,N_23334,N_22477);
nor UO_248 (O_248,N_20336,N_22296);
nor UO_249 (O_249,N_21527,N_21631);
or UO_250 (O_250,N_22995,N_24051);
or UO_251 (O_251,N_24415,N_22048);
and UO_252 (O_252,N_21532,N_21107);
nand UO_253 (O_253,N_22175,N_24942);
and UO_254 (O_254,N_24544,N_21550);
or UO_255 (O_255,N_23114,N_23854);
and UO_256 (O_256,N_20644,N_21284);
nand UO_257 (O_257,N_21237,N_21879);
or UO_258 (O_258,N_20342,N_24405);
and UO_259 (O_259,N_23538,N_22584);
and UO_260 (O_260,N_22059,N_23625);
nor UO_261 (O_261,N_23641,N_20959);
nor UO_262 (O_262,N_23474,N_21984);
nand UO_263 (O_263,N_24812,N_24773);
nand UO_264 (O_264,N_24789,N_21664);
nor UO_265 (O_265,N_24394,N_21669);
and UO_266 (O_266,N_22823,N_21582);
nor UO_267 (O_267,N_23790,N_24623);
nand UO_268 (O_268,N_24363,N_23907);
xor UO_269 (O_269,N_24938,N_23228);
or UO_270 (O_270,N_24872,N_24914);
and UO_271 (O_271,N_23988,N_21445);
nor UO_272 (O_272,N_22394,N_21964);
nand UO_273 (O_273,N_22350,N_21457);
nand UO_274 (O_274,N_23253,N_22648);
nand UO_275 (O_275,N_22250,N_20408);
and UO_276 (O_276,N_20551,N_22044);
nand UO_277 (O_277,N_20677,N_22914);
nand UO_278 (O_278,N_21403,N_24536);
nor UO_279 (O_279,N_20659,N_20453);
or UO_280 (O_280,N_21012,N_23283);
xor UO_281 (O_281,N_23747,N_24618);
or UO_282 (O_282,N_24808,N_23809);
nand UO_283 (O_283,N_21715,N_22066);
nor UO_284 (O_284,N_21410,N_20315);
nand UO_285 (O_285,N_20334,N_20821);
nand UO_286 (O_286,N_24690,N_23484);
nor UO_287 (O_287,N_20048,N_21333);
or UO_288 (O_288,N_21253,N_22202);
and UO_289 (O_289,N_22884,N_22439);
nor UO_290 (O_290,N_20335,N_21868);
and UO_291 (O_291,N_22975,N_22282);
and UO_292 (O_292,N_21040,N_23937);
nand UO_293 (O_293,N_21386,N_22948);
and UO_294 (O_294,N_21590,N_24581);
nor UO_295 (O_295,N_22430,N_22703);
nor UO_296 (O_296,N_23263,N_23065);
nor UO_297 (O_297,N_23573,N_22033);
nor UO_298 (O_298,N_24882,N_20264);
or UO_299 (O_299,N_20274,N_23374);
nor UO_300 (O_300,N_20193,N_20319);
and UO_301 (O_301,N_24287,N_24413);
nor UO_302 (O_302,N_22537,N_20516);
or UO_303 (O_303,N_21630,N_21676);
and UO_304 (O_304,N_24093,N_20532);
nor UO_305 (O_305,N_20378,N_22605);
nand UO_306 (O_306,N_20005,N_21429);
and UO_307 (O_307,N_23035,N_24028);
nand UO_308 (O_308,N_23984,N_24897);
nand UO_309 (O_309,N_22221,N_21578);
nand UO_310 (O_310,N_24894,N_20042);
and UO_311 (O_311,N_22301,N_22168);
nand UO_312 (O_312,N_20397,N_20368);
and UO_313 (O_313,N_20399,N_24044);
nor UO_314 (O_314,N_24166,N_20097);
nor UO_315 (O_315,N_22483,N_21648);
or UO_316 (O_316,N_20754,N_22209);
nor UO_317 (O_317,N_23069,N_24805);
or UO_318 (O_318,N_24390,N_22996);
or UO_319 (O_319,N_20075,N_24609);
nor UO_320 (O_320,N_22512,N_24706);
nand UO_321 (O_321,N_22852,N_24285);
or UO_322 (O_322,N_24620,N_23627);
or UO_323 (O_323,N_21431,N_24280);
and UO_324 (O_324,N_22583,N_24602);
nor UO_325 (O_325,N_24995,N_20360);
and UO_326 (O_326,N_21617,N_20318);
and UO_327 (O_327,N_21489,N_22210);
nor UO_328 (O_328,N_21358,N_22459);
nor UO_329 (O_329,N_20751,N_20059);
or UO_330 (O_330,N_24035,N_24345);
and UO_331 (O_331,N_21231,N_24065);
and UO_332 (O_332,N_21623,N_23403);
nand UO_333 (O_333,N_20542,N_21679);
and UO_334 (O_334,N_20684,N_24462);
or UO_335 (O_335,N_20043,N_20014);
or UO_336 (O_336,N_20060,N_20626);
nand UO_337 (O_337,N_23922,N_21995);
or UO_338 (O_338,N_24824,N_21208);
xor UO_339 (O_339,N_24451,N_20034);
or UO_340 (O_340,N_21008,N_22113);
xnor UO_341 (O_341,N_22620,N_21743);
nor UO_342 (O_342,N_20705,N_23332);
nor UO_343 (O_343,N_21321,N_20015);
nand UO_344 (O_344,N_21597,N_24059);
or UO_345 (O_345,N_23890,N_22077);
nand UO_346 (O_346,N_21232,N_20178);
nand UO_347 (O_347,N_24632,N_24792);
nand UO_348 (O_348,N_22504,N_20849);
or UO_349 (O_349,N_21523,N_20594);
nor UO_350 (O_350,N_24157,N_24591);
nor UO_351 (O_351,N_22086,N_22724);
nand UO_352 (O_352,N_22038,N_23302);
nand UO_353 (O_353,N_21025,N_23836);
and UO_354 (O_354,N_23328,N_24800);
nand UO_355 (O_355,N_24227,N_24440);
nand UO_356 (O_356,N_23244,N_24736);
or UO_357 (O_357,N_20494,N_21427);
or UO_358 (O_358,N_21537,N_20366);
or UO_359 (O_359,N_22667,N_20080);
nor UO_360 (O_360,N_22865,N_22681);
xor UO_361 (O_361,N_20445,N_20482);
and UO_362 (O_362,N_24517,N_21180);
and UO_363 (O_363,N_24504,N_20134);
nand UO_364 (O_364,N_23229,N_20159);
and UO_365 (O_365,N_22018,N_23179);
or UO_366 (O_366,N_24321,N_20549);
xor UO_367 (O_367,N_21186,N_20261);
or UO_368 (O_368,N_24029,N_24837);
and UO_369 (O_369,N_24449,N_22934);
or UO_370 (O_370,N_20617,N_23803);
or UO_371 (O_371,N_22285,N_23313);
nand UO_372 (O_372,N_24972,N_23002);
nand UO_373 (O_373,N_23552,N_22383);
or UO_374 (O_374,N_22859,N_23308);
and UO_375 (O_375,N_24457,N_22373);
and UO_376 (O_376,N_23180,N_21275);
or UO_377 (O_377,N_23542,N_22036);
xor UO_378 (O_378,N_21187,N_21035);
and UO_379 (O_379,N_21046,N_20624);
and UO_380 (O_380,N_20163,N_21173);
xor UO_381 (O_381,N_22629,N_22065);
nor UO_382 (O_382,N_21946,N_22315);
nand UO_383 (O_383,N_22556,N_22327);
nor UO_384 (O_384,N_24670,N_23167);
nand UO_385 (O_385,N_20667,N_21433);
or UO_386 (O_386,N_23386,N_22198);
nor UO_387 (O_387,N_23541,N_22422);
and UO_388 (O_388,N_23380,N_21009);
nand UO_389 (O_389,N_21075,N_21774);
or UO_390 (O_390,N_23117,N_21266);
nor UO_391 (O_391,N_22325,N_22578);
and UO_392 (O_392,N_21058,N_22000);
nor UO_393 (O_393,N_24691,N_24021);
nor UO_394 (O_394,N_24480,N_22156);
or UO_395 (O_395,N_24219,N_23767);
nand UO_396 (O_396,N_21190,N_23454);
or UO_397 (O_397,N_22453,N_24336);
nand UO_398 (O_398,N_20214,N_24332);
and UO_399 (O_399,N_22709,N_23994);
and UO_400 (O_400,N_24732,N_24149);
nand UO_401 (O_401,N_21872,N_22116);
nand UO_402 (O_402,N_20661,N_24297);
or UO_403 (O_403,N_22707,N_20580);
or UO_404 (O_404,N_23558,N_22761);
or UO_405 (O_405,N_20382,N_24041);
nor UO_406 (O_406,N_24919,N_20038);
or UO_407 (O_407,N_20557,N_21484);
nand UO_408 (O_408,N_21225,N_24704);
nor UO_409 (O_409,N_24037,N_23598);
nand UO_410 (O_410,N_23416,N_23147);
nor UO_411 (O_411,N_20800,N_23894);
or UO_412 (O_412,N_23832,N_24410);
and UO_413 (O_413,N_24647,N_20487);
and UO_414 (O_414,N_20729,N_22770);
and UO_415 (O_415,N_23853,N_24512);
nor UO_416 (O_416,N_24172,N_20481);
nor UO_417 (O_417,N_20856,N_24594);
nand UO_418 (O_418,N_22916,N_23300);
or UO_419 (O_419,N_23813,N_21695);
nand UO_420 (O_420,N_23068,N_21125);
and UO_421 (O_421,N_20243,N_24599);
nor UO_422 (O_422,N_23499,N_20225);
or UO_423 (O_423,N_21094,N_22794);
nor UO_424 (O_424,N_21172,N_20924);
nor UO_425 (O_425,N_22693,N_24073);
nand UO_426 (O_426,N_23346,N_24904);
nand UO_427 (O_427,N_20260,N_24362);
nand UO_428 (O_428,N_23338,N_24398);
nor UO_429 (O_429,N_22365,N_20874);
and UO_430 (O_430,N_20699,N_24019);
or UO_431 (O_431,N_20377,N_20308);
nor UO_432 (O_432,N_21661,N_22951);
or UO_433 (O_433,N_21601,N_23174);
or UO_434 (O_434,N_23231,N_24884);
nor UO_435 (O_435,N_21194,N_24269);
nand UO_436 (O_436,N_22345,N_20182);
or UO_437 (O_437,N_22785,N_24106);
or UO_438 (O_438,N_22193,N_21645);
and UO_439 (O_439,N_22446,N_21688);
nand UO_440 (O_440,N_21039,N_23539);
and UO_441 (O_441,N_23040,N_24585);
or UO_442 (O_442,N_24182,N_22739);
nand UO_443 (O_443,N_23693,N_24603);
or UO_444 (O_444,N_24807,N_21299);
nand UO_445 (O_445,N_23185,N_21731);
nor UO_446 (O_446,N_22646,N_24204);
nand UO_447 (O_447,N_24026,N_24467);
and UO_448 (O_448,N_23194,N_20929);
nand UO_449 (O_449,N_22598,N_23381);
and UO_450 (O_450,N_22169,N_22549);
nor UO_451 (O_451,N_21450,N_23778);
or UO_452 (O_452,N_20838,N_22368);
nand UO_453 (O_453,N_21441,N_23995);
and UO_454 (O_454,N_24062,N_23036);
xnor UO_455 (O_455,N_20407,N_23027);
or UO_456 (O_456,N_21943,N_21586);
or UO_457 (O_457,N_22003,N_20810);
and UO_458 (O_458,N_20417,N_23091);
or UO_459 (O_459,N_23398,N_23535);
or UO_460 (O_460,N_20440,N_24668);
and UO_461 (O_461,N_24641,N_23473);
nand UO_462 (O_462,N_20816,N_24116);
nand UO_463 (O_463,N_22690,N_24466);
nand UO_464 (O_464,N_24448,N_22732);
nor UO_465 (O_465,N_22927,N_20200);
xor UO_466 (O_466,N_23657,N_20112);
nand UO_467 (O_467,N_23480,N_23077);
and UO_468 (O_468,N_21467,N_21827);
or UO_469 (O_469,N_22731,N_23098);
or UO_470 (O_470,N_24562,N_21944);
nor UO_471 (O_471,N_23744,N_23335);
or UO_472 (O_472,N_21773,N_24240);
nand UO_473 (O_473,N_22745,N_22753);
and UO_474 (O_474,N_20530,N_23136);
or UO_475 (O_475,N_22395,N_23987);
nand UO_476 (O_476,N_22810,N_20818);
nor UO_477 (O_477,N_23680,N_23029);
or UO_478 (O_478,N_21956,N_20383);
and UO_479 (O_479,N_21320,N_22073);
and UO_480 (O_480,N_22130,N_22427);
nor UO_481 (O_481,N_20784,N_24257);
or UO_482 (O_482,N_20541,N_21504);
and UO_483 (O_483,N_22670,N_21680);
and UO_484 (O_484,N_23282,N_23927);
or UO_485 (O_485,N_21939,N_20326);
and UO_486 (O_486,N_21092,N_22485);
nor UO_487 (O_487,N_21353,N_22390);
and UO_488 (O_488,N_20128,N_24366);
nor UO_489 (O_489,N_24135,N_24309);
and UO_490 (O_490,N_22554,N_23777);
nand UO_491 (O_491,N_23238,N_22717);
nand UO_492 (O_492,N_23333,N_20136);
nand UO_493 (O_493,N_22932,N_23016);
nor UO_494 (O_494,N_23351,N_24043);
and UO_495 (O_495,N_24600,N_21886);
nor UO_496 (O_496,N_22973,N_21280);
or UO_497 (O_497,N_20263,N_21205);
or UO_498 (O_498,N_24264,N_24115);
or UO_499 (O_499,N_20674,N_20609);
nor UO_500 (O_500,N_20219,N_22046);
nand UO_501 (O_501,N_20676,N_23678);
and UO_502 (O_502,N_21256,N_22087);
and UO_503 (O_503,N_22180,N_22665);
or UO_504 (O_504,N_20994,N_22757);
and UO_505 (O_505,N_23808,N_22790);
or UO_506 (O_506,N_24493,N_20570);
nand UO_507 (O_507,N_21038,N_23101);
and UO_508 (O_508,N_21729,N_21497);
nand UO_509 (O_509,N_24248,N_21192);
nor UO_510 (O_510,N_20031,N_23064);
or UO_511 (O_511,N_23290,N_20509);
or UO_512 (O_512,N_22836,N_24236);
nor UO_513 (O_513,N_21826,N_24066);
or UO_514 (O_514,N_23309,N_23659);
and UO_515 (O_515,N_21213,N_24702);
and UO_516 (O_516,N_23042,N_21440);
nor UO_517 (O_517,N_20972,N_22011);
nand UO_518 (O_518,N_22297,N_21105);
nand UO_519 (O_519,N_21473,N_21437);
nor UO_520 (O_520,N_22701,N_20934);
or UO_521 (O_521,N_21456,N_21463);
xnor UO_522 (O_522,N_21355,N_24860);
or UO_523 (O_523,N_24121,N_23881);
or UO_524 (O_524,N_20635,N_23565);
and UO_525 (O_525,N_20988,N_22450);
and UO_526 (O_526,N_24967,N_22470);
nor UO_527 (O_527,N_22879,N_20918);
nor UO_528 (O_528,N_21080,N_22287);
or UO_529 (O_529,N_21349,N_20281);
and UO_530 (O_530,N_24388,N_23533);
xor UO_531 (O_531,N_20518,N_22802);
and UO_532 (O_532,N_20950,N_21050);
xor UO_533 (O_533,N_20974,N_24096);
or UO_534 (O_534,N_22682,N_22307);
nand UO_535 (O_535,N_20969,N_21279);
or UO_536 (O_536,N_21210,N_20369);
nor UO_537 (O_537,N_20033,N_22213);
and UO_538 (O_538,N_20181,N_24646);
nor UO_539 (O_539,N_20602,N_24485);
or UO_540 (O_540,N_24842,N_20296);
or UO_541 (O_541,N_21061,N_24846);
and UO_542 (O_542,N_24369,N_24921);
nand UO_543 (O_543,N_23574,N_23521);
or UO_544 (O_544,N_24569,N_22634);
nand UO_545 (O_545,N_21882,N_23795);
nor UO_546 (O_546,N_20245,N_22219);
and UO_547 (O_547,N_21920,N_24651);
nor UO_548 (O_548,N_23930,N_23634);
and UO_549 (O_549,N_21505,N_21836);
and UO_550 (O_550,N_20750,N_24697);
nand UO_551 (O_551,N_21717,N_21328);
nand UO_552 (O_552,N_22643,N_20471);
nand UO_553 (O_553,N_20204,N_21354);
nand UO_554 (O_554,N_22526,N_22134);
nor UO_555 (O_555,N_24806,N_22170);
nand UO_556 (O_556,N_20848,N_24283);
nand UO_557 (O_557,N_21372,N_21036);
nand UO_558 (O_558,N_23511,N_20999);
nor UO_559 (O_559,N_22843,N_23402);
nor UO_560 (O_560,N_21021,N_22111);
and UO_561 (O_561,N_21155,N_23272);
nand UO_562 (O_562,N_23315,N_21121);
and UO_563 (O_563,N_20629,N_24714);
nand UO_564 (O_564,N_20846,N_23007);
nand UO_565 (O_565,N_20299,N_20879);
and UO_566 (O_566,N_23663,N_20686);
and UO_567 (O_567,N_21163,N_21572);
xnor UO_568 (O_568,N_24452,N_22624);
and UO_569 (O_569,N_24039,N_20992);
nand UO_570 (O_570,N_21885,N_24482);
nand UO_571 (O_571,N_20668,N_23719);
or UO_572 (O_572,N_22433,N_24893);
or UO_573 (O_573,N_22226,N_23183);
and UO_574 (O_574,N_23420,N_21841);
or UO_575 (O_575,N_23551,N_24378);
nor UO_576 (O_576,N_21769,N_23367);
nor UO_577 (O_577,N_20125,N_24936);
and UO_578 (O_578,N_23926,N_20923);
nor UO_579 (O_579,N_22799,N_23866);
nor UO_580 (O_580,N_23105,N_20289);
or UO_581 (O_581,N_21175,N_21500);
nand UO_582 (O_582,N_24099,N_22595);
or UO_583 (O_583,N_22236,N_23998);
nor UO_584 (O_584,N_21698,N_21130);
nand UO_585 (O_585,N_21257,N_20619);
nor UO_586 (O_586,N_23433,N_21719);
and UO_587 (O_587,N_23278,N_22440);
nand UO_588 (O_588,N_24162,N_21341);
and UO_589 (O_589,N_20565,N_23864);
or UO_590 (O_590,N_22958,N_22479);
or UO_591 (O_591,N_24983,N_21499);
and UO_592 (O_592,N_23916,N_24113);
and UO_593 (O_593,N_21751,N_21912);
or UO_594 (O_594,N_21961,N_23782);
nand UO_595 (O_595,N_20257,N_23428);
nand UO_596 (O_596,N_20237,N_21666);
or UO_597 (O_597,N_24943,N_21663);
and UO_598 (O_598,N_24853,N_22093);
nor UO_599 (O_599,N_20436,N_21802);
or UO_600 (O_600,N_24006,N_24521);
and UO_601 (O_601,N_21557,N_24198);
or UO_602 (O_602,N_21332,N_24654);
or UO_603 (O_603,N_24358,N_22416);
nor UO_604 (O_604,N_24988,N_20161);
nor UO_605 (O_605,N_20389,N_21696);
nand UO_606 (O_606,N_23843,N_22569);
nand UO_607 (O_607,N_20643,N_21954);
and UO_608 (O_608,N_24555,N_24488);
or UO_609 (O_609,N_22148,N_20921);
or UO_610 (O_610,N_21498,N_23417);
nor UO_611 (O_611,N_20603,N_23222);
nand UO_612 (O_612,N_20246,N_21334);
nand UO_613 (O_613,N_20757,N_20177);
nor UO_614 (O_614,N_24420,N_24104);
or UO_615 (O_615,N_22849,N_22076);
or UO_616 (O_616,N_21718,N_22766);
nand UO_617 (O_617,N_22853,N_21014);
and UO_618 (O_618,N_24042,N_23012);
nand UO_619 (O_619,N_21893,N_21828);
nand UO_620 (O_620,N_21908,N_20822);
xor UO_621 (O_621,N_24787,N_23715);
or UO_622 (O_622,N_21989,N_24834);
nor UO_623 (O_623,N_22045,N_20024);
nand UO_624 (O_624,N_23083,N_23792);
and UO_625 (O_625,N_20426,N_21196);
and UO_626 (O_626,N_24851,N_22570);
nand UO_627 (O_627,N_22833,N_21976);
nand UO_628 (O_628,N_24997,N_21366);
and UO_629 (O_629,N_21561,N_21338);
and UO_630 (O_630,N_24355,N_20813);
nand UO_631 (O_631,N_24437,N_23193);
or UO_632 (O_632,N_24381,N_22791);
and UO_633 (O_633,N_21579,N_21927);
or UO_634 (O_634,N_20218,N_20490);
nand UO_635 (O_635,N_20051,N_24181);
or UO_636 (O_636,N_22002,N_24675);
or UO_637 (O_637,N_21096,N_20783);
and UO_638 (O_638,N_23515,N_22901);
nand UO_639 (O_639,N_24976,N_20562);
nor UO_640 (O_640,N_22013,N_20732);
and UO_641 (O_641,N_24155,N_22809);
or UO_642 (O_642,N_20148,N_23716);
and UO_643 (O_643,N_20836,N_23195);
nor UO_644 (O_644,N_22351,N_22985);
and UO_645 (O_645,N_21458,N_21652);
nor UO_646 (O_646,N_21426,N_22617);
and UO_647 (O_647,N_24622,N_20637);
or UO_648 (O_648,N_24491,N_20022);
nor UO_649 (O_649,N_24281,N_24564);
and UO_650 (O_650,N_21632,N_24718);
nor UO_651 (O_651,N_20802,N_23134);
nor UO_652 (O_652,N_21048,N_22517);
nand UO_653 (O_653,N_22067,N_21614);
nand UO_654 (O_654,N_23726,N_21981);
nor UO_655 (O_655,N_24611,N_22530);
and UO_656 (O_656,N_23258,N_22923);
xor UO_657 (O_657,N_23437,N_20995);
nor UO_658 (O_658,N_20421,N_23163);
or UO_659 (O_659,N_20275,N_23373);
and UO_660 (O_660,N_21792,N_24385);
or UO_661 (O_661,N_24542,N_21892);
nor UO_662 (O_662,N_24375,N_22016);
nand UO_663 (O_663,N_24503,N_23435);
nand UO_664 (O_664,N_23383,N_21930);
nor UO_665 (O_665,N_21399,N_24045);
nand UO_666 (O_666,N_22051,N_24268);
nand UO_667 (O_667,N_21361,N_24048);
and UO_668 (O_668,N_21135,N_20765);
or UO_669 (O_669,N_24100,N_22780);
and UO_670 (O_670,N_24191,N_22109);
and UO_671 (O_671,N_20117,N_23175);
and UO_672 (O_672,N_22660,N_23635);
and UO_673 (O_673,N_23615,N_23967);
or UO_674 (O_674,N_21336,N_21539);
nand UO_675 (O_675,N_22474,N_23104);
nand UO_676 (O_676,N_22490,N_22966);
nand UO_677 (O_677,N_21917,N_21111);
nor UO_678 (O_678,N_22518,N_22727);
or UO_679 (O_679,N_24981,N_21848);
nor UO_680 (O_680,N_21102,N_21726);
or UO_681 (O_681,N_24434,N_22194);
nand UO_682 (O_682,N_21864,N_22873);
and UO_683 (O_683,N_24401,N_22153);
and UO_684 (O_684,N_21124,N_22402);
nor UO_685 (O_685,N_24565,N_20116);
nand UO_686 (O_686,N_21822,N_23914);
nand UO_687 (O_687,N_23720,N_22861);
nor UO_688 (O_688,N_24058,N_23463);
xor UO_689 (O_689,N_22435,N_24945);
nand UO_690 (O_690,N_21624,N_22494);
nor UO_691 (O_691,N_23976,N_23648);
nor UO_692 (O_692,N_20891,N_21677);
or UO_693 (O_693,N_21026,N_21062);
or UO_694 (O_694,N_23743,N_22316);
nor UO_695 (O_695,N_22922,N_21894);
or UO_696 (O_696,N_22150,N_22069);
nand UO_697 (O_697,N_23997,N_21090);
or UO_698 (O_698,N_24465,N_22704);
nand UO_699 (O_699,N_22826,N_22423);
and UO_700 (O_700,N_23526,N_22410);
nand UO_701 (O_701,N_21273,N_21082);
or UO_702 (O_702,N_21028,N_21543);
and UO_703 (O_703,N_24604,N_21351);
or UO_704 (O_704,N_22895,N_23286);
and UO_705 (O_705,N_24327,N_22920);
or UO_706 (O_706,N_22331,N_22586);
or UO_707 (O_707,N_24423,N_21803);
nor UO_708 (O_708,N_23303,N_20072);
nor UO_709 (O_709,N_21808,N_21980);
nand UO_710 (O_710,N_20514,N_20288);
nand UO_711 (O_711,N_20236,N_21975);
or UO_712 (O_712,N_20224,N_20909);
nand UO_713 (O_713,N_22702,N_24324);
or UO_714 (O_714,N_20916,N_24102);
or UO_715 (O_715,N_24284,N_20122);
nor UO_716 (O_716,N_21304,N_22870);
or UO_717 (O_717,N_22885,N_21999);
or UO_718 (O_718,N_21350,N_20220);
and UO_719 (O_719,N_21602,N_20793);
and UO_720 (O_720,N_23365,N_24057);
nor UO_721 (O_721,N_23122,N_20293);
nor UO_722 (O_722,N_20589,N_22597);
nand UO_723 (O_723,N_21356,N_21662);
and UO_724 (O_724,N_20430,N_22234);
or UO_725 (O_725,N_20110,N_23985);
nor UO_726 (O_726,N_21887,N_21681);
nand UO_727 (O_727,N_22915,N_21285);
or UO_728 (O_728,N_20902,N_20179);
nand UO_729 (O_729,N_23094,N_21503);
and UO_730 (O_730,N_21136,N_21202);
or UO_731 (O_731,N_20446,N_24475);
nand UO_732 (O_732,N_22095,N_23575);
xnor UO_733 (O_733,N_23896,N_24289);
and UO_734 (O_734,N_20465,N_23208);
nand UO_735 (O_735,N_24262,N_23770);
or UO_736 (O_736,N_21034,N_21145);
nor UO_737 (O_737,N_23887,N_22713);
nand UO_738 (O_738,N_20695,N_20427);
nand UO_739 (O_739,N_20406,N_23845);
nand UO_740 (O_740,N_24705,N_21119);
nand UO_741 (O_741,N_24958,N_24000);
nand UO_742 (O_742,N_21701,N_24748);
nor UO_743 (O_743,N_22936,N_23531);
nand UO_744 (O_744,N_24383,N_21970);
and UO_745 (O_745,N_23918,N_21438);
or UO_746 (O_746,N_24396,N_20153);
nand UO_747 (O_747,N_23878,N_21425);
nor UO_748 (O_748,N_20194,N_21739);
or UO_749 (O_749,N_23677,N_20375);
nand UO_750 (O_750,N_24373,N_22208);
nor UO_751 (O_751,N_22165,N_23989);
nor UO_752 (O_752,N_20964,N_22164);
nand UO_753 (O_753,N_20492,N_22881);
and UO_754 (O_754,N_21323,N_22619);
and UO_755 (O_755,N_20249,N_20512);
and UO_756 (O_756,N_23048,N_20428);
nor UO_757 (O_757,N_23651,N_20472);
or UO_758 (O_758,N_23031,N_24250);
nand UO_759 (O_759,N_22762,N_24829);
or UO_760 (O_760,N_21667,N_23694);
nor UO_761 (O_761,N_20865,N_21972);
or UO_762 (O_762,N_20309,N_24888);
nand UO_763 (O_763,N_20965,N_20827);
nand UO_764 (O_764,N_24738,N_22145);
nand UO_765 (O_765,N_22816,N_23468);
nand UO_766 (O_766,N_22759,N_22197);
and UO_767 (O_767,N_24180,N_23645);
and UO_768 (O_768,N_20744,N_23990);
nor UO_769 (O_769,N_21851,N_22415);
or UO_770 (O_770,N_21037,N_24816);
and UO_771 (O_771,N_21554,N_21963);
nor UO_772 (O_772,N_24270,N_20149);
or UO_773 (O_773,N_24163,N_20590);
or UO_774 (O_774,N_22658,N_21288);
nor UO_775 (O_775,N_24524,N_22454);
nand UO_776 (O_776,N_21060,N_23734);
or UO_777 (O_777,N_21177,N_24498);
nor UO_778 (O_778,N_20414,N_24571);
or UO_779 (O_779,N_20569,N_21521);
or UO_780 (O_780,N_20464,N_22542);
nand UO_781 (O_781,N_20937,N_22159);
or UO_782 (O_782,N_22812,N_23216);
or UO_783 (O_783,N_20010,N_23700);
nor UO_784 (O_784,N_22929,N_24864);
nor UO_785 (O_785,N_22393,N_21000);
or UO_786 (O_786,N_22825,N_21516);
nor UO_787 (O_787,N_20317,N_22588);
nand UO_788 (O_788,N_24636,N_23337);
and UO_789 (O_789,N_21223,N_20251);
nand UO_790 (O_790,N_22388,N_20298);
and UO_791 (O_791,N_23721,N_23073);
nor UO_792 (O_792,N_22096,N_22320);
nor UO_793 (O_793,N_24917,N_23284);
and UO_794 (O_794,N_23666,N_23780);
or UO_795 (O_795,N_21276,N_23495);
nand UO_796 (O_796,N_22412,N_23577);
nor UO_797 (O_797,N_20032,N_22131);
nand UO_798 (O_798,N_22206,N_22063);
or UO_799 (O_799,N_23191,N_23921);
or UO_800 (O_800,N_23126,N_22372);
nor UO_801 (O_801,N_21238,N_21781);
nor UO_802 (O_802,N_24534,N_24167);
or UO_803 (O_803,N_23153,N_20521);
nand UO_804 (O_804,N_21948,N_23637);
xnor UO_805 (O_805,N_23923,N_24658);
nor UO_806 (O_806,N_24138,N_20792);
nor UO_807 (O_807,N_24272,N_24303);
and UO_808 (O_808,N_22289,N_22984);
nor UO_809 (O_809,N_24526,N_24147);
or UO_810 (O_810,N_24352,N_20130);
or UO_811 (O_811,N_21570,N_24470);
and UO_812 (O_812,N_24112,N_23277);
and UO_813 (O_813,N_24274,N_24724);
or UO_814 (O_814,N_24196,N_22891);
nor UO_815 (O_815,N_24924,N_24001);
nand UO_816 (O_816,N_23986,N_20171);
nor UO_817 (O_817,N_20459,N_23181);
nand UO_818 (O_818,N_22793,N_23753);
or UO_819 (O_819,N_21493,N_23320);
nand UO_820 (O_820,N_23793,N_24528);
nor UO_821 (O_821,N_22360,N_24598);
nor UO_822 (O_822,N_20241,N_22426);
and UO_823 (O_823,N_20505,N_23932);
or UO_824 (O_824,N_23611,N_20817);
or UO_825 (O_825,N_20155,N_21613);
nor UO_826 (O_826,N_20098,N_20958);
or UO_827 (O_827,N_21720,N_21636);
nor UO_828 (O_828,N_22763,N_21820);
and UO_829 (O_829,N_20145,N_23322);
nor UO_830 (O_830,N_24994,N_23410);
or UO_831 (O_831,N_24117,N_23760);
nand UO_832 (O_832,N_24004,N_20722);
and UO_833 (O_833,N_23877,N_23442);
and UO_834 (O_834,N_22348,N_21243);
or UO_835 (O_835,N_23550,N_20026);
nor UO_836 (O_836,N_23471,N_20401);
nor UO_837 (O_837,N_21486,N_23080);
nand UO_838 (O_838,N_20905,N_23274);
and UO_839 (O_839,N_21643,N_22980);
nor UO_840 (O_840,N_24177,N_21862);
nand UO_841 (O_841,N_22188,N_22172);
nor UO_842 (O_842,N_20634,N_24210);
nand UO_843 (O_843,N_23822,N_22889);
nor UO_844 (O_844,N_23557,N_20118);
and UO_845 (O_845,N_24803,N_23629);
or UO_846 (O_846,N_22559,N_20240);
or UO_847 (O_847,N_23891,N_24980);
or UO_848 (O_848,N_20347,N_22311);
nor UO_849 (O_849,N_21551,N_21116);
or UO_850 (O_850,N_23034,N_20344);
nor UO_851 (O_851,N_24617,N_23704);
nand UO_852 (O_852,N_20679,N_24545);
nor UO_853 (O_853,N_23691,N_20277);
or UO_854 (O_854,N_22405,N_20835);
or UO_855 (O_855,N_20131,N_21470);
or UO_856 (O_856,N_24531,N_20556);
nand UO_857 (O_857,N_21439,N_20093);
or UO_858 (O_858,N_20587,N_22784);
or UO_859 (O_859,N_20788,N_23672);
and UO_860 (O_860,N_23583,N_23512);
and UO_861 (O_861,N_23936,N_20890);
nor UO_862 (O_862,N_23920,N_21922);
and UO_863 (O_863,N_23214,N_22303);
and UO_864 (O_864,N_24431,N_21693);
or UO_865 (O_865,N_21938,N_23528);
nor UO_866 (O_866,N_24131,N_20206);
or UO_867 (O_867,N_23794,N_20611);
xor UO_868 (O_868,N_24184,N_22700);
and UO_869 (O_869,N_23639,N_24441);
xor UO_870 (O_870,N_22626,N_24563);
or UO_871 (O_871,N_24487,N_21377);
xor UO_872 (O_872,N_20535,N_20508);
or UO_873 (O_873,N_21684,N_24552);
nor UO_874 (O_874,N_20912,N_23434);
xnor UO_875 (O_875,N_23232,N_23382);
nand UO_876 (O_876,N_21873,N_24091);
and UO_877 (O_877,N_22956,N_22580);
or UO_878 (O_878,N_22434,N_23791);
xnor UO_879 (O_879,N_24365,N_22178);
nor UO_880 (O_880,N_20013,N_24119);
and UO_881 (O_881,N_21760,N_22935);
and UO_882 (O_882,N_22531,N_24220);
or UO_883 (O_883,N_20989,N_20330);
and UO_884 (O_884,N_21509,N_21289);
nor UO_885 (O_885,N_22893,N_20198);
nand UO_886 (O_886,N_24377,N_21724);
and UO_887 (O_887,N_20633,N_21395);
xor UO_888 (O_888,N_21653,N_22602);
or UO_889 (O_889,N_23019,N_20419);
or UO_890 (O_890,N_22090,N_24887);
or UO_891 (O_891,N_20721,N_24217);
or UO_892 (O_892,N_20648,N_24087);
or UO_893 (O_893,N_21825,N_20100);
and UO_894 (O_894,N_20796,N_22056);
and UO_895 (O_895,N_24719,N_23710);
or UO_896 (O_896,N_24414,N_23737);
and UO_897 (O_897,N_24583,N_23472);
or UO_898 (O_898,N_23831,N_24496);
nor UO_899 (O_899,N_24796,N_22042);
and UO_900 (O_900,N_24903,N_20781);
or UO_901 (O_901,N_22606,N_24089);
and UO_902 (O_902,N_20559,N_23852);
and UO_903 (O_903,N_23591,N_22550);
and UO_904 (O_904,N_24624,N_24189);
or UO_905 (O_905,N_23390,N_24154);
nor UO_906 (O_906,N_24978,N_22910);
nor UO_907 (O_907,N_22933,N_22192);
and UO_908 (O_908,N_20519,N_22355);
nor UO_909 (O_909,N_21252,N_22030);
xor UO_910 (O_910,N_21022,N_24680);
and UO_911 (O_911,N_20618,N_23090);
nand UO_912 (O_912,N_21189,N_21322);
and UO_913 (O_913,N_23205,N_21239);
and UO_914 (O_914,N_24011,N_21391);
nand UO_915 (O_915,N_22419,N_22102);
or UO_916 (O_916,N_22267,N_23486);
xnor UO_917 (O_917,N_24520,N_24689);
nor UO_918 (O_918,N_22779,N_21911);
and UO_919 (O_919,N_24993,N_24759);
nand UO_920 (O_920,N_24607,N_22568);
nor UO_921 (O_921,N_20598,N_24764);
and UO_922 (O_922,N_21544,N_24444);
and UO_923 (O_923,N_21129,N_24395);
nor UO_924 (O_924,N_22878,N_23462);
xnor UO_925 (O_925,N_24353,N_21076);
nor UO_926 (O_926,N_22684,N_23361);
nor UO_927 (O_927,N_20381,N_21211);
nor UO_928 (O_928,N_23584,N_21902);
or UO_929 (O_929,N_22309,N_24862);
nand UO_930 (O_930,N_21644,N_22231);
and UO_931 (O_931,N_21665,N_21766);
or UO_932 (O_932,N_20089,N_23336);
nor UO_933 (O_933,N_21817,N_24379);
and UO_934 (O_934,N_22085,N_24625);
or UO_935 (O_935,N_22564,N_20935);
and UO_936 (O_936,N_20646,N_20248);
and UO_937 (O_937,N_20157,N_24214);
nor UO_938 (O_938,N_23348,N_24975);
and UO_939 (O_939,N_24885,N_20806);
nand UO_940 (O_940,N_23318,N_22445);
or UO_941 (O_941,N_24752,N_21306);
nand UO_942 (O_942,N_23182,N_23701);
nand UO_943 (O_943,N_21838,N_21006);
nor UO_944 (O_944,N_22715,N_20135);
nor UO_945 (O_945,N_22476,N_21314);
and UO_946 (O_946,N_20625,N_24909);
or UO_947 (O_947,N_23948,N_20084);
nand UO_948 (O_948,N_22939,N_20503);
nor UO_949 (O_949,N_23050,N_24661);
nand UO_950 (O_950,N_22986,N_20830);
or UO_951 (O_951,N_23617,N_21277);
nor UO_952 (O_952,N_24729,N_23508);
or UO_953 (O_953,N_23301,N_20169);
nor UO_954 (O_954,N_23725,N_23066);
or UO_955 (O_955,N_23806,N_24674);
or UO_956 (O_956,N_21898,N_24218);
or UO_957 (O_957,N_20952,N_20451);
nand UO_958 (O_958,N_22924,N_22913);
nor UO_959 (O_959,N_23357,N_21629);
or UO_960 (O_960,N_23142,N_22251);
nor UO_961 (O_961,N_23519,N_24911);
or UO_962 (O_962,N_23264,N_23973);
nor UO_963 (O_963,N_20162,N_23265);
or UO_964 (O_964,N_23982,N_21869);
or UO_965 (O_965,N_22406,N_22452);
or UO_966 (O_966,N_21033,N_21517);
and UO_967 (O_967,N_20258,N_24031);
nor UO_968 (O_968,N_21955,N_22190);
and UO_969 (O_969,N_24292,N_22838);
and UO_970 (O_970,N_21600,N_21018);
nand UO_971 (O_971,N_23493,N_22057);
nand UO_972 (O_972,N_20871,N_21154);
nand UO_973 (O_973,N_22265,N_20044);
nor UO_974 (O_974,N_24637,N_20452);
nand UO_975 (O_975,N_20443,N_21371);
nand UO_976 (O_976,N_23427,N_24619);
nor UO_977 (O_977,N_23145,N_22774);
or UO_978 (O_978,N_23686,N_23785);
and UO_979 (O_979,N_20652,N_21605);
nand UO_980 (O_980,N_24225,N_22964);
nand UO_981 (O_981,N_23008,N_21606);
nor UO_982 (O_982,N_21935,N_22627);
nor UO_983 (O_983,N_20878,N_22911);
or UO_984 (O_984,N_22656,N_21245);
nor UO_985 (O_985,N_23966,N_21233);
or UO_986 (O_986,N_24082,N_23917);
xor UO_987 (O_987,N_21528,N_20954);
nand UO_988 (O_988,N_23220,N_20927);
nand UO_989 (O_989,N_24173,N_24016);
and UO_990 (O_990,N_21592,N_22872);
and UO_991 (O_991,N_20392,N_21224);
nand UO_992 (O_992,N_22768,N_22468);
or UO_993 (O_993,N_24277,N_21281);
nand UO_994 (O_994,N_21264,N_23783);
or UO_995 (O_995,N_23840,N_22438);
nor UO_996 (O_996,N_20803,N_20278);
nand UO_997 (O_997,N_24768,N_24582);
nand UO_998 (O_998,N_24916,N_23158);
or UO_999 (O_999,N_22246,N_20470);
nand UO_1000 (O_1000,N_24030,N_20616);
nor UO_1001 (O_1001,N_20906,N_24118);
nor UO_1002 (O_1002,N_23834,N_21552);
nor UO_1003 (O_1003,N_20776,N_22173);
nand UO_1004 (O_1004,N_23047,N_23848);
nor UO_1005 (O_1005,N_20047,N_21296);
nand UO_1006 (O_1006,N_24954,N_23943);
and UO_1007 (O_1007,N_21633,N_23620);
and UO_1008 (O_1008,N_23097,N_22021);
nand UO_1009 (O_1009,N_21673,N_21151);
or UO_1010 (O_1010,N_22214,N_23951);
or UO_1011 (O_1011,N_21857,N_23589);
and UO_1012 (O_1012,N_24406,N_20374);
nand UO_1013 (O_1013,N_22866,N_20151);
nand UO_1014 (O_1014,N_24992,N_20036);
or UO_1015 (O_1015,N_22177,N_23103);
nand UO_1016 (O_1016,N_20450,N_23689);
nand UO_1017 (O_1017,N_23341,N_24778);
nand UO_1018 (O_1018,N_20137,N_23698);
nand UO_1019 (O_1019,N_21584,N_20058);
nor UO_1020 (O_1020,N_22886,N_22252);
nand UO_1021 (O_1021,N_22685,N_24855);
nand UO_1022 (O_1022,N_23148,N_21723);
and UO_1023 (O_1023,N_23476,N_23673);
nor UO_1024 (O_1024,N_22949,N_24753);
nand UO_1025 (O_1025,N_23736,N_21506);
or UO_1026 (O_1026,N_20745,N_22147);
or UO_1027 (O_1027,N_22540,N_21485);
or UO_1028 (O_1028,N_24463,N_24081);
nand UO_1029 (O_1029,N_23655,N_21979);
or UO_1030 (O_1030,N_22357,N_23423);
nand UO_1031 (O_1031,N_20003,N_20692);
or UO_1032 (O_1032,N_20801,N_24960);
nand UO_1033 (O_1033,N_23750,N_24518);
and UO_1034 (O_1034,N_20980,N_20380);
or UO_1035 (O_1035,N_21262,N_23255);
and UO_1036 (O_1036,N_22358,N_21668);
or UO_1037 (O_1037,N_21343,N_23129);
or UO_1038 (O_1038,N_22332,N_20077);
nor UO_1039 (O_1039,N_21044,N_21837);
or UO_1040 (O_1040,N_21079,N_24061);
nand UO_1041 (O_1041,N_23578,N_22129);
and UO_1042 (O_1042,N_20673,N_23690);
and UO_1043 (O_1043,N_24229,N_23053);
xor UO_1044 (O_1044,N_20456,N_23827);
and UO_1045 (O_1045,N_23084,N_21712);
and UO_1046 (O_1046,N_24127,N_20018);
nand UO_1047 (O_1047,N_22189,N_22072);
or UO_1048 (O_1048,N_24587,N_22697);
nand UO_1049 (O_1049,N_24652,N_24123);
and UO_1050 (O_1050,N_20017,N_22819);
nor UO_1051 (O_1051,N_23177,N_20685);
nor UO_1052 (O_1052,N_20195,N_24508);
nand UO_1053 (O_1053,N_24863,N_21287);
xnor UO_1054 (O_1054,N_23273,N_21789);
or UO_1055 (O_1055,N_22451,N_22346);
or UO_1056 (O_1056,N_21844,N_21128);
nor UO_1057 (O_1057,N_21966,N_20292);
or UO_1058 (O_1058,N_22240,N_24713);
nor UO_1059 (O_1059,N_23947,N_22449);
or UO_1060 (O_1060,N_24939,N_23202);
or UO_1061 (O_1061,N_24014,N_24720);
nand UO_1062 (O_1062,N_21553,N_22441);
or UO_1063 (O_1063,N_20504,N_23413);
nor UO_1064 (O_1064,N_23464,N_22647);
nor UO_1065 (O_1065,N_21337,N_23911);
and UO_1066 (O_1066,N_22987,N_23500);
and UO_1067 (O_1067,N_22047,N_24438);
or UO_1068 (O_1068,N_21782,N_23560);
nand UO_1069 (O_1069,N_22493,N_20740);
or UO_1070 (O_1070,N_23450,N_22488);
nand UO_1071 (O_1071,N_20814,N_21880);
nor UO_1072 (O_1072,N_20948,N_20295);
nand UO_1073 (O_1073,N_24962,N_23807);
or UO_1074 (O_1074,N_23446,N_21137);
nor UO_1075 (O_1075,N_20120,N_24160);
nor UO_1076 (O_1076,N_24934,N_23196);
or UO_1077 (O_1077,N_21459,N_22176);
and UO_1078 (O_1078,N_22694,N_22663);
nor UO_1079 (O_1079,N_22039,N_21798);
nand UO_1080 (O_1080,N_24046,N_23025);
nor UO_1081 (O_1081,N_21452,N_21157);
and UO_1082 (O_1082,N_20824,N_24741);
and UO_1083 (O_1083,N_20724,N_21945);
and UO_1084 (O_1084,N_20391,N_24519);
nand UO_1085 (O_1085,N_20405,N_23507);
and UO_1086 (O_1086,N_22380,N_20975);
nand UO_1087 (O_1087,N_21747,N_22877);
nor UO_1088 (O_1088,N_24009,N_24590);
nand UO_1089 (O_1089,N_22765,N_20215);
and UO_1090 (O_1090,N_20774,N_21510);
or UO_1091 (O_1091,N_23596,N_23684);
or UO_1092 (O_1092,N_23079,N_22623);
nand UO_1093 (O_1093,N_22290,N_22216);
or UO_1094 (O_1094,N_22848,N_22132);
nor UO_1095 (O_1095,N_20985,N_21263);
nor UO_1096 (O_1096,N_24347,N_22633);
nor UO_1097 (O_1097,N_22591,N_23607);
nand UO_1098 (O_1098,N_21476,N_24566);
xor UO_1099 (O_1099,N_20837,N_24643);
nor UO_1100 (O_1100,N_23749,N_22796);
and UO_1101 (O_1101,N_22462,N_22091);
and UO_1102 (O_1102,N_24476,N_21468);
nor UO_1103 (O_1103,N_23482,N_20139);
nor UO_1104 (O_1104,N_23152,N_23358);
and UO_1105 (O_1105,N_24259,N_24439);
or UO_1106 (O_1106,N_23828,N_20769);
or UO_1107 (O_1107,N_22912,N_24231);
nor UO_1108 (O_1108,N_24982,N_24193);
and UO_1109 (O_1109,N_24857,N_21479);
nand UO_1110 (O_1110,N_22243,N_24311);
or UO_1111 (O_1111,N_24677,N_20640);
nand UO_1112 (O_1112,N_24060,N_21990);
nor UO_1113 (O_1113,N_21839,N_24168);
nand UO_1114 (O_1114,N_20545,N_22651);
nor UO_1115 (O_1115,N_21858,N_20734);
nor UO_1116 (O_1116,N_21052,N_22114);
and UO_1117 (O_1117,N_24500,N_22769);
nand UO_1118 (O_1118,N_23509,N_23670);
xnor UO_1119 (O_1119,N_24723,N_21380);
and UO_1120 (O_1120,N_20041,N_22547);
nand UO_1121 (O_1121,N_21874,N_20185);
nor UO_1122 (O_1122,N_21501,N_23494);
nor UO_1123 (O_1123,N_22696,N_22689);
nor UO_1124 (O_1124,N_23697,N_23116);
nand UO_1125 (O_1125,N_23751,N_20660);
nand UO_1126 (O_1126,N_24136,N_23561);
nand UO_1127 (O_1127,N_21639,N_22921);
xor UO_1128 (O_1128,N_20641,N_20094);
and UO_1129 (O_1129,N_22466,N_22084);
or UO_1130 (O_1130,N_21512,N_24813);
nor UO_1131 (O_1131,N_23492,N_24692);
nand UO_1132 (O_1132,N_22097,N_20065);
or UO_1133 (O_1133,N_20981,N_23364);
and UO_1134 (O_1134,N_20910,N_24322);
nor UO_1135 (O_1135,N_23046,N_21713);
nand UO_1136 (O_1136,N_24419,N_24263);
or UO_1137 (O_1137,N_20914,N_24169);
nor UO_1138 (O_1138,N_21374,N_20480);
nand UO_1139 (O_1139,N_22377,N_24699);
nor UO_1140 (O_1140,N_23110,N_20771);
and UO_1141 (O_1141,N_20739,N_20968);
and UO_1142 (O_1142,N_20650,N_24492);
nor UO_1143 (O_1143,N_21850,N_21936);
and UO_1144 (O_1144,N_20183,N_23132);
or UO_1145 (O_1145,N_22969,N_20209);
nand UO_1146 (O_1146,N_24843,N_22772);
nor UO_1147 (O_1147,N_24047,N_20353);
nor UO_1148 (O_1148,N_20045,N_20002);
nor UO_1149 (O_1149,N_22064,N_22413);
nand UO_1150 (O_1150,N_23516,N_22959);
and UO_1151 (O_1151,N_20710,N_22481);
nand UO_1152 (O_1152,N_20286,N_21919);
and UO_1153 (O_1153,N_21221,N_20961);
or UO_1154 (O_1154,N_23082,N_24433);
nor UO_1155 (O_1155,N_23133,N_21755);
or UO_1156 (O_1156,N_22242,N_21993);
or UO_1157 (O_1157,N_23198,N_20885);
and UO_1158 (O_1158,N_21241,N_23206);
or UO_1159 (O_1159,N_22712,N_21147);
and UO_1160 (O_1160,N_24348,N_20250);
and UO_1161 (O_1161,N_23978,N_23184);
and UO_1162 (O_1162,N_20291,N_24318);
and UO_1163 (O_1163,N_21906,N_23010);
nand UO_1164 (O_1164,N_22750,N_22312);
nor UO_1165 (O_1165,N_20272,N_24481);
xor UO_1166 (O_1166,N_21895,N_22711);
or UO_1167 (O_1167,N_21565,N_21095);
nand UO_1168 (O_1168,N_21809,N_20006);
or UO_1169 (O_1169,N_23254,N_20186);
nand UO_1170 (O_1170,N_20951,N_24835);
xor UO_1171 (O_1171,N_22029,N_24715);
and UO_1172 (O_1172,N_22551,N_22404);
nor UO_1173 (O_1173,N_22639,N_24380);
and UO_1174 (O_1174,N_21983,N_23419);
and UO_1175 (O_1175,N_24235,N_21915);
nand UO_1176 (O_1176,N_20725,N_21302);
and UO_1177 (O_1177,N_21852,N_24794);
and UO_1178 (O_1178,N_22616,N_24870);
nand UO_1179 (O_1179,N_23456,N_20967);
nor UO_1180 (O_1180,N_22015,N_21951);
nor UO_1181 (O_1181,N_24586,N_23481);
nand UO_1182 (O_1182,N_24350,N_23913);
and UO_1183 (O_1183,N_21115,N_23772);
nand UO_1184 (O_1184,N_23957,N_22378);
xor UO_1185 (O_1185,N_24973,N_24040);
or UO_1186 (O_1186,N_22408,N_24538);
nand UO_1187 (O_1187,N_24337,N_24948);
nand UO_1188 (O_1188,N_21525,N_20279);
or UO_1189 (O_1189,N_24408,N_20620);
or UO_1190 (O_1190,N_23345,N_23111);
nand UO_1191 (O_1191,N_22491,N_23344);
nand UO_1192 (O_1192,N_22710,N_21615);
or UO_1193 (O_1193,N_23979,N_22781);
nand UO_1194 (O_1194,N_21655,N_20701);
or UO_1195 (O_1195,N_22326,N_23013);
and UO_1196 (O_1196,N_23581,N_23165);
and UO_1197 (O_1197,N_24543,N_22882);
nor UO_1198 (O_1198,N_23221,N_21625);
nand UO_1199 (O_1199,N_21335,N_20025);
and UO_1200 (O_1200,N_24328,N_22080);
nand UO_1201 (O_1201,N_23676,N_23384);
nand UO_1202 (O_1202,N_24679,N_21388);
nor UO_1203 (O_1203,N_21815,N_22238);
nand UO_1204 (O_1204,N_23810,N_22464);
and UO_1205 (O_1205,N_23909,N_23590);
or UO_1206 (O_1206,N_23135,N_23682);
and UO_1207 (O_1207,N_24662,N_21761);
xnor UO_1208 (O_1208,N_23143,N_21642);
and UO_1209 (O_1209,N_20173,N_23455);
nor UO_1210 (O_1210,N_23296,N_22807);
and UO_1211 (O_1211,N_24124,N_24296);
and UO_1212 (O_1212,N_23478,N_21813);
nor UO_1213 (O_1213,N_20936,N_23674);
xor UO_1214 (O_1214,N_24331,N_21408);
and UO_1215 (O_1215,N_24858,N_24418);
or UO_1216 (O_1216,N_20982,N_20441);
nor UO_1217 (O_1217,N_21722,N_24211);
nand UO_1218 (O_1218,N_20174,N_20253);
and UO_1219 (O_1219,N_20081,N_22558);
nand UO_1220 (O_1220,N_23139,N_23011);
or UO_1221 (O_1221,N_22981,N_22748);
nor UO_1222 (O_1222,N_22041,N_20707);
nand UO_1223 (O_1223,N_23441,N_22055);
and UO_1224 (O_1224,N_22374,N_24766);
and UO_1225 (O_1225,N_22581,N_21870);
nand UO_1226 (O_1226,N_23113,N_24771);
nor UO_1227 (O_1227,N_22075,N_24412);
nand UO_1228 (O_1228,N_20731,N_21734);
nor UO_1229 (O_1229,N_22946,N_23733);
and UO_1230 (O_1230,N_24254,N_20606);
nor UO_1231 (O_1231,N_20525,N_23411);
nand UO_1232 (O_1232,N_20457,N_23349);
nor UO_1233 (O_1233,N_22903,N_23665);
nand UO_1234 (O_1234,N_24547,N_21368);
nor UO_1235 (O_1235,N_21675,N_22675);
nor UO_1236 (O_1236,N_20867,N_22174);
nor UO_1237 (O_1237,N_21378,N_24215);
or UO_1238 (O_1238,N_23115,N_22222);
or UO_1239 (O_1239,N_22062,N_20911);
nand UO_1240 (O_1240,N_21750,N_22747);
nor UO_1241 (O_1241,N_21067,N_24367);
or UO_1242 (O_1242,N_23477,N_22456);
or UO_1243 (O_1243,N_20636,N_23870);
or UO_1244 (O_1244,N_23833,N_20887);
nor UO_1245 (O_1245,N_20244,N_24913);
and UO_1246 (O_1246,N_20252,N_24927);
nand UO_1247 (O_1247,N_23280,N_21595);
and UO_1248 (O_1248,N_22520,N_24540);
nand UO_1249 (O_1249,N_23219,N_20716);
nand UO_1250 (O_1250,N_22679,N_20763);
xnor UO_1251 (O_1251,N_23058,N_21329);
nand UO_1252 (O_1252,N_24573,N_20499);
and UO_1253 (O_1253,N_23269,N_22856);
nand UO_1254 (O_1254,N_21072,N_20681);
nand UO_1255 (O_1255,N_22133,N_20141);
xor UO_1256 (O_1256,N_24891,N_22022);
and UO_1257 (O_1257,N_22671,N_21757);
nor UO_1258 (O_1258,N_24987,N_23908);
or UO_1259 (O_1259,N_23339,N_22083);
and UO_1260 (O_1260,N_20540,N_20546);
nand UO_1261 (O_1261,N_24549,N_23616);
or UO_1262 (O_1262,N_21316,N_22786);
nor UO_1263 (O_1263,N_23835,N_21738);
and UO_1264 (O_1264,N_21941,N_24793);
and UO_1265 (O_1265,N_24317,N_24743);
nand UO_1266 (O_1266,N_24883,N_22101);
and UO_1267 (O_1267,N_22888,N_23078);
nand UO_1268 (O_1268,N_23658,N_24086);
nand UO_1269 (O_1269,N_23071,N_20582);
and UO_1270 (O_1270,N_20102,N_22523);
nand UO_1271 (O_1271,N_21819,N_22764);
or UO_1272 (O_1272,N_21507,N_20713);
or UO_1273 (O_1273,N_20356,N_24685);
nand UO_1274 (O_1274,N_20688,N_21199);
xor UO_1275 (O_1275,N_21195,N_21754);
and UO_1276 (O_1276,N_22037,N_20460);
nand UO_1277 (O_1277,N_23933,N_22968);
or UO_1278 (O_1278,N_22545,N_23669);
xor UO_1279 (O_1279,N_24791,N_23138);
or UO_1280 (O_1280,N_22543,N_21863);
or UO_1281 (O_1281,N_22511,N_23723);
nor UO_1282 (O_1282,N_20016,N_24224);
nand UO_1283 (O_1283,N_22755,N_23638);
nand UO_1284 (O_1284,N_20889,N_20584);
and UO_1285 (O_1285,N_24817,N_24302);
nor UO_1286 (O_1286,N_20697,N_22308);
and UO_1287 (O_1287,N_24468,N_20168);
and UO_1288 (O_1288,N_21604,N_20690);
nand UO_1289 (O_1289,N_20305,N_22974);
nor UO_1290 (O_1290,N_22507,N_24572);
or UO_1291 (O_1291,N_23051,N_23597);
and UO_1292 (O_1292,N_21198,N_21258);
and UO_1293 (O_1293,N_20866,N_20790);
and UO_1294 (O_1294,N_20316,N_24335);
and UO_1295 (O_1295,N_22457,N_22012);
or UO_1296 (O_1296,N_24717,N_24076);
or UO_1297 (O_1297,N_20176,N_24152);
nand UO_1298 (O_1298,N_21204,N_23888);
and UO_1299 (O_1299,N_24933,N_21934);
nor UO_1300 (O_1300,N_20805,N_20001);
and UO_1301 (O_1301,N_20479,N_20592);
or UO_1302 (O_1302,N_23297,N_21415);
nor UO_1303 (O_1303,N_21714,N_22599);
or UO_1304 (O_1304,N_24085,N_23242);
nor UO_1305 (O_1305,N_22031,N_24839);
nand UO_1306 (O_1306,N_20547,N_21904);
nor UO_1307 (O_1307,N_24114,N_23952);
or UO_1308 (O_1308,N_22215,N_22676);
nor UO_1309 (O_1309,N_22237,N_24239);
or UO_1310 (O_1310,N_23991,N_22333);
nand UO_1311 (O_1311,N_21339,N_20825);
or UO_1312 (O_1312,N_23855,N_21997);
nand UO_1313 (O_1313,N_24023,N_23171);
or UO_1314 (O_1314,N_21998,N_20880);
nand UO_1315 (O_1315,N_20290,N_22589);
or UO_1316 (O_1316,N_23510,N_20384);
nand UO_1317 (O_1317,N_22854,N_24795);
and UO_1318 (O_1318,N_21138,N_22546);
and UO_1319 (O_1319,N_22614,N_20074);
or UO_1320 (O_1320,N_24097,N_20069);
nand UO_1321 (O_1321,N_23405,N_20794);
or UO_1322 (O_1322,N_22840,N_21170);
nand UO_1323 (O_1323,N_23938,N_21913);
and UO_1324 (O_1324,N_20190,N_22957);
nor UO_1325 (O_1325,N_23307,N_24667);
nand UO_1326 (O_1326,N_22204,N_24952);
nor UO_1327 (O_1327,N_24802,N_21118);
xnor UO_1328 (O_1328,N_22403,N_24290);
or UO_1329 (O_1329,N_23668,N_21818);
and UO_1330 (O_1330,N_20829,N_20158);
nand UO_1331 (O_1331,N_23438,N_20395);
and UO_1332 (O_1332,N_20928,N_22004);
nand UO_1333 (O_1333,N_22268,N_22026);
and UO_1334 (O_1334,N_22361,N_24648);
or UO_1335 (O_1335,N_24560,N_21389);
nor UO_1336 (O_1336,N_21446,N_21790);
or UO_1337 (O_1337,N_22112,N_20040);
or UO_1338 (O_1338,N_20448,N_20146);
nand UO_1339 (O_1339,N_21030,N_20332);
or UO_1340 (O_1340,N_20567,N_23057);
and UO_1341 (O_1341,N_23800,N_23123);
and UO_1342 (O_1342,N_20372,N_23306);
nand UO_1343 (O_1343,N_24775,N_24955);
nand UO_1344 (O_1344,N_23014,N_20857);
and UO_1345 (O_1345,N_21899,N_21059);
or UO_1346 (O_1346,N_21422,N_22425);
or UO_1347 (O_1347,N_24050,N_20061);
or UO_1348 (O_1348,N_21435,N_20096);
nor UO_1349 (O_1349,N_22943,N_20919);
and UO_1350 (O_1350,N_20608,N_23465);
and UO_1351 (O_1351,N_21053,N_23514);
nand UO_1352 (O_1352,N_22604,N_24460);
nor UO_1353 (O_1353,N_20247,N_21260);
nand UO_1354 (O_1354,N_22344,N_21744);
and UO_1355 (O_1355,N_22630,N_20585);
and UO_1356 (O_1356,N_20839,N_22071);
nor UO_1357 (O_1357,N_24964,N_20573);
nor UO_1358 (O_1358,N_20770,N_21492);
or UO_1359 (O_1359,N_23650,N_22304);
nand UO_1360 (O_1360,N_23805,N_21795);
and UO_1361 (O_1361,N_20845,N_21859);
nand UO_1362 (O_1362,N_21865,N_22565);
or UO_1363 (O_1363,N_20439,N_24455);
nand UO_1364 (O_1364,N_23385,N_20070);
or UO_1365 (O_1365,N_21248,N_20210);
nand UO_1366 (O_1366,N_22009,N_22396);
nand UO_1367 (O_1367,N_20199,N_24153);
or UO_1368 (O_1368,N_20572,N_23426);
nand UO_1369 (O_1369,N_21740,N_20578);
and UO_1370 (O_1370,N_20738,N_22894);
nor UO_1371 (O_1371,N_21588,N_20329);
and UO_1372 (O_1372,N_20079,N_20861);
and UO_1373 (O_1373,N_20394,N_23902);
or UO_1374 (O_1374,N_20156,N_23369);
nor UO_1375 (O_1375,N_22960,N_24546);
nand UO_1376 (O_1376,N_24707,N_21495);
xnor UO_1377 (O_1377,N_24761,N_21694);
nand UO_1378 (O_1378,N_24575,N_22771);
nand UO_1379 (O_1379,N_24830,N_21417);
nor UO_1380 (O_1380,N_23971,N_23304);
and UO_1381 (O_1381,N_24421,N_20657);
and UO_1382 (O_1382,N_23252,N_21947);
xnor UO_1383 (O_1383,N_24356,N_24338);
or UO_1384 (O_1384,N_22105,N_21149);
nand UO_1385 (O_1385,N_20978,N_23624);
nand UO_1386 (O_1386,N_21101,N_23457);
nand UO_1387 (O_1387,N_23124,N_22965);
nand UO_1388 (O_1388,N_22782,N_23559);
nand UO_1389 (O_1389,N_24923,N_22329);
nand UO_1390 (O_1390,N_23140,N_20029);
xnor UO_1391 (O_1391,N_23317,N_23032);
or UO_1392 (O_1392,N_22678,N_21178);
nor UO_1393 (O_1393,N_21162,N_23108);
nor UO_1394 (O_1394,N_21220,N_24754);
nor UO_1395 (O_1395,N_20533,N_20126);
nand UO_1396 (O_1396,N_20851,N_24313);
nand UO_1397 (O_1397,N_22284,N_21830);
nand UO_1398 (O_1398,N_20717,N_24762);
nor UO_1399 (O_1399,N_20850,N_23729);
nand UO_1400 (O_1400,N_20223,N_22487);
nand UO_1401 (O_1401,N_24694,N_20526);
or UO_1402 (O_1402,N_24357,N_20568);
nand UO_1403 (O_1403,N_20359,N_20313);
nor UO_1404 (O_1404,N_23872,N_23763);
or UO_1405 (O_1405,N_21901,N_23491);
and UO_1406 (O_1406,N_23488,N_21251);
or UO_1407 (O_1407,N_23983,N_20064);
and UO_1408 (O_1408,N_20170,N_23771);
or UO_1409 (O_1409,N_24083,N_21758);
and UO_1410 (O_1410,N_22260,N_22381);
nand UO_1411 (O_1411,N_22137,N_24868);
nor UO_1412 (O_1412,N_21414,N_24090);
nor UO_1413 (O_1413,N_23467,N_20807);
and UO_1414 (O_1414,N_24965,N_23141);
and UO_1415 (O_1415,N_20698,N_22050);
nand UO_1416 (O_1416,N_21488,N_23788);
and UO_1417 (O_1417,N_23204,N_23752);
or UO_1418 (O_1418,N_23292,N_21480);
and UO_1419 (O_1419,N_24499,N_22896);
and UO_1420 (O_1420,N_21546,N_20907);
or UO_1421 (O_1421,N_23062,N_21918);
or UO_1422 (O_1422,N_24698,N_23996);
and UO_1423 (O_1423,N_23475,N_20812);
nand UO_1424 (O_1424,N_20844,N_20203);
or UO_1425 (O_1425,N_20144,N_24055);
or UO_1426 (O_1426,N_24291,N_22612);
and UO_1427 (O_1427,N_24282,N_21359);
nor UO_1428 (O_1428,N_22254,N_24584);
nand UO_1429 (O_1429,N_24098,N_24985);
and UO_1430 (O_1430,N_21821,N_24944);
and UO_1431 (O_1431,N_22152,N_20737);
nor UO_1432 (O_1432,N_21404,N_23173);
nor UO_1433 (O_1433,N_20996,N_24222);
nand UO_1434 (O_1434,N_24245,N_22082);
and UO_1435 (O_1435,N_24101,N_23819);
nor UO_1436 (O_1436,N_23393,N_22842);
nor UO_1437 (O_1437,N_22120,N_24232);
or UO_1438 (O_1438,N_20575,N_21168);
nor UO_1439 (O_1439,N_21029,N_20709);
nand UO_1440 (O_1440,N_24551,N_23885);
nand UO_1441 (O_1441,N_23568,N_20864);
nand UO_1442 (O_1442,N_22917,N_21599);
nor UO_1443 (O_1443,N_20561,N_24221);
nor UO_1444 (O_1444,N_23172,N_23614);
and UO_1445 (O_1445,N_23603,N_23781);
nor UO_1446 (O_1446,N_20528,N_20306);
or UO_1447 (O_1447,N_24486,N_20583);
and UO_1448 (O_1448,N_23527,N_21810);
xor UO_1449 (O_1449,N_23970,N_24012);
nor UO_1450 (O_1450,N_22061,N_22988);
and UO_1451 (O_1451,N_21416,N_20501);
and UO_1452 (O_1452,N_20321,N_20138);
nor UO_1453 (O_1453,N_21200,N_20109);
nand UO_1454 (O_1454,N_21164,N_24529);
and UO_1455 (O_1455,N_24473,N_21845);
nor UO_1456 (O_1456,N_21942,N_20828);
and UO_1457 (O_1457,N_24442,N_21228);
xor UO_1458 (O_1458,N_23236,N_22657);
and UO_1459 (O_1459,N_20979,N_23466);
and UO_1460 (O_1460,N_22621,N_24703);
or UO_1461 (O_1461,N_21235,N_22862);
xnor UO_1462 (O_1462,N_22863,N_23227);
and UO_1463 (O_1463,N_24340,N_24005);
and UO_1464 (O_1464,N_20437,N_21063);
or UO_1465 (O_1465,N_24404,N_24653);
nor UO_1466 (O_1466,N_23421,N_22655);
or UO_1467 (O_1467,N_23681,N_20627);
or UO_1468 (O_1468,N_24339,N_23041);
nor UO_1469 (O_1469,N_23028,N_23356);
nor UO_1470 (O_1470,N_24069,N_20020);
and UO_1471 (O_1471,N_24185,N_24077);
and UO_1472 (O_1472,N_21487,N_21842);
or UO_1473 (O_1473,N_20875,N_20367);
nor UO_1474 (O_1474,N_21514,N_22699);
nor UO_1475 (O_1475,N_20474,N_23223);
or UO_1476 (O_1476,N_22020,N_20520);
and UO_1477 (O_1477,N_21548,N_22058);
nor UO_1478 (O_1478,N_20113,N_22371);
or UO_1479 (O_1479,N_20591,N_20502);
nor UO_1480 (O_1480,N_22744,N_20011);
or UO_1481 (O_1481,N_21678,N_21958);
and UO_1482 (O_1482,N_22005,N_23582);
nand UO_1483 (O_1483,N_20855,N_22952);
or UO_1484 (O_1484,N_23081,N_21110);
nor UO_1485 (O_1485,N_22904,N_21184);
nor UO_1486 (O_1486,N_21247,N_20184);
or UO_1487 (O_1487,N_24553,N_23288);
or UO_1488 (O_1488,N_23631,N_20842);
or UO_1489 (O_1489,N_21811,N_24822);
nand UO_1490 (O_1490,N_22832,N_21434);
and UO_1491 (O_1491,N_24137,N_24915);
nand UO_1492 (O_1492,N_23764,N_21926);
or UO_1493 (O_1493,N_24471,N_23880);
nor UO_1494 (O_1494,N_22978,N_23350);
xnor UO_1495 (O_1495,N_22890,N_24847);
nor UO_1496 (O_1496,N_24036,N_22539);
or UO_1497 (O_1497,N_20683,N_24502);
and UO_1498 (O_1498,N_22317,N_21083);
nand UO_1499 (O_1499,N_24836,N_22736);
xor UO_1500 (O_1500,N_24472,N_24899);
and UO_1501 (O_1501,N_21005,N_23667);
or UO_1502 (O_1502,N_20019,N_24308);
or UO_1503 (O_1503,N_20413,N_21824);
nor UO_1504 (O_1504,N_21041,N_21166);
and UO_1505 (O_1505,N_22171,N_22756);
xor UO_1506 (O_1506,N_21103,N_21443);
nor UO_1507 (O_1507,N_21494,N_21703);
nor UO_1508 (O_1508,N_22283,N_24260);
nor UO_1509 (O_1509,N_23376,N_20991);
or UO_1510 (O_1510,N_24631,N_23661);
and UO_1511 (O_1511,N_21171,N_22167);
and UO_1512 (O_1512,N_20009,N_23610);
or UO_1513 (O_1513,N_23070,N_20325);
nor UO_1514 (O_1514,N_20500,N_21640);
nand UO_1515 (O_1515,N_24971,N_23045);
or UO_1516 (O_1516,N_22467,N_20355);
and UO_1517 (O_1517,N_23226,N_24838);
and UO_1518 (O_1518,N_22868,N_24869);
and UO_1519 (O_1519,N_21442,N_21564);
or UO_1520 (O_1520,N_20164,N_22813);
and UO_1521 (O_1521,N_21971,N_23879);
xor UO_1522 (O_1522,N_22668,N_23844);
nor UO_1523 (O_1523,N_20121,N_22195);
nor UO_1524 (O_1524,N_20753,N_22503);
nand UO_1525 (O_1525,N_23262,N_22841);
nand UO_1526 (O_1526,N_21635,N_21742);
nand UO_1527 (O_1527,N_22561,N_20957);
or UO_1528 (O_1528,N_22313,N_20858);
xnor UO_1529 (O_1529,N_21123,N_20728);
or UO_1530 (O_1530,N_21209,N_20442);
or UO_1531 (O_1531,N_24811,N_21534);
nor UO_1532 (O_1532,N_21003,N_24951);
nor UO_1533 (O_1533,N_21921,N_20945);
nand UO_1534 (O_1534,N_22472,N_23643);
and UO_1535 (O_1535,N_20983,N_24490);
nor UO_1536 (O_1536,N_23518,N_24018);
nor UO_1537 (O_1537,N_24541,N_22442);
nand UO_1538 (O_1538,N_23368,N_24333);
nor UO_1539 (O_1539,N_24015,N_22384);
nand UO_1540 (O_1540,N_23644,N_24845);
and UO_1541 (O_1541,N_20232,N_23406);
and UO_1542 (O_1542,N_24341,N_23534);
nor UO_1543 (O_1543,N_24111,N_20057);
nand UO_1544 (O_1544,N_21390,N_20111);
nor UO_1545 (O_1545,N_21047,N_21628);
nand UO_1546 (O_1546,N_23259,N_20265);
nor UO_1547 (O_1547,N_23294,N_24523);
or UO_1548 (O_1548,N_22855,N_23553);
nor UO_1549 (O_1549,N_22342,N_20090);
or UO_1550 (O_1550,N_22618,N_23711);
or UO_1551 (O_1551,N_23343,N_20749);
and UO_1552 (O_1552,N_20841,N_21952);
nand UO_1553 (O_1553,N_23905,N_21687);
and UO_1554 (O_1554,N_20795,N_22729);
or UO_1555 (O_1555,N_22328,N_20285);
or UO_1556 (O_1556,N_24640,N_22787);
or UO_1557 (O_1557,N_24450,N_24612);
nor UO_1558 (O_1558,N_24484,N_24522);
or UO_1559 (O_1559,N_20671,N_20410);
or UO_1560 (O_1560,N_20463,N_22563);
or UO_1561 (O_1561,N_23599,N_24666);
or UO_1562 (O_1562,N_21641,N_21916);
or UO_1563 (O_1563,N_22302,N_22664);
and UO_1564 (O_1564,N_20208,N_24996);
nand UO_1565 (O_1565,N_23291,N_23377);
nand UO_1566 (O_1566,N_20256,N_24735);
or UO_1567 (O_1567,N_20743,N_23289);
nor UO_1568 (O_1568,N_21759,N_24107);
nor UO_1569 (O_1569,N_24998,N_23160);
and UO_1570 (O_1570,N_23649,N_22143);
xnor UO_1571 (O_1571,N_23498,N_24826);
and UO_1572 (O_1572,N_21637,N_23585);
and UO_1573 (O_1573,N_24017,N_21340);
and UO_1574 (O_1574,N_22596,N_21730);
and UO_1575 (O_1575,N_21560,N_21907);
nand UO_1576 (O_1576,N_20649,N_21428);
nand UO_1577 (O_1577,N_20534,N_24495);
and UO_1578 (O_1578,N_21342,N_20339);
nand UO_1579 (O_1579,N_21763,N_23212);
and UO_1580 (O_1580,N_24212,N_20506);
and UO_1581 (O_1581,N_21814,N_21585);
or UO_1582 (O_1582,N_22399,N_22669);
or UO_1583 (O_1583,N_20963,N_21381);
and UO_1584 (O_1584,N_24200,N_20493);
nand UO_1585 (O_1585,N_24873,N_23815);
nor UO_1586 (O_1586,N_24928,N_21100);
or UO_1587 (O_1587,N_21327,N_21309);
nand UO_1588 (O_1588,N_20269,N_20099);
nor UO_1589 (O_1589,N_21447,N_20600);
nand UO_1590 (O_1590,N_22954,N_21345);
nor UO_1591 (O_1591,N_24722,N_21066);
and UO_1592 (O_1592,N_21784,N_20544);
nand UO_1593 (O_1593,N_21449,N_23085);
and UO_1594 (O_1594,N_22686,N_24684);
xnor UO_1595 (O_1595,N_24527,N_23418);
and UO_1596 (O_1596,N_21311,N_23903);
or UO_1597 (O_1597,N_22900,N_20884);
or UO_1598 (O_1598,N_21562,N_20114);
nand UO_1599 (O_1599,N_23106,N_24568);
and UO_1600 (O_1600,N_24453,N_24417);
and UO_1601 (O_1601,N_23372,N_20523);
or UO_1602 (O_1602,N_20361,N_24080);
or UO_1603 (O_1603,N_22814,N_24946);
nand UO_1604 (O_1604,N_23287,N_24850);
nor UO_1605 (O_1605,N_24399,N_21393);
or UO_1606 (O_1606,N_23120,N_24525);
and UO_1607 (O_1607,N_23235,N_21777);
nand UO_1608 (O_1608,N_22256,N_23359);
or UO_1609 (O_1609,N_24627,N_22110);
and UO_1610 (O_1610,N_23096,N_23128);
and UO_1611 (O_1611,N_20351,N_24686);
or UO_1612 (O_1612,N_22385,N_21994);
nand UO_1613 (O_1613,N_23314,N_22074);
nand UO_1614 (O_1614,N_22225,N_24819);
and UO_1615 (O_1615,N_22804,N_20242);
nor UO_1616 (O_1616,N_21197,N_22635);
nand UO_1617 (O_1617,N_22506,N_22822);
or UO_1618 (O_1618,N_21461,N_22353);
or UO_1619 (O_1619,N_23569,N_20477);
or UO_1620 (O_1620,N_24432,N_24329);
or UO_1621 (O_1621,N_22940,N_21054);
nand UO_1622 (O_1622,N_24226,N_24991);
nor UO_1623 (O_1623,N_20581,N_21188);
nor UO_1624 (O_1624,N_23490,N_22339);
nand UO_1625 (O_1625,N_22592,N_24170);
nor UO_1626 (O_1626,N_23059,N_22126);
or UO_1627 (O_1627,N_21091,N_22019);
and UO_1628 (O_1628,N_21269,N_20622);
nor UO_1629 (O_1629,N_24143,N_20119);
nor UO_1630 (O_1630,N_20675,N_24700);
or UO_1631 (O_1631,N_20287,N_20376);
and UO_1632 (O_1632,N_22733,N_20160);
and UO_1633 (O_1633,N_24301,N_20883);
xnor UO_1634 (O_1634,N_22864,N_20614);
nand UO_1635 (O_1635,N_23146,N_21638);
or UO_1636 (O_1636,N_21950,N_21482);
nand UO_1637 (O_1637,N_22992,N_20621);
nand UO_1638 (O_1638,N_20639,N_21791);
nor UO_1639 (O_1639,N_21325,N_24881);
nor UO_1640 (O_1640,N_20108,N_22389);
or UO_1641 (O_1641,N_22139,N_20892);
or UO_1642 (O_1642,N_24094,N_21363);
nand UO_1643 (O_1643,N_23532,N_21462);
and UO_1644 (O_1644,N_24407,N_23718);
nand UO_1645 (O_1645,N_22369,N_21890);
or UO_1646 (O_1646,N_24650,N_21491);
nor UO_1647 (O_1647,N_22262,N_20496);
or UO_1648 (O_1648,N_24025,N_23882);
and UO_1649 (O_1649,N_22714,N_22971);
or UO_1650 (O_1650,N_24034,N_20387);
and UO_1651 (O_1651,N_21308,N_22053);
and UO_1652 (O_1652,N_23992,N_23742);
or UO_1653 (O_1653,N_23170,N_22541);
or UO_1654 (O_1654,N_24295,N_20656);
nand UO_1655 (O_1655,N_21875,N_23695);
and UO_1656 (O_1656,N_21991,N_20997);
and UO_1657 (O_1657,N_21705,N_22718);
nand UO_1658 (O_1658,N_20904,N_23520);
nor UO_1659 (O_1659,N_23470,N_24249);
nand UO_1660 (O_1660,N_21317,N_21407);
and UO_1661 (O_1661,N_22938,N_20973);
and UO_1662 (O_1662,N_23461,N_21924);
or UO_1663 (O_1663,N_20105,N_23020);
and UO_1664 (O_1664,N_21725,N_22379);
and UO_1665 (O_1665,N_22089,N_23415);
nor UO_1666 (O_1666,N_21856,N_22625);
and UO_1667 (O_1667,N_24071,N_24556);
and UO_1668 (O_1668,N_20478,N_21733);
nand UO_1669 (O_1669,N_23546,N_21706);
nand UO_1670 (O_1670,N_20898,N_21286);
nand UO_1671 (O_1671,N_22522,N_20733);
nor UO_1672 (O_1672,N_24203,N_24592);
and UO_1673 (O_1673,N_23804,N_21444);
nor UO_1674 (O_1674,N_22722,N_21365);
and UO_1675 (O_1675,N_21131,N_20107);
nand UO_1676 (O_1676,N_22199,N_20539);
nand UO_1677 (O_1677,N_21659,N_24342);
and UO_1678 (O_1678,N_23707,N_22993);
and UO_1679 (O_1679,N_24672,N_24436);
and UO_1680 (O_1680,N_24820,N_24757);
nor UO_1681 (O_1681,N_20854,N_22322);
nand UO_1682 (O_1682,N_24139,N_20662);
or UO_1683 (O_1683,N_24393,N_24610);
or UO_1684 (O_1684,N_21545,N_22266);
nor UO_1685 (O_1685,N_22789,N_24906);
nand UO_1686 (O_1686,N_24171,N_24150);
nand UO_1687 (O_1687,N_20853,N_21634);
nor UO_1688 (O_1688,N_21419,N_24711);
nor UO_1689 (O_1689,N_22721,N_22160);
or UO_1690 (O_1690,N_24265,N_20615);
nand UO_1691 (O_1691,N_23030,N_21787);
or UO_1692 (O_1692,N_20718,N_21430);
nor UO_1693 (O_1693,N_23647,N_20354);
and UO_1694 (O_1694,N_22318,N_22386);
or UO_1695 (O_1695,N_23964,N_20766);
nand UO_1696 (O_1696,N_22424,N_24969);
nand UO_1697 (O_1697,N_22867,N_23960);
nand UO_1698 (O_1698,N_20758,N_21412);
and UO_1699 (O_1699,N_20396,N_22860);
or UO_1700 (O_1700,N_22982,N_20166);
nand UO_1701 (O_1701,N_21265,N_21303);
and UO_1702 (O_1702,N_23548,N_22926);
xnor UO_1703 (O_1703,N_22363,N_22638);
and UO_1704 (O_1704,N_23095,N_20596);
nand UO_1705 (O_1705,N_22461,N_20154);
xnor UO_1706 (O_1706,N_23503,N_20103);
or UO_1707 (O_1707,N_24279,N_22687);
xor UO_1708 (O_1708,N_24533,N_24750);
nor UO_1709 (O_1709,N_21344,N_22510);
nor UO_1710 (O_1710,N_20554,N_24589);
nand UO_1711 (O_1711,N_22259,N_22688);
nand UO_1712 (O_1712,N_23340,N_23362);
nand UO_1713 (O_1713,N_22294,N_20270);
nor UO_1714 (O_1714,N_23588,N_24064);
and UO_1715 (O_1715,N_21620,N_21580);
nor UO_1716 (O_1716,N_21524,N_21959);
nand UO_1717 (O_1717,N_21464,N_24892);
and UO_1718 (O_1718,N_20104,N_23342);
or UO_1719 (O_1719,N_20623,N_21405);
and UO_1720 (O_1720,N_22025,N_23021);
and UO_1721 (O_1721,N_23247,N_23642);
xor UO_1722 (O_1722,N_20229,N_23389);
and UO_1723 (O_1723,N_21292,N_20055);
nand UO_1724 (O_1724,N_24645,N_21649);
nor UO_1725 (O_1725,N_22429,N_21846);
nor UO_1726 (O_1726,N_24230,N_20052);
nor UO_1727 (O_1727,N_20895,N_23779);
or UO_1728 (O_1728,N_23439,N_24755);
and UO_1729 (O_1729,N_23329,N_22847);
and UO_1730 (O_1730,N_20931,N_20511);
xnor UO_1731 (O_1731,N_23155,N_20852);
and UO_1732 (O_1732,N_22839,N_24003);
nand UO_1733 (O_1733,N_24669,N_21775);
or UO_1734 (O_1734,N_21367,N_20411);
nand UO_1735 (O_1735,N_22979,N_22628);
and UO_1736 (O_1736,N_22258,N_22692);
nand UO_1737 (O_1737,N_21520,N_21621);
nand UO_1738 (O_1738,N_21324,N_23664);
and UO_1739 (O_1739,N_23839,N_23608);
or UO_1740 (O_1740,N_21674,N_24760);
nor UO_1741 (O_1741,N_23709,N_22144);
nor UO_1742 (O_1742,N_22674,N_22919);
and UO_1743 (O_1743,N_20872,N_24258);
or UO_1744 (O_1744,N_23162,N_21108);
or UO_1745 (O_1745,N_23654,N_23898);
and UO_1746 (O_1746,N_24056,N_20653);
nand UO_1747 (O_1747,N_23121,N_22573);
nand UO_1748 (O_1748,N_24601,N_22907);
and UO_1749 (O_1749,N_22994,N_22844);
nor UO_1750 (O_1750,N_22746,N_24895);
nand UO_1751 (O_1751,N_21282,N_22232);
nand UO_1752 (O_1752,N_20922,N_23713);
nand UO_1753 (O_1753,N_22607,N_23727);
nand UO_1754 (O_1754,N_22455,N_20324);
or UO_1755 (O_1755,N_20647,N_20167);
and UO_1756 (O_1756,N_24683,N_20434);
xnor UO_1757 (O_1757,N_21001,N_21776);
nor UO_1758 (O_1758,N_20761,N_20760);
nor UO_1759 (O_1759,N_21310,N_21176);
and UO_1760 (O_1760,N_24539,N_20008);
and UO_1761 (O_1761,N_24049,N_23501);
or UO_1762 (O_1762,N_22828,N_21581);
and UO_1763 (O_1763,N_23883,N_22829);
nor UO_1764 (O_1764,N_23330,N_24810);
nor UO_1765 (O_1765,N_24400,N_21596);
or UO_1766 (O_1766,N_24725,N_23594);
nand UO_1767 (O_1767,N_24389,N_20211);
nand UO_1768 (O_1768,N_22447,N_23812);
or UO_1769 (O_1769,N_20843,N_21767);
and UO_1770 (O_1770,N_20920,N_22496);
xnor UO_1771 (O_1771,N_20691,N_20564);
and UO_1772 (O_1772,N_23929,N_24010);
nor UO_1773 (O_1773,N_20037,N_20101);
nor UO_1774 (O_1774,N_24990,N_23271);
nor UO_1775 (O_1775,N_22121,N_22502);
or UO_1776 (O_1776,N_21960,N_20302);
nor UO_1777 (O_1777,N_23621,N_23144);
nor UO_1778 (O_1778,N_24781,N_23946);
or UO_1779 (O_1779,N_21903,N_20630);
nand UO_1780 (O_1780,N_21313,N_24605);
nor UO_1781 (O_1781,N_24510,N_21133);
nand UO_1782 (O_1782,N_23268,N_21683);
and UO_1783 (O_1783,N_23679,N_22337);
nor UO_1784 (O_1784,N_21786,N_21226);
nor UO_1785 (O_1785,N_22776,N_24809);
and UO_1786 (O_1786,N_22641,N_23487);
nand UO_1787 (O_1787,N_20877,N_20454);
nor UO_1788 (O_1788,N_23248,N_21397);
and UO_1789 (O_1789,N_20071,N_23859);
nor UO_1790 (O_1790,N_24920,N_24574);
or UO_1791 (O_1791,N_22024,N_21515);
nand UO_1792 (O_1792,N_24376,N_20403);
nand UO_1793 (O_1793,N_20831,N_21049);
nor UO_1794 (O_1794,N_24673,N_20311);
or UO_1795 (O_1795,N_20779,N_21240);
nand UO_1796 (O_1796,N_23556,N_24779);
nor UO_1797 (O_1797,N_22653,N_20748);
and UO_1798 (O_1798,N_20832,N_22778);
and UO_1799 (O_1799,N_23319,N_24088);
or UO_1800 (O_1800,N_20601,N_23370);
and UO_1801 (O_1801,N_22529,N_22366);
or UO_1802 (O_1802,N_20431,N_21531);
nand UO_1803 (O_1803,N_24930,N_22773);
and UO_1804 (O_1804,N_22758,N_20283);
or UO_1805 (O_1805,N_22869,N_23633);
and UO_1806 (O_1806,N_22519,N_20458);
nor UO_1807 (O_1807,N_24515,N_23928);
nand UO_1808 (O_1808,N_23756,N_23489);
nor UO_1809 (O_1809,N_21418,N_20485);
and UO_1810 (O_1810,N_20897,N_20762);
nand UO_1811 (O_1811,N_24782,N_20703);
nand UO_1812 (O_1812,N_21779,N_24316);
nand UO_1813 (O_1813,N_21206,N_20868);
and UO_1814 (O_1814,N_22811,N_20462);
nor UO_1815 (O_1815,N_24146,N_23224);
nand UO_1816 (O_1816,N_22615,N_22261);
and UO_1817 (O_1817,N_21244,N_20416);
nand UO_1818 (O_1818,N_20658,N_21379);
and UO_1819 (O_1819,N_23945,N_21369);
nor UO_1820 (O_1820,N_24105,N_20385);
nor UO_1821 (O_1821,N_21710,N_24797);
or UO_1822 (O_1822,N_21519,N_20714);
nor UO_1823 (O_1823,N_24244,N_21013);
nor UO_1824 (O_1824,N_21847,N_23934);
or UO_1825 (O_1825,N_24237,N_23200);
and UO_1826 (O_1826,N_21540,N_24129);
nand UO_1827 (O_1827,N_20067,N_24426);
or UO_1828 (O_1828,N_23187,N_22293);
nand UO_1829 (O_1829,N_21511,N_22407);
nor UO_1830 (O_1830,N_21538,N_20538);
nand UO_1831 (O_1831,N_23260,N_22314);
nor UO_1832 (O_1832,N_23408,N_22726);
nor UO_1833 (O_1833,N_20507,N_24554);
and UO_1834 (O_1834,N_24142,N_24696);
nand UO_1835 (O_1835,N_22007,N_22601);
nor UO_1836 (O_1836,N_23241,N_21274);
nor UO_1837 (O_1837,N_23536,N_22528);
and UO_1838 (O_1838,N_21004,N_20095);
nor UO_1839 (O_1839,N_21230,N_23687);
and UO_1840 (O_1840,N_23562,N_22279);
or UO_1841 (O_1841,N_24959,N_20398);
or UO_1842 (O_1842,N_23186,N_24253);
nand UO_1843 (O_1843,N_24876,N_24966);
or UO_1844 (O_1844,N_24275,N_22800);
nand UO_1845 (O_1845,N_21384,N_24501);
nand UO_1846 (O_1846,N_20953,N_21409);
and UO_1847 (O_1847,N_23821,N_24739);
and UO_1848 (O_1848,N_24497,N_22123);
and UO_1849 (O_1849,N_21139,N_21536);
nand UO_1850 (O_1850,N_20425,N_21387);
or UO_1851 (O_1851,N_21158,N_22795);
nand UO_1852 (O_1852,N_22183,N_22437);
nand UO_1853 (O_1853,N_23006,N_21064);
or UO_1854 (O_1854,N_21518,N_20669);
or UO_1855 (O_1855,N_23261,N_20742);
and UO_1856 (O_1856,N_21829,N_20307);
nand UO_1857 (O_1857,N_21685,N_21905);
nor UO_1858 (O_1858,N_24201,N_22637);
nor UO_1859 (O_1859,N_23609,N_24278);
and UO_1860 (O_1860,N_24429,N_20498);
and UO_1861 (O_1861,N_20896,N_21823);
xor UO_1862 (O_1862,N_23378,N_23331);
or UO_1863 (O_1863,N_22808,N_22473);
or UO_1864 (O_1864,N_22263,N_20607);
nor UO_1865 (O_1865,N_21577,N_21185);
nor UO_1866 (O_1866,N_23391,N_23151);
or UO_1867 (O_1867,N_23054,N_20706);
nand UO_1868 (O_1868,N_21529,N_22245);
or UO_1869 (O_1869,N_22990,N_23207);
nor UO_1870 (O_1870,N_20230,N_20645);
or UO_1871 (O_1871,N_24678,N_20715);
nor UO_1872 (O_1872,N_23867,N_23895);
nand UO_1873 (O_1873,N_23797,N_20588);
nand UO_1874 (O_1874,N_21816,N_20438);
and UO_1875 (O_1875,N_22719,N_23118);
or UO_1876 (O_1876,N_21583,N_23387);
and UO_1877 (O_1877,N_20736,N_23218);
or UO_1878 (O_1878,N_23570,N_21423);
nand UO_1879 (O_1879,N_20638,N_21732);
or UO_1880 (O_1880,N_21236,N_22270);
or UO_1881 (O_1881,N_24940,N_24314);
or UO_1882 (O_1882,N_23775,N_22288);
nor UO_1883 (O_1883,N_20804,N_22092);
and UO_1884 (O_1884,N_23392,N_22803);
or UO_1885 (O_1885,N_24075,N_22200);
and UO_1886 (O_1886,N_21089,N_23063);
nand UO_1887 (O_1887,N_21982,N_20893);
nor UO_1888 (O_1888,N_22577,N_22469);
nand UO_1889 (O_1889,N_20700,N_20987);
nand UO_1890 (O_1890,N_22989,N_21291);
nor UO_1891 (O_1891,N_21002,N_24027);
nor UO_1892 (O_1892,N_20476,N_20028);
nand UO_1893 (O_1893,N_24422,N_22184);
or UO_1894 (O_1894,N_20599,N_23279);
and UO_1895 (O_1895,N_23863,N_22544);
nand UO_1896 (O_1896,N_22141,N_24681);
and UO_1897 (O_1897,N_21871,N_23211);
xor UO_1898 (O_1898,N_23925,N_24877);
nand UO_1899 (O_1899,N_24130,N_21745);
or UO_1900 (O_1900,N_23285,N_22187);
and UO_1901 (O_1901,N_24742,N_20276);
nand UO_1902 (O_1902,N_20217,N_20004);
nor UO_1903 (O_1903,N_20942,N_24867);
nor UO_1904 (O_1904,N_23363,N_21953);
or UO_1905 (O_1905,N_24639,N_23203);
nor UO_1906 (O_1906,N_24428,N_23371);
nand UO_1907 (O_1907,N_23270,N_21043);
and UO_1908 (O_1908,N_20746,N_20331);
or UO_1909 (O_1909,N_23732,N_20723);
and UO_1910 (O_1910,N_23485,N_20268);
nor UO_1911 (O_1911,N_22492,N_22299);
and UO_1912 (O_1912,N_22820,N_24255);
nand UO_1913 (O_1913,N_21496,N_21272);
nand UO_1914 (O_1914,N_23249,N_22788);
nor UO_1915 (O_1915,N_23825,N_24164);
and UO_1916 (O_1916,N_20782,N_24159);
nand UO_1917 (O_1917,N_21716,N_23765);
nor UO_1918 (O_1918,N_22409,N_22883);
or UO_1919 (O_1919,N_23237,N_21854);
and UO_1920 (O_1920,N_23251,N_20693);
or UO_1921 (O_1921,N_23619,N_23735);
and UO_1922 (O_1922,N_21651,N_20320);
nor UO_1923 (O_1923,N_20926,N_20140);
and UO_1924 (O_1924,N_20267,N_24022);
nor UO_1925 (O_1925,N_24186,N_20035);
nand UO_1926 (O_1926,N_20404,N_24957);
or UO_1927 (O_1927,N_22818,N_20949);
and UO_1928 (O_1928,N_24663,N_22754);
and UO_1929 (O_1929,N_24937,N_23683);
nor UO_1930 (O_1930,N_24986,N_23858);
nor UO_1931 (O_1931,N_22107,N_23395);
xor UO_1932 (O_1932,N_24202,N_24931);
xnor UO_1933 (O_1933,N_23696,N_22645);
nand UO_1934 (O_1934,N_24733,N_22945);
and UO_1935 (O_1935,N_24464,N_23601);
nor UO_1936 (O_1936,N_21612,N_23555);
and UO_1937 (O_1937,N_22489,N_22400);
and UO_1938 (O_1938,N_20418,N_23738);
and UO_1939 (O_1939,N_24608,N_21542);
nand UO_1940 (O_1940,N_23529,N_22930);
and UO_1941 (O_1941,N_23275,N_20007);
nor UO_1942 (O_1942,N_23192,N_24570);
or UO_1943 (O_1943,N_20340,N_24208);
nor UO_1944 (O_1944,N_22224,N_23759);
nand UO_1945 (O_1945,N_23522,N_24368);
xnor UO_1946 (O_1946,N_22767,N_24749);
and UO_1947 (O_1947,N_21070,N_21179);
nor UO_1948 (O_1948,N_23505,N_23234);
and UO_1949 (O_1949,N_24861,N_20491);
and UO_1950 (O_1950,N_21682,N_24312);
nand UO_1951 (O_1951,N_20039,N_23606);
nand UO_1952 (O_1952,N_23524,N_21804);
nand UO_1953 (O_1953,N_20196,N_21229);
or UO_1954 (O_1954,N_23230,N_20150);
and UO_1955 (O_1955,N_24384,N_20205);
nor UO_1956 (O_1956,N_24092,N_21142);
nand UO_1957 (O_1957,N_24351,N_23087);
or UO_1958 (O_1958,N_24315,N_24120);
and UO_1959 (O_1959,N_24132,N_21589);
nand UO_1960 (O_1960,N_24772,N_20338);
nor UO_1961 (O_1961,N_23496,N_21352);
or UO_1962 (O_1962,N_22560,N_20809);
nor UO_1963 (O_1963,N_23017,N_21654);
xor UO_1964 (O_1964,N_22574,N_23748);
and UO_1965 (O_1965,N_22928,N_23267);
nor UO_1966 (O_1966,N_20711,N_20486);
and UO_1967 (O_1967,N_21398,N_21307);
or UO_1968 (O_1968,N_21861,N_24133);
and UO_1969 (O_1969,N_23640,N_23157);
nand UO_1970 (O_1970,N_24783,N_23037);
nor UO_1971 (O_1971,N_24905,N_21611);
and UO_1972 (O_1972,N_22035,N_20834);
and UO_1973 (O_1973,N_23440,N_21362);
or UO_1974 (O_1974,N_23215,N_23919);
or UO_1975 (O_1975,N_23567,N_23612);
and UO_1976 (O_1976,N_23407,N_21099);
nand UO_1977 (O_1977,N_23523,N_24427);
xnor UO_1978 (O_1978,N_21347,N_21593);
or UO_1979 (O_1979,N_24032,N_21011);
or UO_1980 (O_1980,N_20357,N_21112);
or UO_1981 (O_1981,N_24756,N_23886);
or UO_1982 (O_1982,N_24514,N_20543);
nand UO_1983 (O_1983,N_22536,N_21413);
nand UO_1984 (O_1984,N_20786,N_22622);
nor UO_1985 (O_1985,N_21071,N_24751);
nor UO_1986 (O_1986,N_24511,N_23692);
nand UO_1987 (O_1987,N_23746,N_23189);
nand UO_1988 (O_1988,N_22649,N_20328);
and UO_1989 (O_1989,N_24397,N_21084);
or UO_1990 (O_1990,N_22458,N_22642);
and UO_1991 (O_1991,N_22513,N_22876);
nor UO_1992 (O_1992,N_22908,N_24140);
or UO_1993 (O_1993,N_24664,N_24478);
xnor UO_1994 (O_1994,N_24941,N_21312);
or UO_1995 (O_1995,N_21081,N_21156);
nand UO_1996 (O_1996,N_24929,N_24550);
or UO_1997 (O_1997,N_24513,N_20764);
nor UO_1998 (O_1998,N_23266,N_23975);
nand UO_1999 (O_1999,N_22006,N_22535);
or UO_2000 (O_2000,N_20201,N_20333);
and UO_2001 (O_2001,N_20363,N_24902);
nor UO_2002 (O_2002,N_20420,N_20708);
nor UO_2003 (O_2003,N_21746,N_23305);
nor UO_2004 (O_2004,N_22230,N_23906);
and UO_2005 (O_2005,N_22359,N_22448);
nor UO_2006 (O_2006,N_23823,N_21283);
nor UO_2007 (O_2007,N_24649,N_21191);
nand UO_2008 (O_2008,N_22925,N_23875);
nor UO_2009 (O_2009,N_21222,N_23497);
nand UO_2010 (O_2010,N_21400,N_22367);
nor UO_2011 (O_2011,N_23814,N_24033);
or UO_2012 (O_2012,N_21737,N_21923);
nand UO_2013 (O_2013,N_22801,N_22652);
nand UO_2014 (O_2014,N_24535,N_20076);
nor UO_2015 (O_2015,N_23543,N_24815);
nor UO_2016 (O_2016,N_23566,N_22972);
nand UO_2017 (O_2017,N_24804,N_24392);
and UO_2018 (O_2018,N_21772,N_24108);
nor UO_2019 (O_2019,N_24299,N_20227);
and UO_2020 (O_2020,N_21483,N_22497);
nand UO_2021 (O_2021,N_24578,N_20083);
nand UO_2022 (O_2022,N_20365,N_20337);
or UO_2023 (O_2023,N_20402,N_24656);
nand UO_2024 (O_2024,N_20021,N_23632);
and UO_2025 (O_2025,N_22953,N_21957);
nor UO_2026 (O_2026,N_20132,N_21132);
or UO_2027 (O_2027,N_20901,N_22014);
nor UO_2028 (O_2028,N_21165,N_23239);
nand UO_2029 (O_2029,N_22610,N_23703);
or UO_2030 (O_2030,N_24726,N_24110);
xnor UO_2031 (O_2031,N_24078,N_24932);
nor UO_2032 (O_2032,N_24310,N_23656);
nand UO_2033 (O_2033,N_21259,N_20049);
nor UO_2034 (O_2034,N_22375,N_23004);
nor UO_2035 (O_2035,N_24879,N_22247);
and UO_2036 (O_2036,N_22094,N_24516);
nor UO_2037 (O_2037,N_23959,N_21618);
or UO_2038 (O_2038,N_21174,N_21541);
and UO_2039 (O_2039,N_24537,N_24821);
or UO_2040 (O_2040,N_23125,N_20903);
and UO_2041 (O_2041,N_23802,N_21566);
or UO_2042 (O_2042,N_20142,N_24084);
nor UO_2043 (O_2043,N_24874,N_21558);
nor UO_2044 (O_2044,N_24074,N_23052);
or UO_2045 (O_2045,N_20840,N_20202);
nor UO_2046 (O_2046,N_24548,N_20886);
nor UO_2047 (O_2047,N_21143,N_24477);
and UO_2048 (O_2048,N_21513,N_22418);
and UO_2049 (O_2049,N_21290,N_24273);
nand UO_2050 (O_2050,N_24271,N_24949);
nor UO_2051 (O_2051,N_21466,N_24447);
or UO_2052 (O_2052,N_24458,N_24054);
nand UO_2053 (O_2053,N_24947,N_22515);
or UO_2054 (O_2054,N_20312,N_22738);
nand UO_2055 (O_2055,N_21556,N_24763);
nand UO_2056 (O_2056,N_22128,N_21471);
or UO_2057 (O_2057,N_22752,N_23579);
and UO_2058 (O_2058,N_23281,N_23061);
nand UO_2059 (O_2059,N_22269,N_24721);
nor UO_2060 (O_2060,N_20682,N_24968);
and UO_2061 (O_2061,N_20930,N_23000);
and UO_2062 (O_2062,N_24709,N_24597);
and UO_2063 (O_2063,N_22060,N_20938);
nand UO_2064 (O_2064,N_24469,N_23910);
nand UO_2065 (O_2065,N_22460,N_22636);
or UO_2066 (O_2066,N_24910,N_22751);
or UO_2067 (O_2067,N_20323,N_23968);
nand UO_2068 (O_2068,N_23360,N_21650);
nand UO_2069 (O_2069,N_20735,N_21878);
nand UO_2070 (O_2070,N_23626,N_20613);
nor UO_2071 (O_2071,N_24072,N_20823);
nand UO_2072 (O_2072,N_23458,N_23999);
and UO_2073 (O_2073,N_24557,N_24961);
nand UO_2074 (O_2074,N_22376,N_20517);
or UO_2075 (O_2075,N_24174,N_23199);
nor UO_2076 (O_2076,N_24479,N_22743);
nand UO_2077 (O_2077,N_21201,N_24849);
or UO_2078 (O_2078,N_21490,N_23347);
and UO_2079 (O_2079,N_20696,N_22567);
nand UO_2080 (O_2080,N_24896,N_22720);
or UO_2081 (O_2081,N_24213,N_22253);
and UO_2082 (O_2082,N_23009,N_22099);
nor UO_2083 (O_2083,N_21753,N_20435);
and UO_2084 (O_2084,N_23636,N_21250);
nand UO_2085 (O_2085,N_21141,N_21940);
and UO_2086 (O_2086,N_20977,N_21835);
nor UO_2087 (O_2087,N_22324,N_22182);
and UO_2088 (O_2088,N_20913,N_24774);
nand UO_2089 (O_2089,N_20371,N_24530);
nand UO_2090 (O_2090,N_22295,N_20604);
and UO_2091 (O_2091,N_24261,N_24175);
or UO_2092 (O_2092,N_22875,N_23660);
nor UO_2093 (O_2093,N_24799,N_20767);
nand UO_2094 (O_2094,N_20553,N_20023);
and UO_2095 (O_2095,N_23326,N_23969);
nand UO_2096 (O_2096,N_22950,N_20798);
and UO_2097 (O_2097,N_20444,N_21478);
or UO_2098 (O_2098,N_23100,N_24780);
or UO_2099 (O_2099,N_23316,N_24483);
nand UO_2100 (O_2100,N_22229,N_23067);
nand UO_2101 (O_2101,N_23547,N_21217);
nand UO_2102 (O_2102,N_20207,N_24827);
or UO_2103 (O_2103,N_23963,N_22135);
or UO_2104 (O_2104,N_22644,N_23762);
nand UO_2105 (O_2105,N_20086,N_24984);
nand UO_2106 (O_2106,N_20946,N_20863);
nor UO_2107 (O_2107,N_21073,N_21068);
or UO_2108 (O_2108,N_24926,N_22798);
nand UO_2109 (O_2109,N_23425,N_21741);
or UO_2110 (O_2110,N_23941,N_21160);
and UO_2111 (O_2111,N_20484,N_23366);
and UO_2112 (O_2112,N_23787,N_21402);
and UO_2113 (O_2113,N_22103,N_23811);
and UO_2114 (O_2114,N_22341,N_21788);
nor UO_2115 (O_2115,N_20239,N_22500);
nand UO_2116 (O_2116,N_23868,N_23092);
or UO_2117 (O_2117,N_22211,N_24323);
and UO_2118 (O_2118,N_23243,N_23935);
and UO_2119 (O_2119,N_23354,N_21396);
and UO_2120 (O_2120,N_22613,N_21877);
nand UO_2121 (O_2121,N_20409,N_21016);
and UO_2122 (O_2122,N_20469,N_21300);
nor UO_2123 (O_2123,N_22098,N_22008);
nand UO_2124 (O_2124,N_20082,N_20789);
or UO_2125 (O_2125,N_22906,N_22976);
or UO_2126 (O_2126,N_20483,N_21472);
and UO_2127 (O_2127,N_23445,N_23622);
nor UO_2128 (O_2128,N_22140,N_20050);
nand UO_2129 (O_2129,N_22609,N_23075);
nand UO_2130 (O_2130,N_24580,N_23049);
nor UO_2131 (O_2131,N_20172,N_22931);
nand UO_2132 (O_2132,N_20221,N_20280);
nor UO_2133 (O_2133,N_24922,N_21330);
and UO_2134 (O_2134,N_20597,N_24334);
nand UO_2135 (O_2135,N_24507,N_22495);
and UO_2136 (O_2136,N_23958,N_21891);
nor UO_2137 (O_2137,N_20349,N_20548);
nand UO_2138 (O_2138,N_24298,N_20862);
and UO_2139 (O_2139,N_21318,N_22775);
or UO_2140 (O_2140,N_21346,N_23460);
nand UO_2141 (O_2141,N_22498,N_23225);
or UO_2142 (O_2142,N_21702,N_22827);
or UO_2143 (O_2143,N_24319,N_21563);
and UO_2144 (O_2144,N_24918,N_23757);
or UO_2145 (O_2145,N_23605,N_20030);
and UO_2146 (O_2146,N_22576,N_24288);
or UO_2147 (O_2147,N_21215,N_24758);
or UO_2148 (O_2148,N_20730,N_24577);
or UO_2149 (O_2149,N_20350,N_22970);
or UO_2150 (O_2150,N_22463,N_22735);
and UO_2151 (O_2151,N_23838,N_22999);
nor UO_2152 (O_2152,N_21424,N_20386);
or UO_2153 (O_2153,N_21735,N_21888);
nor UO_2154 (O_2154,N_21298,N_22579);
nor UO_2155 (O_2155,N_24307,N_22695);
or UO_2156 (O_2156,N_20768,N_21768);
nor UO_2157 (O_2157,N_20147,N_20560);
nor UO_2158 (O_2158,N_21088,N_22480);
or UO_2159 (O_2159,N_20755,N_21770);
nand UO_2160 (O_2160,N_23602,N_23554);
or UO_2161 (O_2161,N_20087,N_20719);
nor UO_2162 (O_2162,N_21616,N_22023);
nand UO_2163 (O_2163,N_20488,N_24228);
and UO_2164 (O_2164,N_20876,N_22273);
nand UO_2165 (O_2165,N_24629,N_21024);
nand UO_2166 (O_2166,N_20165,N_21797);
and UO_2167 (O_2167,N_23954,N_20772);
nor UO_2168 (O_2168,N_23209,N_21331);
nand UO_2169 (O_2169,N_24326,N_24361);
nand UO_2170 (O_2170,N_23256,N_21749);
nor UO_2171 (O_2171,N_24002,N_21780);
nor UO_2172 (O_2172,N_24638,N_21469);
nand UO_2173 (O_2173,N_22918,N_24206);
nand UO_2174 (O_2174,N_24411,N_24925);
and UO_2175 (O_2175,N_20998,N_20301);
nand UO_2176 (O_2176,N_21807,N_23310);
nand UO_2177 (O_2177,N_23298,N_20962);
or UO_2178 (O_2178,N_21793,N_21153);
or UO_2179 (O_2179,N_21161,N_20056);
and UO_2180 (O_2180,N_22571,N_22977);
or UO_2181 (O_2181,N_24007,N_21475);
nand UO_2182 (O_2182,N_24165,N_21401);
and UO_2183 (O_2183,N_22533,N_24505);
and UO_2184 (O_2184,N_20400,N_21925);
nand UO_2185 (O_2185,N_24747,N_22892);
nand UO_2186 (O_2186,N_20180,N_22815);
nand UO_2187 (O_2187,N_24053,N_22830);
nand UO_2188 (O_2188,N_20304,N_23768);
nor UO_2189 (O_2189,N_20345,N_21436);
nor UO_2190 (O_2190,N_23776,N_23299);
and UO_2191 (O_2191,N_21093,N_20944);
or UO_2192 (O_2192,N_23197,N_20577);
nand UO_2193 (O_2193,N_21690,N_21752);
and UO_2194 (O_2194,N_24187,N_23240);
nand UO_2195 (O_2195,N_22662,N_23860);
nor UO_2196 (O_2196,N_20990,N_24828);
and UO_2197 (O_2197,N_21502,N_20537);
or UO_2198 (O_2198,N_21069,N_23164);
nor UO_2199 (O_2199,N_21376,N_24145);
nand UO_2200 (O_2200,N_24880,N_22417);
or UO_2201 (O_2201,N_20727,N_22797);
nor UO_2202 (O_2202,N_24634,N_21382);
nand UO_2203 (O_2203,N_21530,N_20510);
or UO_2204 (O_2204,N_22017,N_22683);
nor UO_2205 (O_2205,N_24642,N_24387);
nand UO_2206 (O_2206,N_20282,N_24038);
nor UO_2207 (O_2207,N_20970,N_21533);
nand UO_2208 (O_2208,N_24161,N_22783);
nand UO_2209 (O_2209,N_21860,N_24866);
nor UO_2210 (O_2210,N_24848,N_22149);
nor UO_2211 (O_2211,N_23862,N_22391);
nand UO_2212 (O_2212,N_20527,N_20689);
nand UO_2213 (O_2213,N_21900,N_20666);
or UO_2214 (O_2214,N_22411,N_24615);
and UO_2215 (O_2215,N_20054,N_24841);
xnor UO_2216 (O_2216,N_24024,N_21974);
nand UO_2217 (O_2217,N_23961,N_23993);
or UO_2218 (O_2218,N_24391,N_20129);
and UO_2219 (O_2219,N_22040,N_24676);
nor UO_2220 (O_2220,N_24770,N_24716);
and UO_2221 (O_2221,N_21978,N_23981);
or UO_2222 (O_2222,N_20255,N_22205);
nand UO_2223 (O_2223,N_21889,N_22291);
and UO_2224 (O_2224,N_20550,N_23865);
and UO_2225 (O_2225,N_22207,N_22401);
nor UO_2226 (O_2226,N_21608,N_21812);
nor UO_2227 (O_2227,N_20466,N_21297);
nor UO_2228 (O_2228,N_20127,N_22398);
nor UO_2229 (O_2229,N_23604,N_23321);
and UO_2230 (O_2230,N_23837,N_22088);
nor UO_2231 (O_2231,N_20362,N_22680);
and UO_2232 (O_2232,N_23325,N_21097);
and UO_2233 (O_2233,N_21032,N_24786);
and UO_2234 (O_2234,N_22471,N_21756);
nor UO_2235 (O_2235,N_23176,N_21689);
or UO_2236 (O_2236,N_23593,N_21627);
or UO_2237 (O_2237,N_23112,N_24454);
nor UO_2238 (O_2238,N_22837,N_24197);
or UO_2239 (O_2239,N_21152,N_22572);
nor UO_2240 (O_2240,N_21278,N_22962);
nor UO_2241 (O_2241,N_21249,N_24194);
and UO_2242 (O_2242,N_22330,N_22218);
nand UO_2243 (O_2243,N_22027,N_22909);
nand UO_2244 (O_2244,N_22691,N_24657);
and UO_2245 (O_2245,N_21181,N_20555);
nand UO_2246 (O_2246,N_21477,N_24370);
nor UO_2247 (O_2247,N_22749,N_21933);
or UO_2248 (O_2248,N_20294,N_23312);
nor UO_2249 (O_2249,N_20687,N_23412);
or UO_2250 (O_2250,N_21910,N_21707);
and UO_2251 (O_2251,N_22392,N_24158);
and UO_2252 (O_2252,N_22698,N_23401);
or UO_2253 (O_2253,N_22034,N_23154);
or UO_2254 (O_2254,N_22514,N_24823);
nor UO_2255 (O_2255,N_24588,N_21914);
or UO_2256 (O_2256,N_20197,N_21619);
and UO_2257 (O_2257,N_24435,N_20566);
nor UO_2258 (O_2258,N_22146,N_23901);
nor UO_2259 (O_2259,N_23024,N_21271);
nand UO_2260 (O_2260,N_22241,N_22705);
nand UO_2261 (O_2261,N_24665,N_21214);
xnor UO_2262 (O_2262,N_24063,N_24740);
or UO_2263 (O_2263,N_21607,N_23452);
nand UO_2264 (O_2264,N_24242,N_22028);
or UO_2265 (O_2265,N_22382,N_23685);
and UO_2266 (O_2266,N_21227,N_20780);
nor UO_2267 (O_2267,N_23161,N_20053);
nor UO_2268 (O_2268,N_23323,N_24430);
or UO_2269 (O_2269,N_23876,N_24840);
nor UO_2270 (O_2270,N_20415,N_20213);
nand UO_2271 (O_2271,N_24461,N_23816);
or UO_2272 (O_2272,N_20191,N_22998);
nor UO_2273 (O_2273,N_21794,N_24266);
and UO_2274 (O_2274,N_20284,N_24286);
and UO_2275 (O_2275,N_23217,N_20552);
nor UO_2276 (O_2276,N_21575,N_20558);
and UO_2277 (O_2277,N_23766,N_21692);
nand UO_2278 (O_2278,N_21849,N_22203);
nand UO_2279 (O_2279,N_24970,N_23950);
or UO_2280 (O_2280,N_22465,N_23089);
and UO_2281 (O_2281,N_22054,N_22228);
nor UO_2282 (O_2282,N_21432,N_21375);
nand UO_2283 (O_2283,N_22594,N_23026);
xor UO_2284 (O_2284,N_24243,N_24330);
nor UO_2285 (O_2285,N_23525,N_22106);
nor UO_2286 (O_2286,N_22983,N_24109);
nand UO_2287 (O_2287,N_21783,N_20940);
and UO_2288 (O_2288,N_24386,N_22249);
nor UO_2289 (O_2289,N_21711,N_23276);
nor UO_2290 (O_2290,N_22340,N_21967);
nor UO_2291 (O_2291,N_20655,N_22052);
nor UO_2292 (O_2292,N_22524,N_20943);
or UO_2293 (O_2293,N_21764,N_20234);
and UO_2294 (O_2294,N_23502,N_24682);
and UO_2295 (O_2295,N_20869,N_21255);
or UO_2296 (O_2296,N_23353,N_24416);
nor UO_2297 (O_2297,N_20513,N_24776);
or UO_2298 (O_2298,N_22730,N_22276);
or UO_2299 (O_2299,N_20524,N_21973);
nand UO_2300 (O_2300,N_21193,N_21065);
nand UO_2301 (O_2301,N_20579,N_21454);
and UO_2302 (O_2302,N_21728,N_20704);
and UO_2303 (O_2303,N_20300,N_24234);
nand UO_2304 (O_2304,N_23102,N_22806);
nand UO_2305 (O_2305,N_24890,N_21087);
nand UO_2306 (O_2306,N_21219,N_20091);
and UO_2307 (O_2307,N_23388,N_21949);
or UO_2308 (O_2308,N_24595,N_24446);
and UO_2309 (O_2309,N_20915,N_22708);
or UO_2310 (O_2310,N_22608,N_20670);
or UO_2311 (O_2311,N_21104,N_21406);
and UO_2312 (O_2312,N_22157,N_23513);
and UO_2313 (O_2313,N_21762,N_21909);
or UO_2314 (O_2314,N_24865,N_23739);
and UO_2315 (O_2315,N_20747,N_24701);
nand UO_2316 (O_2316,N_22079,N_20941);
nor UO_2317 (O_2317,N_20310,N_23394);
or UO_2318 (O_2318,N_20726,N_23653);
nand UO_2319 (O_2319,N_20819,N_21587);
nor UO_2320 (O_2320,N_22185,N_24276);
and UO_2321 (O_2321,N_21411,N_22286);
nand UO_2322 (O_2322,N_21117,N_21876);
nand UO_2323 (O_2323,N_24209,N_21267);
nor UO_2324 (O_2324,N_23824,N_22654);
nor UO_2325 (O_2325,N_21453,N_24409);
or UO_2326 (O_2326,N_21992,N_20497);
nand UO_2327 (O_2327,N_21609,N_22305);
and UO_2328 (O_2328,N_23168,N_24635);
nand UO_2329 (O_2329,N_24013,N_24871);
nand UO_2330 (O_2330,N_22323,N_23939);
nor UO_2331 (O_2331,N_23431,N_22557);
or UO_2332 (O_2332,N_22239,N_22233);
nand UO_2333 (O_2333,N_21460,N_20468);
nand UO_2334 (O_2334,N_22478,N_21594);
and UO_2335 (O_2335,N_23904,N_22248);
and UO_2336 (O_2336,N_21140,N_21319);
nand UO_2337 (O_2337,N_22575,N_20917);
xor UO_2338 (O_2338,N_22274,N_24247);
nand UO_2339 (O_2339,N_23537,N_23830);
and UO_2340 (O_2340,N_24898,N_24908);
nand UO_2341 (O_2341,N_24199,N_23093);
and UO_2342 (O_2342,N_23586,N_21254);
and UO_2343 (O_2343,N_23761,N_24953);
nor UO_2344 (O_2344,N_24832,N_23088);
or UO_2345 (O_2345,N_22420,N_20412);
nand UO_2346 (O_2346,N_22777,N_22961);
xor UO_2347 (O_2347,N_22151,N_21027);
and UO_2348 (O_2348,N_21051,N_21833);
and UO_2349 (O_2349,N_20720,N_20346);
nor UO_2350 (O_2350,N_22942,N_20536);
or UO_2351 (O_2351,N_20605,N_23789);
or UO_2352 (O_2352,N_22548,N_24252);
nor UO_2353 (O_2353,N_21207,N_24814);
or UO_2354 (O_2354,N_22272,N_22280);
nor UO_2355 (O_2355,N_24628,N_21106);
and UO_2356 (O_2356,N_21686,N_20563);
or UO_2357 (O_2357,N_22723,N_22734);
and UO_2358 (O_2358,N_23409,N_24506);
nand UO_2359 (O_2359,N_22831,N_21455);
xnor UO_2360 (O_2360,N_24070,N_23818);
nor UO_2361 (O_2361,N_24979,N_24558);
nand UO_2362 (O_2362,N_24371,N_20133);
nor UO_2363 (O_2363,N_24730,N_24103);
nand UO_2364 (O_2364,N_24593,N_22115);
and UO_2365 (O_2365,N_24852,N_21748);
and UO_2366 (O_2366,N_20393,N_20187);
nand UO_2367 (O_2367,N_21962,N_21293);
or UO_2368 (O_2368,N_20947,N_23169);
nor UO_2369 (O_2369,N_21535,N_24459);
nor UO_2370 (O_2370,N_20390,N_20678);
or UO_2371 (O_2371,N_22737,N_23563);
and UO_2372 (O_2372,N_22321,N_21017);
nor UO_2373 (O_2373,N_20364,N_20908);
or UO_2374 (O_2374,N_23580,N_23072);
and UO_2375 (O_2375,N_23571,N_20143);
nor UO_2376 (O_2376,N_20986,N_23884);
and UO_2377 (O_2377,N_21996,N_22235);
and UO_2378 (O_2378,N_20791,N_21055);
nor UO_2379 (O_2379,N_23955,N_21928);
or UO_2380 (O_2380,N_20971,N_24141);
and UO_2381 (O_2381,N_23099,N_24349);
nor UO_2382 (O_2382,N_20651,N_21023);
nand UO_2383 (O_2383,N_20756,N_24474);
or UO_2384 (O_2384,N_20775,N_23630);
or UO_2385 (O_2385,N_23953,N_20422);
nand UO_2386 (O_2386,N_20424,N_24889);
or UO_2387 (O_2387,N_21326,N_23022);
nor UO_2388 (O_2388,N_21985,N_22821);
xnor UO_2389 (O_2389,N_22347,N_23842);
and UO_2390 (O_2390,N_24693,N_22142);
and UO_2391 (O_2391,N_20228,N_21547);
or UO_2392 (O_2392,N_20680,N_21881);
xnor UO_2393 (O_2393,N_24126,N_24156);
or UO_2394 (O_2394,N_23459,N_20574);
or UO_2395 (O_2395,N_24859,N_22600);
or UO_2396 (O_2396,N_22944,N_23717);
nor UO_2397 (O_2397,N_22078,N_22336);
nor UO_2398 (O_2398,N_20115,N_21799);
or UO_2399 (O_2399,N_21988,N_22281);
nor UO_2400 (O_2400,N_24785,N_23056);
or UO_2401 (O_2401,N_20066,N_23798);
nand UO_2402 (O_2402,N_20212,N_24935);
nand UO_2403 (O_2403,N_24878,N_23159);
or UO_2404 (O_2404,N_21656,N_21567);
nand UO_2405 (O_2405,N_20576,N_24343);
nor UO_2406 (O_2406,N_24630,N_23977);
nor UO_2407 (O_2407,N_20314,N_23962);
nand UO_2408 (O_2408,N_20882,N_24728);
nand UO_2409 (O_2409,N_22443,N_21727);
and UO_2410 (O_2410,N_24708,N_22155);
or UO_2411 (O_2411,N_24179,N_20808);
nor UO_2412 (O_2412,N_24844,N_22955);
nor UO_2413 (O_2413,N_24875,N_20152);
nor UO_2414 (O_2414,N_20586,N_23731);
or UO_2415 (O_2415,N_23213,N_20467);
nand UO_2416 (O_2416,N_24856,N_23889);
nor UO_2417 (O_2417,N_22677,N_21834);
nor UO_2418 (O_2418,N_22271,N_23829);
nor UO_2419 (O_2419,N_23849,N_22590);
nand UO_2420 (O_2420,N_24148,N_22566);
or UO_2421 (O_2421,N_23755,N_22125);
or UO_2422 (O_2422,N_24977,N_20797);
nand UO_2423 (O_2423,N_21146,N_21937);
and UO_2424 (O_2424,N_21574,N_21968);
nor UO_2425 (O_2425,N_21448,N_21348);
nand UO_2426 (O_2426,N_21691,N_23038);
nand UO_2427 (O_2427,N_21150,N_23730);
or UO_2428 (O_2428,N_24567,N_22334);
and UO_2429 (O_2429,N_24176,N_21626);
nand UO_2430 (O_2430,N_21120,N_22444);
nor UO_2431 (O_2431,N_23949,N_21242);
nand UO_2432 (O_2432,N_24950,N_21771);
nand UO_2433 (O_2433,N_20238,N_23980);
nand UO_2434 (O_2434,N_21373,N_24122);
and UO_2435 (O_2435,N_22899,N_21555);
and UO_2436 (O_2436,N_20352,N_24192);
nand UO_2437 (O_2437,N_20370,N_24532);
nor UO_2438 (O_2438,N_21127,N_23688);
nand UO_2439 (O_2439,N_20088,N_22275);
xnor UO_2440 (O_2440,N_24900,N_20124);
or UO_2441 (O_2441,N_23190,N_21704);
nor UO_2442 (O_2442,N_23324,N_22154);
or UO_2443 (O_2443,N_21234,N_22179);
nand UO_2444 (O_2444,N_22181,N_22362);
nor UO_2445 (O_2445,N_21270,N_21085);
nand UO_2446 (O_2446,N_20373,N_20379);
nor UO_2447 (O_2447,N_23107,N_22582);
nor UO_2448 (O_2448,N_20388,N_21056);
nand UO_2449 (O_2449,N_20235,N_24616);
and UO_2450 (O_2450,N_23074,N_23924);
or UO_2451 (O_2451,N_22068,N_21465);
and UO_2452 (O_2452,N_24744,N_20610);
and UO_2453 (O_2453,N_21010,N_23293);
or UO_2454 (O_2454,N_21610,N_21526);
or UO_2455 (O_2455,N_20222,N_23662);
or UO_2456 (O_2456,N_20712,N_23784);
nand UO_2457 (O_2457,N_21801,N_22081);
nand UO_2458 (O_2458,N_24825,N_22640);
nand UO_2459 (O_2459,N_20859,N_22414);
or UO_2460 (O_2460,N_21364,N_24831);
or UO_2461 (O_2461,N_21086,N_23671);
and UO_2462 (O_2462,N_20785,N_20226);
or UO_2463 (O_2463,N_23851,N_22118);
and UO_2464 (O_2464,N_21148,N_24344);
nor UO_2465 (O_2465,N_23874,N_21853);
and UO_2466 (O_2466,N_20925,N_22672);
and UO_2467 (O_2467,N_20773,N_21305);
xnor UO_2468 (O_2468,N_20078,N_22186);
nand UO_2469 (O_2469,N_24769,N_20939);
xor UO_2470 (O_2470,N_20612,N_23001);
xnor UO_2471 (O_2471,N_22244,N_23166);
or UO_2472 (O_2472,N_24614,N_23449);
and UO_2473 (O_2473,N_22611,N_24306);
nor UO_2474 (O_2474,N_24095,N_24223);
nand UO_2475 (O_2475,N_20106,N_21571);
and UO_2476 (O_2476,N_23801,N_24727);
nor UO_2477 (O_2477,N_21672,N_20432);
xor UO_2478 (O_2478,N_20262,N_23861);
or UO_2479 (O_2479,N_22277,N_21866);
nand UO_2480 (O_2480,N_20254,N_23873);
or UO_2481 (O_2481,N_23156,N_22898);
xor UO_2482 (O_2482,N_23400,N_21831);
nor UO_2483 (O_2483,N_20833,N_23592);
nand UO_2484 (O_2484,N_22527,N_22725);
and UO_2485 (O_2485,N_21778,N_20000);
nand UO_2486 (O_2486,N_22217,N_21474);
and UO_2487 (O_2487,N_23675,N_21765);
nand UO_2488 (O_2488,N_24207,N_20303);
or UO_2489 (O_2489,N_24956,N_20273);
nor UO_2490 (O_2490,N_24777,N_21007);
and UO_2491 (O_2491,N_22792,N_20348);
nand UO_2492 (O_2492,N_24346,N_20571);
or UO_2493 (O_2493,N_23119,N_23396);
nor UO_2494 (O_2494,N_23399,N_24801);
and UO_2495 (O_2495,N_22661,N_23429);
nand UO_2496 (O_2496,N_20092,N_22335);
nor UO_2497 (O_2497,N_22538,N_24633);
or UO_2498 (O_2498,N_20631,N_22278);
and UO_2499 (O_2499,N_24596,N_22834);
or UO_2500 (O_2500,N_23660,N_22284);
nand UO_2501 (O_2501,N_24822,N_21572);
or UO_2502 (O_2502,N_21319,N_22978);
nor UO_2503 (O_2503,N_22409,N_24537);
nor UO_2504 (O_2504,N_22625,N_23918);
nand UO_2505 (O_2505,N_24366,N_24652);
or UO_2506 (O_2506,N_20576,N_21511);
and UO_2507 (O_2507,N_22236,N_23015);
nand UO_2508 (O_2508,N_20683,N_20475);
nand UO_2509 (O_2509,N_24299,N_24669);
nand UO_2510 (O_2510,N_22120,N_22689);
nand UO_2511 (O_2511,N_20902,N_23588);
nand UO_2512 (O_2512,N_24245,N_23448);
and UO_2513 (O_2513,N_21126,N_21224);
or UO_2514 (O_2514,N_21224,N_20949);
and UO_2515 (O_2515,N_21711,N_24096);
nand UO_2516 (O_2516,N_21044,N_23152);
and UO_2517 (O_2517,N_23605,N_24418);
and UO_2518 (O_2518,N_20507,N_24545);
and UO_2519 (O_2519,N_20655,N_23086);
or UO_2520 (O_2520,N_23445,N_20881);
nand UO_2521 (O_2521,N_20641,N_20697);
nor UO_2522 (O_2522,N_23266,N_22854);
and UO_2523 (O_2523,N_23334,N_20824);
nor UO_2524 (O_2524,N_20872,N_23054);
nand UO_2525 (O_2525,N_22772,N_23268);
nand UO_2526 (O_2526,N_20420,N_24175);
or UO_2527 (O_2527,N_20222,N_24670);
nor UO_2528 (O_2528,N_23035,N_21083);
and UO_2529 (O_2529,N_24211,N_24264);
nand UO_2530 (O_2530,N_24046,N_20914);
and UO_2531 (O_2531,N_24599,N_23769);
or UO_2532 (O_2532,N_21388,N_21724);
nor UO_2533 (O_2533,N_24981,N_20419);
nor UO_2534 (O_2534,N_23337,N_23252);
or UO_2535 (O_2535,N_22224,N_20649);
nand UO_2536 (O_2536,N_20306,N_23531);
nand UO_2537 (O_2537,N_20461,N_22342);
or UO_2538 (O_2538,N_22546,N_22608);
and UO_2539 (O_2539,N_22364,N_24357);
or UO_2540 (O_2540,N_22914,N_24721);
and UO_2541 (O_2541,N_23684,N_23015);
nor UO_2542 (O_2542,N_22374,N_21345);
nor UO_2543 (O_2543,N_21961,N_24176);
nor UO_2544 (O_2544,N_20836,N_24999);
nand UO_2545 (O_2545,N_24599,N_24971);
or UO_2546 (O_2546,N_20311,N_21174);
nor UO_2547 (O_2547,N_20119,N_24155);
and UO_2548 (O_2548,N_23075,N_20624);
or UO_2549 (O_2549,N_22990,N_21927);
nand UO_2550 (O_2550,N_21806,N_21830);
or UO_2551 (O_2551,N_24933,N_23720);
nand UO_2552 (O_2552,N_22731,N_20097);
and UO_2553 (O_2553,N_23748,N_20177);
and UO_2554 (O_2554,N_22549,N_24466);
and UO_2555 (O_2555,N_22296,N_21141);
nand UO_2556 (O_2556,N_22902,N_20489);
nor UO_2557 (O_2557,N_22418,N_24722);
or UO_2558 (O_2558,N_24522,N_24084);
or UO_2559 (O_2559,N_23499,N_22958);
nand UO_2560 (O_2560,N_23902,N_24046);
or UO_2561 (O_2561,N_24172,N_24464);
nor UO_2562 (O_2562,N_21344,N_22118);
or UO_2563 (O_2563,N_23486,N_20821);
nor UO_2564 (O_2564,N_23776,N_23425);
nand UO_2565 (O_2565,N_21099,N_21056);
nand UO_2566 (O_2566,N_23174,N_24930);
and UO_2567 (O_2567,N_22962,N_21347);
xor UO_2568 (O_2568,N_21512,N_20221);
nand UO_2569 (O_2569,N_20530,N_21071);
nor UO_2570 (O_2570,N_21233,N_23291);
nand UO_2571 (O_2571,N_23283,N_20800);
nor UO_2572 (O_2572,N_24609,N_24629);
nand UO_2573 (O_2573,N_23782,N_20505);
nand UO_2574 (O_2574,N_24846,N_24984);
or UO_2575 (O_2575,N_20856,N_21553);
nor UO_2576 (O_2576,N_21119,N_20193);
and UO_2577 (O_2577,N_24832,N_20479);
nand UO_2578 (O_2578,N_22076,N_20981);
nand UO_2579 (O_2579,N_23530,N_24736);
or UO_2580 (O_2580,N_24309,N_22359);
or UO_2581 (O_2581,N_22940,N_21423);
nor UO_2582 (O_2582,N_20365,N_23859);
nand UO_2583 (O_2583,N_22737,N_20981);
or UO_2584 (O_2584,N_24312,N_23653);
nand UO_2585 (O_2585,N_24545,N_20976);
and UO_2586 (O_2586,N_24988,N_21769);
nor UO_2587 (O_2587,N_20577,N_21801);
xor UO_2588 (O_2588,N_21340,N_21514);
or UO_2589 (O_2589,N_24064,N_22640);
and UO_2590 (O_2590,N_23967,N_20807);
or UO_2591 (O_2591,N_20437,N_24032);
or UO_2592 (O_2592,N_24422,N_24062);
nand UO_2593 (O_2593,N_23550,N_24254);
nor UO_2594 (O_2594,N_20013,N_22797);
nor UO_2595 (O_2595,N_23648,N_20669);
or UO_2596 (O_2596,N_20430,N_24256);
or UO_2597 (O_2597,N_20300,N_20415);
xor UO_2598 (O_2598,N_23164,N_23450);
nor UO_2599 (O_2599,N_20940,N_20815);
and UO_2600 (O_2600,N_23604,N_23969);
nor UO_2601 (O_2601,N_20190,N_22844);
nor UO_2602 (O_2602,N_23997,N_20262);
and UO_2603 (O_2603,N_20344,N_20472);
nor UO_2604 (O_2604,N_24974,N_22889);
and UO_2605 (O_2605,N_21859,N_20566);
and UO_2606 (O_2606,N_21343,N_24607);
and UO_2607 (O_2607,N_23489,N_20372);
nand UO_2608 (O_2608,N_20229,N_20830);
nor UO_2609 (O_2609,N_20935,N_22358);
nand UO_2610 (O_2610,N_23108,N_21185);
or UO_2611 (O_2611,N_21857,N_21108);
nand UO_2612 (O_2612,N_22228,N_24580);
and UO_2613 (O_2613,N_24896,N_23470);
nor UO_2614 (O_2614,N_24297,N_22513);
nand UO_2615 (O_2615,N_23511,N_23014);
nor UO_2616 (O_2616,N_23615,N_22397);
nand UO_2617 (O_2617,N_23161,N_22900);
or UO_2618 (O_2618,N_21966,N_21081);
nor UO_2619 (O_2619,N_21284,N_22863);
nor UO_2620 (O_2620,N_24726,N_24154);
or UO_2621 (O_2621,N_21353,N_23114);
or UO_2622 (O_2622,N_20227,N_20313);
and UO_2623 (O_2623,N_24580,N_20889);
and UO_2624 (O_2624,N_20204,N_20048);
nand UO_2625 (O_2625,N_20045,N_22450);
nand UO_2626 (O_2626,N_23732,N_21701);
nor UO_2627 (O_2627,N_22588,N_23635);
nand UO_2628 (O_2628,N_20050,N_23035);
nand UO_2629 (O_2629,N_23296,N_20701);
and UO_2630 (O_2630,N_21932,N_22158);
xnor UO_2631 (O_2631,N_22925,N_23504);
and UO_2632 (O_2632,N_23870,N_24960);
or UO_2633 (O_2633,N_20606,N_22299);
or UO_2634 (O_2634,N_23841,N_23593);
and UO_2635 (O_2635,N_20723,N_20925);
nand UO_2636 (O_2636,N_21050,N_23037);
nor UO_2637 (O_2637,N_24251,N_23258);
and UO_2638 (O_2638,N_21096,N_22056);
and UO_2639 (O_2639,N_21116,N_20770);
nor UO_2640 (O_2640,N_21838,N_20895);
nor UO_2641 (O_2641,N_20695,N_24617);
nand UO_2642 (O_2642,N_21688,N_21406);
nand UO_2643 (O_2643,N_20191,N_20975);
nand UO_2644 (O_2644,N_23350,N_22651);
nor UO_2645 (O_2645,N_23442,N_20271);
and UO_2646 (O_2646,N_20903,N_22126);
and UO_2647 (O_2647,N_23140,N_21032);
nor UO_2648 (O_2648,N_23859,N_23176);
nor UO_2649 (O_2649,N_21463,N_20875);
nor UO_2650 (O_2650,N_24652,N_21148);
and UO_2651 (O_2651,N_22203,N_20182);
nand UO_2652 (O_2652,N_20764,N_24129);
or UO_2653 (O_2653,N_22777,N_21364);
or UO_2654 (O_2654,N_20883,N_23333);
and UO_2655 (O_2655,N_21537,N_20632);
nor UO_2656 (O_2656,N_22903,N_23543);
nand UO_2657 (O_2657,N_23979,N_23307);
and UO_2658 (O_2658,N_24443,N_24030);
nand UO_2659 (O_2659,N_21560,N_22827);
or UO_2660 (O_2660,N_22385,N_20404);
nand UO_2661 (O_2661,N_24544,N_20564);
nand UO_2662 (O_2662,N_24060,N_23479);
or UO_2663 (O_2663,N_23979,N_22402);
nand UO_2664 (O_2664,N_24241,N_20628);
or UO_2665 (O_2665,N_20335,N_22782);
nor UO_2666 (O_2666,N_24773,N_24354);
nand UO_2667 (O_2667,N_23559,N_21110);
and UO_2668 (O_2668,N_22058,N_24911);
xor UO_2669 (O_2669,N_21894,N_20399);
and UO_2670 (O_2670,N_20439,N_21686);
or UO_2671 (O_2671,N_23542,N_23484);
nand UO_2672 (O_2672,N_20900,N_21189);
nand UO_2673 (O_2673,N_20636,N_24443);
and UO_2674 (O_2674,N_23550,N_23067);
or UO_2675 (O_2675,N_23277,N_24102);
nor UO_2676 (O_2676,N_21153,N_22002);
or UO_2677 (O_2677,N_23326,N_23444);
or UO_2678 (O_2678,N_20209,N_20131);
nand UO_2679 (O_2679,N_24708,N_20642);
or UO_2680 (O_2680,N_20251,N_22888);
nor UO_2681 (O_2681,N_20473,N_24948);
nand UO_2682 (O_2682,N_23314,N_24030);
and UO_2683 (O_2683,N_20605,N_21982);
or UO_2684 (O_2684,N_24284,N_23074);
and UO_2685 (O_2685,N_20713,N_23260);
nor UO_2686 (O_2686,N_23440,N_24703);
xnor UO_2687 (O_2687,N_21913,N_22915);
nand UO_2688 (O_2688,N_22031,N_23919);
or UO_2689 (O_2689,N_21870,N_20398);
nor UO_2690 (O_2690,N_23151,N_21300);
or UO_2691 (O_2691,N_20665,N_24686);
and UO_2692 (O_2692,N_20204,N_20986);
nand UO_2693 (O_2693,N_22050,N_22021);
xnor UO_2694 (O_2694,N_21120,N_24814);
nor UO_2695 (O_2695,N_20585,N_24812);
or UO_2696 (O_2696,N_23678,N_20974);
and UO_2697 (O_2697,N_21138,N_22295);
nor UO_2698 (O_2698,N_24930,N_21838);
nor UO_2699 (O_2699,N_21731,N_23779);
nor UO_2700 (O_2700,N_21380,N_20426);
and UO_2701 (O_2701,N_22632,N_24736);
and UO_2702 (O_2702,N_20479,N_21781);
or UO_2703 (O_2703,N_24804,N_21698);
nand UO_2704 (O_2704,N_22584,N_22365);
and UO_2705 (O_2705,N_22622,N_21069);
or UO_2706 (O_2706,N_21932,N_22482);
nand UO_2707 (O_2707,N_23800,N_21551);
nand UO_2708 (O_2708,N_20053,N_24978);
nor UO_2709 (O_2709,N_22248,N_22308);
or UO_2710 (O_2710,N_20863,N_23842);
or UO_2711 (O_2711,N_20816,N_22353);
nand UO_2712 (O_2712,N_21740,N_21843);
nor UO_2713 (O_2713,N_24085,N_24189);
nor UO_2714 (O_2714,N_21845,N_21462);
nand UO_2715 (O_2715,N_22155,N_21950);
nor UO_2716 (O_2716,N_20069,N_22582);
nor UO_2717 (O_2717,N_24063,N_21377);
and UO_2718 (O_2718,N_20838,N_21906);
nor UO_2719 (O_2719,N_22592,N_22234);
and UO_2720 (O_2720,N_23074,N_20352);
nand UO_2721 (O_2721,N_23170,N_21376);
nor UO_2722 (O_2722,N_24760,N_20779);
nand UO_2723 (O_2723,N_23685,N_20429);
nor UO_2724 (O_2724,N_23140,N_22292);
nor UO_2725 (O_2725,N_23960,N_21589);
nor UO_2726 (O_2726,N_24733,N_21574);
nor UO_2727 (O_2727,N_23124,N_21056);
nand UO_2728 (O_2728,N_24149,N_23371);
nand UO_2729 (O_2729,N_22380,N_23757);
nand UO_2730 (O_2730,N_22371,N_20256);
or UO_2731 (O_2731,N_22246,N_21712);
nand UO_2732 (O_2732,N_24284,N_23236);
nor UO_2733 (O_2733,N_20379,N_21365);
nor UO_2734 (O_2734,N_22054,N_24367);
or UO_2735 (O_2735,N_23470,N_24255);
nand UO_2736 (O_2736,N_23019,N_20639);
and UO_2737 (O_2737,N_23788,N_20550);
nand UO_2738 (O_2738,N_21674,N_20835);
nand UO_2739 (O_2739,N_20458,N_20195);
xnor UO_2740 (O_2740,N_21495,N_22252);
and UO_2741 (O_2741,N_21355,N_20695);
nand UO_2742 (O_2742,N_24728,N_20286);
or UO_2743 (O_2743,N_21015,N_22748);
xnor UO_2744 (O_2744,N_20547,N_23106);
and UO_2745 (O_2745,N_23818,N_21465);
nor UO_2746 (O_2746,N_21433,N_22324);
nand UO_2747 (O_2747,N_20956,N_20274);
or UO_2748 (O_2748,N_21417,N_20437);
and UO_2749 (O_2749,N_22838,N_20537);
nand UO_2750 (O_2750,N_22625,N_24232);
or UO_2751 (O_2751,N_23070,N_22893);
nor UO_2752 (O_2752,N_20989,N_21685);
nand UO_2753 (O_2753,N_21281,N_24474);
nor UO_2754 (O_2754,N_20705,N_21913);
nor UO_2755 (O_2755,N_22919,N_23214);
or UO_2756 (O_2756,N_21842,N_24357);
or UO_2757 (O_2757,N_24756,N_20762);
nand UO_2758 (O_2758,N_22501,N_24884);
nand UO_2759 (O_2759,N_20086,N_22107);
or UO_2760 (O_2760,N_23943,N_23926);
nor UO_2761 (O_2761,N_20282,N_22161);
nor UO_2762 (O_2762,N_23479,N_20750);
xor UO_2763 (O_2763,N_24302,N_23511);
or UO_2764 (O_2764,N_24664,N_24767);
and UO_2765 (O_2765,N_20699,N_22008);
nand UO_2766 (O_2766,N_24650,N_24341);
and UO_2767 (O_2767,N_20841,N_20347);
or UO_2768 (O_2768,N_24630,N_24320);
nand UO_2769 (O_2769,N_21484,N_24678);
and UO_2770 (O_2770,N_21367,N_22012);
nor UO_2771 (O_2771,N_20304,N_24012);
or UO_2772 (O_2772,N_22876,N_22242);
nor UO_2773 (O_2773,N_20552,N_20240);
and UO_2774 (O_2774,N_23743,N_20755);
or UO_2775 (O_2775,N_20704,N_22288);
nor UO_2776 (O_2776,N_20656,N_22085);
or UO_2777 (O_2777,N_23140,N_24724);
and UO_2778 (O_2778,N_22156,N_24641);
nor UO_2779 (O_2779,N_23241,N_23063);
and UO_2780 (O_2780,N_23583,N_20189);
nand UO_2781 (O_2781,N_22792,N_20721);
and UO_2782 (O_2782,N_21498,N_20779);
nand UO_2783 (O_2783,N_22844,N_24193);
and UO_2784 (O_2784,N_20929,N_22417);
or UO_2785 (O_2785,N_22359,N_23513);
nand UO_2786 (O_2786,N_22269,N_20964);
nor UO_2787 (O_2787,N_22266,N_20517);
xor UO_2788 (O_2788,N_21834,N_24911);
nand UO_2789 (O_2789,N_20170,N_23103);
nand UO_2790 (O_2790,N_22056,N_23777);
or UO_2791 (O_2791,N_22102,N_24830);
or UO_2792 (O_2792,N_22019,N_23358);
or UO_2793 (O_2793,N_24316,N_21554);
nor UO_2794 (O_2794,N_22877,N_21169);
xnor UO_2795 (O_2795,N_20137,N_21707);
and UO_2796 (O_2796,N_23009,N_21363);
and UO_2797 (O_2797,N_23008,N_21035);
or UO_2798 (O_2798,N_22991,N_22684);
nor UO_2799 (O_2799,N_21074,N_23660);
nor UO_2800 (O_2800,N_24421,N_23136);
and UO_2801 (O_2801,N_23176,N_22892);
nor UO_2802 (O_2802,N_20002,N_21068);
or UO_2803 (O_2803,N_20656,N_22662);
or UO_2804 (O_2804,N_24769,N_23205);
or UO_2805 (O_2805,N_20298,N_20936);
nor UO_2806 (O_2806,N_20039,N_21749);
nor UO_2807 (O_2807,N_23943,N_24366);
and UO_2808 (O_2808,N_21420,N_21794);
nor UO_2809 (O_2809,N_21785,N_23103);
nor UO_2810 (O_2810,N_21996,N_22682);
xor UO_2811 (O_2811,N_23207,N_22478);
nor UO_2812 (O_2812,N_20420,N_23555);
xor UO_2813 (O_2813,N_20447,N_23579);
nand UO_2814 (O_2814,N_24843,N_22848);
or UO_2815 (O_2815,N_23645,N_24818);
or UO_2816 (O_2816,N_20257,N_24028);
and UO_2817 (O_2817,N_23789,N_20487);
and UO_2818 (O_2818,N_22607,N_20481);
and UO_2819 (O_2819,N_20270,N_23778);
or UO_2820 (O_2820,N_21636,N_23296);
or UO_2821 (O_2821,N_23888,N_23690);
xnor UO_2822 (O_2822,N_22969,N_23063);
nor UO_2823 (O_2823,N_23639,N_21399);
nor UO_2824 (O_2824,N_24998,N_24808);
and UO_2825 (O_2825,N_22834,N_21972);
nor UO_2826 (O_2826,N_22419,N_24815);
or UO_2827 (O_2827,N_20724,N_20337);
and UO_2828 (O_2828,N_23932,N_22391);
or UO_2829 (O_2829,N_24816,N_20687);
nand UO_2830 (O_2830,N_23014,N_24771);
nand UO_2831 (O_2831,N_22342,N_20229);
and UO_2832 (O_2832,N_23887,N_23794);
nand UO_2833 (O_2833,N_22090,N_20380);
xnor UO_2834 (O_2834,N_21366,N_20327);
nor UO_2835 (O_2835,N_21690,N_23602);
or UO_2836 (O_2836,N_20499,N_20210);
or UO_2837 (O_2837,N_21803,N_23333);
and UO_2838 (O_2838,N_22991,N_24934);
nor UO_2839 (O_2839,N_23290,N_20106);
or UO_2840 (O_2840,N_22744,N_24524);
nand UO_2841 (O_2841,N_21216,N_23539);
nand UO_2842 (O_2842,N_24054,N_21406);
nor UO_2843 (O_2843,N_20725,N_23003);
and UO_2844 (O_2844,N_23054,N_24631);
or UO_2845 (O_2845,N_20147,N_20997);
or UO_2846 (O_2846,N_23039,N_24753);
nand UO_2847 (O_2847,N_24417,N_20393);
and UO_2848 (O_2848,N_24826,N_20905);
nand UO_2849 (O_2849,N_23831,N_24049);
and UO_2850 (O_2850,N_22692,N_20220);
or UO_2851 (O_2851,N_21095,N_21710);
or UO_2852 (O_2852,N_22287,N_21902);
and UO_2853 (O_2853,N_23137,N_23519);
and UO_2854 (O_2854,N_20099,N_22381);
nand UO_2855 (O_2855,N_22757,N_23741);
and UO_2856 (O_2856,N_23944,N_24808);
nor UO_2857 (O_2857,N_21293,N_23333);
nor UO_2858 (O_2858,N_24053,N_23243);
nand UO_2859 (O_2859,N_22410,N_23091);
nand UO_2860 (O_2860,N_24109,N_24083);
nand UO_2861 (O_2861,N_22357,N_23875);
and UO_2862 (O_2862,N_20315,N_21445);
or UO_2863 (O_2863,N_20625,N_20047);
nand UO_2864 (O_2864,N_20967,N_24962);
and UO_2865 (O_2865,N_23462,N_21764);
xor UO_2866 (O_2866,N_23839,N_23952);
or UO_2867 (O_2867,N_21552,N_22867);
nand UO_2868 (O_2868,N_20461,N_21333);
or UO_2869 (O_2869,N_23240,N_21872);
or UO_2870 (O_2870,N_24004,N_23084);
nand UO_2871 (O_2871,N_20757,N_20022);
or UO_2872 (O_2872,N_23957,N_24625);
nor UO_2873 (O_2873,N_23582,N_20719);
or UO_2874 (O_2874,N_21621,N_22228);
or UO_2875 (O_2875,N_24763,N_22321);
nor UO_2876 (O_2876,N_20121,N_24335);
and UO_2877 (O_2877,N_22178,N_22965);
and UO_2878 (O_2878,N_23084,N_22679);
nor UO_2879 (O_2879,N_24937,N_20189);
and UO_2880 (O_2880,N_21005,N_21456);
nor UO_2881 (O_2881,N_24004,N_22803);
nor UO_2882 (O_2882,N_22904,N_20447);
and UO_2883 (O_2883,N_23685,N_22380);
nand UO_2884 (O_2884,N_21534,N_23769);
nor UO_2885 (O_2885,N_23078,N_23411);
or UO_2886 (O_2886,N_23035,N_23917);
nor UO_2887 (O_2887,N_23634,N_24992);
nand UO_2888 (O_2888,N_22192,N_23661);
nand UO_2889 (O_2889,N_23018,N_23994);
and UO_2890 (O_2890,N_22292,N_22240);
nor UO_2891 (O_2891,N_21947,N_21418);
nand UO_2892 (O_2892,N_23242,N_20799);
or UO_2893 (O_2893,N_20607,N_24376);
nand UO_2894 (O_2894,N_23342,N_23765);
nand UO_2895 (O_2895,N_24472,N_21360);
nor UO_2896 (O_2896,N_23563,N_23753);
nor UO_2897 (O_2897,N_20971,N_24786);
nand UO_2898 (O_2898,N_24741,N_20584);
nand UO_2899 (O_2899,N_20051,N_21386);
nor UO_2900 (O_2900,N_20998,N_23678);
nor UO_2901 (O_2901,N_24849,N_22548);
and UO_2902 (O_2902,N_20508,N_21130);
and UO_2903 (O_2903,N_23786,N_21255);
and UO_2904 (O_2904,N_22452,N_23828);
or UO_2905 (O_2905,N_22473,N_21847);
or UO_2906 (O_2906,N_21819,N_24851);
or UO_2907 (O_2907,N_23708,N_23440);
nor UO_2908 (O_2908,N_22965,N_24291);
nor UO_2909 (O_2909,N_21195,N_24824);
and UO_2910 (O_2910,N_23180,N_22207);
or UO_2911 (O_2911,N_23207,N_20221);
nand UO_2912 (O_2912,N_22607,N_24146);
nand UO_2913 (O_2913,N_24312,N_21197);
nor UO_2914 (O_2914,N_24615,N_20223);
and UO_2915 (O_2915,N_20131,N_22077);
nand UO_2916 (O_2916,N_24132,N_20031);
or UO_2917 (O_2917,N_23118,N_24292);
nor UO_2918 (O_2918,N_24061,N_24087);
nand UO_2919 (O_2919,N_24562,N_20415);
or UO_2920 (O_2920,N_21012,N_23995);
and UO_2921 (O_2921,N_24024,N_23661);
or UO_2922 (O_2922,N_22254,N_21632);
nand UO_2923 (O_2923,N_21631,N_21525);
nand UO_2924 (O_2924,N_23822,N_20601);
xnor UO_2925 (O_2925,N_23816,N_20024);
or UO_2926 (O_2926,N_23731,N_22048);
and UO_2927 (O_2927,N_21031,N_23706);
or UO_2928 (O_2928,N_24216,N_20275);
nand UO_2929 (O_2929,N_24176,N_22663);
nand UO_2930 (O_2930,N_24298,N_24994);
nor UO_2931 (O_2931,N_22172,N_21361);
and UO_2932 (O_2932,N_20070,N_20012);
nand UO_2933 (O_2933,N_20697,N_24042);
and UO_2934 (O_2934,N_21634,N_24820);
nand UO_2935 (O_2935,N_20567,N_24794);
and UO_2936 (O_2936,N_20880,N_23334);
and UO_2937 (O_2937,N_20490,N_20867);
nand UO_2938 (O_2938,N_21216,N_21705);
nand UO_2939 (O_2939,N_21837,N_24315);
or UO_2940 (O_2940,N_24529,N_23232);
nor UO_2941 (O_2941,N_22838,N_20936);
or UO_2942 (O_2942,N_24755,N_22488);
or UO_2943 (O_2943,N_20180,N_23746);
nand UO_2944 (O_2944,N_21003,N_22220);
nand UO_2945 (O_2945,N_21726,N_21972);
nor UO_2946 (O_2946,N_21799,N_24023);
nand UO_2947 (O_2947,N_21745,N_22583);
nor UO_2948 (O_2948,N_21454,N_24953);
or UO_2949 (O_2949,N_22085,N_22612);
or UO_2950 (O_2950,N_23980,N_20763);
nand UO_2951 (O_2951,N_21339,N_23987);
nand UO_2952 (O_2952,N_23255,N_21507);
and UO_2953 (O_2953,N_22287,N_24076);
nor UO_2954 (O_2954,N_24808,N_24434);
nor UO_2955 (O_2955,N_20529,N_21509);
and UO_2956 (O_2956,N_24505,N_21719);
nor UO_2957 (O_2957,N_20881,N_22590);
or UO_2958 (O_2958,N_21726,N_21829);
and UO_2959 (O_2959,N_23828,N_24244);
and UO_2960 (O_2960,N_20570,N_21721);
nand UO_2961 (O_2961,N_21594,N_20418);
nor UO_2962 (O_2962,N_24461,N_20643);
and UO_2963 (O_2963,N_22741,N_21785);
and UO_2964 (O_2964,N_23875,N_23383);
and UO_2965 (O_2965,N_21245,N_20048);
nor UO_2966 (O_2966,N_23870,N_23853);
or UO_2967 (O_2967,N_21232,N_21550);
nand UO_2968 (O_2968,N_22813,N_22109);
nor UO_2969 (O_2969,N_20426,N_22137);
or UO_2970 (O_2970,N_24239,N_24975);
or UO_2971 (O_2971,N_23369,N_21330);
and UO_2972 (O_2972,N_21816,N_21430);
nand UO_2973 (O_2973,N_22730,N_20593);
or UO_2974 (O_2974,N_22738,N_21478);
or UO_2975 (O_2975,N_23122,N_23099);
or UO_2976 (O_2976,N_21694,N_23307);
nand UO_2977 (O_2977,N_22630,N_23374);
nand UO_2978 (O_2978,N_23524,N_22645);
xnor UO_2979 (O_2979,N_24060,N_22310);
or UO_2980 (O_2980,N_21153,N_23620);
nand UO_2981 (O_2981,N_22223,N_21201);
or UO_2982 (O_2982,N_20944,N_24324);
nor UO_2983 (O_2983,N_24318,N_21522);
nand UO_2984 (O_2984,N_23543,N_20827);
nor UO_2985 (O_2985,N_21903,N_24121);
and UO_2986 (O_2986,N_23420,N_24548);
xnor UO_2987 (O_2987,N_20634,N_23829);
nand UO_2988 (O_2988,N_21763,N_24500);
nor UO_2989 (O_2989,N_20019,N_24191);
nor UO_2990 (O_2990,N_22857,N_20179);
nand UO_2991 (O_2991,N_23403,N_23452);
nand UO_2992 (O_2992,N_22809,N_21550);
nor UO_2993 (O_2993,N_23984,N_22743);
nor UO_2994 (O_2994,N_23946,N_20308);
nor UO_2995 (O_2995,N_20221,N_21541);
xnor UO_2996 (O_2996,N_22920,N_23466);
nand UO_2997 (O_2997,N_20297,N_23990);
nor UO_2998 (O_2998,N_24043,N_22416);
nand UO_2999 (O_2999,N_22928,N_21429);
endmodule