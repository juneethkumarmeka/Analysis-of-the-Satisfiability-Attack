module basic_5000_50000_5000_50_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_3163,In_1847);
xor U1 (N_1,In_1209,In_1779);
nand U2 (N_2,In_2676,In_235);
nand U3 (N_3,In_3846,In_3862);
nand U4 (N_4,In_830,In_1293);
xnor U5 (N_5,In_2915,In_1201);
and U6 (N_6,In_2924,In_94);
nor U7 (N_7,In_874,In_796);
nand U8 (N_8,In_2316,In_2935);
or U9 (N_9,In_1588,In_629);
nand U10 (N_10,In_284,In_1283);
xor U11 (N_11,In_3430,In_4730);
nor U12 (N_12,In_1336,In_2794);
or U13 (N_13,In_3975,In_1634);
and U14 (N_14,In_1548,In_2402);
and U15 (N_15,In_2582,In_2731);
and U16 (N_16,In_4067,In_2807);
nand U17 (N_17,In_4866,In_2173);
nand U18 (N_18,In_4082,In_2266);
nor U19 (N_19,In_670,In_909);
or U20 (N_20,In_2944,In_2784);
nor U21 (N_21,In_3161,In_3244);
xor U22 (N_22,In_434,In_2526);
or U23 (N_23,In_2626,In_2801);
and U24 (N_24,In_817,In_2346);
xor U25 (N_25,In_387,In_2700);
xor U26 (N_26,In_4898,In_958);
nor U27 (N_27,In_1223,In_1449);
and U28 (N_28,In_1257,In_2713);
and U29 (N_29,In_1113,In_4800);
or U30 (N_30,In_3081,In_4461);
nor U31 (N_31,In_4643,In_3612);
or U32 (N_32,In_13,In_2971);
xnor U33 (N_33,In_3374,In_4709);
or U34 (N_34,In_3656,In_1103);
nand U35 (N_35,In_3921,In_4627);
xnor U36 (N_36,In_2323,In_2991);
and U37 (N_37,In_1076,In_3491);
nand U38 (N_38,In_38,In_2348);
and U39 (N_39,In_3233,In_2992);
nand U40 (N_40,In_2870,In_880);
xor U41 (N_41,In_4687,In_1644);
xor U42 (N_42,In_4137,In_2565);
xor U43 (N_43,In_4167,In_3788);
nand U44 (N_44,In_1082,In_4160);
and U45 (N_45,In_3818,In_3977);
nor U46 (N_46,In_1664,In_3532);
nand U47 (N_47,In_587,In_1185);
nand U48 (N_48,In_3471,In_1682);
or U49 (N_49,In_4396,In_3669);
and U50 (N_50,In_1901,In_1235);
nor U51 (N_51,In_4855,In_3392);
nor U52 (N_52,In_47,In_4758);
xor U53 (N_53,In_4518,In_4099);
or U54 (N_54,In_4216,In_245);
or U55 (N_55,In_2256,In_299);
nor U56 (N_56,In_3222,In_2852);
nor U57 (N_57,In_3727,In_4931);
or U58 (N_58,In_617,In_1470);
xor U59 (N_59,In_288,In_4420);
nand U60 (N_60,In_1582,In_1724);
nand U61 (N_61,In_3900,In_620);
xor U62 (N_62,In_802,In_1893);
or U63 (N_63,In_4839,In_3472);
and U64 (N_64,In_4304,In_2366);
xor U65 (N_65,In_3752,In_3844);
xor U66 (N_66,In_150,In_3484);
nand U67 (N_67,In_4400,In_756);
nand U68 (N_68,In_2524,In_4103);
nor U69 (N_69,In_84,In_3053);
or U70 (N_70,In_4483,In_4163);
nand U71 (N_71,In_2500,In_2043);
xor U72 (N_72,In_142,In_3954);
nor U73 (N_73,In_230,In_1073);
xnor U74 (N_74,In_1921,In_2357);
nand U75 (N_75,In_530,In_3740);
nor U76 (N_76,In_4311,In_4958);
nor U77 (N_77,In_611,In_4006);
nor U78 (N_78,In_3601,In_3774);
nor U79 (N_79,In_1922,In_3200);
xnor U80 (N_80,In_433,In_4437);
xor U81 (N_81,In_4845,In_4531);
nor U82 (N_82,In_3529,In_3040);
or U83 (N_83,In_2920,In_159);
nor U84 (N_84,In_4155,In_1315);
xnor U85 (N_85,In_4057,In_3603);
nor U86 (N_86,In_1729,In_3531);
and U87 (N_87,In_4588,In_3477);
nand U88 (N_88,In_3762,In_183);
or U89 (N_89,In_382,In_411);
nand U90 (N_90,In_103,In_352);
or U91 (N_91,In_4040,In_379);
or U92 (N_92,In_31,In_1062);
or U93 (N_93,In_2377,In_2730);
and U94 (N_94,In_4548,In_4296);
nand U95 (N_95,In_2652,In_3877);
nor U96 (N_96,In_4021,In_373);
and U97 (N_97,In_4278,In_2781);
nor U98 (N_98,In_4092,In_673);
nand U99 (N_99,In_4339,In_307);
nor U100 (N_100,In_3747,In_2650);
and U101 (N_101,In_3409,In_4312);
nand U102 (N_102,In_3434,In_157);
xnor U103 (N_103,In_3453,In_4517);
nand U104 (N_104,In_3613,In_4862);
or U105 (N_105,In_1422,In_4952);
or U106 (N_106,In_4481,In_1690);
and U107 (N_107,In_1743,In_1608);
nor U108 (N_108,In_1983,In_372);
xor U109 (N_109,In_3057,In_2286);
and U110 (N_110,In_1437,In_4540);
and U111 (N_111,In_4847,In_984);
and U112 (N_112,In_3971,In_4796);
nor U113 (N_113,In_4118,In_4392);
or U114 (N_114,In_3843,In_1683);
and U115 (N_115,In_2374,In_4752);
or U116 (N_116,In_3263,In_3940);
xnor U117 (N_117,In_1672,In_374);
xnor U118 (N_118,In_2188,In_4946);
xnor U119 (N_119,In_1280,In_468);
nor U120 (N_120,In_4478,In_3480);
xnor U121 (N_121,In_675,In_4275);
or U122 (N_122,In_1046,In_507);
nor U123 (N_123,In_2169,In_3969);
nor U124 (N_124,In_2831,In_4041);
nand U125 (N_125,In_4843,In_716);
xor U126 (N_126,In_208,In_2670);
nor U127 (N_127,In_3547,In_3391);
and U128 (N_128,In_3456,In_4575);
or U129 (N_129,In_1857,In_3772);
and U130 (N_130,In_1445,In_812);
xor U131 (N_131,In_2958,In_2654);
or U132 (N_132,In_1291,In_4428);
xor U133 (N_133,In_2150,In_3277);
nor U134 (N_134,In_935,In_2176);
xor U135 (N_135,In_128,In_2613);
xnor U136 (N_136,In_2736,In_676);
and U137 (N_137,In_3572,In_4004);
or U138 (N_138,In_3379,In_1090);
or U139 (N_139,In_2985,In_1942);
nand U140 (N_140,In_4723,In_701);
xor U141 (N_141,In_3732,In_1392);
or U142 (N_142,In_3756,In_4161);
or U143 (N_143,In_414,In_349);
xnor U144 (N_144,In_912,In_2957);
xnor U145 (N_145,In_143,In_1428);
nand U146 (N_146,In_3691,In_1190);
or U147 (N_147,In_557,In_118);
or U148 (N_148,In_2548,In_1747);
nand U149 (N_149,In_4525,In_3965);
or U150 (N_150,In_4105,In_4840);
xor U151 (N_151,In_3201,In_2849);
xor U152 (N_152,In_166,In_3111);
or U153 (N_153,In_4008,In_4417);
and U154 (N_154,In_3338,In_1177);
or U155 (N_155,In_4231,In_4317);
nand U156 (N_156,In_3243,In_718);
nor U157 (N_157,In_2139,In_1171);
nor U158 (N_158,In_2035,In_943);
and U159 (N_159,In_1840,In_4642);
nand U160 (N_160,In_1267,In_4712);
and U161 (N_161,In_3696,In_839);
or U162 (N_162,In_4580,In_1850);
or U163 (N_163,In_4554,In_2115);
and U164 (N_164,In_1909,In_3426);
xor U165 (N_165,In_4033,In_879);
or U166 (N_166,In_4301,In_1249);
nand U167 (N_167,In_843,In_290);
or U168 (N_168,In_2232,In_1621);
nand U169 (N_169,In_4268,In_1534);
and U170 (N_170,In_556,In_3319);
and U171 (N_171,In_661,In_81);
and U172 (N_172,In_3036,In_397);
and U173 (N_173,In_3520,In_558);
nand U174 (N_174,In_3675,In_4812);
xor U175 (N_175,In_2235,In_3976);
or U176 (N_176,In_1828,In_2386);
or U177 (N_177,In_1247,In_2273);
nor U178 (N_178,In_2146,In_3079);
xor U179 (N_179,In_1054,In_140);
or U180 (N_180,In_1360,In_1898);
or U181 (N_181,In_4024,In_893);
nand U182 (N_182,In_3488,In_1920);
nor U183 (N_183,In_4562,In_4943);
xor U184 (N_184,In_3194,In_4571);
nor U185 (N_185,In_216,In_4954);
and U186 (N_186,In_1806,In_3982);
nand U187 (N_187,In_4613,In_898);
or U188 (N_188,In_4599,In_1361);
xnor U189 (N_189,In_2279,In_515);
nor U190 (N_190,In_1938,In_1162);
and U191 (N_191,In_4212,In_4508);
nor U192 (N_192,In_4783,In_1492);
and U193 (N_193,In_44,In_2701);
nor U194 (N_194,In_4093,In_2275);
xnor U195 (N_195,In_560,In_4269);
xnor U196 (N_196,In_3497,In_4402);
nand U197 (N_197,In_3284,In_4334);
nand U198 (N_198,In_2056,In_938);
nand U199 (N_199,In_4539,In_3638);
nor U200 (N_200,In_1357,In_516);
or U201 (N_201,In_4373,In_1098);
and U202 (N_202,In_462,In_1302);
xor U203 (N_203,In_4104,In_2726);
nand U204 (N_204,In_4715,In_4754);
xnor U205 (N_205,In_3781,In_1482);
nor U206 (N_206,In_630,In_4115);
xnor U207 (N_207,In_1452,In_933);
and U208 (N_208,In_492,In_4698);
and U209 (N_209,In_1897,In_895);
and U210 (N_210,In_3049,In_1741);
nand U211 (N_211,In_357,In_3265);
nand U212 (N_212,In_4357,In_932);
and U213 (N_213,In_2495,In_1380);
and U214 (N_214,In_4425,In_3294);
xnor U215 (N_215,In_4832,In_2978);
nor U216 (N_216,In_116,In_4462);
nand U217 (N_217,In_1345,In_2682);
xnor U218 (N_218,In_74,In_2536);
or U219 (N_219,In_914,In_4859);
xor U220 (N_220,In_4177,In_4658);
xnor U221 (N_221,In_1862,In_4264);
nand U222 (N_222,In_593,In_3397);
nor U223 (N_223,In_1892,In_3);
nor U224 (N_224,In_4519,In_43);
nand U225 (N_225,In_4767,In_3022);
or U226 (N_226,In_2998,In_3701);
xnor U227 (N_227,In_3678,In_4725);
and U228 (N_228,In_443,In_3330);
and U229 (N_229,In_3981,In_805);
and U230 (N_230,In_732,In_551);
xnor U231 (N_231,In_3168,In_1289);
nor U232 (N_232,In_1958,In_1000);
nand U233 (N_233,In_71,In_1918);
nand U234 (N_234,In_2246,In_613);
xnor U235 (N_235,In_745,In_2274);
nand U236 (N_236,In_2887,In_3867);
nor U237 (N_237,In_336,In_3719);
and U238 (N_238,In_695,In_999);
or U239 (N_239,In_1487,In_2276);
nor U240 (N_240,In_794,In_4852);
nand U241 (N_241,In_1584,In_4565);
or U242 (N_242,In_48,In_4731);
nor U243 (N_243,In_2101,In_552);
and U244 (N_244,In_3512,In_4039);
and U245 (N_245,In_2660,In_4883);
and U246 (N_246,In_1125,In_1028);
xor U247 (N_247,In_700,In_470);
nor U248 (N_248,In_4633,In_3513);
nor U249 (N_249,In_2356,In_2282);
nor U250 (N_250,In_1978,In_4419);
xnor U251 (N_251,In_4998,In_4026);
and U252 (N_252,In_2567,In_2017);
xor U253 (N_253,In_4720,In_1455);
nand U254 (N_254,In_635,In_427);
or U255 (N_255,In_348,In_1144);
or U256 (N_256,In_1870,In_1242);
nor U257 (N_257,In_3619,In_4504);
or U258 (N_258,In_453,In_393);
or U259 (N_259,In_663,In_4434);
nor U260 (N_260,In_1308,In_3348);
or U261 (N_261,In_2010,In_192);
nand U262 (N_262,In_4361,In_1006);
and U263 (N_263,In_3326,In_2866);
xor U264 (N_264,In_1436,In_3645);
or U265 (N_265,In_1085,In_24);
xnor U266 (N_266,In_1593,In_4764);
and U267 (N_267,In_644,In_1513);
xnor U268 (N_268,In_2679,In_2787);
nand U269 (N_269,In_4193,In_1170);
and U270 (N_270,In_2551,In_465);
or U271 (N_271,In_184,In_3879);
nand U272 (N_272,In_748,In_4695);
or U273 (N_273,In_3096,In_197);
nand U274 (N_274,In_4438,In_4779);
or U275 (N_275,In_224,In_2381);
or U276 (N_276,In_3190,In_3058);
nand U277 (N_277,In_1434,In_877);
xor U278 (N_278,In_979,In_369);
xnor U279 (N_279,In_4255,In_3245);
nand U280 (N_280,In_2163,In_3533);
xnor U281 (N_281,In_1488,In_3490);
nor U282 (N_282,In_2623,In_3563);
xnor U283 (N_283,In_3817,In_1860);
xnor U284 (N_284,In_1498,In_2481);
or U285 (N_285,In_321,In_4611);
or U286 (N_286,In_4672,In_870);
nand U287 (N_287,In_5,In_1522);
nor U288 (N_288,In_3511,In_1295);
nor U289 (N_289,In_4607,In_4223);
xnor U290 (N_290,In_650,In_618);
xor U291 (N_291,In_4102,In_4581);
and U292 (N_292,In_211,In_2552);
nand U293 (N_293,In_1216,In_945);
xnor U294 (N_294,In_2543,In_27);
xor U295 (N_295,In_2760,In_182);
or U296 (N_296,In_4684,In_4975);
nand U297 (N_297,In_3254,In_3218);
and U298 (N_298,In_4248,In_4170);
nand U299 (N_299,In_2394,In_2219);
xnor U300 (N_300,In_2504,In_477);
xor U301 (N_301,In_2303,In_1941);
nand U302 (N_302,In_2186,In_2984);
and U303 (N_303,In_1632,In_2953);
nor U304 (N_304,In_3298,In_3083);
nor U305 (N_305,In_4657,In_1719);
and U306 (N_306,In_512,In_4310);
and U307 (N_307,In_1204,In_486);
and U308 (N_308,In_158,In_899);
nand U309 (N_309,In_73,In_2087);
or U310 (N_310,In_2696,In_1238);
xnor U311 (N_311,In_4234,In_1571);
nand U312 (N_312,In_1679,In_3179);
and U313 (N_313,In_1050,In_3112);
xor U314 (N_314,In_3813,In_2969);
xnor U315 (N_315,In_4221,In_4697);
nor U316 (N_316,In_1102,In_2006);
nor U317 (N_317,In_819,In_4964);
nor U318 (N_318,In_862,In_2638);
xnor U319 (N_319,In_161,In_4838);
xor U320 (N_320,In_187,In_4463);
nor U321 (N_321,In_4661,In_3894);
nand U322 (N_322,In_2688,In_647);
nand U323 (N_323,In_937,In_1167);
or U324 (N_324,In_4207,In_3116);
nor U325 (N_325,In_3288,In_2245);
and U326 (N_326,In_3653,In_1335);
and U327 (N_327,In_2860,In_2307);
or U328 (N_328,In_407,In_1025);
nand U329 (N_329,In_2418,In_2349);
xnor U330 (N_330,In_4511,In_1585);
or U331 (N_331,In_4865,In_3560);
or U332 (N_332,In_4919,In_2990);
nand U333 (N_333,In_1301,In_4809);
and U334 (N_334,In_4543,In_3935);
or U335 (N_335,In_3052,In_2370);
xor U336 (N_336,In_1602,In_1970);
and U337 (N_337,In_4176,In_3371);
xnor U338 (N_338,In_3523,In_181);
and U339 (N_339,In_3489,In_589);
nor U340 (N_340,In_3259,In_400);
xnor U341 (N_341,In_3594,In_2624);
and U342 (N_342,In_3717,In_513);
nor U343 (N_343,In_3467,In_3069);
nand U344 (N_344,In_4753,In_2367);
nand U345 (N_345,In_2926,In_2075);
or U346 (N_346,In_2288,In_1936);
xnor U347 (N_347,In_298,In_2155);
or U348 (N_348,In_3147,In_4704);
nand U349 (N_349,In_1476,In_3094);
and U350 (N_350,In_2228,In_2981);
and U351 (N_351,In_1084,In_1788);
nand U352 (N_352,In_1869,In_3346);
nand U353 (N_353,In_2628,In_742);
nor U354 (N_354,In_621,In_3621);
or U355 (N_355,In_1839,In_4619);
or U356 (N_356,In_4716,In_1178);
or U357 (N_357,In_2559,In_2749);
or U358 (N_358,In_2950,In_3431);
nand U359 (N_359,In_2879,In_4646);
or U360 (N_360,In_3904,In_1776);
nor U361 (N_361,In_302,In_4593);
nor U362 (N_362,In_2554,In_241);
and U363 (N_363,In_3009,In_4644);
and U364 (N_364,In_2651,In_860);
nand U365 (N_365,In_2622,In_4046);
nor U366 (N_366,In_2941,In_4356);
or U367 (N_367,In_976,In_3577);
or U368 (N_368,In_129,In_2106);
or U369 (N_369,In_4579,In_3104);
xnor U370 (N_370,In_3987,In_2912);
nor U371 (N_371,In_916,In_3134);
or U372 (N_372,In_1848,In_2812);
or U373 (N_373,In_3249,In_2966);
or U374 (N_374,In_4963,In_4557);
nor U375 (N_375,In_1926,In_170);
nor U376 (N_376,In_3109,In_3041);
nor U377 (N_377,In_3272,In_845);
and U378 (N_378,In_566,In_1798);
and U379 (N_379,In_4666,In_1526);
nand U380 (N_380,In_3798,In_2472);
or U381 (N_381,In_3400,In_3652);
xnor U382 (N_382,In_381,In_3899);
nand U383 (N_383,In_2478,In_2222);
nor U384 (N_384,In_472,In_1056);
nor U385 (N_385,In_1406,In_1974);
or U386 (N_386,In_4533,In_4377);
or U387 (N_387,In_2332,In_1910);
nor U388 (N_388,In_814,In_1555);
or U389 (N_389,In_9,In_2345);
nand U390 (N_390,In_4923,In_1250);
xor U391 (N_391,In_1418,In_714);
nand U392 (N_392,In_1575,In_3293);
xor U393 (N_393,In_2514,In_4464);
nand U394 (N_394,In_3475,In_2782);
or U395 (N_395,In_1141,In_237);
xnor U396 (N_396,In_2886,In_1736);
and U397 (N_397,In_2513,In_3372);
xnor U398 (N_398,In_3558,In_1424);
and U399 (N_399,In_2637,In_4388);
nor U400 (N_400,In_1935,In_4773);
and U401 (N_401,In_919,In_3928);
xnor U402 (N_402,In_2837,In_1221);
and U403 (N_403,In_437,In_97);
or U404 (N_404,In_3639,In_1887);
xor U405 (N_405,In_218,In_1612);
or U406 (N_406,In_3801,In_3731);
xor U407 (N_407,In_2857,In_1902);
xor U408 (N_408,In_1696,In_2502);
nand U409 (N_409,In_1040,In_1309);
nand U410 (N_410,In_596,In_2611);
nand U411 (N_411,In_778,In_994);
or U412 (N_412,In_4492,In_3395);
nand U413 (N_413,In_3256,In_2725);
and U414 (N_414,In_1078,In_3659);
and U415 (N_415,In_4808,In_2758);
nand U416 (N_416,In_137,In_4065);
and U417 (N_417,In_1464,In_2791);
nand U418 (N_418,In_2473,In_2681);
nor U419 (N_419,In_4215,In_2841);
nand U420 (N_420,In_114,In_2104);
or U421 (N_421,In_1230,In_3778);
or U422 (N_422,In_3151,In_982);
nand U423 (N_423,In_3988,In_190);
nor U424 (N_424,In_4078,In_3440);
nand U425 (N_425,In_1614,In_1687);
or U426 (N_426,In_2158,In_4499);
nor U427 (N_427,In_1448,In_2491);
and U428 (N_428,In_4397,In_3321);
nor U429 (N_429,In_1012,In_4950);
nand U430 (N_430,In_599,In_1415);
xor U431 (N_431,In_1229,In_894);
nand U432 (N_432,In_2803,In_2456);
nand U433 (N_433,In_3980,In_765);
nand U434 (N_434,In_693,In_2595);
or U435 (N_435,In_1382,In_4899);
xor U436 (N_436,In_4467,In_1947);
nand U437 (N_437,In_1739,In_4972);
or U438 (N_438,In_1874,In_2532);
or U439 (N_439,In_4894,In_3002);
nor U440 (N_440,In_1479,In_1899);
nand U441 (N_441,In_3852,In_4165);
xnor U442 (N_442,In_1782,In_4708);
and U443 (N_443,In_883,In_3177);
nor U444 (N_444,In_238,In_3016);
xnor U445 (N_445,In_3203,In_4653);
xor U446 (N_446,In_1425,In_3525);
nor U447 (N_447,In_3297,In_293);
nand U448 (N_448,In_1278,In_1883);
or U449 (N_449,In_4776,In_2260);
nor U450 (N_450,In_1419,In_49);
and U451 (N_451,In_2201,In_3310);
nand U452 (N_452,In_3084,In_3367);
or U453 (N_453,In_1663,In_1694);
nor U454 (N_454,In_583,In_4842);
and U455 (N_455,In_1960,In_744);
nor U456 (N_456,In_3253,In_1019);
nor U457 (N_457,In_2250,In_2918);
and U458 (N_458,In_4990,In_4288);
and U459 (N_459,In_3373,In_3470);
nand U460 (N_460,In_4445,In_834);
nand U461 (N_461,In_981,In_3303);
nand U462 (N_462,In_2468,In_4910);
nand U463 (N_463,In_2479,In_2878);
or U464 (N_464,In_1146,In_2973);
nand U465 (N_465,In_1510,In_2751);
nand U466 (N_466,In_3979,In_6);
or U467 (N_467,In_3349,In_416);
and U468 (N_468,In_2946,In_2819);
or U469 (N_469,In_672,In_3869);
or U470 (N_470,In_972,In_2223);
nor U471 (N_471,In_4470,In_2024);
and U472 (N_472,In_2662,In_4053);
and U473 (N_473,In_4335,In_1018);
nor U474 (N_474,In_4594,In_657);
nand U475 (N_475,In_3775,In_2949);
and U476 (N_476,In_347,In_2590);
and U477 (N_477,In_3993,In_3341);
nor U478 (N_478,In_4826,In_2009);
and U479 (N_479,In_2211,In_243);
nor U480 (N_480,In_4787,In_353);
nor U481 (N_481,In_2835,In_2675);
xor U482 (N_482,In_3441,In_523);
or U483 (N_483,In_3699,In_755);
nand U484 (N_484,In_2070,In_4940);
and U485 (N_485,In_1533,In_2207);
or U486 (N_486,In_474,In_4349);
nor U487 (N_487,In_3646,In_4127);
nand U488 (N_488,In_3276,In_1329);
or U489 (N_489,In_2641,In_602);
nor U490 (N_490,In_3290,In_2411);
nand U491 (N_491,In_1486,In_973);
and U492 (N_492,In_4541,In_858);
and U493 (N_493,In_4675,In_1271);
xnor U494 (N_494,In_3354,In_2134);
nand U495 (N_495,In_4825,In_4597);
or U496 (N_496,In_3212,In_482);
nor U497 (N_497,In_2724,In_1531);
or U498 (N_498,In_4768,In_2280);
and U499 (N_499,In_3683,In_1581);
xor U500 (N_500,In_168,In_392);
nand U501 (N_501,In_3251,In_10);
nor U502 (N_502,In_2627,In_2642);
or U503 (N_503,In_1307,In_3402);
nor U504 (N_504,In_4385,In_645);
or U505 (N_505,In_4453,In_2057);
nor U506 (N_506,In_319,In_873);
nor U507 (N_507,In_4079,In_1515);
xor U508 (N_508,In_3421,In_120);
or U509 (N_509,In_3665,In_3502);
nand U510 (N_510,In_4719,In_3792);
or U511 (N_511,In_33,In_1512);
or U512 (N_512,In_2511,In_4522);
and U513 (N_513,In_4226,In_2240);
and U514 (N_514,In_3361,In_4131);
or U515 (N_515,In_250,In_4589);
nor U516 (N_516,In_544,In_997);
and U517 (N_517,In_4934,In_4314);
xor U518 (N_518,In_974,In_4570);
nand U519 (N_519,In_3100,In_2177);
nor U520 (N_520,In_4932,In_4227);
and U521 (N_521,In_1086,In_4371);
or U522 (N_522,In_4376,In_4393);
nor U523 (N_523,In_80,In_2925);
nand U524 (N_524,In_3636,In_3539);
and U525 (N_525,In_1882,In_1379);
and U526 (N_526,In_14,In_508);
or U527 (N_527,In_3758,In_4480);
and U528 (N_528,In_3716,In_126);
or U529 (N_529,In_4906,In_4202);
nand U530 (N_530,In_1175,In_1689);
xnor U531 (N_531,In_1708,In_2436);
and U532 (N_532,In_2234,In_356);
nor U533 (N_533,In_3322,In_2257);
nor U534 (N_534,In_4213,In_1383);
and U535 (N_535,In_761,In_2538);
and U536 (N_536,In_4380,In_4410);
and U537 (N_537,In_731,In_186);
and U538 (N_538,In_2195,In_3712);
xor U539 (N_539,In_1346,In_760);
nand U540 (N_540,In_2102,In_322);
nand U541 (N_541,In_3439,In_801);
nor U542 (N_542,In_3029,In_2980);
nand U543 (N_543,In_3428,In_3056);
and U544 (N_544,In_1945,In_966);
nand U545 (N_545,In_2046,In_4164);
xor U546 (N_546,In_1709,In_1868);
nor U547 (N_547,In_2923,In_884);
and U548 (N_548,In_1398,In_3810);
or U549 (N_549,In_691,In_4407);
and U550 (N_550,In_4660,In_3845);
xor U551 (N_551,In_4512,In_1866);
nand U552 (N_552,In_390,In_2405);
and U553 (N_553,In_3583,In_3575);
or U554 (N_554,In_3450,In_3495);
nand U555 (N_555,In_3469,In_65);
nand U556 (N_556,In_4240,In_3499);
xnor U557 (N_557,In_141,In_2757);
or U558 (N_558,In_4375,In_1023);
nor U559 (N_559,In_1033,In_4230);
or U560 (N_560,In_2261,In_2351);
nand U561 (N_561,In_4797,In_4493);
xnor U562 (N_562,In_3709,In_4225);
and U563 (N_563,In_3114,In_2224);
and U564 (N_564,In_1530,In_2008);
xor U565 (N_565,In_3003,In_3570);
or U566 (N_566,In_204,In_2703);
or U567 (N_567,In_1074,In_4206);
xnor U568 (N_568,In_4369,In_2639);
and U569 (N_569,In_4174,In_4222);
nor U570 (N_570,In_4330,In_3952);
nand U571 (N_571,In_1115,In_2672);
or U572 (N_572,In_3617,In_1931);
and U573 (N_573,In_221,In_4841);
nor U574 (N_574,In_39,In_3406);
nand U575 (N_575,In_3634,In_292);
or U576 (N_576,In_4591,In_3463);
or U577 (N_577,In_3344,In_3211);
nand U578 (N_578,In_688,In_461);
nand U579 (N_579,In_978,In_944);
or U580 (N_580,In_1507,In_3133);
and U581 (N_581,In_1677,In_885);
or U582 (N_582,In_3063,In_1674);
nand U583 (N_583,In_2272,In_1446);
nand U584 (N_584,In_4333,In_1805);
nand U585 (N_585,In_317,In_2471);
nand U586 (N_586,In_4130,In_2640);
nor U587 (N_587,In_4316,In_1094);
nor U588 (N_588,In_821,In_3773);
xnor U589 (N_589,In_942,In_3741);
xor U590 (N_590,In_2304,In_4191);
and U591 (N_591,In_1624,In_651);
or U592 (N_592,In_3632,In_2934);
xor U593 (N_593,In_380,In_4108);
and U594 (N_594,In_2833,In_667);
nand U595 (N_595,In_3388,In_708);
and U596 (N_596,In_3062,In_2586);
nor U597 (N_597,In_496,In_971);
nand U598 (N_598,In_310,In_876);
xnor U599 (N_599,In_571,In_3724);
and U600 (N_600,In_2945,In_1132);
or U601 (N_601,In_2963,In_406);
xor U602 (N_602,In_3018,In_1274);
xor U603 (N_603,In_3552,In_2435);
nand U604 (N_604,In_3688,In_3262);
or U605 (N_605,In_1057,In_471);
and U606 (N_606,In_3213,In_1496);
nand U607 (N_607,In_195,In_2572);
xnor U608 (N_608,In_1959,In_3024);
nor U609 (N_609,In_2785,In_2483);
or U610 (N_610,In_1164,In_4824);
or U611 (N_611,In_1340,In_2719);
nor U612 (N_612,In_3457,In_1962);
xnor U613 (N_613,In_93,In_1213);
nor U614 (N_614,In_4119,In_711);
or U615 (N_615,In_4770,In_4893);
or U616 (N_616,In_4032,In_3157);
or U617 (N_617,In_1128,In_1725);
nand U618 (N_618,In_206,In_1454);
xnor U619 (N_619,In_1,In_3034);
or U620 (N_620,In_4871,In_2691);
nor U621 (N_621,In_3964,In_1472);
and U622 (N_622,In_2856,In_2205);
or U623 (N_623,In_634,In_1511);
xnor U624 (N_624,In_1126,In_698);
or U625 (N_625,In_1813,In_1474);
and U626 (N_626,In_4717,In_2206);
and U627 (N_627,In_1560,In_4818);
nand U628 (N_628,In_1248,In_775);
nor U629 (N_629,In_4784,In_2943);
and U630 (N_630,In_1660,In_2438);
and U631 (N_631,In_2907,In_2633);
and U632 (N_632,In_3771,In_3045);
or U633 (N_633,In_3393,In_4384);
nand U634 (N_634,In_3238,In_337);
nor U635 (N_635,In_3914,In_4782);
nor U636 (N_636,In_521,In_3289);
xnor U637 (N_637,In_3334,In_713);
nor U638 (N_638,In_420,In_3757);
nand U639 (N_639,In_4587,In_4833);
xor U640 (N_640,In_296,In_1055);
nand U641 (N_641,In_1591,In_4995);
nor U642 (N_642,In_1735,In_3258);
xnor U643 (N_643,In_16,In_2930);
nand U644 (N_644,In_2326,In_1119);
xor U645 (N_645,In_270,In_3145);
nand U646 (N_646,In_1438,In_4300);
nand U647 (N_647,In_803,In_2903);
xor U648 (N_648,In_2076,In_4128);
xnor U649 (N_649,In_2135,In_313);
nor U650 (N_650,In_1234,In_281);
nand U651 (N_651,In_444,In_823);
nor U652 (N_652,In_1535,In_332);
nor U653 (N_653,In_3464,In_2507);
xor U654 (N_654,In_3170,In_4874);
nor U655 (N_655,In_4336,In_3459);
xor U656 (N_656,In_2687,In_4036);
nand U657 (N_657,In_1697,In_1728);
nand U658 (N_658,In_2255,In_2734);
nor U659 (N_659,In_4069,In_335);
nand U660 (N_660,In_2484,In_1463);
nor U661 (N_661,In_3291,In_490);
nor U662 (N_662,In_2824,In_1706);
nand U663 (N_663,In_92,In_1698);
nand U664 (N_664,In_3610,In_3822);
xnor U665 (N_665,In_2497,In_4494);
nor U666 (N_666,In_3427,In_4123);
or U667 (N_667,In_2530,In_953);
and U668 (N_668,In_4742,In_1835);
and U669 (N_669,In_2127,In_365);
or U670 (N_670,In_4370,In_52);
nand U671 (N_671,In_3027,In_2125);
xnor U672 (N_672,In_702,In_2952);
or U673 (N_673,In_1997,In_4814);
or U674 (N_674,In_546,In_4887);
and U675 (N_675,In_585,In_3785);
nand U676 (N_676,In_3769,In_2955);
xnor U677 (N_677,In_1097,In_1895);
or U678 (N_678,In_1051,In_246);
or U679 (N_679,In_64,In_4414);
nor U680 (N_680,In_1110,In_1168);
and U681 (N_681,In_4630,In_2790);
nor U682 (N_682,In_1471,In_2917);
nor U683 (N_683,In_527,In_2114);
xnor U684 (N_684,In_1781,In_2327);
xnor U685 (N_685,In_4340,In_1477);
and U686 (N_686,In_1323,In_4332);
or U687 (N_687,In_1397,In_1688);
nor U688 (N_688,In_4320,In_2562);
and U689 (N_689,In_3135,In_248);
nand U690 (N_690,In_2960,In_2376);
xor U691 (N_691,In_2505,In_3364);
nand U692 (N_692,In_1631,In_3791);
and U693 (N_693,In_4495,In_4969);
and U694 (N_694,In_3281,In_366);
nor U695 (N_695,In_3301,In_2026);
and U696 (N_696,In_1802,In_4366);
and U697 (N_697,In_4999,In_286);
nand U698 (N_698,In_3257,In_3485);
xnor U699 (N_699,In_4823,In_259);
nor U700 (N_700,In_340,In_2225);
and U701 (N_701,In_4054,In_537);
and U702 (N_702,In_3180,In_1939);
nand U703 (N_703,In_4281,In_2231);
or U704 (N_704,In_2053,In_2863);
or U705 (N_705,In_22,In_4955);
or U706 (N_706,In_3566,In_1342);
xor U707 (N_707,In_2442,In_4895);
nand U708 (N_708,In_3105,In_3989);
xor U709 (N_709,In_3538,In_4650);
and U710 (N_710,In_1369,In_3728);
nand U711 (N_711,In_4996,In_4981);
and U712 (N_712,In_1460,In_3102);
nand U713 (N_713,In_1034,In_3328);
xnor U714 (N_714,In_3518,In_4220);
and U715 (N_715,In_2052,In_2230);
or U716 (N_716,In_4259,In_3483);
or U717 (N_717,In_1151,In_545);
or U718 (N_718,In_2522,In_345);
nor U719 (N_719,In_1876,In_758);
or U720 (N_720,In_3657,In_4175);
nand U721 (N_721,In_409,In_1778);
or U722 (N_722,In_1553,In_2569);
or U723 (N_723,In_2553,In_1402);
or U724 (N_724,In_3332,In_1226);
nor U725 (N_725,In_66,In_4939);
nor U726 (N_726,In_2084,In_4194);
and U727 (N_727,In_1385,In_3207);
and U728 (N_728,In_3013,In_3386);
nand U729 (N_729,In_595,In_3582);
xor U730 (N_730,In_511,In_1610);
nor U731 (N_731,In_2193,In_2064);
and U732 (N_732,In_145,In_959);
and U733 (N_733,In_3938,In_2993);
nand U734 (N_734,In_4925,In_1079);
nand U735 (N_735,In_1984,In_4573);
nand U736 (N_736,In_127,In_3241);
nor U737 (N_737,In_1744,In_1749);
nand U738 (N_738,In_2598,In_1825);
nor U739 (N_739,In_4345,In_3442);
nor U740 (N_740,In_4465,In_266);
nand U741 (N_741,In_3789,In_4744);
nor U742 (N_742,In_4299,In_131);
nor U743 (N_743,In_1038,In_1065);
nor U744 (N_744,In_301,In_890);
xor U745 (N_745,In_4909,In_4472);
nand U746 (N_746,In_2746,In_2737);
or U747 (N_747,In_3378,In_3048);
and U748 (N_748,In_3682,In_3793);
or U749 (N_749,In_3132,In_1035);
nand U750 (N_750,In_3642,In_2111);
xnor U751 (N_751,In_1058,In_1617);
nor U752 (N_752,In_388,In_4641);
nor U753 (N_753,In_2203,In_1943);
nor U754 (N_754,In_934,In_2765);
or U755 (N_755,In_272,In_1542);
xor U756 (N_756,In_455,In_1305);
nor U757 (N_757,In_3884,In_2625);
and U758 (N_758,In_737,In_3128);
nand U759 (N_759,In_983,In_4831);
nand U760 (N_760,In_2678,In_4951);
or U761 (N_761,In_3602,In_3370);
xor U762 (N_762,In_3508,In_4900);
xnor U763 (N_763,In_1275,In_1648);
or U764 (N_764,In_3270,In_1774);
nor U765 (N_765,In_4291,In_4415);
and U766 (N_766,In_913,In_3947);
nand U767 (N_767,In_4601,In_3723);
and U768 (N_768,In_1253,In_2309);
nand U769 (N_769,In_475,In_3054);
and U770 (N_770,In_1075,In_4718);
or U771 (N_771,In_600,In_3948);
xor U772 (N_772,In_2269,In_2029);
nor U773 (N_773,In_4456,In_1105);
nor U774 (N_774,In_889,In_3744);
nor U775 (N_775,In_2830,In_2913);
nor U776 (N_776,In_2928,In_4125);
nand U777 (N_777,In_291,In_1233);
and U778 (N_778,In_1319,In_3913);
nor U779 (N_779,In_1785,In_2339);
and U780 (N_780,In_4459,In_1347);
nand U781 (N_781,In_1264,In_901);
and U782 (N_782,In_368,In_2694);
or U783 (N_783,In_791,In_1447);
xnor U784 (N_784,In_1721,In_710);
or U785 (N_785,In_2227,In_1521);
and U786 (N_786,In_638,In_4124);
and U787 (N_787,In_4806,In_449);
nor U788 (N_788,In_37,In_829);
nand U789 (N_789,In_610,In_70);
nand U790 (N_790,In_3827,In_325);
nand U791 (N_791,In_2897,In_964);
xnor U792 (N_792,In_4688,In_3279);
or U793 (N_793,In_316,In_4399);
xnor U794 (N_794,In_3626,In_173);
or U795 (N_795,In_4896,In_2236);
nand U796 (N_796,In_2116,In_2417);
and U797 (N_797,In_2293,In_2618);
or U798 (N_798,In_2671,In_4634);
nand U799 (N_799,In_4949,In_3080);
or U800 (N_800,In_3455,In_2310);
and U801 (N_801,In_576,In_4452);
nand U802 (N_802,In_3292,In_2444);
or U803 (N_803,In_2876,In_4664);
and U804 (N_804,In_3417,In_3068);
and U805 (N_805,In_3647,In_3025);
nor U806 (N_806,In_835,In_3950);
and U807 (N_807,In_2994,In_2885);
nor U808 (N_808,In_1298,In_328);
or U809 (N_809,In_1606,In_946);
nand U810 (N_810,In_2972,In_1999);
nor U811 (N_811,In_3885,In_2433);
nand U812 (N_812,In_3749,In_3882);
xnor U813 (N_813,In_3535,In_4089);
nand U814 (N_814,In_3595,In_4071);
or U815 (N_815,In_1635,In_1723);
and U816 (N_816,In_3448,In_247);
or U817 (N_817,In_2220,In_1567);
xnor U818 (N_818,In_4976,In_2686);
nor U819 (N_819,In_3562,In_2519);
nand U820 (N_820,In_4460,In_3324);
nor U821 (N_821,In_275,In_724);
xnor U822 (N_822,In_487,In_3433);
and U823 (N_823,In_3221,In_3410);
nand U824 (N_824,In_2003,In_856);
xor U825 (N_825,In_2549,In_4524);
nand U826 (N_826,In_628,In_2921);
nand U827 (N_827,In_473,In_3823);
nor U828 (N_828,In_816,In_1738);
or U829 (N_829,In_2174,In_3187);
and U830 (N_830,In_2783,In_4577);
nand U831 (N_831,In_277,In_3085);
or U832 (N_832,In_3866,In_3217);
xnor U833 (N_833,In_3504,In_2285);
and U834 (N_834,In_1384,In_3890);
nand U835 (N_835,In_4308,In_3627);
or U836 (N_836,In_4433,In_383);
or U837 (N_837,In_4183,In_2741);
and U838 (N_838,In_2583,In_384);
xnor U839 (N_839,In_2486,In_3745);
xnor U840 (N_840,In_1975,In_41);
nor U841 (N_841,In_4391,In_4190);
nor U842 (N_842,In_1843,In_2982);
nor U843 (N_843,In_1951,In_4274);
or U844 (N_844,In_3795,In_3090);
xor U845 (N_845,In_4387,In_4484);
nand U846 (N_846,In_826,In_2767);
or U847 (N_847,In_1653,In_2154);
and U848 (N_848,In_2461,In_2229);
or U849 (N_849,In_78,In_69);
xor U850 (N_850,In_759,In_4203);
xnor U851 (N_851,In_2853,In_419);
nor U852 (N_852,In_1010,In_1961);
nand U853 (N_853,In_156,In_4544);
nor U854 (N_854,In_4132,In_798);
nand U855 (N_855,In_2181,In_2321);
nor U856 (N_856,In_222,In_820);
nor U857 (N_857,In_637,In_2717);
or U858 (N_858,In_3797,In_4971);
or U859 (N_859,In_2109,In_148);
nor U860 (N_860,In_3436,In_3396);
and U861 (N_861,In_2162,In_355);
and U862 (N_862,In_3942,In_2776);
or U863 (N_863,In_273,In_1968);
and U864 (N_864,In_3872,In_735);
nor U865 (N_865,In_4491,In_4905);
and U866 (N_866,In_2793,In_360);
or U867 (N_867,In_4815,In_305);
or U868 (N_868,In_2085,In_1767);
and U869 (N_869,In_3800,In_3561);
nand U870 (N_870,In_1562,In_2817);
and U871 (N_871,In_2131,In_1403);
xor U872 (N_872,In_1667,In_3750);
or U873 (N_873,In_4398,In_2933);
nor U874 (N_874,In_4500,In_1435);
or U875 (N_875,In_1566,In_1273);
nor U876 (N_876,In_1024,In_538);
nand U877 (N_877,In_117,In_3908);
or U878 (N_878,In_4822,In_2171);
xnor U879 (N_879,In_2126,In_1645);
xnor U880 (N_880,In_121,In_2715);
nor U881 (N_881,In_4978,In_3973);
and U882 (N_882,In_3231,In_2042);
xnor U883 (N_883,In_4439,In_3082);
xor U884 (N_884,In_2695,In_2742);
or U885 (N_885,In_929,In_3300);
xnor U886 (N_886,In_2768,In_3881);
or U887 (N_887,In_1649,In_1184);
or U888 (N_888,In_948,In_2893);
nor U889 (N_889,In_712,In_2434);
xnor U890 (N_890,In_3418,In_3000);
and U891 (N_891,In_3546,In_4618);
nand U892 (N_892,In_450,In_1020);
xnor U893 (N_893,In_1722,In_448);
nand U894 (N_894,In_3329,In_1390);
nand U895 (N_895,In_4694,In_4362);
nor U896 (N_896,In_4294,In_4935);
and U897 (N_897,In_4590,In_2118);
and U898 (N_898,In_754,In_806);
xnor U899 (N_899,In_2107,In_1816);
nor U900 (N_900,In_2550,In_4267);
nand U901 (N_901,In_3697,In_203);
nand U902 (N_902,In_4017,In_4803);
nand U903 (N_903,In_4973,In_1431);
nor U904 (N_904,In_2071,In_79);
xor U905 (N_905,In_2844,In_2846);
xnor U906 (N_906,In_2068,In_426);
nand U907 (N_907,In_4530,In_2896);
xor U908 (N_908,In_4171,In_4087);
or U909 (N_909,In_4648,In_2636);
nor U910 (N_910,In_4875,In_3568);
nand U911 (N_911,In_2337,In_4285);
nand U912 (N_912,In_762,In_1469);
nor U913 (N_913,In_2289,In_4152);
and U914 (N_914,In_1042,In_3687);
and U915 (N_915,In_149,In_2490);
nand U916 (N_916,In_351,In_4112);
nand U917 (N_917,In_4891,In_1215);
and U918 (N_918,In_4705,In_907);
or U919 (N_919,In_3895,In_2832);
or U920 (N_920,In_2954,In_2996);
xor U921 (N_921,In_2786,In_3342);
and U922 (N_922,In_1276,In_3591);
nand U923 (N_923,In_401,In_2465);
nand U924 (N_924,In_4726,In_2380);
or U925 (N_925,In_4056,In_4195);
nor U926 (N_926,In_4315,In_3668);
or U927 (N_927,In_2859,In_3830);
nand U928 (N_928,In_4503,In_2401);
and U929 (N_929,In_1107,In_588);
nor U930 (N_930,In_3821,In_3353);
nor U931 (N_931,In_2447,In_4563);
and U932 (N_932,In_3360,In_2506);
nor U933 (N_933,In_3017,In_998);
or U934 (N_934,In_56,In_3051);
xnor U935 (N_935,In_1245,In_90);
or U936 (N_936,In_987,In_4051);
or U937 (N_937,In_1352,In_3015);
nand U938 (N_938,In_2619,In_295);
and U939 (N_939,In_3202,In_4229);
nor U940 (N_940,In_866,In_3614);
nand U941 (N_941,In_3715,In_1699);
or U942 (N_942,In_282,In_1173);
or U943 (N_943,In_1181,In_878);
nand U944 (N_944,In_3944,In_1139);
and U945 (N_945,In_1819,In_1332);
or U946 (N_946,In_1363,In_3550);
xor U947 (N_947,In_3666,In_3044);
or U948 (N_948,In_3182,In_2459);
nor U949 (N_949,In_1296,In_1953);
xnor U950 (N_950,In_2355,In_1930);
or U951 (N_951,In_1592,In_3748);
and U952 (N_952,In_1572,In_269);
nand U953 (N_953,In_2059,In_2922);
xnor U954 (N_954,In_312,In_343);
nand U955 (N_955,In_3941,In_1516);
nor U956 (N_956,In_900,In_3401);
nor U957 (N_957,In_652,In_2239);
nor U958 (N_958,In_35,In_1561);
nand U959 (N_959,In_2189,In_569);
or U960 (N_960,In_4777,In_4853);
nand U961 (N_961,In_23,In_4970);
or U962 (N_962,In_3286,In_2493);
or U963 (N_963,In_1420,In_29);
nand U964 (N_964,In_1070,In_2704);
nand U965 (N_965,In_1710,In_2883);
or U966 (N_966,In_1327,In_1658);
and U967 (N_967,In_725,In_4886);
and U968 (N_968,In_4114,In_4262);
and U969 (N_969,In_4837,In_1501);
nand U970 (N_970,In_2218,In_624);
nor U971 (N_971,In_1601,In_3580);
or U972 (N_972,In_285,In_2840);
nand U973 (N_973,In_2589,In_4860);
and U974 (N_974,In_3010,In_3606);
nand U975 (N_975,In_4551,In_1001);
and U976 (N_976,In_4977,In_4352);
nor U977 (N_977,In_540,In_4117);
and U978 (N_978,In_1982,In_2167);
xor U979 (N_979,In_3738,In_4941);
or U980 (N_980,In_4034,In_4997);
xor U981 (N_981,In_4014,In_1784);
nand U982 (N_982,In_2190,In_1815);
or U983 (N_983,In_4432,In_4639);
and U984 (N_984,In_2408,In_568);
and U985 (N_985,In_2299,In_223);
nor U986 (N_986,In_1416,In_1091);
or U987 (N_987,In_3878,In_3225);
nor U988 (N_988,In_605,In_892);
nor U989 (N_989,In_185,In_3435);
nor U990 (N_990,In_1981,In_3708);
nand U991 (N_991,In_1796,In_167);
or U992 (N_992,In_491,In_3234);
xor U993 (N_993,In_2602,In_4790);
nand U994 (N_994,In_2137,In_1647);
nand U995 (N_995,In_2489,In_67);
xnor U996 (N_996,In_2191,In_2656);
nor U997 (N_997,In_2267,In_2020);
or U998 (N_998,In_2426,In_3042);
nor U999 (N_999,In_1159,In_996);
or U1000 (N_1000,In_1716,In_2390);
nor U1001 (N_1001,In_2811,In_4960);
nor U1002 (N_1002,In_2533,N_109);
or U1003 (N_1003,In_3107,In_815);
nand U1004 (N_1004,N_496,In_452);
xnor U1005 (N_1005,N_319,N_758);
nand U1006 (N_1006,In_2334,N_972);
and U1007 (N_1007,N_310,In_4141);
nor U1008 (N_1008,N_255,In_2271);
nor U1009 (N_1009,In_4443,In_377);
or U1010 (N_1010,N_898,In_4348);
nor U1011 (N_1011,In_2574,In_3753);
and U1012 (N_1012,N_564,In_1900);
nor U1013 (N_1013,In_2975,In_3840);
xnor U1014 (N_1014,In_2542,In_957);
and U1015 (N_1015,In_4799,In_1772);
xor U1016 (N_1016,In_4450,In_4745);
nor U1017 (N_1017,N_962,In_1426);
and U1018 (N_1018,N_583,In_4740);
nor U1019 (N_1019,In_565,In_2738);
or U1020 (N_1020,In_1071,In_3590);
and U1021 (N_1021,N_172,N_148);
nor U1022 (N_1022,N_276,In_1133);
and U1023 (N_1023,N_949,In_3308);
nor U1024 (N_1024,In_217,In_580);
nor U1025 (N_1025,N_194,N_854);
nand U1026 (N_1026,N_469,In_2521);
nand U1027 (N_1027,In_1138,In_1493);
xnor U1028 (N_1028,In_1905,In_767);
or U1029 (N_1029,In_831,In_2492);
or U1030 (N_1030,N_217,In_4628);
nand U1031 (N_1031,In_2027,In_454);
xor U1032 (N_1032,N_994,In_1800);
nor U1033 (N_1033,In_2128,N_668);
nand U1034 (N_1034,In_445,In_3782);
nand U1035 (N_1035,N_685,In_3239);
xnor U1036 (N_1036,N_48,N_825);
xnor U1037 (N_1037,In_715,In_1626);
nor U1038 (N_1038,In_4785,In_2396);
and U1039 (N_1039,In_3553,In_3375);
xnor U1040 (N_1040,In_3129,N_926);
nand U1041 (N_1041,In_2062,In_3060);
xnor U1042 (N_1042,In_1089,N_42);
nor U1043 (N_1043,N_231,N_902);
nand U1044 (N_1044,In_4793,In_1896);
nand U1045 (N_1045,In_3658,In_2663);
and U1046 (N_1046,In_549,In_4817);
or U1047 (N_1047,N_776,In_3695);
nand U1048 (N_1048,In_3108,N_22);
xnor U1049 (N_1049,In_3479,In_1780);
and U1050 (N_1050,In_4957,In_107);
nand U1051 (N_1051,N_135,In_1714);
nor U1052 (N_1052,N_794,N_99);
nor U1053 (N_1053,In_3311,N_66);
or U1054 (N_1054,In_2939,In_2415);
or U1055 (N_1055,N_763,In_2);
or U1056 (N_1056,N_137,In_2709);
nor U1057 (N_1057,In_4676,In_2032);
xnor U1058 (N_1058,In_726,In_2005);
and U1059 (N_1059,In_4928,In_3223);
and U1060 (N_1060,In_1795,In_4055);
nand U1061 (N_1061,In_4116,In_772);
nand U1062 (N_1062,N_739,In_1466);
nand U1063 (N_1063,In_1540,N_641);
nand U1064 (N_1064,In_896,In_1803);
nor U1065 (N_1065,In_2038,In_1763);
and U1066 (N_1066,In_4681,N_238);
or U1067 (N_1067,In_3460,In_3327);
or U1068 (N_1068,In_1944,In_3925);
nor U1069 (N_1069,In_1155,In_1595);
nor U1070 (N_1070,In_2308,In_2556);
and U1071 (N_1071,In_1462,In_2564);
and U1072 (N_1072,N_486,In_2312);
nor U1073 (N_1073,In_849,In_1003);
or U1074 (N_1074,In_1320,In_3842);
nand U1075 (N_1075,In_751,In_3680);
nand U1076 (N_1076,In_3578,In_36);
nor U1077 (N_1077,N_771,In_1373);
or U1078 (N_1078,In_4075,N_853);
and U1079 (N_1079,N_872,N_702);
and U1080 (N_1080,In_4143,In_1545);
nor U1081 (N_1081,N_807,In_592);
xnor U1082 (N_1082,N_485,N_600);
and U1083 (N_1083,N_932,In_2823);
xor U1084 (N_1084,N_162,In_32);
or U1085 (N_1085,N_330,In_4733);
xor U1086 (N_1086,In_3955,In_1427);
nor U1087 (N_1087,In_3557,N_611);
or U1088 (N_1088,In_1523,In_3077);
nand U1089 (N_1089,In_4626,N_81);
xnor U1090 (N_1090,N_752,In_2383);
xor U1091 (N_1091,In_660,In_1297);
nor U1092 (N_1092,In_1916,In_2072);
xnor U1093 (N_1093,In_3859,N_458);
or U1094 (N_1094,In_395,In_4355);
nand U1095 (N_1095,In_785,In_113);
or U1096 (N_1096,In_46,In_4848);
nor U1097 (N_1097,N_843,In_4359);
nor U1098 (N_1098,In_2983,N_489);
xor U1099 (N_1099,In_1252,In_1957);
and U1100 (N_1100,In_886,In_258);
xor U1101 (N_1101,N_419,In_1718);
nor U1102 (N_1102,In_4586,In_2002);
and U1103 (N_1103,In_1027,N_691);
and U1104 (N_1104,In_165,In_4791);
xor U1105 (N_1105,In_2649,In_4912);
nor U1106 (N_1106,N_785,In_3967);
xnor U1107 (N_1107,In_1712,In_2906);
or U1108 (N_1108,In_100,In_616);
and U1109 (N_1109,N_317,In_2100);
nand U1110 (N_1110,In_3780,N_287);
and U1111 (N_1111,In_19,N_214);
xnor U1112 (N_1112,In_4678,In_233);
and U1113 (N_1113,In_2264,N_335);
and U1114 (N_1114,In_1081,N_415);
xnor U1115 (N_1115,In_609,In_3755);
nand U1116 (N_1116,In_869,N_840);
and U1117 (N_1117,In_2585,In_2936);
nand U1118 (N_1118,In_2539,In_3184);
nand U1119 (N_1119,In_968,N_26);
or U1120 (N_1120,In_459,N_688);
nand U1121 (N_1121,In_2512,In_3677);
and U1122 (N_1122,N_713,In_1727);
nor U1123 (N_1123,In_709,In_3008);
nor U1124 (N_1124,In_2657,In_746);
xnor U1125 (N_1125,In_2212,In_749);
xor U1126 (N_1126,In_2777,In_4514);
or U1127 (N_1127,N_182,N_340);
nand U1128 (N_1128,In_2065,N_211);
xnor U1129 (N_1129,In_1799,In_3275);
xor U1130 (N_1130,In_2196,In_2894);
nand U1131 (N_1131,In_3377,In_3936);
xor U1132 (N_1132,In_3998,N_351);
or U1133 (N_1133,In_253,In_2892);
and U1134 (N_1134,In_705,In_4938);
nand U1135 (N_1135,N_607,In_479);
xor U1136 (N_1136,In_922,In_1183);
xnor U1137 (N_1137,In_1536,In_2361);
or U1138 (N_1138,N_555,N_1);
and U1139 (N_1139,In_1787,N_886);
nor U1140 (N_1140,In_1786,In_4659);
nor U1141 (N_1141,N_422,In_824);
nand U1142 (N_1142,In_2617,In_3242);
xor U1143 (N_1143,In_3101,In_499);
nand U1144 (N_1144,In_771,In_367);
and U1145 (N_1145,In_3794,In_2404);
nand U1146 (N_1146,N_538,N_235);
and U1147 (N_1147,In_779,N_116);
and U1148 (N_1148,In_3644,In_840);
or U1149 (N_1149,In_3686,In_3011);
nand U1150 (N_1150,In_4834,In_4736);
or U1151 (N_1151,In_1281,In_3005);
nor U1152 (N_1152,In_4673,In_1284);
or U1153 (N_1153,In_4892,In_1879);
nor U1154 (N_1154,In_723,In_1195);
and U1155 (N_1155,In_1212,In_1594);
nor U1156 (N_1156,In_3943,In_3169);
xor U1157 (N_1157,N_323,In_2566);
xnor U1158 (N_1158,In_2399,N_759);
or U1159 (N_1159,In_1985,In_1016);
or U1160 (N_1160,In_3839,In_4558);
nand U1161 (N_1161,In_4418,In_3423);
or U1162 (N_1162,In_3706,In_1414);
nand U1163 (N_1163,In_3369,In_790);
nor U1164 (N_1164,In_2733,In_1600);
or U1165 (N_1165,In_171,N_409);
and U1166 (N_1166,In_2121,N_637);
or U1167 (N_1167,In_2510,In_2772);
xor U1168 (N_1168,In_4827,In_3932);
or U1169 (N_1169,N_325,In_699);
nand U1170 (N_1170,N_755,N_876);
or U1171 (N_1171,In_1265,In_4135);
xor U1172 (N_1172,In_3316,In_1457);
nand U1173 (N_1173,In_2213,In_4080);
nand U1174 (N_1174,In_2888,In_4506);
and U1175 (N_1175,In_4737,In_4073);
or U1176 (N_1176,In_2315,N_374);
or U1177 (N_1177,N_855,In_1246);
or U1178 (N_1178,In_872,In_4368);
nand U1179 (N_1179,In_2476,In_2828);
xnor U1180 (N_1180,In_1742,In_2529);
or U1181 (N_1181,In_4070,In_3155);
xnor U1182 (N_1182,N_865,In_3422);
nand U1183 (N_1183,In_4947,In_1908);
and U1184 (N_1184,In_2697,N_121);
nand U1185 (N_1185,N_16,In_261);
or U1186 (N_1186,In_579,In_581);
nand U1187 (N_1187,In_4095,N_880);
or U1188 (N_1188,In_550,In_804);
or U1189 (N_1189,N_944,N_436);
or U1190 (N_1190,In_1381,N_849);
or U1191 (N_1191,N_535,N_603);
and U1192 (N_1192,In_3404,In_4035);
nand U1193 (N_1193,In_4166,In_3006);
or U1194 (N_1194,N_937,N_267);
nand U1195 (N_1195,In_1656,In_1952);
xnor U1196 (N_1196,In_1833,N_64);
nand U1197 (N_1197,In_2557,In_4497);
nor U1198 (N_1198,In_3445,N_184);
nor U1199 (N_1199,In_3496,In_2041);
and U1200 (N_1200,In_1066,In_2096);
or U1201 (N_1201,In_2172,N_515);
nand U1202 (N_1202,In_4596,In_3509);
nand U1203 (N_1203,In_923,In_4734);
and U1204 (N_1204,In_4691,In_111);
nand U1205 (N_1205,In_3766,In_1222);
nor U1206 (N_1206,In_518,N_630);
nor U1207 (N_1207,In_1764,In_1148);
nor U1208 (N_1208,In_2012,In_4913);
or U1209 (N_1209,In_1559,N_711);
xnor U1210 (N_1210,In_4487,In_45);
nand U1211 (N_1211,In_398,In_3227);
and U1212 (N_1212,In_4325,In_3273);
nor U1213 (N_1213,In_2947,In_4870);
and U1214 (N_1214,In_2430,In_4162);
nor U1215 (N_1215,In_2132,In_1558);
xnor U1216 (N_1216,N_553,N_101);
and U1217 (N_1217,In_2712,In_153);
and U1218 (N_1218,In_4772,N_952);
or U1219 (N_1219,N_119,In_3267);
nor U1220 (N_1220,In_4084,N_207);
or U1221 (N_1221,N_918,N_257);
nor U1222 (N_1222,N_10,In_4505);
or U1223 (N_1223,In_4567,N_110);
xor U1224 (N_1224,In_4280,N_656);
and U1225 (N_1225,In_639,In_2620);
xor U1226 (N_1226,In_2520,In_3110);
nand U1227 (N_1227,In_2517,In_3599);
nor U1228 (N_1228,In_4523,N_501);
xor U1229 (N_1229,In_4496,In_3315);
and U1230 (N_1230,N_719,In_3091);
nand U1231 (N_1231,In_1227,N_951);
nor U1232 (N_1232,In_1823,In_3648);
nand U1233 (N_1233,In_4959,N_992);
xnor U1234 (N_1234,In_3854,In_4074);
or U1235 (N_1235,N_869,In_2199);
xnor U1236 (N_1236,In_3248,In_4319);
nand U1237 (N_1237,In_4293,N_585);
nor U1238 (N_1238,In_1666,N_189);
nor U1239 (N_1239,In_274,N_192);
nor U1240 (N_1240,In_2560,In_2744);
nand U1241 (N_1241,In_2023,N_259);
nand U1242 (N_1242,N_655,In_4948);
and U1243 (N_1243,In_3892,In_402);
or U1244 (N_1244,In_947,In_3035);
or U1245 (N_1245,In_4645,In_1210);
and U1246 (N_1246,N_480,N_910);
or U1247 (N_1247,In_2460,In_2439);
or U1248 (N_1248,In_17,In_4536);
nand U1249 (N_1249,In_4595,N_909);
and U1250 (N_1250,In_4623,In_2855);
nand U1251 (N_1251,N_82,In_2049);
and U1252 (N_1252,N_722,In_897);
nor U1253 (N_1253,In_2487,N_834);
xnor U1254 (N_1254,In_4868,In_1807);
xnor U1255 (N_1255,In_3120,In_2328);
and U1256 (N_1256,N_970,In_3734);
nor U1257 (N_1257,In_2347,In_4621);
xnor U1258 (N_1258,N_144,In_677);
nor U1259 (N_1259,In_1826,In_341);
and U1260 (N_1260,In_2735,In_423);
and U1261 (N_1261,In_674,In_2388);
nand U1262 (N_1262,In_2854,In_4106);
and U1263 (N_1263,In_642,In_1520);
and U1264 (N_1264,N_983,In_1759);
and U1265 (N_1265,In_564,In_662);
and U1266 (N_1266,In_20,In_1846);
or U1267 (N_1267,N_912,In_1490);
xnor U1268 (N_1268,N_998,In_1809);
xnor U1269 (N_1269,In_4338,In_231);
nor U1270 (N_1270,In_918,N_930);
or U1271 (N_1271,N_871,In_1740);
nand U1272 (N_1272,In_4091,In_3907);
nor U1273 (N_1273,In_220,In_3871);
and U1274 (N_1274,In_268,N_499);
and U1275 (N_1275,In_410,N_154);
and U1276 (N_1276,N_165,N_979);
and U1277 (N_1277,In_2575,In_2437);
and U1278 (N_1278,N_273,In_1568);
or U1279 (N_1279,N_468,In_3860);
nand U1280 (N_1280,In_3514,N_220);
or U1281 (N_1281,In_3394,In_739);
xor U1282 (N_1282,In_4061,In_3325);
and U1283 (N_1283,In_1505,In_3229);
or U1284 (N_1284,In_1349,In_4612);
xnor U1285 (N_1285,In_4266,In_4850);
or U1286 (N_1286,N_44,In_1410);
or U1287 (N_1287,In_364,In_2297);
nor U1288 (N_1288,N_531,In_2325);
nor U1289 (N_1289,In_1878,In_1707);
and U1290 (N_1290,N_173,In_3743);
xnor U1291 (N_1291,N_728,In_1949);
and U1292 (N_1292,In_4318,In_2215);
nor U1293 (N_1293,In_528,In_3043);
and U1294 (N_1294,N_393,In_234);
nor U1295 (N_1295,N_751,In_2816);
nand U1296 (N_1296,In_2369,In_2838);
nor U1297 (N_1297,In_3587,N_128);
xnor U1298 (N_1298,N_249,In_1160);
nor U1299 (N_1299,In_1979,In_951);
and U1300 (N_1300,In_2466,N_223);
or U1301 (N_1301,In_3336,In_1041);
xor U1302 (N_1302,N_536,In_1092);
xnor U1303 (N_1303,In_3343,In_4097);
xnor U1304 (N_1304,N_559,In_2362);
nand U1305 (N_1305,In_924,N_612);
nand U1306 (N_1306,In_4142,In_1845);
xor U1307 (N_1307,In_2961,In_1554);
nand U1308 (N_1308,In_768,In_851);
nor U1309 (N_1309,In_2728,In_1456);
xor U1310 (N_1310,In_1762,In_1495);
and U1311 (N_1311,N_820,In_4189);
or U1312 (N_1312,In_4327,N_974);
nand U1313 (N_1313,In_3685,In_4090);
xnor U1314 (N_1314,In_3037,In_2762);
nand U1315 (N_1315,In_3733,N_247);
and U1316 (N_1316,N_638,In_2480);
nand U1317 (N_1317,In_136,In_4652);
or U1318 (N_1318,N_17,In_76);
or U1319 (N_1319,N_30,In_3195);
nor U1320 (N_1320,In_2605,In_318);
or U1321 (N_1321,In_928,In_2058);
or U1322 (N_1322,In_4674,In_2606);
or U1323 (N_1323,In_309,In_1443);
nor U1324 (N_1324,In_2142,In_1117);
xnor U1325 (N_1325,In_1059,N_829);
xnor U1326 (N_1326,In_4987,N_753);
nand U1327 (N_1327,In_4696,In_175);
and U1328 (N_1328,In_2152,N_68);
and U1329 (N_1329,In_458,In_3729);
nand U1330 (N_1330,In_2648,In_861);
or U1331 (N_1331,N_34,In_1376);
nand U1332 (N_1332,In_2094,N_471);
nor U1333 (N_1333,In_3494,In_3021);
nor U1334 (N_1334,In_520,In_682);
nand U1335 (N_1335,In_1628,In_3760);
xnor U1336 (N_1336,N_804,In_3206);
and U1337 (N_1337,In_2097,In_2528);
nor U1338 (N_1338,In_865,In_4477);
xnor U1339 (N_1339,In_2788,In_2867);
nand U1340 (N_1340,In_4640,In_1143);
and U1341 (N_1341,In_4578,In_2458);
or U1342 (N_1342,In_3412,In_1589);
or U1343 (N_1343,N_428,In_3551);
or U1344 (N_1344,In_3506,In_1834);
xnor U1345 (N_1345,In_502,In_1546);
and U1346 (N_1346,In_1651,N_326);
or U1347 (N_1347,In_3629,In_2406);
or U1348 (N_1348,In_788,In_2103);
xor U1349 (N_1349,N_460,In_2587);
and U1350 (N_1350,In_3437,In_1485);
nor U1351 (N_1351,In_2822,In_363);
nor U1352 (N_1352,In_2413,In_2821);
nand U1353 (N_1353,N_265,In_3598);
or U1354 (N_1354,In_1334,N_270);
xor U1355 (N_1355,N_47,In_1928);
or U1356 (N_1356,In_1387,N_355);
xor U1357 (N_1357,In_87,In_3828);
nor U1358 (N_1358,In_2797,In_4088);
nor U1359 (N_1359,In_2769,In_4188);
xnor U1360 (N_1360,In_3713,In_833);
and U1361 (N_1361,In_478,In_4205);
nand U1362 (N_1362,In_3559,In_962);
xnor U1363 (N_1363,N_4,In_4656);
nand U1364 (N_1364,N_837,In_4732);
and U1365 (N_1365,In_1818,In_3305);
nor U1366 (N_1366,In_124,In_1702);
or U1367 (N_1367,In_2428,In_58);
nand U1368 (N_1368,In_2714,In_2083);
nor U1369 (N_1369,In_2494,N_730);
or U1370 (N_1370,In_2294,In_308);
and U1371 (N_1371,In_311,In_3920);
and U1372 (N_1372,N_159,In_229);
nor U1373 (N_1373,N_494,In_1963);
xor U1374 (N_1374,In_4788,In_3466);
and U1375 (N_1375,In_1859,N_39);
nor U1376 (N_1376,In_3153,In_4765);
or U1377 (N_1377,In_1095,N_161);
nor U1378 (N_1378,In_435,N_108);
and U1379 (N_1379,In_601,N_961);
or U1380 (N_1380,N_620,N_93);
or U1381 (N_1381,In_404,In_1537);
or U1382 (N_1382,In_40,N_640);
nand U1383 (N_1383,In_4929,N_404);
nor U1384 (N_1384,In_3067,N_497);
and U1385 (N_1385,In_4219,In_152);
and U1386 (N_1386,In_3888,N_580);
and U1387 (N_1387,In_4471,In_4617);
and U1388 (N_1388,N_367,In_0);
or U1389 (N_1389,In_1500,In_4424);
and U1390 (N_1390,In_1641,In_2086);
or U1391 (N_1391,In_4922,In_1394);
and U1392 (N_1392,In_3191,In_202);
and U1393 (N_1393,In_1122,N_975);
nor U1394 (N_1394,In_1263,N_87);
xnor U1395 (N_1395,In_986,In_2570);
or U1396 (N_1396,In_3124,In_50);
and U1397 (N_1397,In_3767,In_2021);
and U1398 (N_1398,In_1578,In_1353);
nand U1399 (N_1399,In_3670,In_1022);
and U1400 (N_1400,N_847,N_901);
nor U1401 (N_1401,In_1946,In_3517);
or U1402 (N_1402,In_4677,In_4520);
or U1403 (N_1403,In_3462,In_4344);
nor U1404 (N_1404,In_2621,In_4877);
xor U1405 (N_1405,In_3023,In_2165);
or U1406 (N_1406,In_3893,In_2707);
nand U1407 (N_1407,In_1061,In_800);
and U1408 (N_1408,In_4598,In_134);
and U1409 (N_1409,In_2938,In_2000);
or U1410 (N_1410,In_2400,In_3376);
or U1411 (N_1411,N_157,In_2185);
xnor U1412 (N_1412,In_1927,In_2976);
and U1413 (N_1413,In_960,N_353);
or U1414 (N_1414,In_3178,N_987);
xor U1415 (N_1415,In_3458,In_795);
and U1416 (N_1416,In_421,N_24);
and U1417 (N_1417,In_386,N_248);
xor U1418 (N_1418,In_2391,In_4431);
and U1419 (N_1419,In_717,In_442);
nand U1420 (N_1420,In_4816,In_1633);
or U1421 (N_1421,In_4158,N_0);
or U1422 (N_1422,In_1539,In_2449);
nor U1423 (N_1423,N_618,N_348);
or U1424 (N_1424,In_63,N_118);
nand U1425 (N_1425,In_1468,N_58);
or U1426 (N_1426,In_4003,In_2204);
nand U1427 (N_1427,In_915,In_4475);
nor U1428 (N_1428,In_553,In_1661);
xor U1429 (N_1429,N_327,In_3957);
or U1430 (N_1430,In_1359,In_3285);
or U1431 (N_1431,N_437,In_11);
and U1432 (N_1432,In_4488,In_2847);
and U1433 (N_1433,In_2848,In_2752);
nor U1434 (N_1434,In_4654,In_4198);
nor U1435 (N_1435,N_617,In_60);
or U1436 (N_1436,N_167,In_1670);
xor U1437 (N_1437,N_948,In_2113);
xor U1438 (N_1438,In_4651,In_1627);
nand U1439 (N_1439,In_297,In_3420);
nand U1440 (N_1440,N_286,In_3237);
nand U1441 (N_1441,N_850,In_4243);
nand U1442 (N_1442,In_2291,In_2501);
and U1443 (N_1443,In_1971,N_729);
xnor U1444 (N_1444,In_2448,In_1991);
xor U1445 (N_1445,N_438,In_4233);
or U1446 (N_1446,In_1343,N_268);
nor U1447 (N_1447,In_2523,N_251);
and U1448 (N_1448,N_112,In_3317);
nor U1449 (N_1449,N_764,In_394);
nor U1450 (N_1450,In_4550,N_520);
nor U1451 (N_1451,N_36,In_497);
nand U1452 (N_1452,In_2313,N_177);
nand U1453 (N_1453,In_105,In_484);
or U1454 (N_1454,In_2680,In_2644);
xnor U1455 (N_1455,In_2965,In_3219);
nor U1456 (N_1456,N_940,N_307);
nand U1457 (N_1457,In_1973,In_1577);
nand U1458 (N_1458,In_3787,In_1804);
and U1459 (N_1459,In_2890,N_543);
or U1460 (N_1460,N_997,In_2184);
or U1461 (N_1461,In_950,In_965);
or U1462 (N_1462,N_5,In_3075);
or U1463 (N_1463,In_389,In_4979);
nand U1464 (N_1464,In_1849,In_2044);
nor U1465 (N_1465,In_2254,N_421);
nand U1466 (N_1466,In_354,In_3995);
and U1467 (N_1467,In_2546,N_838);
xor U1468 (N_1468,In_199,In_213);
nand U1469 (N_1469,In_4986,In_3331);
nor U1470 (N_1470,N_338,N_693);
xor U1471 (N_1471,N_204,In_4921);
or U1472 (N_1472,In_4239,In_4786);
nand U1473 (N_1473,N_94,In_4000);
nand U1474 (N_1474,In_1824,In_582);
nor U1475 (N_1475,N_19,In_283);
and U1476 (N_1476,In_1650,N_703);
nor U1477 (N_1477,In_844,In_4482);
or U1478 (N_1478,In_3399,In_3620);
and U1479 (N_1479,In_4139,N_405);
and U1480 (N_1480,In_3302,In_1890);
and U1481 (N_1481,In_4031,N_245);
xor U1482 (N_1482,In_864,In_3838);
or U1483 (N_1483,N_619,In_2036);
or U1484 (N_1484,N_433,In_15);
or U1485 (N_1485,In_3624,In_640);
nor U1486 (N_1486,In_4322,In_4727);
or U1487 (N_1487,N_462,N_929);
nor U1488 (N_1488,In_4521,In_2001);
nand U1489 (N_1489,In_2054,N_899);
xor U1490 (N_1490,In_3826,In_4374);
nand U1491 (N_1491,In_925,In_3549);
and U1492 (N_1492,In_1856,In_25);
nand U1493 (N_1493,N_989,N_183);
nor U1494 (N_1494,In_4662,In_2098);
xor U1495 (N_1495,In_4993,In_4869);
or U1496 (N_1496,In_2684,N_263);
nor U1497 (N_1497,In_3350,In_431);
and U1498 (N_1498,N_891,N_6);
nand U1499 (N_1499,In_139,In_4751);
and U1500 (N_1500,In_370,In_119);
or U1501 (N_1501,In_2968,In_210);
xor U1502 (N_1502,In_2092,N_801);
xor U1503 (N_1503,In_4005,N_525);
or U1504 (N_1504,In_4241,In_1142);
or U1505 (N_1505,N_229,In_4270);
or U1506 (N_1506,N_188,In_1370);
or U1507 (N_1507,N_567,In_3643);
nand U1508 (N_1508,In_1322,N_492);
xnor U1509 (N_1509,In_3698,In_2763);
xnor U1510 (N_1510,In_4151,In_3522);
xnor U1511 (N_1511,N_963,In_215);
and U1512 (N_1512,In_4936,In_3764);
and U1513 (N_1513,In_125,In_543);
or U1514 (N_1514,N_925,In_227);
or U1515 (N_1515,In_2292,In_921);
nor U1516 (N_1516,In_4378,In_3385);
xnor U1517 (N_1517,In_263,In_1169);
nor U1518 (N_1518,In_1956,In_3649);
nand U1519 (N_1519,In_1048,N_379);
nand U1520 (N_1520,In_4085,In_926);
xnor U1521 (N_1521,In_3387,In_2470);
nor U1522 (N_1522,In_570,In_4682);
and U1523 (N_1523,In_4295,N_572);
nand U1524 (N_1524,N_508,In_3122);
nand U1525 (N_1525,N_599,In_2970);
and U1526 (N_1526,In_3146,In_1430);
xor U1527 (N_1527,In_2354,N_261);
nand U1528 (N_1528,In_1841,In_2563);
nor U1529 (N_1529,In_666,In_4045);
nand U1530 (N_1530,In_3278,In_2645);
nand U1531 (N_1531,In_2175,N_361);
and U1532 (N_1532,In_4256,In_4989);
xor U1533 (N_1533,N_556,N_960);
nor U1534 (N_1534,In_955,In_1333);
and U1535 (N_1535,In_4774,In_3103);
and U1536 (N_1536,In_1844,In_838);
nand U1537 (N_1537,In_3357,In_4018);
xnor U1538 (N_1538,In_3604,N_227);
and U1539 (N_1539,In_2238,In_4100);
nand U1540 (N_1540,N_800,In_4109);
xnor U1541 (N_1541,In_376,In_205);
nor U1542 (N_1542,N_122,In_4988);
and U1543 (N_1543,N_76,In_1044);
and U1544 (N_1544,In_1837,In_2792);
or U1545 (N_1545,In_278,N_455);
or U1546 (N_1546,N_791,In_4667);
and U1547 (N_1547,In_2145,N_453);
nor U1548 (N_1548,In_3710,In_2898);
nor U1549 (N_1549,In_1705,In_2268);
nand U1550 (N_1550,N_674,In_68);
xnor U1551 (N_1551,N_608,In_3162);
and U1552 (N_1552,In_2187,In_4529);
xnor U1553 (N_1553,In_2421,N_79);
and U1554 (N_1554,In_4542,In_3486);
or U1555 (N_1555,In_4455,In_574);
xor U1556 (N_1556,In_1711,In_4110);
xor U1557 (N_1557,N_714,In_4180);
nor U1558 (N_1558,In_3031,In_920);
and U1559 (N_1559,In_2284,In_2858);
or U1560 (N_1560,In_1851,In_3519);
nor U1561 (N_1561,N_848,In_2775);
nand U1562 (N_1562,In_2659,In_1237);
xor U1563 (N_1563,In_3811,In_3089);
or U1564 (N_1564,In_567,In_627);
xnor U1565 (N_1565,In_1270,N_881);
or U1566 (N_1566,In_4029,N_105);
or U1567 (N_1567,In_3736,N_80);
xnor U1568 (N_1568,In_1277,In_3030);
nand U1569 (N_1569,In_2242,N_505);
nand U1570 (N_1570,In_4828,In_4794);
nor U1571 (N_1571,N_735,In_2022);
nand U1572 (N_1572,N_448,In_4917);
nor U1573 (N_1573,In_4287,N_170);
nand U1574 (N_1574,In_2756,In_2632);
nand U1575 (N_1575,In_522,In_625);
nand U1576 (N_1576,In_2845,In_2690);
nand U1577 (N_1577,In_4209,In_4273);
xnor U1578 (N_1578,In_3368,In_908);
nor U1579 (N_1579,In_2584,In_3527);
and U1580 (N_1580,In_3119,In_3992);
xnor U1581 (N_1581,In_4010,In_4944);
or U1582 (N_1582,In_4196,In_2099);
xor U1583 (N_1583,In_4063,In_2407);
or U1584 (N_1584,In_3997,In_1219);
xnor U1585 (N_1585,In_2527,In_2979);
or U1586 (N_1586,In_1049,In_3805);
and U1587 (N_1587,In_2360,N_558);
xor U1588 (N_1588,In_780,In_3073);
or U1589 (N_1589,N_811,In_1502);
nand U1590 (N_1590,In_2814,In_2252);
or U1591 (N_1591,In_3130,In_4615);
xor U1592 (N_1592,N_254,In_2477);
or U1593 (N_1593,In_101,In_2927);
nor U1594 (N_1594,In_339,In_3739);
nand U1595 (N_1595,In_413,In_2011);
or U1596 (N_1596,In_1260,In_1732);
nand U1597 (N_1597,N_795,N_938);
or U1598 (N_1598,In_2834,In_2677);
and U1599 (N_1599,In_4436,In_2631);
or U1600 (N_1600,N_554,In_3530);
or U1601 (N_1601,N_301,In_590);
or U1602 (N_1602,In_671,N_793);
nor U1603 (N_1603,In_2499,In_1367);
nand U1604 (N_1604,N_152,In_1919);
nand U1605 (N_1605,In_619,In_3946);
nand U1606 (N_1606,In_2429,N_482);
and U1607 (N_1607,In_4341,In_3808);
xor U1608 (N_1608,In_3516,In_3574);
nand U1609 (N_1609,In_721,In_327);
nand U1610 (N_1610,In_1285,In_4760);
and U1611 (N_1611,In_4600,In_3352);
nor U1612 (N_1612,In_575,N_953);
xor U1613 (N_1613,In_1812,In_4416);
xnor U1614 (N_1614,N_986,N_343);
nand U1615 (N_1615,In_425,In_4624);
xnor U1616 (N_1616,In_110,In_1556);
or U1617 (N_1617,In_2160,N_230);
and U1618 (N_1618,In_1172,In_359);
xor U1619 (N_1619,In_2305,In_3166);
and U1620 (N_1620,In_1354,In_3214);
nand U1621 (N_1621,In_2359,In_1372);
nand U1622 (N_1622,In_2706,In_209);
xnor U1623 (N_1623,In_818,In_3934);
or U1624 (N_1624,N_54,N_980);
nand U1625 (N_1625,N_858,In_2214);
nand U1626 (N_1626,In_385,N_84);
nand U1627 (N_1627,N_491,In_242);
xnor U1628 (N_1628,In_3465,N_978);
xor U1629 (N_1629,In_4526,In_769);
xor U1630 (N_1630,In_2281,N_606);
and U1631 (N_1631,In_1203,In_2073);
nand U1632 (N_1632,In_2723,In_992);
nand U1633 (N_1633,In_265,In_1642);
and U1634 (N_1634,In_3503,In_28);
nor U1635 (N_1635,In_4,In_4689);
xnor U1636 (N_1636,N_571,In_198);
and U1637 (N_1637,In_3026,N_196);
nor U1638 (N_1638,N_747,In_4911);
xor U1639 (N_1639,In_2616,In_1067);
or U1640 (N_1640,In_3704,In_2643);
or U1641 (N_1641,In_3990,In_3185);
nand U1642 (N_1642,In_658,In_2080);
nand U1643 (N_1643,N_33,In_3487);
nand U1644 (N_1644,In_2718,In_777);
nand U1645 (N_1645,In_4902,In_1700);
nand U1646 (N_1646,In_1639,In_4217);
or U1647 (N_1647,In_3160,In_656);
and U1648 (N_1648,N_864,N_783);
and U1649 (N_1649,In_2568,In_1131);
nor U1650 (N_1650,In_3307,In_1607);
xnor U1651 (N_1651,In_4882,In_770);
and U1652 (N_1652,N_675,In_177);
nand U1653 (N_1653,In_573,In_4901);
nand U1654 (N_1654,In_822,In_649);
nor U1655 (N_1655,In_4759,N_586);
nor U1656 (N_1656,In_4914,In_952);
and U1657 (N_1657,N_475,In_2243);
and U1658 (N_1658,In_1459,In_4421);
or U1659 (N_1659,N_965,In_2110);
xnor U1660 (N_1660,In_4107,In_4346);
nor U1661 (N_1661,In_172,In_2798);
and U1662 (N_1662,In_1251,In_1386);
xnor U1663 (N_1663,In_891,In_848);
xnor U1664 (N_1664,N_866,In_1393);
or U1665 (N_1665,In_1112,In_1894);
xnor U1666 (N_1666,N_966,N_604);
and U1667 (N_1667,In_782,In_1451);
or U1668 (N_1668,N_181,In_2959);
xor U1669 (N_1669,In_1136,N_339);
nor U1670 (N_1670,In_1904,In_3138);
or U1671 (N_1671,N_916,In_1130);
and U1672 (N_1672,In_4168,In_4820);
nor U1673 (N_1673,N_841,N_796);
xor U1674 (N_1674,In_3911,In_2251);
nand U1675 (N_1675,In_4406,In_3597);
nor U1676 (N_1676,In_3679,In_89);
or U1677 (N_1677,In_2371,N_851);
or U1678 (N_1678,In_3615,In_1754);
nor U1679 (N_1679,In_1912,In_4574);
nand U1680 (N_1680,In_3443,In_3586);
nand U1681 (N_1681,In_2850,In_4360);
xor U1682 (N_1682,In_1068,In_3416);
xnor U1683 (N_1683,N_413,In_4532);
nand U1684 (N_1684,In_3183,N_588);
nor U1685 (N_1685,In_669,In_1808);
nand U1686 (N_1686,In_4738,In_2689);
nor U1687 (N_1687,In_4413,In_1986);
and U1688 (N_1688,N_411,In_1244);
xor U1689 (N_1689,In_329,In_1193);
xnor U1690 (N_1690,In_1662,N_232);
or U1691 (N_1691,In_4561,In_1365);
nand U1692 (N_1692,In_306,In_1134);
or U1693 (N_1693,N_915,In_4625);
nor U1694 (N_1694,In_1104,N_21);
nand U1695 (N_1695,In_1198,In_689);
xor U1696 (N_1696,In_1388,In_4411);
nor U1697 (N_1697,In_3863,In_728);
nand U1698 (N_1698,In_1180,In_867);
nand U1699 (N_1699,In_3152,In_1967);
xor U1700 (N_1700,In_1032,In_2398);
nor U1701 (N_1701,In_1199,In_539);
nor U1702 (N_1702,In_664,N_627);
or U1703 (N_1703,In_4120,In_4663);
or U1704 (N_1704,In_4192,In_2708);
and U1705 (N_1705,In_4028,In_3536);
nor U1706 (N_1706,In_1497,In_3661);
nor U1707 (N_1707,In_1955,In_1726);
and U1708 (N_1708,N_516,In_2443);
xor U1709 (N_1709,In_3779,N_364);
nor U1710 (N_1710,N_190,In_1243);
nor U1711 (N_1711,In_3961,N_133);
nand U1712 (N_1712,In_3864,In_903);
and U1713 (N_1713,N_143,In_3339);
or U1714 (N_1714,In_4757,In_4668);
nand U1715 (N_1715,In_4956,N_305);
nor U1716 (N_1716,In_4569,In_1695);
nor U1717 (N_1717,N_291,In_2117);
xor U1718 (N_1718,In_495,In_3949);
xor U1719 (N_1719,In_2591,N_721);
nand U1720 (N_1720,In_4605,In_4961);
nand U1721 (N_1721,In_1541,In_2932);
or U1722 (N_1722,In_1789,N_40);
nor U1723 (N_1723,N_971,In_3389);
nor U1724 (N_1724,In_3125,In_1064);
or U1725 (N_1725,In_429,In_2122);
and U1726 (N_1726,N_67,In_2608);
nor U1727 (N_1727,In_3705,In_4363);
nand U1728 (N_1728,In_3505,In_4498);
nor U1729 (N_1729,In_3208,In_2016);
xnor U1730 (N_1730,In_4111,In_2138);
nand U1731 (N_1731,In_3887,In_399);
or U1732 (N_1732,In_4435,In_4228);
or U1733 (N_1733,In_1611,In_436);
nand U1734 (N_1734,N_483,In_3858);
and U1735 (N_1735,N_518,In_3671);
nand U1736 (N_1736,In_1995,In_1529);
or U1737 (N_1737,N_736,In_4197);
and U1738 (N_1738,In_2525,In_1174);
and U1739 (N_1739,In_4813,In_194);
xor U1740 (N_1740,In_3725,In_1432);
and U1741 (N_1741,In_1317,In_3667);
or U1742 (N_1742,In_1599,In_1618);
nor U1743 (N_1743,In_2039,In_3616);
nand U1744 (N_1744,In_4126,In_2051);
nor U1745 (N_1745,N_228,In_3028);
or U1746 (N_1746,In_1145,In_4404);
and U1747 (N_1747,In_980,N_27);
xnor U1748 (N_1748,In_4365,In_729);
or U1749 (N_1749,In_4966,N_399);
xnor U1750 (N_1750,In_531,N_333);
or U1751 (N_1751,In_927,N_659);
nor U1752 (N_1752,N_827,N_464);
nand U1753 (N_1753,In_2258,In_4873);
or U1754 (N_1754,In_3142,N_645);
or U1755 (N_1755,In_1494,N_790);
and U1756 (N_1756,In_1080,In_2450);
or U1757 (N_1757,N_696,N_941);
nand U1758 (N_1758,In_2630,N_905);
xnor U1759 (N_1759,N_803,In_1405);
and U1760 (N_1760,In_2710,In_2809);
and U1761 (N_1761,N_149,In_2431);
or U1762 (N_1762,In_4693,In_4258);
and U1763 (N_1763,N_373,N_581);
xnor U1764 (N_1764,In_1791,In_4980);
and U1765 (N_1765,In_3407,In_1156);
or U1766 (N_1766,N_176,In_3573);
nor U1767 (N_1767,In_2937,In_1341);
and U1768 (N_1768,N_521,In_2445);
and U1769 (N_1769,In_4042,In_2891);
and U1770 (N_1770,In_2967,In_2168);
or U1771 (N_1771,In_1643,In_1461);
nand U1772 (N_1772,In_3149,N_440);
nor U1773 (N_1773,In_4861,In_3313);
or U1774 (N_1774,In_4620,N_911);
and U1775 (N_1775,In_3363,In_3039);
or U1776 (N_1776,In_3809,In_4486);
or U1777 (N_1777,In_4473,In_4358);
nor U1778 (N_1778,In_3033,In_2540);
nand U1779 (N_1779,In_3446,N_178);
nand U1780 (N_1780,In_1659,N_218);
nor U1781 (N_1781,In_176,N_35);
nor U1782 (N_1782,In_1407,N_141);
nor U1783 (N_1783,In_2581,N_665);
nand U1784 (N_1784,N_400,In_3556);
xor U1785 (N_1785,N_297,In_2594);
nor U1786 (N_1786,In_3209,N_107);
xor U1787 (N_1787,In_424,In_2324);
and U1788 (N_1788,In_4179,In_2661);
xnor U1789 (N_1789,In_1262,In_3521);
xnor U1790 (N_1790,N_197,In_2336);
xnor U1791 (N_1791,In_956,In_4549);
and U1792 (N_1792,In_607,N_579);
xor U1793 (N_1793,In_3059,In_3915);
nand U1794 (N_1794,In_476,In_1777);
nor U1795 (N_1795,N_563,In_910);
xor U1796 (N_1796,In_4713,In_2451);
nand U1797 (N_1797,In_467,N_658);
xor U1798 (N_1798,In_8,N_597);
and U1799 (N_1799,In_697,In_3832);
or U1800 (N_1800,N_391,In_2739);
or U1801 (N_1801,In_685,In_4647);
or U1802 (N_1802,In_3099,N_684);
and U1803 (N_1803,In_1652,N_873);
xnor U1804 (N_1804,In_1783,In_1467);
and U1805 (N_1805,In_4298,In_1100);
xnor U1806 (N_1806,In_3584,In_4616);
or U1807 (N_1807,In_1625,In_1731);
or U1808 (N_1808,In_42,In_4701);
nand U1809 (N_1809,In_2940,N_303);
xnor U1810 (N_1810,N_371,In_4879);
nor U1811 (N_1811,In_1853,In_2453);
nor U1812 (N_1812,N_859,In_2770);
nor U1813 (N_1813,In_4829,In_3945);
nor U1814 (N_1814,In_1636,In_3910);
or U1815 (N_1815,In_72,In_654);
or U1816 (N_1816,In_2516,In_1884);
or U1817 (N_1817,In_846,In_438);
nand U1818 (N_1818,In_911,In_160);
or U1819 (N_1819,In_2153,In_1481);
nor U1820 (N_1820,In_2615,In_494);
or U1821 (N_1821,In_4156,In_4022);
nor U1822 (N_1822,In_4513,N_150);
nand U1823 (N_1823,In_2082,In_3088);
nor U1824 (N_1824,N_423,In_1640);
nor U1825 (N_1825,In_2836,In_1303);
xnor U1826 (N_1826,N_280,In_1217);
and U1827 (N_1827,In_2432,In_3247);
xor U1828 (N_1828,In_1194,In_828);
nor U1829 (N_1829,In_135,N_522);
and U1830 (N_1830,In_4762,In_1586);
or U1831 (N_1831,N_2,In_1196);
or U1832 (N_1832,In_1609,In_1326);
and U1833 (N_1833,In_4367,In_2800);
nor U1834 (N_1834,N_12,In_3076);
and U1835 (N_1835,In_3857,N_566);
xor U1836 (N_1836,In_4147,In_3985);
nand U1837 (N_1837,In_59,In_2358);
or U1838 (N_1838,In_1311,In_212);
nand U1839 (N_1839,In_3783,In_7);
or U1840 (N_1840,In_3295,In_1288);
xor U1841 (N_1841,In_2987,In_3087);
and U1842 (N_1842,In_4249,In_154);
or U1843 (N_1843,In_2509,N_737);
xnor U1844 (N_1844,N_401,N_334);
and U1845 (N_1845,In_832,N_767);
nor U1846 (N_1846,In_3012,In_4169);
nor U1847 (N_1847,N_812,In_315);
nand U1848 (N_1848,In_727,In_1998);
nor U1849 (N_1849,N_70,In_1218);
xnor U1850 (N_1850,In_2077,In_1917);
or U1851 (N_1851,In_4098,In_294);
nand U1852 (N_1852,In_3474,In_2344);
xor U1853 (N_1853,In_1116,N_368);
nor U1854 (N_1854,In_3918,In_1282);
nor U1855 (N_1855,N_75,N_233);
nor U1856 (N_1856,N_950,In_4342);
or U1857 (N_1857,In_4741,In_3816);
and U1858 (N_1858,In_3411,In_4140);
nand U1859 (N_1859,N_826,In_1713);
xnor U1860 (N_1860,In_3700,N_435);
nand U1861 (N_1861,In_4066,N_560);
xor U1862 (N_1862,In_3246,In_3607);
or U1863 (N_1863,In_4945,N_414);
and U1864 (N_1864,In_4242,In_2508);
xnor U1865 (N_1865,N_592,In_1748);
xor U1866 (N_1866,In_3320,In_2119);
and U1867 (N_1867,In_3926,In_417);
xor U1868 (N_1868,In_2869,N_224);
or U1869 (N_1869,In_1182,In_4211);
nand U1870 (N_1870,In_4277,N_724);
xnor U1871 (N_1871,In_1923,In_4703);
xnor U1872 (N_1872,N_835,In_4307);
nor U1873 (N_1873,In_505,In_2720);
and U1874 (N_1874,In_4326,N_593);
or U1875 (N_1875,In_2061,In_2221);
xor U1876 (N_1876,N_632,In_3197);
and U1877 (N_1877,In_3447,N_517);
or U1878 (N_1878,In_115,In_4553);
or U1879 (N_1879,In_3970,In_1734);
or U1880 (N_1880,In_4603,In_3631);
nand U1881 (N_1881,In_4610,In_480);
xnor U1882 (N_1882,In_3438,In_4389);
nand U1883 (N_1883,N_445,In_4856);
and U1884 (N_1884,In_1036,N_352);
xnor U1885 (N_1885,In_123,In_3889);
nor U1886 (N_1886,N_362,In_3847);
or U1887 (N_1887,In_2469,In_3922);
nand U1888 (N_1888,In_1972,N_574);
nand U1889 (N_1889,N_206,N_450);
and U1890 (N_1890,N_757,In_1150);
nand U1891 (N_1891,N_509,In_4789);
xnor U1892 (N_1892,In_632,In_3674);
nor U1893 (N_1893,In_2143,N_917);
and U1894 (N_1894,In_1569,In_1524);
nor U1895 (N_1895,In_488,In_871);
nor U1896 (N_1896,N_465,In_4076);
and U1897 (N_1897,In_2161,N_406);
or U1898 (N_1898,In_2561,N_145);
or U1899 (N_1899,N_577,N_120);
and U1900 (N_1900,In_985,In_1525);
xor U1901 (N_1901,In_2353,In_2095);
nor U1902 (N_1902,In_4150,N_914);
nand U1903 (N_1903,N_629,In_3676);
nand U1904 (N_1904,N_614,In_2729);
xnor U1905 (N_1905,In_1676,In_3269);
nand U1906 (N_1906,In_4350,In_3020);
xor U1907 (N_1907,N_202,N_582);
nor U1908 (N_1908,In_3158,In_346);
xor U1909 (N_1909,In_1527,N_786);
and U1910 (N_1910,In_3196,In_2942);
xor U1911 (N_1911,N_160,In_1598);
xnor U1912 (N_1912,In_3188,In_2750);
nand U1913 (N_1913,In_4763,In_1733);
or U1914 (N_1914,In_440,In_1745);
and U1915 (N_1915,In_163,In_188);
nand U1916 (N_1916,In_1202,In_3318);
xor U1917 (N_1917,In_3383,N_828);
nor U1918 (N_1918,In_3912,In_3380);
xnor U1919 (N_1919,In_1499,In_813);
nand U1920 (N_1920,In_2902,N_893);
nor U1921 (N_1921,N_427,In_3534);
and U1922 (N_1922,N_9,In_2278);
xor U1923 (N_1923,In_3835,In_1002);
or U1924 (N_1924,In_350,N_316);
or U1925 (N_1925,In_2198,N_459);
or U1926 (N_1926,In_4297,In_2668);
and U1927 (N_1927,In_623,N_45);
or U1928 (N_1928,In_1675,N_653);
and U1929 (N_1929,In_4136,N_57);
and U1930 (N_1930,In_4884,N_345);
nand U1931 (N_1931,In_1613,N_631);
nor U1932 (N_1932,In_249,N_727);
xor U1933 (N_1933,N_666,In_1989);
nor U1934 (N_1934,In_1871,In_4144);
nor U1935 (N_1935,In_2373,In_4390);
or U1936 (N_1936,N_132,N_561);
or U1937 (N_1937,N_18,In_4710);
and U1938 (N_1938,In_1940,In_4897);
nand U1939 (N_1939,In_2603,In_463);
nand U1940 (N_1940,In_3126,In_2270);
and U1941 (N_1941,N_595,In_2124);
nand U1942 (N_1942,In_403,In_3473);
nand U1943 (N_1943,In_3174,In_2748);
nand U1944 (N_1944,N_651,In_3730);
nand U1945 (N_1945,In_3856,N_136);
nand U1946 (N_1946,N_386,In_3929);
or U1947 (N_1947,In_1629,N_106);
or U1948 (N_1948,In_314,N_365);
and U1949 (N_1949,In_3681,N_201);
and U1950 (N_1950,In_271,In_1404);
nor U1951 (N_1951,N_38,In_1504);
nand U1952 (N_1952,N_205,In_1187);
nand U1953 (N_1953,In_2929,In_4881);
xor U1954 (N_1954,In_4908,In_323);
xor U1955 (N_1955,In_517,In_1654);
and U1956 (N_1956,In_3408,In_2498);
or U1957 (N_1957,N_903,N_169);
and U1958 (N_1958,In_2090,In_2178);
xor U1959 (N_1959,N_29,In_3655);
and U1960 (N_1960,In_2722,In_1072);
or U1961 (N_1961,In_1872,In_4027);
nand U1962 (N_1962,In_719,In_4724);
nand U1963 (N_1963,In_54,In_3853);
nor U1964 (N_1964,N_447,In_2900);
or U1965 (N_1965,In_4686,In_1863);
nor U1966 (N_1966,N_946,In_1954);
and U1967 (N_1967,N_124,In_3956);
xnor U1968 (N_1968,In_4792,In_939);
nor U1969 (N_1969,In_4474,In_3718);
and U1970 (N_1970,N_718,In_464);
and U1971 (N_1971,In_3071,In_3873);
nor U1972 (N_1972,In_2964,In_3501);
xor U1973 (N_1973,N_700,In_3978);
nand U1974 (N_1974,In_1118,In_4566);
nor U1975 (N_1975,N_426,N_71);
nand U1976 (N_1976,N_213,In_4383);
or U1977 (N_1977,In_1750,In_2740);
nor U1978 (N_1978,N_390,In_489);
xnor U1979 (N_1979,In_2287,N_576);
nand U1980 (N_1980,In_2074,In_2216);
and U1981 (N_1981,In_4904,In_2535);
nand U1982 (N_1982,In_4711,In_4679);
and U1983 (N_1983,In_498,In_2368);
xor U1984 (N_1984,In_2658,In_2482);
xnor U1985 (N_1985,N_272,In_1717);
nor U1986 (N_1986,In_4441,In_643);
or U1987 (N_1987,In_2170,In_842);
or U1988 (N_1988,N_53,In_4756);
or U1989 (N_1989,In_1135,In_1325);
or U1990 (N_1990,In_4044,In_3074);
xor U1991 (N_1991,In_2409,In_2301);
and U1992 (N_1992,In_2588,In_4937);
or U1993 (N_1993,In_4722,In_1154);
nor U1994 (N_1994,N_958,In_4148);
xnor U1995 (N_1995,N_446,In_4232);
nor U1996 (N_1996,In_1475,In_2475);
xor U1997 (N_1997,In_1915,N_740);
nand U1998 (N_1998,In_1576,In_3690);
or U1999 (N_1999,In_180,In_2593);
nand U2000 (N_2000,N_1650,In_4564);
nor U2001 (N_2001,In_1140,N_644);
xor U2002 (N_2002,N_816,N_1495);
xor U2003 (N_2003,N_768,N_1792);
or U2004 (N_2004,N_7,In_4254);
and U2005 (N_2005,In_1630,In_99);
nor U2006 (N_2006,In_2774,N_1084);
xnor U2007 (N_2007,In_1756,N_1514);
xnor U2008 (N_2008,N_1048,In_631);
or U2009 (N_2009,In_4129,In_4250);
xor U2010 (N_2010,N_742,N_1803);
xnor U2011 (N_2011,N_1441,In_4394);
or U2012 (N_2012,N_1298,N_1590);
and U2013 (N_2013,N_1209,N_356);
nor U2014 (N_2014,N_1367,In_2306);
nor U2015 (N_2015,In_730,In_4246);
nor U2016 (N_2016,In_4302,N_1301);
or U2017 (N_2017,N_1314,N_1079);
and U2018 (N_2018,N_636,In_875);
xor U2019 (N_2019,N_1007,N_191);
and U2020 (N_2020,N_1864,N_1361);
nor U2021 (N_2021,N_784,In_3140);
and U2022 (N_2022,In_260,N_870);
nor U2023 (N_2023,N_1954,In_2302);
nand U2024 (N_2024,N_375,N_1745);
and U2025 (N_2025,N_1169,In_1880);
nand U2026 (N_2026,N_687,In_3510);
xor U2027 (N_2027,In_1550,N_1980);
and U2028 (N_2028,N_1641,N_1587);
and U2029 (N_2029,N_1880,N_723);
and U2030 (N_2030,In_3543,N_1718);
and U2031 (N_2031,N_1093,N_709);
nor U2032 (N_2032,N_1645,In_1207);
nor U2033 (N_2033,In_3703,N_889);
nand U2034 (N_2034,N_1941,In_2397);
xnor U2035 (N_2035,N_1001,In_1473);
nand U2036 (N_2036,N_762,In_4584);
and U2037 (N_2037,In_4854,N_1874);
or U2038 (N_2038,N_1646,N_1833);
nor U2039 (N_2039,In_4237,In_469);
xnor U2040 (N_2040,N_806,N_844);
or U2041 (N_2041,In_1411,N_408);
nand U2042 (N_2042,In_4846,In_1337);
xor U2043 (N_2043,N_511,In_4903);
xnor U2044 (N_2044,In_3306,In_1441);
nand U2045 (N_2045,In_4907,N_226);
xor U2046 (N_2046,In_3589,N_1065);
or U2047 (N_2047,N_1281,N_720);
and U2048 (N_2048,N_102,In_1814);
and U2049 (N_2049,N_1290,N_707);
or U2050 (N_2050,N_681,In_4665);
xor U2051 (N_2051,In_1231,In_4690);
nand U2052 (N_2052,N_441,In_3593);
nand U2053 (N_2053,N_1478,In_940);
nand U2054 (N_2054,In_251,N_748);
or U2055 (N_2055,N_1109,N_1154);
and U2056 (N_2056,In_2317,In_344);
nor U2057 (N_2057,In_783,N_1935);
nand U2058 (N_2058,N_1708,In_1864);
nor U2059 (N_2059,N_797,In_2047);
or U2060 (N_2060,In_2745,N_1038);
nand U2061 (N_2061,In_4535,In_1355);
nand U2062 (N_2062,In_254,N_346);
and U2063 (N_2063,N_1611,N_1243);
xnor U2064 (N_2064,In_2014,In_1045);
xor U2065 (N_2065,N_596,N_1624);
nor U2066 (N_2066,N_552,N_760);
nand U2067 (N_2067,N_1932,In_1286);
nor U2068 (N_2068,In_3545,In_707);
nand U2069 (N_2069,N_1508,In_4186);
or U2070 (N_2070,N_1610,In_3991);
xor U2071 (N_2071,N_745,N_1620);
or U2072 (N_2072,N_1526,In_2810);
xnor U2073 (N_2073,In_4984,In_3996);
xor U2074 (N_2074,N_1158,In_2455);
nor U2075 (N_2075,In_1429,N_1688);
or U2076 (N_2076,In_82,N_289);
nor U2077 (N_2077,N_97,In_2485);
nand U2078 (N_2078,In_4962,In_2997);
nor U2079 (N_2079,In_3121,N_1615);
xnor U2080 (N_2080,In_169,In_1906);
nor U2081 (N_2081,In_2771,In_1549);
nand U2082 (N_2082,N_1710,In_408);
and U2083 (N_2083,N_1921,N_895);
xor U2084 (N_2084,N_628,N_1573);
or U2085 (N_2085,N_1012,In_2612);
and U2086 (N_2086,In_1673,In_4279);
nor U2087 (N_2087,N_565,In_4602);
nand U2088 (N_2088,N_295,In_2646);
xor U2089 (N_2089,In_4811,In_4556);
nand U2090 (N_2090,In_3959,In_3742);
and U2091 (N_2091,In_2901,In_1304);
nor U2092 (N_2092,In_4052,N_822);
xnor U2093 (N_2093,N_1550,N_1340);
and U2094 (N_2094,In_2395,In_2698);
nor U2095 (N_2095,N_1265,N_947);
xor U2096 (N_2096,In_722,In_4019);
and U2097 (N_2097,In_4121,N_1876);
xnor U2098 (N_2098,In_988,In_578);
xor U2099 (N_2099,In_3366,In_4888);
or U2100 (N_2100,In_4235,In_1458);
and U2101 (N_2101,N_1999,N_1578);
nand U2102 (N_2102,N_882,In_2463);
and U2103 (N_2103,In_2112,In_653);
or U2104 (N_2104,N_1172,In_1014);
or U2105 (N_2105,In_1433,In_4485);
and U2106 (N_2106,In_4918,N_179);
nor U2107 (N_2107,In_3803,N_1104);
nand U2108 (N_2108,N_1509,In_3167);
and U2109 (N_2109,In_3896,In_2030);
xor U2110 (N_2110,N_1625,N_1156);
nand U2111 (N_2111,In_1206,N_200);
or U2112 (N_2112,N_1837,In_4670);
nand U2113 (N_2113,In_659,In_1440);
nand U2114 (N_2114,N_1966,In_1934);
and U2115 (N_2115,N_25,N_1997);
nand U2116 (N_2116,N_1783,In_1236);
nor U2117 (N_2117,N_1496,N_1548);
and U2118 (N_2118,N_1284,N_1060);
or U2119 (N_2119,In_1161,In_2300);
or U2120 (N_2120,In_757,N_704);
or U2121 (N_2121,In_1969,N_1062);
xnor U2122 (N_2122,In_4915,N_1433);
xnor U2123 (N_2123,N_397,In_4534);
and U2124 (N_2124,N_389,N_50);
xnor U2125 (N_2125,N_1221,N_1175);
nand U2126 (N_2126,In_1491,N_781);
nand U2127 (N_2127,N_1150,In_4077);
or U2128 (N_2128,N_442,N_1998);
or U2129 (N_2129,N_545,In_4178);
xor U2130 (N_2130,N_1438,N_1970);
xnor U2131 (N_2131,N_1727,N_862);
nor U2132 (N_2132,N_1262,N_1075);
xnor U2133 (N_2133,N_1181,N_551);
xnor U2134 (N_2134,N_1824,In_3165);
xor U2135 (N_2135,In_3038,In_4423);
nor U2136 (N_2136,In_2159,In_2019);
xor U2137 (N_2137,In_1932,In_3849);
or U2138 (N_2138,In_2826,In_2338);
xnor U2139 (N_2139,N_100,In_3204);
nand U2140 (N_2140,In_906,N_1195);
or U2141 (N_2141,N_1740,In_799);
or U2142 (N_2142,In_1827,In_338);
nand U2143 (N_2143,In_4282,In_2420);
nand U2144 (N_2144,In_4247,N_885);
or U2145 (N_2145,N_699,N_750);
and U2146 (N_2146,In_4476,In_4747);
nor U2147 (N_2147,In_1620,N_1108);
xor U2148 (N_2148,In_1228,N_91);
nand U2149 (N_2149,In_2331,N_484);
and U2150 (N_2150,N_1771,N_1160);
or U2151 (N_2151,N_890,N_1260);
nor U2152 (N_2152,In_1371,In_4985);
nand U2153 (N_2153,N_1422,N_1388);
xnor U2154 (N_2154,In_4448,N_341);
and U2155 (N_2155,N_1678,N_1991);
xnor U2156 (N_2156,N_744,In_2764);
xor U2157 (N_2157,In_2518,In_1157);
or U2158 (N_2158,N_1378,In_2948);
or U2159 (N_2159,In_3340,In_2614);
nand U2160 (N_2160,In_3693,In_3628);
xor U2161 (N_2161,In_1990,N_1020);
nor U2162 (N_2162,In_1409,In_3419);
nand U2163 (N_2163,N_1859,In_2290);
xnor U2164 (N_2164,In_1881,N_689);
xnor U2165 (N_2165,In_1657,N_1557);
and U2166 (N_2166,In_1442,In_4306);
or U2167 (N_2167,In_3355,In_1854);
nor U2168 (N_2168,N_1787,N_1434);
xnor U2169 (N_2169,N_1237,In_4545);
xor U2170 (N_2170,N_1556,N_1330);
xor U2171 (N_2171,N_1067,In_430);
nor U2172 (N_2172,N_1019,N_1774);
and U2173 (N_2173,In_3461,N_1600);
or U2174 (N_2174,In_3055,In_3897);
nand U2175 (N_2175,In_375,N_761);
xor U2176 (N_2176,N_1746,N_888);
or U2177 (N_2177,N_1705,N_1605);
and U2178 (N_2178,In_3337,N_874);
or U2179 (N_2179,N_1567,N_710);
nand U2180 (N_2180,N_1977,N_846);
xnor U2181 (N_2181,N_117,N_1044);
xnor U2182 (N_2182,In_3072,In_4412);
nand U2183 (N_2183,N_1056,In_1123);
nand U2184 (N_2184,In_1552,N_1955);
xor U2185 (N_2185,N_1407,N_113);
nand U2186 (N_2186,N_1292,In_3865);
xnor U2187 (N_2187,In_4426,In_904);
or U2188 (N_2188,N_1432,In_4154);
xnor U2189 (N_2189,N_1719,N_1720);
nand U2190 (N_2190,N_1054,In_179);
and U2191 (N_2191,N_1647,N_1482);
nor U2192 (N_2192,N_1368,N_1994);
xnor U2193 (N_2193,In_2197,In_3228);
and U2194 (N_2194,N_601,In_4012);
or U2195 (N_2195,In_1165,N_452);
and U2196 (N_2196,In_3171,N_547);
nand U2197 (N_2197,N_570,In_3172);
and U2198 (N_2198,In_320,In_1013);
or U2199 (N_2199,In_280,N_1384);
or U2200 (N_2200,N_1357,In_2322);
and U2201 (N_2201,N_680,N_879);
and U2202 (N_2202,N_15,In_2635);
nor U2203 (N_2203,In_3684,N_1008);
nor U2204 (N_2204,N_1529,In_825);
nor U2205 (N_2205,N_1356,N_1014);
and U2206 (N_2206,In_4381,In_1189);
or U2207 (N_2207,In_219,N_1703);
nand U2208 (N_2208,N_1387,N_1992);
and U2209 (N_2209,N_1850,N_164);
or U2210 (N_2210,In_1746,N_1589);
xor U2211 (N_2211,N_1462,N_1198);
or U2212 (N_2212,N_1964,In_3047);
or U2213 (N_2213,N_498,In_1366);
and U2214 (N_2214,N_1489,N_1831);
xor U2215 (N_2215,N_1847,N_243);
nand U2216 (N_2216,N_1902,In_4538);
nand U2217 (N_2217,N_1155,N_936);
nand U2218 (N_2218,In_2576,In_4468);
or U2219 (N_2219,N_1133,N_306);
nor U2220 (N_2220,N_1974,N_129);
nand U2221 (N_2221,N_290,In_930);
xor U2222 (N_2222,N_1493,N_1956);
or U2223 (N_2223,N_602,N_677);
nand U2224 (N_2224,N_1763,In_3384);
and U2225 (N_2225,In_456,In_2711);
nand U2226 (N_2226,N_1080,N_1677);
nor U2227 (N_2227,In_4685,N_1118);
or U2228 (N_2228,In_2989,N_1338);
and U2229 (N_2229,N_321,In_418);
and U2230 (N_2230,N_1127,N_344);
nor U2231 (N_2231,N_1598,N_96);
nor U2232 (N_2232,In_3714,N_1767);
or U2233 (N_2233,In_1669,In_1259);
xor U2234 (N_2234,N_163,In_2753);
nor U2235 (N_2235,N_236,N_1279);
and U2236 (N_2236,In_3746,In_62);
nand U2237 (N_2237,In_1179,In_4622);
nand U2238 (N_2238,N_1873,N_1969);
xor U2239 (N_2239,In_3660,In_3537);
and U2240 (N_2240,In_2183,N_1738);
xnor U2241 (N_2241,In_3255,N_1409);
nor U2242 (N_2242,In_2889,N_1025);
nand U2243 (N_2243,In_2547,N_1633);
and U2244 (N_2244,N_302,In_4058);
or U2245 (N_2245,In_2911,N_1802);
and U2246 (N_2246,N_1981,In_3050);
nor U2247 (N_2247,In_1005,N_208);
xnor U2248 (N_2248,In_686,In_1948);
nor U2249 (N_2249,N_1782,N_1501);
or U2250 (N_2250,N_1448,In_773);
nand U2251 (N_2251,N_1344,In_2389);
nand U2252 (N_2252,In_4933,N_1764);
or U2253 (N_2253,In_1017,In_1891);
nand U2254 (N_2254,In_2634,N_1293);
xnor U2255 (N_2255,N_530,N_493);
and U2256 (N_2256,N_300,N_1091);
xnor U2257 (N_2257,In_655,In_1313);
nand U2258 (N_2258,In_931,N_1112);
or U2259 (N_2259,In_2410,N_1616);
or U2260 (N_2260,N_256,In_4851);
and U2261 (N_2261,In_3230,In_3837);
and U2262 (N_2262,N_990,In_2813);
or U2263 (N_2263,N_1623,N_667);
and U2264 (N_2264,In_2244,N_1622);
and U2265 (N_2265,In_3824,In_1377);
xnor U2266 (N_2266,In_970,In_4608);
xor U2267 (N_2267,In_2802,N_1389);
xnor U2268 (N_2268,N_1614,In_12);
or U2269 (N_2269,In_3007,In_2880);
or U2270 (N_2270,N_1412,In_752);
nor U2271 (N_2271,N_1463,In_741);
nor U2272 (N_2272,In_1106,In_1886);
xor U2273 (N_2273,In_4501,In_3726);
or U2274 (N_2274,In_4265,N_1652);
xnor U2275 (N_2275,N_1822,In_1152);
and U2276 (N_2276,N_857,N_1535);
nand U2277 (N_2277,N_1100,N_55);
nand U2278 (N_2278,In_1686,In_3507);
nand U2279 (N_2279,In_1030,In_3618);
and U2280 (N_2280,N_1337,N_510);
xnor U2281 (N_2281,In_4490,N_514);
and U2282 (N_2282,In_3903,In_4427);
or U2283 (N_2283,N_221,N_557);
and U2284 (N_2284,N_1437,In_483);
nor U2285 (N_2285,N_1674,In_4328);
xnor U2286 (N_2286,N_1197,N_274);
nor U2287 (N_2287,N_1993,N_743);
xnor U2288 (N_2288,In_3569,In_3692);
or U2289 (N_2289,N_842,N_1263);
xnor U2290 (N_2290,N_1006,N_1444);
and U2291 (N_2291,In_3500,In_859);
xnor U2292 (N_2292,N_697,N_1440);
nand U2293 (N_2293,N_788,In_989);
xor U2294 (N_2294,N_648,In_3358);
xor U2295 (N_2295,In_1821,In_857);
xnor U2296 (N_2296,N_1310,In_2607);
nand U2297 (N_2297,In_4830,In_1768);
xor U2298 (N_2298,In_3673,In_3759);
and U2299 (N_2299,N_734,In_584);
nand U2300 (N_2300,N_1982,In_1820);
nor U2301 (N_2301,N_1903,In_1412);
xnor U2302 (N_2302,In_608,N_1704);
nor U2303 (N_2303,N_1896,In_525);
or U2304 (N_2304,N_449,N_1654);
and U2305 (N_2305,N_584,N_1226);
nand U2306 (N_2306,In_3405,N_1189);
nor U2307 (N_2307,N_1827,N_219);
nand U2308 (N_2308,In_3880,In_4699);
nand U2309 (N_2309,N_1663,In_1573);
nor U2310 (N_2310,N_1403,In_1358);
nand U2311 (N_2311,In_371,In_77);
nand U2312 (N_2312,N_328,In_3974);
xor U2313 (N_2313,N_1806,N_1584);
or U2314 (N_2314,In_4576,N_203);
and U2315 (N_2315,N_209,In_102);
or U2316 (N_2316,N_1073,N_856);
nand U2317 (N_2317,In_1994,N_380);
or U2318 (N_2318,In_626,In_3763);
xnor U2319 (N_2319,In_200,N_1671);
xnor U2320 (N_2320,N_1256,N_1990);
xnor U2321 (N_2321,In_3113,N_329);
nand U2322 (N_2322,In_1378,N_1939);
nor U2323 (N_2323,N_1202,In_2350);
and U2324 (N_2324,N_1607,N_1471);
nor U2325 (N_2325,N_381,In_2747);
xor U2326 (N_2326,In_2851,In_2865);
and U2327 (N_2327,N_1592,N_111);
nor U2328 (N_2328,N_934,In_3274);
nand U2329 (N_2329,N_1809,In_577);
and U2330 (N_2330,N_1031,N_1494);
nand U2331 (N_2331,N_1919,N_1617);
or U2332 (N_2332,N_1479,In_4386);
xor U2333 (N_2333,N_1748,In_3650);
xor U2334 (N_2334,In_2262,N_1454);
or U2335 (N_2335,In_1792,N_451);
or U2336 (N_2336,N_1794,N_1413);
nor U2337 (N_2337,In_1852,N_1327);
xnor U2338 (N_2338,In_4568,In_1692);
or U2339 (N_2339,N_787,N_1664);
or U2340 (N_2340,In_1077,In_3066);
xnor U2341 (N_2341,N_51,In_1794);
and U2342 (N_2342,In_2895,In_2156);
nor U2343 (N_2343,N_1618,In_3623);
nand U2344 (N_2344,N_1341,N_8);
xor U2345 (N_2345,N_1205,N_1032);
nor U2346 (N_2346,N_1336,N_86);
or U2347 (N_2347,In_3633,N_294);
xnor U2348 (N_2348,N_92,In_1356);
or U2349 (N_2349,In_262,N_1658);
or U2350 (N_2350,In_810,N_1242);
nor U2351 (N_2351,N_1015,N_1376);
or U2352 (N_2352,In_3454,N_1326);
xnor U2353 (N_2353,In_1453,In_1364);
xnor U2354 (N_2354,In_993,N_1206);
xor U2355 (N_2355,In_485,N_1096);
or U2356 (N_2356,N_424,In_3252);
and U2357 (N_2357,N_1971,N_1712);
nor U2358 (N_2358,In_4849,In_3622);
nor U2359 (N_2359,N_782,In_3829);
xor U2360 (N_2360,In_736,N_969);
or U2361 (N_2361,N_1165,N_955);
nor U2362 (N_2362,In_4001,N_1443);
xor U2363 (N_2363,N_1307,In_4867);
or U2364 (N_2364,N_479,N_1207);
or U2365 (N_2365,N_252,In_1590);
nand U2366 (N_2366,N_683,N_1322);
and U2367 (N_2367,In_3261,In_1395);
or U2368 (N_2368,N_1694,In_789);
and U2369 (N_2369,N_1061,In_3117);
xnor U2370 (N_2370,N_1758,N_1204);
nand U2371 (N_2371,N_1497,In_4835);
and U2372 (N_2372,N_285,N_1476);
or U2373 (N_2373,N_1306,N_1393);
nand U2374 (N_2374,N_741,N_1419);
xnor U2375 (N_2375,In_678,In_2537);
or U2376 (N_2376,In_4159,In_3966);
nand U2377 (N_2377,N_892,In_1292);
nand U2378 (N_2378,In_572,In_3930);
nor U2379 (N_2379,In_4502,In_4351);
nand U2380 (N_2380,N_1410,N_1846);
nand U2381 (N_2381,In_4528,N_481);
xnor U2382 (N_2382,In_2555,In_4172);
or U2383 (N_2383,In_3139,N_1153);
and U2384 (N_2384,In_991,In_2040);
nand U2385 (N_2385,N_526,N_463);
nor U2386 (N_2386,N_342,In_4798);
xnor U2387 (N_2387,In_1163,In_3924);
nand U2388 (N_2388,N_1588,N_524);
and U2389 (N_2389,In_888,N_1736);
nor U2390 (N_2390,N_1916,In_1483);
and U2391 (N_2391,N_1914,N_1821);
xnor U2392 (N_2392,N_945,In_3933);
or U2393 (N_2393,N_1812,In_91);
nor U2394 (N_2394,N_1095,N_1468);
nand U2395 (N_2395,In_2796,N_708);
and U2396 (N_2396,In_941,N_138);
and U2397 (N_2397,N_860,In_1004);
or U2398 (N_2398,In_1008,N_151);
xor U2399 (N_2399,In_2599,N_1416);
and U2400 (N_2400,N_1791,N_539);
and U2401 (N_2401,N_1670,In_405);
xor U2402 (N_2402,N_1166,N_664);
or U2403 (N_2403,N_1996,N_819);
and U2404 (N_2404,N_377,In_1043);
nand U2405 (N_2405,In_2916,N_661);
nand U2406 (N_2406,In_1374,N_1319);
nor U2407 (N_2407,In_1914,N_1236);
nor U2408 (N_2408,N_1275,In_334);
and U2409 (N_2409,N_546,N_923);
or U2410 (N_2410,N_1034,In_2089);
nor U2411 (N_2411,In_4878,In_3493);
nor U2412 (N_2412,N_1707,N_646);
nor U2413 (N_2413,In_4321,N_1211);
or U2414 (N_2414,In_1111,In_597);
nand U2415 (N_2415,In_1120,In_3232);
nand U2416 (N_2416,N_1343,N_991);
nor U2417 (N_2417,In_4347,In_447);
or U2418 (N_2418,N_799,N_186);
xnor U2419 (N_2419,In_3548,N_378);
nor U2420 (N_2420,In_4403,N_712);
or U2421 (N_2421,In_4967,In_2140);
nor U2422 (N_2422,N_417,N_1485);
or U2423 (N_2423,N_1101,In_4606);
or U2424 (N_2424,In_646,N_98);
nand U2425 (N_2425,In_1678,N_1750);
xnor U2426 (N_2426,N_134,In_1992);
nand U2427 (N_2427,N_1948,N_260);
nor U2428 (N_2428,In_3565,N_967);
or U2429 (N_2429,N_1571,N_85);
xnor U2430 (N_2430,N_1117,N_544);
and U2431 (N_2431,N_1944,In_3118);
or U2432 (N_2432,In_4671,N_1656);
nand U2433 (N_2433,N_1861,N_1568);
and U2434 (N_2434,In_3765,N_432);
nor U2435 (N_2435,In_3833,N_695);
xnor U2436 (N_2436,In_1752,In_34);
nand U2437 (N_2437,In_1623,In_4181);
nand U2438 (N_2438,In_4429,In_2108);
and U2439 (N_2439,In_3004,In_622);
nand U2440 (N_2440,In_2683,N_1212);
xor U2441 (N_2441,In_547,N_1347);
or U2442 (N_2442,N_1978,In_1083);
nand U2443 (N_2443,In_4122,N_1461);
xnor U2444 (N_2444,N_1342,In_4025);
or U2445 (N_2445,N_1234,N_1161);
nand U2446 (N_2446,In_2977,In_1052);
xor U2447 (N_2447,In_1256,In_57);
and U2448 (N_2448,N_1778,N_13);
nand U2449 (N_2449,In_132,In_1200);
nor U2450 (N_2450,N_1762,N_1232);
and U2451 (N_2451,In_4983,In_2248);
and U2452 (N_2452,N_1621,N_1414);
and U2453 (N_2453,N_457,N_1882);
xnor U2454 (N_2454,N_774,In_2018);
nor U2455 (N_2455,N_1458,N_324);
nor U2456 (N_2456,N_1055,In_2806);
nor U2457 (N_2457,In_4187,In_2705);
xor U2458 (N_2458,In_3635,In_326);
nor U2459 (N_2459,N_1820,In_4669);
and U2460 (N_2460,In_3891,In_493);
and U2461 (N_2461,In_3092,In_1551);
xnor U2462 (N_2462,N_1613,In_3567);
nand U2463 (N_2463,In_4555,In_4479);
nand U2464 (N_2464,In_615,In_2133);
xnor U2465 (N_2465,N_1910,In_519);
nand U2466 (N_2466,N_1875,N_1860);
xnor U2467 (N_2467,In_2604,In_2182);
or U2468 (N_2468,N_1987,N_199);
nand U2469 (N_2469,In_4290,In_1760);
nor U2470 (N_2470,N_1315,N_32);
nand U2471 (N_2471,In_1858,N_1952);
xnor U2472 (N_2472,In_2379,In_3751);
nand U2473 (N_2473,In_4761,In_3492);
and U2474 (N_2474,N_1819,N_1223);
xor U2475 (N_2475,In_3542,In_1153);
or U2476 (N_2476,In_2081,In_3672);
xnor U2477 (N_2477,N_1772,In_743);
and U2478 (N_2478,In_3986,N_1349);
or U2479 (N_2479,N_1911,In_2253);
xor U2480 (N_2480,N_1515,N_403);
nand U2481 (N_2481,N_672,In_784);
nand U2482 (N_2482,N_1267,In_1290);
xor U2483 (N_2483,In_734,N_1628);
nand U2484 (N_2484,In_1314,N_615);
nor U2485 (N_2485,N_262,In_1214);
and U2486 (N_2486,N_1883,In_969);
xnor U2487 (N_2487,In_1401,In_535);
xor U2488 (N_2488,In_1665,N_1739);
and U2489 (N_2489,In_2028,In_4449);
xor U2490 (N_2490,N_1768,N_78);
and U2491 (N_2491,In_4283,In_3524);
nor U2492 (N_2492,N_900,N_1466);
or U2493 (N_2493,In_4974,N_500);
and U2494 (N_2494,N_477,In_147);
and U2495 (N_2495,N_1988,In_3333);
or U2496 (N_2496,In_594,In_1312);
and U2497 (N_2497,In_4885,N_1273);
xnor U2498 (N_2498,N_867,In_1622);
or U2499 (N_2499,In_3314,In_2105);
xnor U2500 (N_2500,N_1445,In_533);
nor U2501 (N_2501,N_1576,N_1683);
nand U2502 (N_2502,N_269,In_3544);
and U2503 (N_2503,N_1709,In_3662);
nand U2504 (N_2504,In_3664,N_1085);
and U2505 (N_2505,N_193,N_1644);
nand U2506 (N_2506,In_1191,In_3776);
nand U2507 (N_2507,N_1157,N_813);
or U2508 (N_2508,In_2364,In_2060);
nor U2509 (N_2509,N_1553,N_1922);
nand U2510 (N_2510,N_973,N_312);
nand U2511 (N_2511,N_652,In_3144);
or U2512 (N_2512,N_1131,N_1435);
and U2513 (N_2513,N_939,N_1457);
nor U2514 (N_2514,In_3689,In_4609);
nor U2515 (N_2515,In_1350,N_731);
nand U2516 (N_2516,N_283,In_3721);
nand U2517 (N_2517,N_1271,N_754);
and U2518 (N_2518,In_850,N_1519);
xor U2519 (N_2519,In_750,In_882);
nor U2520 (N_2520,In_4729,N_1408);
xnor U2521 (N_2521,N_1522,N_69);
xor U2522 (N_2522,In_4309,In_2974);
nor U2523 (N_2523,N_1470,In_2015);
xor U2524 (N_2524,In_1543,N_1599);
nor U2525 (N_2525,N_1426,N_732);
xor U2526 (N_2526,In_2884,N_1253);
or U2527 (N_2527,N_1192,In_2778);
and U2528 (N_2528,N_1180,N_1000);
and U2529 (N_2529,N_906,N_1283);
or U2530 (N_2530,N_765,In_3836);
xnor U2531 (N_2531,N_1960,In_4422);
nor U2532 (N_2532,In_2820,N_1544);
nand U2533 (N_2533,In_1224,In_1225);
and U2534 (N_2534,N_852,In_1258);
or U2535 (N_2535,N_1486,In_1478);
xnor U2536 (N_2536,N_821,In_1966);
or U2537 (N_2537,N_1907,N_1597);
nand U2538 (N_2538,N_1968,N_1603);
nor U2539 (N_2539,In_4086,N_650);
nor U2540 (N_2540,N_1852,N_622);
or U2541 (N_2541,In_1579,N_1732);
or U2542 (N_2542,N_1929,In_240);
and U2543 (N_2543,In_3576,In_1691);
nor U2544 (N_2544,In_1861,N_1235);
nand U2545 (N_2545,N_1714,N_1248);
or U2546 (N_2546,In_4253,N_1473);
xnor U2547 (N_2547,In_1255,In_2914);
nand U2548 (N_2548,N_1533,In_4353);
xor U2549 (N_2549,N_467,N_968);
or U2550 (N_2550,In_827,In_1318);
nor U2551 (N_2551,In_112,In_1596);
nor U2552 (N_2552,In_26,N_1170);
nand U2553 (N_2553,N_284,N_1913);
nand U2554 (N_2554,N_643,N_1436);
and U2555 (N_2555,N_956,N_1923);
xor U2556 (N_2556,N_1619,N_1799);
and U2557 (N_2557,N_402,N_1120);
xnor U2558 (N_2558,N_1894,In_2093);
nor U2559 (N_2559,N_1510,N_1586);
xor U2560 (N_2560,In_2164,N_1194);
nor U2561 (N_2561,In_2013,N_1324);
and U2562 (N_2562,N_1430,In_2910);
xnor U2563 (N_2563,In_4096,In_4257);
nand U2564 (N_2564,In_1797,N_1788);
or U2565 (N_2565,In_3870,N_1164);
and U2566 (N_2566,N_1083,N_240);
and U2567 (N_2567,N_20,In_764);
xor U2568 (N_2568,In_1344,In_2877);
nand U2569 (N_2569,In_1964,In_4552);
nor U2570 (N_2570,In_4444,N_370);
nor U2571 (N_2571,N_1751,In_1324);
or U2572 (N_2572,N_1779,In_3098);
nand U2573 (N_2573,N_1321,N_1636);
nand U2574 (N_2574,N_187,In_679);
nor U2575 (N_2575,In_2363,In_1580);
or U2576 (N_2576,N_1277,N_1418);
nand U2577 (N_2577,N_1318,N_1804);
nand U2578 (N_2578,In_2601,In_1693);
xor U2579 (N_2579,N_1023,N_1853);
xnor U2580 (N_2580,N_1163,N_562);
xnor U2581 (N_2581,In_704,N_995);
nand U2582 (N_2582,N_392,In_3999);
xnor U2583 (N_2583,N_61,In_96);
or U2584 (N_2584,N_798,N_1405);
xnor U2585 (N_2585,N_1528,N_407);
nor U2586 (N_2586,In_4968,N_1360);
nor U2587 (N_2587,N_1027,In_2995);
nor U2588 (N_2588,In_683,In_3825);
nand U2589 (N_2589,N_466,In_4236);
and U2590 (N_2590,In_3398,In_4454);
nand U2591 (N_2591,In_961,In_3266);
nand U2592 (N_2592,In_514,N_1475);
and U2593 (N_2593,N_461,N_90);
or U2594 (N_2594,N_354,N_1420);
nor U2595 (N_2595,N_1140,N_1058);
nor U2596 (N_2596,In_3641,In_3414);
nor U2597 (N_2597,N_1602,N_642);
nor U2598 (N_2598,N_616,N_933);
xor U2599 (N_2599,N_1351,N_1449);
or U2600 (N_2600,N_1215,In_963);
nor U2601 (N_2601,N_670,N_715);
nor U2602 (N_2602,In_1316,In_2808);
nor U2603 (N_2603,In_4702,In_214);
or U2604 (N_2604,In_4059,In_4251);
nor U2605 (N_2605,In_4735,N_1269);
nor U2606 (N_2606,In_4331,N_1116);
and U2607 (N_2607,N_130,In_2382);
nor U2608 (N_2608,In_1197,In_428);
or U2609 (N_2609,In_1937,In_3413);
nor U2610 (N_2610,In_331,In_4023);
or U2611 (N_2611,N_1701,In_2795);
nor U2612 (N_2612,In_995,N_28);
nor U2613 (N_2613,N_1097,In_1965);
xnor U2614 (N_2614,In_53,N_1078);
xnor U2615 (N_2615,N_31,N_1173);
nor U2616 (N_2616,N_1374,In_740);
nand U2617 (N_2617,N_495,N_904);
xnor U2618 (N_2618,In_3834,N_1690);
nor U2619 (N_2619,In_2761,N_359);
nor U2620 (N_2620,In_4013,In_4771);
nand U2621 (N_2621,N_1631,In_868);
nor U2622 (N_2622,In_614,N_1046);
nor U2623 (N_2623,In_4631,N_1855);
or U2624 (N_2624,N_1188,In_2033);
or U2625 (N_2625,In_4778,In_905);
nor U2626 (N_2626,In_3761,In_4218);
nand U2627 (N_2627,In_4138,In_837);
nor U2628 (N_2628,N_678,N_43);
xnor U2629 (N_2629,In_534,N_293);
and U2630 (N_2630,In_665,In_4238);
or U2631 (N_2631,In_2149,In_2392);
or U2632 (N_2632,In_1053,In_2699);
nor U2633 (N_2633,In_1489,N_1285);
or U2634 (N_2634,N_1841,N_1680);
nand U2635 (N_2635,In_2141,N_350);
nand U2636 (N_2636,N_1353,N_1813);
nor U2637 (N_2637,In_2296,N_313);
xor U2638 (N_2638,In_252,In_3596);
xnor U2639 (N_2639,In_1421,N_1460);
nand U2640 (N_2640,N_1176,N_913);
xnor U2641 (N_2641,In_1375,N_512);
and U2642 (N_2642,In_3876,In_2004);
nand U2643 (N_2643,In_1338,In_3963);
or U2644 (N_2644,In_422,N_1560);
xnor U2645 (N_2645,In_3131,In_4655);
and U2646 (N_2646,N_824,In_2330);
xor U2647 (N_2647,N_1483,In_1755);
nor U2648 (N_2648,In_3886,N_1518);
nand U2649 (N_2649,N_1626,N_349);
nand U2650 (N_2650,In_559,In_2862);
nor U2651 (N_2651,In_1737,N_1867);
and U2652 (N_2652,In_3468,N_1925);
xor U2653 (N_2653,N_1984,In_4749);
and U2654 (N_2654,N_1184,In_2352);
xor U2655 (N_2655,N_443,In_2531);
and U2656 (N_2656,In_3902,In_902);
nor U2657 (N_2657,N_1370,In_2412);
or U2658 (N_2658,In_606,In_548);
or U2659 (N_2659,In_2827,N_1728);
xor U2660 (N_2660,In_4430,In_4252);
xor U2661 (N_2661,N_1365,N_1938);
nor U2662 (N_2662,N_1961,In_2721);
xor U2663 (N_2663,In_1761,N_626);
xor U2664 (N_2664,In_1684,In_4857);
nor U2665 (N_2665,N_1793,N_1810);
nand U2666 (N_2666,In_4060,In_236);
xor U2667 (N_2667,N_1851,In_3148);
and U2668 (N_2668,In_2419,N_1558);
xor U2669 (N_2669,N_1673,In_3476);
nor U2670 (N_2670,N_1270,N_318);
and U2671 (N_2671,In_2194,N_1381);
nand U2672 (N_2672,In_3994,In_3951);
xor U2673 (N_2673,N_1651,In_4889);
nand U2674 (N_2674,N_778,In_1400);
and U2675 (N_2675,In_1680,In_1615);
xor U2676 (N_2676,In_2839,In_4802);
and U2677 (N_2677,In_3735,In_2873);
nor U2678 (N_2678,In_2545,In_1439);
or U2679 (N_2679,N_1017,N_1963);
nand U2680 (N_2680,N_1857,N_1246);
nor U2681 (N_2681,In_1465,In_2237);
nand U2682 (N_2682,In_532,N_281);
or U2683 (N_2683,N_1286,In_1121);
nor U2684 (N_2684,In_2755,N_1329);
and U2685 (N_2685,In_4101,N_1369);
and U2686 (N_2686,In_4379,N_1141);
xor U2687 (N_2687,N_1834,N_1431);
xnor U2688 (N_2688,N_1258,In_2667);
nand U2689 (N_2689,In_30,N_1464);
nor U2690 (N_2690,In_3958,N_1545);
xor U2691 (N_2691,In_1766,N_725);
and U2692 (N_2692,N_1601,In_4994);
nand U2693 (N_2693,In_3240,In_2179);
xnor U2694 (N_2694,In_561,In_2815);
or U2695 (N_2695,N_1081,In_4289);
xnor U2696 (N_2696,In_1830,N_1313);
xnor U2697 (N_2697,N_369,N_1828);
nand U2698 (N_2698,N_1676,N_1214);
nor U2699 (N_2699,N_215,N_1296);
nand U2700 (N_2700,N_382,In_854);
and U2701 (N_2701,In_1976,N_62);
nor U2702 (N_2702,N_1686,N_1289);
or U2703 (N_2703,N_253,N_1276);
or U2704 (N_2704,In_4372,N_647);
nand U2705 (N_2705,N_1638,N_1983);
nor U2706 (N_2706,N_1415,N_1527);
nand U2707 (N_2707,In_1087,In_1517);
nand U2708 (N_2708,In_1638,In_1339);
nand U2709 (N_2709,In_1391,In_2674);
and U2710 (N_2710,In_881,N_1264);
nor U2711 (N_2711,N_959,In_3815);
and U2712 (N_2712,In_2766,N_1749);
xor U2713 (N_2713,N_1004,In_2727);
or U2714 (N_2714,In_4629,In_4048);
and U2715 (N_2715,In_1261,N_52);
nand U2716 (N_2716,In_1822,N_271);
xor U2717 (N_2717,N_1655,In_3236);
nand U2718 (N_2718,In_1450,N_1241);
and U2719 (N_2719,In_3304,N_212);
and U2720 (N_2720,In_4637,In_1790);
xnor U2721 (N_2721,N_1801,N_1945);
or U2722 (N_2722,In_3323,N_1540);
or U2723 (N_2723,N_1569,N_529);
xor U2724 (N_2724,N_1681,In_4775);
nand U2725 (N_2725,N_166,In_267);
xnor U2726 (N_2726,In_2180,N_1401);
nand U2727 (N_2727,N_416,N_332);
nor U2728 (N_2728,N_1490,In_1408);
xnor U2729 (N_2729,In_3260,N_770);
nand U2730 (N_2730,In_1770,N_673);
nor U2731 (N_2731,In_1306,In_4636);
nor U2732 (N_2732,N_1669,In_3960);
and U2733 (N_2733,In_1603,In_4409);
and U2734 (N_2734,N_1087,In_1911);
nor U2735 (N_2735,N_883,In_378);
or U2736 (N_2736,In_1801,In_2067);
and U2737 (N_2737,In_3861,In_4836);
nor U2738 (N_2738,In_1503,In_1842);
xor U2739 (N_2739,N_1856,N_808);
nand U2740 (N_2740,N_1231,In_3515);
xnor U2741 (N_2741,N_1346,In_1176);
and U2742 (N_2742,In_4149,N_1066);
nand U2743 (N_2743,In_554,In_255);
nor U2744 (N_2744,N_1428,N_1134);
or U2745 (N_2745,In_3919,In_2034);
nor U2746 (N_2746,In_2754,In_4510);
nor U2747 (N_2747,N_1877,In_4224);
nand U2748 (N_2748,N_1417,In_4204);
or U2749 (N_2749,N_1244,N_1931);
or U2750 (N_2750,N_649,In_3585);
or U2751 (N_2751,In_1583,In_4305);
nor U2752 (N_2752,N_1450,N_921);
and U2753 (N_2753,In_3136,In_3702);
or U2754 (N_2754,N_372,N_298);
xor U2755 (N_2755,N_1733,In_4323);
xnor U2756 (N_2756,In_460,N_1053);
nand U2757 (N_2757,In_3640,In_3851);
nand U2758 (N_2758,In_104,N_1844);
xnor U2759 (N_2759,In_3220,In_361);
xnor U2760 (N_2760,N_1908,N_660);
and U2761 (N_2761,N_1572,N_1049);
nand U2762 (N_2762,In_3093,In_690);
nor U2763 (N_2763,N_1920,In_2416);
nand U2764 (N_2764,N_1596,In_4113);
and U2765 (N_2765,In_3264,N_1317);
and U2766 (N_2766,In_2210,In_3592);
or U2767 (N_2767,In_3154,N_1635);
nand U2768 (N_2768,In_2861,In_4509);
xnor U2769 (N_2769,N_1385,N_1776);
nand U2770 (N_2770,In_4746,In_2031);
nor U2771 (N_2771,In_529,N_387);
or U2772 (N_2772,In_3095,N_738);
nor U2773 (N_2773,N_1137,N_277);
xor U2774 (N_2774,N_1829,N_3);
or U2775 (N_2775,N_756,N_1765);
nand U2776 (N_2776,N_1107,N_1606);
and U2777 (N_2777,In_954,In_853);
nor U2778 (N_2778,In_4446,N_1069);
nor U2779 (N_2779,N_1375,In_2780);
and U2780 (N_2780,N_1272,N_527);
nor U2781 (N_2781,In_3786,N_1612);
nor U2782 (N_2782,N_171,N_296);
xor U2783 (N_2783,N_1151,In_75);
nor U2784 (N_2784,N_473,N_1386);
or U2785 (N_2785,In_3429,N_1780);
nand U2786 (N_2786,N_1989,In_1417);
and U2787 (N_2787,In_3268,In_4583);
or U2788 (N_2788,N_322,N_1030);
xor U2789 (N_2789,N_125,In_1108);
or U2790 (N_2790,N_185,N_115);
and U2791 (N_2791,In_668,In_2249);
or U2792 (N_2792,N_1716,N_1796);
xor U2793 (N_2793,In_4515,In_362);
and U2794 (N_2794,N_839,N_478);
or U2795 (N_2795,N_1660,In_391);
nand U2796 (N_2796,In_2732,N_590);
and U2797 (N_2797,In_2825,N_1233);
or U2798 (N_2798,N_1666,N_908);
or U2799 (N_2799,N_1542,In_4016);
nand U2800 (N_2800,N_1126,In_1413);
nand U2801 (N_2801,N_1033,In_2055);
xnor U2802 (N_2802,N_246,In_396);
and U2803 (N_2803,In_3799,N_1332);
nor U2804 (N_2804,In_3819,N_610);
xor U2805 (N_2805,In_3707,N_363);
nor U2806 (N_2806,N_1973,N_1135);
nand U2807 (N_2807,N_1041,N_1467);
nor U2808 (N_2808,In_4780,In_2037);
and U2809 (N_2809,In_4201,In_2123);
nor U2810 (N_2810,In_358,In_4604);
nand U2811 (N_2811,In_633,N_726);
or U2812 (N_2812,N_385,N_1142);
or U2813 (N_2813,N_922,N_1693);
nor U2814 (N_2814,N_634,N_1893);
or U2815 (N_2815,In_2716,In_680);
and U2816 (N_2816,N_802,N_1530);
nand U2817 (N_2817,In_4739,N_174);
xor U2818 (N_2818,N_88,N_1005);
nand U2819 (N_2819,N_1858,In_500);
nor U2820 (N_2820,In_1021,N_1953);
nand U2821 (N_2821,In_763,N_1737);
or U2822 (N_2822,N_1730,N_1872);
or U2823 (N_2823,N_1196,N_621);
and U2824 (N_2824,N_1698,N_1843);
and U2825 (N_2825,In_2333,N_320);
or U2826 (N_2826,In_3608,In_2868);
xor U2827 (N_2827,N_605,N_935);
nand U2828 (N_2828,N_1391,N_1648);
and U2829 (N_2829,In_2129,N_1668);
xor U2830 (N_2830,In_2209,N_1899);
and U2831 (N_2831,In_2665,N_542);
xnor U2832 (N_2832,N_1439,N_523);
nand U2833 (N_2833,In_2515,N_275);
nor U2834 (N_2834,In_3283,In_3296);
xnor U2835 (N_2835,N_1037,N_1250);
nand U2836 (N_2836,In_1330,In_967);
nand U2837 (N_2837,N_654,In_3451);
nor U2838 (N_2838,In_1279,N_175);
xnor U2839 (N_2839,N_1797,In_324);
xor U2840 (N_2840,N_1098,In_4992);
nand U2841 (N_2841,N_1918,N_1564);
and U2842 (N_2842,In_1211,In_855);
nand U2843 (N_2843,N_985,In_2320);
xor U2844 (N_2844,In_2464,N_1302);
and U2845 (N_2845,In_692,In_2384);
nand U2846 (N_2846,In_3526,In_4002);
or U2847 (N_2847,In_696,In_1009);
nor U2848 (N_2848,In_2899,N_1282);
xnor U2849 (N_2849,In_2403,N_1139);
nor U2850 (N_2850,N_1696,N_425);
and U2851 (N_2851,In_155,In_1129);
xor U2852 (N_2852,In_747,N_1002);
or U2853 (N_2853,In_196,N_153);
nand U2854 (N_2854,N_1516,In_2988);
or U2855 (N_2855,N_1760,N_1577);
and U2856 (N_2856,In_4592,N_1106);
xor U2857 (N_2857,In_4146,In_4942);
xnor U2858 (N_2858,N_533,N_1390);
and U2859 (N_2859,In_3215,In_3143);
nand U2860 (N_2860,In_3078,N_575);
xor U2861 (N_2861,N_1397,In_3181);
and U2862 (N_2862,In_1011,N_578);
nor U2863 (N_2863,In_4649,In_4810);
nor U2864 (N_2864,In_733,In_1913);
nor U2865 (N_2865,In_4559,N_180);
or U2866 (N_2866,In_841,N_156);
xor U2867 (N_2867,N_123,N_1735);
xor U2868 (N_2868,In_1331,N_1099);
xnor U2869 (N_2869,N_158,In_4926);
xor U2870 (N_2870,N_868,N_1520);
nor U2871 (N_2871,N_1498,In_720);
xnor U2872 (N_2872,N_1238,In_3498);
or U2873 (N_2873,N_1766,N_1402);
or U2874 (N_2874,In_2882,N_701);
and U2875 (N_2875,N_487,N_1962);
nand U2876 (N_2876,N_1863,N_1559);
or U2877 (N_2877,N_1551,In_4743);
xor U2878 (N_2878,N_705,In_3070);
nand U2879 (N_2879,N_609,In_1509);
nand U2880 (N_2880,N_476,In_51);
xnor U2881 (N_2881,N_686,N_920);
or U2882 (N_2882,N_1278,N_814);
nand U2883 (N_2883,N_1543,N_1193);
nand U2884 (N_2884,N_1114,N_1649);
and U2885 (N_2885,In_2340,N_1711);
nand U2886 (N_2886,N_1366,N_1502);
nor U2887 (N_2887,N_1886,N_1566);
xor U2888 (N_2888,N_1379,N_1316);
nand U2889 (N_2889,In_2579,In_2151);
or U2890 (N_2890,N_1662,N_394);
and U2891 (N_2891,In_3848,In_1423);
or U2892 (N_2892,N_1909,N_1805);
nand U2893 (N_2893,In_3365,N_146);
or U2894 (N_2894,In_3812,N_1177);
or U2895 (N_2895,N_1144,In_4864);
xor U2896 (N_2896,In_3061,N_1456);
nand U2897 (N_2897,In_3972,In_4395);
or U2898 (N_2898,N_308,N_792);
xor U2899 (N_2899,In_2908,N_1136);
and U2900 (N_2900,N_314,In_3630);
nor U2901 (N_2901,In_1029,In_4214);
nand U2902 (N_2902,In_3235,N_749);
xor U2903 (N_2903,In_2842,N_1715);
nor U2904 (N_2904,In_1519,N_694);
nand U2905 (N_2905,In_2263,In_130);
nand U2906 (N_2906,In_1836,N_1311);
nand U2907 (N_2907,N_635,In_1715);
xnor U2908 (N_2908,N_818,N_1362);
xnor U2909 (N_2909,N_1371,N_1630);
and U2910 (N_2910,In_106,N_1836);
xnor U2911 (N_2911,N_1868,In_1903);
xor U2912 (N_2912,N_1532,In_3625);
or U2913 (N_2913,In_3359,In_2342);
nor U2914 (N_2914,In_1266,In_3777);
nor U2915 (N_2915,N_1924,In_1114);
and U2916 (N_2916,In_786,N_127);
or U2917 (N_2917,N_780,N_1427);
nor U2918 (N_2918,In_4920,N_1411);
xor U2919 (N_2919,N_919,N_1308);
nor U2920 (N_2920,In_3637,N_1132);
or U2921 (N_2921,N_671,In_1570);
nand U2922 (N_2922,In_3909,In_3127);
nand U2923 (N_2923,N_1018,N_1835);
or U2924 (N_2924,N_1364,In_703);
xnor U2925 (N_2925,In_1838,N_1513);
nand U2926 (N_2926,In_4068,N_1906);
or U2927 (N_2927,In_441,In_4692);
xor U2928 (N_2928,In_3444,N_1726);
xor U2929 (N_2929,N_502,N_1451);
nor U2930 (N_2930,N_789,N_429);
nand U2931 (N_2931,In_1351,N_897);
nor U2932 (N_2932,In_83,N_1717);
and U2933 (N_2933,N_1848,N_358);
nand U2934 (N_2934,In_256,In_2007);
xor U2935 (N_2935,In_4880,N_977);
and U2936 (N_2936,N_140,In_4343);
and U2937 (N_2937,N_746,In_2578);
xor U2938 (N_2938,N_1643,In_2488);
nand U2939 (N_2939,In_1877,N_1406);
and U2940 (N_2940,N_1123,N_1870);
and U2941 (N_2941,N_587,In_2157);
nor U2942 (N_2942,N_1609,In_4991);
nor U2943 (N_2943,N_996,In_178);
nor U2944 (N_2944,N_1016,In_189);
xnor U2945 (N_2945,N_1934,In_4157);
and U2946 (N_2946,In_1855,In_684);
xor U2947 (N_2947,In_1096,In_2063);
or U2948 (N_2948,N_589,In_2387);
and U2949 (N_2949,N_278,In_4872);
nor U2950 (N_2950,N_1396,N_1741);
xnor U2951 (N_2951,In_807,N_279);
nor U2952 (N_2952,N_1358,In_1933);
xor U2953 (N_2953,In_1885,In_2962);
nand U2954 (N_2954,N_1171,In_2956);
or U2955 (N_2955,N_676,In_3452);
nand U2956 (N_2956,N_1784,In_3046);
xor U2957 (N_2957,N_311,N_1511);
and U2958 (N_2958,In_1047,In_2378);
nand U2959 (N_2959,N_624,In_1771);
nand U2960 (N_2960,N_1682,N_1580);
or U2961 (N_2961,In_836,N_1959);
and U2962 (N_2962,N_1191,In_2069);
or U2963 (N_2963,N_1224,N_984);
nor U2964 (N_2964,In_3611,In_4547);
xor U2965 (N_2965,N_1937,N_1534);
and U2966 (N_2966,N_1775,In_2365);
or U2967 (N_2967,In_2208,In_3968);
or U2968 (N_2968,N_1512,In_3086);
nand U2969 (N_2969,N_1051,In_1088);
and U2970 (N_2970,In_776,N_1239);
and U2971 (N_2971,In_3482,N_1891);
and U2972 (N_2972,N_1816,In_1137);
xor U2973 (N_2973,N_1887,N_1299);
xnor U2974 (N_2974,N_470,In_1254);
and U2975 (N_2975,N_506,In_4083);
or U2976 (N_2976,In_2144,In_591);
nand U2977 (N_2977,In_949,N_210);
or U2978 (N_2978,N_1421,N_1125);
nand U2979 (N_2979,N_1090,In_3768);
or U2980 (N_2980,In_3106,In_3609);
nand U2981 (N_2981,N_1888,N_1499);
nand U2982 (N_2982,In_2372,N_1687);
or U2983 (N_2983,N_1849,N_1121);
xnor U2984 (N_2984,N_376,N_1675);
and U2985 (N_2985,In_1127,N_1723);
or U2986 (N_2986,N_383,In_4442);
xnor U2987 (N_2987,In_4094,In_3939);
nand U2988 (N_2988,In_191,In_506);
nand U2989 (N_2989,N_1138,In_4585);
xor U2990 (N_2990,N_823,In_122);
xnor U2991 (N_2991,N_337,In_811);
xnor U2992 (N_2992,In_3663,In_3019);
xnor U2993 (N_2993,In_4011,N_706);
or U2994 (N_2994,N_1885,In_4072);
and U2995 (N_2995,In_201,N_884);
nand U2996 (N_2996,In_3287,N_573);
nand U2997 (N_2997,N_1965,In_446);
and U2998 (N_2998,N_1288,N_282);
or U2999 (N_2999,N_1825,In_3382);
and U3000 (N_3000,In_481,N_1240);
and U3001 (N_3001,N_2086,In_2871);
or U3002 (N_3002,N_2936,In_4924);
and U3003 (N_3003,N_2476,N_1274);
nand U3004 (N_3004,N_2944,N_2829);
and U3005 (N_3005,N_2432,N_2817);
nor U3006 (N_3006,In_2829,In_4953);
nor U3007 (N_3007,N_2103,N_2460);
nand U3008 (N_3008,N_2478,N_2510);
nand U3009 (N_3009,In_1528,N_2990);
nor U3010 (N_3010,N_2243,N_2521);
nand U3011 (N_3011,In_3335,N_2917);
nor U3012 (N_3012,N_2662,N_1143);
nor U3013 (N_3013,N_2101,N_2902);
nand U3014 (N_3014,N_2104,N_14);
and U3015 (N_3015,N_2100,In_648);
or U3016 (N_3016,N_1076,In_3923);
nand U3017 (N_3017,N_2063,N_2151);
and U3018 (N_3018,N_195,N_2711);
nor U3019 (N_3019,In_4507,N_1201);
nor U3020 (N_3020,N_2287,In_4916);
or U3021 (N_3021,N_2660,N_2049);
and U3022 (N_3022,N_1219,N_2296);
or U3023 (N_3023,In_2446,N_2591);
xor U3024 (N_3024,N_2137,N_2208);
nand U3025 (N_3025,N_2938,N_2387);
or U3026 (N_3026,N_2447,N_1755);
or U3027 (N_3027,N_2642,In_1547);
nand U3028 (N_3028,N_2867,In_542);
nor U3029 (N_3029,N_2117,In_2148);
or U3030 (N_3030,In_3032,N_1245);
xor U3031 (N_3031,N_1072,In_3916);
or U3032 (N_3032,In_3540,N_2233);
or U3033 (N_3033,N_292,In_1829);
xor U3034 (N_3034,N_2808,N_1068);
xnor U3035 (N_3035,N_2009,In_1093);
xor U3036 (N_3036,N_2629,N_1291);
xnor U3037 (N_3037,N_2412,N_2628);
and U3038 (N_3038,N_244,N_2207);
nor U3039 (N_3039,N_2632,In_3571);
or U3040 (N_3040,N_2329,In_138);
or U3041 (N_3041,N_2027,N_2676);
and U3042 (N_3042,In_4208,N_1039);
nor U3043 (N_3043,In_3953,N_2949);
xnor U3044 (N_3044,N_2020,N_1524);
nand U3045 (N_3045,N_1947,N_1363);
xnor U3046 (N_3046,N_1013,N_2888);
nand U3047 (N_3047,In_3001,N_1781);
nor U3048 (N_3048,N_2220,In_85);
and U3049 (N_3049,In_61,N_2360);
xor U3050 (N_3050,N_2280,In_3150);
or U3051 (N_3051,N_2382,N_1424);
xnor U3052 (N_3052,In_2462,N_2038);
or U3053 (N_3053,N_1879,N_2173);
nor U3054 (N_3054,N_1593,N_2349);
or U3055 (N_3055,In_4683,In_4324);
xnor U3056 (N_3056,N_633,N_810);
nor U3057 (N_3057,N_2406,N_924);
and U3058 (N_3058,N_2758,N_1915);
xnor U3059 (N_3059,N_2164,In_586);
or U3060 (N_3060,N_2171,N_2706);
xnor U3061 (N_3061,N_2718,In_264);
nor U3062 (N_3062,N_1488,N_2709);
or U3063 (N_3063,N_2022,N_2627);
and U3064 (N_3064,In_1619,N_2446);
xnor U3065 (N_3065,N_430,N_2177);
nor U3066 (N_3066,In_2702,N_2974);
or U3067 (N_3067,N_2697,N_1897);
nand U3068 (N_3068,N_2138,In_3927);
or U3069 (N_3069,N_2963,N_1325);
and U3070 (N_3070,N_1491,N_2548);
xor U3071 (N_3071,N_2440,In_1069);
xor U3072 (N_3072,N_1933,N_2331);
or U3073 (N_3073,N_2862,N_2613);
and U3074 (N_3074,N_2269,N_1659);
xnor U3075 (N_3075,In_792,In_2217);
nor U3076 (N_3076,N_662,N_2864);
xnor U3077 (N_3077,N_2572,N_1382);
nand U3078 (N_3078,N_1777,N_2680);
nand U3079 (N_3079,In_2422,N_1035);
or U3080 (N_3080,In_146,N_2705);
and U3081 (N_3081,N_528,N_418);
or U3082 (N_3082,N_1113,N_2108);
xor U3083 (N_3083,In_555,N_2954);
or U3084 (N_3084,N_2928,N_1484);
nand U3085 (N_3085,In_2166,N_779);
nand U3086 (N_3086,N_2153,In_4037);
xnor U3087 (N_3087,N_698,N_2135);
xnor U3088 (N_3088,N_2519,N_216);
xor U3089 (N_3089,N_126,In_2629);
xnor U3090 (N_3090,In_2467,N_431);
or U3091 (N_3091,In_1232,In_3280);
or U3092 (N_3092,N_1373,In_4038);
xnor U3093 (N_3093,N_2362,N_2893);
or U3094 (N_3094,In_2693,N_2212);
nor U3095 (N_3095,N_836,N_2696);
xor U3096 (N_3096,N_2007,N_2877);
xnor U3097 (N_3097,In_3555,N_2409);
and U3098 (N_3098,N_2487,In_2666);
nor U3099 (N_3099,N_2782,N_1958);
and U3100 (N_3100,N_2453,N_2196);
xor U3101 (N_3101,In_257,N_1203);
nor U3102 (N_3102,N_2005,N_2126);
or U3103 (N_3103,N_2694,N_1895);
nor U3104 (N_3104,N_2326,In_4965);
or U3105 (N_3105,N_2725,In_2247);
nand U3106 (N_3106,N_2700,N_103);
xnor U3107 (N_3107,In_2200,N_1562);
nor U3108 (N_3108,N_1865,N_2116);
xor U3109 (N_3109,N_2604,N_2494);
or U3110 (N_3110,N_1926,In_766);
xor U3111 (N_3111,N_2091,N_1957);
nor U3112 (N_3112,N_2544,N_2710);
and U3113 (N_3113,In_1399,N_444);
or U3114 (N_3114,N_2707,N_2757);
xnor U3115 (N_3115,N_1105,N_2348);
or U3116 (N_3116,N_1174,N_2573);
nand U3117 (N_3117,N_2770,N_2788);
nor U3118 (N_3118,In_1147,N_2532);
and U3119 (N_3119,In_526,N_2607);
or U3120 (N_3120,In_3654,In_2319);
nand U3121 (N_3121,In_1538,N_2375);
and U3122 (N_3122,N_1943,N_1725);
nand U3123 (N_3123,In_4185,N_2363);
xor U3124 (N_3124,In_2241,N_2291);
or U3125 (N_3125,N_2737,N_2467);
and U3126 (N_3126,In_4284,N_2797);
nand U3127 (N_3127,N_2899,In_917);
nand U3128 (N_3128,N_2549,N_1331);
nor U3129 (N_3129,N_2730,N_2389);
nor U3130 (N_3130,N_550,N_2225);
nand U3131 (N_3131,In_1701,N_1257);
nand U3132 (N_3132,N_2475,N_1927);
nor U3133 (N_3133,In_4927,N_1446);
nor U3134 (N_3134,N_2300,N_2777);
or U3135 (N_3135,N_2172,N_2567);
nand U3136 (N_3136,N_2581,In_3528);
nor U3137 (N_3137,N_1949,N_832);
xnor U3138 (N_3138,N_77,N_1040);
and U3139 (N_3139,N_2297,N_2392);
and U3140 (N_3140,N_63,N_2449);
nor U3141 (N_3141,In_4153,N_2044);
and U3142 (N_3142,In_415,N_2477);
and U3143 (N_3143,N_237,N_2169);
nand U3144 (N_3144,N_474,N_1538);
nor U3145 (N_3145,N_2538,In_193);
or U3146 (N_3146,N_2570,In_1924);
nor U3147 (N_3147,N_2000,N_2920);
xor U3148 (N_3148,N_2474,N_1505);
xor U3149 (N_3149,In_2580,N_2751);
nand U3150 (N_3150,N_2952,N_2930);
and U3151 (N_3151,N_2084,N_2926);
xor U3152 (N_3152,N_2377,In_4015);
nor U3153 (N_3153,In_2558,In_1109);
or U3154 (N_3154,N_1469,In_144);
and U3155 (N_3155,In_541,N_1702);
or U3156 (N_3156,N_2771,N_2011);
xor U3157 (N_3157,N_2623,N_2796);
or U3158 (N_3158,N_2418,N_2371);
xor U3159 (N_3159,N_931,N_1561);
nand U3160 (N_3160,N_2735,N_2699);
xnor U3161 (N_3161,N_2579,In_510);
and U3162 (N_3162,In_2999,In_2452);
or U3163 (N_3163,N_1459,In_4337);
xnor U3164 (N_3164,N_2809,N_2593);
nand U3165 (N_3165,N_2030,N_2033);
or U3166 (N_3166,In_3415,N_2969);
nor U3167 (N_3167,N_1359,N_1807);
nor U3168 (N_3168,N_2583,N_2051);
or U3169 (N_3169,N_2551,N_1045);
and U3170 (N_3170,In_3312,In_3720);
nand U3171 (N_3171,N_2436,N_2041);
and U3172 (N_3172,N_2812,N_2332);
nor U3173 (N_3173,N_2983,N_131);
nor U3174 (N_3174,N_2790,N_2271);
and U3175 (N_3175,In_4182,In_4844);
nand U3176 (N_3176,N_2987,In_287);
nor U3177 (N_3177,N_1695,In_4184);
and U3178 (N_3178,N_1089,N_1355);
or U3179 (N_3179,N_147,N_2299);
or U3180 (N_3180,N_2045,N_2150);
nor U3181 (N_3181,N_2931,In_4750);
nor U3182 (N_3182,In_2664,N_2353);
xor U3183 (N_3183,N_347,In_863);
nand U3184 (N_3184,N_2281,In_4457);
and U3185 (N_3185,N_2290,In_4560);
xnor U3186 (N_3186,In_4009,N_2828);
nand U3187 (N_3187,N_2076,In_990);
and U3188 (N_3188,N_2292,N_2070);
nand U3189 (N_3189,In_2474,In_4199);
nor U3190 (N_3190,In_2427,N_2155);
or U3191 (N_3191,In_2318,N_2247);
nand U3192 (N_3192,N_2719,N_1901);
and U3193 (N_3193,N_2994,N_2999);
nor U3194 (N_3194,N_2541,N_1057);
and U3195 (N_3195,N_2740,N_2772);
nand U3196 (N_3196,N_2473,N_2922);
xnor U3197 (N_3197,N_2731,N_2789);
nor U3198 (N_3198,N_2012,N_1115);
xor U3199 (N_3199,In_694,In_3224);
nand U3200 (N_3200,N_549,N_519);
and U3201 (N_3201,In_1124,N_2679);
nand U3202 (N_3202,N_2596,N_1287);
xnor U3203 (N_3203,In_4982,In_1544);
xnor U3204 (N_3204,N_2034,N_2262);
nand U3205 (N_3205,N_1070,In_3883);
and U3206 (N_3206,N_2183,N_2664);
nor U3207 (N_3207,N_2860,N_2261);
nand U3208 (N_3208,N_2993,N_2461);
and U3209 (N_3209,N_2639,N_2932);
nor U3210 (N_3210,In_3722,In_232);
or U3211 (N_3211,In_4582,N_2924);
nand U3212 (N_3212,N_2161,N_2756);
or U3213 (N_3213,N_2869,N_1216);
and U3214 (N_3214,N_2352,N_1026);
nand U3215 (N_3215,N_1111,In_1574);
or U3216 (N_3216,In_1929,N_2337);
nor U3217 (N_3217,In_4145,In_3579);
nand U3218 (N_3218,In_3097,N_2163);
nand U3219 (N_3219,N_2982,N_1129);
and U3220 (N_3220,N_1657,N_2585);
and U3221 (N_3221,N_1380,N_2335);
and U3222 (N_3222,N_2124,In_681);
or U3223 (N_3223,N_2956,N_2470);
nand U3224 (N_3224,N_1146,N_2955);
or U3225 (N_3225,N_2558,N_2940);
or U3226 (N_3226,In_2045,N_2031);
or U3227 (N_3227,N_1700,N_1672);
or U3228 (N_3228,N_2463,N_2535);
and U3229 (N_3229,In_1907,N_2942);
xnor U3230 (N_3230,N_877,N_1474);
nor U3231 (N_3231,N_2425,N_2444);
xor U3232 (N_3232,N_1684,N_2658);
xor U3233 (N_3233,N_2260,N_2037);
or U3234 (N_3234,N_2612,N_2139);
nand U3235 (N_3235,In_1310,In_4638);
and U3236 (N_3236,N_1345,N_2654);
xor U3237 (N_3237,In_847,N_1574);
nor U3238 (N_3238,N_2670,N_1585);
nor U3239 (N_3239,N_2638,N_2438);
or U3240 (N_3240,N_2222,In_4408);
xnor U3241 (N_3241,N_2681,N_1147);
xnor U3242 (N_3242,N_1830,N_1442);
or U3243 (N_3243,N_2397,N_1200);
and U3244 (N_3244,N_2511,In_2647);
or U3245 (N_3245,N_2754,N_2166);
nor U3246 (N_3246,N_2239,N_2646);
and U3247 (N_3247,N_2911,N_2966);
nand U3248 (N_3248,N_1225,N_2121);
or U3249 (N_3249,In_3984,N_2170);
and U3250 (N_3250,N_2376,N_1537);
nand U3251 (N_3251,In_4043,N_2776);
xor U3252 (N_3252,N_2350,N_1145);
nor U3253 (N_3253,N_878,N_1752);
or U3254 (N_3254,In_3205,N_2912);
and U3255 (N_3255,In_1685,N_2385);
nor U3256 (N_3256,In_4173,N_72);
nor U3257 (N_3257,N_239,N_2102);
or U3258 (N_3258,N_1372,N_2824);
and U3259 (N_3259,In_1605,N_2971);
nor U3260 (N_3260,N_74,N_2148);
nor U3261 (N_3261,N_2464,N_1800);
xor U3262 (N_3262,N_2825,N_2663);
or U3263 (N_3263,In_1751,N_2768);
or U3264 (N_3264,In_1269,In_4245);
and U3265 (N_3265,In_1480,In_3711);
xnor U3266 (N_3266,N_2373,N_2048);
or U3267 (N_3267,N_1230,N_2424);
and U3268 (N_3268,N_454,In_2226);
or U3269 (N_3269,In_2789,N_2534);
or U3270 (N_3270,N_2159,N_2357);
nand U3271 (N_3271,N_2462,N_1595);
or U3272 (N_3272,N_2480,N_2914);
nor U3273 (N_3273,N_2318,N_532);
nor U3274 (N_3274,N_2405,In_2298);
xnor U3275 (N_3275,N_2687,In_164);
nand U3276 (N_3276,In_2496,In_1950);
and U3277 (N_3277,N_1228,In_4286);
nand U3278 (N_3278,N_2420,N_2741);
nor U3279 (N_3279,In_504,N_2764);
xor U3280 (N_3280,In_2393,N_1871);
or U3281 (N_3281,N_2372,N_1769);
xnor U3282 (N_3282,N_2635,N_2620);
nand U3283 (N_3283,N_2514,In_3250);
nand U3284 (N_3284,N_49,In_2066);
or U3285 (N_3285,In_4030,N_1024);
and U3286 (N_3286,N_65,In_2805);
or U3287 (N_3287,N_2267,In_3156);
xnor U3288 (N_3288,In_4781,N_1086);
nand U3289 (N_3289,N_2489,N_2616);
xnor U3290 (N_3290,N_1563,N_2245);
xnor U3291 (N_3291,N_2039,N_2445);
xor U3292 (N_3292,N_2113,N_2619);
or U3293 (N_3293,In_3841,N_2913);
or U3294 (N_3294,N_2105,N_2844);
nor U3295 (N_3295,In_3186,N_845);
or U3296 (N_3296,N_2813,In_3137);
or U3297 (N_3297,N_2490,In_4890);
nor U3298 (N_3298,In_174,In_4706);
or U3299 (N_3299,N_2324,In_4807);
and U3300 (N_3300,In_4007,N_2647);
nand U3301 (N_3301,N_472,N_2129);
nand U3302 (N_3302,In_2881,N_830);
and U3303 (N_3303,N_1869,N_2677);
nor U3304 (N_3304,In_432,In_1396);
nor U3305 (N_3305,In_95,N_2237);
and U3306 (N_3306,N_2400,N_954);
xor U3307 (N_3307,N_1892,N_2252);
nand U3308 (N_3308,N_2204,In_3309);
or U3309 (N_3309,In_1730,N_2122);
or U3310 (N_3310,In_2424,N_2546);
xor U3311 (N_3311,N_2133,In_2685);
and U3312 (N_3312,N_2555,N_2174);
or U3313 (N_3313,N_1555,N_2206);
nor U3314 (N_3314,In_975,N_1985);
nand U3315 (N_3315,N_1743,N_2584);
nand U3316 (N_3316,N_2689,N_2253);
xnor U3317 (N_3317,In_1867,N_717);
nand U3318 (N_3318,N_2053,N_2626);
and U3319 (N_3319,N_2904,N_1904);
or U3320 (N_3320,N_2423,N_2562);
nor U3321 (N_3321,N_2115,N_2650);
or U3322 (N_3322,N_2734,N_2634);
nand U3323 (N_3323,N_2118,In_228);
nor U3324 (N_3324,N_366,N_1220);
nand U3325 (N_3325,N_2780,In_304);
nor U3326 (N_3326,In_3432,N_2242);
or U3327 (N_3327,N_2656,In_781);
nand U3328 (N_3328,In_4292,N_999);
or U3329 (N_3329,In_501,N_2671);
or U3330 (N_3330,N_1128,In_1484);
nor U3331 (N_3331,N_2152,N_773);
nor U3332 (N_3332,N_2112,N_2419);
and U3333 (N_3333,In_3478,In_1321);
and U3334 (N_3334,N_1506,In_279);
nand U3335 (N_3335,In_4804,In_3931);
nand U3336 (N_3336,N_2998,In_4447);
nor U3337 (N_3337,In_3481,N_2036);
nand U3338 (N_3338,N_1010,In_1993);
nand U3339 (N_3339,N_2431,N_114);
nand U3340 (N_3340,N_2224,In_1239);
nand U3341 (N_3341,N_2801,N_1531);
nor U3342 (N_3342,N_2783,In_3906);
xor U3343 (N_3343,In_562,In_4863);
xor U3344 (N_3344,In_2423,N_1917);
or U3345 (N_3345,N_887,N_907);
xnor U3346 (N_3346,In_3605,N_2945);
nor U3347 (N_3347,N_2875,N_1110);
or U3348 (N_3348,N_2536,In_1565);
nor U3349 (N_3349,N_2608,N_2781);
or U3350 (N_3350,In_604,N_2722);
xor U3351 (N_3351,In_563,N_2190);
xnor U3352 (N_3352,N_2810,N_2678);
nor U3353 (N_3353,N_2618,N_2182);
or U3354 (N_3354,N_2525,N_2897);
nor U3355 (N_3355,N_2492,N_2586);
nor U3356 (N_3356,N_2894,N_2876);
xnor U3357 (N_3357,N_1328,N_1582);
nor U3358 (N_3358,In_4537,N_2228);
nand U3359 (N_3359,In_3403,N_2601);
xnor U3360 (N_3360,In_3175,N_2313);
xor U3361 (N_3361,N_2563,N_2219);
nor U3362 (N_3362,N_2767,In_342);
or U3363 (N_3363,N_2211,In_4200);
xnor U3364 (N_3364,N_2187,N_1773);
nor U3365 (N_3365,N_1423,N_1404);
nor U3366 (N_3366,N_2733,In_4821);
nand U3367 (N_3367,N_2417,N_198);
or U3368 (N_3368,N_2580,N_1047);
nand U3369 (N_3369,N_2441,N_2553);
nand U3370 (N_3370,N_2975,N_513);
xnor U3371 (N_3371,N_2319,In_4329);
and U3372 (N_3372,In_2441,N_2197);
or U3373 (N_3373,In_3600,N_1453);
nor U3374 (N_3374,N_398,N_2637);
or U3375 (N_3375,N_1734,N_2625);
and U3376 (N_3376,N_1222,N_2046);
or U3377 (N_3377,N_1011,In_3014);
nor U3378 (N_3378,N_2249,N_2374);
or U3379 (N_3379,N_2804,N_1036);
nand U3380 (N_3380,N_2811,N_1665);
and U3381 (N_3381,N_2042,N_2799);
nor U3382 (N_3382,N_1912,N_2341);
xor U3383 (N_3383,N_2976,N_2631);
xnor U3384 (N_3384,N_2970,N_541);
nor U3385 (N_3385,N_56,In_1039);
xor U3386 (N_3386,In_1773,In_3855);
and U3387 (N_3387,In_451,In_2571);
and U3388 (N_3388,N_2408,N_2130);
or U3389 (N_3389,In_2904,N_2846);
or U3390 (N_3390,N_1305,N_266);
xnor U3391 (N_3391,N_1539,N_2855);
nor U3392 (N_3392,N_2919,N_591);
and U3393 (N_3393,N_548,N_2753);
nand U3394 (N_3394,N_1759,N_1052);
or U3395 (N_3395,In_2457,In_1637);
nand U3396 (N_3396,N_2752,In_3192);
nand U3397 (N_3397,N_2448,N_1309);
or U3398 (N_3398,N_412,N_2359);
and U3399 (N_3399,N_2140,N_2098);
and U3400 (N_3400,N_2131,N_2369);
xnor U3401 (N_3401,In_1240,N_2857);
nor U3402 (N_3402,N_2191,N_2826);
xor U3403 (N_3403,N_1247,N_2069);
xor U3404 (N_3404,N_2488,N_1575);
xor U3405 (N_3405,N_2491,N_2256);
or U3406 (N_3406,N_1333,N_2024);
nand U3407 (N_3407,N_2089,N_2468);
xnor U3408 (N_3408,N_1352,In_2088);
xor U3409 (N_3409,N_1546,N_1565);
or U3410 (N_3410,N_2910,In_4261);
or U3411 (N_3411,N_2981,In_412);
xor U3412 (N_3412,N_981,N_2984);
nand U3413 (N_3413,N_2391,N_2147);
or U3414 (N_3414,N_2240,N_2072);
nand U3415 (N_3415,In_3554,N_2507);
or U3416 (N_3416,N_2229,In_4801);
and U3417 (N_3417,In_4714,In_3065);
xnor U3418 (N_3418,N_2818,N_434);
and U3419 (N_3419,In_3351,N_1487);
nand U3420 (N_3420,In_4469,N_2395);
or U3421 (N_3421,N_2578,In_1557);
or U3422 (N_3422,N_2014,N_2640);
nand U3423 (N_3423,N_2393,N_534);
and U3424 (N_3424,In_2818,In_1563);
and U3425 (N_3425,N_2394,In_1532);
nor U3426 (N_3426,N_2435,N_875);
nand U3427 (N_3427,N_439,N_2272);
and U3428 (N_3428,N_2889,N_2437);
xnor U3429 (N_3429,N_2339,N_2843);
xor U3430 (N_3430,N_1229,N_2427);
nand U3431 (N_3431,N_1890,N_2325);
nor U3432 (N_3432,N_2872,N_2653);
xor U3433 (N_3433,N_1689,N_2892);
or U3434 (N_3434,N_1523,N_2673);
or U3435 (N_3435,N_993,N_2834);
nor U3436 (N_3436,In_1444,N_2992);
and U3437 (N_3437,N_1103,In_2743);
nor U3438 (N_3438,In_977,In_2192);
and U3439 (N_3439,In_1208,N_2890);
or U3440 (N_3440,N_1377,In_3189);
nand U3441 (N_3441,In_1987,N_2188);
xnor U3442 (N_3442,N_2035,N_2516);
and U3443 (N_3443,In_753,N_2274);
nor U3444 (N_3444,N_2901,N_89);
nor U3445 (N_3445,N_2588,In_4313);
nor U3446 (N_3446,N_37,N_1003);
nor U3447 (N_3447,N_2564,In_2440);
xor U3448 (N_3448,N_2749,N_2617);
nand U3449 (N_3449,In_1268,N_2017);
or U3450 (N_3450,In_1508,N_2962);
nor U3451 (N_3451,In_797,In_239);
xnor U3452 (N_3452,N_976,N_2643);
nor U3453 (N_3453,N_2661,In_3425);
nor U3454 (N_3454,N_2870,N_2455);
xor U3455 (N_3455,N_2403,N_1661);
and U3456 (N_3456,In_3983,N_2672);
nor U3457 (N_3457,In_2147,In_4635);
or U3458 (N_3458,N_2214,N_2763);
and U3459 (N_3459,N_2343,N_2156);
xor U3460 (N_3460,N_2951,N_2960);
nand U3461 (N_3461,N_1854,N_11);
and U3462 (N_3462,N_2023,N_2077);
or U3463 (N_3463,N_1503,N_2937);
xor U3464 (N_3464,In_4795,In_4876);
nor U3465 (N_3465,N_2311,In_1389);
xor U3466 (N_3466,N_2837,In_1757);
nor U3467 (N_3467,In_2048,N_1761);
or U3468 (N_3468,N_1059,N_2314);
or U3469 (N_3469,In_1007,In_1300);
nor U3470 (N_3470,N_2266,In_4721);
or U3471 (N_3471,N_1525,In_1996);
nor U3472 (N_3472,N_1162,N_2645);
or U3473 (N_3473,N_2871,N_1261);
and U3474 (N_3474,N_395,N_2315);
and U3475 (N_3475,N_2160,N_2849);
xnor U3476 (N_3476,In_162,N_490);
nand U3477 (N_3477,N_682,In_4680);
or U3478 (N_3478,In_289,In_774);
nand U3479 (N_3479,N_2941,In_1655);
or U3480 (N_3480,N_2574,N_2095);
nor U3481 (N_3481,In_4382,N_942);
and U3482 (N_3482,In_4049,In_2600);
and U3483 (N_3483,N_2667,N_2513);
nor U3484 (N_3484,N_2298,In_1889);
nor U3485 (N_3485,N_2896,N_2606);
xor U3486 (N_3486,N_2127,In_109);
or U3487 (N_3487,N_766,In_1668);
nor U3488 (N_3488,In_4728,N_1218);
or U3489 (N_3489,In_3814,In_4401);
nand U3490 (N_3490,N_2675,N_2905);
nor U3491 (N_3491,N_2702,N_2471);
or U3492 (N_3492,N_2481,N_1979);
nor U3493 (N_3493,In_1769,N_2270);
nor U3494 (N_3494,In_1186,N_2433);
xnor U3495 (N_3495,N_2110,N_2785);
or U3496 (N_3496,In_3449,In_4440);
xnor U3497 (N_3497,N_2304,N_1795);
and U3498 (N_3498,N_155,N_2316);
and U3499 (N_3499,N_2342,In_3159);
or U3500 (N_3500,N_1591,N_2230);
and U3501 (N_3501,N_388,N_2985);
or U3502 (N_3502,In_1101,In_207);
xnor U3503 (N_3503,In_3770,In_1188);
and U3504 (N_3504,N_568,N_2050);
or U3505 (N_3505,In_108,N_2980);
nor U3506 (N_3506,N_1692,N_2961);
xnor U3507 (N_3507,N_2947,In_276);
xor U3508 (N_3508,N_2057,In_2759);
or U3509 (N_3509,N_2176,N_2879);
or U3510 (N_3510,N_2028,In_4047);
and U3511 (N_3511,In_1299,N_896);
or U3512 (N_3512,In_2343,N_2361);
or U3513 (N_3513,N_1179,N_2995);
or U3514 (N_3514,N_2334,N_2762);
or U3515 (N_3515,N_1383,N_2502);
xnor U3516 (N_3516,N_1398,N_1022);
or U3517 (N_3517,In_3390,In_4707);
or U3518 (N_3518,N_2071,N_2178);
xor U3519 (N_3519,N_2010,N_2257);
and U3520 (N_3520,N_1798,N_2598);
xor U3521 (N_3521,N_1928,N_2713);
nand U3522 (N_3522,N_2775,In_4858);
xnor U3523 (N_3523,N_2651,N_2399);
nand U3524 (N_3524,N_1747,N_2997);
or U3525 (N_3525,N_2184,N_2365);
nand U3526 (N_3526,N_1604,N_2263);
xor U3527 (N_3527,N_2388,N_2655);
and U3528 (N_3528,N_1429,N_2231);
or U3529 (N_3529,In_3581,In_3917);
nand U3530 (N_3530,N_2761,N_2096);
nor U3531 (N_3531,N_2531,N_2692);
nand U3532 (N_3532,In_3588,In_4527);
nor U3533 (N_3533,N_1817,In_2335);
and U3534 (N_3534,In_4364,N_2093);
or U3535 (N_3535,In_226,In_3937);
or U3536 (N_3536,In_2544,N_2726);
xnor U3537 (N_3537,In_3226,N_2125);
nand U3538 (N_3538,N_2136,N_2241);
and U3539 (N_3539,N_669,N_2943);
or U3540 (N_3540,N_1930,N_2175);
xor U3541 (N_3541,In_4546,N_2246);
and U3542 (N_3542,N_2097,N_1395);
or U3543 (N_3543,N_2720,N_1691);
xor U3544 (N_3544,N_1122,N_2891);
and U3545 (N_3545,N_1818,N_2732);
nand U3546 (N_3546,N_2554,N_2223);
and U3547 (N_3547,N_2986,N_2001);
xor U3548 (N_3548,N_1187,In_2779);
xnor U3549 (N_3549,N_2279,In_3193);
and U3550 (N_3550,N_1517,In_4700);
xnor U3551 (N_3551,N_2590,In_3345);
xor U3552 (N_3552,N_1889,N_2194);
nand U3553 (N_3553,N_2512,N_2347);
xnor U3554 (N_3554,In_1099,N_1832);
xor U3555 (N_3555,N_2275,N_1862);
nand U3556 (N_3556,N_2186,N_2404);
and U3557 (N_3557,N_2833,N_2518);
nor U3558 (N_3558,In_4272,N_2144);
xor U3559 (N_3559,In_1758,In_1205);
and U3560 (N_3560,N_2285,In_3802);
or U3561 (N_3561,N_2411,N_2456);
and U3562 (N_3562,N_1823,N_1354);
or U3563 (N_3563,N_1579,N_2430);
nor U3564 (N_3564,N_1213,N_2556);
nor U3565 (N_3565,N_2958,N_456);
xor U3566 (N_3566,N_2273,N_2547);
or U3567 (N_3567,In_3541,In_3737);
and U3568 (N_3568,N_2868,N_2201);
nand U3569 (N_3569,N_2227,N_2141);
nor U3570 (N_3570,N_2873,N_2923);
and U3571 (N_3571,N_1785,N_2308);
xnor U3572 (N_3572,In_3807,In_809);
xor U3573 (N_3573,N_2909,In_3754);
nand U3574 (N_3574,In_1564,N_2193);
xnor U3575 (N_3575,N_1881,In_330);
xnor U3576 (N_3576,N_2765,In_2314);
and U3577 (N_3577,N_863,In_1793);
or U3578 (N_3578,In_612,N_2216);
nand U3579 (N_3579,N_2496,N_234);
or U3580 (N_3580,N_2146,N_2577);
xnor U3581 (N_3581,In_2025,N_360);
nand U3582 (N_3582,N_2021,N_2557);
nor U3583 (N_3583,N_2309,N_2221);
or U3584 (N_3584,N_2600,N_1608);
or U3585 (N_3585,In_1294,N_2484);
and U3586 (N_3586,N_1182,N_2466);
or U3587 (N_3587,N_2939,In_3868);
or U3588 (N_3588,N_2384,N_1064);
xor U3589 (N_3589,In_3173,N_2859);
and U3590 (N_3590,In_1616,N_2294);
nor U3591 (N_3591,In_2341,N_2605);
or U3592 (N_3592,N_23,In_4572);
or U3593 (N_3593,In_2079,N_831);
and U3594 (N_3594,N_1639,N_2244);
nor U3595 (N_3595,N_2968,N_2317);
or U3596 (N_3596,N_1905,N_2043);
nand U3597 (N_3597,In_1158,N_2712);
or U3598 (N_3598,N_2996,N_2964);
or U3599 (N_3599,N_2948,N_2192);
xnor U3600 (N_3600,N_264,N_1757);
and U3601 (N_3601,N_2495,In_1348);
xnor U3602 (N_3602,N_2927,N_2668);
or U3603 (N_3603,N_2040,N_2064);
or U3604 (N_3604,In_2875,N_2524);
or U3605 (N_3605,N_2209,N_2321);
nor U3606 (N_3606,N_488,N_2259);
and U3607 (N_3607,N_2288,N_2906);
and U3608 (N_3608,N_2254,N_2268);
or U3609 (N_3609,N_625,N_507);
or U3610 (N_3610,N_2845,In_808);
nor U3611 (N_3611,N_2469,In_4081);
nor U3612 (N_3612,N_2898,In_1646);
or U3613 (N_3613,In_1831,N_2052);
xor U3614 (N_3614,N_2539,N_139);
nor U3615 (N_3615,N_2957,N_2443);
or U3616 (N_3616,In_2655,N_2738);
nand U3617 (N_3617,N_1697,N_2003);
and U3618 (N_3618,N_1679,N_2199);
or U3619 (N_3619,N_1975,In_636);
or U3620 (N_3620,N_2682,N_2836);
and U3621 (N_3621,In_98,N_2886);
nand U3622 (N_3622,N_2615,N_1808);
nor U3623 (N_3623,N_2887,N_1334);
nor U3624 (N_3624,N_1472,In_1765);
nor U3625 (N_3625,N_1465,N_2847);
nor U3626 (N_3626,In_2078,N_1088);
nor U3627 (N_3627,N_2840,N_2908);
nand U3628 (N_3628,N_2185,N_73);
nand U3629 (N_3629,N_2442,N_1477);
xnor U3630 (N_3630,N_2238,N_2203);
xnor U3631 (N_3631,N_2465,N_2132);
xnor U3632 (N_3632,N_2258,N_2058);
xor U3633 (N_3633,N_2526,N_503);
and U3634 (N_3634,In_3216,N_1159);
and U3635 (N_3635,In_1817,In_3875);
nand U3636 (N_3636,In_1704,N_2413);
and U3637 (N_3637,N_815,N_288);
nor U3638 (N_3638,In_3164,In_2130);
and U3639 (N_3639,N_2533,N_2282);
nor U3640 (N_3640,N_2742,N_2454);
xnor U3641 (N_3641,N_1304,N_2791);
nand U3642 (N_3642,In_4244,N_2265);
nor U3643 (N_3643,N_1742,N_2597);
and U3644 (N_3644,N_2232,N_1811);
and U3645 (N_3645,In_936,N_2119);
nand U3646 (N_3646,N_1634,In_86);
xor U3647 (N_3647,N_2307,N_1744);
nor U3648 (N_3648,N_1280,N_2641);
xnor U3649 (N_3649,In_2233,N_1312);
nor U3650 (N_3650,N_1186,N_2065);
and U3651 (N_3651,N_2701,N_2289);
and U3652 (N_3652,N_1294,N_2745);
nor U3653 (N_3653,N_2426,In_2541);
nor U3654 (N_3654,N_1995,N_2784);
nand U3655 (N_3655,N_1814,N_2323);
and U3656 (N_3656,N_1942,N_2472);
nor U3657 (N_3657,N_2415,N_1826);
and U3658 (N_3658,In_2050,N_2895);
and U3659 (N_3659,N_2013,N_2946);
nand U3660 (N_3660,N_2421,N_1536);
nand U3661 (N_3661,In_4134,N_2085);
nor U3662 (N_3662,N_2189,In_3282);
nor U3663 (N_3663,N_2509,In_2919);
or U3664 (N_3664,N_1185,N_396);
xnor U3665 (N_3665,In_2799,N_2614);
nor U3666 (N_3666,In_3362,In_2295);
or U3667 (N_3667,N_309,N_2565);
nand U3668 (N_3668,In_1192,N_2396);
nand U3669 (N_3669,In_151,N_2120);
xnor U3670 (N_3670,In_536,N_1323);
nor U3671 (N_3671,N_2882,In_2375);
or U3672 (N_3672,In_1775,In_4466);
and U3673 (N_3673,N_2002,N_1972);
nand U3674 (N_3674,N_663,N_2842);
xor U3675 (N_3675,N_1754,In_509);
and U3676 (N_3676,N_2061,N_2458);
or U3677 (N_3677,N_1042,N_2099);
nand U3678 (N_3678,N_2595,In_2843);
nand U3679 (N_3679,N_1756,N_1878);
nor U3680 (N_3680,N_2814,In_1368);
nor U3681 (N_3681,N_2721,In_4489);
nor U3682 (N_3682,N_357,In_1031);
or U3683 (N_3683,N_2226,N_2611);
nand U3684 (N_3684,N_1152,N_2723);
nand U3685 (N_3685,In_4303,N_2755);
and U3686 (N_3686,In_3901,N_1394);
or U3687 (N_3687,In_4614,N_2434);
nand U3688 (N_3688,N_2560,In_2610);
or U3689 (N_3689,N_2950,N_331);
and U3690 (N_3690,In_2136,N_2935);
nand U3691 (N_3691,In_3271,N_1167);
or U3692 (N_3692,N_1082,In_4133);
nand U3693 (N_3693,N_2428,N_2505);
and U3694 (N_3694,In_3198,N_1547);
xor U3695 (N_3695,In_2577,N_2766);
xnor U3696 (N_3696,In_1832,N_2747);
nor U3697 (N_3697,N_2881,N_2778);
and U3698 (N_3698,N_2959,N_2370);
xnor U3699 (N_3699,N_2109,N_894);
nand U3700 (N_3700,N_2769,N_2819);
nor U3701 (N_3701,N_104,N_1729);
nor U3702 (N_3702,N_2863,N_2589);
xnor U3703 (N_3703,N_1227,N_2714);
xor U3704 (N_3704,In_1888,N_1295);
xor U3705 (N_3705,In_738,In_2673);
and U3706 (N_3706,N_2149,N_2883);
and U3707 (N_3707,N_1541,N_2306);
xor U3708 (N_3708,N_2180,N_1632);
nor U3709 (N_3709,N_2674,N_1724);
and U3710 (N_3710,N_2165,N_2856);
xnor U3711 (N_3711,N_1842,N_2832);
xnor U3712 (N_3712,N_1640,In_4263);
and U3713 (N_3713,In_2414,N_2355);
nor U3714 (N_3714,N_1667,N_1653);
nand U3715 (N_3715,In_4766,N_2630);
or U3716 (N_3716,N_1028,N_299);
nand U3717 (N_3717,N_83,In_2609);
and U3718 (N_3718,N_2967,In_2872);
or U3719 (N_3719,N_537,N_1452);
or U3720 (N_3720,In_793,In_2592);
xor U3721 (N_3721,In_3831,N_2386);
nand U3722 (N_3722,In_4354,N_2015);
xor U3723 (N_3723,N_733,N_2530);
and U3724 (N_3724,N_2622,N_2340);
xor U3725 (N_3725,N_805,N_2277);
and U3726 (N_3726,In_2596,N_769);
nand U3727 (N_3727,N_2398,In_706);
xor U3728 (N_3728,In_3804,N_2006);
nand U3729 (N_3729,In_4260,N_2018);
and U3730 (N_3730,N_2143,In_3064);
nand U3731 (N_3731,N_861,N_2286);
or U3732 (N_3732,N_2312,N_2062);
and U3733 (N_3733,N_2523,N_315);
nand U3734 (N_3734,N_2047,In_2909);
xor U3735 (N_3735,N_2142,N_2402);
nor U3736 (N_3736,N_927,N_1594);
or U3737 (N_3737,N_2569,In_2259);
and U3738 (N_3738,N_258,N_2691);
nor U3739 (N_3739,N_2545,In_2773);
or U3740 (N_3740,N_1210,N_775);
and U3741 (N_3741,N_2885,N_2179);
or U3742 (N_3742,In_2091,N_1392);
or U3743 (N_3743,N_2695,N_2566);
nor U3744 (N_3744,N_1092,N_2621);
nor U3745 (N_3745,N_1629,N_1268);
nor U3746 (N_3746,N_2841,In_2951);
and U3747 (N_3747,N_1199,In_1220);
nor U3748 (N_3748,N_2503,N_1790);
nor U3749 (N_3749,N_2026,N_2786);
or U3750 (N_3750,N_1866,N_2380);
nand U3751 (N_3751,In_1865,N_2773);
nand U3752 (N_3752,In_2311,In_3123);
nand U3753 (N_3753,N_1043,N_2333);
xnor U3754 (N_3754,N_2060,N_2008);
xor U3755 (N_3755,N_2322,N_2787);
nor U3756 (N_3756,N_2167,N_2527);
xor U3757 (N_3757,N_2884,N_1637);
and U3758 (N_3758,In_887,N_2497);
or U3759 (N_3759,N_2234,N_2302);
xnor U3760 (N_3760,N_928,N_2016);
or U3761 (N_3761,N_1685,In_4210);
xnor U3762 (N_3762,N_1251,In_1166);
nand U3763 (N_3763,In_3424,N_1217);
and U3764 (N_3764,N_1168,N_1077);
nor U3765 (N_3765,N_2528,In_2931);
nor U3766 (N_3766,N_2979,N_2746);
xor U3767 (N_3767,N_1898,In_133);
nand U3768 (N_3768,N_2537,N_2851);
nor U3769 (N_3769,In_1703,N_2145);
or U3770 (N_3770,N_2485,N_2092);
xnor U3771 (N_3771,In_524,N_2529);
xor U3772 (N_3772,In_4516,N_2202);
nand U3773 (N_3773,N_1753,In_300);
nand U3774 (N_3774,In_1597,N_2128);
nand U3775 (N_3775,In_244,N_2114);
nand U3776 (N_3776,In_2669,N_2724);
or U3777 (N_3777,N_2750,N_2900);
xor U3778 (N_3778,N_2798,N_2205);
and U3779 (N_3779,N_2800,N_2075);
and U3780 (N_3780,N_1300,In_1873);
nor U3781 (N_3781,In_852,N_2068);
xnor U3782 (N_3782,N_2345,In_3651);
or U3783 (N_3783,N_1504,N_2988);
xnor U3784 (N_3784,N_142,N_1770);
or U3785 (N_3785,N_1976,N_2451);
xnor U3786 (N_3786,N_1815,In_225);
and U3787 (N_3787,N_2744,In_3898);
or U3788 (N_3788,N_2381,N_60);
xor U3789 (N_3789,N_2977,N_657);
nand U3790 (N_3790,N_2083,N_2822);
and U3791 (N_3791,In_4748,In_1671);
xor U3792 (N_3792,N_1124,N_2559);
xor U3793 (N_3793,N_1900,N_2915);
and U3794 (N_3794,N_2793,N_2933);
nor U3795 (N_3795,N_1789,N_1936);
and U3796 (N_3796,In_1681,In_4405);
or U3797 (N_3797,N_982,N_1951);
nor U3798 (N_3798,N_2978,N_1967);
nor U3799 (N_3799,N_1481,N_2728);
nor U3800 (N_3800,In_3694,N_2688);
or U3801 (N_3801,N_2501,In_18);
and U3802 (N_3802,N_540,In_1810);
or U3803 (N_3803,N_2716,N_2452);
nand U3804 (N_3804,N_2255,N_420);
nor U3805 (N_3805,In_55,N_2264);
xor U3806 (N_3806,N_2594,N_2522);
xor U3807 (N_3807,N_1400,N_1074);
nand U3808 (N_3808,In_2265,N_410);
xnor U3809 (N_3809,N_2652,N_2106);
or U3810 (N_3810,N_2520,In_2202);
xnor U3811 (N_3811,In_303,N_1021);
and U3812 (N_3812,N_2310,In_21);
nand U3813 (N_3813,N_1009,In_3141);
or U3814 (N_3814,N_2835,N_2078);
xnor U3815 (N_3815,N_1946,N_2390);
xor U3816 (N_3816,N_2739,N_2508);
and U3817 (N_3817,In_2573,N_2874);
nor U3818 (N_3818,In_2385,In_1506);
nor U3819 (N_3819,N_2379,N_2934);
and U3820 (N_3820,N_2094,N_2080);
and U3821 (N_3821,N_2367,N_1339);
and U3822 (N_3822,N_2479,N_2759);
or U3823 (N_3823,In_598,N_2055);
xor U3824 (N_3824,N_2748,N_1303);
or U3825 (N_3825,N_1254,N_1102);
or U3826 (N_3826,N_2561,N_2802);
or U3827 (N_3827,N_2698,N_1940);
and U3828 (N_3828,In_603,N_2213);
xnor U3829 (N_3829,In_2692,N_2366);
nand U3830 (N_3830,N_2351,N_1642);
nand U3831 (N_3831,N_2284,N_2729);
xnor U3832 (N_3832,N_2633,In_3874);
xor U3833 (N_3833,N_2158,N_2378);
or U3834 (N_3834,N_1722,N_242);
or U3835 (N_3835,N_2820,In_2120);
xor U3836 (N_3836,In_1988,In_2329);
nor U3837 (N_3837,N_2736,In_1328);
or U3838 (N_3838,N_1183,N_1029);
nand U3839 (N_3839,N_2486,N_1554);
nor U3840 (N_3840,N_2181,N_2907);
and U3841 (N_3841,N_2703,In_3115);
nor U3842 (N_3842,N_2327,N_1521);
nand U3843 (N_3843,N_2368,N_2659);
or U3844 (N_3844,In_466,N_1706);
xnor U3845 (N_3845,N_2683,N_2708);
xnor U3846 (N_3846,N_2669,N_2025);
and U3847 (N_3847,In_2283,N_2838);
xnor U3848 (N_3848,N_2081,N_2295);
xnor U3849 (N_3849,N_2929,N_2649);
nor U3850 (N_3850,N_2157,N_2356);
nor U3851 (N_3851,N_2853,N_2803);
nor U3852 (N_3852,N_2079,In_2864);
nor U3853 (N_3853,In_4062,N_639);
or U3854 (N_3854,N_2301,In_4769);
xor U3855 (N_3855,N_1845,In_3796);
and U3856 (N_3856,In_1272,N_2195);
nand U3857 (N_3857,N_2815,N_2218);
nor U3858 (N_3858,N_2235,In_4276);
nor U3859 (N_3859,In_1063,N_2991);
and U3860 (N_3860,N_679,In_2277);
nor U3861 (N_3861,N_2704,N_2794);
xnor U3862 (N_3862,N_2056,N_2107);
nor U3863 (N_3863,N_2168,N_2482);
and U3864 (N_3864,N_2576,N_1071);
xnor U3865 (N_3865,N_2603,N_1840);
nor U3866 (N_3866,In_1875,N_2401);
or U3867 (N_3867,N_2278,N_1063);
and U3868 (N_3868,N_2989,In_1604);
nor U3869 (N_3869,In_4805,In_3962);
nand U3870 (N_3870,In_88,N_2540);
xor U3871 (N_3871,N_1570,N_2439);
nand U3872 (N_3872,In_4819,N_2499);
and U3873 (N_3873,N_2416,In_333);
or U3874 (N_3874,N_2821,N_250);
and U3875 (N_3875,N_2250,N_594);
nand U3876 (N_3876,In_2905,N_964);
or U3877 (N_3877,N_1259,N_1507);
nor U3878 (N_3878,N_833,N_2953);
xnor U3879 (N_3879,N_1266,In_2874);
or U3880 (N_3880,N_1348,In_3850);
nand U3881 (N_3881,N_2568,N_1552);
nor U3882 (N_3882,N_2457,N_1731);
and U3883 (N_3883,N_2305,In_1037);
xnor U3884 (N_3884,N_2624,N_2921);
xnor U3885 (N_3885,In_3564,In_4020);
or U3886 (N_3886,N_988,N_2090);
or U3887 (N_3887,In_2986,N_2795);
or U3888 (N_3888,N_2866,In_3790);
or U3889 (N_3889,N_2925,In_457);
or U3890 (N_3890,N_1255,N_2123);
xor U3891 (N_3891,In_4755,N_1986);
xor U3892 (N_3892,N_1149,N_2200);
nor U3893 (N_3893,N_1713,N_2410);
and U3894 (N_3894,In_1977,N_2666);
and U3895 (N_3895,N_59,N_1119);
and U3896 (N_3896,In_1980,N_1130);
xor U3897 (N_3897,N_2665,N_2019);
and U3898 (N_3898,N_2422,N_2850);
xor U3899 (N_3899,N_1839,In_2804);
nand U3900 (N_3900,N_2338,N_2609);
and U3901 (N_3901,N_2717,N_2684);
or U3902 (N_3902,N_2727,N_2074);
and U3903 (N_3903,In_3381,N_2657);
nand U3904 (N_3904,N_1627,N_1492);
or U3905 (N_3905,N_2210,N_569);
and U3906 (N_3906,In_1587,N_2217);
xnor U3907 (N_3907,N_623,N_2571);
nor U3908 (N_3908,N_504,N_1455);
xnor U3909 (N_3909,N_2599,N_2830);
or U3910 (N_3910,N_1549,In_3820);
nor U3911 (N_3911,In_1026,N_2575);
nor U3912 (N_3912,N_598,N_2543);
nor U3913 (N_3913,N_1950,In_2425);
nand U3914 (N_3914,N_41,N_2854);
nand U3915 (N_3915,N_2715,N_2504);
nand U3916 (N_3916,N_777,N_2276);
nor U3917 (N_3917,N_2582,N_2865);
and U3918 (N_3918,In_3299,N_2407);
or U3919 (N_3919,In_787,In_2597);
and U3920 (N_3920,N_1335,In_3905);
and U3921 (N_3921,N_2602,N_2831);
nor U3922 (N_3922,N_1208,N_2358);
or U3923 (N_3923,N_2162,N_2066);
and U3924 (N_3924,In_641,N_2054);
xnor U3925 (N_3925,N_2861,N_336);
and U3926 (N_3926,N_2032,N_1721);
and U3927 (N_3927,N_809,N_2483);
or U3928 (N_3928,N_1786,N_2493);
and U3929 (N_3929,N_2459,N_2743);
or U3930 (N_3930,N_613,N_2330);
nor U3931 (N_3931,N_2429,In_3176);
xor U3932 (N_3932,N_168,N_2515);
nand U3933 (N_3933,N_2644,In_3356);
xor U3934 (N_3934,In_4064,N_1425);
or U3935 (N_3935,N_2774,N_241);
or U3936 (N_3936,N_2383,N_2498);
and U3937 (N_3937,N_2215,N_2336);
or U3938 (N_3938,N_1838,N_304);
nand U3939 (N_3939,N_2610,N_2328);
nor U3940 (N_3940,N_2806,N_2816);
and U3941 (N_3941,N_2198,N_2779);
xor U3942 (N_3942,N_2506,N_2134);
nand U3943 (N_3943,In_3199,N_2636);
or U3944 (N_3944,N_1249,In_3806);
or U3945 (N_3945,In_1720,N_2965);
or U3946 (N_3946,N_2517,N_2111);
nor U3947 (N_3947,In_1060,N_2792);
nand U3948 (N_3948,N_2587,N_2073);
xor U3949 (N_3949,N_2690,N_2693);
nor U3950 (N_3950,N_2087,N_2251);
nor U3951 (N_3951,N_2500,N_2852);
nor U3952 (N_3952,N_1320,In_4451);
nor U3953 (N_3953,N_95,N_2880);
nand U3954 (N_3954,In_1287,In_1015);
xnor U3955 (N_3955,In_2503,In_1149);
or U3956 (N_3956,N_2364,In_2534);
or U3957 (N_3957,N_2685,In_1925);
xor U3958 (N_3958,N_1094,In_4930);
or U3959 (N_3959,In_1362,In_439);
or U3960 (N_3960,N_1480,N_1297);
or U3961 (N_3961,In_4271,N_1050);
nor U3962 (N_3962,N_772,In_2454);
nand U3963 (N_3963,N_2973,N_2648);
and U3964 (N_3964,In_4050,N_2029);
or U3965 (N_3965,N_692,N_225);
or U3966 (N_3966,N_2550,In_503);
xor U3967 (N_3967,N_716,N_2346);
nand U3968 (N_3968,N_957,N_2760);
xnor U3969 (N_3969,N_2858,N_2823);
or U3970 (N_3970,N_1252,N_1500);
nand U3971 (N_3971,In_3784,N_222);
nand U3972 (N_3972,In_1811,In_1514);
and U3973 (N_3973,N_1190,N_1178);
nor U3974 (N_3974,N_2248,In_2653);
xor U3975 (N_3975,N_2918,N_1447);
xnor U3976 (N_3976,N_1350,N_817);
nand U3977 (N_3977,In_1241,N_2414);
nand U3978 (N_3978,N_1399,N_1884);
nand U3979 (N_3979,In_687,N_2686);
xor U3980 (N_3980,N_2059,N_2916);
and U3981 (N_3981,N_2805,In_3347);
or U3982 (N_3982,N_384,In_1518);
or U3983 (N_3983,N_2807,N_2827);
or U3984 (N_3984,N_1583,N_2839);
and U3985 (N_3985,N_2354,In_3210);
xor U3986 (N_3986,N_2088,N_1699);
xor U3987 (N_3987,N_1581,N_2542);
or U3988 (N_3988,N_2552,N_690);
xnor U3989 (N_3989,In_4632,N_2320);
xor U3990 (N_3990,N_2450,In_4458);
xnor U3991 (N_3991,In_1753,N_2293);
or U3992 (N_3992,N_2878,N_943);
nor U3993 (N_3993,N_2154,N_46);
xnor U3994 (N_3994,N_2004,N_2344);
or U3995 (N_3995,N_2903,N_2592);
nand U3996 (N_3996,N_2972,N_2067);
nor U3997 (N_3997,N_2303,N_2848);
and U3998 (N_3998,N_2082,N_2283);
xnor U3999 (N_3999,N_2236,N_1148);
nand U4000 (N_4000,N_3804,N_3653);
and U4001 (N_4001,N_3089,N_3142);
nor U4002 (N_4002,N_3594,N_3879);
nand U4003 (N_4003,N_3004,N_3450);
nand U4004 (N_4004,N_3467,N_3953);
nand U4005 (N_4005,N_3486,N_3494);
and U4006 (N_4006,N_3152,N_3661);
xnor U4007 (N_4007,N_3917,N_3565);
nor U4008 (N_4008,N_3331,N_3814);
and U4009 (N_4009,N_3086,N_3737);
or U4010 (N_4010,N_3791,N_3122);
or U4011 (N_4011,N_3926,N_3548);
or U4012 (N_4012,N_3023,N_3051);
and U4013 (N_4013,N_3537,N_3931);
nand U4014 (N_4014,N_3861,N_3496);
nand U4015 (N_4015,N_3560,N_3934);
nor U4016 (N_4016,N_3924,N_3526);
or U4017 (N_4017,N_3624,N_3267);
and U4018 (N_4018,N_3962,N_3612);
and U4019 (N_4019,N_3769,N_3501);
or U4020 (N_4020,N_3754,N_3874);
xnor U4021 (N_4021,N_3684,N_3725);
nand U4022 (N_4022,N_3100,N_3401);
xnor U4023 (N_4023,N_3113,N_3415);
nor U4024 (N_4024,N_3973,N_3287);
nand U4025 (N_4025,N_3951,N_3421);
nor U4026 (N_4026,N_3060,N_3822);
and U4027 (N_4027,N_3422,N_3026);
nor U4028 (N_4028,N_3283,N_3741);
nor U4029 (N_4029,N_3108,N_3528);
xor U4030 (N_4030,N_3904,N_3079);
and U4031 (N_4031,N_3495,N_3868);
and U4032 (N_4032,N_3226,N_3286);
or U4033 (N_4033,N_3853,N_3660);
or U4034 (N_4034,N_3682,N_3590);
and U4035 (N_4035,N_3617,N_3667);
xnor U4036 (N_4036,N_3271,N_3567);
and U4037 (N_4037,N_3394,N_3115);
nand U4038 (N_4038,N_3043,N_3112);
xnor U4039 (N_4039,N_3125,N_3857);
and U4040 (N_4040,N_3118,N_3309);
and U4041 (N_4041,N_3852,N_3451);
or U4042 (N_4042,N_3938,N_3120);
and U4043 (N_4043,N_3793,N_3045);
nand U4044 (N_4044,N_3825,N_3101);
or U4045 (N_4045,N_3581,N_3418);
nand U4046 (N_4046,N_3257,N_3965);
and U4047 (N_4047,N_3385,N_3550);
xor U4048 (N_4048,N_3666,N_3475);
or U4049 (N_4049,N_3747,N_3453);
and U4050 (N_4050,N_3497,N_3658);
nor U4051 (N_4051,N_3439,N_3430);
or U4052 (N_4052,N_3021,N_3277);
nor U4053 (N_4053,N_3176,N_3241);
and U4054 (N_4054,N_3894,N_3716);
nand U4055 (N_4055,N_3136,N_3899);
nand U4056 (N_4056,N_3790,N_3687);
nor U4057 (N_4057,N_3227,N_3464);
xnor U4058 (N_4058,N_3855,N_3523);
nor U4059 (N_4059,N_3189,N_3573);
or U4060 (N_4060,N_3970,N_3145);
xor U4061 (N_4061,N_3155,N_3950);
and U4062 (N_4062,N_3379,N_3482);
or U4063 (N_4063,N_3760,N_3144);
nor U4064 (N_4064,N_3163,N_3206);
nor U4065 (N_4065,N_3476,N_3847);
nor U4066 (N_4066,N_3440,N_3443);
or U4067 (N_4067,N_3381,N_3696);
or U4068 (N_4068,N_3400,N_3748);
and U4069 (N_4069,N_3956,N_3818);
or U4070 (N_4070,N_3355,N_3895);
or U4071 (N_4071,N_3353,N_3382);
nor U4072 (N_4072,N_3489,N_3012);
nand U4073 (N_4073,N_3196,N_3200);
or U4074 (N_4074,N_3637,N_3763);
nand U4075 (N_4075,N_3310,N_3469);
nand U4076 (N_4076,N_3745,N_3568);
nand U4077 (N_4077,N_3860,N_3961);
nor U4078 (N_4078,N_3557,N_3691);
or U4079 (N_4079,N_3941,N_3339);
nand U4080 (N_4080,N_3519,N_3220);
and U4081 (N_4081,N_3466,N_3036);
nand U4082 (N_4082,N_3638,N_3527);
nand U4083 (N_4083,N_3799,N_3222);
xor U4084 (N_4084,N_3652,N_3608);
xor U4085 (N_4085,N_3963,N_3877);
and U4086 (N_4086,N_3240,N_3369);
nor U4087 (N_4087,N_3412,N_3077);
and U4088 (N_4088,N_3727,N_3246);
or U4089 (N_4089,N_3001,N_3172);
and U4090 (N_4090,N_3531,N_3105);
nand U4091 (N_4091,N_3645,N_3611);
nor U4092 (N_4092,N_3920,N_3997);
or U4093 (N_4093,N_3362,N_3303);
or U4094 (N_4094,N_3305,N_3230);
or U4095 (N_4095,N_3485,N_3761);
or U4096 (N_4096,N_3280,N_3873);
nand U4097 (N_4097,N_3830,N_3459);
nand U4098 (N_4098,N_3796,N_3915);
and U4099 (N_4099,N_3455,N_3368);
nand U4100 (N_4100,N_3037,N_3209);
or U4101 (N_4101,N_3933,N_3297);
nand U4102 (N_4102,N_3985,N_3840);
nand U4103 (N_4103,N_3989,N_3402);
nor U4104 (N_4104,N_3504,N_3503);
or U4105 (N_4105,N_3162,N_3153);
nand U4106 (N_4106,N_3185,N_3561);
nand U4107 (N_4107,N_3929,N_3746);
and U4108 (N_4108,N_3649,N_3069);
nor U4109 (N_4109,N_3210,N_3304);
xnor U4110 (N_4110,N_3884,N_3699);
nor U4111 (N_4111,N_3870,N_3740);
and U4112 (N_4112,N_3204,N_3484);
xnor U4113 (N_4113,N_3056,N_3701);
nand U4114 (N_4114,N_3221,N_3111);
and U4115 (N_4115,N_3018,N_3274);
nand U4116 (N_4116,N_3039,N_3128);
or U4117 (N_4117,N_3614,N_3435);
and U4118 (N_4118,N_3330,N_3392);
nand U4119 (N_4119,N_3493,N_3578);
nor U4120 (N_4120,N_3646,N_3092);
and U4121 (N_4121,N_3733,N_3738);
nand U4122 (N_4122,N_3511,N_3832);
xnor U4123 (N_4123,N_3999,N_3454);
nor U4124 (N_4124,N_3258,N_3423);
and U4125 (N_4125,N_3972,N_3964);
or U4126 (N_4126,N_3046,N_3078);
or U4127 (N_4127,N_3481,N_3815);
xnor U4128 (N_4128,N_3869,N_3157);
nand U4129 (N_4129,N_3803,N_3165);
xnor U4130 (N_4130,N_3471,N_3095);
and U4131 (N_4131,N_3199,N_3584);
and U4132 (N_4132,N_3768,N_3912);
xor U4133 (N_4133,N_3538,N_3446);
nor U4134 (N_4134,N_3097,N_3647);
or U4135 (N_4135,N_3452,N_3959);
and U4136 (N_4136,N_3328,N_3117);
nor U4137 (N_4137,N_3758,N_3170);
or U4138 (N_4138,N_3005,N_3689);
and U4139 (N_4139,N_3872,N_3937);
or U4140 (N_4140,N_3576,N_3032);
nand U4141 (N_4141,N_3014,N_3679);
xnor U4142 (N_4142,N_3618,N_3838);
xor U4143 (N_4143,N_3556,N_3384);
xnor U4144 (N_4144,N_3621,N_3308);
xor U4145 (N_4145,N_3087,N_3426);
nor U4146 (N_4146,N_3845,N_3413);
nor U4147 (N_4147,N_3698,N_3514);
and U4148 (N_4148,N_3648,N_3875);
or U4149 (N_4149,N_3098,N_3913);
nor U4150 (N_4150,N_3789,N_3925);
nor U4151 (N_4151,N_3835,N_3859);
xor U4152 (N_4152,N_3694,N_3784);
nor U4153 (N_4153,N_3072,N_3901);
or U4154 (N_4154,N_3752,N_3948);
or U4155 (N_4155,N_3013,N_3191);
or U4156 (N_4156,N_3225,N_3133);
and U4157 (N_4157,N_3891,N_3311);
nor U4158 (N_4158,N_3148,N_3329);
nand U4159 (N_4159,N_3544,N_3290);
and U4160 (N_4160,N_3756,N_3600);
xor U4161 (N_4161,N_3295,N_3842);
or U4162 (N_4162,N_3492,N_3547);
or U4163 (N_4163,N_3778,N_3135);
and U4164 (N_4164,N_3881,N_3187);
or U4165 (N_4165,N_3823,N_3893);
xor U4166 (N_4166,N_3202,N_3301);
xor U4167 (N_4167,N_3850,N_3316);
nor U4168 (N_4168,N_3766,N_3674);
nor U4169 (N_4169,N_3505,N_3055);
nor U4170 (N_4170,N_3319,N_3837);
and U4171 (N_4171,N_3942,N_3866);
or U4172 (N_4172,N_3688,N_3035);
nand U4173 (N_4173,N_3588,N_3030);
xor U4174 (N_4174,N_3006,N_3644);
or U4175 (N_4175,N_3597,N_3007);
or U4176 (N_4176,N_3816,N_3553);
nor U4177 (N_4177,N_3432,N_3054);
or U4178 (N_4178,N_3864,N_3786);
xnor U4179 (N_4179,N_3071,N_3448);
and U4180 (N_4180,N_3254,N_3211);
nand U4181 (N_4181,N_3031,N_3817);
nor U4182 (N_4182,N_3273,N_3143);
or U4183 (N_4183,N_3958,N_3833);
nand U4184 (N_4184,N_3201,N_3347);
nand U4185 (N_4185,N_3671,N_3247);
nand U4186 (N_4186,N_3554,N_3093);
nor U4187 (N_4187,N_3487,N_3902);
nor U4188 (N_4188,N_3322,N_3935);
nand U4189 (N_4189,N_3009,N_3166);
nand U4190 (N_4190,N_3395,N_3708);
or U4191 (N_4191,N_3218,N_3512);
or U4192 (N_4192,N_3722,N_3320);
nand U4193 (N_4193,N_3123,N_3141);
nand U4194 (N_4194,N_3357,N_3260);
xor U4195 (N_4195,N_3288,N_3178);
nor U4196 (N_4196,N_3358,N_3558);
or U4197 (N_4197,N_3132,N_3490);
nor U4198 (N_4198,N_3593,N_3508);
xor U4199 (N_4199,N_3704,N_3721);
nor U4200 (N_4200,N_3672,N_3203);
and U4201 (N_4201,N_3718,N_3000);
and U4202 (N_4202,N_3217,N_3744);
nand U4203 (N_4203,N_3628,N_3762);
and U4204 (N_4204,N_3299,N_3307);
and U4205 (N_4205,N_3373,N_3800);
or U4206 (N_4206,N_3387,N_3739);
or U4207 (N_4207,N_3783,N_3654);
nand U4208 (N_4208,N_3944,N_3545);
and U4209 (N_4209,N_3234,N_3865);
nor U4210 (N_4210,N_3582,N_3264);
nor U4211 (N_4211,N_3732,N_3268);
nand U4212 (N_4212,N_3083,N_3161);
or U4213 (N_4213,N_3619,N_3836);
nand U4214 (N_4214,N_3116,N_3294);
and U4215 (N_4215,N_3910,N_3957);
nand U4216 (N_4216,N_3237,N_3880);
xnor U4217 (N_4217,N_3839,N_3188);
nor U4218 (N_4218,N_3723,N_3930);
or U4219 (N_4219,N_3546,N_3411);
and U4220 (N_4220,N_3470,N_3785);
nand U4221 (N_4221,N_3575,N_3911);
or U4222 (N_4222,N_3552,N_3641);
nor U4223 (N_4223,N_3040,N_3285);
nor U4224 (N_4224,N_3383,N_3428);
nor U4225 (N_4225,N_3376,N_3088);
nor U4226 (N_4226,N_3673,N_3720);
or U4227 (N_4227,N_3326,N_3946);
nand U4228 (N_4228,N_3434,N_3397);
or U4229 (N_4229,N_3982,N_3772);
and U4230 (N_4230,N_3080,N_3140);
nor U4231 (N_4231,N_3350,N_3406);
nor U4232 (N_4232,N_3726,N_3235);
nand U4233 (N_4233,N_3313,N_3248);
or U4234 (N_4234,N_3794,N_3729);
xor U4235 (N_4235,N_3626,N_3896);
nand U4236 (N_4236,N_3498,N_3947);
and U4237 (N_4237,N_3332,N_3377);
nand U4238 (N_4238,N_3341,N_3306);
or U4239 (N_4239,N_3564,N_3625);
xor U4240 (N_4240,N_3813,N_3675);
nor U4241 (N_4241,N_3524,N_3971);
nor U4242 (N_4242,N_3407,N_3502);
or U4243 (N_4243,N_3713,N_3765);
and U4244 (N_4244,N_3585,N_3966);
and U4245 (N_4245,N_3344,N_3577);
nand U4246 (N_4246,N_3650,N_3085);
and U4247 (N_4247,N_3134,N_3167);
nor U4248 (N_4248,N_3927,N_3690);
or U4249 (N_4249,N_3826,N_3631);
xnor U4250 (N_4250,N_3890,N_3084);
xnor U4251 (N_4251,N_3208,N_3507);
nand U4252 (N_4252,N_3775,N_3867);
nand U4253 (N_4253,N_3954,N_3318);
xor U4254 (N_4254,N_3994,N_3159);
and U4255 (N_4255,N_3321,N_3808);
xor U4256 (N_4256,N_3438,N_3119);
and U4257 (N_4257,N_3700,N_3363);
and U4258 (N_4258,N_3580,N_3779);
xor U4259 (N_4259,N_3630,N_3711);
and U4260 (N_4260,N_3404,N_3851);
nor U4261 (N_4261,N_3529,N_3334);
or U4262 (N_4262,N_3710,N_3995);
or U4263 (N_4263,N_3156,N_3149);
or U4264 (N_4264,N_3566,N_3695);
or U4265 (N_4265,N_3062,N_3102);
nor U4266 (N_4266,N_3282,N_3615);
nor U4267 (N_4267,N_3792,N_3370);
nand U4268 (N_4268,N_3536,N_3991);
xor U4269 (N_4269,N_3033,N_3525);
xnor U4270 (N_4270,N_3445,N_3844);
nand U4271 (N_4271,N_3480,N_3888);
or U4272 (N_4272,N_3479,N_3312);
nand U4273 (N_4273,N_3213,N_3916);
xor U4274 (N_4274,N_3250,N_3082);
nor U4275 (N_4275,N_3787,N_3770);
or U4276 (N_4276,N_3427,N_3300);
xnor U4277 (N_4277,N_3598,N_3223);
nor U4278 (N_4278,N_3767,N_3945);
nor U4279 (N_4279,N_3571,N_3103);
nor U4280 (N_4280,N_3639,N_3391);
nand U4281 (N_4281,N_3955,N_3457);
nand U4282 (N_4282,N_3130,N_3366);
nand U4283 (N_4283,N_3436,N_3632);
nor U4284 (N_4284,N_3414,N_3510);
and U4285 (N_4285,N_3532,N_3923);
and U4286 (N_4286,N_3949,N_3885);
or U4287 (N_4287,N_3843,N_3987);
xnor U4288 (N_4288,N_3676,N_3314);
nand U4289 (N_4289,N_3742,N_3714);
xor U4290 (N_4290,N_3182,N_3921);
or U4291 (N_4291,N_3483,N_3233);
and U4292 (N_4292,N_3705,N_3863);
and U4293 (N_4293,N_3245,N_3807);
nand U4294 (N_4294,N_3265,N_3398);
and U4295 (N_4295,N_3591,N_3408);
and U4296 (N_4296,N_3882,N_3841);
nand U4297 (N_4297,N_3419,N_3570);
xnor U4298 (N_4298,N_3622,N_3703);
or U4299 (N_4299,N_3367,N_3656);
xnor U4300 (N_4300,N_3906,N_3610);
or U4301 (N_4301,N_3986,N_3183);
xor U4302 (N_4302,N_3846,N_3261);
nor U4303 (N_4303,N_3296,N_3977);
nor U4304 (N_4304,N_3730,N_3231);
xor U4305 (N_4305,N_3298,N_3812);
nand U4306 (N_4306,N_3635,N_3693);
nor U4307 (N_4307,N_3806,N_3978);
or U4308 (N_4308,N_3146,N_3409);
xor U4309 (N_4309,N_3168,N_3828);
or U4310 (N_4310,N_3249,N_3399);
nand U4311 (N_4311,N_3346,N_3871);
nor U4312 (N_4312,N_3764,N_3735);
nor U4313 (N_4313,N_3669,N_3065);
nand U4314 (N_4314,N_3829,N_3262);
or U4315 (N_4315,N_3539,N_3107);
and U4316 (N_4316,N_3862,N_3848);
and U4317 (N_4317,N_3534,N_3243);
or U4318 (N_4318,N_3919,N_3431);
xor U4319 (N_4319,N_3905,N_3174);
nand U4320 (N_4320,N_3606,N_3044);
and U4321 (N_4321,N_3076,N_3831);
xnor U4322 (N_4322,N_3281,N_3613);
nor U4323 (N_4323,N_3175,N_3016);
nand U4324 (N_4324,N_3456,N_3659);
or U4325 (N_4325,N_3205,N_3052);
and U4326 (N_4326,N_3229,N_3010);
xnor U4327 (N_4327,N_3259,N_3795);
nand U4328 (N_4328,N_3278,N_3976);
nand U4329 (N_4329,N_3662,N_3047);
xor U4330 (N_4330,N_3061,N_3981);
nand U4331 (N_4331,N_3219,N_3743);
nor U4332 (N_4332,N_3541,N_3194);
xor U4333 (N_4333,N_3798,N_3228);
xnor U4334 (N_4334,N_3781,N_3216);
xor U4335 (N_4335,N_3755,N_3491);
and U4336 (N_4336,N_3465,N_3599);
xnor U4337 (N_4337,N_3190,N_3433);
and U4338 (N_4338,N_3025,N_3515);
or U4339 (N_4339,N_3579,N_3887);
nor U4340 (N_4340,N_3731,N_3236);
or U4341 (N_4341,N_3090,N_3940);
and U4342 (N_4342,N_3736,N_3429);
xnor U4343 (N_4343,N_3081,N_3449);
xor U4344 (N_4344,N_3821,N_3390);
nand U4345 (N_4345,N_3636,N_3239);
xor U4346 (N_4346,N_3886,N_3702);
and U4347 (N_4347,N_3717,N_3275);
and U4348 (N_4348,N_3270,N_3988);
and U4349 (N_4349,N_3932,N_3022);
nor U4350 (N_4350,N_3389,N_3193);
nor U4351 (N_4351,N_3160,N_3651);
nand U4352 (N_4352,N_3242,N_3474);
nand U4353 (N_4353,N_3345,N_3131);
nor U4354 (N_4354,N_3151,N_3192);
nor U4355 (N_4355,N_3028,N_3473);
xnor U4356 (N_4356,N_3706,N_3364);
and U4357 (N_4357,N_3244,N_3960);
nand U4358 (N_4358,N_3041,N_3834);
or U4359 (N_4359,N_3996,N_3068);
xnor U4360 (N_4360,N_3405,N_3472);
nand U4361 (N_4361,N_3734,N_3029);
xor U4362 (N_4362,N_3137,N_3011);
xor U4363 (N_4363,N_3158,N_3336);
or U4364 (N_4364,N_3169,N_3049);
nor U4365 (N_4365,N_3343,N_3360);
xor U4366 (N_4366,N_3683,N_3998);
and U4367 (N_4367,N_3255,N_3352);
or U4368 (N_4368,N_3620,N_3540);
and U4369 (N_4369,N_3444,N_3509);
and U4370 (N_4370,N_3291,N_3634);
xnor U4371 (N_4371,N_3354,N_3883);
nor U4372 (N_4372,N_3657,N_3424);
nor U4373 (N_4373,N_3943,N_3121);
and U4374 (N_4374,N_3928,N_3214);
or U4375 (N_4375,N_3892,N_3458);
nor U4376 (N_4376,N_3809,N_3820);
or U4377 (N_4377,N_3075,N_3323);
and U4378 (N_4378,N_3272,N_3447);
and U4379 (N_4379,N_3184,N_3686);
nor U4380 (N_4380,N_3177,N_3066);
xor U4381 (N_4381,N_3333,N_3074);
and U4382 (N_4382,N_3827,N_3810);
nand U4383 (N_4383,N_3640,N_3633);
nand U4384 (N_4384,N_3530,N_3463);
nand U4385 (N_4385,N_3150,N_3984);
nor U4386 (N_4386,N_3340,N_3129);
nand U4387 (N_4387,N_3898,N_3854);
nand U4388 (N_4388,N_3900,N_3759);
or U4389 (N_4389,N_3668,N_3805);
nor U4390 (N_4390,N_3677,N_3096);
xnor U4391 (N_4391,N_3802,N_3596);
nand U4392 (N_4392,N_3276,N_3015);
xor U4393 (N_4393,N_3179,N_3535);
xor U4394 (N_4394,N_3024,N_3064);
or U4395 (N_4395,N_3753,N_3063);
nor U4396 (N_4396,N_3154,N_3050);
xnor U4397 (N_4397,N_3602,N_3990);
xnor U4398 (N_4398,N_3048,N_3315);
nor U4399 (N_4399,N_3788,N_3325);
nor U4400 (N_4400,N_3681,N_3918);
or U4401 (N_4401,N_3609,N_3099);
and U4402 (N_4402,N_3269,N_3563);
nand U4403 (N_4403,N_3215,N_3109);
nor U4404 (N_4404,N_3773,N_3878);
xnor U4405 (N_4405,N_3410,N_3356);
or U4406 (N_4406,N_3067,N_3478);
xnor U4407 (N_4407,N_3388,N_3020);
and U4408 (N_4408,N_3520,N_3342);
and U4409 (N_4409,N_3279,N_3266);
nand U4410 (N_4410,N_3627,N_3338);
nor U4411 (N_4411,N_3057,N_3849);
nor U4412 (N_4412,N_3797,N_3416);
and U4413 (N_4413,N_3207,N_3091);
nand U4414 (N_4414,N_3757,N_3351);
and U4415 (N_4415,N_3147,N_3897);
nand U4416 (N_4416,N_3974,N_3106);
nand U4417 (N_4417,N_3488,N_3461);
xnor U4418 (N_4418,N_3889,N_3750);
nor U4419 (N_4419,N_3462,N_3518);
and U4420 (N_4420,N_3499,N_3903);
or U4421 (N_4421,N_3027,N_3386);
and U4422 (N_4422,N_3909,N_3437);
nand U4423 (N_4423,N_3603,N_3856);
nor U4424 (N_4424,N_3126,N_3138);
nand U4425 (N_4425,N_3002,N_3349);
xor U4426 (N_4426,N_3782,N_3212);
and U4427 (N_4427,N_3042,N_3574);
or U4428 (N_4428,N_3232,N_3604);
nor U4429 (N_4429,N_3375,N_3403);
or U4430 (N_4430,N_3094,N_3969);
and U4431 (N_4431,N_3251,N_3420);
xnor U4432 (N_4432,N_3586,N_3017);
nand U4433 (N_4433,N_3371,N_3801);
and U4434 (N_4434,N_3393,N_3070);
or U4435 (N_4435,N_3302,N_3293);
or U4436 (N_4436,N_3980,N_3256);
and U4437 (N_4437,N_3680,N_3197);
and U4438 (N_4438,N_3587,N_3697);
nor U4439 (N_4439,N_3292,N_3876);
nand U4440 (N_4440,N_3751,N_3059);
nand U4441 (N_4441,N_3749,N_3643);
nor U4442 (N_4442,N_3104,N_3776);
or U4443 (N_4443,N_3034,N_3139);
and U4444 (N_4444,N_3583,N_3907);
or U4445 (N_4445,N_3513,N_3616);
xor U4446 (N_4446,N_3664,N_3551);
nor U4447 (N_4447,N_3317,N_3629);
and U4448 (N_4448,N_3361,N_3127);
and U4449 (N_4449,N_3327,N_3522);
and U4450 (N_4450,N_3908,N_3607);
nor U4451 (N_4451,N_3521,N_3952);
nor U4452 (N_4452,N_3670,N_3500);
and U4453 (N_4453,N_3164,N_3555);
or U4454 (N_4454,N_3936,N_3003);
xnor U4455 (N_4455,N_3252,N_3858);
nand U4456 (N_4456,N_3771,N_3374);
and U4457 (N_4457,N_3559,N_3058);
nand U4458 (N_4458,N_3692,N_3289);
and U4459 (N_4459,N_3967,N_3365);
xor U4460 (N_4460,N_3533,N_3425);
xor U4461 (N_4461,N_3922,N_3372);
and U4462 (N_4462,N_3335,N_3655);
xor U4463 (N_4463,N_3979,N_3180);
and U4464 (N_4464,N_3992,N_3348);
nand U4465 (N_4465,N_3712,N_3811);
nor U4466 (N_4466,N_3589,N_3993);
nand U4467 (N_4467,N_3110,N_3468);
nor U4468 (N_4468,N_3623,N_3198);
xor U4469 (N_4469,N_3195,N_3595);
and U4470 (N_4470,N_3605,N_3601);
nor U4471 (N_4471,N_3724,N_3324);
nor U4472 (N_4472,N_3378,N_3719);
nor U4473 (N_4473,N_3685,N_3263);
xnor U4474 (N_4474,N_3019,N_3053);
or U4475 (N_4475,N_3173,N_3592);
xnor U4476 (N_4476,N_3665,N_3516);
xor U4477 (N_4477,N_3549,N_3124);
or U4478 (N_4478,N_3186,N_3572);
nor U4479 (N_4479,N_3253,N_3642);
nand U4480 (N_4480,N_3707,N_3663);
nand U4481 (N_4481,N_3359,N_3975);
nand U4482 (N_4482,N_3543,N_3380);
nand U4483 (N_4483,N_3460,N_3983);
xor U4484 (N_4484,N_3968,N_3678);
and U4485 (N_4485,N_3441,N_3337);
xnor U4486 (N_4486,N_3542,N_3774);
or U4487 (N_4487,N_3506,N_3038);
nor U4488 (N_4488,N_3284,N_3517);
and U4489 (N_4489,N_3777,N_3181);
nor U4490 (N_4490,N_3728,N_3238);
xor U4491 (N_4491,N_3715,N_3569);
or U4492 (N_4492,N_3114,N_3477);
nor U4493 (N_4493,N_3396,N_3939);
nor U4494 (N_4494,N_3562,N_3824);
nor U4495 (N_4495,N_3819,N_3171);
nand U4496 (N_4496,N_3417,N_3709);
nor U4497 (N_4497,N_3442,N_3914);
nand U4498 (N_4498,N_3224,N_3008);
nor U4499 (N_4499,N_3780,N_3073);
and U4500 (N_4500,N_3279,N_3517);
and U4501 (N_4501,N_3657,N_3593);
or U4502 (N_4502,N_3249,N_3972);
and U4503 (N_4503,N_3929,N_3688);
and U4504 (N_4504,N_3957,N_3248);
nand U4505 (N_4505,N_3223,N_3607);
xnor U4506 (N_4506,N_3968,N_3401);
or U4507 (N_4507,N_3442,N_3260);
nand U4508 (N_4508,N_3330,N_3356);
nor U4509 (N_4509,N_3640,N_3847);
xnor U4510 (N_4510,N_3022,N_3354);
nand U4511 (N_4511,N_3094,N_3983);
or U4512 (N_4512,N_3714,N_3450);
or U4513 (N_4513,N_3227,N_3920);
or U4514 (N_4514,N_3799,N_3328);
xor U4515 (N_4515,N_3104,N_3199);
xor U4516 (N_4516,N_3897,N_3888);
and U4517 (N_4517,N_3823,N_3691);
xnor U4518 (N_4518,N_3296,N_3506);
or U4519 (N_4519,N_3475,N_3076);
nand U4520 (N_4520,N_3005,N_3070);
or U4521 (N_4521,N_3817,N_3004);
nor U4522 (N_4522,N_3059,N_3600);
or U4523 (N_4523,N_3379,N_3999);
xnor U4524 (N_4524,N_3429,N_3767);
and U4525 (N_4525,N_3504,N_3618);
nor U4526 (N_4526,N_3732,N_3287);
xnor U4527 (N_4527,N_3153,N_3296);
nor U4528 (N_4528,N_3665,N_3176);
xnor U4529 (N_4529,N_3469,N_3743);
and U4530 (N_4530,N_3965,N_3484);
xnor U4531 (N_4531,N_3931,N_3298);
nor U4532 (N_4532,N_3591,N_3734);
and U4533 (N_4533,N_3545,N_3349);
xor U4534 (N_4534,N_3280,N_3340);
nand U4535 (N_4535,N_3812,N_3459);
nand U4536 (N_4536,N_3805,N_3518);
nor U4537 (N_4537,N_3239,N_3363);
nor U4538 (N_4538,N_3666,N_3895);
or U4539 (N_4539,N_3076,N_3910);
and U4540 (N_4540,N_3032,N_3772);
or U4541 (N_4541,N_3918,N_3202);
and U4542 (N_4542,N_3061,N_3899);
nor U4543 (N_4543,N_3110,N_3972);
xnor U4544 (N_4544,N_3128,N_3778);
xnor U4545 (N_4545,N_3403,N_3840);
and U4546 (N_4546,N_3957,N_3646);
xor U4547 (N_4547,N_3808,N_3334);
nor U4548 (N_4548,N_3454,N_3489);
nor U4549 (N_4549,N_3806,N_3261);
or U4550 (N_4550,N_3797,N_3913);
and U4551 (N_4551,N_3356,N_3048);
and U4552 (N_4552,N_3062,N_3922);
xor U4553 (N_4553,N_3615,N_3511);
nor U4554 (N_4554,N_3312,N_3973);
xor U4555 (N_4555,N_3260,N_3044);
or U4556 (N_4556,N_3844,N_3593);
xor U4557 (N_4557,N_3672,N_3219);
or U4558 (N_4558,N_3073,N_3539);
and U4559 (N_4559,N_3035,N_3440);
and U4560 (N_4560,N_3063,N_3668);
nand U4561 (N_4561,N_3703,N_3756);
and U4562 (N_4562,N_3468,N_3474);
or U4563 (N_4563,N_3353,N_3519);
nand U4564 (N_4564,N_3077,N_3068);
and U4565 (N_4565,N_3429,N_3060);
and U4566 (N_4566,N_3041,N_3039);
xnor U4567 (N_4567,N_3343,N_3080);
or U4568 (N_4568,N_3875,N_3496);
or U4569 (N_4569,N_3942,N_3663);
xnor U4570 (N_4570,N_3351,N_3245);
nand U4571 (N_4571,N_3574,N_3066);
nand U4572 (N_4572,N_3513,N_3735);
xor U4573 (N_4573,N_3335,N_3165);
nand U4574 (N_4574,N_3736,N_3968);
xor U4575 (N_4575,N_3651,N_3181);
and U4576 (N_4576,N_3530,N_3580);
or U4577 (N_4577,N_3431,N_3502);
or U4578 (N_4578,N_3535,N_3233);
and U4579 (N_4579,N_3901,N_3416);
or U4580 (N_4580,N_3006,N_3787);
or U4581 (N_4581,N_3980,N_3116);
nor U4582 (N_4582,N_3115,N_3493);
or U4583 (N_4583,N_3641,N_3308);
and U4584 (N_4584,N_3085,N_3161);
nor U4585 (N_4585,N_3567,N_3494);
and U4586 (N_4586,N_3496,N_3593);
and U4587 (N_4587,N_3386,N_3907);
xnor U4588 (N_4588,N_3310,N_3315);
and U4589 (N_4589,N_3556,N_3223);
and U4590 (N_4590,N_3449,N_3007);
nor U4591 (N_4591,N_3726,N_3481);
and U4592 (N_4592,N_3120,N_3677);
xnor U4593 (N_4593,N_3386,N_3299);
and U4594 (N_4594,N_3917,N_3829);
xnor U4595 (N_4595,N_3926,N_3802);
xnor U4596 (N_4596,N_3953,N_3232);
nand U4597 (N_4597,N_3682,N_3345);
or U4598 (N_4598,N_3109,N_3602);
xor U4599 (N_4599,N_3578,N_3300);
nor U4600 (N_4600,N_3817,N_3147);
nor U4601 (N_4601,N_3324,N_3881);
and U4602 (N_4602,N_3221,N_3107);
nand U4603 (N_4603,N_3196,N_3214);
and U4604 (N_4604,N_3806,N_3033);
nor U4605 (N_4605,N_3201,N_3317);
nand U4606 (N_4606,N_3816,N_3628);
nor U4607 (N_4607,N_3392,N_3139);
nor U4608 (N_4608,N_3973,N_3893);
xnor U4609 (N_4609,N_3405,N_3387);
nand U4610 (N_4610,N_3921,N_3685);
xor U4611 (N_4611,N_3026,N_3233);
nor U4612 (N_4612,N_3789,N_3912);
and U4613 (N_4613,N_3814,N_3103);
nor U4614 (N_4614,N_3116,N_3093);
nand U4615 (N_4615,N_3608,N_3718);
or U4616 (N_4616,N_3021,N_3483);
xor U4617 (N_4617,N_3353,N_3913);
xnor U4618 (N_4618,N_3442,N_3194);
or U4619 (N_4619,N_3942,N_3941);
and U4620 (N_4620,N_3162,N_3842);
nor U4621 (N_4621,N_3055,N_3289);
or U4622 (N_4622,N_3201,N_3388);
nor U4623 (N_4623,N_3527,N_3436);
and U4624 (N_4624,N_3819,N_3324);
nor U4625 (N_4625,N_3302,N_3193);
xnor U4626 (N_4626,N_3734,N_3494);
nor U4627 (N_4627,N_3739,N_3922);
and U4628 (N_4628,N_3016,N_3322);
nor U4629 (N_4629,N_3112,N_3059);
nand U4630 (N_4630,N_3832,N_3593);
or U4631 (N_4631,N_3048,N_3982);
nor U4632 (N_4632,N_3730,N_3296);
nor U4633 (N_4633,N_3740,N_3178);
xor U4634 (N_4634,N_3264,N_3948);
nor U4635 (N_4635,N_3448,N_3582);
or U4636 (N_4636,N_3643,N_3434);
nor U4637 (N_4637,N_3196,N_3282);
xor U4638 (N_4638,N_3049,N_3358);
nor U4639 (N_4639,N_3087,N_3468);
nand U4640 (N_4640,N_3823,N_3009);
nand U4641 (N_4641,N_3957,N_3876);
and U4642 (N_4642,N_3918,N_3052);
xnor U4643 (N_4643,N_3662,N_3138);
and U4644 (N_4644,N_3753,N_3621);
and U4645 (N_4645,N_3892,N_3023);
and U4646 (N_4646,N_3333,N_3583);
or U4647 (N_4647,N_3298,N_3027);
nand U4648 (N_4648,N_3817,N_3054);
nand U4649 (N_4649,N_3362,N_3929);
xnor U4650 (N_4650,N_3908,N_3989);
nand U4651 (N_4651,N_3826,N_3767);
xnor U4652 (N_4652,N_3201,N_3762);
and U4653 (N_4653,N_3517,N_3095);
xnor U4654 (N_4654,N_3148,N_3574);
and U4655 (N_4655,N_3469,N_3937);
and U4656 (N_4656,N_3798,N_3058);
xor U4657 (N_4657,N_3669,N_3106);
and U4658 (N_4658,N_3370,N_3384);
and U4659 (N_4659,N_3610,N_3526);
nand U4660 (N_4660,N_3011,N_3047);
or U4661 (N_4661,N_3204,N_3180);
or U4662 (N_4662,N_3192,N_3921);
or U4663 (N_4663,N_3275,N_3017);
and U4664 (N_4664,N_3157,N_3010);
nand U4665 (N_4665,N_3224,N_3153);
nor U4666 (N_4666,N_3565,N_3319);
or U4667 (N_4667,N_3154,N_3699);
or U4668 (N_4668,N_3395,N_3344);
nand U4669 (N_4669,N_3476,N_3570);
nand U4670 (N_4670,N_3120,N_3854);
nor U4671 (N_4671,N_3347,N_3356);
nor U4672 (N_4672,N_3360,N_3724);
or U4673 (N_4673,N_3980,N_3437);
and U4674 (N_4674,N_3885,N_3753);
and U4675 (N_4675,N_3190,N_3010);
and U4676 (N_4676,N_3205,N_3838);
or U4677 (N_4677,N_3444,N_3004);
and U4678 (N_4678,N_3588,N_3406);
nand U4679 (N_4679,N_3393,N_3985);
and U4680 (N_4680,N_3514,N_3105);
xor U4681 (N_4681,N_3554,N_3204);
nand U4682 (N_4682,N_3635,N_3867);
xor U4683 (N_4683,N_3684,N_3974);
and U4684 (N_4684,N_3922,N_3908);
xnor U4685 (N_4685,N_3188,N_3485);
or U4686 (N_4686,N_3294,N_3755);
nand U4687 (N_4687,N_3444,N_3463);
or U4688 (N_4688,N_3049,N_3911);
nor U4689 (N_4689,N_3289,N_3837);
nor U4690 (N_4690,N_3480,N_3329);
xor U4691 (N_4691,N_3473,N_3248);
and U4692 (N_4692,N_3484,N_3162);
xor U4693 (N_4693,N_3345,N_3116);
xor U4694 (N_4694,N_3102,N_3949);
nand U4695 (N_4695,N_3565,N_3409);
and U4696 (N_4696,N_3897,N_3768);
and U4697 (N_4697,N_3126,N_3958);
nand U4698 (N_4698,N_3596,N_3455);
and U4699 (N_4699,N_3678,N_3920);
nor U4700 (N_4700,N_3954,N_3005);
nand U4701 (N_4701,N_3157,N_3606);
and U4702 (N_4702,N_3217,N_3370);
or U4703 (N_4703,N_3684,N_3962);
nor U4704 (N_4704,N_3183,N_3304);
nand U4705 (N_4705,N_3862,N_3214);
xnor U4706 (N_4706,N_3955,N_3540);
xnor U4707 (N_4707,N_3875,N_3736);
nor U4708 (N_4708,N_3671,N_3472);
and U4709 (N_4709,N_3613,N_3483);
nor U4710 (N_4710,N_3545,N_3216);
nor U4711 (N_4711,N_3660,N_3103);
nor U4712 (N_4712,N_3830,N_3462);
nand U4713 (N_4713,N_3744,N_3484);
xor U4714 (N_4714,N_3752,N_3391);
or U4715 (N_4715,N_3413,N_3396);
nand U4716 (N_4716,N_3726,N_3045);
nor U4717 (N_4717,N_3241,N_3269);
and U4718 (N_4718,N_3727,N_3677);
or U4719 (N_4719,N_3184,N_3252);
and U4720 (N_4720,N_3303,N_3669);
nor U4721 (N_4721,N_3353,N_3576);
nand U4722 (N_4722,N_3760,N_3611);
nor U4723 (N_4723,N_3224,N_3745);
and U4724 (N_4724,N_3233,N_3041);
and U4725 (N_4725,N_3180,N_3274);
and U4726 (N_4726,N_3418,N_3092);
and U4727 (N_4727,N_3131,N_3224);
and U4728 (N_4728,N_3448,N_3234);
nand U4729 (N_4729,N_3547,N_3198);
xor U4730 (N_4730,N_3118,N_3559);
nand U4731 (N_4731,N_3399,N_3380);
nand U4732 (N_4732,N_3087,N_3139);
nor U4733 (N_4733,N_3310,N_3416);
and U4734 (N_4734,N_3655,N_3639);
or U4735 (N_4735,N_3495,N_3765);
nand U4736 (N_4736,N_3575,N_3735);
nand U4737 (N_4737,N_3196,N_3394);
nand U4738 (N_4738,N_3845,N_3976);
and U4739 (N_4739,N_3462,N_3051);
nand U4740 (N_4740,N_3870,N_3214);
xnor U4741 (N_4741,N_3960,N_3393);
or U4742 (N_4742,N_3034,N_3064);
or U4743 (N_4743,N_3820,N_3559);
xor U4744 (N_4744,N_3843,N_3032);
nand U4745 (N_4745,N_3896,N_3077);
or U4746 (N_4746,N_3242,N_3445);
or U4747 (N_4747,N_3062,N_3868);
xnor U4748 (N_4748,N_3049,N_3241);
or U4749 (N_4749,N_3786,N_3226);
xor U4750 (N_4750,N_3206,N_3481);
or U4751 (N_4751,N_3536,N_3866);
xor U4752 (N_4752,N_3485,N_3561);
nor U4753 (N_4753,N_3423,N_3083);
nor U4754 (N_4754,N_3815,N_3145);
and U4755 (N_4755,N_3220,N_3522);
and U4756 (N_4756,N_3519,N_3037);
or U4757 (N_4757,N_3439,N_3713);
or U4758 (N_4758,N_3866,N_3928);
nand U4759 (N_4759,N_3503,N_3119);
nand U4760 (N_4760,N_3979,N_3114);
nor U4761 (N_4761,N_3883,N_3954);
and U4762 (N_4762,N_3963,N_3762);
or U4763 (N_4763,N_3840,N_3067);
and U4764 (N_4764,N_3807,N_3131);
nor U4765 (N_4765,N_3034,N_3897);
and U4766 (N_4766,N_3131,N_3611);
or U4767 (N_4767,N_3884,N_3561);
nor U4768 (N_4768,N_3955,N_3748);
nand U4769 (N_4769,N_3420,N_3582);
or U4770 (N_4770,N_3681,N_3137);
xnor U4771 (N_4771,N_3303,N_3446);
or U4772 (N_4772,N_3695,N_3625);
nand U4773 (N_4773,N_3795,N_3419);
and U4774 (N_4774,N_3416,N_3969);
nand U4775 (N_4775,N_3177,N_3473);
xnor U4776 (N_4776,N_3717,N_3103);
nor U4777 (N_4777,N_3665,N_3715);
xor U4778 (N_4778,N_3230,N_3371);
and U4779 (N_4779,N_3791,N_3700);
or U4780 (N_4780,N_3085,N_3784);
or U4781 (N_4781,N_3785,N_3965);
or U4782 (N_4782,N_3077,N_3323);
xnor U4783 (N_4783,N_3574,N_3573);
xnor U4784 (N_4784,N_3437,N_3228);
nor U4785 (N_4785,N_3363,N_3137);
or U4786 (N_4786,N_3393,N_3217);
or U4787 (N_4787,N_3057,N_3783);
or U4788 (N_4788,N_3086,N_3152);
xnor U4789 (N_4789,N_3603,N_3389);
or U4790 (N_4790,N_3427,N_3890);
or U4791 (N_4791,N_3528,N_3549);
and U4792 (N_4792,N_3674,N_3042);
and U4793 (N_4793,N_3584,N_3607);
nor U4794 (N_4794,N_3744,N_3062);
nand U4795 (N_4795,N_3531,N_3018);
xor U4796 (N_4796,N_3362,N_3239);
and U4797 (N_4797,N_3251,N_3567);
xnor U4798 (N_4798,N_3482,N_3460);
nand U4799 (N_4799,N_3997,N_3229);
and U4800 (N_4800,N_3440,N_3501);
or U4801 (N_4801,N_3800,N_3969);
or U4802 (N_4802,N_3141,N_3787);
or U4803 (N_4803,N_3617,N_3734);
xnor U4804 (N_4804,N_3372,N_3172);
nor U4805 (N_4805,N_3202,N_3257);
nand U4806 (N_4806,N_3382,N_3681);
xnor U4807 (N_4807,N_3061,N_3708);
and U4808 (N_4808,N_3727,N_3419);
and U4809 (N_4809,N_3720,N_3399);
and U4810 (N_4810,N_3241,N_3299);
xor U4811 (N_4811,N_3918,N_3587);
nor U4812 (N_4812,N_3037,N_3135);
nand U4813 (N_4813,N_3784,N_3259);
nand U4814 (N_4814,N_3569,N_3255);
nand U4815 (N_4815,N_3016,N_3149);
or U4816 (N_4816,N_3909,N_3386);
xor U4817 (N_4817,N_3006,N_3478);
or U4818 (N_4818,N_3794,N_3928);
or U4819 (N_4819,N_3712,N_3007);
nand U4820 (N_4820,N_3961,N_3757);
or U4821 (N_4821,N_3802,N_3008);
xor U4822 (N_4822,N_3478,N_3245);
nor U4823 (N_4823,N_3190,N_3495);
xnor U4824 (N_4824,N_3604,N_3250);
nand U4825 (N_4825,N_3660,N_3381);
nand U4826 (N_4826,N_3054,N_3824);
nand U4827 (N_4827,N_3202,N_3271);
xnor U4828 (N_4828,N_3211,N_3377);
xnor U4829 (N_4829,N_3477,N_3145);
xnor U4830 (N_4830,N_3116,N_3667);
or U4831 (N_4831,N_3707,N_3024);
nand U4832 (N_4832,N_3701,N_3770);
and U4833 (N_4833,N_3169,N_3851);
or U4834 (N_4834,N_3296,N_3774);
xor U4835 (N_4835,N_3527,N_3244);
and U4836 (N_4836,N_3339,N_3074);
and U4837 (N_4837,N_3542,N_3464);
nor U4838 (N_4838,N_3638,N_3205);
nand U4839 (N_4839,N_3619,N_3390);
and U4840 (N_4840,N_3748,N_3102);
xor U4841 (N_4841,N_3617,N_3482);
xor U4842 (N_4842,N_3350,N_3704);
and U4843 (N_4843,N_3428,N_3033);
or U4844 (N_4844,N_3971,N_3594);
nor U4845 (N_4845,N_3388,N_3255);
or U4846 (N_4846,N_3864,N_3383);
nand U4847 (N_4847,N_3283,N_3648);
or U4848 (N_4848,N_3926,N_3405);
xor U4849 (N_4849,N_3918,N_3623);
nor U4850 (N_4850,N_3780,N_3514);
nand U4851 (N_4851,N_3975,N_3093);
and U4852 (N_4852,N_3235,N_3909);
and U4853 (N_4853,N_3747,N_3423);
xor U4854 (N_4854,N_3304,N_3466);
and U4855 (N_4855,N_3049,N_3144);
or U4856 (N_4856,N_3771,N_3536);
nor U4857 (N_4857,N_3322,N_3284);
or U4858 (N_4858,N_3280,N_3727);
or U4859 (N_4859,N_3288,N_3438);
and U4860 (N_4860,N_3873,N_3515);
xor U4861 (N_4861,N_3916,N_3379);
or U4862 (N_4862,N_3529,N_3054);
nand U4863 (N_4863,N_3542,N_3496);
nand U4864 (N_4864,N_3804,N_3092);
or U4865 (N_4865,N_3447,N_3019);
and U4866 (N_4866,N_3635,N_3568);
nor U4867 (N_4867,N_3191,N_3474);
nor U4868 (N_4868,N_3558,N_3430);
and U4869 (N_4869,N_3016,N_3853);
and U4870 (N_4870,N_3841,N_3857);
nand U4871 (N_4871,N_3975,N_3278);
and U4872 (N_4872,N_3000,N_3096);
xor U4873 (N_4873,N_3506,N_3199);
nand U4874 (N_4874,N_3936,N_3729);
or U4875 (N_4875,N_3288,N_3855);
and U4876 (N_4876,N_3217,N_3580);
or U4877 (N_4877,N_3339,N_3231);
xnor U4878 (N_4878,N_3244,N_3582);
nor U4879 (N_4879,N_3084,N_3681);
nor U4880 (N_4880,N_3729,N_3506);
and U4881 (N_4881,N_3316,N_3125);
nor U4882 (N_4882,N_3246,N_3043);
nand U4883 (N_4883,N_3994,N_3255);
xnor U4884 (N_4884,N_3326,N_3287);
nor U4885 (N_4885,N_3651,N_3970);
and U4886 (N_4886,N_3417,N_3461);
nor U4887 (N_4887,N_3465,N_3316);
xnor U4888 (N_4888,N_3528,N_3648);
nor U4889 (N_4889,N_3022,N_3052);
or U4890 (N_4890,N_3452,N_3148);
or U4891 (N_4891,N_3341,N_3725);
nor U4892 (N_4892,N_3822,N_3933);
xnor U4893 (N_4893,N_3168,N_3583);
nand U4894 (N_4894,N_3693,N_3305);
nor U4895 (N_4895,N_3868,N_3506);
and U4896 (N_4896,N_3701,N_3357);
nand U4897 (N_4897,N_3939,N_3808);
or U4898 (N_4898,N_3155,N_3948);
nor U4899 (N_4899,N_3964,N_3246);
xnor U4900 (N_4900,N_3088,N_3785);
and U4901 (N_4901,N_3027,N_3882);
and U4902 (N_4902,N_3772,N_3128);
and U4903 (N_4903,N_3012,N_3577);
xnor U4904 (N_4904,N_3076,N_3300);
and U4905 (N_4905,N_3623,N_3805);
nor U4906 (N_4906,N_3369,N_3820);
xor U4907 (N_4907,N_3311,N_3781);
xnor U4908 (N_4908,N_3766,N_3948);
nand U4909 (N_4909,N_3475,N_3388);
or U4910 (N_4910,N_3245,N_3773);
xnor U4911 (N_4911,N_3289,N_3661);
nand U4912 (N_4912,N_3967,N_3526);
nor U4913 (N_4913,N_3798,N_3743);
nor U4914 (N_4914,N_3573,N_3570);
nand U4915 (N_4915,N_3991,N_3668);
nand U4916 (N_4916,N_3252,N_3720);
and U4917 (N_4917,N_3938,N_3897);
nand U4918 (N_4918,N_3276,N_3214);
or U4919 (N_4919,N_3967,N_3107);
nand U4920 (N_4920,N_3021,N_3646);
or U4921 (N_4921,N_3991,N_3277);
or U4922 (N_4922,N_3942,N_3946);
and U4923 (N_4923,N_3469,N_3065);
nor U4924 (N_4924,N_3701,N_3030);
xnor U4925 (N_4925,N_3703,N_3172);
or U4926 (N_4926,N_3680,N_3014);
and U4927 (N_4927,N_3304,N_3097);
and U4928 (N_4928,N_3757,N_3967);
and U4929 (N_4929,N_3026,N_3235);
nand U4930 (N_4930,N_3951,N_3516);
or U4931 (N_4931,N_3822,N_3261);
nor U4932 (N_4932,N_3089,N_3447);
xnor U4933 (N_4933,N_3610,N_3563);
or U4934 (N_4934,N_3436,N_3663);
nand U4935 (N_4935,N_3828,N_3561);
nand U4936 (N_4936,N_3983,N_3511);
nor U4937 (N_4937,N_3196,N_3314);
nor U4938 (N_4938,N_3061,N_3041);
or U4939 (N_4939,N_3042,N_3024);
or U4940 (N_4940,N_3841,N_3244);
xor U4941 (N_4941,N_3014,N_3184);
and U4942 (N_4942,N_3321,N_3806);
nand U4943 (N_4943,N_3970,N_3542);
and U4944 (N_4944,N_3462,N_3491);
nor U4945 (N_4945,N_3706,N_3521);
or U4946 (N_4946,N_3505,N_3534);
or U4947 (N_4947,N_3626,N_3089);
nand U4948 (N_4948,N_3821,N_3347);
and U4949 (N_4949,N_3703,N_3046);
or U4950 (N_4950,N_3168,N_3851);
nor U4951 (N_4951,N_3773,N_3684);
nor U4952 (N_4952,N_3958,N_3890);
nor U4953 (N_4953,N_3282,N_3520);
xor U4954 (N_4954,N_3942,N_3502);
and U4955 (N_4955,N_3967,N_3190);
nor U4956 (N_4956,N_3819,N_3094);
nand U4957 (N_4957,N_3362,N_3265);
xor U4958 (N_4958,N_3979,N_3157);
nor U4959 (N_4959,N_3178,N_3209);
xor U4960 (N_4960,N_3783,N_3566);
nor U4961 (N_4961,N_3798,N_3183);
or U4962 (N_4962,N_3790,N_3983);
and U4963 (N_4963,N_3701,N_3660);
and U4964 (N_4964,N_3456,N_3963);
or U4965 (N_4965,N_3966,N_3517);
nor U4966 (N_4966,N_3869,N_3711);
nand U4967 (N_4967,N_3810,N_3842);
nand U4968 (N_4968,N_3844,N_3272);
xor U4969 (N_4969,N_3899,N_3015);
nand U4970 (N_4970,N_3774,N_3775);
nor U4971 (N_4971,N_3747,N_3874);
xor U4972 (N_4972,N_3690,N_3777);
or U4973 (N_4973,N_3229,N_3838);
nand U4974 (N_4974,N_3072,N_3332);
nand U4975 (N_4975,N_3844,N_3954);
xnor U4976 (N_4976,N_3886,N_3068);
and U4977 (N_4977,N_3982,N_3700);
or U4978 (N_4978,N_3853,N_3382);
or U4979 (N_4979,N_3729,N_3986);
or U4980 (N_4980,N_3837,N_3788);
or U4981 (N_4981,N_3465,N_3625);
xor U4982 (N_4982,N_3779,N_3120);
nor U4983 (N_4983,N_3901,N_3013);
or U4984 (N_4984,N_3493,N_3300);
xor U4985 (N_4985,N_3509,N_3311);
nor U4986 (N_4986,N_3044,N_3693);
nor U4987 (N_4987,N_3662,N_3021);
or U4988 (N_4988,N_3776,N_3147);
and U4989 (N_4989,N_3835,N_3639);
and U4990 (N_4990,N_3118,N_3836);
nand U4991 (N_4991,N_3912,N_3034);
nand U4992 (N_4992,N_3529,N_3683);
and U4993 (N_4993,N_3750,N_3966);
nor U4994 (N_4994,N_3000,N_3301);
nand U4995 (N_4995,N_3517,N_3674);
or U4996 (N_4996,N_3791,N_3650);
or U4997 (N_4997,N_3704,N_3830);
xnor U4998 (N_4998,N_3608,N_3400);
xnor U4999 (N_4999,N_3862,N_3963);
nand U5000 (N_5000,N_4874,N_4408);
nand U5001 (N_5001,N_4306,N_4495);
and U5002 (N_5002,N_4721,N_4911);
or U5003 (N_5003,N_4844,N_4678);
xnor U5004 (N_5004,N_4694,N_4123);
nand U5005 (N_5005,N_4888,N_4599);
or U5006 (N_5006,N_4717,N_4532);
nand U5007 (N_5007,N_4352,N_4177);
nor U5008 (N_5008,N_4974,N_4530);
and U5009 (N_5009,N_4116,N_4718);
or U5010 (N_5010,N_4422,N_4134);
nor U5011 (N_5011,N_4150,N_4025);
nor U5012 (N_5012,N_4401,N_4867);
nand U5013 (N_5013,N_4549,N_4443);
xor U5014 (N_5014,N_4729,N_4781);
and U5015 (N_5015,N_4388,N_4001);
nand U5016 (N_5016,N_4474,N_4148);
nand U5017 (N_5017,N_4560,N_4818);
or U5018 (N_5018,N_4297,N_4395);
xor U5019 (N_5019,N_4905,N_4108);
and U5020 (N_5020,N_4379,N_4660);
nor U5021 (N_5021,N_4128,N_4575);
or U5022 (N_5022,N_4344,N_4900);
xnor U5023 (N_5023,N_4237,N_4590);
or U5024 (N_5024,N_4954,N_4511);
and U5025 (N_5025,N_4287,N_4830);
and U5026 (N_5026,N_4021,N_4356);
nand U5027 (N_5027,N_4557,N_4853);
nor U5028 (N_5028,N_4630,N_4078);
nor U5029 (N_5029,N_4949,N_4990);
and U5030 (N_5030,N_4671,N_4995);
and U5031 (N_5031,N_4454,N_4597);
nor U5032 (N_5032,N_4200,N_4424);
and U5033 (N_5033,N_4561,N_4886);
and U5034 (N_5034,N_4458,N_4427);
xnor U5035 (N_5035,N_4983,N_4085);
nand U5036 (N_5036,N_4198,N_4171);
nor U5037 (N_5037,N_4228,N_4270);
and U5038 (N_5038,N_4663,N_4908);
xnor U5039 (N_5039,N_4375,N_4684);
and U5040 (N_5040,N_4258,N_4441);
nor U5041 (N_5041,N_4155,N_4508);
nand U5042 (N_5042,N_4505,N_4572);
xnor U5043 (N_5043,N_4756,N_4866);
nand U5044 (N_5044,N_4326,N_4223);
or U5045 (N_5045,N_4858,N_4095);
nand U5046 (N_5046,N_4758,N_4411);
nand U5047 (N_5047,N_4700,N_4725);
and U5048 (N_5048,N_4364,N_4435);
or U5049 (N_5049,N_4952,N_4096);
nand U5050 (N_5050,N_4368,N_4883);
nand U5051 (N_5051,N_4143,N_4436);
nor U5052 (N_5052,N_4604,N_4412);
and U5053 (N_5053,N_4677,N_4767);
and U5054 (N_5054,N_4061,N_4307);
and U5055 (N_5055,N_4340,N_4358);
nor U5056 (N_5056,N_4730,N_4803);
nor U5057 (N_5057,N_4950,N_4323);
xor U5058 (N_5058,N_4314,N_4088);
or U5059 (N_5059,N_4139,N_4529);
and U5060 (N_5060,N_4037,N_4890);
and U5061 (N_5061,N_4914,N_4073);
xnor U5062 (N_5062,N_4426,N_4175);
or U5063 (N_5063,N_4409,N_4159);
nand U5064 (N_5064,N_4434,N_4667);
and U5065 (N_5065,N_4615,N_4606);
nor U5066 (N_5066,N_4945,N_4417);
nand U5067 (N_5067,N_4760,N_4355);
and U5068 (N_5068,N_4673,N_4525);
or U5069 (N_5069,N_4894,N_4849);
nand U5070 (N_5070,N_4790,N_4745);
and U5071 (N_5071,N_4372,N_4608);
nand U5072 (N_5072,N_4014,N_4846);
nor U5073 (N_5073,N_4452,N_4126);
and U5074 (N_5074,N_4842,N_4241);
nor U5075 (N_5075,N_4902,N_4063);
nand U5076 (N_5076,N_4587,N_4211);
and U5077 (N_5077,N_4145,N_4603);
nand U5078 (N_5078,N_4054,N_4629);
nor U5079 (N_5079,N_4782,N_4056);
nor U5080 (N_5080,N_4804,N_4618);
or U5081 (N_5081,N_4705,N_4548);
or U5082 (N_5082,N_4301,N_4715);
nor U5083 (N_5083,N_4045,N_4311);
or U5084 (N_5084,N_4167,N_4492);
xor U5085 (N_5085,N_4584,N_4413);
nand U5086 (N_5086,N_4956,N_4191);
and U5087 (N_5087,N_4591,N_4464);
and U5088 (N_5088,N_4257,N_4278);
xor U5089 (N_5089,N_4656,N_4939);
nand U5090 (N_5090,N_4512,N_4583);
or U5091 (N_5091,N_4967,N_4860);
xnor U5092 (N_5092,N_4166,N_4058);
and U5093 (N_5093,N_4201,N_4196);
xor U5094 (N_5094,N_4710,N_4267);
or U5095 (N_5095,N_4308,N_4205);
nand U5096 (N_5096,N_4770,N_4496);
xor U5097 (N_5097,N_4773,N_4002);
xor U5098 (N_5098,N_4477,N_4927);
nor U5099 (N_5099,N_4796,N_4049);
or U5100 (N_5100,N_4137,N_4224);
or U5101 (N_5101,N_4194,N_4125);
nand U5102 (N_5102,N_4253,N_4944);
or U5103 (N_5103,N_4097,N_4076);
nor U5104 (N_5104,N_4910,N_4231);
xnor U5105 (N_5105,N_4000,N_4923);
or U5106 (N_5106,N_4199,N_4907);
xnor U5107 (N_5107,N_4038,N_4219);
nand U5108 (N_5108,N_4640,N_4397);
nand U5109 (N_5109,N_4517,N_4699);
nand U5110 (N_5110,N_4363,N_4493);
xnor U5111 (N_5111,N_4887,N_4015);
nand U5112 (N_5112,N_4197,N_4947);
or U5113 (N_5113,N_4222,N_4418);
xnor U5114 (N_5114,N_4631,N_4469);
xor U5115 (N_5115,N_4450,N_4940);
xor U5116 (N_5116,N_4659,N_4963);
xor U5117 (N_5117,N_4127,N_4130);
xnor U5118 (N_5118,N_4565,N_4616);
and U5119 (N_5119,N_4103,N_4720);
nand U5120 (N_5120,N_4010,N_4124);
and U5121 (N_5121,N_4724,N_4092);
or U5122 (N_5122,N_4792,N_4925);
or U5123 (N_5123,N_4385,N_4892);
nor U5124 (N_5124,N_4633,N_4786);
nor U5125 (N_5125,N_4672,N_4747);
nand U5126 (N_5126,N_4377,N_4460);
nor U5127 (N_5127,N_4602,N_4751);
and U5128 (N_5128,N_4999,N_4286);
xor U5129 (N_5129,N_4509,N_4765);
xor U5130 (N_5130,N_4321,N_4554);
and U5131 (N_5131,N_4279,N_4537);
and U5132 (N_5132,N_4920,N_4499);
and U5133 (N_5133,N_4689,N_4893);
nor U5134 (N_5134,N_4889,N_4997);
nor U5135 (N_5135,N_4034,N_4733);
or U5136 (N_5136,N_4333,N_4206);
xnor U5137 (N_5137,N_4918,N_4793);
or U5138 (N_5138,N_4467,N_4807);
nand U5139 (N_5139,N_4988,N_4826);
xnor U5140 (N_5140,N_4612,N_4484);
nor U5141 (N_5141,N_4319,N_4518);
and U5142 (N_5142,N_4627,N_4594);
xnor U5143 (N_5143,N_4275,N_4607);
nand U5144 (N_5144,N_4646,N_4144);
xor U5145 (N_5145,N_4107,N_4723);
nand U5146 (N_5146,N_4698,N_4029);
or U5147 (N_5147,N_4683,N_4870);
or U5148 (N_5148,N_4162,N_4055);
nor U5149 (N_5149,N_4421,N_4420);
and U5150 (N_5150,N_4558,N_4979);
xor U5151 (N_5151,N_4614,N_4759);
nor U5152 (N_5152,N_4272,N_4296);
and U5153 (N_5153,N_4843,N_4808);
nor U5154 (N_5154,N_4284,N_4059);
and U5155 (N_5155,N_4716,N_4057);
nor U5156 (N_5156,N_4106,N_4317);
nor U5157 (N_5157,N_4501,N_4789);
and U5158 (N_5158,N_4068,N_4819);
nor U5159 (N_5159,N_4871,N_4938);
nand U5160 (N_5160,N_4556,N_4466);
and U5161 (N_5161,N_4218,N_4252);
xor U5162 (N_5162,N_4519,N_4153);
nor U5163 (N_5163,N_4806,N_4504);
xor U5164 (N_5164,N_4534,N_4650);
nand U5165 (N_5165,N_4996,N_4390);
xor U5166 (N_5166,N_4544,N_4315);
nor U5167 (N_5167,N_4567,N_4090);
or U5168 (N_5168,N_4651,N_4188);
or U5169 (N_5169,N_4432,N_4714);
or U5170 (N_5170,N_4851,N_4405);
nand U5171 (N_5171,N_4625,N_4934);
nand U5172 (N_5172,N_4313,N_4236);
xnor U5173 (N_5173,N_4690,N_4041);
nand U5174 (N_5174,N_4547,N_4491);
nand U5175 (N_5175,N_4884,N_4482);
xnor U5176 (N_5176,N_4332,N_4552);
and U5177 (N_5177,N_4331,N_4098);
or U5178 (N_5178,N_4288,N_4930);
xor U5179 (N_5179,N_4329,N_4449);
xnor U5180 (N_5180,N_4341,N_4245);
xnor U5181 (N_5181,N_4227,N_4741);
and U5182 (N_5182,N_4687,N_4559);
nand U5183 (N_5183,N_4835,N_4220);
or U5184 (N_5184,N_4051,N_4915);
nand U5185 (N_5185,N_4551,N_4328);
nor U5186 (N_5186,N_4665,N_4030);
and U5187 (N_5187,N_4840,N_4813);
and U5188 (N_5188,N_4611,N_4610);
and U5189 (N_5189,N_4254,N_4283);
or U5190 (N_5190,N_4133,N_4815);
xnor U5191 (N_5191,N_4847,N_4681);
nor U5192 (N_5192,N_4935,N_4471);
xor U5193 (N_5193,N_4779,N_4896);
nand U5194 (N_5194,N_4783,N_4566);
and U5195 (N_5195,N_4772,N_4778);
and U5196 (N_5196,N_4291,N_4320);
nand U5197 (N_5197,N_4023,N_4429);
nand U5198 (N_5198,N_4456,N_4662);
xor U5199 (N_5199,N_4248,N_4764);
xor U5200 (N_5200,N_4669,N_4158);
nand U5201 (N_5201,N_4746,N_4780);
xor U5202 (N_5202,N_4136,N_4771);
nor U5203 (N_5203,N_4234,N_4595);
xor U5204 (N_5204,N_4791,N_4406);
nor U5205 (N_5205,N_4868,N_4003);
nor U5206 (N_5206,N_4638,N_4122);
or U5207 (N_5207,N_4634,N_4958);
xnor U5208 (N_5208,N_4811,N_4176);
and U5209 (N_5209,N_4882,N_4213);
nand U5210 (N_5210,N_4969,N_4173);
nor U5211 (N_5211,N_4442,N_4064);
xor U5212 (N_5212,N_4070,N_4500);
xnor U5213 (N_5213,N_4768,N_4322);
nor U5214 (N_5214,N_4138,N_4520);
or U5215 (N_5215,N_4376,N_4336);
nor U5216 (N_5216,N_4109,N_4416);
and U5217 (N_5217,N_4453,N_4816);
nand U5218 (N_5218,N_4837,N_4761);
and U5219 (N_5219,N_4080,N_4648);
and U5220 (N_5220,N_4007,N_4622);
and U5221 (N_5221,N_4675,N_4794);
or U5222 (N_5222,N_4378,N_4393);
and U5223 (N_5223,N_4971,N_4774);
or U5224 (N_5224,N_4214,N_4312);
and U5225 (N_5225,N_4069,N_4465);
nand U5226 (N_5226,N_4906,N_4043);
and U5227 (N_5227,N_4425,N_4281);
nor U5228 (N_5228,N_4289,N_4897);
nor U5229 (N_5229,N_4682,N_4335);
nand U5230 (N_5230,N_4824,N_4250);
nor U5231 (N_5231,N_4169,N_4503);
nand U5232 (N_5232,N_4528,N_4609);
nor U5233 (N_5233,N_4635,N_4457);
nor U5234 (N_5234,N_4265,N_4538);
nor U5235 (N_5235,N_4345,N_4623);
xor U5236 (N_5236,N_4028,N_4309);
nand U5237 (N_5237,N_4506,N_4112);
and U5238 (N_5238,N_4921,N_4749);
or U5239 (N_5239,N_4147,N_4157);
nand U5240 (N_5240,N_4929,N_4362);
nand U5241 (N_5241,N_4415,N_4576);
or U5242 (N_5242,N_4822,N_4719);
or U5243 (N_5243,N_4179,N_4834);
nand U5244 (N_5244,N_4263,N_4926);
and U5245 (N_5245,N_4973,N_4282);
or U5246 (N_5246,N_4238,N_4976);
xor U5247 (N_5247,N_4904,N_4825);
nand U5248 (N_5248,N_4728,N_4298);
or U5249 (N_5249,N_4202,N_4605);
or U5250 (N_5250,N_4991,N_4582);
xnor U5251 (N_5251,N_4367,N_4221);
nand U5252 (N_5252,N_4119,N_4407);
or U5253 (N_5253,N_4722,N_4553);
xnor U5254 (N_5254,N_4664,N_4655);
or U5255 (N_5255,N_4149,N_4354);
nand U5256 (N_5256,N_4451,N_4020);
nor U5257 (N_5257,N_4195,N_4229);
or U5258 (N_5258,N_4304,N_4259);
or U5259 (N_5259,N_4953,N_4463);
nand U5260 (N_5260,N_4637,N_4094);
or U5261 (N_5261,N_4821,N_4346);
nand U5262 (N_5262,N_4711,N_4742);
nor U5263 (N_5263,N_4769,N_4848);
or U5264 (N_5264,N_4255,N_4562);
xor U5265 (N_5265,N_4885,N_4754);
or U5266 (N_5266,N_4012,N_4498);
nand U5267 (N_5267,N_4373,N_4961);
and U5268 (N_5268,N_4353,N_4762);
xor U5269 (N_5269,N_4490,N_4479);
and U5270 (N_5270,N_4545,N_4533);
or U5271 (N_5271,N_4470,N_4643);
nor U5272 (N_5272,N_4881,N_4686);
xnor U5273 (N_5273,N_4878,N_4679);
and U5274 (N_5274,N_4260,N_4299);
and U5275 (N_5275,N_4757,N_4115);
and U5276 (N_5276,N_4271,N_4480);
nor U5277 (N_5277,N_4736,N_4400);
and U5278 (N_5278,N_4246,N_4812);
nand U5279 (N_5279,N_4579,N_4931);
xor U5280 (N_5280,N_4232,N_4242);
and U5281 (N_5281,N_4876,N_4117);
or U5282 (N_5282,N_4713,N_4357);
xor U5283 (N_5283,N_4555,N_4891);
xnor U5284 (N_5284,N_4310,N_4739);
nor U5285 (N_5285,N_4680,N_4172);
or U5286 (N_5286,N_4899,N_4423);
and U5287 (N_5287,N_4540,N_4922);
nand U5288 (N_5288,N_4370,N_4984);
and U5289 (N_5289,N_4476,N_4965);
nand U5290 (N_5290,N_4316,N_4351);
or U5291 (N_5291,N_4586,N_4445);
xor U5292 (N_5292,N_4032,N_4031);
or U5293 (N_5293,N_4181,N_4601);
or U5294 (N_5294,N_4444,N_4744);
or U5295 (N_5295,N_4775,N_4875);
and U5296 (N_5296,N_4797,N_4750);
nor U5297 (N_5297,N_4862,N_4523);
xnor U5298 (N_5298,N_4067,N_4047);
and U5299 (N_5299,N_4752,N_4105);
xnor U5300 (N_5300,N_4391,N_4670);
nor U5301 (N_5301,N_4704,N_4120);
and U5302 (N_5302,N_4183,N_4394);
or U5303 (N_5303,N_4053,N_4430);
or U5304 (N_5304,N_4941,N_4805);
nand U5305 (N_5305,N_4071,N_4022);
xnor U5306 (N_5306,N_4959,N_4083);
or U5307 (N_5307,N_4577,N_4302);
nand U5308 (N_5308,N_4801,N_4027);
nor U5309 (N_5309,N_4349,N_4334);
xnor U5310 (N_5310,N_4802,N_4082);
or U5311 (N_5311,N_4180,N_4598);
nand U5312 (N_5312,N_4809,N_4928);
nor U5313 (N_5313,N_4857,N_4541);
or U5314 (N_5314,N_4657,N_4475);
or U5315 (N_5315,N_4676,N_4343);
or U5316 (N_5316,N_4589,N_4131);
nor U5317 (N_5317,N_4653,N_4981);
nand U5318 (N_5318,N_4734,N_4462);
and U5319 (N_5319,N_4701,N_4104);
nor U5320 (N_5320,N_4668,N_4964);
nand U5321 (N_5321,N_4712,N_4901);
nand U5322 (N_5322,N_4006,N_4235);
or U5323 (N_5323,N_4203,N_4735);
xnor U5324 (N_5324,N_4527,N_4795);
or U5325 (N_5325,N_4692,N_4274);
nor U5326 (N_5326,N_4986,N_4086);
or U5327 (N_5327,N_4140,N_4624);
nand U5328 (N_5328,N_4366,N_4800);
and U5329 (N_5329,N_4596,N_4305);
nand U5330 (N_5330,N_4186,N_4539);
nor U5331 (N_5331,N_4550,N_4072);
xnor U5332 (N_5332,N_4303,N_4455);
xor U5333 (N_5333,N_4564,N_4230);
nor U5334 (N_5334,N_4156,N_4485);
and U5335 (N_5335,N_4865,N_4193);
and U5336 (N_5336,N_4350,N_4152);
and U5337 (N_5337,N_4507,N_4151);
and U5338 (N_5338,N_4182,N_4102);
or U5339 (N_5339,N_4371,N_4392);
and U5340 (N_5340,N_4398,N_4732);
nor U5341 (N_5341,N_4592,N_4285);
nor U5342 (N_5342,N_4318,N_4066);
or U5343 (N_5343,N_4740,N_4688);
nor U5344 (N_5344,N_4661,N_4652);
or U5345 (N_5345,N_4225,N_4428);
nand U5346 (N_5346,N_4276,N_4977);
xnor U5347 (N_5347,N_4563,N_4024);
and U5348 (N_5348,N_4459,N_4062);
xnor U5349 (N_5349,N_4753,N_4748);
nor U5350 (N_5350,N_4052,N_4419);
nor U5351 (N_5351,N_4832,N_4877);
and U5352 (N_5352,N_4515,N_4016);
nand U5353 (N_5353,N_4033,N_4487);
nor U5354 (N_5354,N_4184,N_4766);
and U5355 (N_5355,N_4266,N_4262);
or U5356 (N_5356,N_4960,N_4626);
and U5357 (N_5357,N_4161,N_4948);
xor U5358 (N_5358,N_4483,N_4065);
and U5359 (N_5359,N_4685,N_4946);
xnor U5360 (N_5360,N_4620,N_4924);
nor U5361 (N_5361,N_4982,N_4516);
or U5362 (N_5362,N_4403,N_4251);
xnor U5363 (N_5363,N_4621,N_4017);
and U5364 (N_5364,N_4187,N_4856);
nor U5365 (N_5365,N_4013,N_4113);
and U5366 (N_5366,N_4178,N_4216);
and U5367 (N_5367,N_4204,N_4387);
nand U5368 (N_5368,N_4142,N_4776);
and U5369 (N_5369,N_4864,N_4300);
nor U5370 (N_5370,N_4593,N_4568);
xnor U5371 (N_5371,N_4933,N_4861);
or U5372 (N_5372,N_4208,N_4854);
and U5373 (N_5373,N_4226,N_4042);
nor U5374 (N_5374,N_4707,N_4585);
nor U5375 (N_5375,N_4277,N_4268);
and U5376 (N_5376,N_4074,N_4536);
xor U5377 (N_5377,N_4050,N_4645);
nor U5378 (N_5378,N_4347,N_4828);
and U5379 (N_5379,N_4360,N_4972);
nand U5380 (N_5380,N_4526,N_4039);
nor U5381 (N_5381,N_4135,N_4101);
xnor U5382 (N_5382,N_4190,N_4233);
or U5383 (N_5383,N_4833,N_4581);
nand U5384 (N_5384,N_4644,N_4936);
or U5385 (N_5385,N_4695,N_4209);
nor U5386 (N_5386,N_4075,N_4290);
xnor U5387 (N_5387,N_4438,N_4461);
nor U5388 (N_5388,N_4210,N_4481);
nor U5389 (N_5389,N_4374,N_4146);
xor U5390 (N_5390,N_4005,N_4641);
xnor U5391 (N_5391,N_4932,N_4524);
and U5392 (N_5392,N_4666,N_4040);
nor U5393 (N_5393,N_4011,N_4799);
or U5394 (N_5394,N_4863,N_4693);
nor U5395 (N_5395,N_4348,N_4845);
xnor U5396 (N_5396,N_4962,N_4359);
nand U5397 (N_5397,N_4957,N_4365);
nor U5398 (N_5398,N_4118,N_4110);
and U5399 (N_5399,N_4448,N_4573);
xor U5400 (N_5400,N_4035,N_4836);
nor U5401 (N_5401,N_4600,N_4829);
nand U5402 (N_5402,N_4571,N_4099);
or U5403 (N_5403,N_4838,N_4613);
nand U5404 (N_5404,N_4987,N_4580);
or U5405 (N_5405,N_4261,N_4817);
and U5406 (N_5406,N_4447,N_4046);
nor U5407 (N_5407,N_4174,N_4189);
or U5408 (N_5408,N_4384,N_4814);
nor U5409 (N_5409,N_4570,N_4619);
or U5410 (N_5410,N_4502,N_4446);
and U5411 (N_5411,N_4240,N_4141);
xor U5412 (N_5412,N_4968,N_4998);
xor U5413 (N_5413,N_4087,N_4414);
xor U5414 (N_5414,N_4244,N_4535);
or U5415 (N_5415,N_4036,N_4743);
nor U5416 (N_5416,N_4823,N_4970);
nor U5417 (N_5417,N_4903,N_4787);
and U5418 (N_5418,N_4325,N_4164);
xor U5419 (N_5419,N_4339,N_4636);
and U5420 (N_5420,N_4247,N_4361);
nand U5421 (N_5421,N_4111,N_4943);
or U5422 (N_5422,N_4895,N_4978);
xor U5423 (N_5423,N_4026,N_4295);
nand U5424 (N_5424,N_4256,N_4292);
xor U5425 (N_5425,N_4569,N_4079);
nand U5426 (N_5426,N_4831,N_4489);
xor U5427 (N_5427,N_4628,N_4873);
and U5428 (N_5428,N_4132,N_4992);
nor U5429 (N_5429,N_4737,N_4898);
nand U5430 (N_5430,N_4522,N_4249);
or U5431 (N_5431,N_4521,N_4989);
nand U5432 (N_5432,N_4018,N_4004);
xnor U5433 (N_5433,N_4588,N_4763);
xnor U5434 (N_5434,N_4942,N_4497);
nor U5435 (N_5435,N_4755,N_4165);
or U5436 (N_5436,N_4859,N_4985);
and U5437 (N_5437,N_4514,N_4009);
and U5438 (N_5438,N_4154,N_4100);
nor U5439 (N_5439,N_4702,N_4337);
nand U5440 (N_5440,N_4543,N_4658);
and U5441 (N_5441,N_4478,N_4513);
xor U5442 (N_5442,N_4207,N_4966);
and U5443 (N_5443,N_4185,N_4880);
xor U5444 (N_5444,N_4820,N_4574);
nand U5445 (N_5445,N_4163,N_4916);
nor U5446 (N_5446,N_4473,N_4827);
and U5447 (N_5447,N_4089,N_4654);
xnor U5448 (N_5448,N_4855,N_4674);
nand U5449 (N_5449,N_4044,N_4488);
or U5450 (N_5450,N_4168,N_4327);
nand U5451 (N_5451,N_4852,N_4951);
nor U5452 (N_5452,N_4917,N_4383);
and U5453 (N_5453,N_4632,N_4330);
and U5454 (N_5454,N_4546,N_4531);
nor U5455 (N_5455,N_4788,N_4994);
xor U5456 (N_5456,N_4810,N_4909);
xor U5457 (N_5457,N_4264,N_4324);
or U5458 (N_5458,N_4879,N_4839);
nand U5459 (N_5459,N_4975,N_4121);
or U5460 (N_5460,N_4510,N_4731);
or U5461 (N_5461,N_4280,N_4937);
xnor U5462 (N_5462,N_4396,N_4431);
or U5463 (N_5463,N_4269,N_4486);
nor U5464 (N_5464,N_4993,N_4696);
or U5465 (N_5465,N_4192,N_4382);
xor U5466 (N_5466,N_4798,N_4472);
and U5467 (N_5467,N_4440,N_4114);
nor U5468 (N_5468,N_4955,N_4170);
and U5469 (N_5469,N_4494,N_4399);
nand U5470 (N_5470,N_4980,N_4691);
and U5471 (N_5471,N_4709,N_4404);
nand U5472 (N_5472,N_4273,N_4912);
or U5473 (N_5473,N_4437,N_4212);
and U5474 (N_5474,N_4243,N_4703);
and U5475 (N_5475,N_4215,N_4129);
xnor U5476 (N_5476,N_4785,N_4919);
nand U5477 (N_5477,N_4342,N_4439);
nor U5478 (N_5478,N_4649,N_4468);
xor U5479 (N_5479,N_4077,N_4019);
nand U5480 (N_5480,N_4913,N_4726);
and U5481 (N_5481,N_4647,N_4160);
and U5482 (N_5482,N_4389,N_4738);
nand U5483 (N_5483,N_4706,N_4008);
nor U5484 (N_5484,N_4708,N_4433);
and U5485 (N_5485,N_4872,N_4784);
nand U5486 (N_5486,N_4697,N_4081);
nor U5487 (N_5487,N_4294,N_4727);
or U5488 (N_5488,N_4850,N_4410);
xor U5489 (N_5489,N_4402,N_4084);
nor U5490 (N_5490,N_4091,N_4381);
nor U5491 (N_5491,N_4617,N_4338);
or U5492 (N_5492,N_4217,N_4369);
or U5493 (N_5493,N_4386,N_4093);
nand U5494 (N_5494,N_4642,N_4048);
xnor U5495 (N_5495,N_4578,N_4239);
and U5496 (N_5496,N_4777,N_4869);
or U5497 (N_5497,N_4639,N_4542);
and U5498 (N_5498,N_4060,N_4293);
xor U5499 (N_5499,N_4380,N_4841);
or U5500 (N_5500,N_4074,N_4022);
and U5501 (N_5501,N_4846,N_4063);
xnor U5502 (N_5502,N_4264,N_4329);
or U5503 (N_5503,N_4876,N_4768);
nand U5504 (N_5504,N_4742,N_4616);
or U5505 (N_5505,N_4197,N_4798);
nand U5506 (N_5506,N_4467,N_4729);
and U5507 (N_5507,N_4404,N_4172);
and U5508 (N_5508,N_4448,N_4644);
and U5509 (N_5509,N_4669,N_4068);
nor U5510 (N_5510,N_4285,N_4470);
xnor U5511 (N_5511,N_4987,N_4600);
and U5512 (N_5512,N_4101,N_4675);
or U5513 (N_5513,N_4277,N_4294);
nor U5514 (N_5514,N_4841,N_4951);
nor U5515 (N_5515,N_4500,N_4052);
xnor U5516 (N_5516,N_4741,N_4681);
and U5517 (N_5517,N_4418,N_4505);
xor U5518 (N_5518,N_4787,N_4163);
nor U5519 (N_5519,N_4017,N_4565);
or U5520 (N_5520,N_4338,N_4832);
nor U5521 (N_5521,N_4827,N_4804);
xnor U5522 (N_5522,N_4815,N_4297);
nor U5523 (N_5523,N_4463,N_4334);
or U5524 (N_5524,N_4230,N_4396);
nand U5525 (N_5525,N_4416,N_4245);
nand U5526 (N_5526,N_4504,N_4874);
nand U5527 (N_5527,N_4064,N_4266);
xor U5528 (N_5528,N_4208,N_4365);
and U5529 (N_5529,N_4732,N_4222);
nand U5530 (N_5530,N_4531,N_4573);
nor U5531 (N_5531,N_4441,N_4107);
xor U5532 (N_5532,N_4602,N_4288);
xor U5533 (N_5533,N_4318,N_4718);
xnor U5534 (N_5534,N_4093,N_4957);
nor U5535 (N_5535,N_4714,N_4221);
nor U5536 (N_5536,N_4181,N_4234);
or U5537 (N_5537,N_4247,N_4471);
or U5538 (N_5538,N_4241,N_4261);
nor U5539 (N_5539,N_4273,N_4718);
nor U5540 (N_5540,N_4185,N_4916);
xnor U5541 (N_5541,N_4900,N_4197);
and U5542 (N_5542,N_4365,N_4360);
xor U5543 (N_5543,N_4577,N_4775);
xor U5544 (N_5544,N_4240,N_4634);
xnor U5545 (N_5545,N_4700,N_4679);
nor U5546 (N_5546,N_4735,N_4690);
nand U5547 (N_5547,N_4116,N_4604);
or U5548 (N_5548,N_4995,N_4048);
nor U5549 (N_5549,N_4808,N_4012);
nand U5550 (N_5550,N_4724,N_4224);
nor U5551 (N_5551,N_4320,N_4322);
nor U5552 (N_5552,N_4689,N_4347);
nor U5553 (N_5553,N_4535,N_4328);
and U5554 (N_5554,N_4307,N_4164);
and U5555 (N_5555,N_4795,N_4104);
nor U5556 (N_5556,N_4252,N_4083);
nor U5557 (N_5557,N_4607,N_4977);
nor U5558 (N_5558,N_4673,N_4911);
and U5559 (N_5559,N_4594,N_4033);
xor U5560 (N_5560,N_4028,N_4137);
and U5561 (N_5561,N_4727,N_4205);
nand U5562 (N_5562,N_4567,N_4504);
nand U5563 (N_5563,N_4833,N_4039);
or U5564 (N_5564,N_4290,N_4989);
xnor U5565 (N_5565,N_4211,N_4664);
or U5566 (N_5566,N_4155,N_4018);
nand U5567 (N_5567,N_4835,N_4356);
nor U5568 (N_5568,N_4793,N_4718);
xor U5569 (N_5569,N_4804,N_4632);
nand U5570 (N_5570,N_4353,N_4184);
nor U5571 (N_5571,N_4228,N_4646);
nor U5572 (N_5572,N_4806,N_4893);
nor U5573 (N_5573,N_4424,N_4317);
and U5574 (N_5574,N_4936,N_4765);
or U5575 (N_5575,N_4746,N_4171);
nor U5576 (N_5576,N_4981,N_4608);
nor U5577 (N_5577,N_4288,N_4607);
xnor U5578 (N_5578,N_4203,N_4652);
or U5579 (N_5579,N_4550,N_4439);
nand U5580 (N_5580,N_4672,N_4210);
nor U5581 (N_5581,N_4233,N_4813);
or U5582 (N_5582,N_4240,N_4492);
xor U5583 (N_5583,N_4385,N_4624);
nand U5584 (N_5584,N_4454,N_4183);
xnor U5585 (N_5585,N_4748,N_4849);
or U5586 (N_5586,N_4735,N_4020);
nor U5587 (N_5587,N_4737,N_4722);
and U5588 (N_5588,N_4536,N_4712);
or U5589 (N_5589,N_4754,N_4115);
xor U5590 (N_5590,N_4436,N_4316);
nor U5591 (N_5591,N_4270,N_4134);
xor U5592 (N_5592,N_4516,N_4533);
nor U5593 (N_5593,N_4357,N_4925);
and U5594 (N_5594,N_4714,N_4676);
nand U5595 (N_5595,N_4498,N_4429);
and U5596 (N_5596,N_4887,N_4176);
xnor U5597 (N_5597,N_4054,N_4812);
nor U5598 (N_5598,N_4818,N_4606);
xnor U5599 (N_5599,N_4927,N_4233);
or U5600 (N_5600,N_4349,N_4140);
nand U5601 (N_5601,N_4856,N_4595);
nand U5602 (N_5602,N_4855,N_4374);
nand U5603 (N_5603,N_4086,N_4195);
or U5604 (N_5604,N_4934,N_4931);
and U5605 (N_5605,N_4082,N_4045);
xnor U5606 (N_5606,N_4554,N_4264);
nand U5607 (N_5607,N_4502,N_4633);
and U5608 (N_5608,N_4496,N_4349);
nand U5609 (N_5609,N_4803,N_4633);
nand U5610 (N_5610,N_4092,N_4022);
nor U5611 (N_5611,N_4837,N_4916);
nor U5612 (N_5612,N_4099,N_4467);
and U5613 (N_5613,N_4324,N_4596);
or U5614 (N_5614,N_4708,N_4908);
nand U5615 (N_5615,N_4682,N_4001);
xor U5616 (N_5616,N_4256,N_4664);
nor U5617 (N_5617,N_4811,N_4515);
or U5618 (N_5618,N_4104,N_4131);
nor U5619 (N_5619,N_4033,N_4396);
xnor U5620 (N_5620,N_4994,N_4707);
and U5621 (N_5621,N_4335,N_4907);
xnor U5622 (N_5622,N_4687,N_4623);
nand U5623 (N_5623,N_4536,N_4880);
or U5624 (N_5624,N_4250,N_4649);
and U5625 (N_5625,N_4864,N_4236);
nor U5626 (N_5626,N_4274,N_4807);
nor U5627 (N_5627,N_4746,N_4449);
and U5628 (N_5628,N_4093,N_4204);
xor U5629 (N_5629,N_4484,N_4581);
nand U5630 (N_5630,N_4885,N_4648);
xnor U5631 (N_5631,N_4213,N_4591);
xor U5632 (N_5632,N_4208,N_4653);
nand U5633 (N_5633,N_4931,N_4366);
nor U5634 (N_5634,N_4052,N_4024);
or U5635 (N_5635,N_4865,N_4710);
xor U5636 (N_5636,N_4288,N_4473);
nor U5637 (N_5637,N_4539,N_4446);
or U5638 (N_5638,N_4553,N_4489);
nor U5639 (N_5639,N_4838,N_4494);
or U5640 (N_5640,N_4543,N_4108);
nor U5641 (N_5641,N_4183,N_4675);
and U5642 (N_5642,N_4196,N_4724);
nand U5643 (N_5643,N_4878,N_4198);
and U5644 (N_5644,N_4039,N_4262);
xor U5645 (N_5645,N_4054,N_4351);
or U5646 (N_5646,N_4492,N_4980);
or U5647 (N_5647,N_4609,N_4420);
and U5648 (N_5648,N_4107,N_4885);
nor U5649 (N_5649,N_4612,N_4773);
nor U5650 (N_5650,N_4714,N_4433);
and U5651 (N_5651,N_4611,N_4432);
nand U5652 (N_5652,N_4235,N_4377);
nor U5653 (N_5653,N_4212,N_4230);
or U5654 (N_5654,N_4367,N_4241);
xnor U5655 (N_5655,N_4625,N_4515);
and U5656 (N_5656,N_4786,N_4798);
xor U5657 (N_5657,N_4268,N_4858);
xor U5658 (N_5658,N_4815,N_4236);
and U5659 (N_5659,N_4250,N_4837);
nor U5660 (N_5660,N_4030,N_4079);
nand U5661 (N_5661,N_4261,N_4086);
xnor U5662 (N_5662,N_4130,N_4683);
nor U5663 (N_5663,N_4893,N_4554);
and U5664 (N_5664,N_4394,N_4258);
and U5665 (N_5665,N_4444,N_4318);
or U5666 (N_5666,N_4830,N_4276);
and U5667 (N_5667,N_4446,N_4953);
nor U5668 (N_5668,N_4497,N_4007);
xor U5669 (N_5669,N_4501,N_4248);
nand U5670 (N_5670,N_4288,N_4203);
and U5671 (N_5671,N_4948,N_4479);
or U5672 (N_5672,N_4594,N_4086);
nand U5673 (N_5673,N_4847,N_4902);
xnor U5674 (N_5674,N_4798,N_4484);
xnor U5675 (N_5675,N_4500,N_4060);
or U5676 (N_5676,N_4026,N_4287);
or U5677 (N_5677,N_4733,N_4234);
and U5678 (N_5678,N_4167,N_4687);
or U5679 (N_5679,N_4618,N_4680);
nand U5680 (N_5680,N_4525,N_4528);
and U5681 (N_5681,N_4010,N_4986);
and U5682 (N_5682,N_4331,N_4682);
xnor U5683 (N_5683,N_4597,N_4524);
nand U5684 (N_5684,N_4859,N_4328);
and U5685 (N_5685,N_4545,N_4184);
and U5686 (N_5686,N_4880,N_4902);
nor U5687 (N_5687,N_4962,N_4014);
nand U5688 (N_5688,N_4652,N_4082);
or U5689 (N_5689,N_4436,N_4726);
nand U5690 (N_5690,N_4846,N_4602);
xnor U5691 (N_5691,N_4278,N_4056);
nor U5692 (N_5692,N_4395,N_4176);
or U5693 (N_5693,N_4616,N_4198);
nand U5694 (N_5694,N_4851,N_4719);
xor U5695 (N_5695,N_4598,N_4769);
nand U5696 (N_5696,N_4820,N_4388);
nor U5697 (N_5697,N_4553,N_4282);
nand U5698 (N_5698,N_4987,N_4848);
nor U5699 (N_5699,N_4194,N_4503);
nand U5700 (N_5700,N_4370,N_4735);
nor U5701 (N_5701,N_4304,N_4808);
and U5702 (N_5702,N_4916,N_4062);
nor U5703 (N_5703,N_4701,N_4694);
nor U5704 (N_5704,N_4553,N_4849);
and U5705 (N_5705,N_4702,N_4348);
nor U5706 (N_5706,N_4865,N_4382);
or U5707 (N_5707,N_4596,N_4068);
and U5708 (N_5708,N_4723,N_4287);
or U5709 (N_5709,N_4199,N_4770);
xnor U5710 (N_5710,N_4839,N_4426);
nor U5711 (N_5711,N_4313,N_4971);
and U5712 (N_5712,N_4416,N_4697);
and U5713 (N_5713,N_4370,N_4122);
xnor U5714 (N_5714,N_4891,N_4943);
xnor U5715 (N_5715,N_4007,N_4267);
and U5716 (N_5716,N_4903,N_4187);
xnor U5717 (N_5717,N_4302,N_4162);
nor U5718 (N_5718,N_4025,N_4895);
nand U5719 (N_5719,N_4610,N_4928);
xnor U5720 (N_5720,N_4535,N_4166);
and U5721 (N_5721,N_4178,N_4428);
nand U5722 (N_5722,N_4022,N_4776);
xor U5723 (N_5723,N_4824,N_4403);
and U5724 (N_5724,N_4056,N_4994);
or U5725 (N_5725,N_4655,N_4351);
nand U5726 (N_5726,N_4107,N_4658);
and U5727 (N_5727,N_4807,N_4148);
nand U5728 (N_5728,N_4920,N_4510);
xor U5729 (N_5729,N_4732,N_4902);
nand U5730 (N_5730,N_4690,N_4479);
or U5731 (N_5731,N_4887,N_4470);
xor U5732 (N_5732,N_4128,N_4974);
xor U5733 (N_5733,N_4081,N_4635);
and U5734 (N_5734,N_4225,N_4148);
nor U5735 (N_5735,N_4539,N_4714);
or U5736 (N_5736,N_4261,N_4156);
nand U5737 (N_5737,N_4691,N_4907);
or U5738 (N_5738,N_4830,N_4709);
nand U5739 (N_5739,N_4804,N_4227);
xnor U5740 (N_5740,N_4923,N_4053);
nor U5741 (N_5741,N_4177,N_4193);
or U5742 (N_5742,N_4165,N_4150);
nor U5743 (N_5743,N_4031,N_4672);
nor U5744 (N_5744,N_4563,N_4650);
and U5745 (N_5745,N_4941,N_4301);
nand U5746 (N_5746,N_4638,N_4457);
nand U5747 (N_5747,N_4533,N_4961);
and U5748 (N_5748,N_4860,N_4249);
xnor U5749 (N_5749,N_4683,N_4899);
xor U5750 (N_5750,N_4053,N_4806);
nand U5751 (N_5751,N_4086,N_4821);
and U5752 (N_5752,N_4715,N_4658);
nand U5753 (N_5753,N_4788,N_4052);
nor U5754 (N_5754,N_4526,N_4147);
nor U5755 (N_5755,N_4196,N_4132);
or U5756 (N_5756,N_4500,N_4991);
nand U5757 (N_5757,N_4374,N_4657);
nor U5758 (N_5758,N_4603,N_4730);
nor U5759 (N_5759,N_4682,N_4466);
xor U5760 (N_5760,N_4107,N_4781);
nand U5761 (N_5761,N_4447,N_4926);
or U5762 (N_5762,N_4274,N_4088);
nand U5763 (N_5763,N_4775,N_4718);
nand U5764 (N_5764,N_4877,N_4178);
xnor U5765 (N_5765,N_4541,N_4459);
and U5766 (N_5766,N_4346,N_4043);
and U5767 (N_5767,N_4053,N_4193);
and U5768 (N_5768,N_4586,N_4008);
or U5769 (N_5769,N_4485,N_4273);
or U5770 (N_5770,N_4225,N_4850);
nand U5771 (N_5771,N_4389,N_4592);
or U5772 (N_5772,N_4126,N_4141);
nor U5773 (N_5773,N_4860,N_4192);
nor U5774 (N_5774,N_4134,N_4553);
and U5775 (N_5775,N_4496,N_4847);
nor U5776 (N_5776,N_4091,N_4754);
nor U5777 (N_5777,N_4669,N_4661);
xnor U5778 (N_5778,N_4965,N_4330);
nand U5779 (N_5779,N_4592,N_4037);
nor U5780 (N_5780,N_4228,N_4802);
and U5781 (N_5781,N_4563,N_4755);
xnor U5782 (N_5782,N_4174,N_4295);
nor U5783 (N_5783,N_4891,N_4996);
xor U5784 (N_5784,N_4307,N_4442);
or U5785 (N_5785,N_4938,N_4441);
nor U5786 (N_5786,N_4248,N_4486);
nor U5787 (N_5787,N_4678,N_4326);
nand U5788 (N_5788,N_4548,N_4302);
xnor U5789 (N_5789,N_4504,N_4810);
or U5790 (N_5790,N_4101,N_4578);
nand U5791 (N_5791,N_4502,N_4744);
and U5792 (N_5792,N_4456,N_4069);
and U5793 (N_5793,N_4875,N_4502);
nand U5794 (N_5794,N_4422,N_4432);
nand U5795 (N_5795,N_4701,N_4697);
nand U5796 (N_5796,N_4958,N_4710);
and U5797 (N_5797,N_4018,N_4532);
nand U5798 (N_5798,N_4503,N_4267);
or U5799 (N_5799,N_4479,N_4015);
nor U5800 (N_5800,N_4710,N_4062);
nand U5801 (N_5801,N_4763,N_4820);
xnor U5802 (N_5802,N_4121,N_4419);
and U5803 (N_5803,N_4521,N_4282);
xnor U5804 (N_5804,N_4670,N_4448);
xor U5805 (N_5805,N_4643,N_4602);
xnor U5806 (N_5806,N_4698,N_4592);
or U5807 (N_5807,N_4893,N_4268);
or U5808 (N_5808,N_4753,N_4357);
and U5809 (N_5809,N_4272,N_4521);
nand U5810 (N_5810,N_4778,N_4686);
nand U5811 (N_5811,N_4470,N_4386);
nor U5812 (N_5812,N_4267,N_4143);
or U5813 (N_5813,N_4513,N_4841);
xnor U5814 (N_5814,N_4455,N_4397);
and U5815 (N_5815,N_4590,N_4455);
and U5816 (N_5816,N_4456,N_4887);
xor U5817 (N_5817,N_4348,N_4517);
nand U5818 (N_5818,N_4166,N_4574);
nand U5819 (N_5819,N_4137,N_4647);
nor U5820 (N_5820,N_4455,N_4613);
xnor U5821 (N_5821,N_4348,N_4803);
or U5822 (N_5822,N_4930,N_4911);
nand U5823 (N_5823,N_4008,N_4990);
nor U5824 (N_5824,N_4723,N_4877);
and U5825 (N_5825,N_4032,N_4670);
xnor U5826 (N_5826,N_4382,N_4309);
and U5827 (N_5827,N_4458,N_4366);
or U5828 (N_5828,N_4921,N_4525);
and U5829 (N_5829,N_4890,N_4768);
or U5830 (N_5830,N_4654,N_4004);
nand U5831 (N_5831,N_4884,N_4639);
or U5832 (N_5832,N_4032,N_4966);
or U5833 (N_5833,N_4985,N_4190);
or U5834 (N_5834,N_4574,N_4859);
and U5835 (N_5835,N_4572,N_4131);
and U5836 (N_5836,N_4953,N_4023);
and U5837 (N_5837,N_4969,N_4484);
nand U5838 (N_5838,N_4039,N_4708);
or U5839 (N_5839,N_4039,N_4127);
nand U5840 (N_5840,N_4897,N_4886);
xnor U5841 (N_5841,N_4264,N_4986);
or U5842 (N_5842,N_4684,N_4857);
or U5843 (N_5843,N_4635,N_4155);
xnor U5844 (N_5844,N_4825,N_4579);
xor U5845 (N_5845,N_4039,N_4981);
nand U5846 (N_5846,N_4088,N_4722);
nand U5847 (N_5847,N_4713,N_4797);
xor U5848 (N_5848,N_4928,N_4676);
nor U5849 (N_5849,N_4244,N_4784);
and U5850 (N_5850,N_4636,N_4253);
or U5851 (N_5851,N_4900,N_4550);
or U5852 (N_5852,N_4041,N_4232);
and U5853 (N_5853,N_4510,N_4164);
nor U5854 (N_5854,N_4685,N_4301);
nor U5855 (N_5855,N_4913,N_4084);
or U5856 (N_5856,N_4587,N_4905);
and U5857 (N_5857,N_4585,N_4002);
or U5858 (N_5858,N_4071,N_4597);
nand U5859 (N_5859,N_4662,N_4999);
xor U5860 (N_5860,N_4631,N_4425);
xor U5861 (N_5861,N_4710,N_4395);
or U5862 (N_5862,N_4140,N_4802);
and U5863 (N_5863,N_4611,N_4167);
xor U5864 (N_5864,N_4946,N_4042);
or U5865 (N_5865,N_4941,N_4526);
nand U5866 (N_5866,N_4997,N_4915);
nor U5867 (N_5867,N_4380,N_4981);
and U5868 (N_5868,N_4293,N_4471);
nand U5869 (N_5869,N_4634,N_4032);
nor U5870 (N_5870,N_4685,N_4454);
nand U5871 (N_5871,N_4615,N_4305);
nor U5872 (N_5872,N_4273,N_4198);
xor U5873 (N_5873,N_4930,N_4886);
nor U5874 (N_5874,N_4248,N_4053);
xor U5875 (N_5875,N_4428,N_4672);
xor U5876 (N_5876,N_4775,N_4079);
nor U5877 (N_5877,N_4302,N_4034);
nor U5878 (N_5878,N_4190,N_4253);
xnor U5879 (N_5879,N_4278,N_4052);
and U5880 (N_5880,N_4339,N_4453);
xnor U5881 (N_5881,N_4289,N_4477);
nand U5882 (N_5882,N_4216,N_4734);
nand U5883 (N_5883,N_4335,N_4766);
xnor U5884 (N_5884,N_4538,N_4579);
and U5885 (N_5885,N_4301,N_4604);
or U5886 (N_5886,N_4482,N_4822);
nand U5887 (N_5887,N_4128,N_4927);
nor U5888 (N_5888,N_4233,N_4300);
nor U5889 (N_5889,N_4635,N_4791);
or U5890 (N_5890,N_4628,N_4332);
nand U5891 (N_5891,N_4104,N_4988);
nor U5892 (N_5892,N_4092,N_4718);
nor U5893 (N_5893,N_4578,N_4958);
xnor U5894 (N_5894,N_4064,N_4859);
xnor U5895 (N_5895,N_4056,N_4347);
nand U5896 (N_5896,N_4418,N_4387);
or U5897 (N_5897,N_4806,N_4479);
xor U5898 (N_5898,N_4636,N_4182);
nand U5899 (N_5899,N_4547,N_4590);
and U5900 (N_5900,N_4494,N_4928);
xnor U5901 (N_5901,N_4302,N_4659);
xor U5902 (N_5902,N_4813,N_4255);
and U5903 (N_5903,N_4760,N_4856);
nand U5904 (N_5904,N_4937,N_4612);
and U5905 (N_5905,N_4552,N_4054);
xor U5906 (N_5906,N_4291,N_4693);
nand U5907 (N_5907,N_4989,N_4804);
nor U5908 (N_5908,N_4032,N_4453);
xor U5909 (N_5909,N_4948,N_4219);
nand U5910 (N_5910,N_4204,N_4117);
nand U5911 (N_5911,N_4476,N_4668);
and U5912 (N_5912,N_4927,N_4146);
or U5913 (N_5913,N_4096,N_4975);
nor U5914 (N_5914,N_4947,N_4932);
nor U5915 (N_5915,N_4677,N_4582);
and U5916 (N_5916,N_4515,N_4420);
or U5917 (N_5917,N_4348,N_4707);
nor U5918 (N_5918,N_4759,N_4658);
xnor U5919 (N_5919,N_4894,N_4310);
or U5920 (N_5920,N_4637,N_4051);
or U5921 (N_5921,N_4736,N_4347);
nand U5922 (N_5922,N_4617,N_4999);
nor U5923 (N_5923,N_4427,N_4230);
and U5924 (N_5924,N_4591,N_4548);
and U5925 (N_5925,N_4029,N_4476);
nand U5926 (N_5926,N_4588,N_4129);
or U5927 (N_5927,N_4187,N_4589);
xor U5928 (N_5928,N_4746,N_4936);
and U5929 (N_5929,N_4188,N_4400);
and U5930 (N_5930,N_4564,N_4319);
or U5931 (N_5931,N_4417,N_4036);
xnor U5932 (N_5932,N_4910,N_4550);
nand U5933 (N_5933,N_4398,N_4982);
or U5934 (N_5934,N_4586,N_4701);
nand U5935 (N_5935,N_4353,N_4282);
xor U5936 (N_5936,N_4927,N_4075);
xnor U5937 (N_5937,N_4312,N_4174);
nand U5938 (N_5938,N_4776,N_4257);
nor U5939 (N_5939,N_4233,N_4480);
xnor U5940 (N_5940,N_4566,N_4922);
and U5941 (N_5941,N_4570,N_4799);
nand U5942 (N_5942,N_4341,N_4166);
nand U5943 (N_5943,N_4037,N_4656);
or U5944 (N_5944,N_4991,N_4792);
nor U5945 (N_5945,N_4221,N_4879);
or U5946 (N_5946,N_4557,N_4001);
or U5947 (N_5947,N_4710,N_4877);
or U5948 (N_5948,N_4730,N_4388);
nor U5949 (N_5949,N_4266,N_4101);
or U5950 (N_5950,N_4469,N_4170);
xnor U5951 (N_5951,N_4202,N_4317);
or U5952 (N_5952,N_4038,N_4325);
and U5953 (N_5953,N_4780,N_4757);
xnor U5954 (N_5954,N_4398,N_4563);
nor U5955 (N_5955,N_4524,N_4925);
or U5956 (N_5956,N_4892,N_4182);
nand U5957 (N_5957,N_4939,N_4632);
xor U5958 (N_5958,N_4905,N_4377);
xnor U5959 (N_5959,N_4911,N_4515);
or U5960 (N_5960,N_4281,N_4276);
nor U5961 (N_5961,N_4183,N_4206);
nand U5962 (N_5962,N_4827,N_4162);
and U5963 (N_5963,N_4548,N_4592);
nor U5964 (N_5964,N_4619,N_4756);
or U5965 (N_5965,N_4037,N_4821);
nand U5966 (N_5966,N_4129,N_4792);
or U5967 (N_5967,N_4944,N_4076);
and U5968 (N_5968,N_4068,N_4920);
xor U5969 (N_5969,N_4563,N_4345);
nor U5970 (N_5970,N_4168,N_4964);
and U5971 (N_5971,N_4144,N_4758);
nor U5972 (N_5972,N_4932,N_4441);
nor U5973 (N_5973,N_4570,N_4454);
and U5974 (N_5974,N_4118,N_4691);
or U5975 (N_5975,N_4655,N_4524);
xor U5976 (N_5976,N_4547,N_4264);
nor U5977 (N_5977,N_4469,N_4544);
or U5978 (N_5978,N_4821,N_4678);
nand U5979 (N_5979,N_4564,N_4138);
nand U5980 (N_5980,N_4686,N_4136);
nor U5981 (N_5981,N_4265,N_4250);
xnor U5982 (N_5982,N_4499,N_4075);
nand U5983 (N_5983,N_4763,N_4682);
nor U5984 (N_5984,N_4065,N_4188);
or U5985 (N_5985,N_4486,N_4471);
nor U5986 (N_5986,N_4534,N_4591);
or U5987 (N_5987,N_4608,N_4587);
nor U5988 (N_5988,N_4371,N_4064);
nand U5989 (N_5989,N_4349,N_4540);
or U5990 (N_5990,N_4253,N_4496);
and U5991 (N_5991,N_4943,N_4654);
and U5992 (N_5992,N_4071,N_4358);
and U5993 (N_5993,N_4662,N_4290);
and U5994 (N_5994,N_4401,N_4458);
or U5995 (N_5995,N_4612,N_4226);
xor U5996 (N_5996,N_4767,N_4186);
nor U5997 (N_5997,N_4605,N_4585);
nand U5998 (N_5998,N_4630,N_4069);
xor U5999 (N_5999,N_4647,N_4885);
and U6000 (N_6000,N_5481,N_5822);
or U6001 (N_6001,N_5299,N_5503);
or U6002 (N_6002,N_5614,N_5146);
xor U6003 (N_6003,N_5958,N_5625);
nor U6004 (N_6004,N_5566,N_5303);
nor U6005 (N_6005,N_5137,N_5794);
xnor U6006 (N_6006,N_5559,N_5834);
nor U6007 (N_6007,N_5861,N_5500);
xor U6008 (N_6008,N_5925,N_5831);
nor U6009 (N_6009,N_5067,N_5611);
or U6010 (N_6010,N_5434,N_5106);
xor U6011 (N_6011,N_5134,N_5766);
and U6012 (N_6012,N_5962,N_5363);
and U6013 (N_6013,N_5360,N_5804);
nor U6014 (N_6014,N_5180,N_5882);
nor U6015 (N_6015,N_5581,N_5410);
xor U6016 (N_6016,N_5467,N_5632);
and U6017 (N_6017,N_5194,N_5457);
xnor U6018 (N_6018,N_5189,N_5668);
xor U6019 (N_6019,N_5000,N_5098);
or U6020 (N_6020,N_5842,N_5331);
nand U6021 (N_6021,N_5865,N_5480);
nand U6022 (N_6022,N_5791,N_5589);
nand U6023 (N_6023,N_5102,N_5319);
xor U6024 (N_6024,N_5711,N_5395);
xnor U6025 (N_6025,N_5693,N_5095);
xnor U6026 (N_6026,N_5600,N_5411);
and U6027 (N_6027,N_5918,N_5291);
nand U6028 (N_6028,N_5634,N_5305);
and U6029 (N_6029,N_5704,N_5629);
nand U6030 (N_6030,N_5343,N_5317);
nand U6031 (N_6031,N_5728,N_5264);
nor U6032 (N_6032,N_5252,N_5341);
or U6033 (N_6033,N_5933,N_5857);
nand U6034 (N_6034,N_5033,N_5565);
nor U6035 (N_6035,N_5945,N_5090);
or U6036 (N_6036,N_5475,N_5825);
nand U6037 (N_6037,N_5172,N_5263);
nor U6038 (N_6038,N_5655,N_5531);
nand U6039 (N_6039,N_5409,N_5726);
and U6040 (N_6040,N_5368,N_5162);
xnor U6041 (N_6041,N_5056,N_5024);
nor U6042 (N_6042,N_5673,N_5029);
and U6043 (N_6043,N_5876,N_5860);
and U6044 (N_6044,N_5519,N_5008);
xor U6045 (N_6045,N_5312,N_5381);
xor U6046 (N_6046,N_5406,N_5851);
or U6047 (N_6047,N_5687,N_5462);
nand U6048 (N_6048,N_5883,N_5520);
nand U6049 (N_6049,N_5719,N_5278);
or U6050 (N_6050,N_5710,N_5377);
nand U6051 (N_6051,N_5209,N_5088);
xnor U6052 (N_6052,N_5809,N_5929);
xor U6053 (N_6053,N_5890,N_5778);
and U6054 (N_6054,N_5070,N_5646);
xnor U6055 (N_6055,N_5679,N_5527);
xnor U6056 (N_6056,N_5229,N_5853);
and U6057 (N_6057,N_5960,N_5402);
nor U6058 (N_6058,N_5613,N_5157);
xor U6059 (N_6059,N_5554,N_5714);
or U6060 (N_6060,N_5596,N_5562);
or U6061 (N_6061,N_5703,N_5281);
nand U6062 (N_6062,N_5751,N_5866);
nand U6063 (N_6063,N_5709,N_5142);
nand U6064 (N_6064,N_5366,N_5170);
nor U6065 (N_6065,N_5132,N_5147);
nand U6066 (N_6066,N_5222,N_5574);
and U6067 (N_6067,N_5419,N_5228);
or U6068 (N_6068,N_5980,N_5570);
xor U6069 (N_6069,N_5948,N_5082);
and U6070 (N_6070,N_5805,N_5294);
nand U6071 (N_6071,N_5062,N_5735);
and U6072 (N_6072,N_5760,N_5211);
nand U6073 (N_6073,N_5010,N_5824);
and U6074 (N_6074,N_5885,N_5829);
or U6075 (N_6075,N_5666,N_5014);
and U6076 (N_6076,N_5595,N_5028);
nand U6077 (N_6077,N_5961,N_5894);
and U6078 (N_6078,N_5425,N_5167);
or U6079 (N_6079,N_5682,N_5889);
nor U6080 (N_6080,N_5787,N_5260);
xor U6081 (N_6081,N_5548,N_5997);
xnor U6082 (N_6082,N_5196,N_5237);
xnor U6083 (N_6083,N_5799,N_5350);
nor U6084 (N_6084,N_5064,N_5922);
nand U6085 (N_6085,N_5286,N_5854);
xor U6086 (N_6086,N_5987,N_5205);
nand U6087 (N_6087,N_5226,N_5455);
nor U6088 (N_6088,N_5351,N_5964);
xnor U6089 (N_6089,N_5246,N_5768);
xnor U6090 (N_6090,N_5466,N_5207);
and U6091 (N_6091,N_5145,N_5645);
xnor U6092 (N_6092,N_5727,N_5582);
nand U6093 (N_6093,N_5275,N_5869);
nand U6094 (N_6094,N_5521,N_5685);
or U6095 (N_6095,N_5290,N_5542);
xor U6096 (N_6096,N_5654,N_5561);
xor U6097 (N_6097,N_5691,N_5387);
xnor U6098 (N_6098,N_5598,N_5620);
and U6099 (N_6099,N_5392,N_5848);
or U6100 (N_6100,N_5050,N_5659);
nand U6101 (N_6101,N_5233,N_5111);
and U6102 (N_6102,N_5692,N_5470);
or U6103 (N_6103,N_5524,N_5605);
and U6104 (N_6104,N_5790,N_5285);
xor U6105 (N_6105,N_5255,N_5954);
or U6106 (N_6106,N_5405,N_5909);
and U6107 (N_6107,N_5585,N_5742);
xnor U6108 (N_6108,N_5274,N_5946);
nand U6109 (N_6109,N_5429,N_5713);
nor U6110 (N_6110,N_5232,N_5543);
or U6111 (N_6111,N_5269,N_5238);
nor U6112 (N_6112,N_5720,N_5849);
nor U6113 (N_6113,N_5771,N_5583);
xnor U6114 (N_6114,N_5783,N_5204);
xor U6115 (N_6115,N_5210,N_5136);
and U6116 (N_6116,N_5268,N_5875);
and U6117 (N_6117,N_5036,N_5432);
nand U6118 (N_6118,N_5427,N_5642);
and U6119 (N_6119,N_5151,N_5117);
nor U6120 (N_6120,N_5216,N_5374);
xor U6121 (N_6121,N_5532,N_5996);
nand U6122 (N_6122,N_5840,N_5079);
and U6123 (N_6123,N_5498,N_5337);
xnor U6124 (N_6124,N_5287,N_5575);
or U6125 (N_6125,N_5573,N_5253);
xor U6126 (N_6126,N_5934,N_5115);
nor U6127 (N_6127,N_5820,N_5164);
and U6128 (N_6128,N_5324,N_5176);
nor U6129 (N_6129,N_5459,N_5345);
nand U6130 (N_6130,N_5049,N_5334);
nand U6131 (N_6131,N_5579,N_5318);
or U6132 (N_6132,N_5718,N_5731);
nor U6133 (N_6133,N_5295,N_5073);
or U6134 (N_6134,N_5746,N_5065);
xnor U6135 (N_6135,N_5097,N_5414);
or U6136 (N_6136,N_5843,N_5203);
xor U6137 (N_6137,N_5112,N_5956);
xnor U6138 (N_6138,N_5775,N_5418);
and U6139 (N_6139,N_5915,N_5650);
nor U6140 (N_6140,N_5302,N_5638);
nor U6141 (N_6141,N_5917,N_5523);
and U6142 (N_6142,N_5931,N_5884);
xnor U6143 (N_6143,N_5382,N_5332);
or U6144 (N_6144,N_5362,N_5221);
nand U6145 (N_6145,N_5160,N_5072);
and U6146 (N_6146,N_5227,N_5348);
nor U6147 (N_6147,N_5386,N_5688);
and U6148 (N_6148,N_5636,N_5124);
nor U6149 (N_6149,N_5725,N_5802);
nand U6150 (N_6150,N_5603,N_5389);
or U6151 (N_6151,N_5431,N_5150);
and U6152 (N_6152,N_5712,N_5335);
or U6153 (N_6153,N_5858,N_5670);
and U6154 (N_6154,N_5896,N_5533);
nor U6155 (N_6155,N_5702,N_5320);
nor U6156 (N_6156,N_5732,N_5736);
and U6157 (N_6157,N_5902,N_5506);
nor U6158 (N_6158,N_5208,N_5384);
and U6159 (N_6159,N_5900,N_5743);
or U6160 (N_6160,N_5747,N_5830);
xor U6161 (N_6161,N_5789,N_5880);
and U6162 (N_6162,N_5788,N_5501);
or U6163 (N_6163,N_5174,N_5623);
nand U6164 (N_6164,N_5104,N_5738);
nand U6165 (N_6165,N_5510,N_5639);
or U6166 (N_6166,N_5779,N_5445);
and U6167 (N_6167,N_5930,N_5708);
or U6168 (N_6168,N_5927,N_5017);
and U6169 (N_6169,N_5982,N_5141);
nand U6170 (N_6170,N_5950,N_5616);
nand U6171 (N_6171,N_5754,N_5576);
xnor U6172 (N_6172,N_5259,N_5539);
nor U6173 (N_6173,N_5753,N_5247);
and U6174 (N_6174,N_5085,N_5535);
xnor U6175 (N_6175,N_5367,N_5109);
and U6176 (N_6176,N_5606,N_5555);
xnor U6177 (N_6177,N_5206,N_5947);
xor U6178 (N_6178,N_5154,N_5664);
xor U6179 (N_6179,N_5817,N_5344);
and U6180 (N_6180,N_5378,N_5422);
nor U6181 (N_6181,N_5936,N_5550);
nand U6182 (N_6182,N_5737,N_5558);
or U6183 (N_6183,N_5383,N_5248);
and U6184 (N_6184,N_5499,N_5235);
or U6185 (N_6185,N_5144,N_5156);
nor U6186 (N_6186,N_5618,N_5730);
xor U6187 (N_6187,N_5800,N_5676);
nor U6188 (N_6188,N_5166,N_5298);
xnor U6189 (N_6189,N_5888,N_5647);
or U6190 (N_6190,N_5450,N_5877);
and U6191 (N_6191,N_5916,N_5163);
xor U6192 (N_6192,N_5356,N_5069);
xnor U6193 (N_6193,N_5035,N_5213);
nand U6194 (N_6194,N_5919,N_5796);
xor U6195 (N_6195,N_5135,N_5179);
xnor U6196 (N_6196,N_5224,N_5546);
and U6197 (N_6197,N_5453,N_5258);
xnor U6198 (N_6198,N_5031,N_5644);
and U6199 (N_6199,N_5155,N_5949);
or U6200 (N_6200,N_5507,N_5012);
nand U6201 (N_6201,N_5850,N_5397);
nand U6202 (N_6202,N_5741,N_5953);
and U6203 (N_6203,N_5214,N_5610);
xor U6204 (N_6204,N_5188,N_5630);
and U6205 (N_6205,N_5801,N_5707);
nor U6206 (N_6206,N_5110,N_5828);
xor U6207 (N_6207,N_5242,N_5143);
xnor U6208 (N_6208,N_5631,N_5340);
and U6209 (N_6209,N_5966,N_5261);
xnor U6210 (N_6210,N_5841,N_5806);
and U6211 (N_6211,N_5512,N_5046);
nand U6212 (N_6212,N_5185,N_5973);
or U6213 (N_6213,N_5059,N_5477);
and U6214 (N_6214,N_5119,N_5832);
xnor U6215 (N_6215,N_5476,N_5123);
nor U6216 (N_6216,N_5231,N_5084);
and U6217 (N_6217,N_5451,N_5182);
and U6218 (N_6218,N_5094,N_5473);
nor U6219 (N_6219,N_5458,N_5895);
nor U6220 (N_6220,N_5680,N_5417);
nand U6221 (N_6221,N_5637,N_5080);
nand U6222 (N_6222,N_5810,N_5016);
nand U6223 (N_6223,N_5525,N_5391);
nand U6224 (N_6224,N_5826,N_5990);
and U6225 (N_6225,N_5026,N_5325);
or U6226 (N_6226,N_5752,N_5364);
nand U6227 (N_6227,N_5131,N_5460);
or U6228 (N_6228,N_5549,N_5660);
or U6229 (N_6229,N_5672,N_5159);
xor U6230 (N_6230,N_5483,N_5923);
and U6231 (N_6231,N_5358,N_5745);
nand U6232 (N_6232,N_5717,N_5552);
nor U6233 (N_6233,N_5300,N_5484);
and U6234 (N_6234,N_5288,N_5590);
and U6235 (N_6235,N_5140,N_5905);
and U6236 (N_6236,N_5813,N_5836);
nand U6237 (N_6237,N_5497,N_5658);
and U6238 (N_6238,N_5058,N_5441);
and U6239 (N_6239,N_5403,N_5330);
nand U6240 (N_6240,N_5436,N_5492);
nor U6241 (N_6241,N_5220,N_5128);
xor U6242 (N_6242,N_5764,N_5283);
nor U6243 (N_6243,N_5706,N_5812);
nor U6244 (N_6244,N_5744,N_5852);
or U6245 (N_6245,N_5514,N_5133);
nor U6246 (N_6246,N_5906,N_5551);
nand U6247 (N_6247,N_5357,N_5149);
nor U6248 (N_6248,N_5308,N_5661);
and U6249 (N_6249,N_5273,N_5845);
and U6250 (N_6250,N_5592,N_5380);
nor U6251 (N_6251,N_5243,N_5969);
and U6252 (N_6252,N_5886,N_5025);
nand U6253 (N_6253,N_5011,N_5602);
or U6254 (N_6254,N_5505,N_5517);
and U6255 (N_6255,N_5249,N_5700);
or U6256 (N_6256,N_5002,N_5256);
xnor U6257 (N_6257,N_5023,N_5584);
or U6258 (N_6258,N_5939,N_5859);
or U6259 (N_6259,N_5621,N_5161);
or U6260 (N_6260,N_5926,N_5245);
nor U6261 (N_6261,N_5393,N_5201);
nor U6262 (N_6262,N_5547,N_5669);
nand U6263 (N_6263,N_5994,N_5667);
xnor U6264 (N_6264,N_5018,N_5270);
xor U6265 (N_6265,N_5433,N_5986);
or U6266 (N_6266,N_5729,N_5045);
and U6267 (N_6267,N_5974,N_5093);
or U6268 (N_6268,N_5001,N_5219);
and U6269 (N_6269,N_5438,N_5478);
and U6270 (N_6270,N_5536,N_5911);
or U6271 (N_6271,N_5495,N_5296);
nor U6272 (N_6272,N_5597,N_5217);
and U6273 (N_6273,N_5181,N_5626);
and U6274 (N_6274,N_5178,N_5758);
or U6275 (N_6275,N_5336,N_5165);
nor U6276 (N_6276,N_5284,N_5148);
or U6277 (N_6277,N_5988,N_5773);
or U6278 (N_6278,N_5469,N_5716);
and U6279 (N_6279,N_5041,N_5116);
nor U6280 (N_6280,N_5223,N_5254);
and U6281 (N_6281,N_5599,N_5624);
nand U6282 (N_6282,N_5657,N_5797);
and U6283 (N_6283,N_5516,N_5748);
or U6284 (N_6284,N_5421,N_5957);
or U6285 (N_6285,N_5092,N_5347);
or U6286 (N_6286,N_5656,N_5490);
nand U6287 (N_6287,N_5793,N_5370);
nand U6288 (N_6288,N_5617,N_5904);
xor U6289 (N_6289,N_5122,N_5442);
nand U6290 (N_6290,N_5424,N_5540);
and U6291 (N_6291,N_5127,N_5100);
or U6292 (N_6292,N_5329,N_5267);
and U6293 (N_6293,N_5870,N_5928);
nor U6294 (N_6294,N_5769,N_5282);
or U6295 (N_6295,N_5463,N_5169);
or U6296 (N_6296,N_5408,N_5833);
or U6297 (N_6297,N_5053,N_5563);
or U6298 (N_6298,N_5030,N_5932);
nor U6299 (N_6299,N_5091,N_5975);
nand U6300 (N_6300,N_5914,N_5239);
and U6301 (N_6301,N_5983,N_5878);
nand U6302 (N_6302,N_5578,N_5042);
nor U6303 (N_6303,N_5724,N_5921);
or U6304 (N_6304,N_5564,N_5407);
nand U6305 (N_6305,N_5199,N_5907);
or U6306 (N_6306,N_5537,N_5591);
xnor U6307 (N_6307,N_5643,N_5734);
xor U6308 (N_6308,N_5837,N_5153);
nor U6309 (N_6309,N_5952,N_5215);
or U6310 (N_6310,N_5971,N_5815);
nand U6311 (N_6311,N_5464,N_5272);
or U6312 (N_6312,N_5040,N_5819);
nor U6313 (N_6313,N_5529,N_5967);
or U6314 (N_6314,N_5013,N_5695);
nand U6315 (N_6315,N_5862,N_5998);
or U6316 (N_6316,N_5874,N_5435);
and U6317 (N_6317,N_5125,N_5494);
nor U6318 (N_6318,N_5782,N_5355);
xnor U6319 (N_6319,N_5863,N_5444);
nand U6320 (N_6320,N_5202,N_5635);
nor U6321 (N_6321,N_5474,N_5057);
nor U6322 (N_6322,N_5781,N_5081);
nand U6323 (N_6323,N_5037,N_5349);
nand U6324 (N_6324,N_5200,N_5675);
and U6325 (N_6325,N_5899,N_5003);
nand U6326 (N_6326,N_5177,N_5633);
nor U6327 (N_6327,N_5439,N_5640);
nand U6328 (N_6328,N_5394,N_5043);
or U6329 (N_6329,N_5047,N_5063);
or U6330 (N_6330,N_5118,N_5452);
xnor U6331 (N_6331,N_5965,N_5601);
nor U6332 (N_6332,N_5485,N_5423);
and U6333 (N_6333,N_5105,N_5129);
and U6334 (N_6334,N_5901,N_5981);
xor U6335 (N_6335,N_5006,N_5310);
xor U6336 (N_6336,N_5653,N_5152);
xnor U6337 (N_6337,N_5293,N_5491);
nand U6338 (N_6338,N_5019,N_5416);
xnor U6339 (N_6339,N_5471,N_5504);
or U6340 (N_6340,N_5526,N_5289);
and U6341 (N_6341,N_5066,N_5762);
and U6342 (N_6342,N_5044,N_5353);
or U6343 (N_6343,N_5847,N_5379);
or U6344 (N_6344,N_5671,N_5749);
xor U6345 (N_6345,N_5765,N_5985);
and U6346 (N_6346,N_5075,N_5039);
or U6347 (N_6347,N_5086,N_5587);
nand U6348 (N_6348,N_5448,N_5937);
and U6349 (N_6349,N_5912,N_5580);
or U6350 (N_6350,N_5972,N_5241);
nor U6351 (N_6351,N_5942,N_5257);
xor U6352 (N_6352,N_5530,N_5756);
xnor U6353 (N_6353,N_5995,N_5191);
and U6354 (N_6354,N_5114,N_5054);
and U6355 (N_6355,N_5686,N_5993);
and U6356 (N_6356,N_5944,N_5301);
or U6357 (N_6357,N_5184,N_5328);
and U6358 (N_6358,N_5113,N_5893);
xor U6359 (N_6359,N_5489,N_5440);
xnor U6360 (N_6360,N_5678,N_5398);
nand U6361 (N_6361,N_5622,N_5311);
or U6362 (N_6362,N_5873,N_5770);
nor U6363 (N_6363,N_5087,N_5404);
xnor U6364 (N_6364,N_5823,N_5887);
nand U6365 (N_6365,N_5327,N_5426);
and U6366 (N_6366,N_5354,N_5814);
and U6367 (N_6367,N_5486,N_5430);
and U6368 (N_6368,N_5138,N_5924);
or U6369 (N_6369,N_5538,N_5487);
nor U6370 (N_6370,N_5891,N_5681);
xnor U6371 (N_6371,N_5197,N_5342);
nand U6372 (N_6372,N_5609,N_5941);
nor U6373 (N_6373,N_5545,N_5651);
or U6374 (N_6374,N_5428,N_5740);
nand U6375 (N_6375,N_5662,N_5420);
xnor U6376 (N_6376,N_5557,N_5544);
nor U6377 (N_6377,N_5401,N_5715);
or U6378 (N_6378,N_5313,N_5465);
nand U6379 (N_6379,N_5007,N_5694);
nand U6380 (N_6380,N_5192,N_5352);
and U6381 (N_6381,N_5641,N_5868);
nor U6382 (N_6382,N_5615,N_5101);
xnor U6383 (N_6383,N_5415,N_5846);
xor U6384 (N_6384,N_5456,N_5195);
or U6385 (N_6385,N_5984,N_5339);
nand U6386 (N_6386,N_5078,N_5560);
or U6387 (N_6387,N_5071,N_5385);
and U6388 (N_6388,N_5240,N_5628);
nor U6389 (N_6389,N_5977,N_5761);
nor U6390 (N_6390,N_5183,N_5627);
nor U6391 (N_6391,N_5186,N_5277);
xor U6392 (N_6392,N_5276,N_5951);
or U6393 (N_6393,N_5055,N_5472);
xor U6394 (N_6394,N_5786,N_5292);
xnor U6395 (N_6395,N_5107,N_5307);
xor U6396 (N_6396,N_5879,N_5032);
nand U6397 (N_6397,N_5665,N_5777);
and U6398 (N_6398,N_5321,N_5060);
or U6399 (N_6399,N_5371,N_5004);
nor U6400 (N_6400,N_5103,N_5594);
xnor U6401 (N_6401,N_5897,N_5326);
xnor U6402 (N_6402,N_5443,N_5607);
xor U6403 (N_6403,N_5588,N_5571);
xnor U6404 (N_6404,N_5513,N_5808);
nand U6405 (N_6405,N_5772,N_5757);
nor U6406 (N_6406,N_5038,N_5864);
or U6407 (N_6407,N_5068,N_5586);
or U6408 (N_6408,N_5373,N_5970);
nor U6409 (N_6409,N_5322,N_5022);
xor U6410 (N_6410,N_5236,N_5612);
nor U6411 (N_6411,N_5839,N_5304);
and U6412 (N_6412,N_5396,N_5696);
or U6413 (N_6413,N_5187,N_5399);
xor U6414 (N_6414,N_5750,N_5314);
or U6415 (N_6415,N_5992,N_5976);
nor U6416 (N_6416,N_5803,N_5978);
nand U6417 (N_6417,N_5935,N_5323);
xnor U6418 (N_6418,N_5881,N_5908);
xnor U6419 (N_6419,N_5333,N_5158);
or U6420 (N_6420,N_5698,N_5785);
nor U6421 (N_6421,N_5518,N_5061);
nor U6422 (N_6422,N_5898,N_5999);
nor U6423 (N_6423,N_5556,N_5955);
or U6424 (N_6424,N_5774,N_5963);
xor U6425 (N_6425,N_5701,N_5509);
xnor U6426 (N_6426,N_5739,N_5528);
xnor U6427 (N_6427,N_5683,N_5684);
nand U6428 (N_6428,N_5892,N_5511);
xor U6429 (N_6429,N_5315,N_5938);
nor U6430 (N_6430,N_5173,N_5051);
xor U6431 (N_6431,N_5619,N_5234);
nor U6432 (N_6432,N_5108,N_5021);
nand U6433 (N_6433,N_5212,N_5130);
nor U6434 (N_6434,N_5569,N_5316);
or U6435 (N_6435,N_5541,N_5979);
xnor U6436 (N_6436,N_5346,N_5390);
and U6437 (N_6437,N_5674,N_5872);
or U6438 (N_6438,N_5991,N_5502);
nand U6439 (N_6439,N_5309,N_5076);
nor U6440 (N_6440,N_5297,N_5780);
nor U6441 (N_6441,N_5577,N_5369);
or U6442 (N_6442,N_5855,N_5365);
xnor U6443 (N_6443,N_5126,N_5871);
xor U6444 (N_6444,N_5005,N_5496);
nor U6445 (N_6445,N_5265,N_5723);
nand U6446 (N_6446,N_5856,N_5795);
nor U6447 (N_6447,N_5568,N_5910);
nor U6448 (N_6448,N_5722,N_5077);
and U6449 (N_6449,N_5608,N_5818);
or U6450 (N_6450,N_5776,N_5454);
nor U6451 (N_6451,N_5792,N_5649);
nor U6452 (N_6452,N_5461,N_5375);
xor U6453 (N_6453,N_5171,N_5361);
nand U6454 (N_6454,N_5811,N_5663);
xnor U6455 (N_6455,N_5553,N_5400);
nor U6456 (N_6456,N_5827,N_5755);
and U6457 (N_6457,N_5020,N_5244);
nor U6458 (N_6458,N_5677,N_5705);
nor U6459 (N_6459,N_5230,N_5593);
nand U6460 (N_6460,N_5648,N_5920);
nand U6461 (N_6461,N_5376,N_5689);
and U6462 (N_6462,N_5412,N_5493);
nor U6463 (N_6463,N_5652,N_5468);
or U6464 (N_6464,N_5096,N_5567);
or U6465 (N_6465,N_5388,N_5604);
xor U6466 (N_6466,N_5048,N_5074);
or U6467 (N_6467,N_5522,N_5218);
and U6468 (N_6468,N_5251,N_5437);
nand U6469 (N_6469,N_5099,N_5250);
nand U6470 (N_6470,N_5733,N_5446);
and U6471 (N_6471,N_5190,N_5359);
or U6472 (N_6472,N_5413,N_5015);
nor U6473 (N_6473,N_5534,N_5767);
and U6474 (N_6474,N_5844,N_5968);
nand U6475 (N_6475,N_5052,N_5449);
and U6476 (N_6476,N_5697,N_5508);
or U6477 (N_6477,N_5759,N_5798);
nand U6478 (N_6478,N_5479,N_5372);
or U6479 (N_6479,N_5262,N_5515);
nor U6480 (N_6480,N_5271,N_5083);
nor U6481 (N_6481,N_5784,N_5034);
nand U6482 (N_6482,N_5175,N_5821);
xor U6483 (N_6483,N_5338,N_5121);
nor U6484 (N_6484,N_5721,N_5198);
and U6485 (N_6485,N_5266,N_5488);
nor U6486 (N_6486,N_5572,N_5835);
and U6487 (N_6487,N_5838,N_5027);
nor U6488 (N_6488,N_5225,N_5306);
xor U6489 (N_6489,N_5690,N_5943);
xor U6490 (N_6490,N_5989,N_5168);
nor U6491 (N_6491,N_5009,N_5807);
or U6492 (N_6492,N_5280,N_5940);
and U6493 (N_6493,N_5482,N_5959);
nor U6494 (N_6494,N_5816,N_5763);
nor U6495 (N_6495,N_5139,N_5447);
and U6496 (N_6496,N_5867,N_5279);
xnor U6497 (N_6497,N_5120,N_5089);
xnor U6498 (N_6498,N_5699,N_5913);
and U6499 (N_6499,N_5903,N_5193);
and U6500 (N_6500,N_5999,N_5236);
xnor U6501 (N_6501,N_5351,N_5393);
nor U6502 (N_6502,N_5285,N_5337);
xor U6503 (N_6503,N_5015,N_5025);
and U6504 (N_6504,N_5642,N_5033);
nand U6505 (N_6505,N_5670,N_5309);
or U6506 (N_6506,N_5938,N_5773);
and U6507 (N_6507,N_5839,N_5342);
nor U6508 (N_6508,N_5496,N_5771);
or U6509 (N_6509,N_5457,N_5307);
and U6510 (N_6510,N_5571,N_5513);
or U6511 (N_6511,N_5928,N_5377);
xnor U6512 (N_6512,N_5550,N_5985);
xor U6513 (N_6513,N_5296,N_5790);
or U6514 (N_6514,N_5519,N_5407);
xnor U6515 (N_6515,N_5982,N_5339);
and U6516 (N_6516,N_5048,N_5383);
and U6517 (N_6517,N_5260,N_5386);
nor U6518 (N_6518,N_5804,N_5729);
nand U6519 (N_6519,N_5972,N_5588);
and U6520 (N_6520,N_5436,N_5254);
nor U6521 (N_6521,N_5946,N_5751);
nand U6522 (N_6522,N_5068,N_5679);
or U6523 (N_6523,N_5626,N_5341);
or U6524 (N_6524,N_5967,N_5610);
nand U6525 (N_6525,N_5570,N_5918);
nor U6526 (N_6526,N_5785,N_5399);
nor U6527 (N_6527,N_5643,N_5263);
nand U6528 (N_6528,N_5284,N_5323);
nor U6529 (N_6529,N_5942,N_5029);
or U6530 (N_6530,N_5947,N_5157);
nand U6531 (N_6531,N_5660,N_5731);
and U6532 (N_6532,N_5929,N_5402);
and U6533 (N_6533,N_5596,N_5929);
or U6534 (N_6534,N_5633,N_5252);
nor U6535 (N_6535,N_5927,N_5328);
or U6536 (N_6536,N_5913,N_5215);
xnor U6537 (N_6537,N_5141,N_5879);
nor U6538 (N_6538,N_5470,N_5724);
or U6539 (N_6539,N_5317,N_5843);
nand U6540 (N_6540,N_5155,N_5819);
nor U6541 (N_6541,N_5899,N_5805);
and U6542 (N_6542,N_5053,N_5690);
xor U6543 (N_6543,N_5604,N_5208);
and U6544 (N_6544,N_5641,N_5888);
or U6545 (N_6545,N_5630,N_5185);
or U6546 (N_6546,N_5650,N_5092);
nand U6547 (N_6547,N_5019,N_5434);
nand U6548 (N_6548,N_5922,N_5490);
xor U6549 (N_6549,N_5678,N_5672);
nand U6550 (N_6550,N_5927,N_5406);
or U6551 (N_6551,N_5810,N_5960);
xor U6552 (N_6552,N_5437,N_5404);
and U6553 (N_6553,N_5020,N_5842);
xor U6554 (N_6554,N_5789,N_5895);
xor U6555 (N_6555,N_5258,N_5995);
nand U6556 (N_6556,N_5763,N_5384);
and U6557 (N_6557,N_5494,N_5858);
nor U6558 (N_6558,N_5731,N_5056);
xor U6559 (N_6559,N_5087,N_5451);
nand U6560 (N_6560,N_5646,N_5297);
or U6561 (N_6561,N_5028,N_5729);
and U6562 (N_6562,N_5292,N_5804);
nand U6563 (N_6563,N_5930,N_5497);
or U6564 (N_6564,N_5941,N_5870);
and U6565 (N_6565,N_5375,N_5594);
and U6566 (N_6566,N_5573,N_5882);
xor U6567 (N_6567,N_5367,N_5172);
and U6568 (N_6568,N_5471,N_5161);
nor U6569 (N_6569,N_5460,N_5450);
xnor U6570 (N_6570,N_5091,N_5731);
or U6571 (N_6571,N_5181,N_5470);
nand U6572 (N_6572,N_5094,N_5176);
nand U6573 (N_6573,N_5688,N_5331);
xor U6574 (N_6574,N_5087,N_5574);
nor U6575 (N_6575,N_5956,N_5453);
nand U6576 (N_6576,N_5568,N_5641);
xor U6577 (N_6577,N_5949,N_5892);
xor U6578 (N_6578,N_5542,N_5540);
or U6579 (N_6579,N_5563,N_5329);
nand U6580 (N_6580,N_5583,N_5312);
and U6581 (N_6581,N_5881,N_5938);
or U6582 (N_6582,N_5175,N_5617);
nor U6583 (N_6583,N_5454,N_5742);
xor U6584 (N_6584,N_5674,N_5039);
nor U6585 (N_6585,N_5335,N_5325);
or U6586 (N_6586,N_5956,N_5200);
nand U6587 (N_6587,N_5753,N_5601);
nand U6588 (N_6588,N_5870,N_5998);
or U6589 (N_6589,N_5772,N_5341);
nor U6590 (N_6590,N_5935,N_5580);
xor U6591 (N_6591,N_5934,N_5167);
nor U6592 (N_6592,N_5854,N_5761);
or U6593 (N_6593,N_5671,N_5151);
or U6594 (N_6594,N_5291,N_5481);
and U6595 (N_6595,N_5046,N_5753);
xor U6596 (N_6596,N_5177,N_5002);
xor U6597 (N_6597,N_5163,N_5654);
nand U6598 (N_6598,N_5956,N_5185);
nor U6599 (N_6599,N_5379,N_5687);
or U6600 (N_6600,N_5868,N_5993);
nor U6601 (N_6601,N_5316,N_5829);
or U6602 (N_6602,N_5653,N_5971);
nor U6603 (N_6603,N_5040,N_5110);
or U6604 (N_6604,N_5311,N_5670);
and U6605 (N_6605,N_5278,N_5612);
nand U6606 (N_6606,N_5113,N_5010);
nor U6607 (N_6607,N_5849,N_5196);
nand U6608 (N_6608,N_5853,N_5625);
nor U6609 (N_6609,N_5529,N_5245);
or U6610 (N_6610,N_5740,N_5642);
and U6611 (N_6611,N_5288,N_5786);
nor U6612 (N_6612,N_5673,N_5724);
and U6613 (N_6613,N_5889,N_5550);
nand U6614 (N_6614,N_5758,N_5967);
xor U6615 (N_6615,N_5297,N_5248);
nor U6616 (N_6616,N_5595,N_5210);
nor U6617 (N_6617,N_5313,N_5909);
nand U6618 (N_6618,N_5913,N_5071);
xor U6619 (N_6619,N_5660,N_5411);
and U6620 (N_6620,N_5031,N_5447);
or U6621 (N_6621,N_5442,N_5918);
nor U6622 (N_6622,N_5704,N_5154);
xnor U6623 (N_6623,N_5440,N_5821);
xnor U6624 (N_6624,N_5718,N_5948);
nand U6625 (N_6625,N_5928,N_5231);
nand U6626 (N_6626,N_5600,N_5250);
and U6627 (N_6627,N_5895,N_5511);
xnor U6628 (N_6628,N_5620,N_5496);
and U6629 (N_6629,N_5246,N_5613);
xor U6630 (N_6630,N_5350,N_5994);
xor U6631 (N_6631,N_5787,N_5189);
nand U6632 (N_6632,N_5877,N_5191);
or U6633 (N_6633,N_5712,N_5683);
nand U6634 (N_6634,N_5213,N_5752);
nor U6635 (N_6635,N_5894,N_5011);
or U6636 (N_6636,N_5258,N_5097);
or U6637 (N_6637,N_5365,N_5081);
or U6638 (N_6638,N_5665,N_5575);
nor U6639 (N_6639,N_5892,N_5174);
and U6640 (N_6640,N_5624,N_5305);
nor U6641 (N_6641,N_5672,N_5077);
nor U6642 (N_6642,N_5082,N_5045);
nor U6643 (N_6643,N_5346,N_5196);
and U6644 (N_6644,N_5271,N_5626);
nand U6645 (N_6645,N_5885,N_5079);
nor U6646 (N_6646,N_5447,N_5039);
xor U6647 (N_6647,N_5601,N_5962);
or U6648 (N_6648,N_5017,N_5814);
and U6649 (N_6649,N_5844,N_5575);
xnor U6650 (N_6650,N_5132,N_5158);
and U6651 (N_6651,N_5730,N_5602);
nor U6652 (N_6652,N_5599,N_5435);
or U6653 (N_6653,N_5424,N_5415);
xor U6654 (N_6654,N_5358,N_5861);
and U6655 (N_6655,N_5059,N_5265);
nand U6656 (N_6656,N_5441,N_5874);
and U6657 (N_6657,N_5312,N_5833);
or U6658 (N_6658,N_5394,N_5279);
nand U6659 (N_6659,N_5950,N_5575);
nor U6660 (N_6660,N_5057,N_5283);
xnor U6661 (N_6661,N_5405,N_5231);
or U6662 (N_6662,N_5864,N_5006);
nand U6663 (N_6663,N_5911,N_5223);
or U6664 (N_6664,N_5217,N_5620);
nand U6665 (N_6665,N_5858,N_5291);
nor U6666 (N_6666,N_5977,N_5930);
or U6667 (N_6667,N_5831,N_5653);
and U6668 (N_6668,N_5990,N_5570);
xnor U6669 (N_6669,N_5244,N_5847);
nor U6670 (N_6670,N_5779,N_5725);
and U6671 (N_6671,N_5405,N_5426);
nand U6672 (N_6672,N_5023,N_5740);
or U6673 (N_6673,N_5141,N_5405);
nand U6674 (N_6674,N_5922,N_5176);
xor U6675 (N_6675,N_5707,N_5334);
and U6676 (N_6676,N_5931,N_5918);
and U6677 (N_6677,N_5843,N_5404);
and U6678 (N_6678,N_5145,N_5096);
nand U6679 (N_6679,N_5395,N_5177);
or U6680 (N_6680,N_5840,N_5127);
nand U6681 (N_6681,N_5652,N_5853);
xnor U6682 (N_6682,N_5492,N_5696);
nor U6683 (N_6683,N_5933,N_5639);
nor U6684 (N_6684,N_5538,N_5009);
nand U6685 (N_6685,N_5635,N_5868);
nor U6686 (N_6686,N_5833,N_5064);
xor U6687 (N_6687,N_5561,N_5069);
or U6688 (N_6688,N_5458,N_5869);
nor U6689 (N_6689,N_5930,N_5012);
and U6690 (N_6690,N_5581,N_5573);
nor U6691 (N_6691,N_5932,N_5131);
nor U6692 (N_6692,N_5819,N_5295);
xor U6693 (N_6693,N_5562,N_5108);
nor U6694 (N_6694,N_5802,N_5441);
xnor U6695 (N_6695,N_5105,N_5540);
or U6696 (N_6696,N_5497,N_5635);
and U6697 (N_6697,N_5152,N_5406);
nor U6698 (N_6698,N_5701,N_5144);
nor U6699 (N_6699,N_5327,N_5192);
xnor U6700 (N_6700,N_5869,N_5048);
or U6701 (N_6701,N_5013,N_5269);
and U6702 (N_6702,N_5943,N_5200);
and U6703 (N_6703,N_5407,N_5192);
or U6704 (N_6704,N_5101,N_5386);
or U6705 (N_6705,N_5664,N_5679);
xor U6706 (N_6706,N_5686,N_5189);
xor U6707 (N_6707,N_5355,N_5904);
xnor U6708 (N_6708,N_5468,N_5258);
and U6709 (N_6709,N_5182,N_5031);
nor U6710 (N_6710,N_5928,N_5483);
xnor U6711 (N_6711,N_5087,N_5695);
nand U6712 (N_6712,N_5829,N_5162);
and U6713 (N_6713,N_5783,N_5799);
or U6714 (N_6714,N_5222,N_5760);
nand U6715 (N_6715,N_5624,N_5793);
and U6716 (N_6716,N_5808,N_5816);
nand U6717 (N_6717,N_5014,N_5952);
and U6718 (N_6718,N_5323,N_5887);
or U6719 (N_6719,N_5038,N_5848);
or U6720 (N_6720,N_5951,N_5485);
nor U6721 (N_6721,N_5209,N_5978);
nor U6722 (N_6722,N_5692,N_5080);
and U6723 (N_6723,N_5074,N_5416);
nor U6724 (N_6724,N_5400,N_5089);
xor U6725 (N_6725,N_5376,N_5757);
xnor U6726 (N_6726,N_5966,N_5390);
xnor U6727 (N_6727,N_5687,N_5151);
or U6728 (N_6728,N_5766,N_5631);
or U6729 (N_6729,N_5833,N_5669);
xnor U6730 (N_6730,N_5790,N_5458);
nor U6731 (N_6731,N_5766,N_5654);
and U6732 (N_6732,N_5723,N_5518);
and U6733 (N_6733,N_5776,N_5185);
xnor U6734 (N_6734,N_5214,N_5729);
xor U6735 (N_6735,N_5385,N_5565);
and U6736 (N_6736,N_5099,N_5057);
or U6737 (N_6737,N_5754,N_5086);
or U6738 (N_6738,N_5612,N_5583);
and U6739 (N_6739,N_5804,N_5386);
or U6740 (N_6740,N_5255,N_5935);
nor U6741 (N_6741,N_5197,N_5401);
nand U6742 (N_6742,N_5776,N_5985);
nor U6743 (N_6743,N_5426,N_5370);
or U6744 (N_6744,N_5750,N_5289);
or U6745 (N_6745,N_5119,N_5922);
and U6746 (N_6746,N_5118,N_5611);
nand U6747 (N_6747,N_5644,N_5477);
and U6748 (N_6748,N_5054,N_5840);
and U6749 (N_6749,N_5791,N_5034);
and U6750 (N_6750,N_5723,N_5934);
or U6751 (N_6751,N_5216,N_5150);
or U6752 (N_6752,N_5634,N_5386);
or U6753 (N_6753,N_5795,N_5836);
nor U6754 (N_6754,N_5198,N_5404);
or U6755 (N_6755,N_5519,N_5170);
xnor U6756 (N_6756,N_5469,N_5020);
xor U6757 (N_6757,N_5825,N_5965);
xor U6758 (N_6758,N_5361,N_5353);
xnor U6759 (N_6759,N_5437,N_5689);
or U6760 (N_6760,N_5098,N_5078);
xnor U6761 (N_6761,N_5480,N_5511);
or U6762 (N_6762,N_5749,N_5949);
or U6763 (N_6763,N_5966,N_5042);
and U6764 (N_6764,N_5972,N_5133);
nor U6765 (N_6765,N_5531,N_5274);
or U6766 (N_6766,N_5028,N_5678);
or U6767 (N_6767,N_5854,N_5866);
nor U6768 (N_6768,N_5575,N_5823);
and U6769 (N_6769,N_5313,N_5316);
nand U6770 (N_6770,N_5524,N_5976);
or U6771 (N_6771,N_5761,N_5381);
or U6772 (N_6772,N_5660,N_5496);
and U6773 (N_6773,N_5578,N_5196);
nand U6774 (N_6774,N_5885,N_5901);
xor U6775 (N_6775,N_5081,N_5956);
nand U6776 (N_6776,N_5067,N_5428);
and U6777 (N_6777,N_5244,N_5953);
nor U6778 (N_6778,N_5293,N_5939);
xnor U6779 (N_6779,N_5980,N_5657);
or U6780 (N_6780,N_5264,N_5483);
and U6781 (N_6781,N_5108,N_5472);
xnor U6782 (N_6782,N_5016,N_5048);
xor U6783 (N_6783,N_5630,N_5724);
or U6784 (N_6784,N_5970,N_5167);
and U6785 (N_6785,N_5161,N_5958);
nor U6786 (N_6786,N_5443,N_5739);
nand U6787 (N_6787,N_5043,N_5292);
xor U6788 (N_6788,N_5979,N_5908);
or U6789 (N_6789,N_5434,N_5650);
or U6790 (N_6790,N_5203,N_5816);
and U6791 (N_6791,N_5078,N_5771);
nor U6792 (N_6792,N_5126,N_5553);
nand U6793 (N_6793,N_5980,N_5061);
nor U6794 (N_6794,N_5015,N_5539);
and U6795 (N_6795,N_5905,N_5263);
and U6796 (N_6796,N_5231,N_5269);
nor U6797 (N_6797,N_5577,N_5133);
nor U6798 (N_6798,N_5170,N_5168);
or U6799 (N_6799,N_5505,N_5567);
and U6800 (N_6800,N_5803,N_5408);
nand U6801 (N_6801,N_5768,N_5271);
nand U6802 (N_6802,N_5708,N_5992);
or U6803 (N_6803,N_5884,N_5138);
nand U6804 (N_6804,N_5108,N_5463);
or U6805 (N_6805,N_5591,N_5862);
nor U6806 (N_6806,N_5832,N_5055);
nor U6807 (N_6807,N_5622,N_5525);
xnor U6808 (N_6808,N_5035,N_5624);
nand U6809 (N_6809,N_5793,N_5781);
nor U6810 (N_6810,N_5450,N_5840);
xor U6811 (N_6811,N_5940,N_5748);
or U6812 (N_6812,N_5923,N_5608);
and U6813 (N_6813,N_5922,N_5139);
nor U6814 (N_6814,N_5106,N_5596);
nor U6815 (N_6815,N_5512,N_5944);
nand U6816 (N_6816,N_5257,N_5162);
and U6817 (N_6817,N_5148,N_5169);
nand U6818 (N_6818,N_5357,N_5037);
and U6819 (N_6819,N_5837,N_5875);
xor U6820 (N_6820,N_5434,N_5989);
or U6821 (N_6821,N_5666,N_5804);
xnor U6822 (N_6822,N_5676,N_5422);
nor U6823 (N_6823,N_5238,N_5010);
nor U6824 (N_6824,N_5776,N_5408);
nand U6825 (N_6825,N_5822,N_5597);
nor U6826 (N_6826,N_5529,N_5258);
xor U6827 (N_6827,N_5469,N_5912);
xor U6828 (N_6828,N_5314,N_5430);
or U6829 (N_6829,N_5427,N_5454);
and U6830 (N_6830,N_5549,N_5934);
and U6831 (N_6831,N_5656,N_5723);
nand U6832 (N_6832,N_5770,N_5376);
nor U6833 (N_6833,N_5055,N_5614);
or U6834 (N_6834,N_5580,N_5278);
and U6835 (N_6835,N_5709,N_5863);
xnor U6836 (N_6836,N_5698,N_5592);
or U6837 (N_6837,N_5524,N_5511);
xnor U6838 (N_6838,N_5576,N_5078);
nor U6839 (N_6839,N_5922,N_5391);
nand U6840 (N_6840,N_5426,N_5211);
xnor U6841 (N_6841,N_5856,N_5924);
nand U6842 (N_6842,N_5692,N_5982);
nand U6843 (N_6843,N_5206,N_5507);
xor U6844 (N_6844,N_5899,N_5329);
nand U6845 (N_6845,N_5292,N_5509);
or U6846 (N_6846,N_5424,N_5773);
or U6847 (N_6847,N_5570,N_5478);
nor U6848 (N_6848,N_5153,N_5957);
or U6849 (N_6849,N_5014,N_5080);
or U6850 (N_6850,N_5575,N_5813);
xor U6851 (N_6851,N_5217,N_5337);
nand U6852 (N_6852,N_5145,N_5513);
and U6853 (N_6853,N_5757,N_5220);
xnor U6854 (N_6854,N_5619,N_5514);
and U6855 (N_6855,N_5246,N_5430);
nor U6856 (N_6856,N_5618,N_5927);
nand U6857 (N_6857,N_5698,N_5023);
nand U6858 (N_6858,N_5604,N_5310);
and U6859 (N_6859,N_5579,N_5497);
and U6860 (N_6860,N_5506,N_5057);
and U6861 (N_6861,N_5407,N_5084);
nor U6862 (N_6862,N_5306,N_5470);
and U6863 (N_6863,N_5365,N_5953);
and U6864 (N_6864,N_5230,N_5194);
xnor U6865 (N_6865,N_5737,N_5406);
or U6866 (N_6866,N_5160,N_5331);
nor U6867 (N_6867,N_5901,N_5466);
and U6868 (N_6868,N_5737,N_5080);
xnor U6869 (N_6869,N_5227,N_5336);
or U6870 (N_6870,N_5043,N_5949);
and U6871 (N_6871,N_5621,N_5365);
nand U6872 (N_6872,N_5617,N_5449);
or U6873 (N_6873,N_5075,N_5702);
or U6874 (N_6874,N_5049,N_5132);
nand U6875 (N_6875,N_5851,N_5550);
or U6876 (N_6876,N_5818,N_5795);
and U6877 (N_6877,N_5977,N_5260);
xor U6878 (N_6878,N_5931,N_5704);
or U6879 (N_6879,N_5874,N_5305);
and U6880 (N_6880,N_5314,N_5929);
nand U6881 (N_6881,N_5200,N_5713);
nand U6882 (N_6882,N_5075,N_5899);
nand U6883 (N_6883,N_5943,N_5245);
and U6884 (N_6884,N_5666,N_5656);
nand U6885 (N_6885,N_5512,N_5430);
xor U6886 (N_6886,N_5888,N_5563);
or U6887 (N_6887,N_5495,N_5498);
xnor U6888 (N_6888,N_5208,N_5764);
nor U6889 (N_6889,N_5216,N_5499);
nor U6890 (N_6890,N_5397,N_5919);
or U6891 (N_6891,N_5671,N_5094);
nor U6892 (N_6892,N_5181,N_5645);
nand U6893 (N_6893,N_5640,N_5978);
nand U6894 (N_6894,N_5450,N_5632);
xnor U6895 (N_6895,N_5286,N_5593);
nor U6896 (N_6896,N_5948,N_5135);
or U6897 (N_6897,N_5342,N_5409);
nand U6898 (N_6898,N_5563,N_5156);
or U6899 (N_6899,N_5929,N_5779);
xor U6900 (N_6900,N_5624,N_5823);
or U6901 (N_6901,N_5760,N_5428);
or U6902 (N_6902,N_5949,N_5633);
nand U6903 (N_6903,N_5778,N_5106);
xnor U6904 (N_6904,N_5773,N_5199);
or U6905 (N_6905,N_5164,N_5339);
xnor U6906 (N_6906,N_5592,N_5004);
xor U6907 (N_6907,N_5040,N_5759);
nor U6908 (N_6908,N_5261,N_5986);
xnor U6909 (N_6909,N_5909,N_5066);
or U6910 (N_6910,N_5527,N_5199);
xnor U6911 (N_6911,N_5554,N_5055);
nor U6912 (N_6912,N_5199,N_5076);
xnor U6913 (N_6913,N_5840,N_5075);
xor U6914 (N_6914,N_5228,N_5140);
or U6915 (N_6915,N_5503,N_5011);
xor U6916 (N_6916,N_5067,N_5081);
nor U6917 (N_6917,N_5822,N_5341);
nand U6918 (N_6918,N_5195,N_5568);
nor U6919 (N_6919,N_5888,N_5653);
xor U6920 (N_6920,N_5720,N_5553);
nor U6921 (N_6921,N_5270,N_5187);
nand U6922 (N_6922,N_5153,N_5416);
and U6923 (N_6923,N_5257,N_5893);
nand U6924 (N_6924,N_5464,N_5488);
nand U6925 (N_6925,N_5952,N_5098);
and U6926 (N_6926,N_5078,N_5934);
or U6927 (N_6927,N_5948,N_5247);
or U6928 (N_6928,N_5566,N_5077);
xor U6929 (N_6929,N_5402,N_5286);
nor U6930 (N_6930,N_5481,N_5068);
or U6931 (N_6931,N_5394,N_5864);
xnor U6932 (N_6932,N_5824,N_5611);
nand U6933 (N_6933,N_5534,N_5484);
and U6934 (N_6934,N_5547,N_5260);
nor U6935 (N_6935,N_5314,N_5344);
and U6936 (N_6936,N_5945,N_5673);
and U6937 (N_6937,N_5172,N_5326);
nor U6938 (N_6938,N_5492,N_5917);
nand U6939 (N_6939,N_5249,N_5513);
or U6940 (N_6940,N_5767,N_5015);
or U6941 (N_6941,N_5835,N_5076);
and U6942 (N_6942,N_5283,N_5586);
nand U6943 (N_6943,N_5263,N_5386);
nand U6944 (N_6944,N_5690,N_5387);
xor U6945 (N_6945,N_5099,N_5301);
xnor U6946 (N_6946,N_5141,N_5537);
or U6947 (N_6947,N_5749,N_5576);
or U6948 (N_6948,N_5556,N_5339);
and U6949 (N_6949,N_5292,N_5794);
and U6950 (N_6950,N_5261,N_5735);
nor U6951 (N_6951,N_5766,N_5196);
and U6952 (N_6952,N_5950,N_5990);
nor U6953 (N_6953,N_5197,N_5667);
xor U6954 (N_6954,N_5509,N_5533);
or U6955 (N_6955,N_5146,N_5058);
nor U6956 (N_6956,N_5049,N_5973);
nor U6957 (N_6957,N_5647,N_5840);
nand U6958 (N_6958,N_5088,N_5802);
nand U6959 (N_6959,N_5279,N_5413);
or U6960 (N_6960,N_5140,N_5889);
xnor U6961 (N_6961,N_5089,N_5862);
and U6962 (N_6962,N_5397,N_5095);
xor U6963 (N_6963,N_5330,N_5643);
or U6964 (N_6964,N_5268,N_5904);
or U6965 (N_6965,N_5090,N_5667);
nand U6966 (N_6966,N_5888,N_5128);
xnor U6967 (N_6967,N_5680,N_5966);
nor U6968 (N_6968,N_5309,N_5980);
nor U6969 (N_6969,N_5908,N_5737);
xnor U6970 (N_6970,N_5355,N_5066);
xor U6971 (N_6971,N_5885,N_5650);
xor U6972 (N_6972,N_5701,N_5603);
nor U6973 (N_6973,N_5294,N_5184);
nand U6974 (N_6974,N_5262,N_5774);
xor U6975 (N_6975,N_5298,N_5994);
nor U6976 (N_6976,N_5710,N_5808);
and U6977 (N_6977,N_5776,N_5807);
or U6978 (N_6978,N_5168,N_5499);
xnor U6979 (N_6979,N_5129,N_5046);
or U6980 (N_6980,N_5169,N_5097);
xnor U6981 (N_6981,N_5700,N_5061);
nand U6982 (N_6982,N_5739,N_5516);
and U6983 (N_6983,N_5684,N_5892);
nand U6984 (N_6984,N_5756,N_5675);
nor U6985 (N_6985,N_5070,N_5512);
xor U6986 (N_6986,N_5395,N_5797);
nand U6987 (N_6987,N_5062,N_5760);
nor U6988 (N_6988,N_5555,N_5682);
nand U6989 (N_6989,N_5484,N_5935);
xnor U6990 (N_6990,N_5317,N_5040);
or U6991 (N_6991,N_5059,N_5587);
and U6992 (N_6992,N_5759,N_5611);
nand U6993 (N_6993,N_5894,N_5412);
or U6994 (N_6994,N_5557,N_5031);
and U6995 (N_6995,N_5531,N_5381);
nand U6996 (N_6996,N_5255,N_5102);
and U6997 (N_6997,N_5364,N_5885);
nand U6998 (N_6998,N_5048,N_5440);
nand U6999 (N_6999,N_5308,N_5762);
nand U7000 (N_7000,N_6727,N_6916);
nor U7001 (N_7001,N_6329,N_6277);
nand U7002 (N_7002,N_6926,N_6894);
or U7003 (N_7003,N_6480,N_6920);
nor U7004 (N_7004,N_6025,N_6590);
or U7005 (N_7005,N_6158,N_6192);
nand U7006 (N_7006,N_6600,N_6587);
nand U7007 (N_7007,N_6406,N_6165);
and U7008 (N_7008,N_6751,N_6606);
or U7009 (N_7009,N_6239,N_6998);
and U7010 (N_7010,N_6750,N_6911);
nor U7011 (N_7011,N_6665,N_6537);
xnor U7012 (N_7012,N_6095,N_6126);
nand U7013 (N_7013,N_6686,N_6097);
and U7014 (N_7014,N_6357,N_6919);
xnor U7015 (N_7015,N_6236,N_6993);
or U7016 (N_7016,N_6575,N_6623);
nand U7017 (N_7017,N_6147,N_6545);
nand U7018 (N_7018,N_6792,N_6736);
nor U7019 (N_7019,N_6882,N_6666);
xor U7020 (N_7020,N_6956,N_6457);
and U7021 (N_7021,N_6383,N_6682);
and U7022 (N_7022,N_6464,N_6586);
nand U7023 (N_7023,N_6511,N_6285);
nand U7024 (N_7024,N_6753,N_6468);
nor U7025 (N_7025,N_6034,N_6805);
or U7026 (N_7026,N_6044,N_6931);
xor U7027 (N_7027,N_6324,N_6243);
nor U7028 (N_7028,N_6513,N_6597);
nand U7029 (N_7029,N_6502,N_6759);
nor U7030 (N_7030,N_6426,N_6091);
or U7031 (N_7031,N_6704,N_6966);
nor U7032 (N_7032,N_6381,N_6626);
nand U7033 (N_7033,N_6201,N_6227);
nand U7034 (N_7034,N_6535,N_6720);
or U7035 (N_7035,N_6829,N_6046);
nand U7036 (N_7036,N_6083,N_6065);
or U7037 (N_7037,N_6059,N_6117);
nor U7038 (N_7038,N_6265,N_6644);
or U7039 (N_7039,N_6207,N_6278);
nand U7040 (N_7040,N_6144,N_6523);
and U7041 (N_7041,N_6768,N_6295);
nand U7042 (N_7042,N_6678,N_6865);
nor U7043 (N_7043,N_6087,N_6215);
xor U7044 (N_7044,N_6553,N_6818);
nand U7045 (N_7045,N_6416,N_6143);
or U7046 (N_7046,N_6456,N_6863);
nand U7047 (N_7047,N_6057,N_6868);
xnor U7048 (N_7048,N_6862,N_6465);
xnor U7049 (N_7049,N_6099,N_6249);
nand U7050 (N_7050,N_6790,N_6194);
nor U7051 (N_7051,N_6020,N_6155);
and U7052 (N_7052,N_6519,N_6417);
nand U7053 (N_7053,N_6237,N_6858);
and U7054 (N_7054,N_6145,N_6771);
nand U7055 (N_7055,N_6887,N_6128);
and U7056 (N_7056,N_6267,N_6199);
xnor U7057 (N_7057,N_6820,N_6892);
nor U7058 (N_7058,N_6177,N_6161);
nor U7059 (N_7059,N_6755,N_6262);
xnor U7060 (N_7060,N_6330,N_6967);
or U7061 (N_7061,N_6048,N_6156);
nor U7062 (N_7062,N_6189,N_6467);
and U7063 (N_7063,N_6387,N_6289);
xnor U7064 (N_7064,N_6430,N_6905);
nand U7065 (N_7065,N_6047,N_6717);
or U7066 (N_7066,N_6029,N_6801);
nor U7067 (N_7067,N_6670,N_6675);
nand U7068 (N_7068,N_6499,N_6404);
or U7069 (N_7069,N_6743,N_6784);
or U7070 (N_7070,N_6811,N_6127);
xor U7071 (N_7071,N_6347,N_6006);
xnor U7072 (N_7072,N_6725,N_6138);
and U7073 (N_7073,N_6737,N_6162);
and U7074 (N_7074,N_6847,N_6134);
and U7075 (N_7075,N_6974,N_6546);
nor U7076 (N_7076,N_6504,N_6853);
and U7077 (N_7077,N_6851,N_6536);
xor U7078 (N_7078,N_6420,N_6185);
and U7079 (N_7079,N_6779,N_6995);
or U7080 (N_7080,N_6634,N_6925);
or U7081 (N_7081,N_6409,N_6361);
nor U7082 (N_7082,N_6191,N_6290);
xnor U7083 (N_7083,N_6166,N_6242);
nand U7084 (N_7084,N_6184,N_6170);
nand U7085 (N_7085,N_6832,N_6338);
and U7086 (N_7086,N_6870,N_6578);
xor U7087 (N_7087,N_6867,N_6848);
xnor U7088 (N_7088,N_6284,N_6757);
or U7089 (N_7089,N_6209,N_6819);
or U7090 (N_7090,N_6306,N_6729);
and U7091 (N_7091,N_6945,N_6951);
nor U7092 (N_7092,N_6241,N_6496);
or U7093 (N_7093,N_6451,N_6258);
nand U7094 (N_7094,N_6061,N_6680);
and U7095 (N_7095,N_6726,N_6076);
nor U7096 (N_7096,N_6445,N_6049);
xor U7097 (N_7097,N_6923,N_6021);
xor U7098 (N_7098,N_6385,N_6313);
or U7099 (N_7099,N_6431,N_6749);
nor U7100 (N_7100,N_6261,N_6762);
nand U7101 (N_7101,N_6875,N_6981);
xor U7102 (N_7102,N_6159,N_6078);
and U7103 (N_7103,N_6731,N_6062);
xor U7104 (N_7104,N_6529,N_6478);
nor U7105 (N_7105,N_6410,N_6983);
nand U7106 (N_7106,N_6558,N_6681);
nor U7107 (N_7107,N_6937,N_6141);
or U7108 (N_7108,N_6205,N_6621);
and U7109 (N_7109,N_6474,N_6627);
nand U7110 (N_7110,N_6498,N_6343);
and U7111 (N_7111,N_6589,N_6092);
xor U7112 (N_7112,N_6171,N_6527);
nor U7113 (N_7113,N_6673,N_6948);
nor U7114 (N_7114,N_6799,N_6655);
xnor U7115 (N_7115,N_6024,N_6425);
nor U7116 (N_7116,N_6372,N_6696);
nor U7117 (N_7117,N_6494,N_6386);
nor U7118 (N_7118,N_6257,N_6331);
nor U7119 (N_7119,N_6100,N_6524);
or U7120 (N_7120,N_6233,N_6287);
xnor U7121 (N_7121,N_6533,N_6893);
nor U7122 (N_7122,N_6714,N_6598);
xnor U7123 (N_7123,N_6214,N_6517);
or U7124 (N_7124,N_6946,N_6958);
or U7125 (N_7125,N_6119,N_6971);
and U7126 (N_7126,N_6777,N_6809);
xor U7127 (N_7127,N_6924,N_6667);
xor U7128 (N_7128,N_6448,N_6140);
and U7129 (N_7129,N_6580,N_6392);
xor U7130 (N_7130,N_6637,N_6460);
xnor U7131 (N_7131,N_6556,N_6316);
and U7132 (N_7132,N_6113,N_6953);
or U7133 (N_7133,N_6884,N_6602);
nand U7134 (N_7134,N_6897,N_6719);
xnor U7135 (N_7135,N_6073,N_6964);
nor U7136 (N_7136,N_6312,N_6611);
nand U7137 (N_7137,N_6407,N_6272);
and U7138 (N_7138,N_6608,N_6573);
and U7139 (N_7139,N_6568,N_6668);
nor U7140 (N_7140,N_6561,N_6772);
nand U7141 (N_7141,N_6785,N_6074);
and U7142 (N_7142,N_6326,N_6336);
xnor U7143 (N_7143,N_6217,N_6271);
and U7144 (N_7144,N_6534,N_6601);
and U7145 (N_7145,N_6222,N_6856);
or U7146 (N_7146,N_6268,N_6797);
nor U7147 (N_7147,N_6154,N_6173);
or U7148 (N_7148,N_6012,N_6936);
nor U7149 (N_7149,N_6015,N_6514);
or U7150 (N_7150,N_6228,N_6403);
and U7151 (N_7151,N_6137,N_6056);
nand U7152 (N_7152,N_6365,N_6512);
nand U7153 (N_7153,N_6572,N_6695);
xor U7154 (N_7154,N_6179,N_6669);
nor U7155 (N_7155,N_6987,N_6742);
nand U7156 (N_7156,N_6356,N_6636);
nand U7157 (N_7157,N_6240,N_6320);
nand U7158 (N_7158,N_6551,N_6421);
or U7159 (N_7159,N_6888,N_6297);
nor U7160 (N_7160,N_6007,N_6857);
nand U7161 (N_7161,N_6291,N_6370);
and U7162 (N_7162,N_6193,N_6618);
nor U7163 (N_7163,N_6789,N_6615);
nor U7164 (N_7164,N_6461,N_6234);
or U7165 (N_7165,N_6830,N_6827);
nor U7166 (N_7166,N_6470,N_6874);
xor U7167 (N_7167,N_6160,N_6813);
and U7168 (N_7168,N_6307,N_6518);
xnor U7169 (N_7169,N_6732,N_6849);
nand U7170 (N_7170,N_6939,N_6379);
nand U7171 (N_7171,N_6027,N_6999);
or U7172 (N_7172,N_6622,N_6965);
xor U7173 (N_7173,N_6219,N_6501);
and U7174 (N_7174,N_6142,N_6439);
nor U7175 (N_7175,N_6877,N_6042);
nand U7176 (N_7176,N_6549,N_6133);
xor U7177 (N_7177,N_6656,N_6345);
xor U7178 (N_7178,N_6836,N_6283);
or U7179 (N_7179,N_6394,N_6715);
xnor U7180 (N_7180,N_6664,N_6082);
xnor U7181 (N_7181,N_6315,N_6642);
and U7182 (N_7182,N_6839,N_6515);
nand U7183 (N_7183,N_6860,N_6859);
nand U7184 (N_7184,N_6220,N_6067);
xnor U7185 (N_7185,N_6908,N_6794);
nor U7186 (N_7186,N_6148,N_6226);
or U7187 (N_7187,N_6593,N_6619);
or U7188 (N_7188,N_6703,N_6775);
or U7189 (N_7189,N_6235,N_6840);
xnor U7190 (N_7190,N_6175,N_6210);
or U7191 (N_7191,N_6221,N_6299);
nor U7192 (N_7192,N_6730,N_6308);
xor U7193 (N_7193,N_6835,N_6872);
or U7194 (N_7194,N_6344,N_6918);
or U7195 (N_7195,N_6699,N_6541);
nor U7196 (N_7196,N_6202,N_6053);
and U7197 (N_7197,N_6068,N_6910);
xnor U7198 (N_7198,N_6052,N_6722);
nand U7199 (N_7199,N_6850,N_6321);
and U7200 (N_7200,N_6774,N_6756);
nand U7201 (N_7201,N_6604,N_6563);
xnor U7202 (N_7202,N_6505,N_6866);
nand U7203 (N_7203,N_6351,N_6674);
nor U7204 (N_7204,N_6585,N_6683);
or U7205 (N_7205,N_6253,N_6274);
xor U7206 (N_7206,N_6028,N_6429);
nor U7207 (N_7207,N_6982,N_6060);
and U7208 (N_7208,N_6869,N_6400);
nor U7209 (N_7209,N_6491,N_6218);
and U7210 (N_7210,N_6019,N_6001);
nor U7211 (N_7211,N_6571,N_6167);
and U7212 (N_7212,N_6102,N_6023);
and U7213 (N_7213,N_6190,N_6639);
and U7214 (N_7214,N_6441,N_6728);
nand U7215 (N_7215,N_6108,N_6116);
nor U7216 (N_7216,N_6466,N_6488);
nor U7217 (N_7217,N_6933,N_6079);
nor U7218 (N_7218,N_6773,N_6990);
nor U7219 (N_7219,N_6935,N_6913);
xor U7220 (N_7220,N_6603,N_6943);
xor U7221 (N_7221,N_6748,N_6638);
and U7222 (N_7222,N_6340,N_6917);
xor U7223 (N_7223,N_6776,N_6952);
and U7224 (N_7224,N_6438,N_6374);
nor U7225 (N_7225,N_6927,N_6906);
xnor U7226 (N_7226,N_6596,N_6463);
or U7227 (N_7227,N_6831,N_6876);
and U7228 (N_7228,N_6098,N_6823);
nor U7229 (N_7229,N_6758,N_6035);
or U7230 (N_7230,N_6708,N_6591);
nor U7231 (N_7231,N_6497,N_6399);
and U7232 (N_7232,N_6994,N_6500);
nor U7233 (N_7233,N_6168,N_6413);
nand U7234 (N_7234,N_6803,N_6816);
nand U7235 (N_7235,N_6396,N_6435);
nor U7236 (N_7236,N_6928,N_6146);
xor U7237 (N_7237,N_6689,N_6090);
and U7238 (N_7238,N_6979,N_6390);
and U7239 (N_7239,N_6206,N_6845);
nor U7240 (N_7240,N_6938,N_6954);
nand U7241 (N_7241,N_6716,N_6462);
nand U7242 (N_7242,N_6968,N_6802);
or U7243 (N_7243,N_6934,N_6051);
nand U7244 (N_7244,N_6106,N_6486);
xor U7245 (N_7245,N_6036,N_6010);
xnor U7246 (N_7246,N_6349,N_6705);
nor U7247 (N_7247,N_6609,N_6692);
nand U7248 (N_7248,N_6211,N_6713);
nand U7249 (N_7249,N_6369,N_6122);
and U7250 (N_7250,N_6280,N_6635);
or U7251 (N_7251,N_6436,N_6094);
nor U7252 (N_7252,N_6475,N_6625);
and U7253 (N_7253,N_6879,N_6111);
nor U7254 (N_7254,N_6229,N_6570);
or U7255 (N_7255,N_6332,N_6806);
or U7256 (N_7256,N_6795,N_6972);
xnor U7257 (N_7257,N_6245,N_6389);
xor U7258 (N_7258,N_6139,N_6889);
xor U7259 (N_7259,N_6969,N_6016);
nor U7260 (N_7260,N_6481,N_6903);
nor U7261 (N_7261,N_6018,N_6341);
xor U7262 (N_7262,N_6907,N_6531);
or U7263 (N_7263,N_6780,N_6296);
and U7264 (N_7264,N_6398,N_6781);
nand U7265 (N_7265,N_6855,N_6616);
xnor U7266 (N_7266,N_6004,N_6579);
nand U7267 (N_7267,N_6030,N_6382);
nor U7268 (N_7268,N_6922,N_6594);
and U7269 (N_7269,N_6411,N_6084);
or U7270 (N_7270,N_6255,N_6124);
xnor U7271 (N_7271,N_6914,N_6883);
or U7272 (N_7272,N_6150,N_6458);
nor U7273 (N_7273,N_6443,N_6476);
and U7274 (N_7274,N_6520,N_6401);
and U7275 (N_7275,N_6899,N_6783);
or U7276 (N_7276,N_6747,N_6101);
nor U7277 (N_7277,N_6352,N_6477);
xnor U7278 (N_7278,N_6978,N_6550);
or U7279 (N_7279,N_6640,N_6033);
nand U7280 (N_7280,N_6086,N_6017);
xor U7281 (N_7281,N_6450,N_6614);
or U7282 (N_7282,N_6292,N_6157);
xor U7283 (N_7283,N_6649,N_6418);
nor U7284 (N_7284,N_6471,N_6348);
nor U7285 (N_7285,N_6940,N_6495);
and U7286 (N_7286,N_6328,N_6373);
nand U7287 (N_7287,N_6564,N_6125);
xor U7288 (N_7288,N_6960,N_6852);
nor U7289 (N_7289,N_6013,N_6377);
nand U7290 (N_7290,N_6317,N_6688);
nand U7291 (N_7291,N_6454,N_6055);
nor U7292 (N_7292,N_6815,N_6066);
nand U7293 (N_7293,N_6810,N_6424);
or U7294 (N_7294,N_6230,N_6539);
nor U7295 (N_7295,N_6522,N_6962);
nand U7296 (N_7296,N_6828,N_6198);
xor U7297 (N_7297,N_6181,N_6654);
xnor U7298 (N_7298,N_6281,N_6698);
or U7299 (N_7299,N_6764,N_6694);
nor U7300 (N_7300,N_6131,N_6197);
xor U7301 (N_7301,N_6959,N_6921);
nor U7302 (N_7302,N_6547,N_6043);
nor U7303 (N_7303,N_6485,N_6391);
nor U7304 (N_7304,N_6452,N_6873);
nor U7305 (N_7305,N_6453,N_6355);
nand U7306 (N_7306,N_6507,N_6358);
and U7307 (N_7307,N_6322,N_6367);
nor U7308 (N_7308,N_6294,N_6212);
nor U7309 (N_7309,N_6402,N_6264);
nor U7310 (N_7310,N_6256,N_6364);
nand U7311 (N_7311,N_6112,N_6796);
nand U7312 (N_7312,N_6200,N_6005);
and U7313 (N_7313,N_6647,N_6648);
or U7314 (N_7314,N_6592,N_6260);
nand U7315 (N_7315,N_6447,N_6878);
or U7316 (N_7316,N_6300,N_6629);
and U7317 (N_7317,N_6949,N_6444);
and U7318 (N_7318,N_6003,N_6031);
or U7319 (N_7319,N_6318,N_6807);
or U7320 (N_7320,N_6977,N_6808);
and U7321 (N_7321,N_6581,N_6375);
and U7322 (N_7322,N_6405,N_6760);
or U7323 (N_7323,N_6787,N_6992);
and U7324 (N_7324,N_6895,N_6838);
nor U7325 (N_7325,N_6309,N_6479);
and U7326 (N_7326,N_6216,N_6130);
xnor U7327 (N_7327,N_6740,N_6991);
or U7328 (N_7328,N_6380,N_6252);
nor U7329 (N_7329,N_6415,N_6788);
nand U7330 (N_7330,N_6103,N_6449);
or U7331 (N_7331,N_6339,N_6980);
nor U7332 (N_7332,N_6660,N_6037);
nand U7333 (N_7333,N_6251,N_6069);
nor U7334 (N_7334,N_6187,N_6250);
or U7335 (N_7335,N_6890,N_6302);
and U7336 (N_7336,N_6841,N_6039);
xnor U7337 (N_7337,N_6080,N_6123);
xnor U7338 (N_7338,N_6651,N_6746);
nor U7339 (N_7339,N_6081,N_6718);
or U7340 (N_7340,N_6770,N_6528);
or U7341 (N_7341,N_6040,N_6473);
and U7342 (N_7342,N_6008,N_6266);
xor U7343 (N_7343,N_6428,N_6842);
xnor U7344 (N_7344,N_6089,N_6293);
nor U7345 (N_7345,N_6490,N_6607);
or U7346 (N_7346,N_6371,N_6038);
xnor U7347 (N_7347,N_6697,N_6325);
and U7348 (N_7348,N_6393,N_6822);
and U7349 (N_7349,N_6837,N_6767);
nor U7350 (N_7350,N_6153,N_6950);
and U7351 (N_7351,N_6136,N_6532);
nor U7352 (N_7352,N_6186,N_6885);
xor U7353 (N_7353,N_6483,N_6432);
xnor U7354 (N_7354,N_6632,N_6800);
and U7355 (N_7355,N_6555,N_6833);
or U7356 (N_7356,N_6213,N_6645);
or U7357 (N_7357,N_6576,N_6440);
and U7358 (N_7358,N_6691,N_6246);
xnor U7359 (N_7359,N_6433,N_6880);
xnor U7360 (N_7360,N_6419,N_6963);
and U7361 (N_7361,N_6584,N_6273);
xnor U7362 (N_7362,N_6864,N_6088);
or U7363 (N_7363,N_6196,N_6304);
and U7364 (N_7364,N_6985,N_6957);
nor U7365 (N_7365,N_6814,N_6070);
nand U7366 (N_7366,N_6151,N_6854);
nand U7367 (N_7367,N_6804,N_6172);
nor U7368 (N_7368,N_6350,N_6254);
xnor U7369 (N_7369,N_6085,N_6305);
nor U7370 (N_7370,N_6687,N_6763);
xnor U7371 (N_7371,N_6509,N_6798);
and U7372 (N_7372,N_6929,N_6702);
and U7373 (N_7373,N_6050,N_6739);
or U7374 (N_7374,N_6263,N_6359);
or U7375 (N_7375,N_6548,N_6817);
and U7376 (N_7376,N_6932,N_6077);
xor U7377 (N_7377,N_6752,N_6628);
xor U7378 (N_7378,N_6354,N_6861);
xnor U7379 (N_7379,N_6169,N_6650);
nor U7380 (N_7380,N_6427,N_6489);
nand U7381 (N_7381,N_6135,N_6121);
xnor U7382 (N_7382,N_6279,N_6902);
and U7383 (N_7383,N_6973,N_6286);
or U7384 (N_7384,N_6521,N_6824);
nor U7385 (N_7385,N_6685,N_6032);
nor U7386 (N_7386,N_6583,N_6275);
or U7387 (N_7387,N_6516,N_6118);
nand U7388 (N_7388,N_6132,N_6530);
and U7389 (N_7389,N_6323,N_6333);
xnor U7390 (N_7390,N_6723,N_6064);
and U7391 (N_7391,N_6011,N_6000);
and U7392 (N_7392,N_6653,N_6912);
and U7393 (N_7393,N_6552,N_6093);
and U7394 (N_7394,N_6363,N_6671);
xnor U7395 (N_7395,N_6301,N_6569);
or U7396 (N_7396,N_6314,N_6303);
nor U7397 (N_7397,N_6026,N_6542);
nor U7398 (N_7398,N_6009,N_6577);
or U7399 (N_7399,N_6909,N_6395);
nand U7400 (N_7400,N_6582,N_6412);
nor U7401 (N_7401,N_6605,N_6821);
or U7402 (N_7402,N_6672,N_6744);
xor U7403 (N_7403,N_6540,N_6559);
nand U7404 (N_7404,N_6711,N_6298);
xor U7405 (N_7405,N_6288,N_6701);
or U7406 (N_7406,N_6188,N_6225);
xnor U7407 (N_7407,N_6506,N_6754);
xor U7408 (N_7408,N_6469,N_6707);
nor U7409 (N_7409,N_6276,N_6346);
and U7410 (N_7410,N_6204,N_6662);
nand U7411 (N_7411,N_6896,N_6846);
or U7412 (N_7412,N_6741,N_6129);
nor U7413 (N_7413,N_6944,N_6712);
nor U7414 (N_7414,N_6989,N_6791);
nor U7415 (N_7415,N_6930,N_6310);
nand U7416 (N_7416,N_6658,N_6996);
or U7417 (N_7417,N_6182,N_6544);
nor U7418 (N_7418,N_6208,N_6376);
nor U7419 (N_7419,N_6643,N_6360);
nand U7420 (N_7420,N_6915,N_6734);
nand U7421 (N_7421,N_6384,N_6075);
xor U7422 (N_7422,N_6397,N_6163);
nand U7423 (N_7423,N_6492,N_6612);
nor U7424 (N_7424,N_6526,N_6901);
xor U7425 (N_7425,N_6633,N_6180);
and U7426 (N_7426,N_6109,N_6107);
nor U7427 (N_7427,N_6472,N_6721);
nand U7428 (N_7428,N_6975,N_6041);
nor U7429 (N_7429,N_6482,N_6248);
or U7430 (N_7430,N_6567,N_6149);
nor U7431 (N_7431,N_6114,N_6022);
nand U7432 (N_7432,N_6709,N_6437);
nor U7433 (N_7433,N_6110,N_6613);
nor U7434 (N_7434,N_6105,N_6423);
nand U7435 (N_7435,N_6947,N_6826);
or U7436 (N_7436,N_6566,N_6319);
nand U7437 (N_7437,N_6484,N_6388);
xor U7438 (N_7438,N_6588,N_6766);
nand U7439 (N_7439,N_6843,N_6898);
nand U7440 (N_7440,N_6414,N_6652);
xor U7441 (N_7441,N_6231,N_6942);
or U7442 (N_7442,N_6844,N_6232);
nand U7443 (N_7443,N_6422,N_6891);
nor U7444 (N_7444,N_6624,N_6631);
nand U7445 (N_7445,N_6493,N_6014);
nand U7446 (N_7446,N_6508,N_6164);
or U7447 (N_7447,N_6152,N_6045);
or U7448 (N_7448,N_6976,N_6054);
nor U7449 (N_7449,N_6574,N_6071);
nor U7450 (N_7450,N_6178,N_6562);
nor U7451 (N_7451,N_6543,N_6557);
nand U7452 (N_7452,N_6247,N_6986);
nand U7453 (N_7453,N_6334,N_6311);
nor U7454 (N_7454,N_6335,N_6104);
xnor U7455 (N_7455,N_6565,N_6176);
nand U7456 (N_7456,N_6684,N_6679);
xnor U7457 (N_7457,N_6259,N_6282);
nand U7458 (N_7458,N_6058,N_6970);
or U7459 (N_7459,N_6442,N_6337);
nand U7460 (N_7460,N_6342,N_6676);
nand U7461 (N_7461,N_6238,N_6778);
nor U7462 (N_7462,N_6244,N_6735);
nand U7463 (N_7463,N_6904,N_6269);
and U7464 (N_7464,N_6812,N_6063);
or U7465 (N_7465,N_6353,N_6002);
xnor U7466 (N_7466,N_6997,N_6620);
and U7467 (N_7467,N_6661,N_6503);
and U7468 (N_7468,N_6120,N_6677);
or U7469 (N_7469,N_6710,N_6174);
and U7470 (N_7470,N_6941,N_6362);
and U7471 (N_7471,N_6738,N_6327);
nor U7472 (N_7472,N_6881,N_6871);
xnor U7473 (N_7473,N_6641,N_6487);
nand U7474 (N_7474,N_6657,N_6834);
nor U7475 (N_7475,N_6700,N_6825);
nor U7476 (N_7476,N_6368,N_6724);
nor U7477 (N_7477,N_6096,N_6733);
xnor U7478 (N_7478,N_6203,N_6599);
xnor U7479 (N_7479,N_6525,N_6610);
nand U7480 (N_7480,N_6538,N_6786);
nand U7481 (N_7481,N_6455,N_6984);
and U7482 (N_7482,N_6595,N_6510);
or U7483 (N_7483,N_6769,N_6646);
xnor U7484 (N_7484,N_6224,N_6886);
and U7485 (N_7485,N_6378,N_6745);
and U7486 (N_7486,N_6782,N_6366);
xnor U7487 (N_7487,N_6630,N_6223);
or U7488 (N_7488,N_6554,N_6706);
nand U7489 (N_7489,N_6183,N_6195);
or U7490 (N_7490,N_6955,N_6560);
nand U7491 (N_7491,N_6663,N_6459);
xor U7492 (N_7492,N_6988,N_6900);
or U7493 (N_7493,N_6446,N_6617);
nand U7494 (N_7494,N_6690,N_6270);
xor U7495 (N_7495,N_6408,N_6659);
or U7496 (N_7496,N_6765,N_6072);
xor U7497 (N_7497,N_6115,N_6793);
nand U7498 (N_7498,N_6434,N_6761);
nor U7499 (N_7499,N_6961,N_6693);
nand U7500 (N_7500,N_6151,N_6968);
nand U7501 (N_7501,N_6292,N_6323);
nand U7502 (N_7502,N_6397,N_6954);
or U7503 (N_7503,N_6606,N_6192);
and U7504 (N_7504,N_6496,N_6438);
and U7505 (N_7505,N_6148,N_6003);
xor U7506 (N_7506,N_6874,N_6509);
nor U7507 (N_7507,N_6752,N_6615);
nand U7508 (N_7508,N_6274,N_6738);
xor U7509 (N_7509,N_6741,N_6458);
and U7510 (N_7510,N_6328,N_6926);
nor U7511 (N_7511,N_6777,N_6274);
xnor U7512 (N_7512,N_6434,N_6149);
or U7513 (N_7513,N_6568,N_6639);
and U7514 (N_7514,N_6278,N_6564);
xnor U7515 (N_7515,N_6753,N_6781);
nor U7516 (N_7516,N_6826,N_6812);
xor U7517 (N_7517,N_6079,N_6592);
nor U7518 (N_7518,N_6964,N_6716);
nor U7519 (N_7519,N_6651,N_6668);
or U7520 (N_7520,N_6896,N_6384);
or U7521 (N_7521,N_6125,N_6855);
xnor U7522 (N_7522,N_6201,N_6690);
xnor U7523 (N_7523,N_6133,N_6883);
and U7524 (N_7524,N_6487,N_6822);
or U7525 (N_7525,N_6261,N_6485);
and U7526 (N_7526,N_6434,N_6290);
xor U7527 (N_7527,N_6074,N_6759);
nor U7528 (N_7528,N_6287,N_6255);
nand U7529 (N_7529,N_6644,N_6013);
and U7530 (N_7530,N_6260,N_6168);
nand U7531 (N_7531,N_6021,N_6332);
nand U7532 (N_7532,N_6307,N_6244);
nand U7533 (N_7533,N_6110,N_6938);
nor U7534 (N_7534,N_6802,N_6147);
nand U7535 (N_7535,N_6615,N_6895);
nor U7536 (N_7536,N_6356,N_6830);
nand U7537 (N_7537,N_6592,N_6962);
nand U7538 (N_7538,N_6520,N_6595);
nor U7539 (N_7539,N_6966,N_6705);
xnor U7540 (N_7540,N_6407,N_6853);
or U7541 (N_7541,N_6588,N_6439);
or U7542 (N_7542,N_6061,N_6711);
or U7543 (N_7543,N_6099,N_6369);
xnor U7544 (N_7544,N_6258,N_6414);
nor U7545 (N_7545,N_6955,N_6566);
nor U7546 (N_7546,N_6079,N_6547);
or U7547 (N_7547,N_6342,N_6248);
nand U7548 (N_7548,N_6979,N_6046);
or U7549 (N_7549,N_6066,N_6537);
nand U7550 (N_7550,N_6858,N_6844);
nand U7551 (N_7551,N_6180,N_6140);
nand U7552 (N_7552,N_6415,N_6548);
nor U7553 (N_7553,N_6447,N_6581);
and U7554 (N_7554,N_6295,N_6077);
or U7555 (N_7555,N_6415,N_6816);
and U7556 (N_7556,N_6272,N_6147);
nor U7557 (N_7557,N_6831,N_6248);
xor U7558 (N_7558,N_6161,N_6955);
nor U7559 (N_7559,N_6358,N_6338);
nor U7560 (N_7560,N_6981,N_6916);
xnor U7561 (N_7561,N_6425,N_6286);
nand U7562 (N_7562,N_6366,N_6564);
nor U7563 (N_7563,N_6221,N_6974);
or U7564 (N_7564,N_6885,N_6786);
and U7565 (N_7565,N_6620,N_6626);
xor U7566 (N_7566,N_6589,N_6677);
nor U7567 (N_7567,N_6420,N_6843);
nand U7568 (N_7568,N_6767,N_6730);
or U7569 (N_7569,N_6674,N_6884);
and U7570 (N_7570,N_6906,N_6041);
nor U7571 (N_7571,N_6275,N_6744);
xor U7572 (N_7572,N_6381,N_6424);
or U7573 (N_7573,N_6063,N_6115);
nor U7574 (N_7574,N_6791,N_6546);
xor U7575 (N_7575,N_6532,N_6139);
nor U7576 (N_7576,N_6675,N_6678);
nand U7577 (N_7577,N_6081,N_6519);
and U7578 (N_7578,N_6650,N_6048);
or U7579 (N_7579,N_6210,N_6589);
nor U7580 (N_7580,N_6569,N_6618);
nand U7581 (N_7581,N_6132,N_6996);
nor U7582 (N_7582,N_6473,N_6078);
xnor U7583 (N_7583,N_6159,N_6093);
and U7584 (N_7584,N_6476,N_6469);
and U7585 (N_7585,N_6409,N_6168);
and U7586 (N_7586,N_6495,N_6871);
and U7587 (N_7587,N_6820,N_6205);
xnor U7588 (N_7588,N_6266,N_6346);
xor U7589 (N_7589,N_6285,N_6617);
or U7590 (N_7590,N_6247,N_6719);
and U7591 (N_7591,N_6536,N_6730);
xor U7592 (N_7592,N_6426,N_6305);
xnor U7593 (N_7593,N_6661,N_6668);
nand U7594 (N_7594,N_6556,N_6958);
nand U7595 (N_7595,N_6085,N_6222);
and U7596 (N_7596,N_6288,N_6763);
and U7597 (N_7597,N_6226,N_6416);
xnor U7598 (N_7598,N_6274,N_6573);
nor U7599 (N_7599,N_6563,N_6048);
or U7600 (N_7600,N_6349,N_6039);
nor U7601 (N_7601,N_6377,N_6482);
nand U7602 (N_7602,N_6647,N_6976);
xnor U7603 (N_7603,N_6081,N_6805);
xor U7604 (N_7604,N_6570,N_6169);
or U7605 (N_7605,N_6187,N_6984);
nand U7606 (N_7606,N_6899,N_6622);
or U7607 (N_7607,N_6393,N_6177);
or U7608 (N_7608,N_6828,N_6431);
nor U7609 (N_7609,N_6808,N_6014);
nor U7610 (N_7610,N_6180,N_6201);
nor U7611 (N_7611,N_6790,N_6621);
nor U7612 (N_7612,N_6048,N_6658);
or U7613 (N_7613,N_6688,N_6796);
xnor U7614 (N_7614,N_6337,N_6850);
xnor U7615 (N_7615,N_6433,N_6923);
xnor U7616 (N_7616,N_6570,N_6618);
and U7617 (N_7617,N_6224,N_6549);
xor U7618 (N_7618,N_6128,N_6682);
and U7619 (N_7619,N_6206,N_6043);
and U7620 (N_7620,N_6059,N_6017);
and U7621 (N_7621,N_6131,N_6656);
xor U7622 (N_7622,N_6447,N_6685);
nand U7623 (N_7623,N_6448,N_6532);
xor U7624 (N_7624,N_6039,N_6091);
nor U7625 (N_7625,N_6524,N_6173);
and U7626 (N_7626,N_6625,N_6097);
xnor U7627 (N_7627,N_6310,N_6085);
xor U7628 (N_7628,N_6342,N_6977);
nor U7629 (N_7629,N_6598,N_6554);
and U7630 (N_7630,N_6491,N_6361);
nor U7631 (N_7631,N_6810,N_6722);
and U7632 (N_7632,N_6459,N_6834);
xor U7633 (N_7633,N_6732,N_6413);
nand U7634 (N_7634,N_6836,N_6460);
nor U7635 (N_7635,N_6866,N_6714);
nor U7636 (N_7636,N_6265,N_6564);
nand U7637 (N_7637,N_6363,N_6438);
or U7638 (N_7638,N_6725,N_6600);
nor U7639 (N_7639,N_6394,N_6112);
and U7640 (N_7640,N_6594,N_6629);
nand U7641 (N_7641,N_6060,N_6336);
nand U7642 (N_7642,N_6434,N_6810);
nor U7643 (N_7643,N_6836,N_6473);
or U7644 (N_7644,N_6732,N_6966);
nor U7645 (N_7645,N_6124,N_6523);
nor U7646 (N_7646,N_6544,N_6629);
nand U7647 (N_7647,N_6641,N_6133);
nor U7648 (N_7648,N_6835,N_6690);
and U7649 (N_7649,N_6832,N_6993);
and U7650 (N_7650,N_6938,N_6244);
nor U7651 (N_7651,N_6821,N_6967);
nand U7652 (N_7652,N_6643,N_6083);
and U7653 (N_7653,N_6942,N_6494);
and U7654 (N_7654,N_6550,N_6328);
and U7655 (N_7655,N_6260,N_6082);
or U7656 (N_7656,N_6400,N_6352);
and U7657 (N_7657,N_6890,N_6553);
nor U7658 (N_7658,N_6988,N_6910);
nand U7659 (N_7659,N_6401,N_6450);
xor U7660 (N_7660,N_6144,N_6147);
nor U7661 (N_7661,N_6900,N_6070);
or U7662 (N_7662,N_6643,N_6133);
nand U7663 (N_7663,N_6042,N_6201);
or U7664 (N_7664,N_6737,N_6449);
xor U7665 (N_7665,N_6078,N_6444);
xnor U7666 (N_7666,N_6757,N_6477);
nand U7667 (N_7667,N_6732,N_6101);
or U7668 (N_7668,N_6817,N_6553);
and U7669 (N_7669,N_6900,N_6143);
or U7670 (N_7670,N_6006,N_6560);
xor U7671 (N_7671,N_6278,N_6961);
xnor U7672 (N_7672,N_6068,N_6405);
or U7673 (N_7673,N_6602,N_6933);
and U7674 (N_7674,N_6815,N_6131);
or U7675 (N_7675,N_6890,N_6862);
xor U7676 (N_7676,N_6701,N_6900);
xnor U7677 (N_7677,N_6150,N_6836);
xor U7678 (N_7678,N_6630,N_6509);
xnor U7679 (N_7679,N_6120,N_6479);
nand U7680 (N_7680,N_6907,N_6645);
or U7681 (N_7681,N_6323,N_6679);
or U7682 (N_7682,N_6211,N_6028);
and U7683 (N_7683,N_6637,N_6170);
nand U7684 (N_7684,N_6330,N_6028);
nand U7685 (N_7685,N_6835,N_6614);
nor U7686 (N_7686,N_6573,N_6530);
nand U7687 (N_7687,N_6350,N_6798);
nor U7688 (N_7688,N_6250,N_6492);
xnor U7689 (N_7689,N_6757,N_6221);
nor U7690 (N_7690,N_6551,N_6522);
or U7691 (N_7691,N_6426,N_6075);
nand U7692 (N_7692,N_6841,N_6042);
xnor U7693 (N_7693,N_6864,N_6113);
nor U7694 (N_7694,N_6661,N_6434);
and U7695 (N_7695,N_6494,N_6304);
or U7696 (N_7696,N_6325,N_6757);
nand U7697 (N_7697,N_6338,N_6604);
xor U7698 (N_7698,N_6620,N_6354);
nand U7699 (N_7699,N_6210,N_6078);
and U7700 (N_7700,N_6558,N_6519);
nand U7701 (N_7701,N_6912,N_6079);
or U7702 (N_7702,N_6668,N_6551);
xor U7703 (N_7703,N_6082,N_6949);
and U7704 (N_7704,N_6618,N_6012);
nor U7705 (N_7705,N_6085,N_6238);
nor U7706 (N_7706,N_6994,N_6444);
or U7707 (N_7707,N_6831,N_6250);
or U7708 (N_7708,N_6559,N_6077);
nor U7709 (N_7709,N_6959,N_6976);
nor U7710 (N_7710,N_6905,N_6264);
and U7711 (N_7711,N_6981,N_6515);
nor U7712 (N_7712,N_6552,N_6920);
or U7713 (N_7713,N_6590,N_6035);
or U7714 (N_7714,N_6141,N_6279);
or U7715 (N_7715,N_6891,N_6290);
xor U7716 (N_7716,N_6099,N_6738);
xnor U7717 (N_7717,N_6482,N_6968);
nor U7718 (N_7718,N_6188,N_6868);
nor U7719 (N_7719,N_6310,N_6866);
nand U7720 (N_7720,N_6321,N_6236);
or U7721 (N_7721,N_6341,N_6858);
and U7722 (N_7722,N_6805,N_6672);
nand U7723 (N_7723,N_6029,N_6770);
nand U7724 (N_7724,N_6986,N_6814);
and U7725 (N_7725,N_6188,N_6316);
and U7726 (N_7726,N_6583,N_6286);
and U7727 (N_7727,N_6637,N_6809);
nand U7728 (N_7728,N_6263,N_6041);
or U7729 (N_7729,N_6141,N_6595);
and U7730 (N_7730,N_6045,N_6762);
nand U7731 (N_7731,N_6601,N_6597);
and U7732 (N_7732,N_6251,N_6494);
xnor U7733 (N_7733,N_6544,N_6219);
nand U7734 (N_7734,N_6489,N_6683);
or U7735 (N_7735,N_6092,N_6128);
and U7736 (N_7736,N_6584,N_6474);
nor U7737 (N_7737,N_6098,N_6924);
or U7738 (N_7738,N_6105,N_6402);
and U7739 (N_7739,N_6909,N_6777);
nor U7740 (N_7740,N_6348,N_6931);
or U7741 (N_7741,N_6747,N_6645);
nand U7742 (N_7742,N_6617,N_6502);
or U7743 (N_7743,N_6632,N_6742);
xor U7744 (N_7744,N_6837,N_6095);
nor U7745 (N_7745,N_6901,N_6637);
and U7746 (N_7746,N_6988,N_6946);
nor U7747 (N_7747,N_6118,N_6880);
and U7748 (N_7748,N_6207,N_6255);
xor U7749 (N_7749,N_6842,N_6983);
and U7750 (N_7750,N_6360,N_6188);
or U7751 (N_7751,N_6925,N_6357);
xor U7752 (N_7752,N_6302,N_6453);
nor U7753 (N_7753,N_6570,N_6001);
nand U7754 (N_7754,N_6785,N_6425);
nand U7755 (N_7755,N_6310,N_6755);
nand U7756 (N_7756,N_6647,N_6763);
xor U7757 (N_7757,N_6610,N_6685);
nor U7758 (N_7758,N_6194,N_6687);
or U7759 (N_7759,N_6435,N_6290);
xor U7760 (N_7760,N_6323,N_6597);
and U7761 (N_7761,N_6963,N_6528);
xor U7762 (N_7762,N_6978,N_6244);
nor U7763 (N_7763,N_6897,N_6962);
or U7764 (N_7764,N_6739,N_6328);
nand U7765 (N_7765,N_6287,N_6564);
nand U7766 (N_7766,N_6655,N_6972);
or U7767 (N_7767,N_6291,N_6092);
xnor U7768 (N_7768,N_6590,N_6862);
nand U7769 (N_7769,N_6863,N_6557);
and U7770 (N_7770,N_6287,N_6718);
xnor U7771 (N_7771,N_6330,N_6447);
or U7772 (N_7772,N_6060,N_6912);
and U7773 (N_7773,N_6843,N_6571);
and U7774 (N_7774,N_6051,N_6935);
nand U7775 (N_7775,N_6222,N_6537);
nor U7776 (N_7776,N_6404,N_6624);
and U7777 (N_7777,N_6857,N_6130);
and U7778 (N_7778,N_6816,N_6335);
nand U7779 (N_7779,N_6926,N_6314);
xor U7780 (N_7780,N_6840,N_6509);
or U7781 (N_7781,N_6054,N_6205);
xnor U7782 (N_7782,N_6113,N_6933);
xnor U7783 (N_7783,N_6146,N_6600);
nand U7784 (N_7784,N_6850,N_6685);
xnor U7785 (N_7785,N_6077,N_6584);
and U7786 (N_7786,N_6003,N_6776);
nor U7787 (N_7787,N_6856,N_6000);
and U7788 (N_7788,N_6184,N_6732);
and U7789 (N_7789,N_6577,N_6966);
nand U7790 (N_7790,N_6478,N_6025);
and U7791 (N_7791,N_6996,N_6306);
xnor U7792 (N_7792,N_6219,N_6943);
nand U7793 (N_7793,N_6853,N_6756);
or U7794 (N_7794,N_6129,N_6925);
xnor U7795 (N_7795,N_6364,N_6313);
nand U7796 (N_7796,N_6956,N_6674);
nand U7797 (N_7797,N_6223,N_6326);
xnor U7798 (N_7798,N_6226,N_6116);
nand U7799 (N_7799,N_6364,N_6659);
and U7800 (N_7800,N_6315,N_6022);
xor U7801 (N_7801,N_6961,N_6270);
nor U7802 (N_7802,N_6533,N_6965);
and U7803 (N_7803,N_6381,N_6904);
and U7804 (N_7804,N_6524,N_6276);
xnor U7805 (N_7805,N_6027,N_6531);
or U7806 (N_7806,N_6098,N_6310);
nor U7807 (N_7807,N_6021,N_6396);
nand U7808 (N_7808,N_6955,N_6356);
nor U7809 (N_7809,N_6824,N_6339);
nor U7810 (N_7810,N_6112,N_6888);
or U7811 (N_7811,N_6516,N_6495);
or U7812 (N_7812,N_6027,N_6077);
or U7813 (N_7813,N_6164,N_6980);
or U7814 (N_7814,N_6064,N_6599);
nor U7815 (N_7815,N_6652,N_6167);
nor U7816 (N_7816,N_6542,N_6377);
and U7817 (N_7817,N_6486,N_6647);
nand U7818 (N_7818,N_6918,N_6795);
nor U7819 (N_7819,N_6486,N_6576);
nor U7820 (N_7820,N_6467,N_6016);
or U7821 (N_7821,N_6669,N_6643);
xor U7822 (N_7822,N_6023,N_6114);
and U7823 (N_7823,N_6418,N_6613);
nand U7824 (N_7824,N_6309,N_6626);
nand U7825 (N_7825,N_6497,N_6580);
or U7826 (N_7826,N_6697,N_6977);
and U7827 (N_7827,N_6027,N_6114);
xor U7828 (N_7828,N_6683,N_6543);
xor U7829 (N_7829,N_6100,N_6659);
nor U7830 (N_7830,N_6303,N_6430);
xnor U7831 (N_7831,N_6130,N_6723);
xor U7832 (N_7832,N_6982,N_6365);
and U7833 (N_7833,N_6185,N_6750);
nand U7834 (N_7834,N_6816,N_6951);
nor U7835 (N_7835,N_6407,N_6919);
or U7836 (N_7836,N_6689,N_6721);
xnor U7837 (N_7837,N_6565,N_6462);
nor U7838 (N_7838,N_6652,N_6927);
and U7839 (N_7839,N_6827,N_6938);
xnor U7840 (N_7840,N_6361,N_6824);
and U7841 (N_7841,N_6930,N_6016);
nor U7842 (N_7842,N_6068,N_6211);
xnor U7843 (N_7843,N_6075,N_6222);
and U7844 (N_7844,N_6455,N_6322);
xnor U7845 (N_7845,N_6534,N_6389);
nor U7846 (N_7846,N_6349,N_6283);
nand U7847 (N_7847,N_6651,N_6546);
nor U7848 (N_7848,N_6611,N_6371);
nor U7849 (N_7849,N_6074,N_6607);
nand U7850 (N_7850,N_6792,N_6391);
xnor U7851 (N_7851,N_6863,N_6247);
and U7852 (N_7852,N_6666,N_6383);
nand U7853 (N_7853,N_6913,N_6005);
nand U7854 (N_7854,N_6412,N_6821);
xnor U7855 (N_7855,N_6571,N_6085);
and U7856 (N_7856,N_6640,N_6116);
or U7857 (N_7857,N_6361,N_6509);
and U7858 (N_7858,N_6100,N_6579);
and U7859 (N_7859,N_6447,N_6704);
xor U7860 (N_7860,N_6782,N_6023);
nand U7861 (N_7861,N_6985,N_6295);
xnor U7862 (N_7862,N_6961,N_6701);
and U7863 (N_7863,N_6477,N_6778);
xor U7864 (N_7864,N_6767,N_6019);
xor U7865 (N_7865,N_6763,N_6919);
and U7866 (N_7866,N_6019,N_6323);
nand U7867 (N_7867,N_6210,N_6760);
nor U7868 (N_7868,N_6093,N_6164);
and U7869 (N_7869,N_6742,N_6538);
nand U7870 (N_7870,N_6351,N_6079);
nor U7871 (N_7871,N_6036,N_6833);
or U7872 (N_7872,N_6227,N_6246);
xnor U7873 (N_7873,N_6342,N_6557);
nand U7874 (N_7874,N_6549,N_6146);
or U7875 (N_7875,N_6790,N_6892);
nor U7876 (N_7876,N_6691,N_6291);
nor U7877 (N_7877,N_6272,N_6974);
xnor U7878 (N_7878,N_6689,N_6994);
xnor U7879 (N_7879,N_6307,N_6968);
and U7880 (N_7880,N_6931,N_6785);
nor U7881 (N_7881,N_6431,N_6615);
or U7882 (N_7882,N_6869,N_6818);
or U7883 (N_7883,N_6299,N_6296);
nor U7884 (N_7884,N_6370,N_6598);
xor U7885 (N_7885,N_6256,N_6219);
or U7886 (N_7886,N_6412,N_6922);
nand U7887 (N_7887,N_6174,N_6876);
xnor U7888 (N_7888,N_6812,N_6461);
nor U7889 (N_7889,N_6402,N_6311);
or U7890 (N_7890,N_6282,N_6643);
and U7891 (N_7891,N_6733,N_6367);
or U7892 (N_7892,N_6808,N_6250);
nor U7893 (N_7893,N_6470,N_6594);
nand U7894 (N_7894,N_6132,N_6918);
nand U7895 (N_7895,N_6711,N_6260);
and U7896 (N_7896,N_6077,N_6521);
xnor U7897 (N_7897,N_6491,N_6266);
or U7898 (N_7898,N_6300,N_6822);
nor U7899 (N_7899,N_6856,N_6163);
nor U7900 (N_7900,N_6725,N_6614);
and U7901 (N_7901,N_6224,N_6152);
nand U7902 (N_7902,N_6120,N_6829);
or U7903 (N_7903,N_6185,N_6719);
nand U7904 (N_7904,N_6757,N_6931);
nand U7905 (N_7905,N_6691,N_6672);
or U7906 (N_7906,N_6463,N_6923);
and U7907 (N_7907,N_6561,N_6243);
xnor U7908 (N_7908,N_6731,N_6942);
nor U7909 (N_7909,N_6850,N_6627);
nand U7910 (N_7910,N_6656,N_6058);
nor U7911 (N_7911,N_6496,N_6191);
nand U7912 (N_7912,N_6992,N_6306);
nor U7913 (N_7913,N_6901,N_6171);
and U7914 (N_7914,N_6403,N_6324);
or U7915 (N_7915,N_6959,N_6138);
nand U7916 (N_7916,N_6853,N_6431);
nor U7917 (N_7917,N_6520,N_6126);
xnor U7918 (N_7918,N_6139,N_6581);
and U7919 (N_7919,N_6389,N_6834);
xnor U7920 (N_7920,N_6202,N_6198);
or U7921 (N_7921,N_6362,N_6612);
or U7922 (N_7922,N_6533,N_6826);
nand U7923 (N_7923,N_6863,N_6391);
xnor U7924 (N_7924,N_6282,N_6037);
or U7925 (N_7925,N_6700,N_6278);
nor U7926 (N_7926,N_6790,N_6943);
nand U7927 (N_7927,N_6274,N_6996);
and U7928 (N_7928,N_6477,N_6221);
or U7929 (N_7929,N_6444,N_6353);
and U7930 (N_7930,N_6012,N_6785);
xor U7931 (N_7931,N_6473,N_6796);
xnor U7932 (N_7932,N_6800,N_6250);
and U7933 (N_7933,N_6299,N_6631);
and U7934 (N_7934,N_6610,N_6384);
xor U7935 (N_7935,N_6566,N_6968);
nand U7936 (N_7936,N_6535,N_6848);
xnor U7937 (N_7937,N_6555,N_6313);
xor U7938 (N_7938,N_6373,N_6178);
or U7939 (N_7939,N_6458,N_6173);
xnor U7940 (N_7940,N_6236,N_6665);
or U7941 (N_7941,N_6424,N_6612);
nand U7942 (N_7942,N_6739,N_6245);
or U7943 (N_7943,N_6774,N_6358);
nand U7944 (N_7944,N_6184,N_6584);
or U7945 (N_7945,N_6313,N_6760);
nand U7946 (N_7946,N_6901,N_6152);
or U7947 (N_7947,N_6650,N_6643);
and U7948 (N_7948,N_6391,N_6678);
or U7949 (N_7949,N_6759,N_6973);
nand U7950 (N_7950,N_6748,N_6597);
nand U7951 (N_7951,N_6832,N_6530);
and U7952 (N_7952,N_6882,N_6199);
and U7953 (N_7953,N_6419,N_6274);
nand U7954 (N_7954,N_6963,N_6443);
nor U7955 (N_7955,N_6524,N_6762);
and U7956 (N_7956,N_6430,N_6887);
and U7957 (N_7957,N_6167,N_6634);
nand U7958 (N_7958,N_6392,N_6618);
xor U7959 (N_7959,N_6847,N_6007);
nand U7960 (N_7960,N_6539,N_6254);
nor U7961 (N_7961,N_6973,N_6179);
or U7962 (N_7962,N_6715,N_6379);
nand U7963 (N_7963,N_6456,N_6769);
xor U7964 (N_7964,N_6901,N_6266);
or U7965 (N_7965,N_6749,N_6309);
and U7966 (N_7966,N_6105,N_6099);
xnor U7967 (N_7967,N_6566,N_6639);
nand U7968 (N_7968,N_6577,N_6151);
nor U7969 (N_7969,N_6844,N_6276);
xor U7970 (N_7970,N_6588,N_6147);
xnor U7971 (N_7971,N_6694,N_6756);
and U7972 (N_7972,N_6077,N_6850);
nor U7973 (N_7973,N_6947,N_6545);
xor U7974 (N_7974,N_6113,N_6402);
and U7975 (N_7975,N_6896,N_6162);
and U7976 (N_7976,N_6245,N_6668);
and U7977 (N_7977,N_6046,N_6172);
nand U7978 (N_7978,N_6303,N_6305);
and U7979 (N_7979,N_6740,N_6670);
or U7980 (N_7980,N_6119,N_6951);
xnor U7981 (N_7981,N_6012,N_6729);
nand U7982 (N_7982,N_6361,N_6369);
or U7983 (N_7983,N_6931,N_6037);
and U7984 (N_7984,N_6447,N_6096);
nor U7985 (N_7985,N_6969,N_6006);
or U7986 (N_7986,N_6297,N_6540);
and U7987 (N_7987,N_6735,N_6367);
nor U7988 (N_7988,N_6221,N_6761);
nand U7989 (N_7989,N_6848,N_6386);
and U7990 (N_7990,N_6339,N_6585);
nand U7991 (N_7991,N_6706,N_6261);
nor U7992 (N_7992,N_6030,N_6994);
and U7993 (N_7993,N_6635,N_6602);
and U7994 (N_7994,N_6604,N_6550);
xor U7995 (N_7995,N_6448,N_6575);
xor U7996 (N_7996,N_6957,N_6615);
nand U7997 (N_7997,N_6977,N_6884);
nand U7998 (N_7998,N_6224,N_6500);
xor U7999 (N_7999,N_6793,N_6569);
or U8000 (N_8000,N_7457,N_7084);
nand U8001 (N_8001,N_7267,N_7953);
nor U8002 (N_8002,N_7619,N_7799);
nor U8003 (N_8003,N_7256,N_7897);
and U8004 (N_8004,N_7978,N_7017);
nand U8005 (N_8005,N_7542,N_7821);
and U8006 (N_8006,N_7390,N_7153);
xor U8007 (N_8007,N_7810,N_7329);
and U8008 (N_8008,N_7307,N_7512);
nand U8009 (N_8009,N_7890,N_7187);
nor U8010 (N_8010,N_7046,N_7221);
nor U8011 (N_8011,N_7475,N_7443);
nand U8012 (N_8012,N_7743,N_7868);
and U8013 (N_8013,N_7614,N_7081);
or U8014 (N_8014,N_7060,N_7927);
nor U8015 (N_8015,N_7131,N_7013);
nand U8016 (N_8016,N_7015,N_7887);
and U8017 (N_8017,N_7739,N_7867);
nand U8018 (N_8018,N_7637,N_7128);
and U8019 (N_8019,N_7011,N_7252);
or U8020 (N_8020,N_7848,N_7106);
or U8021 (N_8021,N_7581,N_7695);
and U8022 (N_8022,N_7892,N_7566);
or U8023 (N_8023,N_7056,N_7444);
and U8024 (N_8024,N_7731,N_7213);
nand U8025 (N_8025,N_7946,N_7020);
nand U8026 (N_8026,N_7723,N_7853);
nand U8027 (N_8027,N_7157,N_7211);
or U8028 (N_8028,N_7682,N_7005);
nor U8029 (N_8029,N_7163,N_7206);
and U8030 (N_8030,N_7369,N_7626);
nor U8031 (N_8031,N_7347,N_7819);
nand U8032 (N_8032,N_7415,N_7171);
nor U8033 (N_8033,N_7126,N_7753);
nand U8034 (N_8034,N_7006,N_7893);
and U8035 (N_8035,N_7125,N_7918);
nand U8036 (N_8036,N_7939,N_7297);
and U8037 (N_8037,N_7662,N_7716);
nor U8038 (N_8038,N_7782,N_7485);
xnor U8039 (N_8039,N_7278,N_7790);
or U8040 (N_8040,N_7822,N_7676);
nand U8041 (N_8041,N_7098,N_7692);
or U8042 (N_8042,N_7580,N_7730);
nor U8043 (N_8043,N_7228,N_7570);
or U8044 (N_8044,N_7969,N_7933);
or U8045 (N_8045,N_7191,N_7697);
xor U8046 (N_8046,N_7551,N_7370);
and U8047 (N_8047,N_7332,N_7247);
or U8048 (N_8048,N_7384,N_7631);
xor U8049 (N_8049,N_7660,N_7583);
and U8050 (N_8050,N_7378,N_7207);
xor U8051 (N_8051,N_7504,N_7104);
or U8052 (N_8052,N_7036,N_7321);
and U8053 (N_8053,N_7272,N_7747);
nand U8054 (N_8054,N_7667,N_7983);
or U8055 (N_8055,N_7497,N_7507);
and U8056 (N_8056,N_7473,N_7411);
or U8057 (N_8057,N_7041,N_7913);
nor U8058 (N_8058,N_7845,N_7721);
nand U8059 (N_8059,N_7051,N_7879);
xor U8060 (N_8060,N_7413,N_7296);
and U8061 (N_8061,N_7623,N_7405);
or U8062 (N_8062,N_7494,N_7178);
nand U8063 (N_8063,N_7082,N_7419);
nand U8064 (N_8064,N_7711,N_7737);
or U8065 (N_8065,N_7410,N_7803);
nor U8066 (N_8066,N_7699,N_7679);
and U8067 (N_8067,N_7266,N_7458);
xnor U8068 (N_8068,N_7154,N_7009);
and U8069 (N_8069,N_7857,N_7592);
xnor U8070 (N_8070,N_7740,N_7186);
and U8071 (N_8071,N_7787,N_7688);
xor U8072 (N_8072,N_7397,N_7764);
xnor U8073 (N_8073,N_7495,N_7996);
xor U8074 (N_8074,N_7701,N_7994);
nand U8075 (N_8075,N_7998,N_7238);
xnor U8076 (N_8076,N_7963,N_7896);
nor U8077 (N_8077,N_7536,N_7102);
xnor U8078 (N_8078,N_7841,N_7801);
nand U8079 (N_8079,N_7630,N_7816);
xnor U8080 (N_8080,N_7330,N_7085);
and U8081 (N_8081,N_7044,N_7202);
or U8082 (N_8082,N_7487,N_7677);
nand U8083 (N_8083,N_7094,N_7377);
and U8084 (N_8084,N_7018,N_7218);
xnor U8085 (N_8085,N_7000,N_7120);
nand U8086 (N_8086,N_7791,N_7636);
and U8087 (N_8087,N_7331,N_7964);
nor U8088 (N_8088,N_7024,N_7026);
nand U8089 (N_8089,N_7204,N_7649);
nor U8090 (N_8090,N_7869,N_7729);
nand U8091 (N_8091,N_7759,N_7883);
or U8092 (N_8092,N_7260,N_7048);
xnor U8093 (N_8093,N_7517,N_7972);
and U8094 (N_8094,N_7573,N_7875);
xor U8095 (N_8095,N_7601,N_7563);
nand U8096 (N_8096,N_7030,N_7261);
and U8097 (N_8097,N_7847,N_7664);
or U8098 (N_8098,N_7290,N_7921);
xnor U8099 (N_8099,N_7926,N_7451);
or U8100 (N_8100,N_7138,N_7426);
nor U8101 (N_8101,N_7915,N_7889);
and U8102 (N_8102,N_7912,N_7249);
xor U8103 (N_8103,N_7170,N_7696);
xor U8104 (N_8104,N_7123,N_7609);
and U8105 (N_8105,N_7666,N_7292);
or U8106 (N_8106,N_7680,N_7454);
or U8107 (N_8107,N_7312,N_7161);
and U8108 (N_8108,N_7217,N_7076);
nand U8109 (N_8109,N_7836,N_7949);
xnor U8110 (N_8110,N_7670,N_7728);
nand U8111 (N_8111,N_7245,N_7529);
xnor U8112 (N_8112,N_7557,N_7093);
nor U8113 (N_8113,N_7143,N_7371);
and U8114 (N_8114,N_7865,N_7718);
and U8115 (N_8115,N_7302,N_7834);
xnor U8116 (N_8116,N_7546,N_7215);
or U8117 (N_8117,N_7966,N_7936);
and U8118 (N_8118,N_7886,N_7045);
and U8119 (N_8119,N_7306,N_7641);
and U8120 (N_8120,N_7486,N_7310);
nand U8121 (N_8121,N_7379,N_7977);
nor U8122 (N_8122,N_7083,N_7356);
and U8123 (N_8123,N_7406,N_7422);
nand U8124 (N_8124,N_7719,N_7663);
and U8125 (N_8125,N_7057,N_7155);
nor U8126 (N_8126,N_7785,N_7600);
or U8127 (N_8127,N_7577,N_7770);
xnor U8128 (N_8128,N_7885,N_7201);
xor U8129 (N_8129,N_7383,N_7941);
or U8130 (N_8130,N_7337,N_7254);
nor U8131 (N_8131,N_7476,N_7944);
and U8132 (N_8132,N_7638,N_7672);
nand U8133 (N_8133,N_7762,N_7979);
nor U8134 (N_8134,N_7610,N_7109);
xnor U8135 (N_8135,N_7483,N_7802);
or U8136 (N_8136,N_7985,N_7856);
xnor U8137 (N_8137,N_7545,N_7231);
and U8138 (N_8138,N_7814,N_7535);
xnor U8139 (N_8139,N_7295,N_7352);
or U8140 (N_8140,N_7558,N_7524);
and U8141 (N_8141,N_7174,N_7427);
nor U8142 (N_8142,N_7940,N_7930);
and U8143 (N_8143,N_7008,N_7991);
or U8144 (N_8144,N_7040,N_7779);
nand U8145 (N_8145,N_7327,N_7523);
nor U8146 (N_8146,N_7172,N_7665);
nand U8147 (N_8147,N_7981,N_7830);
or U8148 (N_8148,N_7070,N_7360);
or U8149 (N_8149,N_7544,N_7771);
nor U8150 (N_8150,N_7162,N_7090);
and U8151 (N_8151,N_7250,N_7815);
and U8152 (N_8152,N_7077,N_7960);
nor U8153 (N_8153,N_7068,N_7804);
and U8154 (N_8154,N_7796,N_7831);
nor U8155 (N_8155,N_7606,N_7734);
or U8156 (N_8156,N_7611,N_7698);
or U8157 (N_8157,N_7904,N_7243);
or U8158 (N_8158,N_7744,N_7358);
nor U8159 (N_8159,N_7222,N_7756);
xor U8160 (N_8160,N_7087,N_7388);
and U8161 (N_8161,N_7055,N_7033);
xnor U8162 (N_8162,N_7229,N_7992);
or U8163 (N_8163,N_7633,N_7603);
nand U8164 (N_8164,N_7907,N_7112);
and U8165 (N_8165,N_7279,N_7361);
and U8166 (N_8166,N_7277,N_7318);
nand U8167 (N_8167,N_7226,N_7501);
nor U8168 (N_8168,N_7074,N_7767);
nand U8169 (N_8169,N_7237,N_7514);
nand U8170 (N_8170,N_7565,N_7835);
or U8171 (N_8171,N_7287,N_7351);
xor U8172 (N_8172,N_7141,N_7488);
nor U8173 (N_8173,N_7643,N_7425);
or U8174 (N_8174,N_7300,N_7876);
nor U8175 (N_8175,N_7525,N_7590);
nand U8176 (N_8176,N_7144,N_7653);
nor U8177 (N_8177,N_7650,N_7552);
nand U8178 (N_8178,N_7707,N_7119);
and U8179 (N_8179,N_7466,N_7188);
and U8180 (N_8180,N_7837,N_7232);
xor U8181 (N_8181,N_7066,N_7291);
nand U8182 (N_8182,N_7725,N_7530);
nor U8183 (N_8183,N_7655,N_7987);
nor U8184 (N_8184,N_7807,N_7965);
xnor U8185 (N_8185,N_7099,N_7346);
nor U8186 (N_8186,N_7812,N_7971);
or U8187 (N_8187,N_7160,N_7735);
nor U8188 (N_8188,N_7596,N_7622);
nor U8189 (N_8189,N_7608,N_7268);
xor U8190 (N_8190,N_7851,N_7948);
nand U8191 (N_8191,N_7850,N_7934);
and U8192 (N_8192,N_7414,N_7528);
nand U8193 (N_8193,N_7645,N_7316);
nor U8194 (N_8194,N_7304,N_7447);
nand U8195 (N_8195,N_7955,N_7103);
nand U8196 (N_8196,N_7129,N_7334);
xor U8197 (N_8197,N_7986,N_7298);
and U8198 (N_8198,N_7047,N_7362);
and U8199 (N_8199,N_7647,N_7895);
or U8200 (N_8200,N_7148,N_7537);
xnor U8201 (N_8201,N_7381,N_7811);
and U8202 (N_8202,N_7203,N_7449);
or U8203 (N_8203,N_7973,N_7441);
and U8204 (N_8204,N_7396,N_7309);
or U8205 (N_8205,N_7880,N_7715);
xnor U8206 (N_8206,N_7661,N_7825);
nor U8207 (N_8207,N_7429,N_7588);
or U8208 (N_8208,N_7092,N_7858);
nor U8209 (N_8209,N_7308,N_7374);
nand U8210 (N_8210,N_7866,N_7982);
xor U8211 (N_8211,N_7693,N_7271);
or U8212 (N_8212,N_7540,N_7617);
and U8213 (N_8213,N_7319,N_7376);
and U8214 (N_8214,N_7687,N_7209);
and U8215 (N_8215,N_7929,N_7548);
and U8216 (N_8216,N_7754,N_7627);
and U8217 (N_8217,N_7389,N_7673);
xnor U8218 (N_8218,N_7355,N_7002);
or U8219 (N_8219,N_7765,N_7065);
nor U8220 (N_8220,N_7958,N_7793);
nor U8221 (N_8221,N_7824,N_7763);
xnor U8222 (N_8222,N_7829,N_7445);
nand U8223 (N_8223,N_7169,N_7669);
and U8224 (N_8224,N_7778,N_7301);
or U8225 (N_8225,N_7274,N_7902);
nand U8226 (N_8226,N_7416,N_7976);
or U8227 (N_8227,N_7373,N_7937);
or U8228 (N_8228,N_7846,N_7962);
nor U8229 (N_8229,N_7299,N_7430);
xnor U8230 (N_8230,N_7380,N_7513);
nand U8231 (N_8231,N_7136,N_7532);
or U8232 (N_8232,N_7342,N_7648);
nand U8233 (N_8233,N_7919,N_7714);
and U8234 (N_8234,N_7181,N_7158);
and U8235 (N_8235,N_7736,N_7789);
nor U8236 (N_8236,N_7062,N_7275);
xnor U8237 (N_8237,N_7945,N_7959);
xor U8238 (N_8238,N_7881,N_7196);
nor U8239 (N_8239,N_7175,N_7950);
or U8240 (N_8240,N_7114,N_7900);
and U8241 (N_8241,N_7016,N_7724);
or U8242 (N_8242,N_7184,N_7738);
xor U8243 (N_8243,N_7364,N_7363);
or U8244 (N_8244,N_7111,N_7431);
and U8245 (N_8245,N_7792,N_7244);
nand U8246 (N_8246,N_7391,N_7854);
nand U8247 (N_8247,N_7461,N_7654);
xnor U8248 (N_8248,N_7042,N_7500);
xor U8249 (N_8249,N_7385,N_7280);
and U8250 (N_8250,N_7898,N_7255);
nor U8251 (N_8251,N_7025,N_7780);
xnor U8252 (N_8252,N_7100,N_7012);
nor U8253 (N_8253,N_7481,N_7855);
or U8254 (N_8254,N_7560,N_7720);
and U8255 (N_8255,N_7709,N_7489);
or U8256 (N_8256,N_7727,N_7624);
nor U8257 (N_8257,N_7039,N_7568);
xnor U8258 (N_8258,N_7906,N_7574);
xnor U8259 (N_8259,N_7579,N_7348);
and U8260 (N_8260,N_7700,N_7598);
nand U8261 (N_8261,N_7684,N_7997);
nand U8262 (N_8262,N_7233,N_7442);
or U8263 (N_8263,N_7561,N_7165);
and U8264 (N_8264,N_7484,N_7455);
and U8265 (N_8265,N_7285,N_7127);
xor U8266 (N_8266,N_7095,N_7938);
or U8267 (N_8267,N_7354,N_7368);
nand U8268 (N_8268,N_7200,N_7465);
and U8269 (N_8269,N_7974,N_7589);
xor U8270 (N_8270,N_7826,N_7818);
and U8271 (N_8271,N_7903,N_7021);
and U8272 (N_8272,N_7432,N_7531);
nor U8273 (N_8273,N_7185,N_7079);
xor U8274 (N_8274,N_7616,N_7452);
xnor U8275 (N_8275,N_7073,N_7943);
nor U8276 (N_8276,N_7311,N_7527);
and U8277 (N_8277,N_7409,N_7145);
or U8278 (N_8278,N_7935,N_7220);
or U8279 (N_8279,N_7151,N_7556);
or U8280 (N_8280,N_7706,N_7671);
and U8281 (N_8281,N_7061,N_7493);
and U8282 (N_8282,N_7198,N_7176);
or U8283 (N_8283,N_7899,N_7263);
and U8284 (N_8284,N_7491,N_7553);
nor U8285 (N_8285,N_7407,N_7597);
xor U8286 (N_8286,N_7757,N_7620);
nand U8287 (N_8287,N_7262,N_7450);
xnor U8288 (N_8288,N_7156,N_7599);
and U8289 (N_8289,N_7035,N_7418);
nor U8290 (N_8290,N_7269,N_7420);
or U8291 (N_8291,N_7058,N_7506);
nor U8292 (N_8292,N_7490,N_7505);
xnor U8293 (N_8293,N_7224,N_7468);
or U8294 (N_8294,N_7794,N_7547);
xor U8295 (N_8295,N_7216,N_7519);
and U8296 (N_8296,N_7089,N_7951);
xnor U8297 (N_8297,N_7894,N_7192);
nand U8298 (N_8298,N_7205,N_7795);
nand U8299 (N_8299,N_7908,N_7336);
xnor U8300 (N_8300,N_7595,N_7550);
nand U8301 (N_8301,N_7375,N_7434);
and U8302 (N_8302,N_7503,N_7054);
nor U8303 (N_8303,N_7417,N_7022);
or U8304 (N_8304,N_7014,N_7132);
xor U8305 (N_8305,N_7859,N_7395);
or U8306 (N_8306,N_7080,N_7587);
and U8307 (N_8307,N_7947,N_7117);
nand U8308 (N_8308,N_7471,N_7029);
nand U8309 (N_8309,N_7717,N_7652);
and U8310 (N_8310,N_7572,N_7146);
and U8311 (N_8311,N_7844,N_7852);
and U8312 (N_8312,N_7477,N_7694);
nand U8313 (N_8313,N_7251,N_7710);
nand U8314 (N_8314,N_7382,N_7223);
nand U8315 (N_8315,N_7349,N_7028);
xnor U8316 (N_8316,N_7635,N_7657);
nor U8317 (N_8317,N_7871,N_7877);
nor U8318 (N_8318,N_7980,N_7862);
nor U8319 (N_8319,N_7179,N_7470);
xnor U8320 (N_8320,N_7359,N_7408);
nor U8321 (N_8321,N_7428,N_7783);
and U8322 (N_8322,N_7562,N_7931);
xnor U8323 (N_8323,N_7511,N_7554);
and U8324 (N_8324,N_7078,N_7708);
nand U8325 (N_8325,N_7387,N_7571);
or U8326 (N_8326,N_7928,N_7340);
nand U8327 (N_8327,N_7402,N_7833);
nand U8328 (N_8328,N_7464,N_7303);
and U8329 (N_8329,N_7874,N_7448);
nor U8330 (N_8330,N_7462,N_7400);
xor U8331 (N_8331,N_7433,N_7576);
or U8332 (N_8332,N_7970,N_7749);
and U8333 (N_8333,N_7122,N_7745);
xor U8334 (N_8334,N_7543,N_7777);
xor U8335 (N_8335,N_7001,N_7164);
nor U8336 (N_8336,N_7037,N_7492);
nand U8337 (N_8337,N_7242,N_7108);
or U8338 (N_8338,N_7878,N_7999);
or U8339 (N_8339,N_7197,N_7173);
and U8340 (N_8340,N_7742,N_7870);
xor U8341 (N_8341,N_7586,N_7459);
or U8342 (N_8342,N_7265,N_7518);
nor U8343 (N_8343,N_7118,N_7975);
and U8344 (N_8344,N_7726,N_7788);
and U8345 (N_8345,N_7317,N_7957);
nand U8346 (N_8346,N_7607,N_7393);
nand U8347 (N_8347,N_7798,N_7593);
nand U8348 (N_8348,N_7049,N_7520);
nand U8349 (N_8349,N_7281,N_7526);
xor U8350 (N_8350,N_7235,N_7605);
nor U8351 (N_8351,N_7088,N_7861);
nor U8352 (N_8352,N_7195,N_7463);
nor U8353 (N_8353,N_7366,N_7335);
nand U8354 (N_8354,N_7843,N_7456);
nor U8355 (N_8355,N_7225,N_7258);
or U8356 (N_8356,N_7967,N_7293);
nand U8357 (N_8357,N_7690,N_7472);
nor U8358 (N_8358,N_7584,N_7559);
nor U8359 (N_8359,N_7282,N_7704);
nor U8360 (N_8360,N_7142,N_7618);
or U8361 (N_8361,N_7863,N_7133);
nand U8362 (N_8362,N_7421,N_7043);
or U8363 (N_8363,N_7681,N_7350);
or U8364 (N_8364,N_7034,N_7032);
nand U8365 (N_8365,N_7467,N_7167);
and U8366 (N_8366,N_7817,N_7403);
xor U8367 (N_8367,N_7923,N_7438);
nor U8368 (N_8368,N_7091,N_7924);
nor U8369 (N_8369,N_7784,N_7343);
xor U8370 (N_8370,N_7678,N_7773);
xor U8371 (N_8371,N_7901,N_7023);
nor U8372 (N_8372,N_7910,N_7806);
and U8373 (N_8373,N_7440,N_7686);
or U8374 (N_8374,N_7236,N_7639);
xor U8375 (N_8375,N_7642,N_7446);
xnor U8376 (N_8376,N_7555,N_7479);
and U8377 (N_8377,N_7404,N_7294);
xnor U8378 (N_8378,N_7193,N_7752);
nand U8379 (N_8379,N_7152,N_7072);
or U8380 (N_8380,N_7139,N_7864);
or U8381 (N_8381,N_7702,N_7071);
or U8382 (N_8382,N_7180,N_7344);
or U8383 (N_8383,N_7110,N_7199);
nor U8384 (N_8384,N_7741,N_7732);
nor U8385 (N_8385,N_7832,N_7038);
nand U8386 (N_8386,N_7137,N_7594);
nand U8387 (N_8387,N_7629,N_7140);
or U8388 (N_8388,N_7917,N_7283);
nor U8389 (N_8389,N_7827,N_7190);
or U8390 (N_8390,N_7891,N_7534);
nand U8391 (N_8391,N_7365,N_7713);
nand U8392 (N_8392,N_7182,N_7659);
nor U8393 (N_8393,N_7988,N_7746);
and U8394 (N_8394,N_7345,N_7750);
and U8395 (N_8395,N_7952,N_7149);
or U8396 (N_8396,N_7257,N_7888);
xnor U8397 (N_8397,N_7183,N_7159);
or U8398 (N_8398,N_7423,N_7766);
nand U8399 (N_8399,N_7840,N_7989);
nand U8400 (N_8400,N_7474,N_7357);
or U8401 (N_8401,N_7984,N_7401);
and U8402 (N_8402,N_7809,N_7634);
and U8403 (N_8403,N_7240,N_7480);
and U8404 (N_8404,N_7027,N_7394);
nand U8405 (N_8405,N_7932,N_7842);
nor U8406 (N_8406,N_7478,N_7961);
nand U8407 (N_8407,N_7567,N_7115);
xor U8408 (N_8408,N_7063,N_7135);
xnor U8409 (N_8409,N_7805,N_7632);
nand U8410 (N_8410,N_7499,N_7284);
and U8411 (N_8411,N_7691,N_7776);
xor U8412 (N_8412,N_7522,N_7651);
nand U8413 (N_8413,N_7230,N_7786);
xnor U8414 (N_8414,N_7323,N_7305);
or U8415 (N_8415,N_7675,N_7640);
xnor U8416 (N_8416,N_7482,N_7105);
and U8417 (N_8417,N_7591,N_7575);
nor U8418 (N_8418,N_7498,N_7733);
xnor U8419 (N_8419,N_7515,N_7769);
nand U8420 (N_8420,N_7124,N_7496);
and U8421 (N_8421,N_7705,N_7516);
nor U8422 (N_8422,N_7121,N_7399);
xor U8423 (N_8423,N_7234,N_7521);
nand U8424 (N_8424,N_7166,N_7813);
nor U8425 (N_8425,N_7549,N_7270);
nand U8426 (N_8426,N_7147,N_7069);
nor U8427 (N_8427,N_7324,N_7541);
xnor U8428 (N_8428,N_7905,N_7656);
and U8429 (N_8429,N_7050,N_7194);
nand U8430 (N_8430,N_7797,N_7644);
nor U8431 (N_8431,N_7758,N_7621);
nand U8432 (N_8432,N_7774,N_7510);
nand U8433 (N_8433,N_7398,N_7322);
and U8434 (N_8434,N_7003,N_7392);
xor U8435 (N_8435,N_7059,N_7315);
or U8436 (N_8436,N_7538,N_7646);
nor U8437 (N_8437,N_7925,N_7189);
nand U8438 (N_8438,N_7276,N_7683);
or U8439 (N_8439,N_7004,N_7435);
and U8440 (N_8440,N_7314,N_7031);
xnor U8441 (N_8441,N_7968,N_7075);
xnor U8442 (N_8442,N_7751,N_7007);
nor U8443 (N_8443,N_7722,N_7772);
nor U8444 (N_8444,N_7674,N_7097);
xnor U8445 (N_8445,N_7325,N_7320);
and U8446 (N_8446,N_7286,N_7882);
nor U8447 (N_8447,N_7253,N_7820);
xnor U8448 (N_8448,N_7689,N_7755);
and U8449 (N_8449,N_7239,N_7386);
or U8450 (N_8450,N_7326,N_7439);
and U8451 (N_8451,N_7338,N_7838);
nor U8452 (N_8452,N_7096,N_7177);
or U8453 (N_8453,N_7585,N_7502);
or U8454 (N_8454,N_7288,N_7911);
nand U8455 (N_8455,N_7839,N_7508);
and U8456 (N_8456,N_7768,N_7703);
nand U8457 (N_8457,N_7509,N_7064);
nor U8458 (N_8458,N_7248,N_7437);
or U8459 (N_8459,N_7067,N_7922);
or U8460 (N_8460,N_7412,N_7101);
nor U8461 (N_8461,N_7273,N_7849);
nor U8462 (N_8462,N_7993,N_7625);
and U8463 (N_8463,N_7328,N_7712);
or U8464 (N_8464,N_7914,N_7134);
nor U8465 (N_8465,N_7341,N_7353);
xnor U8466 (N_8466,N_7613,N_7995);
xor U8467 (N_8467,N_7289,N_7920);
xor U8468 (N_8468,N_7685,N_7564);
and U8469 (N_8469,N_7533,N_7052);
and U8470 (N_8470,N_7872,N_7246);
nor U8471 (N_8471,N_7942,N_7264);
nor U8472 (N_8472,N_7113,N_7775);
and U8473 (N_8473,N_7219,N_7241);
nor U8474 (N_8474,N_7873,N_7168);
or U8475 (N_8475,N_7990,N_7916);
or U8476 (N_8476,N_7010,N_7612);
nor U8477 (N_8477,N_7053,N_7823);
or U8478 (N_8478,N_7259,N_7453);
nand U8479 (N_8479,N_7615,N_7628);
and U8480 (N_8480,N_7760,N_7086);
xnor U8481 (N_8481,N_7469,N_7860);
nor U8482 (N_8482,N_7954,N_7436);
nor U8483 (N_8483,N_7828,N_7748);
xnor U8484 (N_8484,N_7116,N_7212);
nand U8485 (N_8485,N_7150,N_7582);
nor U8486 (N_8486,N_7227,N_7214);
nand U8487 (N_8487,N_7424,N_7130);
or U8488 (N_8488,N_7578,N_7333);
nor U8489 (N_8489,N_7107,N_7210);
nor U8490 (N_8490,N_7800,N_7569);
nand U8491 (N_8491,N_7761,N_7604);
nor U8492 (N_8492,N_7956,N_7884);
nor U8493 (N_8493,N_7658,N_7781);
xor U8494 (N_8494,N_7808,N_7539);
xnor U8495 (N_8495,N_7367,N_7208);
xor U8496 (N_8496,N_7602,N_7019);
and U8497 (N_8497,N_7339,N_7668);
nand U8498 (N_8498,N_7909,N_7372);
nor U8499 (N_8499,N_7313,N_7460);
nor U8500 (N_8500,N_7558,N_7525);
xnor U8501 (N_8501,N_7380,N_7761);
xnor U8502 (N_8502,N_7974,N_7952);
nor U8503 (N_8503,N_7975,N_7727);
xnor U8504 (N_8504,N_7446,N_7026);
nand U8505 (N_8505,N_7621,N_7823);
xor U8506 (N_8506,N_7367,N_7773);
or U8507 (N_8507,N_7211,N_7455);
nor U8508 (N_8508,N_7565,N_7878);
or U8509 (N_8509,N_7690,N_7340);
nor U8510 (N_8510,N_7525,N_7574);
or U8511 (N_8511,N_7300,N_7827);
or U8512 (N_8512,N_7010,N_7751);
or U8513 (N_8513,N_7340,N_7610);
and U8514 (N_8514,N_7598,N_7459);
nor U8515 (N_8515,N_7803,N_7683);
and U8516 (N_8516,N_7734,N_7781);
nand U8517 (N_8517,N_7604,N_7431);
or U8518 (N_8518,N_7254,N_7298);
or U8519 (N_8519,N_7169,N_7208);
or U8520 (N_8520,N_7914,N_7718);
nand U8521 (N_8521,N_7132,N_7004);
nand U8522 (N_8522,N_7086,N_7745);
and U8523 (N_8523,N_7781,N_7196);
and U8524 (N_8524,N_7800,N_7657);
nand U8525 (N_8525,N_7763,N_7157);
or U8526 (N_8526,N_7520,N_7613);
nand U8527 (N_8527,N_7075,N_7638);
xnor U8528 (N_8528,N_7990,N_7039);
or U8529 (N_8529,N_7890,N_7651);
nand U8530 (N_8530,N_7571,N_7317);
or U8531 (N_8531,N_7102,N_7092);
xor U8532 (N_8532,N_7787,N_7488);
nand U8533 (N_8533,N_7157,N_7874);
xor U8534 (N_8534,N_7842,N_7334);
nand U8535 (N_8535,N_7994,N_7179);
nand U8536 (N_8536,N_7038,N_7796);
xnor U8537 (N_8537,N_7897,N_7133);
xor U8538 (N_8538,N_7688,N_7092);
nand U8539 (N_8539,N_7837,N_7936);
or U8540 (N_8540,N_7005,N_7527);
nand U8541 (N_8541,N_7887,N_7670);
xor U8542 (N_8542,N_7248,N_7533);
nand U8543 (N_8543,N_7267,N_7883);
or U8544 (N_8544,N_7824,N_7042);
and U8545 (N_8545,N_7126,N_7277);
or U8546 (N_8546,N_7575,N_7219);
nand U8547 (N_8547,N_7135,N_7875);
and U8548 (N_8548,N_7271,N_7651);
and U8549 (N_8549,N_7696,N_7133);
nor U8550 (N_8550,N_7173,N_7328);
nand U8551 (N_8551,N_7915,N_7725);
xor U8552 (N_8552,N_7910,N_7496);
xor U8553 (N_8553,N_7196,N_7551);
and U8554 (N_8554,N_7467,N_7903);
nand U8555 (N_8555,N_7528,N_7669);
or U8556 (N_8556,N_7464,N_7099);
nand U8557 (N_8557,N_7839,N_7524);
nor U8558 (N_8558,N_7493,N_7157);
or U8559 (N_8559,N_7205,N_7682);
xnor U8560 (N_8560,N_7610,N_7626);
nor U8561 (N_8561,N_7566,N_7228);
nand U8562 (N_8562,N_7957,N_7442);
xnor U8563 (N_8563,N_7255,N_7955);
xor U8564 (N_8564,N_7827,N_7442);
nor U8565 (N_8565,N_7748,N_7322);
xor U8566 (N_8566,N_7411,N_7968);
nor U8567 (N_8567,N_7121,N_7545);
nand U8568 (N_8568,N_7767,N_7500);
nor U8569 (N_8569,N_7905,N_7495);
nand U8570 (N_8570,N_7752,N_7879);
nor U8571 (N_8571,N_7527,N_7328);
nor U8572 (N_8572,N_7299,N_7203);
nand U8573 (N_8573,N_7771,N_7022);
nand U8574 (N_8574,N_7977,N_7378);
nand U8575 (N_8575,N_7109,N_7650);
xnor U8576 (N_8576,N_7467,N_7230);
nand U8577 (N_8577,N_7328,N_7450);
nor U8578 (N_8578,N_7623,N_7118);
or U8579 (N_8579,N_7851,N_7906);
or U8580 (N_8580,N_7795,N_7143);
or U8581 (N_8581,N_7316,N_7819);
and U8582 (N_8582,N_7081,N_7745);
and U8583 (N_8583,N_7682,N_7776);
and U8584 (N_8584,N_7880,N_7717);
or U8585 (N_8585,N_7732,N_7195);
nand U8586 (N_8586,N_7149,N_7741);
nor U8587 (N_8587,N_7207,N_7092);
and U8588 (N_8588,N_7711,N_7742);
nand U8589 (N_8589,N_7778,N_7772);
xnor U8590 (N_8590,N_7601,N_7412);
and U8591 (N_8591,N_7468,N_7699);
and U8592 (N_8592,N_7444,N_7017);
nor U8593 (N_8593,N_7536,N_7942);
or U8594 (N_8594,N_7195,N_7814);
nor U8595 (N_8595,N_7166,N_7745);
nand U8596 (N_8596,N_7245,N_7026);
xor U8597 (N_8597,N_7333,N_7432);
nand U8598 (N_8598,N_7991,N_7870);
or U8599 (N_8599,N_7593,N_7632);
and U8600 (N_8600,N_7526,N_7369);
nor U8601 (N_8601,N_7710,N_7169);
and U8602 (N_8602,N_7383,N_7376);
nor U8603 (N_8603,N_7382,N_7899);
xor U8604 (N_8604,N_7078,N_7221);
nand U8605 (N_8605,N_7742,N_7739);
or U8606 (N_8606,N_7097,N_7149);
nor U8607 (N_8607,N_7324,N_7926);
nor U8608 (N_8608,N_7052,N_7726);
nand U8609 (N_8609,N_7664,N_7566);
nand U8610 (N_8610,N_7845,N_7675);
or U8611 (N_8611,N_7268,N_7632);
nand U8612 (N_8612,N_7270,N_7726);
and U8613 (N_8613,N_7467,N_7551);
and U8614 (N_8614,N_7446,N_7897);
xnor U8615 (N_8615,N_7847,N_7071);
nand U8616 (N_8616,N_7953,N_7580);
nor U8617 (N_8617,N_7136,N_7086);
and U8618 (N_8618,N_7305,N_7853);
or U8619 (N_8619,N_7868,N_7628);
nor U8620 (N_8620,N_7457,N_7462);
or U8621 (N_8621,N_7486,N_7480);
nand U8622 (N_8622,N_7743,N_7105);
and U8623 (N_8623,N_7569,N_7281);
nand U8624 (N_8624,N_7371,N_7081);
xor U8625 (N_8625,N_7092,N_7613);
xor U8626 (N_8626,N_7722,N_7506);
nand U8627 (N_8627,N_7064,N_7740);
xor U8628 (N_8628,N_7296,N_7424);
nand U8629 (N_8629,N_7067,N_7422);
nand U8630 (N_8630,N_7862,N_7021);
or U8631 (N_8631,N_7765,N_7738);
and U8632 (N_8632,N_7607,N_7495);
nor U8633 (N_8633,N_7614,N_7430);
or U8634 (N_8634,N_7883,N_7918);
nand U8635 (N_8635,N_7041,N_7856);
xor U8636 (N_8636,N_7917,N_7839);
nand U8637 (N_8637,N_7788,N_7920);
and U8638 (N_8638,N_7000,N_7560);
xor U8639 (N_8639,N_7642,N_7149);
and U8640 (N_8640,N_7154,N_7312);
and U8641 (N_8641,N_7354,N_7503);
and U8642 (N_8642,N_7336,N_7945);
xnor U8643 (N_8643,N_7365,N_7049);
nand U8644 (N_8644,N_7619,N_7060);
and U8645 (N_8645,N_7323,N_7967);
or U8646 (N_8646,N_7268,N_7702);
and U8647 (N_8647,N_7620,N_7231);
nand U8648 (N_8648,N_7798,N_7425);
and U8649 (N_8649,N_7670,N_7969);
and U8650 (N_8650,N_7870,N_7225);
nor U8651 (N_8651,N_7341,N_7494);
and U8652 (N_8652,N_7383,N_7774);
nor U8653 (N_8653,N_7989,N_7157);
xor U8654 (N_8654,N_7489,N_7667);
nor U8655 (N_8655,N_7376,N_7943);
and U8656 (N_8656,N_7137,N_7150);
and U8657 (N_8657,N_7285,N_7723);
and U8658 (N_8658,N_7939,N_7096);
nor U8659 (N_8659,N_7199,N_7590);
or U8660 (N_8660,N_7870,N_7070);
xnor U8661 (N_8661,N_7165,N_7668);
nor U8662 (N_8662,N_7936,N_7980);
xnor U8663 (N_8663,N_7142,N_7379);
or U8664 (N_8664,N_7593,N_7962);
nor U8665 (N_8665,N_7968,N_7352);
and U8666 (N_8666,N_7174,N_7142);
nand U8667 (N_8667,N_7654,N_7209);
and U8668 (N_8668,N_7739,N_7898);
xnor U8669 (N_8669,N_7217,N_7519);
and U8670 (N_8670,N_7030,N_7077);
or U8671 (N_8671,N_7097,N_7210);
xnor U8672 (N_8672,N_7657,N_7490);
xnor U8673 (N_8673,N_7855,N_7745);
or U8674 (N_8674,N_7134,N_7671);
or U8675 (N_8675,N_7754,N_7148);
xor U8676 (N_8676,N_7076,N_7424);
nor U8677 (N_8677,N_7892,N_7849);
nand U8678 (N_8678,N_7855,N_7131);
nor U8679 (N_8679,N_7088,N_7397);
xor U8680 (N_8680,N_7915,N_7319);
xor U8681 (N_8681,N_7134,N_7681);
or U8682 (N_8682,N_7620,N_7599);
and U8683 (N_8683,N_7183,N_7505);
or U8684 (N_8684,N_7517,N_7767);
and U8685 (N_8685,N_7008,N_7582);
or U8686 (N_8686,N_7109,N_7009);
and U8687 (N_8687,N_7090,N_7264);
xor U8688 (N_8688,N_7475,N_7886);
xnor U8689 (N_8689,N_7787,N_7693);
nor U8690 (N_8690,N_7441,N_7924);
xor U8691 (N_8691,N_7869,N_7551);
xor U8692 (N_8692,N_7730,N_7415);
nand U8693 (N_8693,N_7771,N_7595);
and U8694 (N_8694,N_7267,N_7012);
or U8695 (N_8695,N_7883,N_7611);
and U8696 (N_8696,N_7633,N_7689);
xor U8697 (N_8697,N_7149,N_7981);
or U8698 (N_8698,N_7441,N_7112);
and U8699 (N_8699,N_7788,N_7089);
nand U8700 (N_8700,N_7854,N_7201);
or U8701 (N_8701,N_7531,N_7614);
or U8702 (N_8702,N_7318,N_7585);
and U8703 (N_8703,N_7112,N_7923);
nor U8704 (N_8704,N_7523,N_7881);
nor U8705 (N_8705,N_7778,N_7653);
and U8706 (N_8706,N_7226,N_7344);
xor U8707 (N_8707,N_7803,N_7312);
and U8708 (N_8708,N_7080,N_7586);
and U8709 (N_8709,N_7810,N_7780);
nor U8710 (N_8710,N_7078,N_7050);
nand U8711 (N_8711,N_7599,N_7799);
nor U8712 (N_8712,N_7132,N_7556);
or U8713 (N_8713,N_7726,N_7072);
and U8714 (N_8714,N_7179,N_7316);
xor U8715 (N_8715,N_7216,N_7643);
xnor U8716 (N_8716,N_7226,N_7173);
nor U8717 (N_8717,N_7598,N_7134);
nand U8718 (N_8718,N_7088,N_7588);
nor U8719 (N_8719,N_7197,N_7256);
nand U8720 (N_8720,N_7990,N_7811);
and U8721 (N_8721,N_7304,N_7989);
and U8722 (N_8722,N_7012,N_7508);
or U8723 (N_8723,N_7739,N_7914);
xnor U8724 (N_8724,N_7373,N_7528);
and U8725 (N_8725,N_7299,N_7467);
xor U8726 (N_8726,N_7591,N_7134);
and U8727 (N_8727,N_7931,N_7469);
xnor U8728 (N_8728,N_7116,N_7181);
nand U8729 (N_8729,N_7462,N_7829);
and U8730 (N_8730,N_7357,N_7580);
and U8731 (N_8731,N_7219,N_7521);
xnor U8732 (N_8732,N_7174,N_7020);
and U8733 (N_8733,N_7016,N_7787);
nand U8734 (N_8734,N_7387,N_7493);
and U8735 (N_8735,N_7027,N_7143);
xnor U8736 (N_8736,N_7028,N_7553);
nor U8737 (N_8737,N_7767,N_7523);
xor U8738 (N_8738,N_7875,N_7619);
nor U8739 (N_8739,N_7102,N_7469);
xnor U8740 (N_8740,N_7822,N_7265);
nor U8741 (N_8741,N_7254,N_7353);
and U8742 (N_8742,N_7666,N_7647);
nand U8743 (N_8743,N_7133,N_7522);
xnor U8744 (N_8744,N_7838,N_7693);
nand U8745 (N_8745,N_7215,N_7284);
nor U8746 (N_8746,N_7045,N_7656);
or U8747 (N_8747,N_7856,N_7639);
xor U8748 (N_8748,N_7515,N_7690);
xnor U8749 (N_8749,N_7680,N_7573);
nor U8750 (N_8750,N_7951,N_7221);
or U8751 (N_8751,N_7620,N_7364);
xnor U8752 (N_8752,N_7238,N_7106);
or U8753 (N_8753,N_7877,N_7625);
and U8754 (N_8754,N_7049,N_7797);
nand U8755 (N_8755,N_7546,N_7566);
nor U8756 (N_8756,N_7448,N_7932);
xnor U8757 (N_8757,N_7182,N_7569);
nor U8758 (N_8758,N_7986,N_7962);
nand U8759 (N_8759,N_7182,N_7663);
and U8760 (N_8760,N_7867,N_7030);
and U8761 (N_8761,N_7512,N_7133);
nor U8762 (N_8762,N_7622,N_7161);
nor U8763 (N_8763,N_7097,N_7826);
nand U8764 (N_8764,N_7995,N_7439);
or U8765 (N_8765,N_7975,N_7181);
or U8766 (N_8766,N_7551,N_7067);
nor U8767 (N_8767,N_7079,N_7280);
or U8768 (N_8768,N_7440,N_7894);
xor U8769 (N_8769,N_7791,N_7044);
nand U8770 (N_8770,N_7779,N_7095);
xor U8771 (N_8771,N_7711,N_7376);
or U8772 (N_8772,N_7142,N_7230);
xor U8773 (N_8773,N_7178,N_7649);
nand U8774 (N_8774,N_7629,N_7013);
nor U8775 (N_8775,N_7980,N_7059);
or U8776 (N_8776,N_7714,N_7510);
xor U8777 (N_8777,N_7420,N_7364);
nand U8778 (N_8778,N_7239,N_7120);
xor U8779 (N_8779,N_7872,N_7559);
nor U8780 (N_8780,N_7669,N_7137);
nor U8781 (N_8781,N_7954,N_7281);
or U8782 (N_8782,N_7089,N_7559);
nand U8783 (N_8783,N_7804,N_7764);
xor U8784 (N_8784,N_7104,N_7491);
xnor U8785 (N_8785,N_7045,N_7016);
or U8786 (N_8786,N_7323,N_7186);
nor U8787 (N_8787,N_7103,N_7529);
xor U8788 (N_8788,N_7015,N_7441);
and U8789 (N_8789,N_7842,N_7636);
nor U8790 (N_8790,N_7970,N_7126);
or U8791 (N_8791,N_7058,N_7681);
or U8792 (N_8792,N_7279,N_7351);
and U8793 (N_8793,N_7234,N_7491);
or U8794 (N_8794,N_7636,N_7023);
xor U8795 (N_8795,N_7635,N_7444);
xnor U8796 (N_8796,N_7989,N_7527);
xor U8797 (N_8797,N_7375,N_7611);
xor U8798 (N_8798,N_7330,N_7446);
xnor U8799 (N_8799,N_7221,N_7092);
nor U8800 (N_8800,N_7484,N_7159);
or U8801 (N_8801,N_7786,N_7273);
nor U8802 (N_8802,N_7633,N_7926);
nor U8803 (N_8803,N_7413,N_7454);
nand U8804 (N_8804,N_7411,N_7793);
nor U8805 (N_8805,N_7864,N_7327);
nand U8806 (N_8806,N_7383,N_7871);
or U8807 (N_8807,N_7130,N_7553);
and U8808 (N_8808,N_7695,N_7312);
or U8809 (N_8809,N_7374,N_7319);
or U8810 (N_8810,N_7504,N_7667);
or U8811 (N_8811,N_7518,N_7357);
nor U8812 (N_8812,N_7944,N_7618);
nor U8813 (N_8813,N_7525,N_7439);
nor U8814 (N_8814,N_7007,N_7793);
nor U8815 (N_8815,N_7638,N_7348);
nor U8816 (N_8816,N_7001,N_7479);
and U8817 (N_8817,N_7365,N_7915);
and U8818 (N_8818,N_7701,N_7922);
xnor U8819 (N_8819,N_7960,N_7775);
or U8820 (N_8820,N_7284,N_7308);
and U8821 (N_8821,N_7482,N_7442);
nor U8822 (N_8822,N_7963,N_7695);
and U8823 (N_8823,N_7478,N_7850);
nand U8824 (N_8824,N_7435,N_7747);
xor U8825 (N_8825,N_7800,N_7367);
xor U8826 (N_8826,N_7591,N_7879);
xor U8827 (N_8827,N_7573,N_7822);
or U8828 (N_8828,N_7441,N_7104);
or U8829 (N_8829,N_7903,N_7426);
and U8830 (N_8830,N_7093,N_7027);
and U8831 (N_8831,N_7587,N_7982);
nor U8832 (N_8832,N_7569,N_7536);
nand U8833 (N_8833,N_7423,N_7717);
nor U8834 (N_8834,N_7725,N_7078);
nor U8835 (N_8835,N_7038,N_7143);
nand U8836 (N_8836,N_7925,N_7403);
or U8837 (N_8837,N_7497,N_7868);
and U8838 (N_8838,N_7843,N_7951);
and U8839 (N_8839,N_7229,N_7847);
nor U8840 (N_8840,N_7691,N_7857);
nor U8841 (N_8841,N_7957,N_7173);
nand U8842 (N_8842,N_7847,N_7136);
and U8843 (N_8843,N_7365,N_7497);
and U8844 (N_8844,N_7459,N_7412);
or U8845 (N_8845,N_7103,N_7178);
or U8846 (N_8846,N_7111,N_7145);
xnor U8847 (N_8847,N_7658,N_7007);
xor U8848 (N_8848,N_7494,N_7828);
or U8849 (N_8849,N_7148,N_7634);
and U8850 (N_8850,N_7191,N_7198);
nand U8851 (N_8851,N_7050,N_7801);
or U8852 (N_8852,N_7920,N_7284);
xor U8853 (N_8853,N_7304,N_7727);
or U8854 (N_8854,N_7488,N_7539);
nand U8855 (N_8855,N_7741,N_7461);
nand U8856 (N_8856,N_7236,N_7352);
and U8857 (N_8857,N_7139,N_7587);
nand U8858 (N_8858,N_7955,N_7180);
and U8859 (N_8859,N_7323,N_7713);
xor U8860 (N_8860,N_7629,N_7068);
xnor U8861 (N_8861,N_7595,N_7526);
nand U8862 (N_8862,N_7277,N_7279);
or U8863 (N_8863,N_7398,N_7331);
nor U8864 (N_8864,N_7808,N_7787);
and U8865 (N_8865,N_7416,N_7494);
nand U8866 (N_8866,N_7275,N_7492);
nand U8867 (N_8867,N_7601,N_7152);
nor U8868 (N_8868,N_7887,N_7328);
nor U8869 (N_8869,N_7354,N_7598);
and U8870 (N_8870,N_7918,N_7492);
nand U8871 (N_8871,N_7041,N_7465);
xor U8872 (N_8872,N_7882,N_7576);
nand U8873 (N_8873,N_7369,N_7939);
or U8874 (N_8874,N_7750,N_7254);
nor U8875 (N_8875,N_7693,N_7295);
nor U8876 (N_8876,N_7672,N_7446);
nand U8877 (N_8877,N_7537,N_7214);
nand U8878 (N_8878,N_7487,N_7745);
nand U8879 (N_8879,N_7748,N_7377);
and U8880 (N_8880,N_7361,N_7198);
or U8881 (N_8881,N_7817,N_7327);
or U8882 (N_8882,N_7825,N_7187);
nor U8883 (N_8883,N_7695,N_7757);
nor U8884 (N_8884,N_7942,N_7542);
nor U8885 (N_8885,N_7814,N_7895);
nand U8886 (N_8886,N_7774,N_7078);
nand U8887 (N_8887,N_7468,N_7151);
and U8888 (N_8888,N_7505,N_7736);
xor U8889 (N_8889,N_7713,N_7672);
nor U8890 (N_8890,N_7608,N_7527);
xor U8891 (N_8891,N_7266,N_7692);
nand U8892 (N_8892,N_7271,N_7536);
xor U8893 (N_8893,N_7008,N_7771);
and U8894 (N_8894,N_7276,N_7941);
nand U8895 (N_8895,N_7514,N_7773);
nor U8896 (N_8896,N_7757,N_7224);
and U8897 (N_8897,N_7098,N_7776);
nor U8898 (N_8898,N_7220,N_7979);
nand U8899 (N_8899,N_7373,N_7393);
xor U8900 (N_8900,N_7871,N_7025);
and U8901 (N_8901,N_7825,N_7483);
xnor U8902 (N_8902,N_7444,N_7878);
nand U8903 (N_8903,N_7658,N_7229);
or U8904 (N_8904,N_7825,N_7088);
xor U8905 (N_8905,N_7029,N_7732);
xnor U8906 (N_8906,N_7662,N_7503);
nor U8907 (N_8907,N_7809,N_7021);
or U8908 (N_8908,N_7077,N_7677);
nand U8909 (N_8909,N_7720,N_7593);
and U8910 (N_8910,N_7123,N_7043);
nor U8911 (N_8911,N_7191,N_7178);
or U8912 (N_8912,N_7479,N_7180);
xnor U8913 (N_8913,N_7787,N_7674);
or U8914 (N_8914,N_7861,N_7247);
xor U8915 (N_8915,N_7251,N_7537);
xnor U8916 (N_8916,N_7752,N_7019);
xor U8917 (N_8917,N_7909,N_7401);
xor U8918 (N_8918,N_7962,N_7927);
nand U8919 (N_8919,N_7550,N_7394);
xnor U8920 (N_8920,N_7966,N_7953);
or U8921 (N_8921,N_7698,N_7994);
nor U8922 (N_8922,N_7467,N_7870);
nand U8923 (N_8923,N_7021,N_7064);
xnor U8924 (N_8924,N_7574,N_7110);
nand U8925 (N_8925,N_7227,N_7281);
nand U8926 (N_8926,N_7648,N_7176);
nand U8927 (N_8927,N_7001,N_7387);
and U8928 (N_8928,N_7503,N_7658);
nor U8929 (N_8929,N_7080,N_7379);
xor U8930 (N_8930,N_7983,N_7652);
xnor U8931 (N_8931,N_7544,N_7610);
or U8932 (N_8932,N_7477,N_7757);
xor U8933 (N_8933,N_7120,N_7274);
xnor U8934 (N_8934,N_7474,N_7142);
xor U8935 (N_8935,N_7562,N_7738);
nor U8936 (N_8936,N_7207,N_7265);
and U8937 (N_8937,N_7210,N_7606);
or U8938 (N_8938,N_7410,N_7036);
nor U8939 (N_8939,N_7916,N_7176);
or U8940 (N_8940,N_7148,N_7625);
xnor U8941 (N_8941,N_7488,N_7750);
xnor U8942 (N_8942,N_7837,N_7017);
and U8943 (N_8943,N_7355,N_7695);
xor U8944 (N_8944,N_7869,N_7807);
nor U8945 (N_8945,N_7697,N_7729);
nand U8946 (N_8946,N_7771,N_7700);
nor U8947 (N_8947,N_7240,N_7710);
xor U8948 (N_8948,N_7749,N_7711);
and U8949 (N_8949,N_7762,N_7730);
xor U8950 (N_8950,N_7857,N_7777);
or U8951 (N_8951,N_7513,N_7135);
nor U8952 (N_8952,N_7516,N_7807);
nor U8953 (N_8953,N_7712,N_7682);
and U8954 (N_8954,N_7262,N_7081);
nand U8955 (N_8955,N_7137,N_7460);
xnor U8956 (N_8956,N_7082,N_7562);
xor U8957 (N_8957,N_7680,N_7028);
or U8958 (N_8958,N_7666,N_7274);
or U8959 (N_8959,N_7949,N_7722);
nor U8960 (N_8960,N_7539,N_7896);
nand U8961 (N_8961,N_7065,N_7135);
xnor U8962 (N_8962,N_7059,N_7368);
nor U8963 (N_8963,N_7642,N_7045);
nor U8964 (N_8964,N_7173,N_7053);
or U8965 (N_8965,N_7869,N_7087);
xor U8966 (N_8966,N_7064,N_7550);
nand U8967 (N_8967,N_7420,N_7468);
or U8968 (N_8968,N_7007,N_7815);
nand U8969 (N_8969,N_7780,N_7472);
or U8970 (N_8970,N_7199,N_7004);
or U8971 (N_8971,N_7639,N_7962);
xor U8972 (N_8972,N_7124,N_7524);
and U8973 (N_8973,N_7865,N_7627);
nor U8974 (N_8974,N_7881,N_7955);
and U8975 (N_8975,N_7777,N_7443);
nor U8976 (N_8976,N_7413,N_7027);
nand U8977 (N_8977,N_7621,N_7265);
and U8978 (N_8978,N_7587,N_7204);
xnor U8979 (N_8979,N_7698,N_7108);
or U8980 (N_8980,N_7870,N_7978);
and U8981 (N_8981,N_7716,N_7179);
and U8982 (N_8982,N_7670,N_7896);
nand U8983 (N_8983,N_7058,N_7930);
or U8984 (N_8984,N_7311,N_7797);
nand U8985 (N_8985,N_7767,N_7836);
nor U8986 (N_8986,N_7899,N_7279);
or U8987 (N_8987,N_7814,N_7609);
or U8988 (N_8988,N_7453,N_7495);
and U8989 (N_8989,N_7589,N_7089);
or U8990 (N_8990,N_7539,N_7147);
or U8991 (N_8991,N_7438,N_7615);
nor U8992 (N_8992,N_7571,N_7489);
or U8993 (N_8993,N_7530,N_7495);
or U8994 (N_8994,N_7686,N_7959);
nand U8995 (N_8995,N_7620,N_7046);
nand U8996 (N_8996,N_7711,N_7754);
nor U8997 (N_8997,N_7548,N_7887);
or U8998 (N_8998,N_7062,N_7031);
or U8999 (N_8999,N_7269,N_7470);
nor U9000 (N_9000,N_8241,N_8889);
xnor U9001 (N_9001,N_8101,N_8834);
nor U9002 (N_9002,N_8956,N_8179);
or U9003 (N_9003,N_8347,N_8167);
and U9004 (N_9004,N_8686,N_8535);
nand U9005 (N_9005,N_8166,N_8439);
nand U9006 (N_9006,N_8835,N_8692);
and U9007 (N_9007,N_8119,N_8572);
or U9008 (N_9008,N_8429,N_8557);
xnor U9009 (N_9009,N_8622,N_8646);
nor U9010 (N_9010,N_8096,N_8174);
and U9011 (N_9011,N_8123,N_8201);
xor U9012 (N_9012,N_8820,N_8004);
xor U9013 (N_9013,N_8726,N_8163);
nor U9014 (N_9014,N_8003,N_8411);
or U9015 (N_9015,N_8407,N_8814);
nor U9016 (N_9016,N_8006,N_8806);
xor U9017 (N_9017,N_8129,N_8419);
and U9018 (N_9018,N_8478,N_8178);
and U9019 (N_9019,N_8950,N_8769);
and U9020 (N_9020,N_8410,N_8741);
nor U9021 (N_9021,N_8609,N_8306);
nand U9022 (N_9022,N_8169,N_8848);
and U9023 (N_9023,N_8768,N_8857);
and U9024 (N_9024,N_8892,N_8063);
nand U9025 (N_9025,N_8093,N_8332);
and U9026 (N_9026,N_8902,N_8470);
xnor U9027 (N_9027,N_8699,N_8250);
nand U9028 (N_9028,N_8265,N_8369);
xnor U9029 (N_9029,N_8448,N_8222);
or U9030 (N_9030,N_8334,N_8841);
or U9031 (N_9031,N_8349,N_8426);
nor U9032 (N_9032,N_8357,N_8958);
nor U9033 (N_9033,N_8148,N_8711);
or U9034 (N_9034,N_8882,N_8353);
and U9035 (N_9035,N_8531,N_8431);
nand U9036 (N_9036,N_8716,N_8977);
nand U9037 (N_9037,N_8939,N_8420);
xor U9038 (N_9038,N_8521,N_8135);
nand U9039 (N_9039,N_8738,N_8386);
nand U9040 (N_9040,N_8682,N_8099);
nand U9041 (N_9041,N_8731,N_8679);
nand U9042 (N_9042,N_8839,N_8243);
nand U9043 (N_9043,N_8788,N_8136);
or U9044 (N_9044,N_8678,N_8864);
or U9045 (N_9045,N_8971,N_8601);
or U9046 (N_9046,N_8016,N_8913);
or U9047 (N_9047,N_8724,N_8672);
or U9048 (N_9048,N_8229,N_8967);
or U9049 (N_9049,N_8673,N_8651);
or U9050 (N_9050,N_8271,N_8295);
or U9051 (N_9051,N_8712,N_8563);
xnor U9052 (N_9052,N_8255,N_8638);
or U9053 (N_9053,N_8631,N_8746);
xor U9054 (N_9054,N_8773,N_8995);
xor U9055 (N_9055,N_8213,N_8268);
nand U9056 (N_9056,N_8514,N_8182);
nor U9057 (N_9057,N_8062,N_8813);
or U9058 (N_9058,N_8574,N_8454);
or U9059 (N_9059,N_8542,N_8970);
nor U9060 (N_9060,N_8309,N_8816);
xor U9061 (N_9061,N_8840,N_8377);
nand U9062 (N_9062,N_8888,N_8954);
nor U9063 (N_9063,N_8367,N_8885);
or U9064 (N_9064,N_8031,N_8983);
and U9065 (N_9065,N_8056,N_8641);
nor U9066 (N_9066,N_8088,N_8170);
nor U9067 (N_9067,N_8125,N_8138);
nor U9068 (N_9068,N_8078,N_8636);
xor U9069 (N_9069,N_8903,N_8482);
and U9070 (N_9070,N_8073,N_8160);
and U9071 (N_9071,N_8851,N_8727);
nand U9072 (N_9072,N_8149,N_8610);
or U9073 (N_9073,N_8628,N_8378);
and U9074 (N_9074,N_8822,N_8336);
xor U9075 (N_9075,N_8126,N_8944);
nand U9076 (N_9076,N_8674,N_8748);
and U9077 (N_9077,N_8142,N_8914);
nor U9078 (N_9078,N_8952,N_8918);
xnor U9079 (N_9079,N_8035,N_8931);
or U9080 (N_9080,N_8786,N_8547);
xnor U9081 (N_9081,N_8489,N_8462);
nor U9082 (N_9082,N_8591,N_8934);
nand U9083 (N_9083,N_8210,N_8643);
and U9084 (N_9084,N_8779,N_8592);
xor U9085 (N_9085,N_8249,N_8577);
and U9086 (N_9086,N_8463,N_8024);
xnor U9087 (N_9087,N_8204,N_8013);
nand U9088 (N_9088,N_8171,N_8141);
nor U9089 (N_9089,N_8460,N_8758);
nor U9090 (N_9090,N_8272,N_8642);
nand U9091 (N_9091,N_8040,N_8286);
nor U9092 (N_9092,N_8373,N_8434);
and U9093 (N_9093,N_8812,N_8085);
or U9094 (N_9094,N_8940,N_8886);
xnor U9095 (N_9095,N_8270,N_8365);
xor U9096 (N_9096,N_8059,N_8630);
and U9097 (N_9097,N_8790,N_8703);
and U9098 (N_9098,N_8384,N_8767);
nand U9099 (N_9099,N_8134,N_8990);
nor U9100 (N_9100,N_8202,N_8621);
and U9101 (N_9101,N_8856,N_8963);
nand U9102 (N_9102,N_8875,N_8829);
nand U9103 (N_9103,N_8067,N_8828);
and U9104 (N_9104,N_8831,N_8394);
and U9105 (N_9105,N_8528,N_8484);
or U9106 (N_9106,N_8909,N_8754);
or U9107 (N_9107,N_8810,N_8915);
nand U9108 (N_9108,N_8140,N_8261);
and U9109 (N_9109,N_8038,N_8897);
nor U9110 (N_9110,N_8865,N_8842);
nand U9111 (N_9111,N_8433,N_8957);
nand U9112 (N_9112,N_8532,N_8804);
xnor U9113 (N_9113,N_8105,N_8663);
nor U9114 (N_9114,N_8916,N_8743);
nand U9115 (N_9115,N_8449,N_8198);
nor U9116 (N_9116,N_8154,N_8020);
nor U9117 (N_9117,N_8304,N_8879);
xnor U9118 (N_9118,N_8186,N_8089);
and U9119 (N_9119,N_8193,N_8965);
xnor U9120 (N_9120,N_8279,N_8736);
or U9121 (N_9121,N_8585,N_8240);
xor U9122 (N_9122,N_8799,N_8668);
nand U9123 (N_9123,N_8147,N_8504);
and U9124 (N_9124,N_8905,N_8706);
nand U9125 (N_9125,N_8280,N_8273);
or U9126 (N_9126,N_8285,N_8849);
or U9127 (N_9127,N_8103,N_8553);
xor U9128 (N_9128,N_8620,N_8608);
nand U9129 (N_9129,N_8978,N_8314);
xnor U9130 (N_9130,N_8069,N_8480);
or U9131 (N_9131,N_8092,N_8298);
and U9132 (N_9132,N_8032,N_8007);
nand U9133 (N_9133,N_8765,N_8570);
or U9134 (N_9134,N_8108,N_8595);
nand U9135 (N_9135,N_8605,N_8606);
and U9136 (N_9136,N_8614,N_8759);
or U9137 (N_9137,N_8122,N_8805);
nor U9138 (N_9138,N_8556,N_8308);
nand U9139 (N_9139,N_8029,N_8517);
xnor U9140 (N_9140,N_8825,N_8361);
or U9141 (N_9141,N_8852,N_8742);
nor U9142 (N_9142,N_8127,N_8284);
nor U9143 (N_9143,N_8991,N_8391);
or U9144 (N_9144,N_8720,N_8387);
xor U9145 (N_9145,N_8132,N_8018);
xnor U9146 (N_9146,N_8499,N_8869);
and U9147 (N_9147,N_8729,N_8143);
and U9148 (N_9148,N_8060,N_8569);
nand U9149 (N_9149,N_8095,N_8015);
xor U9150 (N_9150,N_8087,N_8675);
nand U9151 (N_9151,N_8259,N_8587);
or U9152 (N_9152,N_8844,N_8988);
nor U9153 (N_9153,N_8113,N_8581);
or U9154 (N_9154,N_8576,N_8305);
and U9155 (N_9155,N_8333,N_8486);
nand U9156 (N_9156,N_8872,N_8156);
and U9157 (N_9157,N_8976,N_8926);
or U9158 (N_9158,N_8231,N_8248);
and U9159 (N_9159,N_8502,N_8091);
nor U9160 (N_9160,N_8074,N_8492);
xnor U9161 (N_9161,N_8066,N_8026);
and U9162 (N_9162,N_8982,N_8808);
nand U9163 (N_9163,N_8055,N_8941);
nand U9164 (N_9164,N_8838,N_8946);
xnor U9165 (N_9165,N_8511,N_8766);
nor U9166 (N_9166,N_8802,N_8413);
nand U9167 (N_9167,N_8194,N_8968);
or U9168 (N_9168,N_8697,N_8320);
xnor U9169 (N_9169,N_8552,N_8770);
and U9170 (N_9170,N_8269,N_8847);
nand U9171 (N_9171,N_8604,N_8155);
nand U9172 (N_9172,N_8145,N_8376);
xor U9173 (N_9173,N_8153,N_8760);
nand U9174 (N_9174,N_8818,N_8562);
nand U9175 (N_9175,N_8447,N_8942);
and U9176 (N_9176,N_8870,N_8104);
and U9177 (N_9177,N_8709,N_8393);
or U9178 (N_9178,N_8246,N_8961);
nor U9179 (N_9179,N_8012,N_8263);
xor U9180 (N_9180,N_8588,N_8212);
nand U9181 (N_9181,N_8100,N_8501);
nor U9182 (N_9182,N_8477,N_8745);
xor U9183 (N_9183,N_8516,N_8177);
xnor U9184 (N_9184,N_8803,N_8874);
nand U9185 (N_9185,N_8043,N_8625);
nand U9186 (N_9186,N_8283,N_8560);
nor U9187 (N_9187,N_8589,N_8415);
nand U9188 (N_9188,N_8654,N_8649);
nand U9189 (N_9189,N_8948,N_8901);
nor U9190 (N_9190,N_8994,N_8809);
and U9191 (N_9191,N_8019,N_8695);
nor U9192 (N_9192,N_8493,N_8761);
or U9193 (N_9193,N_8986,N_8900);
nand U9194 (N_9194,N_8301,N_8371);
or U9195 (N_9195,N_8262,N_8000);
or U9196 (N_9196,N_8685,N_8208);
or U9197 (N_9197,N_8680,N_8181);
and U9198 (N_9198,N_8039,N_8877);
xor U9199 (N_9199,N_8302,N_8794);
xnor U9200 (N_9200,N_8432,N_8054);
xnor U9201 (N_9201,N_8190,N_8688);
or U9202 (N_9202,N_8500,N_8467);
xnor U9203 (N_9203,N_8616,N_8070);
xor U9204 (N_9204,N_8352,N_8236);
or U9205 (N_9205,N_8498,N_8564);
and U9206 (N_9206,N_8076,N_8634);
nand U9207 (N_9207,N_8597,N_8853);
xor U9208 (N_9208,N_8701,N_8833);
nor U9209 (N_9209,N_8951,N_8922);
nor U9210 (N_9210,N_8356,N_8795);
or U9211 (N_9211,N_8578,N_8519);
and U9212 (N_9212,N_8859,N_8188);
nand U9213 (N_9213,N_8895,N_8645);
and U9214 (N_9214,N_8893,N_8996);
and U9215 (N_9215,N_8910,N_8550);
xnor U9216 (N_9216,N_8217,N_8526);
and U9217 (N_9217,N_8081,N_8929);
xnor U9218 (N_9218,N_8571,N_8200);
xnor U9219 (N_9219,N_8730,N_8549);
or U9220 (N_9220,N_8811,N_8666);
nand U9221 (N_9221,N_8107,N_8121);
nand U9222 (N_9222,N_8962,N_8707);
nand U9223 (N_9223,N_8536,N_8771);
and U9224 (N_9224,N_8586,N_8600);
nor U9225 (N_9225,N_8021,N_8216);
and U9226 (N_9226,N_8529,N_8046);
or U9227 (N_9227,N_8254,N_8704);
nand U9228 (N_9228,N_8281,N_8800);
nor U9229 (N_9229,N_8339,N_8045);
nand U9230 (N_9230,N_8647,N_8894);
xor U9231 (N_9231,N_8209,N_8331);
nor U9232 (N_9232,N_8323,N_8436);
and U9233 (N_9233,N_8541,N_8797);
and U9234 (N_9234,N_8580,N_8445);
nor U9235 (N_9235,N_8955,N_8772);
nand U9236 (N_9236,N_8251,N_8010);
or U9237 (N_9237,N_8898,N_8617);
and U9238 (N_9238,N_8278,N_8774);
and U9239 (N_9239,N_8947,N_8162);
and U9240 (N_9240,N_8335,N_8400);
nand U9241 (N_9241,N_8830,N_8165);
nand U9242 (N_9242,N_8094,N_8739);
and U9243 (N_9243,N_8530,N_8418);
nand U9244 (N_9244,N_8777,N_8052);
nor U9245 (N_9245,N_8923,N_8025);
xnor U9246 (N_9246,N_8057,N_8292);
xnor U9247 (N_9247,N_8446,N_8881);
nand U9248 (N_9248,N_8997,N_8382);
xor U9249 (N_9249,N_8972,N_8466);
or U9250 (N_9250,N_8253,N_8611);
nor U9251 (N_9251,N_8317,N_8753);
or U9252 (N_9252,N_8061,N_8161);
or U9253 (N_9253,N_8047,N_8363);
xor U9254 (N_9254,N_8086,N_8664);
xor U9255 (N_9255,N_8257,N_8546);
nor U9256 (N_9256,N_8681,N_8311);
nor U9257 (N_9257,N_8884,N_8346);
and U9258 (N_9258,N_8959,N_8490);
and U9259 (N_9259,N_8694,N_8689);
xor U9260 (N_9260,N_8868,N_8206);
xnor U9261 (N_9261,N_8896,N_8408);
nor U9262 (N_9262,N_8544,N_8687);
nand U9263 (N_9263,N_8291,N_8303);
and U9264 (N_9264,N_8505,N_8538);
nand U9265 (N_9265,N_8033,N_8583);
xnor U9266 (N_9266,N_8602,N_8474);
xnor U9267 (N_9267,N_8041,N_8590);
xnor U9268 (N_9268,N_8639,N_8110);
nand U9269 (N_9269,N_8599,N_8487);
xor U9270 (N_9270,N_8423,N_8203);
or U9271 (N_9271,N_8579,N_8328);
xor U9272 (N_9272,N_8476,N_8082);
nor U9273 (N_9273,N_8215,N_8315);
and U9274 (N_9274,N_8551,N_8665);
nand U9275 (N_9275,N_8388,N_8558);
and U9276 (N_9276,N_8329,N_8710);
nor U9277 (N_9277,N_8722,N_8960);
xor U9278 (N_9278,N_8798,N_8780);
nor U9279 (N_9279,N_8824,N_8455);
nor U9280 (N_9280,N_8801,N_8044);
or U9281 (N_9281,N_8998,N_8366);
nor U9282 (N_9282,N_8219,N_8992);
xor U9283 (N_9283,N_8949,N_8252);
nand U9284 (N_9284,N_8933,N_8392);
or U9285 (N_9285,N_8930,N_8150);
xnor U9286 (N_9286,N_8533,N_8290);
and U9287 (N_9287,N_8379,N_8380);
or U9288 (N_9288,N_8027,N_8507);
nand U9289 (N_9289,N_8691,N_8633);
nand U9290 (N_9290,N_8719,N_8593);
nor U9291 (N_9291,N_8435,N_8358);
nor U9292 (N_9292,N_8444,N_8050);
nor U9293 (N_9293,N_8227,N_8116);
and U9294 (N_9294,N_8974,N_8464);
and U9295 (N_9295,N_8539,N_8655);
and U9296 (N_9296,N_8921,N_8566);
or U9297 (N_9297,N_8624,N_8428);
and U9298 (N_9298,N_8827,N_8629);
nand U9299 (N_9299,N_8383,N_8671);
nor U9300 (N_9300,N_8935,N_8226);
or U9301 (N_9301,N_8168,N_8635);
and U9302 (N_9302,N_8266,N_8778);
nor U9303 (N_9303,N_8751,N_8028);
or U9304 (N_9304,N_8911,N_8205);
xnor U9305 (N_9305,N_8402,N_8863);
nand U9306 (N_9306,N_8296,N_8855);
or U9307 (N_9307,N_8496,N_8565);
nor U9308 (N_9308,N_8244,N_8164);
nor U9309 (N_9309,N_8071,N_8115);
xnor U9310 (N_9310,N_8659,N_8372);
nand U9311 (N_9311,N_8700,N_8422);
xnor U9312 (N_9312,N_8891,N_8981);
xor U9313 (N_9313,N_8749,N_8937);
and U9314 (N_9314,N_8385,N_8399);
nand U9315 (N_9315,N_8159,N_8065);
xor U9316 (N_9316,N_8485,N_8294);
and U9317 (N_9317,N_8715,N_8669);
or U9318 (N_9318,N_8740,N_8618);
xor U9319 (N_9319,N_8396,N_8503);
or U9320 (N_9320,N_8508,N_8953);
xor U9321 (N_9321,N_8293,N_8008);
nand U9322 (N_9322,N_8737,N_8300);
nor U9323 (N_9323,N_8098,N_8453);
and U9324 (N_9324,N_8404,N_8523);
and U9325 (N_9325,N_8316,N_8427);
nand U9326 (N_9326,N_8696,N_8354);
nand U9327 (N_9327,N_8370,N_8005);
nand U9328 (N_9328,N_8211,N_8999);
nor U9329 (N_9329,N_8932,N_8267);
xor U9330 (N_9330,N_8483,N_8807);
xor U9331 (N_9331,N_8854,N_8693);
xnor U9332 (N_9332,N_8189,N_8648);
or U9333 (N_9333,N_8185,N_8355);
nor U9334 (N_9334,N_8375,N_8979);
and U9335 (N_9335,N_8559,N_8728);
xnor U9336 (N_9336,N_8878,N_8702);
xor U9337 (N_9337,N_8117,N_8661);
or U9338 (N_9338,N_8755,N_8235);
nor U9339 (N_9339,N_8657,N_8796);
xnor U9340 (N_9340,N_8723,N_8175);
or U9341 (N_9341,N_8424,N_8350);
xor U9342 (N_9342,N_8757,N_8318);
nor U9343 (N_9343,N_8573,N_8924);
xnor U9344 (N_9344,N_8525,N_8327);
xnor U9345 (N_9345,N_8792,N_8381);
xnor U9346 (N_9346,N_8360,N_8247);
and U9347 (N_9347,N_8144,N_8718);
or U9348 (N_9348,N_8049,N_8157);
and U9349 (N_9349,N_8130,N_8223);
nand U9350 (N_9350,N_8481,N_8124);
nand U9351 (N_9351,N_8397,N_8491);
xor U9352 (N_9352,N_8890,N_8776);
nand U9353 (N_9353,N_8324,N_8184);
nor U9354 (N_9354,N_8850,N_8058);
xor U9355 (N_9355,N_8139,N_8389);
and U9356 (N_9356,N_8619,N_8936);
nor U9357 (N_9357,N_8907,N_8214);
or U9358 (N_9358,N_8173,N_8456);
nor U9359 (N_9359,N_8919,N_8051);
nand U9360 (N_9360,N_8242,N_8938);
or U9361 (N_9361,N_8543,N_8348);
nor U9362 (N_9362,N_8845,N_8980);
and U9363 (N_9363,N_8465,N_8964);
xnor U9364 (N_9364,N_8555,N_8713);
xor U9365 (N_9365,N_8109,N_8416);
xnor U9366 (N_9366,N_8207,N_8861);
and U9367 (N_9367,N_8826,N_8819);
nand U9368 (N_9368,N_8405,N_8338);
or U9369 (N_9369,N_8783,N_8321);
or U9370 (N_9370,N_8342,N_8943);
nand U9371 (N_9371,N_8866,N_8014);
and U9372 (N_9372,N_8787,N_8112);
xnor U9373 (N_9373,N_8714,N_8858);
and U9374 (N_9374,N_8196,N_8079);
nor U9375 (N_9375,N_8414,N_8920);
nor U9376 (N_9376,N_8345,N_8846);
xnor U9377 (N_9377,N_8417,N_8359);
and U9378 (N_9378,N_8077,N_8734);
nor U9379 (N_9379,N_8183,N_8725);
nor U9380 (N_9380,N_8313,N_8717);
nand U9381 (N_9381,N_8750,N_8471);
nand U9382 (N_9382,N_8684,N_8667);
nor U9383 (N_9383,N_8660,N_8128);
nand U9384 (N_9384,N_8509,N_8191);
nor U9385 (N_9385,N_8756,N_8596);
nor U9386 (N_9386,N_8001,N_8969);
nor U9387 (N_9387,N_8337,N_8945);
or U9388 (N_9388,N_8120,N_8048);
and U9389 (N_9389,N_8537,N_8218);
nand U9390 (N_9390,N_8409,N_8118);
or U9391 (N_9391,N_8002,N_8966);
or U9392 (N_9392,N_8698,N_8036);
nand U9393 (N_9393,N_8258,N_8705);
nor U9394 (N_9394,N_8843,N_8137);
nand U9395 (N_9395,N_8452,N_8662);
nor U9396 (N_9396,N_8322,N_8494);
and U9397 (N_9397,N_8683,N_8022);
nor U9398 (N_9398,N_8437,N_8925);
and U9399 (N_9399,N_8993,N_8518);
and U9400 (N_9400,N_8114,N_8561);
and U9401 (N_9401,N_8495,N_8545);
or U9402 (N_9402,N_8276,N_8042);
nand U9403 (N_9403,N_8899,N_8351);
and U9404 (N_9404,N_8459,N_8823);
xnor U9405 (N_9405,N_8401,N_8195);
or U9406 (N_9406,N_8912,N_8260);
nor U9407 (N_9407,N_8862,N_8904);
xnor U9408 (N_9408,N_8876,N_8199);
and U9409 (N_9409,N_8582,N_8721);
or U9410 (N_9410,N_8747,N_8053);
xnor U9411 (N_9411,N_8017,N_8403);
and U9412 (N_9412,N_8873,N_8009);
or U9413 (N_9413,N_8187,N_8763);
or U9414 (N_9414,N_8228,N_8364);
nor U9415 (N_9415,N_8374,N_8652);
xnor U9416 (N_9416,N_8880,N_8152);
nor U9417 (N_9417,N_8233,N_8412);
and U9418 (N_9418,N_8083,N_8764);
and U9419 (N_9419,N_8330,N_8479);
and U9420 (N_9420,N_8656,N_8612);
nor U9421 (N_9421,N_8817,N_8461);
or U9422 (N_9422,N_8887,N_8821);
nor U9423 (N_9423,N_8837,N_8615);
nand U9424 (N_9424,N_8475,N_8172);
xor U9425 (N_9425,N_8917,N_8438);
nor U9426 (N_9426,N_8232,N_8644);
nor U9427 (N_9427,N_8442,N_8287);
nand U9428 (N_9428,N_8406,N_8744);
xor U9429 (N_9429,N_8245,N_8430);
nand U9430 (N_9430,N_8623,N_8037);
or U9431 (N_9431,N_8928,N_8782);
nor U9432 (N_9432,N_8275,N_8548);
or U9433 (N_9433,N_8472,N_8488);
nor U9434 (N_9434,N_8030,N_8398);
nor U9435 (N_9435,N_8341,N_8594);
nor U9436 (N_9436,N_8282,N_8264);
nor U9437 (N_9437,N_8158,N_8640);
and U9438 (N_9438,N_8784,N_8815);
and U9439 (N_9439,N_8084,N_8762);
or U9440 (N_9440,N_8984,N_8450);
nand U9441 (N_9441,N_8192,N_8584);
nand U9442 (N_9442,N_8225,N_8220);
nor U9443 (N_9443,N_8344,N_8151);
nor U9444 (N_9444,N_8133,N_8515);
and U9445 (N_9445,N_8473,N_8368);
or U9446 (N_9446,N_8575,N_8554);
xor U9447 (N_9447,N_8650,N_8297);
xnor U9448 (N_9448,N_8288,N_8224);
nor U9449 (N_9449,N_8234,N_8627);
or U9450 (N_9450,N_8072,N_8534);
and U9451 (N_9451,N_8908,N_8441);
nor U9452 (N_9452,N_8034,N_8421);
nand U9453 (N_9453,N_8527,N_8064);
nand U9454 (N_9454,N_8326,N_8237);
and U9455 (N_9455,N_8708,N_8732);
or U9456 (N_9456,N_8340,N_8111);
or U9457 (N_9457,N_8607,N_8860);
nand U9458 (N_9458,N_8468,N_8102);
nor U9459 (N_9459,N_8632,N_8927);
or U9460 (N_9460,N_8906,N_8080);
and U9461 (N_9461,N_8319,N_8781);
or U9462 (N_9462,N_8883,N_8513);
and U9463 (N_9463,N_8637,N_8568);
nand U9464 (N_9464,N_8310,N_8146);
and U9465 (N_9465,N_8457,N_8735);
or U9466 (N_9466,N_8512,N_8524);
or U9467 (N_9467,N_8307,N_8097);
xor U9468 (N_9468,N_8299,N_8011);
nor U9469 (N_9469,N_8975,N_8221);
nor U9470 (N_9470,N_8312,N_8598);
nor U9471 (N_9471,N_8670,N_8390);
nor U9472 (N_9472,N_8733,N_8068);
and U9473 (N_9473,N_8469,N_8362);
nand U9474 (N_9474,N_8789,N_8277);
or U9475 (N_9475,N_8775,N_8987);
or U9476 (N_9476,N_8793,N_8090);
and U9477 (N_9477,N_8989,N_8075);
nand U9478 (N_9478,N_8256,N_8510);
nor U9479 (N_9479,N_8613,N_8871);
or U9480 (N_9480,N_8506,N_8867);
nand U9481 (N_9481,N_8131,N_8023);
xnor U9482 (N_9482,N_8690,N_8238);
xor U9483 (N_9483,N_8497,N_8567);
xnor U9484 (N_9484,N_8603,N_8395);
xnor U9485 (N_9485,N_8836,N_8658);
and U9486 (N_9486,N_8106,N_8985);
and U9487 (N_9487,N_8676,N_8197);
and U9488 (N_9488,N_8520,N_8522);
and U9489 (N_9489,N_8425,N_8791);
nand U9490 (N_9490,N_8540,N_8325);
nand U9491 (N_9491,N_8458,N_8440);
nor U9492 (N_9492,N_8752,N_8239);
nor U9493 (N_9493,N_8626,N_8451);
nand U9494 (N_9494,N_8443,N_8343);
nand U9495 (N_9495,N_8180,N_8653);
xnor U9496 (N_9496,N_8176,N_8274);
xor U9497 (N_9497,N_8230,N_8973);
xor U9498 (N_9498,N_8785,N_8677);
and U9499 (N_9499,N_8832,N_8289);
xor U9500 (N_9500,N_8808,N_8714);
xnor U9501 (N_9501,N_8772,N_8893);
and U9502 (N_9502,N_8558,N_8954);
or U9503 (N_9503,N_8879,N_8835);
and U9504 (N_9504,N_8432,N_8575);
nor U9505 (N_9505,N_8571,N_8875);
nor U9506 (N_9506,N_8121,N_8987);
or U9507 (N_9507,N_8333,N_8100);
nor U9508 (N_9508,N_8815,N_8067);
nand U9509 (N_9509,N_8435,N_8015);
nor U9510 (N_9510,N_8042,N_8625);
or U9511 (N_9511,N_8990,N_8052);
nor U9512 (N_9512,N_8324,N_8141);
xnor U9513 (N_9513,N_8793,N_8939);
xnor U9514 (N_9514,N_8297,N_8262);
and U9515 (N_9515,N_8299,N_8350);
and U9516 (N_9516,N_8708,N_8460);
xor U9517 (N_9517,N_8096,N_8496);
or U9518 (N_9518,N_8623,N_8502);
xnor U9519 (N_9519,N_8004,N_8950);
nor U9520 (N_9520,N_8450,N_8735);
nand U9521 (N_9521,N_8475,N_8964);
xnor U9522 (N_9522,N_8767,N_8137);
and U9523 (N_9523,N_8706,N_8683);
or U9524 (N_9524,N_8331,N_8531);
and U9525 (N_9525,N_8796,N_8418);
or U9526 (N_9526,N_8955,N_8813);
nor U9527 (N_9527,N_8762,N_8637);
and U9528 (N_9528,N_8613,N_8299);
nor U9529 (N_9529,N_8036,N_8281);
xnor U9530 (N_9530,N_8466,N_8714);
nor U9531 (N_9531,N_8596,N_8331);
or U9532 (N_9532,N_8090,N_8986);
xnor U9533 (N_9533,N_8642,N_8005);
xnor U9534 (N_9534,N_8269,N_8654);
nand U9535 (N_9535,N_8367,N_8432);
or U9536 (N_9536,N_8723,N_8883);
xnor U9537 (N_9537,N_8168,N_8576);
or U9538 (N_9538,N_8054,N_8908);
and U9539 (N_9539,N_8007,N_8378);
nand U9540 (N_9540,N_8034,N_8127);
xnor U9541 (N_9541,N_8698,N_8352);
nor U9542 (N_9542,N_8621,N_8005);
xor U9543 (N_9543,N_8021,N_8400);
xnor U9544 (N_9544,N_8536,N_8156);
and U9545 (N_9545,N_8422,N_8981);
or U9546 (N_9546,N_8914,N_8834);
or U9547 (N_9547,N_8423,N_8327);
and U9548 (N_9548,N_8199,N_8337);
xnor U9549 (N_9549,N_8011,N_8427);
and U9550 (N_9550,N_8184,N_8427);
nor U9551 (N_9551,N_8303,N_8200);
xnor U9552 (N_9552,N_8649,N_8552);
xnor U9553 (N_9553,N_8832,N_8083);
and U9554 (N_9554,N_8926,N_8183);
and U9555 (N_9555,N_8466,N_8040);
or U9556 (N_9556,N_8176,N_8877);
nor U9557 (N_9557,N_8740,N_8987);
or U9558 (N_9558,N_8947,N_8451);
nand U9559 (N_9559,N_8070,N_8976);
xnor U9560 (N_9560,N_8239,N_8829);
nor U9561 (N_9561,N_8440,N_8397);
and U9562 (N_9562,N_8162,N_8477);
or U9563 (N_9563,N_8125,N_8593);
xnor U9564 (N_9564,N_8417,N_8807);
nand U9565 (N_9565,N_8879,N_8854);
xnor U9566 (N_9566,N_8567,N_8628);
or U9567 (N_9567,N_8790,N_8135);
nand U9568 (N_9568,N_8827,N_8508);
and U9569 (N_9569,N_8250,N_8434);
xnor U9570 (N_9570,N_8904,N_8344);
and U9571 (N_9571,N_8963,N_8112);
nand U9572 (N_9572,N_8310,N_8847);
xnor U9573 (N_9573,N_8410,N_8789);
nand U9574 (N_9574,N_8623,N_8071);
and U9575 (N_9575,N_8503,N_8384);
or U9576 (N_9576,N_8610,N_8005);
nand U9577 (N_9577,N_8639,N_8907);
xnor U9578 (N_9578,N_8305,N_8720);
or U9579 (N_9579,N_8255,N_8811);
xnor U9580 (N_9580,N_8440,N_8133);
and U9581 (N_9581,N_8769,N_8459);
nand U9582 (N_9582,N_8898,N_8427);
nor U9583 (N_9583,N_8173,N_8411);
nor U9584 (N_9584,N_8883,N_8031);
and U9585 (N_9585,N_8454,N_8698);
or U9586 (N_9586,N_8904,N_8383);
and U9587 (N_9587,N_8047,N_8116);
nor U9588 (N_9588,N_8730,N_8755);
nand U9589 (N_9589,N_8833,N_8150);
or U9590 (N_9590,N_8652,N_8542);
or U9591 (N_9591,N_8896,N_8607);
or U9592 (N_9592,N_8866,N_8879);
nor U9593 (N_9593,N_8014,N_8741);
nand U9594 (N_9594,N_8972,N_8080);
nor U9595 (N_9595,N_8093,N_8963);
or U9596 (N_9596,N_8057,N_8275);
and U9597 (N_9597,N_8436,N_8096);
nor U9598 (N_9598,N_8138,N_8794);
nand U9599 (N_9599,N_8214,N_8697);
nand U9600 (N_9600,N_8998,N_8655);
xor U9601 (N_9601,N_8988,N_8353);
nor U9602 (N_9602,N_8514,N_8052);
and U9603 (N_9603,N_8222,N_8979);
xnor U9604 (N_9604,N_8547,N_8470);
xnor U9605 (N_9605,N_8297,N_8502);
and U9606 (N_9606,N_8825,N_8556);
nor U9607 (N_9607,N_8136,N_8825);
or U9608 (N_9608,N_8103,N_8702);
nand U9609 (N_9609,N_8964,N_8164);
xnor U9610 (N_9610,N_8515,N_8699);
xor U9611 (N_9611,N_8440,N_8960);
nand U9612 (N_9612,N_8959,N_8525);
nand U9613 (N_9613,N_8114,N_8461);
nand U9614 (N_9614,N_8845,N_8399);
or U9615 (N_9615,N_8856,N_8030);
nor U9616 (N_9616,N_8000,N_8332);
nor U9617 (N_9617,N_8534,N_8330);
xnor U9618 (N_9618,N_8665,N_8427);
or U9619 (N_9619,N_8245,N_8158);
and U9620 (N_9620,N_8417,N_8928);
nand U9621 (N_9621,N_8431,N_8790);
or U9622 (N_9622,N_8766,N_8543);
xnor U9623 (N_9623,N_8677,N_8060);
nand U9624 (N_9624,N_8149,N_8409);
nor U9625 (N_9625,N_8564,N_8207);
or U9626 (N_9626,N_8785,N_8512);
nor U9627 (N_9627,N_8896,N_8048);
or U9628 (N_9628,N_8694,N_8893);
or U9629 (N_9629,N_8649,N_8228);
nor U9630 (N_9630,N_8499,N_8716);
xnor U9631 (N_9631,N_8786,N_8879);
or U9632 (N_9632,N_8365,N_8011);
nand U9633 (N_9633,N_8143,N_8592);
nor U9634 (N_9634,N_8491,N_8898);
nand U9635 (N_9635,N_8433,N_8626);
and U9636 (N_9636,N_8765,N_8306);
xor U9637 (N_9637,N_8680,N_8869);
and U9638 (N_9638,N_8290,N_8226);
nand U9639 (N_9639,N_8455,N_8988);
and U9640 (N_9640,N_8301,N_8665);
nor U9641 (N_9641,N_8860,N_8193);
nor U9642 (N_9642,N_8562,N_8493);
nor U9643 (N_9643,N_8811,N_8745);
or U9644 (N_9644,N_8561,N_8804);
nor U9645 (N_9645,N_8715,N_8764);
and U9646 (N_9646,N_8782,N_8476);
and U9647 (N_9647,N_8224,N_8514);
and U9648 (N_9648,N_8051,N_8312);
and U9649 (N_9649,N_8798,N_8905);
or U9650 (N_9650,N_8091,N_8988);
and U9651 (N_9651,N_8232,N_8224);
nand U9652 (N_9652,N_8834,N_8337);
and U9653 (N_9653,N_8591,N_8788);
nand U9654 (N_9654,N_8750,N_8295);
or U9655 (N_9655,N_8204,N_8225);
nor U9656 (N_9656,N_8750,N_8764);
xnor U9657 (N_9657,N_8411,N_8422);
xnor U9658 (N_9658,N_8085,N_8005);
or U9659 (N_9659,N_8098,N_8363);
and U9660 (N_9660,N_8443,N_8981);
nand U9661 (N_9661,N_8799,N_8194);
nor U9662 (N_9662,N_8603,N_8244);
nand U9663 (N_9663,N_8042,N_8819);
xor U9664 (N_9664,N_8118,N_8307);
nand U9665 (N_9665,N_8518,N_8448);
nand U9666 (N_9666,N_8426,N_8589);
and U9667 (N_9667,N_8937,N_8350);
xor U9668 (N_9668,N_8741,N_8703);
nand U9669 (N_9669,N_8867,N_8537);
nor U9670 (N_9670,N_8068,N_8642);
nand U9671 (N_9671,N_8648,N_8090);
and U9672 (N_9672,N_8517,N_8879);
nand U9673 (N_9673,N_8942,N_8725);
nor U9674 (N_9674,N_8785,N_8850);
or U9675 (N_9675,N_8677,N_8697);
nand U9676 (N_9676,N_8262,N_8908);
and U9677 (N_9677,N_8256,N_8571);
nand U9678 (N_9678,N_8099,N_8211);
nand U9679 (N_9679,N_8411,N_8684);
or U9680 (N_9680,N_8761,N_8133);
nand U9681 (N_9681,N_8974,N_8103);
and U9682 (N_9682,N_8394,N_8095);
or U9683 (N_9683,N_8051,N_8588);
and U9684 (N_9684,N_8422,N_8294);
nor U9685 (N_9685,N_8617,N_8179);
or U9686 (N_9686,N_8276,N_8421);
xnor U9687 (N_9687,N_8843,N_8116);
nand U9688 (N_9688,N_8535,N_8945);
nand U9689 (N_9689,N_8691,N_8844);
xnor U9690 (N_9690,N_8490,N_8155);
and U9691 (N_9691,N_8527,N_8343);
xor U9692 (N_9692,N_8039,N_8883);
xor U9693 (N_9693,N_8607,N_8321);
or U9694 (N_9694,N_8119,N_8320);
and U9695 (N_9695,N_8328,N_8686);
nand U9696 (N_9696,N_8285,N_8019);
and U9697 (N_9697,N_8415,N_8446);
xnor U9698 (N_9698,N_8207,N_8373);
and U9699 (N_9699,N_8635,N_8014);
xnor U9700 (N_9700,N_8666,N_8915);
or U9701 (N_9701,N_8760,N_8344);
or U9702 (N_9702,N_8713,N_8804);
and U9703 (N_9703,N_8910,N_8856);
nor U9704 (N_9704,N_8865,N_8724);
and U9705 (N_9705,N_8294,N_8577);
or U9706 (N_9706,N_8733,N_8028);
nor U9707 (N_9707,N_8899,N_8132);
and U9708 (N_9708,N_8577,N_8381);
or U9709 (N_9709,N_8670,N_8292);
or U9710 (N_9710,N_8558,N_8455);
nand U9711 (N_9711,N_8793,N_8224);
xor U9712 (N_9712,N_8792,N_8378);
and U9713 (N_9713,N_8182,N_8336);
and U9714 (N_9714,N_8081,N_8342);
xnor U9715 (N_9715,N_8055,N_8847);
or U9716 (N_9716,N_8481,N_8546);
nor U9717 (N_9717,N_8988,N_8181);
and U9718 (N_9718,N_8287,N_8345);
and U9719 (N_9719,N_8773,N_8826);
or U9720 (N_9720,N_8103,N_8447);
xnor U9721 (N_9721,N_8249,N_8578);
or U9722 (N_9722,N_8900,N_8767);
or U9723 (N_9723,N_8966,N_8951);
or U9724 (N_9724,N_8542,N_8769);
or U9725 (N_9725,N_8719,N_8810);
or U9726 (N_9726,N_8099,N_8056);
nand U9727 (N_9727,N_8750,N_8027);
or U9728 (N_9728,N_8642,N_8950);
xor U9729 (N_9729,N_8527,N_8339);
and U9730 (N_9730,N_8493,N_8770);
nor U9731 (N_9731,N_8008,N_8470);
or U9732 (N_9732,N_8513,N_8555);
nand U9733 (N_9733,N_8697,N_8798);
or U9734 (N_9734,N_8718,N_8621);
xor U9735 (N_9735,N_8737,N_8061);
nor U9736 (N_9736,N_8472,N_8492);
and U9737 (N_9737,N_8734,N_8186);
and U9738 (N_9738,N_8973,N_8703);
and U9739 (N_9739,N_8049,N_8367);
or U9740 (N_9740,N_8878,N_8112);
xor U9741 (N_9741,N_8404,N_8690);
nand U9742 (N_9742,N_8007,N_8147);
xnor U9743 (N_9743,N_8238,N_8039);
xnor U9744 (N_9744,N_8466,N_8178);
and U9745 (N_9745,N_8375,N_8661);
or U9746 (N_9746,N_8797,N_8795);
nand U9747 (N_9747,N_8139,N_8419);
nor U9748 (N_9748,N_8494,N_8818);
nor U9749 (N_9749,N_8670,N_8344);
and U9750 (N_9750,N_8388,N_8101);
nor U9751 (N_9751,N_8256,N_8144);
nand U9752 (N_9752,N_8465,N_8133);
nor U9753 (N_9753,N_8518,N_8229);
nand U9754 (N_9754,N_8724,N_8539);
nor U9755 (N_9755,N_8416,N_8108);
or U9756 (N_9756,N_8434,N_8252);
nand U9757 (N_9757,N_8919,N_8938);
or U9758 (N_9758,N_8406,N_8598);
nand U9759 (N_9759,N_8814,N_8742);
nor U9760 (N_9760,N_8899,N_8595);
nand U9761 (N_9761,N_8205,N_8667);
or U9762 (N_9762,N_8005,N_8593);
nand U9763 (N_9763,N_8785,N_8971);
and U9764 (N_9764,N_8788,N_8054);
nor U9765 (N_9765,N_8574,N_8402);
nor U9766 (N_9766,N_8625,N_8511);
nand U9767 (N_9767,N_8887,N_8551);
or U9768 (N_9768,N_8938,N_8294);
nand U9769 (N_9769,N_8581,N_8231);
nor U9770 (N_9770,N_8616,N_8906);
nand U9771 (N_9771,N_8900,N_8785);
nand U9772 (N_9772,N_8660,N_8546);
nand U9773 (N_9773,N_8662,N_8787);
nor U9774 (N_9774,N_8853,N_8633);
xnor U9775 (N_9775,N_8214,N_8572);
xnor U9776 (N_9776,N_8486,N_8563);
and U9777 (N_9777,N_8519,N_8143);
xnor U9778 (N_9778,N_8242,N_8563);
nor U9779 (N_9779,N_8106,N_8794);
xor U9780 (N_9780,N_8632,N_8407);
or U9781 (N_9781,N_8319,N_8079);
nand U9782 (N_9782,N_8198,N_8357);
or U9783 (N_9783,N_8293,N_8781);
xor U9784 (N_9784,N_8038,N_8504);
nand U9785 (N_9785,N_8816,N_8457);
xnor U9786 (N_9786,N_8791,N_8751);
nor U9787 (N_9787,N_8427,N_8994);
and U9788 (N_9788,N_8589,N_8339);
or U9789 (N_9789,N_8776,N_8357);
and U9790 (N_9790,N_8813,N_8817);
or U9791 (N_9791,N_8932,N_8170);
and U9792 (N_9792,N_8017,N_8348);
xor U9793 (N_9793,N_8949,N_8621);
xnor U9794 (N_9794,N_8255,N_8988);
and U9795 (N_9795,N_8995,N_8670);
and U9796 (N_9796,N_8586,N_8884);
nand U9797 (N_9797,N_8380,N_8668);
or U9798 (N_9798,N_8544,N_8703);
nand U9799 (N_9799,N_8464,N_8327);
xnor U9800 (N_9800,N_8437,N_8794);
nor U9801 (N_9801,N_8776,N_8589);
xnor U9802 (N_9802,N_8800,N_8252);
nor U9803 (N_9803,N_8571,N_8194);
or U9804 (N_9804,N_8879,N_8862);
nor U9805 (N_9805,N_8839,N_8548);
nor U9806 (N_9806,N_8497,N_8082);
or U9807 (N_9807,N_8194,N_8986);
nor U9808 (N_9808,N_8414,N_8717);
nand U9809 (N_9809,N_8687,N_8374);
or U9810 (N_9810,N_8130,N_8726);
xnor U9811 (N_9811,N_8060,N_8178);
and U9812 (N_9812,N_8939,N_8745);
and U9813 (N_9813,N_8747,N_8284);
or U9814 (N_9814,N_8866,N_8768);
or U9815 (N_9815,N_8070,N_8157);
nand U9816 (N_9816,N_8461,N_8058);
nand U9817 (N_9817,N_8930,N_8891);
nor U9818 (N_9818,N_8166,N_8767);
and U9819 (N_9819,N_8499,N_8545);
xor U9820 (N_9820,N_8889,N_8972);
nor U9821 (N_9821,N_8228,N_8441);
nor U9822 (N_9822,N_8365,N_8172);
and U9823 (N_9823,N_8339,N_8879);
or U9824 (N_9824,N_8942,N_8936);
nand U9825 (N_9825,N_8059,N_8691);
nand U9826 (N_9826,N_8093,N_8469);
nand U9827 (N_9827,N_8201,N_8567);
nand U9828 (N_9828,N_8629,N_8883);
xnor U9829 (N_9829,N_8233,N_8616);
nand U9830 (N_9830,N_8836,N_8968);
and U9831 (N_9831,N_8017,N_8976);
nor U9832 (N_9832,N_8326,N_8914);
and U9833 (N_9833,N_8659,N_8468);
and U9834 (N_9834,N_8480,N_8052);
nor U9835 (N_9835,N_8036,N_8136);
nor U9836 (N_9836,N_8294,N_8352);
or U9837 (N_9837,N_8977,N_8246);
nand U9838 (N_9838,N_8076,N_8085);
nor U9839 (N_9839,N_8999,N_8245);
xnor U9840 (N_9840,N_8381,N_8956);
nor U9841 (N_9841,N_8578,N_8759);
and U9842 (N_9842,N_8046,N_8566);
xor U9843 (N_9843,N_8503,N_8671);
xnor U9844 (N_9844,N_8275,N_8056);
nand U9845 (N_9845,N_8337,N_8258);
and U9846 (N_9846,N_8982,N_8526);
xor U9847 (N_9847,N_8419,N_8423);
or U9848 (N_9848,N_8506,N_8437);
nand U9849 (N_9849,N_8717,N_8211);
xor U9850 (N_9850,N_8361,N_8895);
xor U9851 (N_9851,N_8417,N_8108);
nand U9852 (N_9852,N_8318,N_8302);
or U9853 (N_9853,N_8003,N_8242);
nand U9854 (N_9854,N_8060,N_8249);
and U9855 (N_9855,N_8342,N_8827);
nor U9856 (N_9856,N_8563,N_8848);
xor U9857 (N_9857,N_8838,N_8209);
nor U9858 (N_9858,N_8062,N_8511);
nor U9859 (N_9859,N_8946,N_8055);
xnor U9860 (N_9860,N_8746,N_8538);
xnor U9861 (N_9861,N_8421,N_8797);
and U9862 (N_9862,N_8263,N_8068);
and U9863 (N_9863,N_8388,N_8860);
nand U9864 (N_9864,N_8702,N_8286);
xnor U9865 (N_9865,N_8542,N_8029);
nand U9866 (N_9866,N_8646,N_8308);
and U9867 (N_9867,N_8178,N_8268);
nand U9868 (N_9868,N_8146,N_8136);
or U9869 (N_9869,N_8383,N_8443);
and U9870 (N_9870,N_8788,N_8172);
and U9871 (N_9871,N_8992,N_8848);
and U9872 (N_9872,N_8521,N_8176);
or U9873 (N_9873,N_8509,N_8373);
nor U9874 (N_9874,N_8646,N_8218);
or U9875 (N_9875,N_8430,N_8008);
nor U9876 (N_9876,N_8507,N_8437);
and U9877 (N_9877,N_8193,N_8214);
nand U9878 (N_9878,N_8106,N_8956);
and U9879 (N_9879,N_8312,N_8434);
or U9880 (N_9880,N_8968,N_8307);
or U9881 (N_9881,N_8169,N_8724);
nand U9882 (N_9882,N_8919,N_8959);
or U9883 (N_9883,N_8968,N_8985);
nor U9884 (N_9884,N_8587,N_8443);
or U9885 (N_9885,N_8759,N_8968);
xor U9886 (N_9886,N_8434,N_8301);
and U9887 (N_9887,N_8826,N_8694);
and U9888 (N_9888,N_8699,N_8669);
or U9889 (N_9889,N_8898,N_8853);
nand U9890 (N_9890,N_8859,N_8540);
nand U9891 (N_9891,N_8685,N_8178);
nor U9892 (N_9892,N_8256,N_8299);
and U9893 (N_9893,N_8467,N_8419);
xnor U9894 (N_9894,N_8834,N_8187);
or U9895 (N_9895,N_8659,N_8950);
and U9896 (N_9896,N_8570,N_8426);
and U9897 (N_9897,N_8027,N_8140);
nor U9898 (N_9898,N_8816,N_8234);
or U9899 (N_9899,N_8863,N_8912);
xor U9900 (N_9900,N_8733,N_8154);
and U9901 (N_9901,N_8895,N_8019);
or U9902 (N_9902,N_8301,N_8118);
xor U9903 (N_9903,N_8165,N_8539);
xnor U9904 (N_9904,N_8190,N_8249);
nand U9905 (N_9905,N_8341,N_8787);
nor U9906 (N_9906,N_8716,N_8754);
nand U9907 (N_9907,N_8781,N_8211);
or U9908 (N_9908,N_8612,N_8601);
or U9909 (N_9909,N_8405,N_8677);
nand U9910 (N_9910,N_8665,N_8524);
nor U9911 (N_9911,N_8430,N_8664);
or U9912 (N_9912,N_8735,N_8923);
xnor U9913 (N_9913,N_8659,N_8399);
and U9914 (N_9914,N_8328,N_8175);
and U9915 (N_9915,N_8348,N_8189);
or U9916 (N_9916,N_8792,N_8068);
nand U9917 (N_9917,N_8067,N_8859);
xor U9918 (N_9918,N_8755,N_8396);
nand U9919 (N_9919,N_8925,N_8918);
nor U9920 (N_9920,N_8893,N_8857);
xnor U9921 (N_9921,N_8999,N_8992);
nor U9922 (N_9922,N_8569,N_8663);
and U9923 (N_9923,N_8107,N_8885);
or U9924 (N_9924,N_8519,N_8113);
and U9925 (N_9925,N_8331,N_8002);
and U9926 (N_9926,N_8568,N_8961);
nand U9927 (N_9927,N_8533,N_8244);
or U9928 (N_9928,N_8314,N_8938);
and U9929 (N_9929,N_8362,N_8379);
nor U9930 (N_9930,N_8195,N_8688);
nor U9931 (N_9931,N_8074,N_8962);
nor U9932 (N_9932,N_8759,N_8062);
or U9933 (N_9933,N_8025,N_8220);
xor U9934 (N_9934,N_8851,N_8923);
nand U9935 (N_9935,N_8730,N_8012);
and U9936 (N_9936,N_8811,N_8578);
and U9937 (N_9937,N_8594,N_8382);
nor U9938 (N_9938,N_8629,N_8912);
and U9939 (N_9939,N_8509,N_8512);
nor U9940 (N_9940,N_8379,N_8587);
xnor U9941 (N_9941,N_8827,N_8822);
or U9942 (N_9942,N_8707,N_8659);
or U9943 (N_9943,N_8521,N_8857);
and U9944 (N_9944,N_8309,N_8938);
or U9945 (N_9945,N_8620,N_8384);
xnor U9946 (N_9946,N_8473,N_8329);
nor U9947 (N_9947,N_8941,N_8363);
xor U9948 (N_9948,N_8209,N_8848);
or U9949 (N_9949,N_8488,N_8067);
nor U9950 (N_9950,N_8767,N_8272);
nor U9951 (N_9951,N_8781,N_8440);
and U9952 (N_9952,N_8598,N_8149);
nor U9953 (N_9953,N_8536,N_8191);
and U9954 (N_9954,N_8287,N_8965);
nand U9955 (N_9955,N_8373,N_8116);
nand U9956 (N_9956,N_8370,N_8782);
and U9957 (N_9957,N_8484,N_8646);
and U9958 (N_9958,N_8830,N_8052);
xor U9959 (N_9959,N_8612,N_8810);
xor U9960 (N_9960,N_8971,N_8890);
nor U9961 (N_9961,N_8416,N_8175);
nand U9962 (N_9962,N_8773,N_8555);
xor U9963 (N_9963,N_8981,N_8354);
and U9964 (N_9964,N_8558,N_8381);
nor U9965 (N_9965,N_8488,N_8462);
nor U9966 (N_9966,N_8528,N_8995);
nand U9967 (N_9967,N_8611,N_8726);
nor U9968 (N_9968,N_8423,N_8692);
xnor U9969 (N_9969,N_8705,N_8440);
or U9970 (N_9970,N_8278,N_8366);
xnor U9971 (N_9971,N_8277,N_8136);
nor U9972 (N_9972,N_8936,N_8241);
or U9973 (N_9973,N_8530,N_8086);
and U9974 (N_9974,N_8843,N_8533);
nand U9975 (N_9975,N_8372,N_8069);
xnor U9976 (N_9976,N_8610,N_8088);
xor U9977 (N_9977,N_8086,N_8163);
xor U9978 (N_9978,N_8975,N_8548);
or U9979 (N_9979,N_8671,N_8320);
and U9980 (N_9980,N_8637,N_8486);
nor U9981 (N_9981,N_8115,N_8566);
nand U9982 (N_9982,N_8507,N_8969);
and U9983 (N_9983,N_8583,N_8246);
or U9984 (N_9984,N_8702,N_8879);
or U9985 (N_9985,N_8533,N_8251);
or U9986 (N_9986,N_8538,N_8580);
and U9987 (N_9987,N_8632,N_8803);
xor U9988 (N_9988,N_8523,N_8596);
and U9989 (N_9989,N_8169,N_8930);
xor U9990 (N_9990,N_8862,N_8774);
and U9991 (N_9991,N_8781,N_8164);
nor U9992 (N_9992,N_8835,N_8585);
xnor U9993 (N_9993,N_8121,N_8737);
nor U9994 (N_9994,N_8049,N_8469);
nand U9995 (N_9995,N_8381,N_8391);
or U9996 (N_9996,N_8886,N_8519);
nor U9997 (N_9997,N_8484,N_8248);
nand U9998 (N_9998,N_8240,N_8204);
nand U9999 (N_9999,N_8031,N_8823);
nor U10000 (N_10000,N_9861,N_9790);
and U10001 (N_10001,N_9287,N_9275);
nor U10002 (N_10002,N_9923,N_9847);
nor U10003 (N_10003,N_9495,N_9663);
nor U10004 (N_10004,N_9160,N_9122);
nand U10005 (N_10005,N_9000,N_9124);
xnor U10006 (N_10006,N_9992,N_9588);
or U10007 (N_10007,N_9474,N_9027);
xnor U10008 (N_10008,N_9263,N_9099);
nor U10009 (N_10009,N_9039,N_9153);
and U10010 (N_10010,N_9497,N_9491);
nand U10011 (N_10011,N_9824,N_9567);
and U10012 (N_10012,N_9305,N_9919);
xor U10013 (N_10013,N_9737,N_9545);
and U10014 (N_10014,N_9937,N_9139);
nand U10015 (N_10015,N_9557,N_9765);
and U10016 (N_10016,N_9306,N_9309);
nand U10017 (N_10017,N_9354,N_9433);
and U10018 (N_10018,N_9386,N_9652);
nor U10019 (N_10019,N_9860,N_9047);
or U10020 (N_10020,N_9524,N_9964);
nor U10021 (N_10021,N_9719,N_9402);
nand U10022 (N_10022,N_9628,N_9695);
or U10023 (N_10023,N_9585,N_9600);
or U10024 (N_10024,N_9704,N_9133);
nor U10025 (N_10025,N_9336,N_9261);
and U10026 (N_10026,N_9269,N_9262);
nor U10027 (N_10027,N_9953,N_9101);
or U10028 (N_10028,N_9839,N_9978);
nand U10029 (N_10029,N_9996,N_9137);
xnor U10030 (N_10030,N_9375,N_9237);
and U10031 (N_10031,N_9449,N_9519);
and U10032 (N_10032,N_9598,N_9615);
nor U10033 (N_10033,N_9014,N_9098);
or U10034 (N_10034,N_9035,N_9420);
xor U10035 (N_10035,N_9258,N_9845);
nand U10036 (N_10036,N_9869,N_9983);
nor U10037 (N_10037,N_9674,N_9412);
or U10038 (N_10038,N_9537,N_9738);
nand U10039 (N_10039,N_9076,N_9288);
and U10040 (N_10040,N_9390,N_9095);
xor U10041 (N_10041,N_9142,N_9686);
xnor U10042 (N_10042,N_9225,N_9195);
xnor U10043 (N_10043,N_9882,N_9163);
and U10044 (N_10044,N_9389,N_9709);
xor U10045 (N_10045,N_9618,N_9363);
or U10046 (N_10046,N_9979,N_9054);
and U10047 (N_10047,N_9427,N_9013);
xor U10048 (N_10048,N_9611,N_9104);
or U10049 (N_10049,N_9779,N_9702);
or U10050 (N_10050,N_9636,N_9460);
or U10051 (N_10051,N_9612,N_9894);
nor U10052 (N_10052,N_9121,N_9453);
and U10053 (N_10053,N_9362,N_9659);
nor U10054 (N_10054,N_9494,N_9568);
nand U10055 (N_10055,N_9602,N_9909);
nand U10056 (N_10056,N_9310,N_9543);
or U10057 (N_10057,N_9048,N_9271);
nor U10058 (N_10058,N_9194,N_9821);
or U10059 (N_10059,N_9823,N_9374);
xnor U10060 (N_10060,N_9204,N_9871);
or U10061 (N_10061,N_9769,N_9883);
or U10062 (N_10062,N_9081,N_9028);
nor U10063 (N_10063,N_9538,N_9623);
xor U10064 (N_10064,N_9743,N_9371);
nand U10065 (N_10065,N_9378,N_9658);
xnor U10066 (N_10066,N_9346,N_9555);
nand U10067 (N_10067,N_9967,N_9084);
or U10068 (N_10068,N_9185,N_9068);
and U10069 (N_10069,N_9107,N_9925);
nor U10070 (N_10070,N_9922,N_9757);
xor U10071 (N_10071,N_9850,N_9958);
nor U10072 (N_10072,N_9862,N_9172);
nor U10073 (N_10073,N_9653,N_9228);
nand U10074 (N_10074,N_9630,N_9140);
and U10075 (N_10075,N_9733,N_9739);
and U10076 (N_10076,N_9638,N_9289);
nand U10077 (N_10077,N_9096,N_9024);
or U10078 (N_10078,N_9029,N_9146);
and U10079 (N_10079,N_9514,N_9441);
nor U10080 (N_10080,N_9498,N_9637);
nand U10081 (N_10081,N_9331,N_9404);
nor U10082 (N_10082,N_9298,N_9102);
nand U10083 (N_10083,N_9956,N_9209);
nand U10084 (N_10084,N_9428,N_9866);
xnor U10085 (N_10085,N_9665,N_9946);
and U10086 (N_10086,N_9754,N_9459);
and U10087 (N_10087,N_9949,N_9191);
nor U10088 (N_10088,N_9462,N_9587);
or U10089 (N_10089,N_9252,N_9670);
nand U10090 (N_10090,N_9347,N_9961);
or U10091 (N_10091,N_9372,N_9406);
and U10092 (N_10092,N_9534,N_9301);
or U10093 (N_10093,N_9985,N_9432);
nand U10094 (N_10094,N_9912,N_9721);
and U10095 (N_10095,N_9994,N_9166);
xnor U10096 (N_10096,N_9234,N_9276);
xnor U10097 (N_10097,N_9804,N_9466);
and U10098 (N_10098,N_9905,N_9025);
nand U10099 (N_10099,N_9669,N_9945);
nand U10100 (N_10100,N_9577,N_9808);
and U10101 (N_10101,N_9890,N_9312);
and U10102 (N_10102,N_9936,N_9366);
nand U10103 (N_10103,N_9679,N_9118);
nand U10104 (N_10104,N_9279,N_9159);
and U10105 (N_10105,N_9734,N_9328);
xor U10106 (N_10106,N_9868,N_9929);
nand U10107 (N_10107,N_9859,N_9988);
nor U10108 (N_10108,N_9852,N_9960);
or U10109 (N_10109,N_9499,N_9316);
nor U10110 (N_10110,N_9536,N_9162);
and U10111 (N_10111,N_9833,N_9640);
and U10112 (N_10112,N_9878,N_9771);
nor U10113 (N_10113,N_9840,N_9671);
nor U10114 (N_10114,N_9250,N_9317);
or U10115 (N_10115,N_9981,N_9214);
or U10116 (N_10116,N_9717,N_9751);
xnor U10117 (N_10117,N_9435,N_9512);
xor U10118 (N_10118,N_9535,N_9277);
nor U10119 (N_10119,N_9812,N_9976);
nand U10120 (N_10120,N_9626,N_9016);
and U10121 (N_10121,N_9339,N_9240);
or U10122 (N_10122,N_9093,N_9530);
nand U10123 (N_10123,N_9801,N_9542);
nand U10124 (N_10124,N_9415,N_9825);
nor U10125 (N_10125,N_9780,N_9110);
or U10126 (N_10126,N_9716,N_9675);
and U10127 (N_10127,N_9888,N_9711);
or U10128 (N_10128,N_9791,N_9583);
nor U10129 (N_10129,N_9643,N_9832);
nor U10130 (N_10130,N_9473,N_9006);
or U10131 (N_10131,N_9792,N_9188);
or U10132 (N_10132,N_9338,N_9179);
xnor U10133 (N_10133,N_9184,N_9731);
and U10134 (N_10134,N_9323,N_9421);
or U10135 (N_10135,N_9863,N_9220);
or U10136 (N_10136,N_9603,N_9759);
nand U10137 (N_10137,N_9877,N_9785);
and U10138 (N_10138,N_9827,N_9294);
nor U10139 (N_10139,N_9297,N_9423);
or U10140 (N_10140,N_9073,N_9710);
xnor U10141 (N_10141,N_9573,N_9311);
xor U10142 (N_10142,N_9224,N_9489);
and U10143 (N_10143,N_9436,N_9383);
xor U10144 (N_10144,N_9503,N_9798);
or U10145 (N_10145,N_9931,N_9395);
nor U10146 (N_10146,N_9198,N_9472);
nor U10147 (N_10147,N_9405,N_9400);
xnor U10148 (N_10148,N_9770,N_9954);
nor U10149 (N_10149,N_9112,N_9767);
and U10150 (N_10150,N_9930,N_9515);
or U10151 (N_10151,N_9712,N_9464);
and U10152 (N_10152,N_9174,N_9642);
and U10153 (N_10153,N_9203,N_9033);
and U10154 (N_10154,N_9126,N_9886);
nand U10155 (N_10155,N_9511,N_9008);
or U10156 (N_10156,N_9571,N_9049);
xnor U10157 (N_10157,N_9351,N_9062);
nand U10158 (N_10158,N_9274,N_9947);
xor U10159 (N_10159,N_9607,N_9553);
and U10160 (N_10160,N_9259,N_9501);
or U10161 (N_10161,N_9896,N_9962);
or U10162 (N_10162,N_9022,N_9678);
nor U10163 (N_10163,N_9797,N_9778);
and U10164 (N_10164,N_9111,N_9060);
nand U10165 (N_10165,N_9321,N_9278);
nor U10166 (N_10166,N_9307,N_9326);
xnor U10167 (N_10167,N_9736,N_9058);
nand U10168 (N_10168,N_9273,N_9546);
nor U10169 (N_10169,N_9693,N_9963);
nor U10170 (N_10170,N_9470,N_9606);
nor U10171 (N_10171,N_9270,N_9044);
nor U10172 (N_10172,N_9452,N_9249);
xor U10173 (N_10173,N_9186,N_9264);
nor U10174 (N_10174,N_9613,N_9345);
and U10175 (N_10175,N_9621,N_9566);
nor U10176 (N_10176,N_9318,N_9722);
xor U10177 (N_10177,N_9071,N_9023);
nor U10178 (N_10178,N_9496,N_9079);
or U10179 (N_10179,N_9714,N_9753);
nand U10180 (N_10180,N_9899,N_9820);
xor U10181 (N_10181,N_9192,N_9619);
and U10182 (N_10182,N_9744,N_9382);
nor U10183 (N_10183,N_9493,N_9291);
nand U10184 (N_10184,N_9350,N_9763);
or U10185 (N_10185,N_9826,N_9810);
or U10186 (N_10186,N_9902,N_9819);
or U10187 (N_10187,N_9007,N_9924);
or U10188 (N_10188,N_9380,N_9768);
nand U10189 (N_10189,N_9520,N_9189);
nor U10190 (N_10190,N_9698,N_9487);
or U10191 (N_10191,N_9418,N_9468);
or U10192 (N_10192,N_9564,N_9236);
or U10193 (N_10193,N_9835,N_9397);
and U10194 (N_10194,N_9181,N_9772);
xor U10195 (N_10195,N_9706,N_9943);
nand U10196 (N_10196,N_9088,N_9015);
nand U10197 (N_10197,N_9916,N_9213);
nor U10198 (N_10198,N_9756,N_9822);
or U10199 (N_10199,N_9300,N_9451);
nor U10200 (N_10200,N_9851,N_9340);
or U10201 (N_10201,N_9687,N_9781);
nor U10202 (N_10202,N_9986,N_9541);
nand U10203 (N_10203,N_9548,N_9115);
nor U10204 (N_10204,N_9841,N_9726);
nor U10205 (N_10205,N_9083,N_9647);
xor U10206 (N_10206,N_9149,N_9900);
or U10207 (N_10207,N_9425,N_9447);
nand U10208 (N_10208,N_9001,N_9408);
or U10209 (N_10209,N_9517,N_9881);
nor U10210 (N_10210,N_9199,N_9117);
nor U10211 (N_10211,N_9855,N_9265);
or U10212 (N_10212,N_9074,N_9042);
xnor U10213 (N_10213,N_9917,N_9525);
or U10214 (N_10214,N_9103,N_9685);
xnor U10215 (N_10215,N_9399,N_9657);
xnor U10216 (N_10216,N_9631,N_9718);
xor U10217 (N_10217,N_9951,N_9786);
nand U10218 (N_10218,N_9304,N_9446);
or U10219 (N_10219,N_9668,N_9795);
and U10220 (N_10220,N_9907,N_9941);
and U10221 (N_10221,N_9673,N_9552);
nor U10222 (N_10222,N_9993,N_9794);
or U10223 (N_10223,N_9867,N_9041);
nand U10224 (N_10224,N_9982,N_9085);
and U10225 (N_10225,N_9471,N_9217);
nand U10226 (N_10226,N_9620,N_9782);
nand U10227 (N_10227,N_9341,N_9703);
or U10228 (N_10228,N_9559,N_9507);
nor U10229 (N_10229,N_9950,N_9639);
xnor U10230 (N_10230,N_9901,N_9222);
xor U10231 (N_10231,N_9616,N_9151);
nor U10232 (N_10232,N_9991,N_9513);
xor U10233 (N_10233,N_9476,N_9752);
nand U10234 (N_10234,N_9522,N_9144);
nand U10235 (N_10235,N_9036,N_9777);
nor U10236 (N_10236,N_9388,N_9556);
or U10237 (N_10237,N_9504,N_9248);
and U10238 (N_10238,N_9742,N_9729);
or U10239 (N_10239,N_9226,N_9125);
nand U10240 (N_10240,N_9429,N_9461);
nand U10241 (N_10241,N_9903,N_9002);
nand U10242 (N_10242,N_9809,N_9957);
xor U10243 (N_10243,N_9987,N_9865);
or U10244 (N_10244,N_9582,N_9648);
and U10245 (N_10245,N_9268,N_9677);
xor U10246 (N_10246,N_9183,N_9565);
and U10247 (N_10247,N_9135,N_9417);
nand U10248 (N_10248,N_9651,N_9244);
nor U10249 (N_10249,N_9562,N_9385);
nand U10250 (N_10250,N_9486,N_9972);
or U10251 (N_10251,N_9688,N_9359);
nor U10252 (N_10252,N_9034,N_9356);
xor U10253 (N_10253,N_9296,N_9070);
nor U10254 (N_10254,N_9131,N_9691);
and U10255 (N_10255,N_9773,N_9529);
nand U10256 (N_10256,N_9330,N_9599);
nand U10257 (N_10257,N_9509,N_9523);
xnor U10258 (N_10258,N_9010,N_9128);
nor U10259 (N_10259,N_9342,N_9325);
xor U10260 (N_10260,N_9510,N_9200);
or U10261 (N_10261,N_9069,N_9828);
or U10262 (N_10262,N_9885,N_9431);
xor U10263 (N_10263,N_9457,N_9313);
xnor U10264 (N_10264,N_9114,N_9784);
nor U10265 (N_10265,N_9176,N_9935);
nand U10266 (N_10266,N_9239,N_9683);
or U10267 (N_10267,N_9030,N_9168);
or U10268 (N_10268,N_9539,N_9290);
xor U10269 (N_10269,N_9660,N_9020);
or U10270 (N_10270,N_9066,N_9077);
or U10271 (N_10271,N_9796,N_9662);
or U10272 (N_10272,N_9177,N_9123);
nand U10273 (N_10273,N_9910,N_9829);
or U10274 (N_10274,N_9971,N_9051);
or U10275 (N_10275,N_9701,N_9257);
or U10276 (N_10276,N_9959,N_9202);
or U10277 (N_10277,N_9045,N_9046);
and U10278 (N_10278,N_9880,N_9879);
xnor U10279 (N_10279,N_9645,N_9141);
nor U10280 (N_10280,N_9260,N_9700);
nor U10281 (N_10281,N_9082,N_9764);
xnor U10282 (N_10282,N_9834,N_9094);
nor U10283 (N_10283,N_9377,N_9891);
and U10284 (N_10284,N_9403,N_9550);
xnor U10285 (N_10285,N_9940,N_9358);
nor U10286 (N_10286,N_9218,N_9370);
and U10287 (N_10287,N_9134,N_9246);
and U10288 (N_10288,N_9018,N_9438);
or U10289 (N_10289,N_9267,N_9800);
nand U10290 (N_10290,N_9465,N_9109);
nand U10291 (N_10291,N_9629,N_9622);
nand U10292 (N_10292,N_9641,N_9748);
nor U10293 (N_10293,N_9672,N_9857);
or U10294 (N_10294,N_9696,N_9995);
nand U10295 (N_10295,N_9817,N_9019);
nor U10296 (N_10296,N_9059,N_9989);
nand U10297 (N_10297,N_9968,N_9811);
or U10298 (N_10298,N_9970,N_9337);
and U10299 (N_10299,N_9130,N_9975);
nor U10300 (N_10300,N_9575,N_9167);
or U10301 (N_10301,N_9928,N_9038);
or U10302 (N_10302,N_9627,N_9661);
xnor U10303 (N_10303,N_9597,N_9254);
nor U10304 (N_10304,N_9776,N_9352);
or U10305 (N_10305,N_9915,N_9610);
nand U10306 (N_10306,N_9143,N_9939);
and U10307 (N_10307,N_9387,N_9732);
nand U10308 (N_10308,N_9938,N_9170);
and U10309 (N_10309,N_9327,N_9369);
nor U10310 (N_10310,N_9761,N_9596);
and U10311 (N_10311,N_9895,N_9361);
nor U10312 (N_10312,N_9031,N_9157);
or U10313 (N_10313,N_9419,N_9984);
xnor U10314 (N_10314,N_9223,N_9303);
nor U10315 (N_10315,N_9502,N_9911);
nand U10316 (N_10316,N_9478,N_9649);
xnor U10317 (N_10317,N_9450,N_9087);
and U10318 (N_10318,N_9171,N_9707);
and U10319 (N_10319,N_9475,N_9766);
and U10320 (N_10320,N_9793,N_9805);
or U10321 (N_10321,N_9293,N_9414);
nand U10322 (N_10322,N_9547,N_9724);
and U10323 (N_10323,N_9136,N_9091);
nor U10324 (N_10324,N_9664,N_9040);
and U10325 (N_10325,N_9154,N_9818);
xnor U10326 (N_10326,N_9032,N_9723);
or U10327 (N_10327,N_9479,N_9830);
nand U10328 (N_10328,N_9333,N_9578);
xor U10329 (N_10329,N_9241,N_9009);
and U10330 (N_10330,N_9646,N_9760);
and U10331 (N_10331,N_9526,N_9201);
nand U10332 (N_10332,N_9758,N_9974);
and U10333 (N_10333,N_9212,N_9591);
xnor U10334 (N_10334,N_9365,N_9516);
nand U10335 (N_10335,N_9158,N_9017);
xor U10336 (N_10336,N_9918,N_9196);
xnor U10337 (N_10337,N_9579,N_9676);
and U10338 (N_10338,N_9283,N_9601);
nor U10339 (N_10339,N_9814,N_9178);
and U10340 (N_10340,N_9500,N_9614);
nand U10341 (N_10341,N_9454,N_9593);
xor U10342 (N_10342,N_9853,N_9393);
nor U10343 (N_10343,N_9344,N_9266);
and U10344 (N_10344,N_9799,N_9965);
nor U10345 (N_10345,N_9926,N_9242);
and U10346 (N_10346,N_9803,N_9576);
nor U10347 (N_10347,N_9286,N_9355);
or U10348 (N_10348,N_9531,N_9373);
and U10349 (N_10349,N_9381,N_9842);
nand U10350 (N_10350,N_9063,N_9667);
nand U10351 (N_10351,N_9934,N_9870);
xor U10352 (N_10352,N_9745,N_9207);
and U10353 (N_10353,N_9343,N_9119);
nor U10354 (N_10354,N_9401,N_9132);
or U10355 (N_10355,N_9376,N_9332);
xnor U10356 (N_10356,N_9836,N_9854);
nand U10357 (N_10357,N_9229,N_9540);
xnor U10358 (N_10358,N_9043,N_9708);
and U10359 (N_10359,N_9353,N_9394);
nand U10360 (N_10360,N_9874,N_9889);
nor U10361 (N_10361,N_9413,N_9872);
nor U10362 (N_10362,N_9011,N_9424);
and U10363 (N_10363,N_9904,N_9057);
or U10364 (N_10364,N_9692,N_9302);
and U10365 (N_10365,N_9713,N_9080);
nand U10366 (N_10366,N_9092,N_9998);
xor U10367 (N_10367,N_9072,N_9608);
nand U10368 (N_10368,N_9990,N_9730);
or U10369 (N_10369,N_9532,N_9884);
nor U10370 (N_10370,N_9584,N_9442);
xnor U10371 (N_10371,N_9064,N_9815);
nand U10372 (N_10372,N_9205,N_9272);
xnor U10373 (N_10373,N_9741,N_9521);
and U10374 (N_10374,N_9161,N_9314);
and U10375 (N_10375,N_9148,N_9893);
and U10376 (N_10376,N_9284,N_9997);
and U10377 (N_10377,N_9831,N_9368);
nand U10378 (N_10378,N_9238,N_9021);
or U10379 (N_10379,N_9586,N_9292);
nand U10380 (N_10380,N_9156,N_9458);
and U10381 (N_10381,N_9746,N_9106);
nand U10382 (N_10382,N_9783,N_9255);
nor U10383 (N_10383,N_9078,N_9426);
and U10384 (N_10384,N_9913,N_9506);
or U10385 (N_10385,N_9280,N_9595);
nand U10386 (N_10386,N_9589,N_9747);
xnor U10387 (N_10387,N_9681,N_9933);
or U10388 (N_10388,N_9319,N_9129);
or U10389 (N_10389,N_9392,N_9299);
or U10390 (N_10390,N_9789,N_9409);
xnor U10391 (N_10391,N_9053,N_9802);
and U10392 (N_10392,N_9334,N_9230);
xnor U10393 (N_10393,N_9108,N_9480);
and U10394 (N_10394,N_9838,N_9398);
or U10395 (N_10395,N_9469,N_9697);
or U10396 (N_10396,N_9210,N_9012);
xnor U10397 (N_10397,N_9594,N_9282);
and U10398 (N_10398,N_9492,N_9843);
and U10399 (N_10399,N_9897,N_9164);
or U10400 (N_10400,N_9689,N_9285);
nor U10401 (N_10401,N_9206,N_9624);
and U10402 (N_10402,N_9580,N_9932);
nand U10403 (N_10403,N_9320,N_9533);
and U10404 (N_10404,N_9256,N_9705);
and U10405 (N_10405,N_9243,N_9921);
nand U10406 (N_10406,N_9774,N_9856);
and U10407 (N_10407,N_9357,N_9037);
nor U10408 (N_10408,N_9065,N_9050);
or U10409 (N_10409,N_9977,N_9527);
nor U10410 (N_10410,N_9221,N_9251);
nand U10411 (N_10411,N_9656,N_9120);
or U10412 (N_10412,N_9873,N_9097);
nand U10413 (N_10413,N_9898,N_9490);
nand U10414 (N_10414,N_9145,N_9335);
and U10415 (N_10415,N_9384,N_9407);
xor U10416 (N_10416,N_9560,N_9090);
or U10417 (N_10417,N_9633,N_9914);
nor U10418 (N_10418,N_9849,N_9755);
nor U10419 (N_10419,N_9360,N_9574);
nand U10420 (N_10420,N_9349,N_9684);
xnor U10421 (N_10421,N_9563,N_9806);
nand U10422 (N_10422,N_9906,N_9155);
or U10423 (N_10423,N_9253,N_9422);
nand U10424 (N_10424,N_9245,N_9682);
nand U10425 (N_10425,N_9089,N_9813);
or U10426 (N_10426,N_9483,N_9680);
nand U10427 (N_10427,N_9175,N_9655);
and U10428 (N_10428,N_9650,N_9484);
xor U10429 (N_10429,N_9455,N_9942);
xnor U10430 (N_10430,N_9232,N_9544);
nand U10431 (N_10431,N_9569,N_9440);
and U10432 (N_10432,N_9572,N_9026);
nand U10433 (N_10433,N_9367,N_9443);
nand U10434 (N_10434,N_9056,N_9208);
and U10435 (N_10435,N_9235,N_9105);
xnor U10436 (N_10436,N_9694,N_9138);
xnor U10437 (N_10437,N_9750,N_9590);
or U10438 (N_10438,N_9625,N_9528);
xor U10439 (N_10439,N_9481,N_9182);
nor U10440 (N_10440,N_9690,N_9837);
nor U10441 (N_10441,N_9324,N_9379);
xnor U10442 (N_10442,N_9948,N_9762);
or U10443 (N_10443,N_9444,N_9980);
xnor U10444 (N_10444,N_9570,N_9448);
nand U10445 (N_10445,N_9875,N_9396);
xnor U10446 (N_10446,N_9604,N_9720);
and U10447 (N_10447,N_9920,N_9434);
or U10448 (N_10448,N_9100,N_9086);
xnor U10449 (N_10449,N_9807,N_9439);
nand U10450 (N_10450,N_9052,N_9113);
nand U10451 (N_10451,N_9999,N_9190);
nor U10452 (N_10452,N_9848,N_9281);
or U10453 (N_10453,N_9219,N_9635);
xor U10454 (N_10454,N_9617,N_9554);
nor U10455 (N_10455,N_9348,N_9699);
or U10456 (N_10456,N_9952,N_9846);
and U10457 (N_10457,N_9445,N_9116);
and U10458 (N_10458,N_9955,N_9715);
or U10459 (N_10459,N_9322,N_9416);
xor U10460 (N_10460,N_9127,N_9727);
nor U10461 (N_10461,N_9644,N_9927);
xnor U10462 (N_10462,N_9463,N_9969);
and U10463 (N_10463,N_9308,N_9061);
nand U10464 (N_10464,N_9654,N_9315);
xor U10465 (N_10465,N_9561,N_9467);
nor U10466 (N_10466,N_9634,N_9632);
nand U10467 (N_10467,N_9966,N_9728);
or U10468 (N_10468,N_9482,N_9165);
and U10469 (N_10469,N_9787,N_9816);
nor U10470 (N_10470,N_9067,N_9003);
and U10471 (N_10471,N_9892,N_9551);
nor U10472 (N_10472,N_9505,N_9055);
nor U10473 (N_10473,N_9197,N_9558);
or U10474 (N_10474,N_9187,N_9147);
or U10475 (N_10475,N_9740,N_9609);
nand U10476 (N_10476,N_9887,N_9216);
and U10477 (N_10477,N_9666,N_9150);
and U10478 (N_10478,N_9169,N_9908);
nor U10479 (N_10479,N_9391,N_9477);
nand U10480 (N_10480,N_9876,N_9233);
and U10481 (N_10481,N_9152,N_9410);
nor U10482 (N_10482,N_9973,N_9247);
and U10483 (N_10483,N_9004,N_9488);
xor U10484 (N_10484,N_9518,N_9605);
xor U10485 (N_10485,N_9844,N_9549);
nor U10486 (N_10486,N_9592,N_9211);
nor U10487 (N_10487,N_9788,N_9193);
nor U10488 (N_10488,N_9364,N_9858);
nand U10489 (N_10489,N_9430,N_9456);
or U10490 (N_10490,N_9005,N_9329);
nand U10491 (N_10491,N_9180,N_9173);
or U10492 (N_10492,N_9437,N_9295);
or U10493 (N_10493,N_9075,N_9944);
xnor U10494 (N_10494,N_9864,N_9231);
and U10495 (N_10495,N_9581,N_9485);
xnor U10496 (N_10496,N_9725,N_9227);
xnor U10497 (N_10497,N_9508,N_9735);
nor U10498 (N_10498,N_9775,N_9215);
and U10499 (N_10499,N_9749,N_9411);
nor U10500 (N_10500,N_9344,N_9194);
xor U10501 (N_10501,N_9691,N_9359);
nor U10502 (N_10502,N_9811,N_9652);
and U10503 (N_10503,N_9919,N_9713);
or U10504 (N_10504,N_9064,N_9237);
and U10505 (N_10505,N_9696,N_9312);
nor U10506 (N_10506,N_9461,N_9075);
xor U10507 (N_10507,N_9992,N_9175);
and U10508 (N_10508,N_9788,N_9508);
and U10509 (N_10509,N_9257,N_9411);
xor U10510 (N_10510,N_9476,N_9758);
and U10511 (N_10511,N_9805,N_9728);
xor U10512 (N_10512,N_9401,N_9970);
xor U10513 (N_10513,N_9611,N_9399);
xor U10514 (N_10514,N_9525,N_9598);
xnor U10515 (N_10515,N_9899,N_9872);
xor U10516 (N_10516,N_9860,N_9171);
or U10517 (N_10517,N_9791,N_9189);
xor U10518 (N_10518,N_9394,N_9465);
nor U10519 (N_10519,N_9084,N_9600);
and U10520 (N_10520,N_9306,N_9991);
and U10521 (N_10521,N_9716,N_9925);
nand U10522 (N_10522,N_9403,N_9107);
and U10523 (N_10523,N_9947,N_9873);
or U10524 (N_10524,N_9877,N_9249);
xor U10525 (N_10525,N_9752,N_9347);
nor U10526 (N_10526,N_9426,N_9457);
nor U10527 (N_10527,N_9596,N_9472);
or U10528 (N_10528,N_9327,N_9921);
xnor U10529 (N_10529,N_9370,N_9153);
and U10530 (N_10530,N_9044,N_9473);
nor U10531 (N_10531,N_9419,N_9231);
nor U10532 (N_10532,N_9131,N_9950);
xor U10533 (N_10533,N_9205,N_9640);
xor U10534 (N_10534,N_9080,N_9698);
nand U10535 (N_10535,N_9394,N_9219);
or U10536 (N_10536,N_9908,N_9624);
and U10537 (N_10537,N_9008,N_9130);
nand U10538 (N_10538,N_9583,N_9495);
xor U10539 (N_10539,N_9859,N_9704);
and U10540 (N_10540,N_9433,N_9025);
xnor U10541 (N_10541,N_9812,N_9409);
or U10542 (N_10542,N_9857,N_9878);
and U10543 (N_10543,N_9765,N_9790);
nor U10544 (N_10544,N_9634,N_9001);
xor U10545 (N_10545,N_9520,N_9444);
nand U10546 (N_10546,N_9265,N_9374);
nor U10547 (N_10547,N_9055,N_9375);
nor U10548 (N_10548,N_9807,N_9253);
nand U10549 (N_10549,N_9518,N_9330);
xor U10550 (N_10550,N_9328,N_9256);
nor U10551 (N_10551,N_9081,N_9335);
nand U10552 (N_10552,N_9803,N_9286);
or U10553 (N_10553,N_9175,N_9695);
xnor U10554 (N_10554,N_9893,N_9315);
and U10555 (N_10555,N_9908,N_9590);
nor U10556 (N_10556,N_9238,N_9357);
xor U10557 (N_10557,N_9368,N_9400);
xnor U10558 (N_10558,N_9207,N_9181);
and U10559 (N_10559,N_9547,N_9400);
xnor U10560 (N_10560,N_9040,N_9908);
or U10561 (N_10561,N_9200,N_9942);
nand U10562 (N_10562,N_9497,N_9346);
xor U10563 (N_10563,N_9708,N_9996);
and U10564 (N_10564,N_9778,N_9175);
xor U10565 (N_10565,N_9543,N_9112);
and U10566 (N_10566,N_9714,N_9833);
nand U10567 (N_10567,N_9649,N_9531);
nand U10568 (N_10568,N_9343,N_9496);
xor U10569 (N_10569,N_9778,N_9043);
or U10570 (N_10570,N_9452,N_9172);
xnor U10571 (N_10571,N_9150,N_9476);
or U10572 (N_10572,N_9002,N_9895);
nand U10573 (N_10573,N_9184,N_9779);
nor U10574 (N_10574,N_9257,N_9663);
and U10575 (N_10575,N_9640,N_9720);
or U10576 (N_10576,N_9536,N_9100);
or U10577 (N_10577,N_9244,N_9457);
xnor U10578 (N_10578,N_9942,N_9215);
and U10579 (N_10579,N_9774,N_9458);
xnor U10580 (N_10580,N_9492,N_9917);
nand U10581 (N_10581,N_9357,N_9905);
nand U10582 (N_10582,N_9786,N_9192);
and U10583 (N_10583,N_9911,N_9697);
or U10584 (N_10584,N_9048,N_9868);
nand U10585 (N_10585,N_9779,N_9128);
nand U10586 (N_10586,N_9449,N_9549);
and U10587 (N_10587,N_9323,N_9973);
xnor U10588 (N_10588,N_9692,N_9189);
nor U10589 (N_10589,N_9554,N_9129);
nand U10590 (N_10590,N_9342,N_9062);
nor U10591 (N_10591,N_9790,N_9593);
or U10592 (N_10592,N_9311,N_9556);
and U10593 (N_10593,N_9801,N_9612);
nor U10594 (N_10594,N_9380,N_9239);
and U10595 (N_10595,N_9499,N_9577);
or U10596 (N_10596,N_9045,N_9910);
and U10597 (N_10597,N_9225,N_9177);
nand U10598 (N_10598,N_9827,N_9442);
nand U10599 (N_10599,N_9530,N_9627);
nand U10600 (N_10600,N_9129,N_9251);
or U10601 (N_10601,N_9249,N_9815);
or U10602 (N_10602,N_9807,N_9906);
xor U10603 (N_10603,N_9343,N_9702);
nor U10604 (N_10604,N_9901,N_9898);
and U10605 (N_10605,N_9842,N_9034);
and U10606 (N_10606,N_9295,N_9214);
and U10607 (N_10607,N_9112,N_9758);
or U10608 (N_10608,N_9899,N_9161);
xnor U10609 (N_10609,N_9630,N_9022);
and U10610 (N_10610,N_9016,N_9655);
xnor U10611 (N_10611,N_9377,N_9129);
xnor U10612 (N_10612,N_9952,N_9378);
nor U10613 (N_10613,N_9536,N_9386);
nor U10614 (N_10614,N_9263,N_9337);
and U10615 (N_10615,N_9230,N_9995);
nand U10616 (N_10616,N_9517,N_9443);
xnor U10617 (N_10617,N_9885,N_9779);
xnor U10618 (N_10618,N_9339,N_9736);
and U10619 (N_10619,N_9366,N_9910);
or U10620 (N_10620,N_9590,N_9471);
xor U10621 (N_10621,N_9595,N_9271);
or U10622 (N_10622,N_9612,N_9653);
or U10623 (N_10623,N_9286,N_9296);
nand U10624 (N_10624,N_9190,N_9221);
nor U10625 (N_10625,N_9450,N_9602);
or U10626 (N_10626,N_9915,N_9447);
xnor U10627 (N_10627,N_9023,N_9333);
xnor U10628 (N_10628,N_9570,N_9805);
or U10629 (N_10629,N_9111,N_9471);
xor U10630 (N_10630,N_9166,N_9098);
nand U10631 (N_10631,N_9864,N_9811);
or U10632 (N_10632,N_9851,N_9529);
xnor U10633 (N_10633,N_9118,N_9501);
xnor U10634 (N_10634,N_9418,N_9423);
nand U10635 (N_10635,N_9581,N_9982);
nand U10636 (N_10636,N_9648,N_9572);
or U10637 (N_10637,N_9475,N_9997);
xnor U10638 (N_10638,N_9750,N_9929);
or U10639 (N_10639,N_9593,N_9846);
and U10640 (N_10640,N_9917,N_9395);
and U10641 (N_10641,N_9726,N_9757);
and U10642 (N_10642,N_9633,N_9261);
and U10643 (N_10643,N_9101,N_9886);
nand U10644 (N_10644,N_9861,N_9761);
nand U10645 (N_10645,N_9774,N_9119);
and U10646 (N_10646,N_9546,N_9169);
nand U10647 (N_10647,N_9434,N_9674);
and U10648 (N_10648,N_9654,N_9080);
xor U10649 (N_10649,N_9660,N_9206);
nand U10650 (N_10650,N_9800,N_9125);
nand U10651 (N_10651,N_9990,N_9149);
and U10652 (N_10652,N_9932,N_9618);
nand U10653 (N_10653,N_9759,N_9134);
and U10654 (N_10654,N_9518,N_9282);
and U10655 (N_10655,N_9806,N_9512);
and U10656 (N_10656,N_9447,N_9635);
or U10657 (N_10657,N_9445,N_9396);
and U10658 (N_10658,N_9586,N_9860);
or U10659 (N_10659,N_9835,N_9010);
nor U10660 (N_10660,N_9607,N_9443);
and U10661 (N_10661,N_9536,N_9848);
nand U10662 (N_10662,N_9840,N_9264);
nor U10663 (N_10663,N_9927,N_9494);
xor U10664 (N_10664,N_9559,N_9269);
nor U10665 (N_10665,N_9463,N_9807);
and U10666 (N_10666,N_9981,N_9038);
nor U10667 (N_10667,N_9257,N_9096);
xnor U10668 (N_10668,N_9339,N_9462);
and U10669 (N_10669,N_9877,N_9567);
and U10670 (N_10670,N_9404,N_9530);
xor U10671 (N_10671,N_9839,N_9530);
and U10672 (N_10672,N_9286,N_9343);
nand U10673 (N_10673,N_9260,N_9905);
and U10674 (N_10674,N_9070,N_9294);
or U10675 (N_10675,N_9957,N_9206);
nand U10676 (N_10676,N_9747,N_9877);
nand U10677 (N_10677,N_9673,N_9454);
and U10678 (N_10678,N_9760,N_9966);
xnor U10679 (N_10679,N_9261,N_9413);
nand U10680 (N_10680,N_9711,N_9237);
xnor U10681 (N_10681,N_9605,N_9438);
xor U10682 (N_10682,N_9932,N_9082);
nand U10683 (N_10683,N_9951,N_9089);
nand U10684 (N_10684,N_9929,N_9416);
or U10685 (N_10685,N_9804,N_9584);
or U10686 (N_10686,N_9246,N_9046);
nand U10687 (N_10687,N_9005,N_9357);
or U10688 (N_10688,N_9510,N_9625);
xor U10689 (N_10689,N_9797,N_9457);
nor U10690 (N_10690,N_9328,N_9749);
nor U10691 (N_10691,N_9777,N_9837);
xnor U10692 (N_10692,N_9640,N_9086);
and U10693 (N_10693,N_9298,N_9163);
nor U10694 (N_10694,N_9418,N_9907);
xnor U10695 (N_10695,N_9923,N_9943);
nand U10696 (N_10696,N_9812,N_9098);
and U10697 (N_10697,N_9126,N_9350);
nand U10698 (N_10698,N_9782,N_9734);
or U10699 (N_10699,N_9114,N_9166);
xor U10700 (N_10700,N_9932,N_9640);
nor U10701 (N_10701,N_9052,N_9849);
and U10702 (N_10702,N_9289,N_9821);
nor U10703 (N_10703,N_9728,N_9091);
nand U10704 (N_10704,N_9865,N_9711);
and U10705 (N_10705,N_9679,N_9884);
nor U10706 (N_10706,N_9285,N_9021);
xnor U10707 (N_10707,N_9500,N_9460);
nor U10708 (N_10708,N_9721,N_9437);
nor U10709 (N_10709,N_9269,N_9697);
and U10710 (N_10710,N_9298,N_9666);
nand U10711 (N_10711,N_9265,N_9002);
nor U10712 (N_10712,N_9769,N_9798);
nand U10713 (N_10713,N_9546,N_9494);
nor U10714 (N_10714,N_9908,N_9800);
xor U10715 (N_10715,N_9070,N_9334);
and U10716 (N_10716,N_9301,N_9055);
or U10717 (N_10717,N_9600,N_9489);
or U10718 (N_10718,N_9304,N_9010);
or U10719 (N_10719,N_9684,N_9551);
xor U10720 (N_10720,N_9744,N_9638);
xnor U10721 (N_10721,N_9334,N_9537);
nand U10722 (N_10722,N_9037,N_9871);
or U10723 (N_10723,N_9008,N_9972);
nand U10724 (N_10724,N_9334,N_9999);
or U10725 (N_10725,N_9909,N_9490);
nor U10726 (N_10726,N_9468,N_9714);
and U10727 (N_10727,N_9908,N_9551);
and U10728 (N_10728,N_9371,N_9194);
xor U10729 (N_10729,N_9056,N_9518);
or U10730 (N_10730,N_9270,N_9569);
or U10731 (N_10731,N_9385,N_9867);
nor U10732 (N_10732,N_9955,N_9545);
nand U10733 (N_10733,N_9450,N_9074);
xnor U10734 (N_10734,N_9177,N_9597);
nand U10735 (N_10735,N_9118,N_9131);
xor U10736 (N_10736,N_9611,N_9634);
nand U10737 (N_10737,N_9117,N_9204);
nand U10738 (N_10738,N_9764,N_9695);
or U10739 (N_10739,N_9988,N_9609);
and U10740 (N_10740,N_9833,N_9630);
or U10741 (N_10741,N_9049,N_9320);
xor U10742 (N_10742,N_9913,N_9370);
and U10743 (N_10743,N_9289,N_9499);
xor U10744 (N_10744,N_9445,N_9309);
nor U10745 (N_10745,N_9111,N_9188);
or U10746 (N_10746,N_9881,N_9987);
or U10747 (N_10747,N_9178,N_9926);
nand U10748 (N_10748,N_9893,N_9681);
xnor U10749 (N_10749,N_9284,N_9765);
and U10750 (N_10750,N_9280,N_9213);
nor U10751 (N_10751,N_9835,N_9221);
nand U10752 (N_10752,N_9549,N_9672);
nand U10753 (N_10753,N_9270,N_9633);
xnor U10754 (N_10754,N_9451,N_9262);
nor U10755 (N_10755,N_9310,N_9210);
xnor U10756 (N_10756,N_9340,N_9365);
xor U10757 (N_10757,N_9321,N_9989);
nand U10758 (N_10758,N_9644,N_9453);
nand U10759 (N_10759,N_9910,N_9838);
or U10760 (N_10760,N_9622,N_9501);
xor U10761 (N_10761,N_9676,N_9942);
xnor U10762 (N_10762,N_9472,N_9625);
and U10763 (N_10763,N_9182,N_9458);
nor U10764 (N_10764,N_9819,N_9989);
and U10765 (N_10765,N_9455,N_9741);
and U10766 (N_10766,N_9638,N_9207);
xnor U10767 (N_10767,N_9757,N_9860);
and U10768 (N_10768,N_9242,N_9869);
xor U10769 (N_10769,N_9193,N_9295);
or U10770 (N_10770,N_9366,N_9656);
xor U10771 (N_10771,N_9005,N_9064);
or U10772 (N_10772,N_9823,N_9629);
nand U10773 (N_10773,N_9511,N_9289);
or U10774 (N_10774,N_9092,N_9899);
or U10775 (N_10775,N_9285,N_9956);
or U10776 (N_10776,N_9175,N_9708);
xnor U10777 (N_10777,N_9176,N_9275);
nand U10778 (N_10778,N_9389,N_9468);
and U10779 (N_10779,N_9310,N_9368);
xnor U10780 (N_10780,N_9631,N_9895);
or U10781 (N_10781,N_9133,N_9684);
xnor U10782 (N_10782,N_9824,N_9548);
nor U10783 (N_10783,N_9813,N_9230);
or U10784 (N_10784,N_9716,N_9753);
or U10785 (N_10785,N_9232,N_9265);
nor U10786 (N_10786,N_9089,N_9426);
xor U10787 (N_10787,N_9371,N_9921);
and U10788 (N_10788,N_9323,N_9769);
xor U10789 (N_10789,N_9606,N_9643);
nor U10790 (N_10790,N_9774,N_9046);
and U10791 (N_10791,N_9438,N_9293);
xnor U10792 (N_10792,N_9456,N_9004);
or U10793 (N_10793,N_9313,N_9676);
or U10794 (N_10794,N_9492,N_9966);
and U10795 (N_10795,N_9757,N_9938);
and U10796 (N_10796,N_9663,N_9068);
nand U10797 (N_10797,N_9460,N_9689);
xor U10798 (N_10798,N_9056,N_9958);
or U10799 (N_10799,N_9644,N_9195);
and U10800 (N_10800,N_9940,N_9482);
nand U10801 (N_10801,N_9086,N_9868);
xnor U10802 (N_10802,N_9569,N_9095);
nor U10803 (N_10803,N_9615,N_9178);
xnor U10804 (N_10804,N_9202,N_9932);
xnor U10805 (N_10805,N_9482,N_9671);
xor U10806 (N_10806,N_9063,N_9673);
and U10807 (N_10807,N_9497,N_9799);
nand U10808 (N_10808,N_9002,N_9509);
nand U10809 (N_10809,N_9186,N_9256);
or U10810 (N_10810,N_9360,N_9657);
xnor U10811 (N_10811,N_9805,N_9862);
nand U10812 (N_10812,N_9186,N_9851);
and U10813 (N_10813,N_9322,N_9835);
xor U10814 (N_10814,N_9182,N_9657);
and U10815 (N_10815,N_9156,N_9085);
or U10816 (N_10816,N_9472,N_9457);
xor U10817 (N_10817,N_9632,N_9062);
xor U10818 (N_10818,N_9104,N_9624);
nand U10819 (N_10819,N_9457,N_9536);
and U10820 (N_10820,N_9645,N_9677);
xnor U10821 (N_10821,N_9148,N_9865);
and U10822 (N_10822,N_9589,N_9549);
or U10823 (N_10823,N_9640,N_9437);
or U10824 (N_10824,N_9379,N_9650);
or U10825 (N_10825,N_9842,N_9248);
nand U10826 (N_10826,N_9274,N_9621);
or U10827 (N_10827,N_9896,N_9140);
nand U10828 (N_10828,N_9713,N_9209);
xor U10829 (N_10829,N_9803,N_9482);
xor U10830 (N_10830,N_9675,N_9393);
and U10831 (N_10831,N_9422,N_9177);
or U10832 (N_10832,N_9727,N_9508);
nand U10833 (N_10833,N_9527,N_9694);
nand U10834 (N_10834,N_9524,N_9203);
and U10835 (N_10835,N_9304,N_9469);
or U10836 (N_10836,N_9566,N_9433);
and U10837 (N_10837,N_9872,N_9440);
and U10838 (N_10838,N_9256,N_9486);
nor U10839 (N_10839,N_9139,N_9520);
nor U10840 (N_10840,N_9210,N_9801);
nor U10841 (N_10841,N_9813,N_9796);
nor U10842 (N_10842,N_9885,N_9778);
nor U10843 (N_10843,N_9968,N_9150);
nand U10844 (N_10844,N_9568,N_9065);
and U10845 (N_10845,N_9981,N_9127);
nor U10846 (N_10846,N_9703,N_9932);
xnor U10847 (N_10847,N_9461,N_9899);
xnor U10848 (N_10848,N_9996,N_9238);
xnor U10849 (N_10849,N_9204,N_9994);
and U10850 (N_10850,N_9876,N_9900);
and U10851 (N_10851,N_9773,N_9595);
nand U10852 (N_10852,N_9395,N_9337);
or U10853 (N_10853,N_9459,N_9708);
or U10854 (N_10854,N_9691,N_9881);
nor U10855 (N_10855,N_9747,N_9592);
nor U10856 (N_10856,N_9984,N_9616);
xor U10857 (N_10857,N_9418,N_9084);
and U10858 (N_10858,N_9995,N_9397);
xor U10859 (N_10859,N_9758,N_9724);
xor U10860 (N_10860,N_9235,N_9672);
nor U10861 (N_10861,N_9881,N_9039);
nor U10862 (N_10862,N_9936,N_9094);
or U10863 (N_10863,N_9375,N_9685);
xnor U10864 (N_10864,N_9031,N_9304);
or U10865 (N_10865,N_9258,N_9904);
or U10866 (N_10866,N_9387,N_9474);
nand U10867 (N_10867,N_9108,N_9813);
nand U10868 (N_10868,N_9778,N_9290);
xor U10869 (N_10869,N_9626,N_9375);
nor U10870 (N_10870,N_9169,N_9487);
nor U10871 (N_10871,N_9353,N_9429);
nor U10872 (N_10872,N_9353,N_9784);
xor U10873 (N_10873,N_9592,N_9582);
nand U10874 (N_10874,N_9570,N_9824);
nand U10875 (N_10875,N_9457,N_9855);
nand U10876 (N_10876,N_9183,N_9648);
nor U10877 (N_10877,N_9643,N_9647);
xor U10878 (N_10878,N_9679,N_9545);
nor U10879 (N_10879,N_9225,N_9074);
nand U10880 (N_10880,N_9450,N_9169);
xor U10881 (N_10881,N_9098,N_9435);
nor U10882 (N_10882,N_9878,N_9371);
and U10883 (N_10883,N_9237,N_9042);
nor U10884 (N_10884,N_9278,N_9037);
and U10885 (N_10885,N_9318,N_9852);
xor U10886 (N_10886,N_9459,N_9181);
nand U10887 (N_10887,N_9526,N_9986);
and U10888 (N_10888,N_9268,N_9283);
and U10889 (N_10889,N_9414,N_9276);
nor U10890 (N_10890,N_9170,N_9733);
xnor U10891 (N_10891,N_9406,N_9308);
xnor U10892 (N_10892,N_9716,N_9004);
nand U10893 (N_10893,N_9919,N_9094);
nor U10894 (N_10894,N_9152,N_9411);
nor U10895 (N_10895,N_9101,N_9990);
nand U10896 (N_10896,N_9377,N_9965);
xnor U10897 (N_10897,N_9637,N_9321);
xor U10898 (N_10898,N_9149,N_9895);
and U10899 (N_10899,N_9245,N_9615);
xor U10900 (N_10900,N_9865,N_9961);
xnor U10901 (N_10901,N_9811,N_9758);
nor U10902 (N_10902,N_9316,N_9238);
and U10903 (N_10903,N_9910,N_9414);
and U10904 (N_10904,N_9597,N_9523);
nand U10905 (N_10905,N_9237,N_9528);
and U10906 (N_10906,N_9858,N_9216);
nand U10907 (N_10907,N_9706,N_9957);
nor U10908 (N_10908,N_9685,N_9540);
nor U10909 (N_10909,N_9049,N_9220);
or U10910 (N_10910,N_9155,N_9947);
or U10911 (N_10911,N_9530,N_9815);
nand U10912 (N_10912,N_9705,N_9722);
nor U10913 (N_10913,N_9185,N_9365);
nand U10914 (N_10914,N_9876,N_9933);
and U10915 (N_10915,N_9842,N_9872);
nor U10916 (N_10916,N_9683,N_9726);
nor U10917 (N_10917,N_9483,N_9777);
or U10918 (N_10918,N_9994,N_9745);
nor U10919 (N_10919,N_9467,N_9072);
and U10920 (N_10920,N_9168,N_9290);
xor U10921 (N_10921,N_9435,N_9876);
nand U10922 (N_10922,N_9384,N_9387);
xnor U10923 (N_10923,N_9292,N_9303);
and U10924 (N_10924,N_9569,N_9196);
nand U10925 (N_10925,N_9669,N_9204);
and U10926 (N_10926,N_9411,N_9393);
or U10927 (N_10927,N_9482,N_9079);
xor U10928 (N_10928,N_9237,N_9736);
or U10929 (N_10929,N_9852,N_9786);
and U10930 (N_10930,N_9275,N_9903);
nor U10931 (N_10931,N_9441,N_9279);
and U10932 (N_10932,N_9120,N_9118);
nor U10933 (N_10933,N_9273,N_9035);
nand U10934 (N_10934,N_9319,N_9810);
or U10935 (N_10935,N_9586,N_9932);
and U10936 (N_10936,N_9730,N_9064);
or U10937 (N_10937,N_9986,N_9358);
nor U10938 (N_10938,N_9238,N_9832);
or U10939 (N_10939,N_9797,N_9346);
nor U10940 (N_10940,N_9217,N_9375);
or U10941 (N_10941,N_9499,N_9308);
or U10942 (N_10942,N_9821,N_9663);
xnor U10943 (N_10943,N_9440,N_9184);
and U10944 (N_10944,N_9751,N_9564);
nand U10945 (N_10945,N_9739,N_9891);
and U10946 (N_10946,N_9973,N_9678);
xor U10947 (N_10947,N_9666,N_9295);
or U10948 (N_10948,N_9589,N_9612);
nand U10949 (N_10949,N_9415,N_9943);
xnor U10950 (N_10950,N_9052,N_9579);
nor U10951 (N_10951,N_9886,N_9263);
or U10952 (N_10952,N_9872,N_9508);
xnor U10953 (N_10953,N_9668,N_9451);
or U10954 (N_10954,N_9097,N_9720);
and U10955 (N_10955,N_9361,N_9246);
nand U10956 (N_10956,N_9605,N_9192);
xnor U10957 (N_10957,N_9135,N_9082);
and U10958 (N_10958,N_9706,N_9100);
nor U10959 (N_10959,N_9751,N_9839);
xnor U10960 (N_10960,N_9269,N_9839);
and U10961 (N_10961,N_9552,N_9492);
nor U10962 (N_10962,N_9367,N_9717);
xnor U10963 (N_10963,N_9026,N_9593);
xor U10964 (N_10964,N_9376,N_9224);
nand U10965 (N_10965,N_9980,N_9339);
nor U10966 (N_10966,N_9669,N_9513);
nor U10967 (N_10967,N_9003,N_9861);
or U10968 (N_10968,N_9938,N_9358);
or U10969 (N_10969,N_9364,N_9691);
or U10970 (N_10970,N_9069,N_9595);
xor U10971 (N_10971,N_9547,N_9221);
nand U10972 (N_10972,N_9999,N_9039);
or U10973 (N_10973,N_9101,N_9314);
nor U10974 (N_10974,N_9971,N_9687);
nor U10975 (N_10975,N_9686,N_9214);
or U10976 (N_10976,N_9963,N_9167);
xor U10977 (N_10977,N_9205,N_9057);
or U10978 (N_10978,N_9201,N_9355);
nor U10979 (N_10979,N_9156,N_9097);
nor U10980 (N_10980,N_9683,N_9464);
nand U10981 (N_10981,N_9437,N_9203);
nand U10982 (N_10982,N_9084,N_9920);
nor U10983 (N_10983,N_9848,N_9791);
nor U10984 (N_10984,N_9344,N_9160);
or U10985 (N_10985,N_9434,N_9034);
or U10986 (N_10986,N_9932,N_9543);
xor U10987 (N_10987,N_9586,N_9342);
xnor U10988 (N_10988,N_9375,N_9413);
xor U10989 (N_10989,N_9608,N_9162);
nor U10990 (N_10990,N_9676,N_9003);
nor U10991 (N_10991,N_9151,N_9006);
nor U10992 (N_10992,N_9665,N_9199);
or U10993 (N_10993,N_9414,N_9799);
or U10994 (N_10994,N_9863,N_9987);
nor U10995 (N_10995,N_9529,N_9455);
or U10996 (N_10996,N_9034,N_9240);
and U10997 (N_10997,N_9207,N_9037);
nand U10998 (N_10998,N_9577,N_9124);
or U10999 (N_10999,N_9907,N_9812);
and U11000 (N_11000,N_10416,N_10743);
xor U11001 (N_11001,N_10224,N_10360);
nand U11002 (N_11002,N_10796,N_10203);
or U11003 (N_11003,N_10495,N_10273);
and U11004 (N_11004,N_10401,N_10666);
nor U11005 (N_11005,N_10391,N_10990);
xnor U11006 (N_11006,N_10600,N_10361);
or U11007 (N_11007,N_10583,N_10109);
nor U11008 (N_11008,N_10425,N_10342);
nor U11009 (N_11009,N_10005,N_10143);
xor U11010 (N_11010,N_10722,N_10853);
xnor U11011 (N_11011,N_10013,N_10619);
or U11012 (N_11012,N_10841,N_10556);
xor U11013 (N_11013,N_10314,N_10376);
nor U11014 (N_11014,N_10855,N_10441);
or U11015 (N_11015,N_10698,N_10971);
xor U11016 (N_11016,N_10467,N_10091);
and U11017 (N_11017,N_10780,N_10587);
nand U11018 (N_11018,N_10106,N_10998);
and U11019 (N_11019,N_10799,N_10606);
and U11020 (N_11020,N_10813,N_10744);
nor U11021 (N_11021,N_10792,N_10029);
xor U11022 (N_11022,N_10649,N_10035);
xnor U11023 (N_11023,N_10565,N_10231);
nor U11024 (N_11024,N_10635,N_10573);
xnor U11025 (N_11025,N_10031,N_10329);
and U11026 (N_11026,N_10704,N_10118);
or U11027 (N_11027,N_10579,N_10580);
xor U11028 (N_11028,N_10161,N_10043);
or U11029 (N_11029,N_10122,N_10330);
and U11030 (N_11030,N_10087,N_10969);
and U11031 (N_11031,N_10067,N_10967);
xor U11032 (N_11032,N_10907,N_10303);
nand U11033 (N_11033,N_10693,N_10520);
xor U11034 (N_11034,N_10584,N_10269);
or U11035 (N_11035,N_10147,N_10589);
nand U11036 (N_11036,N_10006,N_10321);
and U11037 (N_11037,N_10253,N_10896);
nor U11038 (N_11038,N_10047,N_10760);
nand U11039 (N_11039,N_10810,N_10854);
xnor U11040 (N_11040,N_10605,N_10478);
nand U11041 (N_11041,N_10207,N_10137);
nand U11042 (N_11042,N_10383,N_10954);
or U11043 (N_11043,N_10826,N_10458);
xnor U11044 (N_11044,N_10912,N_10774);
and U11045 (N_11045,N_10513,N_10599);
nor U11046 (N_11046,N_10621,N_10811);
or U11047 (N_11047,N_10663,N_10468);
nand U11048 (N_11048,N_10536,N_10681);
nor U11049 (N_11049,N_10095,N_10222);
nand U11050 (N_11050,N_10604,N_10772);
or U11051 (N_11051,N_10687,N_10262);
or U11052 (N_11052,N_10252,N_10485);
nor U11053 (N_11053,N_10429,N_10756);
and U11054 (N_11054,N_10749,N_10643);
nand U11055 (N_11055,N_10205,N_10461);
nand U11056 (N_11056,N_10412,N_10977);
nor U11057 (N_11057,N_10845,N_10612);
nand U11058 (N_11058,N_10163,N_10966);
nor U11059 (N_11059,N_10084,N_10713);
nor U11060 (N_11060,N_10221,N_10011);
nand U11061 (N_11061,N_10922,N_10153);
or U11062 (N_11062,N_10973,N_10403);
and U11063 (N_11063,N_10070,N_10724);
and U11064 (N_11064,N_10155,N_10994);
and U11065 (N_11065,N_10530,N_10914);
nand U11066 (N_11066,N_10918,N_10846);
or U11067 (N_11067,N_10276,N_10246);
xor U11068 (N_11068,N_10823,N_10630);
or U11069 (N_11069,N_10627,N_10219);
or U11070 (N_11070,N_10673,N_10941);
xor U11071 (N_11071,N_10884,N_10754);
nor U11072 (N_11072,N_10484,N_10284);
nor U11073 (N_11073,N_10256,N_10025);
or U11074 (N_11074,N_10240,N_10509);
or U11075 (N_11075,N_10665,N_10036);
or U11076 (N_11076,N_10173,N_10209);
nand U11077 (N_11077,N_10558,N_10065);
nor U11078 (N_11078,N_10308,N_10568);
nor U11079 (N_11079,N_10229,N_10661);
or U11080 (N_11080,N_10124,N_10825);
and U11081 (N_11081,N_10697,N_10545);
xnor U11082 (N_11082,N_10156,N_10261);
or U11083 (N_11083,N_10519,N_10968);
xor U11084 (N_11084,N_10806,N_10088);
or U11085 (N_11085,N_10063,N_10232);
xnor U11086 (N_11086,N_10551,N_10432);
or U11087 (N_11087,N_10571,N_10911);
nor U11088 (N_11088,N_10422,N_10553);
or U11089 (N_11089,N_10542,N_10102);
and U11090 (N_11090,N_10936,N_10268);
nor U11091 (N_11091,N_10089,N_10337);
nand U11092 (N_11092,N_10861,N_10508);
nor U11093 (N_11093,N_10415,N_10367);
and U11094 (N_11094,N_10712,N_10370);
nand U11095 (N_11095,N_10313,N_10198);
nor U11096 (N_11096,N_10032,N_10591);
xor U11097 (N_11097,N_10493,N_10181);
and U11098 (N_11098,N_10510,N_10257);
or U11099 (N_11099,N_10372,N_10684);
nand U11100 (N_11100,N_10332,N_10081);
nor U11101 (N_11101,N_10214,N_10164);
or U11102 (N_11102,N_10647,N_10059);
or U11103 (N_11103,N_10608,N_10499);
or U11104 (N_11104,N_10932,N_10560);
nor U11105 (N_11105,N_10945,N_10236);
xnor U11106 (N_11106,N_10857,N_10856);
nor U11107 (N_11107,N_10529,N_10135);
nor U11108 (N_11108,N_10525,N_10909);
xor U11109 (N_11109,N_10593,N_10533);
xor U11110 (N_11110,N_10714,N_10325);
xnor U11111 (N_11111,N_10396,N_10201);
or U11112 (N_11112,N_10312,N_10935);
xor U11113 (N_11113,N_10588,N_10905);
xor U11114 (N_11114,N_10187,N_10271);
or U11115 (N_11115,N_10414,N_10944);
xor U11116 (N_11116,N_10386,N_10547);
nand U11117 (N_11117,N_10052,N_10993);
nor U11118 (N_11118,N_10477,N_10211);
nor U11119 (N_11119,N_10292,N_10819);
and U11120 (N_11120,N_10777,N_10265);
nor U11121 (N_11121,N_10715,N_10514);
nand U11122 (N_11122,N_10335,N_10624);
nor U11123 (N_11123,N_10549,N_10259);
xor U11124 (N_11124,N_10957,N_10557);
and U11125 (N_11125,N_10836,N_10516);
xnor U11126 (N_11126,N_10940,N_10294);
nand U11127 (N_11127,N_10931,N_10185);
nor U11128 (N_11128,N_10404,N_10097);
nor U11129 (N_11129,N_10788,N_10334);
or U11130 (N_11130,N_10601,N_10385);
nand U11131 (N_11131,N_10729,N_10505);
nor U11132 (N_11132,N_10778,N_10578);
and U11133 (N_11133,N_10389,N_10701);
or U11134 (N_11134,N_10498,N_10012);
nand U11135 (N_11135,N_10033,N_10920);
or U11136 (N_11136,N_10677,N_10476);
nand U11137 (N_11137,N_10730,N_10149);
nand U11138 (N_11138,N_10691,N_10466);
nand U11139 (N_11139,N_10829,N_10837);
nand U11140 (N_11140,N_10138,N_10597);
nor U11141 (N_11141,N_10742,N_10139);
and U11142 (N_11142,N_10355,N_10208);
nor U11143 (N_11143,N_10311,N_10787);
nor U11144 (N_11144,N_10368,N_10798);
nor U11145 (N_11145,N_10650,N_10460);
nor U11146 (N_11146,N_10528,N_10480);
nor U11147 (N_11147,N_10674,N_10289);
nor U11148 (N_11148,N_10518,N_10282);
xor U11149 (N_11149,N_10628,N_10042);
xor U11150 (N_11150,N_10781,N_10145);
nand U11151 (N_11151,N_10615,N_10379);
xnor U11152 (N_11152,N_10976,N_10763);
and U11153 (N_11153,N_10641,N_10077);
or U11154 (N_11154,N_10058,N_10226);
nand U11155 (N_11155,N_10668,N_10919);
xnor U11156 (N_11156,N_10475,N_10079);
nand U11157 (N_11157,N_10771,N_10353);
nor U11158 (N_11158,N_10879,N_10929);
and U11159 (N_11159,N_10115,N_10989);
nor U11160 (N_11160,N_10500,N_10487);
or U11161 (N_11161,N_10101,N_10793);
or U11162 (N_11162,N_10610,N_10297);
xnor U11163 (N_11163,N_10393,N_10183);
nand U11164 (N_11164,N_10288,N_10706);
and U11165 (N_11165,N_10891,N_10134);
nor U11166 (N_11166,N_10894,N_10463);
xnor U11167 (N_11167,N_10123,N_10490);
and U11168 (N_11168,N_10347,N_10263);
and U11169 (N_11169,N_10357,N_10725);
and U11170 (N_11170,N_10609,N_10535);
xnor U11171 (N_11171,N_10866,N_10318);
or U11172 (N_11172,N_10675,N_10200);
and U11173 (N_11173,N_10030,N_10167);
xor U11174 (N_11174,N_10769,N_10822);
or U11175 (N_11175,N_10595,N_10260);
and U11176 (N_11176,N_10291,N_10157);
and U11177 (N_11177,N_10670,N_10344);
nor U11178 (N_11178,N_10913,N_10373);
or U11179 (N_11179,N_10801,N_10045);
xnor U11180 (N_11180,N_10875,N_10794);
and U11181 (N_11181,N_10574,N_10930);
xnor U11182 (N_11182,N_10125,N_10340);
xor U11183 (N_11183,N_10924,N_10281);
xnor U11184 (N_11184,N_10119,N_10021);
and U11185 (N_11185,N_10820,N_10278);
nand U11186 (N_11186,N_10948,N_10305);
xnor U11187 (N_11187,N_10411,N_10504);
and U11188 (N_11188,N_10705,N_10864);
and U11189 (N_11189,N_10426,N_10522);
or U11190 (N_11190,N_10544,N_10274);
or U11191 (N_11191,N_10474,N_10680);
and U11192 (N_11192,N_10465,N_10096);
nor U11193 (N_11193,N_10803,N_10501);
nand U11194 (N_11194,N_10366,N_10204);
nor U11195 (N_11195,N_10152,N_10092);
nand U11196 (N_11196,N_10721,N_10451);
and U11197 (N_11197,N_10916,N_10479);
and U11198 (N_11198,N_10682,N_10953);
or U11199 (N_11199,N_10450,N_10765);
xnor U11200 (N_11200,N_10860,N_10423);
nor U11201 (N_11201,N_10105,N_10572);
and U11202 (N_11202,N_10736,N_10093);
nor U11203 (N_11203,N_10162,N_10108);
or U11204 (N_11204,N_10146,N_10975);
or U11205 (N_11205,N_10515,N_10443);
xnor U11206 (N_11206,N_10795,N_10452);
and U11207 (N_11207,N_10534,N_10060);
or U11208 (N_11208,N_10700,N_10507);
or U11209 (N_11209,N_10442,N_10992);
nor U11210 (N_11210,N_10345,N_10702);
xor U11211 (N_11211,N_10764,N_10655);
or U11212 (N_11212,N_10407,N_10054);
xnor U11213 (N_11213,N_10766,N_10188);
xor U11214 (N_11214,N_10020,N_10120);
or U11215 (N_11215,N_10223,N_10925);
xor U11216 (N_11216,N_10358,N_10494);
nand U11217 (N_11217,N_10885,N_10175);
and U11218 (N_11218,N_10759,N_10440);
xnor U11219 (N_11219,N_10306,N_10235);
nor U11220 (N_11220,N_10324,N_10503);
xnor U11221 (N_11221,N_10817,N_10662);
or U11222 (N_11222,N_10865,N_10350);
and U11223 (N_11223,N_10267,N_10327);
xor U11224 (N_11224,N_10692,N_10646);
nor U11225 (N_11225,N_10195,N_10398);
and U11226 (N_11226,N_10527,N_10094);
xor U11227 (N_11227,N_10618,N_10651);
xnor U11228 (N_11228,N_10934,N_10755);
xnor U11229 (N_11229,N_10238,N_10028);
nor U11230 (N_11230,N_10947,N_10242);
nand U11231 (N_11231,N_10116,N_10707);
or U11232 (N_11232,N_10511,N_10850);
or U11233 (N_11233,N_10076,N_10160);
xnor U11234 (N_11234,N_10319,N_10356);
and U11235 (N_11235,N_10815,N_10972);
nor U11236 (N_11236,N_10678,N_10351);
xnor U11237 (N_11237,N_10191,N_10171);
nand U11238 (N_11238,N_10409,N_10015);
nor U11239 (N_11239,N_10695,N_10981);
xor U11240 (N_11240,N_10293,N_10938);
xnor U11241 (N_11241,N_10213,N_10359);
nor U11242 (N_11242,N_10481,N_10720);
nand U11243 (N_11243,N_10166,N_10295);
nor U11244 (N_11244,N_10392,N_10645);
and U11245 (N_11245,N_10538,N_10038);
and U11246 (N_11246,N_10039,N_10014);
or U11247 (N_11247,N_10809,N_10377);
nand U11248 (N_11248,N_10464,N_10307);
xnor U11249 (N_11249,N_10085,N_10148);
xnor U11250 (N_11250,N_10943,N_10080);
xor U11251 (N_11251,N_10397,N_10824);
nor U11252 (N_11252,N_10168,N_10708);
nand U11253 (N_11253,N_10107,N_10550);
or U11254 (N_11254,N_10874,N_10113);
nand U11255 (N_11255,N_10083,N_10814);
nor U11256 (N_11256,N_10346,N_10978);
or U11257 (N_11257,N_10928,N_10979);
or U11258 (N_11258,N_10300,N_10199);
or U11259 (N_11259,N_10427,N_10838);
nor U11260 (N_11260,N_10672,N_10898);
or U11261 (N_11261,N_10064,N_10783);
or U11262 (N_11262,N_10197,N_10915);
and U11263 (N_11263,N_10394,N_10762);
and U11264 (N_11264,N_10245,N_10910);
or U11265 (N_11265,N_10354,N_10384);
or U11266 (N_11266,N_10473,N_10285);
and U11267 (N_11267,N_10046,N_10598);
and U11268 (N_11268,N_10927,N_10026);
and U11269 (N_11269,N_10950,N_10444);
or U11270 (N_11270,N_10362,N_10629);
or U11271 (N_11271,N_10322,N_10339);
nand U11272 (N_11272,N_10456,N_10985);
nand U11273 (N_11273,N_10952,N_10390);
nor U11274 (N_11274,N_10581,N_10380);
nand U11275 (N_11275,N_10051,N_10835);
and U11276 (N_11276,N_10387,N_10876);
or U11277 (N_11277,N_10055,N_10986);
nor U11278 (N_11278,N_10078,N_10683);
and U11279 (N_11279,N_10179,N_10893);
xnor U11280 (N_11280,N_10375,N_10531);
nand U11281 (N_11281,N_10402,N_10984);
nor U11282 (N_11282,N_10636,N_10196);
nor U11283 (N_11283,N_10867,N_10471);
nand U11284 (N_11284,N_10563,N_10997);
or U11285 (N_11285,N_10888,N_10159);
nor U11286 (N_11286,N_10165,N_10048);
xnor U11287 (N_11287,N_10174,N_10024);
nand U11288 (N_11288,N_10727,N_10903);
and U11289 (N_11289,N_10136,N_10939);
xnor U11290 (N_11290,N_10186,N_10694);
nor U11291 (N_11291,N_10616,N_10802);
or U11292 (N_11292,N_10142,N_10190);
or U11293 (N_11293,N_10454,N_10326);
and U11294 (N_11294,N_10892,N_10254);
nor U11295 (N_11295,N_10216,N_10577);
or U11296 (N_11296,N_10566,N_10594);
nor U11297 (N_11297,N_10099,N_10447);
nor U11298 (N_11298,N_10233,N_10842);
xor U11299 (N_11299,N_10982,N_10328);
and U11300 (N_11300,N_10170,N_10521);
nor U11301 (N_11301,N_10652,N_10352);
and U11302 (N_11302,N_10496,N_10056);
xnor U11303 (N_11303,N_10298,N_10667);
and U11304 (N_11304,N_10926,N_10686);
xnor U11305 (N_11305,N_10104,N_10082);
or U11306 (N_11306,N_10277,N_10689);
xnor U11307 (N_11307,N_10717,N_10061);
nor U11308 (N_11308,N_10239,N_10955);
xnor U11309 (N_11309,N_10506,N_10805);
or U11310 (N_11310,N_10625,N_10457);
and U11311 (N_11311,N_10215,N_10103);
and U11312 (N_11312,N_10831,N_10469);
and U11313 (N_11313,N_10654,N_10719);
nor U11314 (N_11314,N_10004,N_10585);
nor U11315 (N_11315,N_10299,N_10182);
and U11316 (N_11316,N_10000,N_10603);
xnor U11317 (N_11317,N_10336,N_10212);
nand U11318 (N_11318,N_10453,N_10758);
nor U11319 (N_11319,N_10150,N_10839);
nand U11320 (N_11320,N_10546,N_10739);
and U11321 (N_11321,N_10617,N_10037);
nand U11322 (N_11322,N_10247,N_10323);
xor U11323 (N_11323,N_10374,N_10483);
nand U11324 (N_11324,N_10685,N_10847);
or U11325 (N_11325,N_10991,N_10034);
nand U11326 (N_11326,N_10317,N_10596);
nor U11327 (N_11327,N_10679,N_10676);
nor U11328 (N_11328,N_10750,N_10671);
or U11329 (N_11329,N_10863,N_10614);
or U11330 (N_11330,N_10816,N_10069);
or U11331 (N_11331,N_10988,N_10633);
nor U11332 (N_11332,N_10331,N_10225);
or U11333 (N_11333,N_10237,N_10420);
nor U11334 (N_11334,N_10901,N_10178);
or U11335 (N_11335,N_10877,N_10741);
or U11336 (N_11336,N_10711,N_10851);
or U11337 (N_11337,N_10890,N_10250);
or U11338 (N_11338,N_10592,N_10309);
or U11339 (N_11339,N_10192,N_10539);
xnor U11340 (N_11340,N_10887,N_10017);
and U11341 (N_11341,N_10937,N_10648);
and U11342 (N_11342,N_10111,N_10868);
or U11343 (N_11343,N_10283,N_10275);
nand U11344 (N_11344,N_10923,N_10900);
nand U11345 (N_11345,N_10400,N_10644);
and U11346 (N_11346,N_10623,N_10746);
or U11347 (N_11347,N_10880,N_10255);
or U11348 (N_11348,N_10942,N_10446);
xor U11349 (N_11349,N_10602,N_10488);
and U11350 (N_11350,N_10002,N_10752);
or U11351 (N_11351,N_10859,N_10001);
xor U11352 (N_11352,N_10779,N_10388);
nor U11353 (N_11353,N_10830,N_10963);
and U11354 (N_11354,N_10249,N_10439);
nand U11355 (N_11355,N_10956,N_10959);
nor U11356 (N_11356,N_10540,N_10421);
or U11357 (N_11357,N_10569,N_10062);
and U11358 (N_11358,N_10517,N_10669);
nand U11359 (N_11359,N_10007,N_10382);
nor U11360 (N_11360,N_10008,N_10041);
nor U11361 (N_11361,N_10220,N_10127);
xor U11362 (N_11362,N_10638,N_10537);
nor U11363 (N_11363,N_10431,N_10405);
xor U11364 (N_11364,N_10709,N_10027);
xor U11365 (N_11365,N_10970,N_10050);
xor U11366 (N_11366,N_10491,N_10206);
nor U11367 (N_11367,N_10620,N_10369);
nand U11368 (N_11368,N_10761,N_10270);
nand U11369 (N_11369,N_10151,N_10117);
and U11370 (N_11370,N_10455,N_10657);
or U11371 (N_11371,N_10266,N_10999);
nor U11372 (N_11372,N_10492,N_10996);
nand U11373 (N_11373,N_10044,N_10555);
xor U11374 (N_11374,N_10889,N_10789);
or U11375 (N_11375,N_10974,N_10417);
or U11376 (N_11376,N_10995,N_10753);
and U11377 (N_11377,N_10902,N_10552);
and U11378 (N_11378,N_10497,N_10009);
and U11379 (N_11379,N_10631,N_10818);
or U11380 (N_11380,N_10406,N_10098);
nand U11381 (N_11381,N_10734,N_10878);
nand U11382 (N_11382,N_10074,N_10897);
nand U11383 (N_11383,N_10960,N_10184);
xor U11384 (N_11384,N_10886,N_10751);
or U11385 (N_11385,N_10541,N_10862);
nand U11386 (N_11386,N_10410,N_10251);
or U11387 (N_11387,N_10797,N_10140);
nor U11388 (N_11388,N_10272,N_10244);
and U11389 (N_11389,N_10304,N_10726);
and U11390 (N_11390,N_10193,N_10433);
nor U11391 (N_11391,N_10234,N_10664);
or U11392 (N_11392,N_10296,N_10424);
or U11393 (N_11393,N_10637,N_10873);
nor U11394 (N_11394,N_10784,N_10110);
nand U11395 (N_11395,N_10341,N_10696);
or U11396 (N_11396,N_10642,N_10228);
and U11397 (N_11397,N_10189,N_10395);
nand U11398 (N_11398,N_10858,N_10172);
or U11399 (N_11399,N_10010,N_10016);
xor U11400 (N_11400,N_10129,N_10333);
xor U11401 (N_11401,N_10567,N_10690);
nor U11402 (N_11402,N_10782,N_10634);
nand U11403 (N_11403,N_10154,N_10248);
xor U11404 (N_11404,N_10286,N_10848);
or U11405 (N_11405,N_10438,N_10315);
nand U11406 (N_11406,N_10302,N_10144);
xnor U11407 (N_11407,N_10962,N_10899);
and U11408 (N_11408,N_10365,N_10987);
nor U11409 (N_11409,N_10243,N_10489);
or U11410 (N_11410,N_10176,N_10965);
xor U11411 (N_11411,N_10023,N_10632);
nand U11412 (N_11412,N_10906,N_10320);
nor U11413 (N_11413,N_10775,N_10871);
or U11414 (N_11414,N_10194,N_10611);
nor U11415 (N_11415,N_10728,N_10951);
nand U11416 (N_11416,N_10121,N_10019);
and U11417 (N_11417,N_10745,N_10881);
or U11418 (N_11418,N_10126,N_10718);
xor U11419 (N_11419,N_10436,N_10053);
nand U11420 (N_11420,N_10716,N_10582);
and U11421 (N_11421,N_10946,N_10723);
nand U11422 (N_11422,N_10921,N_10470);
nand U11423 (N_11423,N_10449,N_10659);
nor U11424 (N_11424,N_10158,N_10949);
nand U11425 (N_11425,N_10003,N_10435);
xor U11426 (N_11426,N_10576,N_10378);
or U11427 (N_11427,N_10462,N_10622);
or U11428 (N_11428,N_10210,N_10790);
or U11429 (N_11429,N_10980,N_10626);
or U11430 (N_11430,N_10280,N_10348);
and U11431 (N_11431,N_10800,N_10869);
nor U11432 (N_11432,N_10776,N_10731);
xnor U11433 (N_11433,N_10738,N_10852);
nor U11434 (N_11434,N_10073,N_10732);
and U11435 (N_11435,N_10434,N_10057);
or U11436 (N_11436,N_10445,N_10371);
or U11437 (N_11437,N_10791,N_10486);
and U11438 (N_11438,N_10523,N_10133);
xor U11439 (N_11439,N_10613,N_10430);
nand U11440 (N_11440,N_10958,N_10287);
nor U11441 (N_11441,N_10258,N_10747);
nor U11442 (N_11442,N_10786,N_10141);
xor U11443 (N_11443,N_10660,N_10472);
xnor U11444 (N_11444,N_10658,N_10524);
xnor U11445 (N_11445,N_10870,N_10482);
xor U11446 (N_11446,N_10843,N_10437);
and U11447 (N_11447,N_10264,N_10072);
nor U11448 (N_11448,N_10459,N_10639);
and U11449 (N_11449,N_10699,N_10737);
nand U11450 (N_11450,N_10656,N_10381);
nand U11451 (N_11451,N_10640,N_10040);
and U11452 (N_11452,N_10022,N_10364);
xor U11453 (N_11453,N_10872,N_10833);
and U11454 (N_11454,N_10301,N_10090);
and U11455 (N_11455,N_10049,N_10290);
and U11456 (N_11456,N_10241,N_10363);
xor U11457 (N_11457,N_10904,N_10128);
and U11458 (N_11458,N_10218,N_10590);
or U11459 (N_11459,N_10770,N_10834);
nand U11460 (N_11460,N_10828,N_10112);
or U11461 (N_11461,N_10844,N_10807);
and U11462 (N_11462,N_10883,N_10227);
xnor U11463 (N_11463,N_10785,N_10559);
xor U11464 (N_11464,N_10177,N_10310);
or U11465 (N_11465,N_10688,N_10526);
and U11466 (N_11466,N_10418,N_10740);
and U11467 (N_11467,N_10512,N_10804);
nand U11468 (N_11468,N_10983,N_10448);
nor U11469 (N_11469,N_10502,N_10933);
and U11470 (N_11470,N_10917,N_10202);
and U11471 (N_11471,N_10548,N_10180);
and U11472 (N_11472,N_10964,N_10895);
nand U11473 (N_11473,N_10413,N_10349);
xnor U11474 (N_11474,N_10653,N_10773);
nor U11475 (N_11475,N_10554,N_10575);
xor U11476 (N_11476,N_10562,N_10832);
nor U11477 (N_11477,N_10338,N_10882);
xor U11478 (N_11478,N_10703,N_10075);
nand U11479 (N_11479,N_10408,N_10808);
nand U11480 (N_11480,N_10169,N_10066);
nand U11481 (N_11481,N_10086,N_10849);
or U11482 (N_11482,N_10071,N_10130);
xor U11483 (N_11483,N_10018,N_10564);
or U11484 (N_11484,N_10561,N_10419);
xor U11485 (N_11485,N_10840,N_10733);
and U11486 (N_11486,N_10570,N_10767);
or U11487 (N_11487,N_10586,N_10132);
xor U11488 (N_11488,N_10812,N_10230);
or U11489 (N_11489,N_10821,N_10428);
xnor U11490 (N_11490,N_10735,N_10757);
nor U11491 (N_11491,N_10068,N_10399);
or U11492 (N_11492,N_10827,N_10710);
nand U11493 (N_11493,N_10961,N_10217);
xor U11494 (N_11494,N_10607,N_10768);
and U11495 (N_11495,N_10100,N_10532);
nand U11496 (N_11496,N_10131,N_10908);
nor U11497 (N_11497,N_10316,N_10543);
nor U11498 (N_11498,N_10343,N_10748);
nor U11499 (N_11499,N_10279,N_10114);
nor U11500 (N_11500,N_10465,N_10263);
xor U11501 (N_11501,N_10166,N_10034);
nor U11502 (N_11502,N_10541,N_10763);
and U11503 (N_11503,N_10085,N_10591);
xnor U11504 (N_11504,N_10682,N_10524);
xor U11505 (N_11505,N_10355,N_10623);
and U11506 (N_11506,N_10979,N_10461);
nor U11507 (N_11507,N_10679,N_10192);
nand U11508 (N_11508,N_10496,N_10435);
nand U11509 (N_11509,N_10354,N_10038);
nand U11510 (N_11510,N_10631,N_10023);
or U11511 (N_11511,N_10850,N_10766);
or U11512 (N_11512,N_10634,N_10916);
and U11513 (N_11513,N_10991,N_10561);
nor U11514 (N_11514,N_10221,N_10723);
or U11515 (N_11515,N_10107,N_10726);
nand U11516 (N_11516,N_10806,N_10422);
nor U11517 (N_11517,N_10245,N_10422);
nand U11518 (N_11518,N_10435,N_10262);
or U11519 (N_11519,N_10090,N_10324);
nand U11520 (N_11520,N_10811,N_10695);
and U11521 (N_11521,N_10091,N_10019);
xor U11522 (N_11522,N_10766,N_10556);
or U11523 (N_11523,N_10955,N_10669);
or U11524 (N_11524,N_10653,N_10153);
xor U11525 (N_11525,N_10380,N_10421);
nand U11526 (N_11526,N_10205,N_10755);
or U11527 (N_11527,N_10775,N_10266);
and U11528 (N_11528,N_10506,N_10241);
xnor U11529 (N_11529,N_10979,N_10468);
xor U11530 (N_11530,N_10689,N_10535);
nand U11531 (N_11531,N_10226,N_10771);
or U11532 (N_11532,N_10970,N_10431);
nand U11533 (N_11533,N_10209,N_10696);
nand U11534 (N_11534,N_10237,N_10699);
xor U11535 (N_11535,N_10456,N_10706);
or U11536 (N_11536,N_10438,N_10386);
xnor U11537 (N_11537,N_10312,N_10687);
nand U11538 (N_11538,N_10737,N_10978);
and U11539 (N_11539,N_10777,N_10355);
or U11540 (N_11540,N_10701,N_10922);
and U11541 (N_11541,N_10873,N_10446);
xnor U11542 (N_11542,N_10687,N_10799);
or U11543 (N_11543,N_10111,N_10397);
nand U11544 (N_11544,N_10473,N_10982);
and U11545 (N_11545,N_10726,N_10933);
nand U11546 (N_11546,N_10292,N_10782);
xnor U11547 (N_11547,N_10180,N_10055);
nand U11548 (N_11548,N_10766,N_10640);
nor U11549 (N_11549,N_10831,N_10862);
and U11550 (N_11550,N_10819,N_10334);
nor U11551 (N_11551,N_10416,N_10805);
nand U11552 (N_11552,N_10425,N_10017);
nor U11553 (N_11553,N_10790,N_10792);
and U11554 (N_11554,N_10761,N_10956);
nand U11555 (N_11555,N_10052,N_10989);
or U11556 (N_11556,N_10677,N_10260);
nor U11557 (N_11557,N_10666,N_10140);
nand U11558 (N_11558,N_10484,N_10430);
or U11559 (N_11559,N_10298,N_10973);
xnor U11560 (N_11560,N_10457,N_10114);
and U11561 (N_11561,N_10204,N_10647);
nand U11562 (N_11562,N_10864,N_10796);
and U11563 (N_11563,N_10304,N_10753);
or U11564 (N_11564,N_10962,N_10405);
nor U11565 (N_11565,N_10727,N_10741);
nand U11566 (N_11566,N_10849,N_10124);
or U11567 (N_11567,N_10585,N_10264);
or U11568 (N_11568,N_10735,N_10673);
nand U11569 (N_11569,N_10988,N_10430);
xnor U11570 (N_11570,N_10278,N_10934);
xnor U11571 (N_11571,N_10271,N_10820);
or U11572 (N_11572,N_10790,N_10925);
xor U11573 (N_11573,N_10558,N_10354);
xnor U11574 (N_11574,N_10403,N_10985);
and U11575 (N_11575,N_10944,N_10577);
or U11576 (N_11576,N_10421,N_10065);
and U11577 (N_11577,N_10477,N_10934);
and U11578 (N_11578,N_10272,N_10448);
nor U11579 (N_11579,N_10631,N_10270);
nand U11580 (N_11580,N_10290,N_10503);
nor U11581 (N_11581,N_10159,N_10004);
and U11582 (N_11582,N_10735,N_10785);
nor U11583 (N_11583,N_10436,N_10070);
nor U11584 (N_11584,N_10377,N_10954);
xnor U11585 (N_11585,N_10683,N_10336);
nand U11586 (N_11586,N_10985,N_10296);
xor U11587 (N_11587,N_10177,N_10415);
xnor U11588 (N_11588,N_10831,N_10736);
xor U11589 (N_11589,N_10456,N_10396);
nor U11590 (N_11590,N_10526,N_10508);
or U11591 (N_11591,N_10457,N_10324);
nor U11592 (N_11592,N_10428,N_10717);
xor U11593 (N_11593,N_10528,N_10164);
nor U11594 (N_11594,N_10201,N_10653);
and U11595 (N_11595,N_10744,N_10630);
xor U11596 (N_11596,N_10111,N_10005);
xnor U11597 (N_11597,N_10352,N_10904);
and U11598 (N_11598,N_10617,N_10775);
xnor U11599 (N_11599,N_10895,N_10540);
or U11600 (N_11600,N_10996,N_10852);
and U11601 (N_11601,N_10895,N_10458);
nand U11602 (N_11602,N_10960,N_10026);
nor U11603 (N_11603,N_10123,N_10441);
xnor U11604 (N_11604,N_10482,N_10779);
or U11605 (N_11605,N_10591,N_10713);
or U11606 (N_11606,N_10301,N_10944);
or U11607 (N_11607,N_10098,N_10028);
nand U11608 (N_11608,N_10975,N_10564);
nor U11609 (N_11609,N_10964,N_10561);
nor U11610 (N_11610,N_10469,N_10743);
nor U11611 (N_11611,N_10364,N_10308);
nor U11612 (N_11612,N_10413,N_10817);
or U11613 (N_11613,N_10292,N_10415);
nor U11614 (N_11614,N_10761,N_10821);
xnor U11615 (N_11615,N_10430,N_10345);
and U11616 (N_11616,N_10344,N_10672);
nor U11617 (N_11617,N_10508,N_10468);
xor U11618 (N_11618,N_10328,N_10281);
or U11619 (N_11619,N_10016,N_10948);
and U11620 (N_11620,N_10156,N_10500);
nor U11621 (N_11621,N_10137,N_10176);
nor U11622 (N_11622,N_10160,N_10033);
nand U11623 (N_11623,N_10664,N_10195);
nand U11624 (N_11624,N_10910,N_10291);
nand U11625 (N_11625,N_10076,N_10090);
nor U11626 (N_11626,N_10853,N_10267);
xnor U11627 (N_11627,N_10893,N_10976);
and U11628 (N_11628,N_10529,N_10605);
and U11629 (N_11629,N_10517,N_10888);
and U11630 (N_11630,N_10060,N_10813);
xnor U11631 (N_11631,N_10872,N_10405);
nor U11632 (N_11632,N_10445,N_10144);
nand U11633 (N_11633,N_10392,N_10563);
and U11634 (N_11634,N_10286,N_10120);
nor U11635 (N_11635,N_10854,N_10249);
or U11636 (N_11636,N_10559,N_10784);
nor U11637 (N_11637,N_10901,N_10478);
nor U11638 (N_11638,N_10549,N_10413);
or U11639 (N_11639,N_10095,N_10262);
and U11640 (N_11640,N_10151,N_10730);
xnor U11641 (N_11641,N_10205,N_10229);
nor U11642 (N_11642,N_10482,N_10639);
and U11643 (N_11643,N_10063,N_10673);
or U11644 (N_11644,N_10826,N_10159);
nor U11645 (N_11645,N_10263,N_10204);
or U11646 (N_11646,N_10938,N_10557);
nand U11647 (N_11647,N_10688,N_10006);
and U11648 (N_11648,N_10088,N_10878);
nand U11649 (N_11649,N_10908,N_10037);
or U11650 (N_11650,N_10444,N_10722);
and U11651 (N_11651,N_10574,N_10234);
xor U11652 (N_11652,N_10862,N_10413);
or U11653 (N_11653,N_10730,N_10685);
nor U11654 (N_11654,N_10864,N_10179);
or U11655 (N_11655,N_10238,N_10822);
and U11656 (N_11656,N_10517,N_10587);
xor U11657 (N_11657,N_10034,N_10033);
nor U11658 (N_11658,N_10946,N_10005);
xnor U11659 (N_11659,N_10699,N_10883);
nand U11660 (N_11660,N_10546,N_10623);
xnor U11661 (N_11661,N_10119,N_10860);
nand U11662 (N_11662,N_10799,N_10600);
xor U11663 (N_11663,N_10049,N_10599);
nand U11664 (N_11664,N_10603,N_10074);
or U11665 (N_11665,N_10966,N_10079);
nor U11666 (N_11666,N_10052,N_10160);
nand U11667 (N_11667,N_10669,N_10355);
nor U11668 (N_11668,N_10837,N_10269);
nand U11669 (N_11669,N_10127,N_10839);
and U11670 (N_11670,N_10085,N_10072);
or U11671 (N_11671,N_10060,N_10854);
nand U11672 (N_11672,N_10640,N_10627);
nand U11673 (N_11673,N_10312,N_10878);
and U11674 (N_11674,N_10586,N_10009);
nor U11675 (N_11675,N_10678,N_10145);
nand U11676 (N_11676,N_10377,N_10200);
nand U11677 (N_11677,N_10995,N_10168);
xnor U11678 (N_11678,N_10530,N_10528);
nand U11679 (N_11679,N_10039,N_10972);
or U11680 (N_11680,N_10057,N_10017);
or U11681 (N_11681,N_10705,N_10314);
xnor U11682 (N_11682,N_10361,N_10800);
and U11683 (N_11683,N_10325,N_10146);
or U11684 (N_11684,N_10623,N_10966);
nor U11685 (N_11685,N_10755,N_10398);
nand U11686 (N_11686,N_10163,N_10204);
nor U11687 (N_11687,N_10781,N_10682);
nand U11688 (N_11688,N_10270,N_10357);
nor U11689 (N_11689,N_10574,N_10749);
nor U11690 (N_11690,N_10173,N_10563);
or U11691 (N_11691,N_10510,N_10670);
and U11692 (N_11692,N_10432,N_10343);
nor U11693 (N_11693,N_10143,N_10518);
and U11694 (N_11694,N_10106,N_10826);
xnor U11695 (N_11695,N_10564,N_10760);
or U11696 (N_11696,N_10458,N_10272);
nor U11697 (N_11697,N_10192,N_10628);
nand U11698 (N_11698,N_10856,N_10453);
xor U11699 (N_11699,N_10095,N_10670);
xnor U11700 (N_11700,N_10727,N_10793);
or U11701 (N_11701,N_10947,N_10793);
and U11702 (N_11702,N_10894,N_10294);
and U11703 (N_11703,N_10495,N_10394);
nand U11704 (N_11704,N_10783,N_10231);
and U11705 (N_11705,N_10914,N_10514);
nand U11706 (N_11706,N_10408,N_10663);
or U11707 (N_11707,N_10694,N_10460);
xnor U11708 (N_11708,N_10710,N_10913);
nand U11709 (N_11709,N_10674,N_10637);
or U11710 (N_11710,N_10914,N_10674);
and U11711 (N_11711,N_10927,N_10905);
nand U11712 (N_11712,N_10910,N_10386);
or U11713 (N_11713,N_10192,N_10973);
or U11714 (N_11714,N_10052,N_10352);
nor U11715 (N_11715,N_10326,N_10075);
nor U11716 (N_11716,N_10313,N_10462);
nand U11717 (N_11717,N_10713,N_10232);
and U11718 (N_11718,N_10984,N_10193);
and U11719 (N_11719,N_10303,N_10415);
nand U11720 (N_11720,N_10561,N_10744);
or U11721 (N_11721,N_10403,N_10362);
or U11722 (N_11722,N_10212,N_10057);
xor U11723 (N_11723,N_10998,N_10444);
nand U11724 (N_11724,N_10937,N_10503);
nand U11725 (N_11725,N_10901,N_10870);
nor U11726 (N_11726,N_10601,N_10276);
or U11727 (N_11727,N_10597,N_10021);
nor U11728 (N_11728,N_10781,N_10620);
and U11729 (N_11729,N_10847,N_10571);
and U11730 (N_11730,N_10214,N_10240);
and U11731 (N_11731,N_10404,N_10438);
and U11732 (N_11732,N_10194,N_10122);
or U11733 (N_11733,N_10011,N_10471);
nor U11734 (N_11734,N_10227,N_10249);
nor U11735 (N_11735,N_10516,N_10200);
xnor U11736 (N_11736,N_10263,N_10616);
xor U11737 (N_11737,N_10101,N_10644);
nand U11738 (N_11738,N_10695,N_10873);
xor U11739 (N_11739,N_10664,N_10681);
or U11740 (N_11740,N_10507,N_10142);
or U11741 (N_11741,N_10525,N_10170);
xnor U11742 (N_11742,N_10323,N_10611);
nor U11743 (N_11743,N_10130,N_10867);
nand U11744 (N_11744,N_10181,N_10644);
and U11745 (N_11745,N_10421,N_10462);
nor U11746 (N_11746,N_10238,N_10824);
and U11747 (N_11747,N_10624,N_10686);
nor U11748 (N_11748,N_10211,N_10147);
xnor U11749 (N_11749,N_10282,N_10224);
or U11750 (N_11750,N_10632,N_10308);
and U11751 (N_11751,N_10673,N_10402);
and U11752 (N_11752,N_10228,N_10476);
or U11753 (N_11753,N_10448,N_10745);
nor U11754 (N_11754,N_10566,N_10298);
xor U11755 (N_11755,N_10151,N_10096);
nand U11756 (N_11756,N_10758,N_10846);
nor U11757 (N_11757,N_10130,N_10774);
nand U11758 (N_11758,N_10824,N_10862);
nand U11759 (N_11759,N_10826,N_10799);
nand U11760 (N_11760,N_10417,N_10148);
nor U11761 (N_11761,N_10032,N_10926);
nand U11762 (N_11762,N_10769,N_10873);
nor U11763 (N_11763,N_10437,N_10124);
nand U11764 (N_11764,N_10230,N_10752);
xor U11765 (N_11765,N_10775,N_10416);
nand U11766 (N_11766,N_10097,N_10459);
nand U11767 (N_11767,N_10924,N_10833);
and U11768 (N_11768,N_10125,N_10575);
nor U11769 (N_11769,N_10925,N_10243);
xor U11770 (N_11770,N_10347,N_10605);
nand U11771 (N_11771,N_10768,N_10215);
and U11772 (N_11772,N_10688,N_10197);
nand U11773 (N_11773,N_10957,N_10455);
nor U11774 (N_11774,N_10531,N_10281);
or U11775 (N_11775,N_10807,N_10904);
xnor U11776 (N_11776,N_10920,N_10909);
xnor U11777 (N_11777,N_10518,N_10770);
nand U11778 (N_11778,N_10175,N_10465);
xor U11779 (N_11779,N_10201,N_10467);
xor U11780 (N_11780,N_10220,N_10197);
or U11781 (N_11781,N_10808,N_10847);
nand U11782 (N_11782,N_10819,N_10738);
nand U11783 (N_11783,N_10350,N_10282);
and U11784 (N_11784,N_10224,N_10650);
nor U11785 (N_11785,N_10199,N_10034);
nor U11786 (N_11786,N_10430,N_10483);
xor U11787 (N_11787,N_10820,N_10772);
xnor U11788 (N_11788,N_10235,N_10267);
and U11789 (N_11789,N_10807,N_10278);
nand U11790 (N_11790,N_10402,N_10706);
nand U11791 (N_11791,N_10817,N_10644);
xnor U11792 (N_11792,N_10410,N_10276);
xor U11793 (N_11793,N_10749,N_10457);
nand U11794 (N_11794,N_10633,N_10833);
or U11795 (N_11795,N_10637,N_10422);
or U11796 (N_11796,N_10376,N_10167);
nor U11797 (N_11797,N_10360,N_10241);
or U11798 (N_11798,N_10250,N_10816);
and U11799 (N_11799,N_10165,N_10718);
or U11800 (N_11800,N_10479,N_10592);
or U11801 (N_11801,N_10317,N_10359);
and U11802 (N_11802,N_10908,N_10050);
or U11803 (N_11803,N_10883,N_10687);
nand U11804 (N_11804,N_10157,N_10561);
xor U11805 (N_11805,N_10151,N_10511);
or U11806 (N_11806,N_10203,N_10738);
or U11807 (N_11807,N_10775,N_10884);
nor U11808 (N_11808,N_10901,N_10915);
nand U11809 (N_11809,N_10166,N_10066);
and U11810 (N_11810,N_10140,N_10589);
or U11811 (N_11811,N_10775,N_10338);
nor U11812 (N_11812,N_10423,N_10133);
nand U11813 (N_11813,N_10444,N_10084);
or U11814 (N_11814,N_10597,N_10164);
or U11815 (N_11815,N_10100,N_10114);
xor U11816 (N_11816,N_10172,N_10953);
xor U11817 (N_11817,N_10709,N_10771);
and U11818 (N_11818,N_10142,N_10476);
or U11819 (N_11819,N_10334,N_10839);
xor U11820 (N_11820,N_10995,N_10752);
or U11821 (N_11821,N_10842,N_10969);
or U11822 (N_11822,N_10797,N_10428);
nand U11823 (N_11823,N_10373,N_10500);
nor U11824 (N_11824,N_10749,N_10077);
nand U11825 (N_11825,N_10638,N_10932);
xnor U11826 (N_11826,N_10864,N_10959);
nor U11827 (N_11827,N_10954,N_10061);
or U11828 (N_11828,N_10552,N_10875);
xnor U11829 (N_11829,N_10935,N_10536);
or U11830 (N_11830,N_10523,N_10387);
nor U11831 (N_11831,N_10145,N_10928);
nand U11832 (N_11832,N_10758,N_10151);
or U11833 (N_11833,N_10632,N_10685);
xor U11834 (N_11834,N_10111,N_10622);
xor U11835 (N_11835,N_10970,N_10817);
and U11836 (N_11836,N_10472,N_10174);
nand U11837 (N_11837,N_10058,N_10274);
nor U11838 (N_11838,N_10716,N_10038);
xnor U11839 (N_11839,N_10608,N_10368);
xor U11840 (N_11840,N_10314,N_10541);
nor U11841 (N_11841,N_10455,N_10735);
or U11842 (N_11842,N_10303,N_10906);
nor U11843 (N_11843,N_10568,N_10378);
xnor U11844 (N_11844,N_10311,N_10029);
nand U11845 (N_11845,N_10925,N_10022);
nor U11846 (N_11846,N_10639,N_10024);
xor U11847 (N_11847,N_10869,N_10477);
nor U11848 (N_11848,N_10481,N_10848);
and U11849 (N_11849,N_10465,N_10542);
nand U11850 (N_11850,N_10986,N_10783);
xor U11851 (N_11851,N_10646,N_10660);
and U11852 (N_11852,N_10850,N_10411);
xor U11853 (N_11853,N_10205,N_10250);
and U11854 (N_11854,N_10801,N_10675);
xor U11855 (N_11855,N_10645,N_10138);
or U11856 (N_11856,N_10015,N_10142);
nor U11857 (N_11857,N_10213,N_10720);
nor U11858 (N_11858,N_10722,N_10769);
and U11859 (N_11859,N_10996,N_10701);
nand U11860 (N_11860,N_10053,N_10589);
or U11861 (N_11861,N_10465,N_10400);
and U11862 (N_11862,N_10646,N_10618);
nand U11863 (N_11863,N_10318,N_10143);
or U11864 (N_11864,N_10131,N_10099);
or U11865 (N_11865,N_10696,N_10197);
nand U11866 (N_11866,N_10366,N_10624);
or U11867 (N_11867,N_10738,N_10610);
nand U11868 (N_11868,N_10983,N_10905);
and U11869 (N_11869,N_10184,N_10047);
nor U11870 (N_11870,N_10793,N_10798);
xor U11871 (N_11871,N_10844,N_10641);
xnor U11872 (N_11872,N_10282,N_10929);
nand U11873 (N_11873,N_10336,N_10512);
nor U11874 (N_11874,N_10879,N_10186);
nor U11875 (N_11875,N_10463,N_10248);
nand U11876 (N_11876,N_10455,N_10312);
and U11877 (N_11877,N_10808,N_10127);
and U11878 (N_11878,N_10625,N_10263);
nor U11879 (N_11879,N_10286,N_10913);
nor U11880 (N_11880,N_10780,N_10541);
nand U11881 (N_11881,N_10294,N_10843);
and U11882 (N_11882,N_10108,N_10456);
or U11883 (N_11883,N_10968,N_10716);
or U11884 (N_11884,N_10888,N_10980);
xnor U11885 (N_11885,N_10272,N_10652);
and U11886 (N_11886,N_10897,N_10059);
nand U11887 (N_11887,N_10794,N_10485);
nor U11888 (N_11888,N_10202,N_10739);
nor U11889 (N_11889,N_10861,N_10248);
and U11890 (N_11890,N_10495,N_10266);
or U11891 (N_11891,N_10361,N_10025);
nand U11892 (N_11892,N_10614,N_10110);
xnor U11893 (N_11893,N_10203,N_10845);
nand U11894 (N_11894,N_10264,N_10837);
or U11895 (N_11895,N_10648,N_10774);
and U11896 (N_11896,N_10631,N_10443);
nor U11897 (N_11897,N_10674,N_10467);
xor U11898 (N_11898,N_10376,N_10612);
nor U11899 (N_11899,N_10820,N_10084);
xnor U11900 (N_11900,N_10019,N_10654);
and U11901 (N_11901,N_10247,N_10606);
nand U11902 (N_11902,N_10352,N_10079);
xnor U11903 (N_11903,N_10284,N_10753);
or U11904 (N_11904,N_10387,N_10861);
or U11905 (N_11905,N_10142,N_10969);
nand U11906 (N_11906,N_10765,N_10306);
xnor U11907 (N_11907,N_10038,N_10012);
and U11908 (N_11908,N_10124,N_10990);
or U11909 (N_11909,N_10884,N_10358);
nand U11910 (N_11910,N_10655,N_10965);
xor U11911 (N_11911,N_10392,N_10244);
and U11912 (N_11912,N_10526,N_10689);
and U11913 (N_11913,N_10401,N_10193);
nand U11914 (N_11914,N_10149,N_10480);
xor U11915 (N_11915,N_10822,N_10546);
and U11916 (N_11916,N_10611,N_10203);
nand U11917 (N_11917,N_10258,N_10033);
nand U11918 (N_11918,N_10394,N_10486);
xnor U11919 (N_11919,N_10062,N_10013);
xnor U11920 (N_11920,N_10296,N_10873);
xnor U11921 (N_11921,N_10300,N_10707);
nor U11922 (N_11922,N_10483,N_10941);
or U11923 (N_11923,N_10362,N_10273);
nor U11924 (N_11924,N_10602,N_10774);
nand U11925 (N_11925,N_10895,N_10070);
nor U11926 (N_11926,N_10571,N_10073);
nor U11927 (N_11927,N_10259,N_10908);
or U11928 (N_11928,N_10689,N_10832);
xor U11929 (N_11929,N_10105,N_10237);
or U11930 (N_11930,N_10716,N_10560);
nand U11931 (N_11931,N_10445,N_10562);
nand U11932 (N_11932,N_10480,N_10550);
xor U11933 (N_11933,N_10476,N_10215);
xnor U11934 (N_11934,N_10277,N_10928);
nand U11935 (N_11935,N_10821,N_10009);
and U11936 (N_11936,N_10977,N_10859);
nand U11937 (N_11937,N_10316,N_10458);
nor U11938 (N_11938,N_10773,N_10651);
or U11939 (N_11939,N_10225,N_10099);
nor U11940 (N_11940,N_10999,N_10611);
nor U11941 (N_11941,N_10681,N_10167);
and U11942 (N_11942,N_10210,N_10020);
or U11943 (N_11943,N_10323,N_10204);
nand U11944 (N_11944,N_10889,N_10391);
or U11945 (N_11945,N_10249,N_10430);
and U11946 (N_11946,N_10520,N_10865);
or U11947 (N_11947,N_10445,N_10218);
nor U11948 (N_11948,N_10762,N_10808);
or U11949 (N_11949,N_10444,N_10944);
xor U11950 (N_11950,N_10082,N_10240);
and U11951 (N_11951,N_10824,N_10661);
xor U11952 (N_11952,N_10675,N_10734);
xnor U11953 (N_11953,N_10702,N_10765);
xor U11954 (N_11954,N_10842,N_10966);
nand U11955 (N_11955,N_10514,N_10706);
nand U11956 (N_11956,N_10866,N_10295);
or U11957 (N_11957,N_10574,N_10249);
and U11958 (N_11958,N_10764,N_10401);
nor U11959 (N_11959,N_10907,N_10657);
and U11960 (N_11960,N_10331,N_10594);
and U11961 (N_11961,N_10931,N_10810);
or U11962 (N_11962,N_10337,N_10890);
nand U11963 (N_11963,N_10539,N_10628);
and U11964 (N_11964,N_10148,N_10550);
nand U11965 (N_11965,N_10690,N_10545);
or U11966 (N_11966,N_10275,N_10847);
or U11967 (N_11967,N_10263,N_10415);
or U11968 (N_11968,N_10750,N_10292);
xor U11969 (N_11969,N_10350,N_10628);
nor U11970 (N_11970,N_10434,N_10698);
nand U11971 (N_11971,N_10187,N_10496);
nand U11972 (N_11972,N_10220,N_10587);
xor U11973 (N_11973,N_10439,N_10754);
nand U11974 (N_11974,N_10614,N_10822);
or U11975 (N_11975,N_10042,N_10090);
xnor U11976 (N_11976,N_10774,N_10040);
nor U11977 (N_11977,N_10491,N_10245);
nor U11978 (N_11978,N_10710,N_10959);
xor U11979 (N_11979,N_10568,N_10916);
xnor U11980 (N_11980,N_10492,N_10121);
or U11981 (N_11981,N_10179,N_10074);
nor U11982 (N_11982,N_10728,N_10766);
nand U11983 (N_11983,N_10297,N_10849);
nand U11984 (N_11984,N_10011,N_10957);
and U11985 (N_11985,N_10202,N_10217);
and U11986 (N_11986,N_10840,N_10808);
and U11987 (N_11987,N_10478,N_10430);
nor U11988 (N_11988,N_10976,N_10576);
xnor U11989 (N_11989,N_10869,N_10471);
xor U11990 (N_11990,N_10169,N_10429);
nor U11991 (N_11991,N_10746,N_10407);
and U11992 (N_11992,N_10218,N_10487);
xor U11993 (N_11993,N_10985,N_10712);
and U11994 (N_11994,N_10533,N_10560);
nor U11995 (N_11995,N_10226,N_10125);
and U11996 (N_11996,N_10855,N_10095);
nor U11997 (N_11997,N_10652,N_10817);
nor U11998 (N_11998,N_10174,N_10947);
nand U11999 (N_11999,N_10197,N_10548);
nor U12000 (N_12000,N_11482,N_11773);
or U12001 (N_12001,N_11040,N_11736);
xor U12002 (N_12002,N_11515,N_11004);
or U12003 (N_12003,N_11357,N_11119);
xor U12004 (N_12004,N_11355,N_11408);
xor U12005 (N_12005,N_11940,N_11218);
nor U12006 (N_12006,N_11972,N_11808);
nand U12007 (N_12007,N_11688,N_11265);
nor U12008 (N_12008,N_11652,N_11693);
xnor U12009 (N_12009,N_11700,N_11985);
nor U12010 (N_12010,N_11673,N_11026);
nand U12011 (N_12011,N_11557,N_11713);
xor U12012 (N_12012,N_11551,N_11781);
or U12013 (N_12013,N_11451,N_11181);
and U12014 (N_12014,N_11588,N_11734);
nand U12015 (N_12015,N_11943,N_11749);
and U12016 (N_12016,N_11886,N_11827);
nor U12017 (N_12017,N_11592,N_11829);
nand U12018 (N_12018,N_11891,N_11812);
or U12019 (N_12019,N_11223,N_11144);
or U12020 (N_12020,N_11718,N_11473);
nand U12021 (N_12021,N_11686,N_11976);
nand U12022 (N_12022,N_11330,N_11431);
or U12023 (N_12023,N_11619,N_11702);
nand U12024 (N_12024,N_11649,N_11971);
and U12025 (N_12025,N_11798,N_11082);
nand U12026 (N_12026,N_11487,N_11175);
nand U12027 (N_12027,N_11504,N_11725);
and U12028 (N_12028,N_11080,N_11358);
and U12029 (N_12029,N_11994,N_11521);
or U12030 (N_12030,N_11574,N_11010);
or U12031 (N_12031,N_11951,N_11429);
or U12032 (N_12032,N_11348,N_11782);
xnor U12033 (N_12033,N_11586,N_11165);
or U12034 (N_12034,N_11529,N_11347);
or U12035 (N_12035,N_11623,N_11655);
nand U12036 (N_12036,N_11048,N_11785);
xnor U12037 (N_12037,N_11635,N_11682);
or U12038 (N_12038,N_11957,N_11792);
nand U12039 (N_12039,N_11836,N_11484);
and U12040 (N_12040,N_11721,N_11398);
xnor U12041 (N_12041,N_11579,N_11290);
nand U12042 (N_12042,N_11367,N_11970);
or U12043 (N_12043,N_11411,N_11662);
and U12044 (N_12044,N_11853,N_11434);
and U12045 (N_12045,N_11488,N_11661);
nor U12046 (N_12046,N_11747,N_11844);
nand U12047 (N_12047,N_11818,N_11506);
nand U12048 (N_12048,N_11240,N_11717);
xnor U12049 (N_12049,N_11086,N_11560);
xor U12050 (N_12050,N_11025,N_11136);
nand U12051 (N_12051,N_11415,N_11980);
or U12052 (N_12052,N_11116,N_11227);
nor U12053 (N_12053,N_11149,N_11877);
xnor U12054 (N_12054,N_11582,N_11556);
or U12055 (N_12055,N_11780,N_11385);
and U12056 (N_12056,N_11069,N_11106);
nand U12057 (N_12057,N_11340,N_11778);
or U12058 (N_12058,N_11030,N_11637);
nor U12059 (N_12059,N_11044,N_11805);
xnor U12060 (N_12060,N_11728,N_11407);
nor U12061 (N_12061,N_11283,N_11452);
xnor U12062 (N_12062,N_11685,N_11823);
xnor U12063 (N_12063,N_11032,N_11413);
nand U12064 (N_12064,N_11249,N_11930);
xnor U12065 (N_12065,N_11237,N_11189);
nand U12066 (N_12066,N_11102,N_11876);
or U12067 (N_12067,N_11199,N_11169);
xnor U12068 (N_12068,N_11672,N_11308);
xnor U12069 (N_12069,N_11809,N_11097);
nand U12070 (N_12070,N_11883,N_11268);
and U12071 (N_12071,N_11936,N_11578);
and U12072 (N_12072,N_11183,N_11027);
or U12073 (N_12073,N_11915,N_11279);
xnor U12074 (N_12074,N_11111,N_11335);
nand U12075 (N_12075,N_11628,N_11790);
nor U12076 (N_12076,N_11042,N_11210);
nand U12077 (N_12077,N_11527,N_11548);
or U12078 (N_12078,N_11315,N_11377);
and U12079 (N_12079,N_11676,N_11599);
nand U12080 (N_12080,N_11061,N_11365);
nor U12081 (N_12081,N_11570,N_11863);
xnor U12082 (N_12082,N_11336,N_11703);
nand U12083 (N_12083,N_11595,N_11138);
or U12084 (N_12084,N_11674,N_11607);
or U12085 (N_12085,N_11076,N_11437);
nand U12086 (N_12086,N_11494,N_11624);
nand U12087 (N_12087,N_11765,N_11617);
xnor U12088 (N_12088,N_11612,N_11501);
xnor U12089 (N_12089,N_11948,N_11726);
nand U12090 (N_12090,N_11945,N_11788);
and U12091 (N_12091,N_11926,N_11650);
nand U12092 (N_12092,N_11294,N_11195);
or U12093 (N_12093,N_11744,N_11067);
xnor U12094 (N_12094,N_11046,N_11857);
and U12095 (N_12095,N_11850,N_11982);
or U12096 (N_12096,N_11689,N_11735);
and U12097 (N_12097,N_11796,N_11683);
nor U12098 (N_12098,N_11397,N_11271);
nor U12099 (N_12099,N_11799,N_11510);
nor U12100 (N_12100,N_11309,N_11284);
xor U12101 (N_12101,N_11239,N_11803);
nor U12102 (N_12102,N_11854,N_11573);
nand U12103 (N_12103,N_11432,N_11712);
xor U12104 (N_12104,N_11167,N_11896);
or U12105 (N_12105,N_11626,N_11561);
nor U12106 (N_12106,N_11889,N_11491);
or U12107 (N_12107,N_11225,N_11420);
nor U12108 (N_12108,N_11015,N_11742);
nand U12109 (N_12109,N_11000,N_11485);
nand U12110 (N_12110,N_11659,N_11384);
or U12111 (N_12111,N_11601,N_11632);
nor U12112 (N_12112,N_11989,N_11990);
nor U12113 (N_12113,N_11418,N_11478);
xnor U12114 (N_12114,N_11641,N_11691);
nor U12115 (N_12115,N_11993,N_11983);
xor U12116 (N_12116,N_11421,N_11664);
or U12117 (N_12117,N_11344,N_11159);
nand U12118 (N_12118,N_11648,N_11060);
nand U12119 (N_12119,N_11255,N_11250);
nand U12120 (N_12120,N_11304,N_11753);
and U12121 (N_12121,N_11852,N_11746);
or U12122 (N_12122,N_11419,N_11562);
nor U12123 (N_12123,N_11401,N_11963);
nor U12124 (N_12124,N_11145,N_11459);
nor U12125 (N_12125,N_11122,N_11640);
and U12126 (N_12126,N_11558,N_11550);
nor U12127 (N_12127,N_11858,N_11542);
nand U12128 (N_12128,N_11848,N_11037);
nor U12129 (N_12129,N_11366,N_11028);
nor U12130 (N_12130,N_11467,N_11709);
nand U12131 (N_12131,N_11953,N_11197);
or U12132 (N_12132,N_11179,N_11811);
nand U12133 (N_12133,N_11828,N_11361);
xor U12134 (N_12134,N_11532,N_11156);
xnor U12135 (N_12135,N_11687,N_11492);
xnor U12136 (N_12136,N_11834,N_11651);
xor U12137 (N_12137,N_11740,N_11902);
and U12138 (N_12138,N_11621,N_11928);
or U12139 (N_12139,N_11656,N_11139);
xnor U12140 (N_12140,N_11133,N_11598);
or U12141 (N_12141,N_11405,N_11517);
nand U12142 (N_12142,N_11207,N_11666);
or U12143 (N_12143,N_11203,N_11917);
or U12144 (N_12144,N_11302,N_11898);
xor U12145 (N_12145,N_11813,N_11938);
nand U12146 (N_12146,N_11722,N_11113);
and U12147 (N_12147,N_11184,N_11233);
nor U12148 (N_12148,N_11056,N_11444);
nor U12149 (N_12149,N_11552,N_11751);
nor U12150 (N_12150,N_11826,N_11801);
and U12151 (N_12151,N_11705,N_11738);
nor U12152 (N_12152,N_11150,N_11732);
nand U12153 (N_12153,N_11918,N_11331);
xor U12154 (N_12154,N_11312,N_11049);
nand U12155 (N_12155,N_11380,N_11777);
or U12156 (N_12156,N_11600,N_11499);
nor U12157 (N_12157,N_11537,N_11988);
or U12158 (N_12158,N_11837,N_11845);
and U12159 (N_12159,N_11232,N_11081);
nor U12160 (N_12160,N_11404,N_11412);
xor U12161 (N_12161,N_11849,N_11638);
nor U12162 (N_12162,N_11514,N_11783);
and U12163 (N_12163,N_11533,N_11229);
nor U12164 (N_12164,N_11320,N_11645);
nand U12165 (N_12165,N_11329,N_11003);
and U12166 (N_12166,N_11422,N_11544);
or U12167 (N_12167,N_11964,N_11314);
nand U12168 (N_12168,N_11919,N_11436);
xnor U12169 (N_12169,N_11251,N_11425);
and U12170 (N_12170,N_11956,N_11791);
and U12171 (N_12171,N_11878,N_11226);
xnor U12172 (N_12172,N_11142,N_11318);
nor U12173 (N_12173,N_11675,N_11966);
and U12174 (N_12174,N_11341,N_11523);
xor U12175 (N_12175,N_11285,N_11440);
or U12176 (N_12176,N_11757,N_11643);
and U12177 (N_12177,N_11841,N_11368);
and U12178 (N_12178,N_11298,N_11117);
or U12179 (N_12179,N_11921,N_11961);
and U12180 (N_12180,N_11430,N_11319);
and U12181 (N_12181,N_11224,N_11190);
nand U12182 (N_12182,N_11870,N_11062);
or U12183 (N_12183,N_11545,N_11282);
or U12184 (N_12184,N_11900,N_11525);
nor U12185 (N_12185,N_11470,N_11952);
nand U12186 (N_12186,N_11804,N_11280);
nor U12187 (N_12187,N_11843,N_11604);
nand U12188 (N_12188,N_11005,N_11088);
and U12189 (N_12189,N_11755,N_11105);
nor U12190 (N_12190,N_11914,N_11608);
nor U12191 (N_12191,N_11057,N_11091);
nor U12192 (N_12192,N_11678,N_11495);
and U12193 (N_12193,N_11126,N_11831);
nor U12194 (N_12194,N_11731,N_11092);
xnor U12195 (N_12195,N_11512,N_11653);
nand U12196 (N_12196,N_11814,N_11575);
or U12197 (N_12197,N_11029,N_11480);
nor U12198 (N_12198,N_11584,N_11051);
nand U12199 (N_12199,N_11093,N_11263);
nand U12200 (N_12200,N_11720,N_11571);
nor U12201 (N_12201,N_11241,N_11486);
nor U12202 (N_12202,N_11438,N_11359);
or U12203 (N_12203,N_11786,N_11449);
and U12204 (N_12204,N_11034,N_11085);
xnor U12205 (N_12205,N_11893,N_11072);
nor U12206 (N_12206,N_11833,N_11301);
or U12207 (N_12207,N_11191,N_11995);
or U12208 (N_12208,N_11855,N_11892);
xor U12209 (N_12209,N_11497,N_11847);
nor U12210 (N_12210,N_11262,N_11427);
and U12211 (N_12211,N_11955,N_11193);
or U12212 (N_12212,N_11171,N_11198);
nor U12213 (N_12213,N_11458,N_11866);
or U12214 (N_12214,N_11213,N_11987);
or U12215 (N_12215,N_11597,N_11007);
or U12216 (N_12216,N_11932,N_11647);
xor U12217 (N_12217,N_11311,N_11291);
nand U12218 (N_12218,N_11762,N_11821);
nand U12219 (N_12219,N_11094,N_11944);
nand U12220 (N_12220,N_11068,N_11381);
xor U12221 (N_12221,N_11825,N_11172);
or U12222 (N_12222,N_11018,N_11526);
or U12223 (N_12223,N_11130,N_11924);
nand U12224 (N_12224,N_11922,N_11148);
or U12225 (N_12225,N_11869,N_11180);
and U12226 (N_12226,N_11824,N_11238);
nand U12227 (N_12227,N_11110,N_11031);
nor U12228 (N_12228,N_11694,N_11351);
xor U12229 (N_12229,N_11657,N_11563);
xor U12230 (N_12230,N_11055,N_11644);
nand U12231 (N_12231,N_11011,N_11243);
nor U12232 (N_12232,N_11748,N_11699);
or U12233 (N_12233,N_11100,N_11382);
or U12234 (N_12234,N_11729,N_11447);
or U12235 (N_12235,N_11806,N_11194);
nor U12236 (N_12236,N_11730,N_11505);
xor U12237 (N_12237,N_11038,N_11503);
nand U12238 (N_12238,N_11242,N_11297);
or U12239 (N_12239,N_11390,N_11045);
xor U12240 (N_12240,N_11904,N_11151);
xnor U12241 (N_12241,N_11173,N_11196);
or U12242 (N_12242,N_11220,N_11681);
nand U12243 (N_12243,N_11764,N_11779);
xor U12244 (N_12244,N_11129,N_11392);
or U12245 (N_12245,N_11576,N_11246);
xnor U12246 (N_12246,N_11041,N_11202);
xnor U12247 (N_12247,N_11152,N_11325);
and U12248 (N_12248,N_11474,N_11353);
nand U12249 (N_12249,N_11770,N_11937);
nand U12250 (N_12250,N_11417,N_11083);
or U12251 (N_12251,N_11939,N_11864);
and U12252 (N_12252,N_11114,N_11927);
nand U12253 (N_12253,N_11903,N_11154);
xor U12254 (N_12254,N_11760,N_11310);
nand U12255 (N_12255,N_11230,N_11614);
xnor U12256 (N_12256,N_11134,N_11206);
and U12257 (N_12257,N_11200,N_11168);
xor U12258 (N_12258,N_11454,N_11743);
and U12259 (N_12259,N_11991,N_11274);
nor U12260 (N_12260,N_11547,N_11816);
nand U12261 (N_12261,N_11934,N_11912);
nand U12262 (N_12262,N_11679,N_11949);
nand U12263 (N_12263,N_11609,N_11535);
xnor U12264 (N_12264,N_11009,N_11797);
and U12265 (N_12265,N_11594,N_11723);
and U12266 (N_12266,N_11433,N_11112);
or U12267 (N_12267,N_11231,N_11235);
nor U12268 (N_12268,N_11901,N_11324);
xnor U12269 (N_12269,N_11109,N_11008);
and U12270 (N_12270,N_11345,N_11278);
nand U12271 (N_12271,N_11715,N_11615);
xor U12272 (N_12272,N_11021,N_11252);
xnor U12273 (N_12273,N_11186,N_11822);
nand U12274 (N_12274,N_11606,N_11909);
and U12275 (N_12275,N_11006,N_11121);
xnor U12276 (N_12276,N_11669,N_11445);
nor U12277 (N_12277,N_11307,N_11910);
xor U12278 (N_12278,N_11457,N_11369);
and U12279 (N_12279,N_11695,N_11832);
nor U12280 (N_12280,N_11933,N_11063);
or U12281 (N_12281,N_11020,N_11750);
nand U12282 (N_12282,N_11920,N_11104);
nand U12283 (N_12283,N_11087,N_11118);
and U12284 (N_12284,N_11929,N_11977);
and U12285 (N_12285,N_11332,N_11639);
nor U12286 (N_12286,N_11388,N_11880);
xnor U12287 (N_12287,N_11591,N_11270);
and U12288 (N_12288,N_11326,N_11399);
xnor U12289 (N_12289,N_11569,N_11981);
nand U12290 (N_12290,N_11911,N_11605);
nand U12291 (N_12291,N_11153,N_11146);
and U12292 (N_12292,N_11327,N_11103);
nand U12293 (N_12293,N_11942,N_11176);
and U12294 (N_12294,N_11524,N_11567);
and U12295 (N_12295,N_11216,N_11708);
nor U12296 (N_12296,N_11602,N_11516);
or U12297 (N_12297,N_11667,N_11724);
nor U12298 (N_12298,N_11453,N_11328);
or U12299 (N_12299,N_11089,N_11039);
xor U12300 (N_12300,N_11140,N_11646);
or U12301 (N_12301,N_11670,N_11553);
xor U12302 (N_12302,N_11756,N_11899);
nor U12303 (N_12303,N_11620,N_11158);
xnor U12304 (N_12304,N_11300,N_11162);
nand U12305 (N_12305,N_11387,N_11095);
nand U12306 (N_12306,N_11531,N_11984);
nor U12307 (N_12307,N_11120,N_11817);
or U12308 (N_12308,N_11905,N_11745);
and U12309 (N_12309,N_11170,N_11618);
and U12310 (N_12310,N_11838,N_11555);
nand U12311 (N_12311,N_11339,N_11568);
nor U12312 (N_12312,N_11469,N_11663);
nand U12313 (N_12313,N_11214,N_11477);
xor U12314 (N_12314,N_11631,N_11541);
or U12315 (N_12315,N_11528,N_11337);
nand U12316 (N_12316,N_11543,N_11394);
xnor U12317 (N_12317,N_11064,N_11287);
or U12318 (N_12318,N_11894,N_11931);
or U12319 (N_12319,N_11259,N_11099);
or U12320 (N_12320,N_11967,N_11012);
nand U12321 (N_12321,N_11802,N_11215);
xor U12322 (N_12322,N_11462,N_11128);
nand U12323 (N_12323,N_11716,N_11733);
nand U12324 (N_12324,N_11334,N_11520);
nor U12325 (N_12325,N_11389,N_11634);
xor U12326 (N_12326,N_11446,N_11079);
and U12327 (N_12327,N_11839,N_11819);
nor U12328 (N_12328,N_11098,N_11277);
xor U12329 (N_12329,N_11860,N_11406);
xnor U12330 (N_12330,N_11035,N_11974);
and U12331 (N_12331,N_11941,N_11954);
nand U12332 (N_12332,N_11379,N_11840);
nand U12333 (N_12333,N_11101,N_11959);
or U12334 (N_12334,N_11800,N_11289);
nor U12335 (N_12335,N_11177,N_11611);
or U12336 (N_12336,N_11185,N_11247);
nand U12337 (N_12337,N_11316,N_11395);
xor U12338 (N_12338,N_11383,N_11589);
nor U12339 (N_12339,N_11070,N_11108);
xor U12340 (N_12340,N_11986,N_11992);
and U12341 (N_12341,N_11442,N_11947);
nand U12342 (N_12342,N_11461,N_11248);
xnor U12343 (N_12343,N_11572,N_11507);
and U12344 (N_12344,N_11164,N_11522);
or U12345 (N_12345,N_11580,N_11997);
and U12346 (N_12346,N_11519,N_11074);
nand U12347 (N_12347,N_11356,N_11508);
xor U12348 (N_12348,N_11460,N_11124);
xnor U12349 (N_12349,N_11763,N_11017);
xor U12350 (N_12350,N_11616,N_11884);
nand U12351 (N_12351,N_11636,N_11475);
nand U12352 (N_12352,N_11443,N_11767);
nor U12353 (N_12353,N_11776,N_11424);
xnor U12354 (N_12354,N_11132,N_11897);
xnor U12355 (N_12355,N_11851,N_11625);
nor U12356 (N_12356,N_11769,N_11680);
nand U12357 (N_12357,N_11166,N_11665);
nand U12358 (N_12358,N_11856,N_11204);
nand U12359 (N_12359,N_11378,N_11490);
nand U12360 (N_12360,N_11275,N_11071);
and U12361 (N_12361,N_11370,N_11013);
xnor U12362 (N_12362,N_11741,N_11881);
or U12363 (N_12363,N_11962,N_11131);
nand U12364 (N_12364,N_11272,N_11794);
or U12365 (N_12365,N_11273,N_11610);
nand U12366 (N_12366,N_11157,N_11727);
and U12367 (N_12367,N_11842,N_11019);
xnor U12368 (N_12368,N_11209,N_11228);
xnor U12369 (N_12369,N_11002,N_11603);
nor U12370 (N_12370,N_11895,N_11364);
and U12371 (N_12371,N_11143,N_11772);
or U12372 (N_12372,N_11400,N_11671);
nor U12373 (N_12373,N_11182,N_11867);
or U12374 (N_12374,N_11739,N_11024);
or U12375 (N_12375,N_11630,N_11761);
xnor U12376 (N_12376,N_11303,N_11428);
or U12377 (N_12377,N_11913,N_11423);
nor U12378 (N_12378,N_11321,N_11774);
or U12379 (N_12379,N_11489,N_11965);
and U12380 (N_12380,N_11692,N_11254);
nor U12381 (N_12381,N_11257,N_11187);
nand U12382 (N_12382,N_11998,N_11286);
and U12383 (N_12383,N_11217,N_11306);
and U12384 (N_12384,N_11053,N_11868);
or U12385 (N_12385,N_11201,N_11861);
and U12386 (N_12386,N_11887,N_11292);
or U12387 (N_12387,N_11323,N_11054);
and U12388 (N_12388,N_11968,N_11701);
nor U12389 (N_12389,N_11222,N_11036);
nand U12390 (N_12390,N_11058,N_11219);
nand U12391 (N_12391,N_11710,N_11435);
or U12392 (N_12392,N_11078,N_11916);
nor U12393 (N_12393,N_11978,N_11043);
nand U12394 (N_12394,N_11236,N_11752);
nand U12395 (N_12395,N_11882,N_11771);
nand U12396 (N_12396,N_11698,N_11871);
nand U12397 (N_12397,N_11875,N_11362);
or U12398 (N_12398,N_11016,N_11221);
and U12399 (N_12399,N_11950,N_11737);
nand U12400 (N_12400,N_11346,N_11059);
nand U12401 (N_12401,N_11299,N_11975);
xnor U12402 (N_12402,N_11846,N_11141);
nand U12403 (N_12403,N_11979,N_11066);
xnor U12404 (N_12404,N_11498,N_11810);
nor U12405 (N_12405,N_11613,N_11023);
nand U12406 (N_12406,N_11295,N_11075);
nand U12407 (N_12407,N_11807,N_11360);
nor U12408 (N_12408,N_11642,N_11178);
nand U12409 (N_12409,N_11518,N_11455);
nand U12410 (N_12410,N_11759,N_11014);
nor U12411 (N_12411,N_11590,N_11372);
or U12412 (N_12412,N_11958,N_11448);
xnor U12413 (N_12413,N_11416,N_11343);
and U12414 (N_12414,N_11441,N_11260);
and U12415 (N_12415,N_11244,N_11410);
and U12416 (N_12416,N_11374,N_11677);
and U12417 (N_12417,N_11787,N_11084);
nor U12418 (N_12418,N_11999,N_11288);
nand U12419 (N_12419,N_11322,N_11338);
or U12420 (N_12420,N_11373,N_11865);
nand U12421 (N_12421,N_11393,N_11996);
nor U12422 (N_12422,N_11538,N_11192);
and U12423 (N_12423,N_11690,N_11596);
and U12424 (N_12424,N_11559,N_11946);
or U12425 (N_12425,N_11073,N_11317);
nor U12426 (N_12426,N_11188,N_11795);
and U12427 (N_12427,N_11660,N_11784);
or U12428 (N_12428,N_11513,N_11511);
nand U12429 (N_12429,N_11629,N_11546);
xnor U12430 (N_12430,N_11960,N_11593);
nor U12431 (N_12431,N_11754,N_11789);
nor U12432 (N_12432,N_11123,N_11566);
xor U12433 (N_12433,N_11684,N_11305);
xnor U12434 (N_12434,N_11633,N_11500);
xor U12435 (N_12435,N_11135,N_11585);
and U12436 (N_12436,N_11472,N_11565);
nand U12437 (N_12437,N_11859,N_11815);
nand U12438 (N_12438,N_11402,N_11872);
and U12439 (N_12439,N_11386,N_11065);
nand U12440 (N_12440,N_11654,N_11391);
or U12441 (N_12441,N_11234,N_11581);
and U12442 (N_12442,N_11456,N_11719);
and U12443 (N_12443,N_11409,N_11775);
nor U12444 (N_12444,N_11342,N_11293);
xor U12445 (N_12445,N_11161,N_11536);
or U12446 (N_12446,N_11468,N_11925);
xnor U12447 (N_12447,N_11115,N_11704);
or U12448 (N_12448,N_11466,N_11147);
or U12449 (N_12449,N_11205,N_11696);
and U12450 (N_12450,N_11627,N_11047);
nor U12451 (N_12451,N_11481,N_11363);
nor U12452 (N_12452,N_11211,N_11371);
nand U12453 (N_12453,N_11969,N_11907);
xnor U12454 (N_12454,N_11539,N_11050);
nand U12455 (N_12455,N_11155,N_11888);
and U12456 (N_12456,N_11439,N_11908);
nor U12457 (N_12457,N_11414,N_11577);
nand U12458 (N_12458,N_11711,N_11403);
or U12459 (N_12459,N_11267,N_11396);
nand U12460 (N_12460,N_11281,N_11879);
nor U12461 (N_12461,N_11350,N_11137);
and U12462 (N_12462,N_11583,N_11476);
and U12463 (N_12463,N_11906,N_11313);
or U12464 (N_12464,N_11471,N_11697);
and U12465 (N_12465,N_11001,N_11212);
and U12466 (N_12466,N_11873,N_11349);
and U12467 (N_12467,N_11587,N_11174);
nor U12468 (N_12468,N_11820,N_11375);
xor U12469 (N_12469,N_11935,N_11714);
or U12470 (N_12470,N_11768,N_11706);
and U12471 (N_12471,N_11874,N_11245);
xnor U12472 (N_12472,N_11463,N_11163);
or U12473 (N_12473,N_11352,N_11022);
nor U12474 (N_12474,N_11668,N_11835);
xor U12475 (N_12475,N_11554,N_11450);
or U12476 (N_12476,N_11973,N_11766);
or U12477 (N_12477,N_11354,N_11269);
nand U12478 (N_12478,N_11885,N_11033);
xor U12479 (N_12479,N_11127,N_11496);
xor U12480 (N_12480,N_11862,N_11258);
nand U12481 (N_12481,N_11333,N_11376);
xnor U12482 (N_12482,N_11276,N_11256);
nand U12483 (N_12483,N_11530,N_11465);
nand U12484 (N_12484,N_11622,N_11830);
xnor U12485 (N_12485,N_11534,N_11658);
and U12486 (N_12486,N_11253,N_11107);
nor U12487 (N_12487,N_11090,N_11502);
xnor U12488 (N_12488,N_11540,N_11208);
and U12489 (N_12489,N_11464,N_11890);
xor U12490 (N_12490,N_11052,N_11564);
nor U12491 (N_12491,N_11549,N_11793);
nand U12492 (N_12492,N_11296,N_11261);
nand U12493 (N_12493,N_11096,N_11758);
xnor U12494 (N_12494,N_11160,N_11077);
xor U12495 (N_12495,N_11264,N_11426);
or U12496 (N_12496,N_11923,N_11707);
nand U12497 (N_12497,N_11125,N_11266);
nand U12498 (N_12498,N_11479,N_11509);
nand U12499 (N_12499,N_11493,N_11483);
xor U12500 (N_12500,N_11012,N_11912);
nand U12501 (N_12501,N_11751,N_11871);
and U12502 (N_12502,N_11127,N_11380);
or U12503 (N_12503,N_11481,N_11517);
nand U12504 (N_12504,N_11291,N_11061);
nand U12505 (N_12505,N_11107,N_11815);
nand U12506 (N_12506,N_11218,N_11931);
xnor U12507 (N_12507,N_11386,N_11971);
nand U12508 (N_12508,N_11975,N_11719);
nand U12509 (N_12509,N_11007,N_11773);
nand U12510 (N_12510,N_11133,N_11029);
and U12511 (N_12511,N_11518,N_11916);
nand U12512 (N_12512,N_11799,N_11125);
and U12513 (N_12513,N_11731,N_11201);
nand U12514 (N_12514,N_11073,N_11153);
nand U12515 (N_12515,N_11934,N_11304);
xor U12516 (N_12516,N_11307,N_11259);
nor U12517 (N_12517,N_11537,N_11173);
and U12518 (N_12518,N_11825,N_11053);
or U12519 (N_12519,N_11514,N_11806);
nor U12520 (N_12520,N_11993,N_11289);
xnor U12521 (N_12521,N_11783,N_11026);
xnor U12522 (N_12522,N_11955,N_11040);
nor U12523 (N_12523,N_11948,N_11038);
or U12524 (N_12524,N_11385,N_11499);
nand U12525 (N_12525,N_11422,N_11051);
nand U12526 (N_12526,N_11274,N_11807);
xor U12527 (N_12527,N_11935,N_11908);
xnor U12528 (N_12528,N_11162,N_11239);
nor U12529 (N_12529,N_11062,N_11842);
xor U12530 (N_12530,N_11343,N_11387);
or U12531 (N_12531,N_11663,N_11225);
and U12532 (N_12532,N_11413,N_11141);
nor U12533 (N_12533,N_11672,N_11882);
nand U12534 (N_12534,N_11726,N_11937);
nand U12535 (N_12535,N_11905,N_11588);
xor U12536 (N_12536,N_11129,N_11875);
or U12537 (N_12537,N_11108,N_11297);
or U12538 (N_12538,N_11346,N_11336);
nor U12539 (N_12539,N_11636,N_11444);
or U12540 (N_12540,N_11525,N_11375);
xor U12541 (N_12541,N_11774,N_11732);
nand U12542 (N_12542,N_11671,N_11814);
nand U12543 (N_12543,N_11680,N_11426);
nand U12544 (N_12544,N_11850,N_11718);
or U12545 (N_12545,N_11982,N_11060);
and U12546 (N_12546,N_11091,N_11935);
nor U12547 (N_12547,N_11938,N_11669);
or U12548 (N_12548,N_11049,N_11274);
nand U12549 (N_12549,N_11291,N_11954);
and U12550 (N_12550,N_11271,N_11890);
nand U12551 (N_12551,N_11732,N_11897);
nor U12552 (N_12552,N_11097,N_11507);
nor U12553 (N_12553,N_11077,N_11414);
and U12554 (N_12554,N_11421,N_11546);
xor U12555 (N_12555,N_11243,N_11239);
xor U12556 (N_12556,N_11546,N_11219);
or U12557 (N_12557,N_11443,N_11226);
xor U12558 (N_12558,N_11611,N_11805);
and U12559 (N_12559,N_11842,N_11190);
nand U12560 (N_12560,N_11620,N_11509);
nand U12561 (N_12561,N_11851,N_11972);
xor U12562 (N_12562,N_11334,N_11174);
and U12563 (N_12563,N_11777,N_11036);
or U12564 (N_12564,N_11808,N_11894);
or U12565 (N_12565,N_11236,N_11198);
xnor U12566 (N_12566,N_11814,N_11263);
xor U12567 (N_12567,N_11136,N_11493);
or U12568 (N_12568,N_11830,N_11282);
and U12569 (N_12569,N_11186,N_11927);
nor U12570 (N_12570,N_11005,N_11327);
or U12571 (N_12571,N_11281,N_11006);
and U12572 (N_12572,N_11418,N_11650);
nand U12573 (N_12573,N_11925,N_11495);
nor U12574 (N_12574,N_11366,N_11036);
and U12575 (N_12575,N_11922,N_11056);
xor U12576 (N_12576,N_11758,N_11064);
and U12577 (N_12577,N_11627,N_11197);
nor U12578 (N_12578,N_11810,N_11942);
nor U12579 (N_12579,N_11294,N_11554);
nand U12580 (N_12580,N_11565,N_11390);
and U12581 (N_12581,N_11611,N_11637);
xor U12582 (N_12582,N_11529,N_11481);
and U12583 (N_12583,N_11175,N_11895);
and U12584 (N_12584,N_11808,N_11381);
and U12585 (N_12585,N_11101,N_11972);
nor U12586 (N_12586,N_11305,N_11301);
nor U12587 (N_12587,N_11630,N_11620);
xor U12588 (N_12588,N_11546,N_11661);
nor U12589 (N_12589,N_11360,N_11236);
xnor U12590 (N_12590,N_11950,N_11217);
xor U12591 (N_12591,N_11382,N_11839);
nor U12592 (N_12592,N_11103,N_11938);
nand U12593 (N_12593,N_11135,N_11485);
or U12594 (N_12594,N_11311,N_11983);
and U12595 (N_12595,N_11329,N_11246);
or U12596 (N_12596,N_11886,N_11283);
nand U12597 (N_12597,N_11162,N_11513);
nand U12598 (N_12598,N_11346,N_11446);
nand U12599 (N_12599,N_11152,N_11052);
nand U12600 (N_12600,N_11306,N_11173);
or U12601 (N_12601,N_11769,N_11564);
xor U12602 (N_12602,N_11222,N_11132);
or U12603 (N_12603,N_11884,N_11613);
or U12604 (N_12604,N_11369,N_11249);
nor U12605 (N_12605,N_11429,N_11127);
nand U12606 (N_12606,N_11606,N_11945);
and U12607 (N_12607,N_11766,N_11085);
and U12608 (N_12608,N_11866,N_11742);
and U12609 (N_12609,N_11901,N_11382);
nand U12610 (N_12610,N_11076,N_11750);
xnor U12611 (N_12611,N_11120,N_11702);
or U12612 (N_12612,N_11898,N_11421);
nand U12613 (N_12613,N_11502,N_11683);
nor U12614 (N_12614,N_11608,N_11715);
nand U12615 (N_12615,N_11339,N_11509);
or U12616 (N_12616,N_11689,N_11441);
nand U12617 (N_12617,N_11292,N_11152);
or U12618 (N_12618,N_11299,N_11443);
nand U12619 (N_12619,N_11964,N_11954);
nor U12620 (N_12620,N_11411,N_11027);
and U12621 (N_12621,N_11139,N_11308);
or U12622 (N_12622,N_11354,N_11202);
and U12623 (N_12623,N_11094,N_11469);
or U12624 (N_12624,N_11213,N_11767);
nor U12625 (N_12625,N_11670,N_11949);
xor U12626 (N_12626,N_11134,N_11244);
or U12627 (N_12627,N_11327,N_11932);
and U12628 (N_12628,N_11190,N_11408);
xor U12629 (N_12629,N_11196,N_11953);
xor U12630 (N_12630,N_11347,N_11712);
nand U12631 (N_12631,N_11669,N_11726);
or U12632 (N_12632,N_11347,N_11817);
or U12633 (N_12633,N_11038,N_11341);
and U12634 (N_12634,N_11541,N_11254);
and U12635 (N_12635,N_11764,N_11737);
nand U12636 (N_12636,N_11971,N_11007);
nand U12637 (N_12637,N_11057,N_11151);
nand U12638 (N_12638,N_11748,N_11666);
nand U12639 (N_12639,N_11017,N_11533);
nand U12640 (N_12640,N_11581,N_11384);
xor U12641 (N_12641,N_11015,N_11445);
or U12642 (N_12642,N_11690,N_11663);
and U12643 (N_12643,N_11075,N_11959);
xor U12644 (N_12644,N_11039,N_11980);
or U12645 (N_12645,N_11671,N_11802);
or U12646 (N_12646,N_11166,N_11183);
or U12647 (N_12647,N_11490,N_11400);
and U12648 (N_12648,N_11834,N_11998);
xnor U12649 (N_12649,N_11719,N_11098);
xnor U12650 (N_12650,N_11969,N_11626);
or U12651 (N_12651,N_11840,N_11151);
and U12652 (N_12652,N_11422,N_11484);
and U12653 (N_12653,N_11695,N_11748);
or U12654 (N_12654,N_11105,N_11290);
xor U12655 (N_12655,N_11208,N_11443);
nor U12656 (N_12656,N_11674,N_11499);
xor U12657 (N_12657,N_11052,N_11395);
and U12658 (N_12658,N_11039,N_11637);
xnor U12659 (N_12659,N_11977,N_11914);
nand U12660 (N_12660,N_11523,N_11463);
xnor U12661 (N_12661,N_11882,N_11581);
nor U12662 (N_12662,N_11655,N_11183);
nand U12663 (N_12663,N_11030,N_11853);
and U12664 (N_12664,N_11328,N_11483);
or U12665 (N_12665,N_11632,N_11628);
nor U12666 (N_12666,N_11131,N_11237);
xor U12667 (N_12667,N_11913,N_11907);
nor U12668 (N_12668,N_11464,N_11646);
nor U12669 (N_12669,N_11044,N_11063);
and U12670 (N_12670,N_11895,N_11225);
xor U12671 (N_12671,N_11271,N_11660);
or U12672 (N_12672,N_11092,N_11948);
nand U12673 (N_12673,N_11207,N_11355);
nand U12674 (N_12674,N_11979,N_11718);
and U12675 (N_12675,N_11688,N_11133);
nor U12676 (N_12676,N_11519,N_11207);
or U12677 (N_12677,N_11210,N_11144);
nand U12678 (N_12678,N_11226,N_11880);
xnor U12679 (N_12679,N_11561,N_11070);
and U12680 (N_12680,N_11739,N_11302);
or U12681 (N_12681,N_11069,N_11254);
nand U12682 (N_12682,N_11083,N_11656);
and U12683 (N_12683,N_11551,N_11909);
xnor U12684 (N_12684,N_11382,N_11837);
and U12685 (N_12685,N_11516,N_11246);
xor U12686 (N_12686,N_11301,N_11053);
and U12687 (N_12687,N_11776,N_11113);
and U12688 (N_12688,N_11320,N_11957);
xor U12689 (N_12689,N_11079,N_11697);
nand U12690 (N_12690,N_11275,N_11355);
xnor U12691 (N_12691,N_11051,N_11303);
nand U12692 (N_12692,N_11269,N_11587);
and U12693 (N_12693,N_11644,N_11343);
nand U12694 (N_12694,N_11748,N_11893);
nand U12695 (N_12695,N_11821,N_11380);
nor U12696 (N_12696,N_11380,N_11537);
and U12697 (N_12697,N_11504,N_11716);
xnor U12698 (N_12698,N_11468,N_11873);
and U12699 (N_12699,N_11125,N_11942);
or U12700 (N_12700,N_11007,N_11290);
xnor U12701 (N_12701,N_11173,N_11770);
and U12702 (N_12702,N_11902,N_11176);
nor U12703 (N_12703,N_11018,N_11282);
or U12704 (N_12704,N_11904,N_11126);
or U12705 (N_12705,N_11751,N_11343);
nor U12706 (N_12706,N_11671,N_11153);
or U12707 (N_12707,N_11157,N_11857);
and U12708 (N_12708,N_11132,N_11490);
nand U12709 (N_12709,N_11906,N_11094);
or U12710 (N_12710,N_11667,N_11375);
nand U12711 (N_12711,N_11384,N_11881);
nand U12712 (N_12712,N_11337,N_11138);
or U12713 (N_12713,N_11327,N_11930);
xnor U12714 (N_12714,N_11280,N_11606);
or U12715 (N_12715,N_11964,N_11802);
or U12716 (N_12716,N_11651,N_11381);
nand U12717 (N_12717,N_11119,N_11196);
nor U12718 (N_12718,N_11029,N_11831);
or U12719 (N_12719,N_11229,N_11077);
nor U12720 (N_12720,N_11487,N_11896);
or U12721 (N_12721,N_11138,N_11503);
and U12722 (N_12722,N_11700,N_11755);
and U12723 (N_12723,N_11192,N_11616);
xnor U12724 (N_12724,N_11688,N_11197);
xnor U12725 (N_12725,N_11874,N_11622);
or U12726 (N_12726,N_11531,N_11566);
or U12727 (N_12727,N_11800,N_11188);
nor U12728 (N_12728,N_11896,N_11679);
or U12729 (N_12729,N_11484,N_11054);
or U12730 (N_12730,N_11131,N_11568);
nor U12731 (N_12731,N_11718,N_11486);
or U12732 (N_12732,N_11836,N_11702);
and U12733 (N_12733,N_11034,N_11599);
and U12734 (N_12734,N_11698,N_11923);
nand U12735 (N_12735,N_11074,N_11048);
nor U12736 (N_12736,N_11853,N_11779);
xnor U12737 (N_12737,N_11123,N_11306);
nor U12738 (N_12738,N_11278,N_11521);
or U12739 (N_12739,N_11583,N_11985);
or U12740 (N_12740,N_11934,N_11377);
nor U12741 (N_12741,N_11862,N_11484);
nor U12742 (N_12742,N_11656,N_11983);
nor U12743 (N_12743,N_11574,N_11650);
xnor U12744 (N_12744,N_11571,N_11813);
or U12745 (N_12745,N_11517,N_11496);
and U12746 (N_12746,N_11329,N_11416);
xor U12747 (N_12747,N_11719,N_11482);
nor U12748 (N_12748,N_11396,N_11903);
nor U12749 (N_12749,N_11047,N_11564);
nor U12750 (N_12750,N_11426,N_11131);
or U12751 (N_12751,N_11585,N_11321);
nand U12752 (N_12752,N_11780,N_11333);
xor U12753 (N_12753,N_11954,N_11419);
and U12754 (N_12754,N_11024,N_11795);
nand U12755 (N_12755,N_11914,N_11582);
xor U12756 (N_12756,N_11390,N_11457);
nor U12757 (N_12757,N_11709,N_11843);
nand U12758 (N_12758,N_11439,N_11467);
and U12759 (N_12759,N_11548,N_11311);
and U12760 (N_12760,N_11423,N_11341);
xnor U12761 (N_12761,N_11514,N_11379);
nand U12762 (N_12762,N_11340,N_11608);
xor U12763 (N_12763,N_11959,N_11932);
and U12764 (N_12764,N_11913,N_11335);
or U12765 (N_12765,N_11064,N_11668);
and U12766 (N_12766,N_11644,N_11483);
nor U12767 (N_12767,N_11905,N_11790);
or U12768 (N_12768,N_11335,N_11082);
or U12769 (N_12769,N_11053,N_11607);
or U12770 (N_12770,N_11035,N_11595);
and U12771 (N_12771,N_11654,N_11327);
and U12772 (N_12772,N_11467,N_11860);
nand U12773 (N_12773,N_11097,N_11136);
nor U12774 (N_12774,N_11970,N_11800);
and U12775 (N_12775,N_11665,N_11802);
xor U12776 (N_12776,N_11584,N_11139);
nor U12777 (N_12777,N_11161,N_11810);
nand U12778 (N_12778,N_11499,N_11260);
or U12779 (N_12779,N_11926,N_11582);
nand U12780 (N_12780,N_11711,N_11913);
or U12781 (N_12781,N_11998,N_11291);
xor U12782 (N_12782,N_11383,N_11988);
or U12783 (N_12783,N_11185,N_11517);
nand U12784 (N_12784,N_11423,N_11184);
or U12785 (N_12785,N_11037,N_11146);
or U12786 (N_12786,N_11211,N_11433);
or U12787 (N_12787,N_11745,N_11512);
or U12788 (N_12788,N_11057,N_11260);
nand U12789 (N_12789,N_11706,N_11666);
nor U12790 (N_12790,N_11150,N_11587);
nor U12791 (N_12791,N_11022,N_11063);
or U12792 (N_12792,N_11739,N_11725);
nand U12793 (N_12793,N_11654,N_11918);
nor U12794 (N_12794,N_11954,N_11044);
and U12795 (N_12795,N_11994,N_11693);
and U12796 (N_12796,N_11121,N_11303);
or U12797 (N_12797,N_11865,N_11976);
xnor U12798 (N_12798,N_11673,N_11415);
xor U12799 (N_12799,N_11078,N_11069);
nor U12800 (N_12800,N_11249,N_11374);
nor U12801 (N_12801,N_11049,N_11023);
or U12802 (N_12802,N_11736,N_11001);
nor U12803 (N_12803,N_11936,N_11589);
xor U12804 (N_12804,N_11679,N_11668);
nor U12805 (N_12805,N_11234,N_11149);
and U12806 (N_12806,N_11184,N_11900);
nand U12807 (N_12807,N_11381,N_11767);
nand U12808 (N_12808,N_11621,N_11961);
xor U12809 (N_12809,N_11098,N_11996);
xor U12810 (N_12810,N_11326,N_11807);
and U12811 (N_12811,N_11235,N_11441);
or U12812 (N_12812,N_11516,N_11009);
nor U12813 (N_12813,N_11172,N_11186);
or U12814 (N_12814,N_11821,N_11869);
nand U12815 (N_12815,N_11041,N_11416);
and U12816 (N_12816,N_11576,N_11683);
nand U12817 (N_12817,N_11305,N_11972);
and U12818 (N_12818,N_11416,N_11726);
and U12819 (N_12819,N_11619,N_11705);
nand U12820 (N_12820,N_11525,N_11557);
or U12821 (N_12821,N_11244,N_11369);
and U12822 (N_12822,N_11689,N_11911);
xor U12823 (N_12823,N_11399,N_11584);
nand U12824 (N_12824,N_11308,N_11255);
nor U12825 (N_12825,N_11585,N_11594);
or U12826 (N_12826,N_11201,N_11598);
nor U12827 (N_12827,N_11141,N_11584);
and U12828 (N_12828,N_11068,N_11842);
nor U12829 (N_12829,N_11398,N_11332);
xnor U12830 (N_12830,N_11027,N_11867);
nor U12831 (N_12831,N_11125,N_11788);
nand U12832 (N_12832,N_11922,N_11379);
or U12833 (N_12833,N_11664,N_11680);
nor U12834 (N_12834,N_11312,N_11648);
and U12835 (N_12835,N_11473,N_11249);
nand U12836 (N_12836,N_11571,N_11497);
or U12837 (N_12837,N_11994,N_11533);
nor U12838 (N_12838,N_11293,N_11391);
or U12839 (N_12839,N_11300,N_11378);
or U12840 (N_12840,N_11639,N_11007);
or U12841 (N_12841,N_11683,N_11272);
or U12842 (N_12842,N_11494,N_11839);
and U12843 (N_12843,N_11442,N_11172);
or U12844 (N_12844,N_11068,N_11582);
nor U12845 (N_12845,N_11188,N_11709);
xor U12846 (N_12846,N_11024,N_11282);
or U12847 (N_12847,N_11681,N_11711);
nand U12848 (N_12848,N_11535,N_11990);
xor U12849 (N_12849,N_11088,N_11027);
or U12850 (N_12850,N_11972,N_11942);
nor U12851 (N_12851,N_11435,N_11752);
nand U12852 (N_12852,N_11341,N_11813);
or U12853 (N_12853,N_11123,N_11708);
and U12854 (N_12854,N_11265,N_11799);
xor U12855 (N_12855,N_11548,N_11821);
and U12856 (N_12856,N_11403,N_11280);
and U12857 (N_12857,N_11623,N_11025);
nand U12858 (N_12858,N_11816,N_11118);
nand U12859 (N_12859,N_11563,N_11431);
and U12860 (N_12860,N_11568,N_11836);
or U12861 (N_12861,N_11523,N_11546);
nor U12862 (N_12862,N_11896,N_11138);
xor U12863 (N_12863,N_11073,N_11371);
nor U12864 (N_12864,N_11345,N_11220);
or U12865 (N_12865,N_11015,N_11497);
nand U12866 (N_12866,N_11366,N_11772);
or U12867 (N_12867,N_11973,N_11462);
or U12868 (N_12868,N_11329,N_11612);
nor U12869 (N_12869,N_11482,N_11946);
xor U12870 (N_12870,N_11737,N_11120);
nand U12871 (N_12871,N_11038,N_11188);
nand U12872 (N_12872,N_11095,N_11241);
and U12873 (N_12873,N_11282,N_11230);
or U12874 (N_12874,N_11837,N_11559);
nand U12875 (N_12875,N_11731,N_11788);
nor U12876 (N_12876,N_11444,N_11470);
and U12877 (N_12877,N_11596,N_11939);
nor U12878 (N_12878,N_11139,N_11543);
nor U12879 (N_12879,N_11200,N_11383);
nand U12880 (N_12880,N_11269,N_11301);
and U12881 (N_12881,N_11525,N_11418);
xnor U12882 (N_12882,N_11686,N_11989);
nor U12883 (N_12883,N_11203,N_11959);
and U12884 (N_12884,N_11576,N_11276);
and U12885 (N_12885,N_11837,N_11486);
xnor U12886 (N_12886,N_11823,N_11656);
xnor U12887 (N_12887,N_11257,N_11218);
and U12888 (N_12888,N_11159,N_11167);
or U12889 (N_12889,N_11995,N_11597);
nand U12890 (N_12890,N_11710,N_11281);
or U12891 (N_12891,N_11938,N_11685);
xor U12892 (N_12892,N_11079,N_11771);
or U12893 (N_12893,N_11075,N_11586);
xnor U12894 (N_12894,N_11687,N_11299);
nand U12895 (N_12895,N_11464,N_11521);
nand U12896 (N_12896,N_11802,N_11391);
nand U12897 (N_12897,N_11880,N_11354);
xnor U12898 (N_12898,N_11256,N_11617);
nor U12899 (N_12899,N_11132,N_11740);
and U12900 (N_12900,N_11353,N_11379);
and U12901 (N_12901,N_11292,N_11785);
nand U12902 (N_12902,N_11607,N_11102);
nor U12903 (N_12903,N_11991,N_11529);
xnor U12904 (N_12904,N_11773,N_11818);
xnor U12905 (N_12905,N_11088,N_11266);
or U12906 (N_12906,N_11055,N_11196);
nor U12907 (N_12907,N_11113,N_11076);
and U12908 (N_12908,N_11425,N_11194);
nor U12909 (N_12909,N_11684,N_11099);
and U12910 (N_12910,N_11785,N_11278);
or U12911 (N_12911,N_11337,N_11583);
or U12912 (N_12912,N_11146,N_11750);
and U12913 (N_12913,N_11117,N_11360);
and U12914 (N_12914,N_11701,N_11007);
nand U12915 (N_12915,N_11646,N_11090);
or U12916 (N_12916,N_11651,N_11582);
and U12917 (N_12917,N_11218,N_11752);
xnor U12918 (N_12918,N_11918,N_11915);
and U12919 (N_12919,N_11482,N_11136);
and U12920 (N_12920,N_11417,N_11099);
nor U12921 (N_12921,N_11395,N_11824);
xor U12922 (N_12922,N_11790,N_11113);
or U12923 (N_12923,N_11444,N_11985);
nand U12924 (N_12924,N_11371,N_11659);
nand U12925 (N_12925,N_11890,N_11266);
nand U12926 (N_12926,N_11994,N_11666);
nand U12927 (N_12927,N_11922,N_11453);
xor U12928 (N_12928,N_11968,N_11141);
xor U12929 (N_12929,N_11050,N_11046);
or U12930 (N_12930,N_11474,N_11665);
xor U12931 (N_12931,N_11117,N_11207);
and U12932 (N_12932,N_11557,N_11043);
xnor U12933 (N_12933,N_11851,N_11047);
and U12934 (N_12934,N_11976,N_11860);
nand U12935 (N_12935,N_11579,N_11234);
or U12936 (N_12936,N_11404,N_11588);
and U12937 (N_12937,N_11395,N_11794);
xnor U12938 (N_12938,N_11503,N_11127);
and U12939 (N_12939,N_11385,N_11893);
nor U12940 (N_12940,N_11407,N_11471);
or U12941 (N_12941,N_11270,N_11149);
xnor U12942 (N_12942,N_11882,N_11529);
nand U12943 (N_12943,N_11309,N_11915);
or U12944 (N_12944,N_11373,N_11174);
xnor U12945 (N_12945,N_11338,N_11610);
nor U12946 (N_12946,N_11419,N_11050);
xnor U12947 (N_12947,N_11560,N_11413);
nor U12948 (N_12948,N_11226,N_11196);
or U12949 (N_12949,N_11944,N_11783);
or U12950 (N_12950,N_11751,N_11794);
or U12951 (N_12951,N_11079,N_11919);
nand U12952 (N_12952,N_11737,N_11828);
or U12953 (N_12953,N_11853,N_11244);
nor U12954 (N_12954,N_11648,N_11129);
nor U12955 (N_12955,N_11729,N_11521);
xor U12956 (N_12956,N_11126,N_11284);
or U12957 (N_12957,N_11737,N_11309);
xor U12958 (N_12958,N_11116,N_11439);
xor U12959 (N_12959,N_11482,N_11683);
xnor U12960 (N_12960,N_11868,N_11065);
or U12961 (N_12961,N_11715,N_11524);
nand U12962 (N_12962,N_11562,N_11334);
nand U12963 (N_12963,N_11513,N_11526);
or U12964 (N_12964,N_11512,N_11451);
nand U12965 (N_12965,N_11767,N_11874);
nor U12966 (N_12966,N_11996,N_11717);
nand U12967 (N_12967,N_11207,N_11627);
nor U12968 (N_12968,N_11790,N_11336);
and U12969 (N_12969,N_11787,N_11917);
xnor U12970 (N_12970,N_11021,N_11555);
xor U12971 (N_12971,N_11596,N_11069);
or U12972 (N_12972,N_11638,N_11704);
nand U12973 (N_12973,N_11227,N_11846);
nand U12974 (N_12974,N_11692,N_11546);
nand U12975 (N_12975,N_11939,N_11763);
nor U12976 (N_12976,N_11547,N_11492);
nand U12977 (N_12977,N_11443,N_11651);
nand U12978 (N_12978,N_11769,N_11159);
or U12979 (N_12979,N_11563,N_11084);
or U12980 (N_12980,N_11617,N_11641);
nor U12981 (N_12981,N_11889,N_11060);
and U12982 (N_12982,N_11489,N_11612);
xor U12983 (N_12983,N_11850,N_11383);
xor U12984 (N_12984,N_11723,N_11767);
nand U12985 (N_12985,N_11826,N_11289);
nor U12986 (N_12986,N_11597,N_11641);
xnor U12987 (N_12987,N_11597,N_11414);
nand U12988 (N_12988,N_11737,N_11702);
or U12989 (N_12989,N_11405,N_11360);
xor U12990 (N_12990,N_11180,N_11265);
xnor U12991 (N_12991,N_11208,N_11422);
and U12992 (N_12992,N_11447,N_11503);
nor U12993 (N_12993,N_11318,N_11442);
or U12994 (N_12994,N_11196,N_11812);
and U12995 (N_12995,N_11580,N_11519);
or U12996 (N_12996,N_11185,N_11096);
and U12997 (N_12997,N_11134,N_11998);
and U12998 (N_12998,N_11565,N_11623);
nor U12999 (N_12999,N_11651,N_11791);
nor U13000 (N_13000,N_12763,N_12971);
nand U13001 (N_13001,N_12806,N_12455);
xnor U13002 (N_13002,N_12324,N_12101);
and U13003 (N_13003,N_12362,N_12798);
xnor U13004 (N_13004,N_12283,N_12855);
and U13005 (N_13005,N_12964,N_12249);
nand U13006 (N_13006,N_12134,N_12412);
or U13007 (N_13007,N_12478,N_12114);
xor U13008 (N_13008,N_12409,N_12642);
nor U13009 (N_13009,N_12269,N_12557);
nor U13010 (N_13010,N_12127,N_12054);
xnor U13011 (N_13011,N_12172,N_12709);
or U13012 (N_13012,N_12427,N_12107);
or U13013 (N_13013,N_12947,N_12193);
nand U13014 (N_13014,N_12475,N_12446);
and U13015 (N_13015,N_12527,N_12816);
and U13016 (N_13016,N_12915,N_12242);
nand U13017 (N_13017,N_12080,N_12065);
xnor U13018 (N_13018,N_12335,N_12442);
nor U13019 (N_13019,N_12733,N_12079);
xnor U13020 (N_13020,N_12483,N_12801);
and U13021 (N_13021,N_12099,N_12364);
nor U13022 (N_13022,N_12055,N_12960);
nand U13023 (N_13023,N_12706,N_12875);
or U13024 (N_13024,N_12687,N_12419);
and U13025 (N_13025,N_12753,N_12067);
and U13026 (N_13026,N_12985,N_12363);
nor U13027 (N_13027,N_12370,N_12568);
xor U13028 (N_13028,N_12423,N_12639);
nor U13029 (N_13029,N_12145,N_12760);
or U13030 (N_13030,N_12720,N_12053);
nor U13031 (N_13031,N_12002,N_12360);
and U13032 (N_13032,N_12481,N_12043);
nor U13033 (N_13033,N_12644,N_12774);
nand U13034 (N_13034,N_12573,N_12980);
nor U13035 (N_13035,N_12815,N_12896);
nand U13036 (N_13036,N_12197,N_12665);
xnor U13037 (N_13037,N_12930,N_12317);
xnor U13038 (N_13038,N_12461,N_12117);
or U13039 (N_13039,N_12656,N_12630);
nand U13040 (N_13040,N_12589,N_12584);
nor U13041 (N_13041,N_12281,N_12789);
nand U13042 (N_13042,N_12693,N_12883);
or U13043 (N_13043,N_12426,N_12983);
nor U13044 (N_13044,N_12682,N_12035);
nand U13045 (N_13045,N_12070,N_12711);
xor U13046 (N_13046,N_12950,N_12521);
nor U13047 (N_13047,N_12981,N_12278);
and U13048 (N_13048,N_12390,N_12371);
nor U13049 (N_13049,N_12128,N_12498);
xnor U13050 (N_13050,N_12480,N_12357);
and U13051 (N_13051,N_12177,N_12492);
or U13052 (N_13052,N_12803,N_12617);
or U13053 (N_13053,N_12543,N_12171);
nor U13054 (N_13054,N_12619,N_12895);
xor U13055 (N_13055,N_12474,N_12424);
nand U13056 (N_13056,N_12247,N_12635);
and U13057 (N_13057,N_12230,N_12661);
and U13058 (N_13058,N_12306,N_12150);
and U13059 (N_13059,N_12032,N_12702);
nand U13060 (N_13060,N_12751,N_12392);
or U13061 (N_13061,N_12927,N_12141);
nand U13062 (N_13062,N_12995,N_12185);
xnor U13063 (N_13063,N_12484,N_12976);
xnor U13064 (N_13064,N_12119,N_12092);
nor U13065 (N_13065,N_12776,N_12533);
nand U13066 (N_13066,N_12777,N_12962);
and U13067 (N_13067,N_12076,N_12752);
or U13068 (N_13068,N_12041,N_12365);
or U13069 (N_13069,N_12603,N_12289);
or U13070 (N_13070,N_12571,N_12633);
or U13071 (N_13071,N_12257,N_12137);
nor U13072 (N_13072,N_12063,N_12116);
xnor U13073 (N_13073,N_12519,N_12946);
nor U13074 (N_13074,N_12270,N_12914);
xnor U13075 (N_13075,N_12704,N_12576);
nor U13076 (N_13076,N_12579,N_12515);
nand U13077 (N_13077,N_12337,N_12773);
and U13078 (N_13078,N_12325,N_12315);
nand U13079 (N_13079,N_12613,N_12098);
nand U13080 (N_13080,N_12303,N_12192);
nor U13081 (N_13081,N_12266,N_12856);
nand U13082 (N_13082,N_12183,N_12597);
nor U13083 (N_13083,N_12651,N_12731);
xnor U13084 (N_13084,N_12404,N_12788);
or U13085 (N_13085,N_12186,N_12354);
xor U13086 (N_13086,N_12330,N_12332);
nor U13087 (N_13087,N_12061,N_12372);
xnor U13088 (N_13088,N_12085,N_12545);
xnor U13089 (N_13089,N_12487,N_12434);
nor U13090 (N_13090,N_12871,N_12184);
xnor U13091 (N_13091,N_12277,N_12508);
or U13092 (N_13092,N_12583,N_12612);
nand U13093 (N_13093,N_12326,N_12444);
nand U13094 (N_13094,N_12842,N_12033);
nand U13095 (N_13095,N_12282,N_12955);
xnor U13096 (N_13096,N_12321,N_12645);
nor U13097 (N_13097,N_12808,N_12944);
xor U13098 (N_13098,N_12724,N_12825);
and U13099 (N_13099,N_12929,N_12958);
and U13100 (N_13100,N_12491,N_12493);
nand U13101 (N_13101,N_12695,N_12380);
nor U13102 (N_13102,N_12744,N_12523);
nor U13103 (N_13103,N_12859,N_12712);
and U13104 (N_13104,N_12292,N_12361);
nor U13105 (N_13105,N_12485,N_12236);
xnor U13106 (N_13106,N_12677,N_12046);
nand U13107 (N_13107,N_12003,N_12221);
xnor U13108 (N_13108,N_12708,N_12403);
and U13109 (N_13109,N_12530,N_12304);
nor U13110 (N_13110,N_12987,N_12050);
nand U13111 (N_13111,N_12738,N_12464);
xor U13112 (N_13112,N_12599,N_12758);
nand U13113 (N_13113,N_12268,N_12624);
and U13114 (N_13114,N_12389,N_12840);
nor U13115 (N_13115,N_12863,N_12699);
xnor U13116 (N_13116,N_12919,N_12714);
and U13117 (N_13117,N_12340,N_12428);
xnor U13118 (N_13118,N_12564,N_12157);
nand U13119 (N_13119,N_12587,N_12582);
xor U13120 (N_13120,N_12298,N_12060);
xor U13121 (N_13121,N_12894,N_12334);
and U13122 (N_13122,N_12507,N_12903);
nor U13123 (N_13123,N_12254,N_12078);
and U13124 (N_13124,N_12989,N_12386);
and U13125 (N_13125,N_12263,N_12122);
xnor U13126 (N_13126,N_12472,N_12328);
or U13127 (N_13127,N_12234,N_12727);
xnor U13128 (N_13128,N_12465,N_12796);
or U13129 (N_13129,N_12213,N_12187);
nand U13130 (N_13130,N_12432,N_12740);
xor U13131 (N_13131,N_12591,N_12473);
and U13132 (N_13132,N_12820,N_12295);
or U13133 (N_13133,N_12174,N_12666);
and U13134 (N_13134,N_12986,N_12025);
and U13135 (N_13135,N_12378,N_12662);
and U13136 (N_13136,N_12548,N_12433);
and U13137 (N_13137,N_12160,N_12531);
xor U13138 (N_13138,N_12565,N_12074);
nor U13139 (N_13139,N_12316,N_12113);
xnor U13140 (N_13140,N_12880,N_12688);
xor U13141 (N_13141,N_12497,N_12482);
xor U13142 (N_13142,N_12488,N_12348);
nor U13143 (N_13143,N_12541,N_12147);
nor U13144 (N_13144,N_12713,N_12844);
nand U13145 (N_13145,N_12105,N_12590);
and U13146 (N_13146,N_12463,N_12600);
nand U13147 (N_13147,N_12671,N_12072);
xor U13148 (N_13148,N_12504,N_12867);
and U13149 (N_13149,N_12089,N_12313);
or U13150 (N_13150,N_12761,N_12908);
nor U13151 (N_13151,N_12349,N_12745);
or U13152 (N_13152,N_12346,N_12961);
and U13153 (N_13153,N_12151,N_12874);
nand U13154 (N_13154,N_12934,N_12500);
or U13155 (N_13155,N_12440,N_12553);
nand U13156 (N_13156,N_12144,N_12764);
and U13157 (N_13157,N_12652,N_12786);
and U13158 (N_13158,N_12299,N_12732);
and U13159 (N_13159,N_12848,N_12581);
or U13160 (N_13160,N_12766,N_12931);
nand U13161 (N_13161,N_12209,N_12200);
and U13162 (N_13162,N_12814,N_12809);
and U13163 (N_13163,N_12280,N_12047);
nor U13164 (N_13164,N_12861,N_12648);
or U13165 (N_13165,N_12800,N_12302);
and U13166 (N_13166,N_12634,N_12938);
or U13167 (N_13167,N_12218,N_12979);
xor U13168 (N_13168,N_12018,N_12715);
nand U13169 (N_13169,N_12196,N_12836);
nand U13170 (N_13170,N_12159,N_12574);
xnor U13171 (N_13171,N_12837,N_12351);
and U13172 (N_13172,N_12593,N_12486);
or U13173 (N_13173,N_12968,N_12609);
or U13174 (N_13174,N_12296,N_12009);
and U13175 (N_13175,N_12872,N_12957);
xor U13176 (N_13176,N_12982,N_12918);
xnor U13177 (N_13177,N_12802,N_12112);
or U13178 (N_13178,N_12772,N_12700);
or U13179 (N_13179,N_12139,N_12454);
xnor U13180 (N_13180,N_12676,N_12069);
nand U13181 (N_13181,N_12245,N_12992);
xor U13182 (N_13182,N_12344,N_12835);
and U13183 (N_13183,N_12211,N_12376);
nand U13184 (N_13184,N_12120,N_12225);
xnor U13185 (N_13185,N_12625,N_12984);
and U13186 (N_13186,N_12747,N_12096);
xnor U13187 (N_13187,N_12275,N_12084);
nand U13188 (N_13188,N_12264,N_12954);
or U13189 (N_13189,N_12385,N_12743);
or U13190 (N_13190,N_12108,N_12686);
xor U13191 (N_13191,N_12407,N_12300);
xor U13192 (N_13192,N_12023,N_12650);
nand U13193 (N_13193,N_12723,N_12717);
or U13194 (N_13194,N_12963,N_12350);
or U13195 (N_13195,N_12922,N_12594);
or U13196 (N_13196,N_12606,N_12754);
xnor U13197 (N_13197,N_12308,N_12595);
nand U13198 (N_13198,N_12851,N_12857);
or U13199 (N_13199,N_12529,N_12019);
and U13200 (N_13200,N_12191,N_12860);
and U13201 (N_13201,N_12536,N_12008);
or U13202 (N_13202,N_12058,N_12601);
nor U13203 (N_13203,N_12347,N_12158);
nor U13204 (N_13204,N_12629,N_12237);
xnor U13205 (N_13205,N_12399,N_12907);
nand U13206 (N_13206,N_12605,N_12244);
xnor U13207 (N_13207,N_12830,N_12966);
nand U13208 (N_13208,N_12767,N_12179);
xnor U13209 (N_13209,N_12062,N_12336);
xor U13210 (N_13210,N_12517,N_12679);
xor U13211 (N_13211,N_12276,N_12034);
xnor U13212 (N_13212,N_12694,N_12036);
or U13213 (N_13213,N_12794,N_12828);
nor U13214 (N_13214,N_12294,N_12087);
xnor U13215 (N_13215,N_12017,N_12692);
nor U13216 (N_13216,N_12458,N_12164);
or U13217 (N_13217,N_12439,N_12673);
and U13218 (N_13218,N_12208,N_12792);
nand U13219 (N_13219,N_12524,N_12878);
nor U13220 (N_13220,N_12022,N_12106);
nand U13221 (N_13221,N_12598,N_12554);
or U13222 (N_13222,N_12217,N_12479);
nand U13223 (N_13223,N_12621,N_12445);
nand U13224 (N_13224,N_12260,N_12812);
nand U13225 (N_13225,N_12924,N_12779);
nor U13226 (N_13226,N_12216,N_12226);
nor U13227 (N_13227,N_12222,N_12626);
xor U13228 (N_13228,N_12567,N_12140);
nand U13229 (N_13229,N_12510,N_12819);
and U13230 (N_13230,N_12735,N_12616);
nor U13231 (N_13231,N_12799,N_12014);
nor U13232 (N_13232,N_12900,N_12885);
and U13233 (N_13233,N_12251,N_12450);
and U13234 (N_13234,N_12569,N_12750);
and U13235 (N_13235,N_12866,N_12004);
xor U13236 (N_13236,N_12572,N_12869);
nor U13237 (N_13237,N_12707,N_12130);
xnor U13238 (N_13238,N_12395,N_12675);
and U13239 (N_13239,N_12663,N_12864);
xnor U13240 (N_13240,N_12398,N_12301);
xor U13241 (N_13241,N_12411,N_12559);
xnor U13242 (N_13242,N_12839,N_12026);
xnor U13243 (N_13243,N_12467,N_12996);
or U13244 (N_13244,N_12307,N_12821);
or U13245 (N_13245,N_12212,N_12771);
nand U13246 (N_13246,N_12015,N_12791);
or U13247 (N_13247,N_12932,N_12604);
nand U13248 (N_13248,N_12448,N_12575);
or U13249 (N_13249,N_12341,N_12180);
nor U13250 (N_13250,N_12318,N_12373);
nor U13251 (N_13251,N_12933,N_12259);
or U13252 (N_13252,N_12161,N_12782);
or U13253 (N_13253,N_12312,N_12188);
or U13254 (N_13254,N_12494,N_12358);
nand U13255 (N_13255,N_12170,N_12056);
and U13256 (N_13256,N_12207,N_12006);
nor U13257 (N_13257,N_12807,N_12066);
and U13258 (N_13258,N_12255,N_12719);
nor U13259 (N_13259,N_12558,N_12476);
or U13260 (N_13260,N_12417,N_12031);
nand U13261 (N_13261,N_12797,N_12876);
nand U13262 (N_13262,N_12670,N_12870);
and U13263 (N_13263,N_12990,N_12462);
and U13264 (N_13264,N_12829,N_12012);
nor U13265 (N_13265,N_12865,N_12853);
xnor U13266 (N_13266,N_12082,N_12503);
nand U13267 (N_13267,N_12974,N_12024);
xor U13268 (N_13268,N_12627,N_12383);
nand U13269 (N_13269,N_12355,N_12369);
xor U13270 (N_13270,N_12956,N_12381);
or U13271 (N_13271,N_12173,N_12231);
xnor U13272 (N_13272,N_12608,N_12387);
or U13273 (N_13273,N_12506,N_12415);
nand U13274 (N_13274,N_12739,N_12149);
xnor U13275 (N_13275,N_12997,N_12401);
and U13276 (N_13276,N_12854,N_12452);
and U13277 (N_13277,N_12535,N_12831);
nor U13278 (N_13278,N_12729,N_12248);
nand U13279 (N_13279,N_12832,N_12843);
nand U13280 (N_13280,N_12091,N_12272);
xor U13281 (N_13281,N_12939,N_12333);
xnor U13282 (N_13282,N_12095,N_12397);
nand U13283 (N_13283,N_12311,N_12429);
xnor U13284 (N_13284,N_12538,N_12001);
or U13285 (N_13285,N_12391,N_12416);
or U13286 (N_13286,N_12680,N_12265);
or U13287 (N_13287,N_12978,N_12285);
nor U13288 (N_13288,N_12881,N_12672);
nand U13289 (N_13289,N_12586,N_12356);
nor U13290 (N_13290,N_12215,N_12468);
xnor U13291 (N_13291,N_12273,N_12827);
or U13292 (N_13292,N_12102,N_12852);
and U13293 (N_13293,N_12038,N_12252);
nand U13294 (N_13294,N_12512,N_12516);
and U13295 (N_13295,N_12288,N_12129);
nand U13296 (N_13296,N_12522,N_12400);
or U13297 (N_13297,N_12042,N_12267);
and U13298 (N_13298,N_12850,N_12256);
nor U13299 (N_13299,N_12610,N_12804);
and U13300 (N_13300,N_12028,N_12090);
or U13301 (N_13301,N_12556,N_12124);
or U13302 (N_13302,N_12889,N_12722);
and U13303 (N_13303,N_12734,N_12240);
xor U13304 (N_13304,N_12741,N_12000);
or U13305 (N_13305,N_12413,N_12297);
nor U13306 (N_13306,N_12641,N_12115);
nor U13307 (N_13307,N_12121,N_12097);
and U13308 (N_13308,N_12988,N_12528);
nand U13309 (N_13309,N_12893,N_12195);
or U13310 (N_13310,N_12201,N_12921);
nor U13311 (N_13311,N_12525,N_12262);
or U13312 (N_13312,N_12847,N_12243);
or U13313 (N_13313,N_12884,N_12570);
nor U13314 (N_13314,N_12620,N_12011);
or U13315 (N_13315,N_12705,N_12071);
or U13316 (N_13316,N_12109,N_12746);
xor U13317 (N_13317,N_12466,N_12951);
nand U13318 (N_13318,N_12394,N_12970);
nor U13319 (N_13319,N_12345,N_12783);
nand U13320 (N_13320,N_12905,N_12916);
and U13321 (N_13321,N_12646,N_12873);
and U13322 (N_13322,N_12029,N_12909);
nor U13323 (N_13323,N_12913,N_12214);
nor U13324 (N_13324,N_12897,N_12379);
xor U13325 (N_13325,N_12975,N_12994);
xnor U13326 (N_13326,N_12681,N_12199);
xor U13327 (N_13327,N_12622,N_12375);
or U13328 (N_13328,N_12937,N_12892);
or U13329 (N_13329,N_12410,N_12759);
xnor U13330 (N_13330,N_12178,N_12737);
xor U13331 (N_13331,N_12678,N_12689);
and U13332 (N_13332,N_12784,N_12136);
nor U13333 (N_13333,N_12703,N_12813);
and U13334 (N_13334,N_12882,N_12143);
nor U13335 (N_13335,N_12817,N_12366);
or U13336 (N_13336,N_12206,N_12659);
xnor U13337 (N_13337,N_12431,N_12765);
and U13338 (N_13338,N_12886,N_12632);
nand U13339 (N_13339,N_12948,N_12368);
or U13340 (N_13340,N_12636,N_12155);
nor U13341 (N_13341,N_12040,N_12169);
nand U13342 (N_13342,N_12945,N_12175);
xor U13343 (N_13343,N_12756,N_12953);
nand U13344 (N_13344,N_12064,N_12329);
and U13345 (N_13345,N_12238,N_12685);
or U13346 (N_13346,N_12075,N_12104);
nand U13347 (N_13347,N_12451,N_12396);
nand U13348 (N_13348,N_12279,N_12716);
xnor U13349 (N_13349,N_12563,N_12331);
and U13350 (N_13350,N_12323,N_12618);
and U13351 (N_13351,N_12027,N_12239);
xor U13352 (N_13352,N_12668,N_12406);
nor U13353 (N_13353,N_12901,N_12291);
nand U13354 (N_13354,N_12198,N_12822);
nor U13355 (N_13355,N_12100,N_12749);
xor U13356 (N_13356,N_12585,N_12010);
nand U13357 (N_13357,N_12841,N_12936);
nand U13358 (N_13358,N_12405,N_12623);
xor U13359 (N_13359,N_12438,N_12030);
and U13360 (N_13360,N_12602,N_12258);
or U13361 (N_13361,N_12210,N_12890);
nor U13362 (N_13362,N_12923,N_12305);
nand U13363 (N_13363,N_12441,N_12877);
xnor U13364 (N_13364,N_12224,N_12615);
and U13365 (N_13365,N_12422,N_12049);
or U13366 (N_13366,N_12135,N_12189);
and U13367 (N_13367,N_12470,N_12220);
xnor U13368 (N_13368,N_12898,N_12935);
nor U13369 (N_13369,N_12787,N_12502);
or U13370 (N_13370,N_12460,N_12414);
xnor U13371 (N_13371,N_12920,N_12549);
xnor U13372 (N_13372,N_12314,N_12167);
xnor U13373 (N_13373,N_12421,N_12941);
xnor U13374 (N_13374,N_12596,N_12785);
nand U13375 (N_13375,N_12657,N_12123);
and U13376 (N_13376,N_12544,N_12770);
and U13377 (N_13377,N_12628,N_12284);
and U13378 (N_13378,N_12862,N_12736);
and U13379 (N_13379,N_12654,N_12088);
and U13380 (N_13380,N_12578,N_12156);
nand U13381 (N_13381,N_12943,N_12233);
xnor U13382 (N_13382,N_12457,N_12021);
nor U13383 (N_13383,N_12176,N_12781);
nand U13384 (N_13384,N_12228,N_12834);
or U13385 (N_13385,N_12942,N_12562);
nor U13386 (N_13386,N_12477,N_12999);
xnor U13387 (N_13387,N_12219,N_12696);
nor U13388 (N_13388,N_12505,N_12437);
xnor U13389 (N_13389,N_12780,N_12153);
and U13390 (N_13390,N_12887,N_12138);
and U13391 (N_13391,N_12967,N_12327);
xnor U13392 (N_13392,N_12742,N_12310);
xnor U13393 (N_13393,N_12910,N_12838);
nor U13394 (N_13394,N_12588,N_12182);
nor U13395 (N_13395,N_12367,N_12132);
nor U13396 (N_13396,N_12805,N_12204);
nand U13397 (N_13397,N_12833,N_12194);
or U13398 (N_13398,N_12499,N_12181);
and U13399 (N_13399,N_12637,N_12952);
or U13400 (N_13400,N_12489,N_12142);
xnor U13401 (N_13401,N_12081,N_12094);
and U13402 (N_13402,N_12227,N_12664);
nand U13403 (N_13403,N_12125,N_12402);
or U13404 (N_13404,N_12229,N_12342);
xor U13405 (N_13405,N_12246,N_12007);
xnor U13406 (N_13406,N_12110,N_12902);
or U13407 (N_13407,N_12718,N_12879);
xnor U13408 (N_13408,N_12534,N_12039);
xor U13409 (N_13409,N_12550,N_12166);
or U13410 (N_13410,N_12725,N_12148);
or U13411 (N_13411,N_12730,N_12203);
and U13412 (N_13412,N_12514,N_12093);
or U13413 (N_13413,N_12647,N_12501);
or U13414 (N_13414,N_12925,N_12755);
nor U13415 (N_13415,N_12691,N_12511);
nand U13416 (N_13416,N_12775,N_12388);
nand U13417 (N_13417,N_12698,N_12449);
or U13418 (N_13418,N_12631,N_12607);
xor U13419 (N_13419,N_12352,N_12162);
nand U13420 (N_13420,N_12845,N_12778);
and U13421 (N_13421,N_12762,N_12768);
and U13422 (N_13422,N_12048,N_12205);
nand U13423 (N_13423,N_12701,N_12555);
nor U13424 (N_13424,N_12888,N_12359);
nor U13425 (N_13425,N_12435,N_12846);
nand U13426 (N_13426,N_12826,N_12849);
nand U13427 (N_13427,N_12532,N_12660);
nor U13428 (N_13428,N_12261,N_12382);
nand U13429 (N_13429,N_12051,N_12163);
nand U13430 (N_13430,N_12490,N_12377);
nor U13431 (N_13431,N_12057,N_12152);
or U13432 (N_13432,N_12459,N_12520);
or U13433 (N_13433,N_12393,N_12669);
and U13434 (N_13434,N_12537,N_12131);
and U13435 (N_13435,N_12690,N_12045);
xnor U13436 (N_13436,N_12940,N_12374);
nand U13437 (N_13437,N_12253,N_12287);
or U13438 (N_13438,N_12899,N_12103);
nor U13439 (N_13439,N_12223,N_12456);
nand U13440 (N_13440,N_12338,N_12638);
nand U13441 (N_13441,N_12823,N_12322);
or U13442 (N_13442,N_12769,N_12858);
xor U13443 (N_13443,N_12309,N_12949);
and U13444 (N_13444,N_12447,N_12710);
nor U13445 (N_13445,N_12810,N_12928);
or U13446 (N_13446,N_12509,N_12667);
nand U13447 (N_13447,N_12977,N_12697);
xnor U13448 (N_13448,N_12972,N_12118);
nor U13449 (N_13449,N_12793,N_12674);
and U13450 (N_13450,N_12561,N_12546);
and U13451 (N_13451,N_12146,N_12235);
nand U13452 (N_13452,N_12926,N_12513);
or U13453 (N_13453,N_12993,N_12526);
xnor U13454 (N_13454,N_12684,N_12016);
and U13455 (N_13455,N_12912,N_12552);
or U13456 (N_13456,N_12748,N_12320);
nor U13457 (N_13457,N_12592,N_12518);
nor U13458 (N_13458,N_12539,N_12073);
nand U13459 (N_13459,N_12168,N_12649);
xnor U13460 (N_13460,N_12190,N_12551);
or U13461 (N_13461,N_12353,N_12436);
xnor U13462 (N_13462,N_12640,N_12757);
nor U13463 (N_13463,N_12965,N_12453);
nand U13464 (N_13464,N_12241,N_12293);
or U13465 (N_13465,N_12154,N_12969);
and U13466 (N_13466,N_12086,N_12250);
or U13467 (N_13467,N_12973,N_12290);
xor U13468 (N_13468,N_12202,N_12726);
or U13469 (N_13469,N_12560,N_12077);
and U13470 (N_13470,N_12469,N_12540);
nor U13471 (N_13471,N_12286,N_12418);
nor U13472 (N_13472,N_12232,N_12911);
nor U13473 (N_13473,N_12384,N_12443);
xnor U13474 (N_13474,N_12408,N_12339);
nor U13475 (N_13475,N_12998,N_12013);
nand U13476 (N_13476,N_12083,N_12037);
or U13477 (N_13477,N_12904,N_12655);
nor U13478 (N_13478,N_12111,N_12611);
nand U13479 (N_13479,N_12566,N_12059);
or U13480 (N_13480,N_12319,N_12020);
and U13481 (N_13481,N_12165,N_12577);
xnor U13482 (N_13482,N_12133,N_12683);
and U13483 (N_13483,N_12790,N_12868);
or U13484 (N_13484,N_12824,N_12580);
or U13485 (N_13485,N_12430,N_12721);
nand U13486 (N_13486,N_12495,N_12547);
nor U13487 (N_13487,N_12906,N_12068);
nor U13488 (N_13488,N_12728,N_12274);
nand U13489 (N_13489,N_12126,N_12044);
nand U13490 (N_13490,N_12959,N_12991);
and U13491 (N_13491,N_12658,N_12343);
nand U13492 (N_13492,N_12653,N_12811);
nand U13493 (N_13493,N_12420,N_12795);
or U13494 (N_13494,N_12052,N_12496);
nand U13495 (N_13495,N_12425,N_12891);
and U13496 (N_13496,N_12271,N_12614);
nor U13497 (N_13497,N_12643,N_12471);
or U13498 (N_13498,N_12542,N_12917);
nor U13499 (N_13499,N_12818,N_12005);
nand U13500 (N_13500,N_12364,N_12404);
nand U13501 (N_13501,N_12047,N_12116);
nor U13502 (N_13502,N_12583,N_12004);
nand U13503 (N_13503,N_12483,N_12269);
xor U13504 (N_13504,N_12634,N_12165);
nand U13505 (N_13505,N_12435,N_12791);
or U13506 (N_13506,N_12465,N_12100);
nand U13507 (N_13507,N_12835,N_12097);
nand U13508 (N_13508,N_12445,N_12001);
nor U13509 (N_13509,N_12923,N_12025);
xnor U13510 (N_13510,N_12918,N_12533);
xnor U13511 (N_13511,N_12525,N_12367);
nor U13512 (N_13512,N_12143,N_12339);
xnor U13513 (N_13513,N_12954,N_12936);
xor U13514 (N_13514,N_12961,N_12102);
xnor U13515 (N_13515,N_12836,N_12924);
nor U13516 (N_13516,N_12550,N_12416);
nor U13517 (N_13517,N_12414,N_12508);
nor U13518 (N_13518,N_12227,N_12630);
nor U13519 (N_13519,N_12534,N_12790);
nand U13520 (N_13520,N_12590,N_12366);
and U13521 (N_13521,N_12768,N_12208);
xnor U13522 (N_13522,N_12981,N_12680);
and U13523 (N_13523,N_12736,N_12984);
nand U13524 (N_13524,N_12951,N_12665);
nor U13525 (N_13525,N_12582,N_12468);
or U13526 (N_13526,N_12502,N_12857);
or U13527 (N_13527,N_12251,N_12709);
xnor U13528 (N_13528,N_12775,N_12591);
xor U13529 (N_13529,N_12785,N_12727);
nor U13530 (N_13530,N_12918,N_12736);
xnor U13531 (N_13531,N_12045,N_12604);
nand U13532 (N_13532,N_12337,N_12059);
xor U13533 (N_13533,N_12868,N_12883);
and U13534 (N_13534,N_12943,N_12968);
xor U13535 (N_13535,N_12084,N_12947);
or U13536 (N_13536,N_12575,N_12568);
nor U13537 (N_13537,N_12312,N_12400);
nor U13538 (N_13538,N_12376,N_12232);
xnor U13539 (N_13539,N_12589,N_12378);
nor U13540 (N_13540,N_12877,N_12516);
or U13541 (N_13541,N_12871,N_12514);
nor U13542 (N_13542,N_12223,N_12347);
nor U13543 (N_13543,N_12641,N_12155);
nor U13544 (N_13544,N_12183,N_12519);
or U13545 (N_13545,N_12917,N_12960);
nand U13546 (N_13546,N_12444,N_12882);
nor U13547 (N_13547,N_12357,N_12149);
or U13548 (N_13548,N_12510,N_12508);
nand U13549 (N_13549,N_12624,N_12958);
nand U13550 (N_13550,N_12781,N_12026);
nand U13551 (N_13551,N_12028,N_12403);
nand U13552 (N_13552,N_12083,N_12664);
or U13553 (N_13553,N_12264,N_12584);
and U13554 (N_13554,N_12922,N_12136);
and U13555 (N_13555,N_12284,N_12996);
nand U13556 (N_13556,N_12951,N_12144);
or U13557 (N_13557,N_12321,N_12881);
and U13558 (N_13558,N_12380,N_12752);
nor U13559 (N_13559,N_12331,N_12302);
nand U13560 (N_13560,N_12311,N_12769);
xnor U13561 (N_13561,N_12217,N_12453);
nor U13562 (N_13562,N_12570,N_12477);
and U13563 (N_13563,N_12267,N_12646);
xnor U13564 (N_13564,N_12182,N_12843);
or U13565 (N_13565,N_12871,N_12003);
and U13566 (N_13566,N_12652,N_12842);
nor U13567 (N_13567,N_12577,N_12585);
xor U13568 (N_13568,N_12445,N_12590);
or U13569 (N_13569,N_12094,N_12037);
nand U13570 (N_13570,N_12304,N_12649);
nor U13571 (N_13571,N_12469,N_12321);
nor U13572 (N_13572,N_12631,N_12918);
and U13573 (N_13573,N_12283,N_12543);
nor U13574 (N_13574,N_12799,N_12752);
and U13575 (N_13575,N_12095,N_12377);
and U13576 (N_13576,N_12266,N_12013);
nand U13577 (N_13577,N_12261,N_12917);
and U13578 (N_13578,N_12408,N_12352);
xor U13579 (N_13579,N_12038,N_12986);
nor U13580 (N_13580,N_12240,N_12440);
nor U13581 (N_13581,N_12561,N_12352);
nand U13582 (N_13582,N_12957,N_12296);
nand U13583 (N_13583,N_12036,N_12770);
or U13584 (N_13584,N_12469,N_12954);
and U13585 (N_13585,N_12190,N_12269);
and U13586 (N_13586,N_12025,N_12170);
xor U13587 (N_13587,N_12775,N_12924);
nor U13588 (N_13588,N_12904,N_12861);
nand U13589 (N_13589,N_12178,N_12720);
and U13590 (N_13590,N_12607,N_12138);
and U13591 (N_13591,N_12250,N_12611);
nor U13592 (N_13592,N_12591,N_12321);
nor U13593 (N_13593,N_12799,N_12464);
xor U13594 (N_13594,N_12114,N_12960);
xnor U13595 (N_13595,N_12787,N_12334);
nand U13596 (N_13596,N_12405,N_12622);
nand U13597 (N_13597,N_12851,N_12951);
or U13598 (N_13598,N_12909,N_12722);
xor U13599 (N_13599,N_12312,N_12332);
or U13600 (N_13600,N_12214,N_12729);
nor U13601 (N_13601,N_12021,N_12353);
or U13602 (N_13602,N_12615,N_12906);
xor U13603 (N_13603,N_12881,N_12779);
and U13604 (N_13604,N_12251,N_12610);
and U13605 (N_13605,N_12534,N_12182);
nand U13606 (N_13606,N_12743,N_12180);
or U13607 (N_13607,N_12297,N_12764);
nand U13608 (N_13608,N_12892,N_12438);
or U13609 (N_13609,N_12425,N_12012);
xnor U13610 (N_13610,N_12261,N_12246);
xnor U13611 (N_13611,N_12733,N_12238);
and U13612 (N_13612,N_12228,N_12648);
xnor U13613 (N_13613,N_12992,N_12540);
nand U13614 (N_13614,N_12415,N_12935);
or U13615 (N_13615,N_12459,N_12222);
and U13616 (N_13616,N_12811,N_12576);
nand U13617 (N_13617,N_12905,N_12884);
nand U13618 (N_13618,N_12425,N_12382);
nor U13619 (N_13619,N_12496,N_12393);
nor U13620 (N_13620,N_12316,N_12749);
nand U13621 (N_13621,N_12948,N_12870);
nor U13622 (N_13622,N_12909,N_12531);
or U13623 (N_13623,N_12209,N_12625);
or U13624 (N_13624,N_12611,N_12666);
xnor U13625 (N_13625,N_12347,N_12606);
nor U13626 (N_13626,N_12450,N_12572);
xnor U13627 (N_13627,N_12453,N_12976);
and U13628 (N_13628,N_12351,N_12885);
xnor U13629 (N_13629,N_12426,N_12006);
or U13630 (N_13630,N_12605,N_12538);
and U13631 (N_13631,N_12553,N_12836);
and U13632 (N_13632,N_12318,N_12075);
and U13633 (N_13633,N_12596,N_12690);
and U13634 (N_13634,N_12134,N_12681);
or U13635 (N_13635,N_12646,N_12179);
nor U13636 (N_13636,N_12717,N_12508);
or U13637 (N_13637,N_12940,N_12932);
xnor U13638 (N_13638,N_12275,N_12870);
or U13639 (N_13639,N_12536,N_12403);
and U13640 (N_13640,N_12061,N_12636);
and U13641 (N_13641,N_12560,N_12908);
and U13642 (N_13642,N_12688,N_12150);
or U13643 (N_13643,N_12561,N_12849);
nor U13644 (N_13644,N_12646,N_12560);
nor U13645 (N_13645,N_12904,N_12971);
nand U13646 (N_13646,N_12754,N_12036);
or U13647 (N_13647,N_12709,N_12420);
and U13648 (N_13648,N_12182,N_12157);
and U13649 (N_13649,N_12675,N_12204);
and U13650 (N_13650,N_12178,N_12022);
nor U13651 (N_13651,N_12177,N_12253);
and U13652 (N_13652,N_12170,N_12735);
nand U13653 (N_13653,N_12714,N_12759);
or U13654 (N_13654,N_12066,N_12023);
xnor U13655 (N_13655,N_12386,N_12162);
and U13656 (N_13656,N_12294,N_12979);
xor U13657 (N_13657,N_12651,N_12709);
nor U13658 (N_13658,N_12901,N_12452);
xor U13659 (N_13659,N_12392,N_12665);
and U13660 (N_13660,N_12735,N_12145);
or U13661 (N_13661,N_12348,N_12428);
or U13662 (N_13662,N_12994,N_12992);
nand U13663 (N_13663,N_12148,N_12731);
nand U13664 (N_13664,N_12917,N_12797);
or U13665 (N_13665,N_12471,N_12934);
and U13666 (N_13666,N_12063,N_12171);
nand U13667 (N_13667,N_12281,N_12617);
nand U13668 (N_13668,N_12582,N_12947);
and U13669 (N_13669,N_12660,N_12515);
and U13670 (N_13670,N_12671,N_12685);
xnor U13671 (N_13671,N_12688,N_12643);
nor U13672 (N_13672,N_12313,N_12162);
or U13673 (N_13673,N_12486,N_12250);
nor U13674 (N_13674,N_12063,N_12360);
xnor U13675 (N_13675,N_12228,N_12142);
nand U13676 (N_13676,N_12000,N_12492);
nand U13677 (N_13677,N_12437,N_12810);
and U13678 (N_13678,N_12653,N_12989);
and U13679 (N_13679,N_12944,N_12080);
nand U13680 (N_13680,N_12169,N_12151);
xnor U13681 (N_13681,N_12073,N_12117);
and U13682 (N_13682,N_12220,N_12668);
or U13683 (N_13683,N_12032,N_12603);
nor U13684 (N_13684,N_12908,N_12549);
nand U13685 (N_13685,N_12315,N_12794);
nand U13686 (N_13686,N_12956,N_12691);
or U13687 (N_13687,N_12798,N_12308);
or U13688 (N_13688,N_12919,N_12276);
or U13689 (N_13689,N_12813,N_12828);
nor U13690 (N_13690,N_12741,N_12286);
or U13691 (N_13691,N_12788,N_12662);
and U13692 (N_13692,N_12251,N_12194);
nand U13693 (N_13693,N_12550,N_12779);
nand U13694 (N_13694,N_12761,N_12658);
nand U13695 (N_13695,N_12235,N_12976);
nand U13696 (N_13696,N_12628,N_12186);
nand U13697 (N_13697,N_12845,N_12449);
nand U13698 (N_13698,N_12512,N_12502);
nor U13699 (N_13699,N_12974,N_12062);
nand U13700 (N_13700,N_12572,N_12885);
xnor U13701 (N_13701,N_12752,N_12288);
and U13702 (N_13702,N_12246,N_12999);
or U13703 (N_13703,N_12792,N_12719);
nor U13704 (N_13704,N_12887,N_12120);
xnor U13705 (N_13705,N_12817,N_12863);
nor U13706 (N_13706,N_12262,N_12694);
and U13707 (N_13707,N_12222,N_12889);
nand U13708 (N_13708,N_12250,N_12561);
nand U13709 (N_13709,N_12961,N_12004);
and U13710 (N_13710,N_12234,N_12475);
or U13711 (N_13711,N_12256,N_12209);
nor U13712 (N_13712,N_12450,N_12555);
and U13713 (N_13713,N_12116,N_12831);
nor U13714 (N_13714,N_12466,N_12162);
xor U13715 (N_13715,N_12977,N_12123);
xor U13716 (N_13716,N_12833,N_12265);
nor U13717 (N_13717,N_12311,N_12976);
nor U13718 (N_13718,N_12137,N_12110);
nor U13719 (N_13719,N_12159,N_12755);
or U13720 (N_13720,N_12580,N_12594);
or U13721 (N_13721,N_12642,N_12303);
or U13722 (N_13722,N_12132,N_12381);
or U13723 (N_13723,N_12704,N_12804);
and U13724 (N_13724,N_12268,N_12550);
or U13725 (N_13725,N_12299,N_12917);
nor U13726 (N_13726,N_12774,N_12942);
nand U13727 (N_13727,N_12143,N_12227);
nor U13728 (N_13728,N_12567,N_12633);
xor U13729 (N_13729,N_12724,N_12008);
nor U13730 (N_13730,N_12531,N_12630);
nand U13731 (N_13731,N_12021,N_12999);
and U13732 (N_13732,N_12239,N_12736);
or U13733 (N_13733,N_12941,N_12730);
or U13734 (N_13734,N_12712,N_12729);
and U13735 (N_13735,N_12967,N_12517);
or U13736 (N_13736,N_12419,N_12110);
and U13737 (N_13737,N_12876,N_12834);
nand U13738 (N_13738,N_12953,N_12970);
or U13739 (N_13739,N_12699,N_12234);
nor U13740 (N_13740,N_12617,N_12662);
or U13741 (N_13741,N_12695,N_12541);
and U13742 (N_13742,N_12720,N_12523);
xor U13743 (N_13743,N_12053,N_12049);
nor U13744 (N_13744,N_12127,N_12866);
and U13745 (N_13745,N_12438,N_12139);
xor U13746 (N_13746,N_12185,N_12798);
nand U13747 (N_13747,N_12514,N_12557);
and U13748 (N_13748,N_12263,N_12583);
xor U13749 (N_13749,N_12218,N_12484);
nand U13750 (N_13750,N_12493,N_12411);
nand U13751 (N_13751,N_12178,N_12710);
nand U13752 (N_13752,N_12953,N_12744);
and U13753 (N_13753,N_12480,N_12966);
or U13754 (N_13754,N_12097,N_12762);
xnor U13755 (N_13755,N_12121,N_12567);
or U13756 (N_13756,N_12323,N_12962);
xnor U13757 (N_13757,N_12667,N_12059);
xnor U13758 (N_13758,N_12567,N_12571);
and U13759 (N_13759,N_12026,N_12449);
or U13760 (N_13760,N_12382,N_12398);
xor U13761 (N_13761,N_12341,N_12812);
and U13762 (N_13762,N_12774,N_12579);
and U13763 (N_13763,N_12782,N_12686);
or U13764 (N_13764,N_12446,N_12490);
and U13765 (N_13765,N_12575,N_12745);
or U13766 (N_13766,N_12350,N_12179);
nor U13767 (N_13767,N_12249,N_12474);
and U13768 (N_13768,N_12971,N_12374);
nor U13769 (N_13769,N_12501,N_12261);
and U13770 (N_13770,N_12479,N_12763);
or U13771 (N_13771,N_12869,N_12317);
or U13772 (N_13772,N_12459,N_12211);
and U13773 (N_13773,N_12975,N_12463);
nand U13774 (N_13774,N_12678,N_12918);
nand U13775 (N_13775,N_12012,N_12524);
or U13776 (N_13776,N_12931,N_12995);
or U13777 (N_13777,N_12859,N_12143);
or U13778 (N_13778,N_12656,N_12357);
and U13779 (N_13779,N_12338,N_12685);
xor U13780 (N_13780,N_12035,N_12474);
nor U13781 (N_13781,N_12247,N_12930);
xnor U13782 (N_13782,N_12414,N_12502);
xor U13783 (N_13783,N_12081,N_12164);
nand U13784 (N_13784,N_12867,N_12321);
nand U13785 (N_13785,N_12928,N_12663);
or U13786 (N_13786,N_12448,N_12393);
xor U13787 (N_13787,N_12300,N_12474);
nor U13788 (N_13788,N_12576,N_12425);
nor U13789 (N_13789,N_12468,N_12314);
nand U13790 (N_13790,N_12975,N_12909);
nand U13791 (N_13791,N_12544,N_12905);
and U13792 (N_13792,N_12939,N_12359);
and U13793 (N_13793,N_12758,N_12404);
and U13794 (N_13794,N_12560,N_12549);
xor U13795 (N_13795,N_12913,N_12515);
xnor U13796 (N_13796,N_12114,N_12057);
or U13797 (N_13797,N_12704,N_12882);
and U13798 (N_13798,N_12411,N_12653);
or U13799 (N_13799,N_12209,N_12847);
nand U13800 (N_13800,N_12785,N_12220);
nand U13801 (N_13801,N_12778,N_12091);
nand U13802 (N_13802,N_12479,N_12881);
or U13803 (N_13803,N_12543,N_12324);
nor U13804 (N_13804,N_12477,N_12410);
nand U13805 (N_13805,N_12531,N_12078);
nor U13806 (N_13806,N_12752,N_12500);
nand U13807 (N_13807,N_12203,N_12928);
nor U13808 (N_13808,N_12812,N_12593);
nor U13809 (N_13809,N_12200,N_12547);
nand U13810 (N_13810,N_12160,N_12515);
nor U13811 (N_13811,N_12231,N_12406);
and U13812 (N_13812,N_12352,N_12032);
nand U13813 (N_13813,N_12400,N_12663);
and U13814 (N_13814,N_12855,N_12319);
xnor U13815 (N_13815,N_12805,N_12519);
nor U13816 (N_13816,N_12906,N_12612);
nand U13817 (N_13817,N_12132,N_12077);
xor U13818 (N_13818,N_12030,N_12788);
nand U13819 (N_13819,N_12263,N_12018);
xor U13820 (N_13820,N_12575,N_12596);
nand U13821 (N_13821,N_12788,N_12383);
and U13822 (N_13822,N_12467,N_12669);
xnor U13823 (N_13823,N_12779,N_12826);
xnor U13824 (N_13824,N_12443,N_12078);
nor U13825 (N_13825,N_12633,N_12436);
nor U13826 (N_13826,N_12187,N_12373);
xor U13827 (N_13827,N_12509,N_12665);
nand U13828 (N_13828,N_12058,N_12256);
xor U13829 (N_13829,N_12674,N_12588);
or U13830 (N_13830,N_12076,N_12945);
and U13831 (N_13831,N_12204,N_12018);
nand U13832 (N_13832,N_12762,N_12793);
nor U13833 (N_13833,N_12416,N_12673);
nand U13834 (N_13834,N_12154,N_12490);
xor U13835 (N_13835,N_12234,N_12314);
xnor U13836 (N_13836,N_12661,N_12308);
xor U13837 (N_13837,N_12868,N_12983);
xor U13838 (N_13838,N_12878,N_12340);
nor U13839 (N_13839,N_12687,N_12617);
and U13840 (N_13840,N_12106,N_12477);
and U13841 (N_13841,N_12004,N_12314);
or U13842 (N_13842,N_12182,N_12329);
and U13843 (N_13843,N_12437,N_12502);
and U13844 (N_13844,N_12063,N_12177);
xnor U13845 (N_13845,N_12594,N_12095);
nand U13846 (N_13846,N_12267,N_12526);
nand U13847 (N_13847,N_12572,N_12189);
nor U13848 (N_13848,N_12929,N_12538);
or U13849 (N_13849,N_12772,N_12050);
xnor U13850 (N_13850,N_12306,N_12643);
xor U13851 (N_13851,N_12189,N_12070);
nand U13852 (N_13852,N_12360,N_12762);
nor U13853 (N_13853,N_12730,N_12711);
nand U13854 (N_13854,N_12659,N_12079);
nand U13855 (N_13855,N_12747,N_12020);
and U13856 (N_13856,N_12196,N_12104);
and U13857 (N_13857,N_12319,N_12619);
or U13858 (N_13858,N_12846,N_12555);
nor U13859 (N_13859,N_12820,N_12088);
and U13860 (N_13860,N_12415,N_12101);
nand U13861 (N_13861,N_12510,N_12525);
nand U13862 (N_13862,N_12722,N_12665);
nand U13863 (N_13863,N_12075,N_12409);
nor U13864 (N_13864,N_12640,N_12963);
nor U13865 (N_13865,N_12608,N_12124);
nand U13866 (N_13866,N_12337,N_12618);
and U13867 (N_13867,N_12660,N_12969);
or U13868 (N_13868,N_12770,N_12383);
nor U13869 (N_13869,N_12905,N_12279);
nor U13870 (N_13870,N_12507,N_12950);
and U13871 (N_13871,N_12737,N_12398);
or U13872 (N_13872,N_12446,N_12149);
nor U13873 (N_13873,N_12933,N_12947);
or U13874 (N_13874,N_12383,N_12630);
nand U13875 (N_13875,N_12326,N_12389);
nand U13876 (N_13876,N_12239,N_12523);
and U13877 (N_13877,N_12337,N_12767);
nor U13878 (N_13878,N_12346,N_12937);
nand U13879 (N_13879,N_12409,N_12441);
xnor U13880 (N_13880,N_12147,N_12714);
and U13881 (N_13881,N_12248,N_12754);
and U13882 (N_13882,N_12066,N_12141);
nor U13883 (N_13883,N_12095,N_12195);
and U13884 (N_13884,N_12749,N_12486);
nand U13885 (N_13885,N_12172,N_12986);
nand U13886 (N_13886,N_12683,N_12453);
nor U13887 (N_13887,N_12174,N_12222);
nor U13888 (N_13888,N_12746,N_12704);
and U13889 (N_13889,N_12963,N_12508);
and U13890 (N_13890,N_12517,N_12422);
or U13891 (N_13891,N_12138,N_12557);
nor U13892 (N_13892,N_12991,N_12865);
or U13893 (N_13893,N_12116,N_12746);
nand U13894 (N_13894,N_12313,N_12538);
nand U13895 (N_13895,N_12953,N_12388);
xnor U13896 (N_13896,N_12530,N_12697);
nor U13897 (N_13897,N_12733,N_12118);
or U13898 (N_13898,N_12948,N_12812);
xor U13899 (N_13899,N_12420,N_12189);
or U13900 (N_13900,N_12130,N_12544);
nor U13901 (N_13901,N_12279,N_12189);
xor U13902 (N_13902,N_12993,N_12687);
or U13903 (N_13903,N_12464,N_12572);
nor U13904 (N_13904,N_12573,N_12287);
or U13905 (N_13905,N_12533,N_12100);
and U13906 (N_13906,N_12767,N_12505);
and U13907 (N_13907,N_12900,N_12476);
and U13908 (N_13908,N_12448,N_12503);
nand U13909 (N_13909,N_12144,N_12277);
xor U13910 (N_13910,N_12826,N_12592);
nor U13911 (N_13911,N_12743,N_12868);
xnor U13912 (N_13912,N_12690,N_12171);
xor U13913 (N_13913,N_12026,N_12334);
and U13914 (N_13914,N_12380,N_12734);
and U13915 (N_13915,N_12238,N_12634);
nor U13916 (N_13916,N_12511,N_12726);
nand U13917 (N_13917,N_12908,N_12730);
nor U13918 (N_13918,N_12174,N_12912);
or U13919 (N_13919,N_12351,N_12592);
xor U13920 (N_13920,N_12189,N_12169);
and U13921 (N_13921,N_12596,N_12086);
and U13922 (N_13922,N_12475,N_12330);
nand U13923 (N_13923,N_12148,N_12358);
nand U13924 (N_13924,N_12097,N_12333);
nand U13925 (N_13925,N_12880,N_12067);
and U13926 (N_13926,N_12787,N_12962);
and U13927 (N_13927,N_12788,N_12007);
or U13928 (N_13928,N_12890,N_12768);
and U13929 (N_13929,N_12653,N_12658);
xnor U13930 (N_13930,N_12880,N_12881);
nand U13931 (N_13931,N_12896,N_12016);
nand U13932 (N_13932,N_12414,N_12366);
and U13933 (N_13933,N_12489,N_12018);
or U13934 (N_13934,N_12917,N_12320);
and U13935 (N_13935,N_12793,N_12825);
xnor U13936 (N_13936,N_12848,N_12409);
or U13937 (N_13937,N_12159,N_12110);
or U13938 (N_13938,N_12118,N_12732);
or U13939 (N_13939,N_12569,N_12972);
xnor U13940 (N_13940,N_12517,N_12380);
nand U13941 (N_13941,N_12782,N_12077);
and U13942 (N_13942,N_12757,N_12391);
nor U13943 (N_13943,N_12824,N_12197);
nor U13944 (N_13944,N_12082,N_12411);
xnor U13945 (N_13945,N_12202,N_12255);
xnor U13946 (N_13946,N_12617,N_12088);
or U13947 (N_13947,N_12036,N_12409);
or U13948 (N_13948,N_12742,N_12297);
and U13949 (N_13949,N_12153,N_12831);
nand U13950 (N_13950,N_12350,N_12400);
nor U13951 (N_13951,N_12237,N_12621);
or U13952 (N_13952,N_12086,N_12091);
or U13953 (N_13953,N_12557,N_12352);
and U13954 (N_13954,N_12223,N_12446);
and U13955 (N_13955,N_12552,N_12777);
xor U13956 (N_13956,N_12167,N_12224);
xor U13957 (N_13957,N_12790,N_12949);
xor U13958 (N_13958,N_12562,N_12844);
or U13959 (N_13959,N_12513,N_12322);
xnor U13960 (N_13960,N_12352,N_12133);
nor U13961 (N_13961,N_12761,N_12237);
xnor U13962 (N_13962,N_12184,N_12695);
and U13963 (N_13963,N_12004,N_12398);
or U13964 (N_13964,N_12956,N_12116);
xor U13965 (N_13965,N_12311,N_12739);
nand U13966 (N_13966,N_12098,N_12560);
nand U13967 (N_13967,N_12644,N_12913);
or U13968 (N_13968,N_12773,N_12998);
or U13969 (N_13969,N_12250,N_12638);
or U13970 (N_13970,N_12463,N_12715);
nand U13971 (N_13971,N_12658,N_12037);
xor U13972 (N_13972,N_12737,N_12341);
nor U13973 (N_13973,N_12289,N_12709);
nand U13974 (N_13974,N_12276,N_12433);
nand U13975 (N_13975,N_12637,N_12615);
nor U13976 (N_13976,N_12324,N_12317);
nand U13977 (N_13977,N_12835,N_12629);
nor U13978 (N_13978,N_12342,N_12277);
xor U13979 (N_13979,N_12878,N_12619);
nor U13980 (N_13980,N_12139,N_12107);
nand U13981 (N_13981,N_12365,N_12377);
xor U13982 (N_13982,N_12726,N_12821);
or U13983 (N_13983,N_12093,N_12263);
and U13984 (N_13984,N_12685,N_12221);
xor U13985 (N_13985,N_12406,N_12544);
and U13986 (N_13986,N_12950,N_12044);
xnor U13987 (N_13987,N_12570,N_12376);
nor U13988 (N_13988,N_12286,N_12607);
and U13989 (N_13989,N_12685,N_12034);
nand U13990 (N_13990,N_12179,N_12122);
or U13991 (N_13991,N_12872,N_12203);
and U13992 (N_13992,N_12218,N_12859);
nor U13993 (N_13993,N_12841,N_12811);
xnor U13994 (N_13994,N_12064,N_12431);
or U13995 (N_13995,N_12151,N_12963);
nor U13996 (N_13996,N_12382,N_12482);
nand U13997 (N_13997,N_12627,N_12785);
nor U13998 (N_13998,N_12062,N_12604);
and U13999 (N_13999,N_12031,N_12826);
xnor U14000 (N_14000,N_13598,N_13038);
nand U14001 (N_14001,N_13166,N_13670);
nand U14002 (N_14002,N_13990,N_13701);
xnor U14003 (N_14003,N_13618,N_13815);
or U14004 (N_14004,N_13274,N_13703);
or U14005 (N_14005,N_13557,N_13828);
and U14006 (N_14006,N_13860,N_13468);
and U14007 (N_14007,N_13880,N_13039);
nor U14008 (N_14008,N_13222,N_13732);
or U14009 (N_14009,N_13040,N_13961);
nor U14010 (N_14010,N_13717,N_13532);
xnor U14011 (N_14011,N_13268,N_13134);
or U14012 (N_14012,N_13693,N_13918);
xnor U14013 (N_14013,N_13839,N_13147);
xnor U14014 (N_14014,N_13031,N_13731);
xor U14015 (N_14015,N_13533,N_13639);
nand U14016 (N_14016,N_13373,N_13615);
nor U14017 (N_14017,N_13509,N_13167);
nor U14018 (N_14018,N_13446,N_13277);
and U14019 (N_14019,N_13762,N_13710);
or U14020 (N_14020,N_13255,N_13494);
nand U14021 (N_14021,N_13515,N_13625);
nand U14022 (N_14022,N_13803,N_13911);
nor U14023 (N_14023,N_13844,N_13170);
or U14024 (N_14024,N_13993,N_13376);
nand U14025 (N_14025,N_13303,N_13979);
xor U14026 (N_14026,N_13884,N_13594);
nand U14027 (N_14027,N_13913,N_13048);
xor U14028 (N_14028,N_13840,N_13435);
or U14029 (N_14029,N_13651,N_13195);
xnor U14030 (N_14030,N_13954,N_13278);
nand U14031 (N_14031,N_13610,N_13320);
and U14032 (N_14032,N_13239,N_13846);
and U14033 (N_14033,N_13292,N_13280);
nor U14034 (N_14034,N_13802,N_13797);
nand U14035 (N_14035,N_13083,N_13930);
nand U14036 (N_14036,N_13460,N_13207);
nand U14037 (N_14037,N_13480,N_13151);
and U14038 (N_14038,N_13978,N_13986);
xor U14039 (N_14039,N_13261,N_13008);
nor U14040 (N_14040,N_13381,N_13496);
nor U14041 (N_14041,N_13365,N_13213);
xor U14042 (N_14042,N_13910,N_13902);
nor U14043 (N_14043,N_13635,N_13115);
nor U14044 (N_14044,N_13069,N_13395);
xor U14045 (N_14045,N_13089,N_13582);
or U14046 (N_14046,N_13872,N_13046);
or U14047 (N_14047,N_13461,N_13338);
nor U14048 (N_14048,N_13003,N_13694);
and U14049 (N_14049,N_13737,N_13560);
or U14050 (N_14050,N_13778,N_13283);
or U14051 (N_14051,N_13226,N_13485);
nand U14052 (N_14052,N_13248,N_13103);
or U14053 (N_14053,N_13223,N_13758);
nor U14054 (N_14054,N_13102,N_13090);
nor U14055 (N_14055,N_13919,N_13956);
nand U14056 (N_14056,N_13315,N_13398);
nor U14057 (N_14057,N_13606,N_13275);
and U14058 (N_14058,N_13153,N_13005);
nor U14059 (N_14059,N_13149,N_13484);
nand U14060 (N_14060,N_13951,N_13947);
and U14061 (N_14061,N_13366,N_13503);
or U14062 (N_14062,N_13835,N_13770);
nor U14063 (N_14063,N_13305,N_13238);
xor U14064 (N_14064,N_13228,N_13440);
and U14065 (N_14065,N_13780,N_13660);
and U14066 (N_14066,N_13209,N_13953);
xor U14067 (N_14067,N_13759,N_13029);
and U14068 (N_14068,N_13092,N_13889);
xnor U14069 (N_14069,N_13112,N_13071);
xnor U14070 (N_14070,N_13895,N_13114);
nor U14071 (N_14071,N_13906,N_13377);
or U14072 (N_14072,N_13413,N_13499);
nor U14073 (N_14073,N_13612,N_13721);
and U14074 (N_14074,N_13129,N_13179);
or U14075 (N_14075,N_13857,N_13944);
or U14076 (N_14076,N_13434,N_13028);
nand U14077 (N_14077,N_13516,N_13536);
nand U14078 (N_14078,N_13394,N_13599);
nor U14079 (N_14079,N_13330,N_13386);
and U14080 (N_14080,N_13804,N_13611);
and U14081 (N_14081,N_13596,N_13816);
xnor U14082 (N_14082,N_13353,N_13309);
or U14083 (N_14083,N_13608,N_13851);
nor U14084 (N_14084,N_13544,N_13357);
nand U14085 (N_14085,N_13319,N_13165);
xnor U14086 (N_14086,N_13959,N_13963);
or U14087 (N_14087,N_13649,N_13314);
xor U14088 (N_14088,N_13010,N_13970);
xnor U14089 (N_14089,N_13571,N_13042);
nand U14090 (N_14090,N_13697,N_13224);
nand U14091 (N_14091,N_13405,N_13217);
nand U14092 (N_14092,N_13080,N_13237);
xnor U14093 (N_14093,N_13367,N_13276);
xor U14094 (N_14094,N_13487,N_13106);
nand U14095 (N_14095,N_13637,N_13766);
nor U14096 (N_14096,N_13297,N_13137);
nor U14097 (N_14097,N_13850,N_13310);
and U14098 (N_14098,N_13282,N_13619);
nand U14099 (N_14099,N_13510,N_13118);
nand U14100 (N_14100,N_13754,N_13871);
nand U14101 (N_14101,N_13156,N_13858);
nor U14102 (N_14102,N_13655,N_13645);
nand U14103 (N_14103,N_13148,N_13643);
and U14104 (N_14104,N_13441,N_13987);
nor U14105 (N_14105,N_13316,N_13519);
or U14106 (N_14106,N_13617,N_13350);
and U14107 (N_14107,N_13502,N_13924);
and U14108 (N_14108,N_13879,N_13359);
and U14109 (N_14109,N_13511,N_13450);
xor U14110 (N_14110,N_13144,N_13836);
or U14111 (N_14111,N_13327,N_13627);
and U14112 (N_14112,N_13607,N_13416);
xor U14113 (N_14113,N_13874,N_13750);
nor U14114 (N_14114,N_13719,N_13454);
xor U14115 (N_14115,N_13541,N_13925);
or U14116 (N_14116,N_13968,N_13425);
nand U14117 (N_14117,N_13231,N_13622);
xnor U14118 (N_14118,N_13674,N_13926);
nor U14119 (N_14119,N_13812,N_13943);
and U14120 (N_14120,N_13855,N_13225);
or U14121 (N_14121,N_13066,N_13025);
nand U14122 (N_14122,N_13734,N_13568);
nand U14123 (N_14123,N_13585,N_13991);
and U14124 (N_14124,N_13623,N_13246);
xor U14125 (N_14125,N_13988,N_13996);
xor U14126 (N_14126,N_13583,N_13322);
xor U14127 (N_14127,N_13154,N_13638);
nor U14128 (N_14128,N_13579,N_13791);
xnor U14129 (N_14129,N_13286,N_13390);
nand U14130 (N_14130,N_13108,N_13837);
nor U14131 (N_14131,N_13853,N_13668);
xnor U14132 (N_14132,N_13636,N_13186);
nand U14133 (N_14133,N_13885,N_13730);
or U14134 (N_14134,N_13937,N_13935);
or U14135 (N_14135,N_13065,N_13783);
nor U14136 (N_14136,N_13894,N_13404);
and U14137 (N_14137,N_13400,N_13244);
xnor U14138 (N_14138,N_13325,N_13577);
and U14139 (N_14139,N_13486,N_13989);
nand U14140 (N_14140,N_13295,N_13574);
or U14141 (N_14141,N_13356,N_13070);
and U14142 (N_14142,N_13540,N_13182);
and U14143 (N_14143,N_13088,N_13145);
and U14144 (N_14144,N_13426,N_13015);
and U14145 (N_14145,N_13584,N_13591);
nor U14146 (N_14146,N_13997,N_13662);
or U14147 (N_14147,N_13221,N_13388);
nor U14148 (N_14148,N_13026,N_13044);
and U14149 (N_14149,N_13266,N_13279);
and U14150 (N_14150,N_13489,N_13210);
nand U14151 (N_14151,N_13984,N_13269);
and U14152 (N_14152,N_13832,N_13698);
or U14153 (N_14153,N_13146,N_13705);
and U14154 (N_14154,N_13001,N_13476);
and U14155 (N_14155,N_13431,N_13795);
xnor U14156 (N_14156,N_13600,N_13251);
or U14157 (N_14157,N_13914,N_13321);
or U14158 (N_14158,N_13392,N_13189);
xnor U14159 (N_14159,N_13604,N_13672);
xor U14160 (N_14160,N_13813,N_13328);
xnor U14161 (N_14161,N_13014,N_13774);
and U14162 (N_14162,N_13477,N_13856);
or U14163 (N_14163,N_13180,N_13825);
xnor U14164 (N_14164,N_13983,N_13899);
nand U14165 (N_14165,N_13686,N_13082);
xnor U14166 (N_14166,N_13534,N_13423);
xnor U14167 (N_14167,N_13401,N_13634);
nand U14168 (N_14168,N_13518,N_13415);
nor U14169 (N_14169,N_13027,N_13666);
nand U14170 (N_14170,N_13708,N_13729);
or U14171 (N_14171,N_13202,N_13587);
and U14172 (N_14172,N_13807,N_13957);
nor U14173 (N_14173,N_13535,N_13669);
and U14174 (N_14174,N_13054,N_13525);
nand U14175 (N_14175,N_13692,N_13427);
nand U14176 (N_14176,N_13863,N_13784);
nand U14177 (N_14177,N_13234,N_13020);
nor U14178 (N_14178,N_13036,N_13301);
nor U14179 (N_14179,N_13445,N_13652);
and U14180 (N_14180,N_13363,N_13581);
or U14181 (N_14181,N_13420,N_13590);
or U14182 (N_14182,N_13756,N_13138);
nand U14183 (N_14183,N_13539,N_13051);
or U14184 (N_14184,N_13827,N_13869);
or U14185 (N_14185,N_13281,N_13861);
and U14186 (N_14186,N_13826,N_13626);
or U14187 (N_14187,N_13616,N_13449);
xor U14188 (N_14188,N_13785,N_13007);
nand U14189 (N_14189,N_13592,N_13665);
nand U14190 (N_14190,N_13247,N_13702);
or U14191 (N_14191,N_13892,N_13467);
or U14192 (N_14192,N_13849,N_13272);
xor U14193 (N_14193,N_13142,N_13864);
nand U14194 (N_14194,N_13972,N_13820);
nor U14195 (N_14195,N_13459,N_13941);
or U14196 (N_14196,N_13776,N_13444);
xnor U14197 (N_14197,N_13707,N_13341);
nor U14198 (N_14198,N_13706,N_13862);
and U14199 (N_14199,N_13677,N_13260);
xnor U14200 (N_14200,N_13883,N_13160);
or U14201 (N_14201,N_13920,N_13609);
and U14202 (N_14202,N_13829,N_13249);
and U14203 (N_14203,N_13308,N_13159);
or U14204 (N_14204,N_13663,N_13412);
nand U14205 (N_14205,N_13973,N_13999);
or U14206 (N_14206,N_13746,N_13220);
and U14207 (N_14207,N_13346,N_13464);
nor U14208 (N_14208,N_13399,N_13711);
xnor U14209 (N_14209,N_13075,N_13882);
xor U14210 (N_14210,N_13688,N_13173);
nor U14211 (N_14211,N_13447,N_13546);
nor U14212 (N_14212,N_13448,N_13200);
xor U14213 (N_14213,N_13822,N_13418);
and U14214 (N_14214,N_13201,N_13374);
xnor U14215 (N_14215,N_13466,N_13128);
nor U14216 (N_14216,N_13021,N_13901);
xor U14217 (N_14217,N_13417,N_13263);
nor U14218 (N_14218,N_13504,N_13945);
nor U14219 (N_14219,N_13903,N_13424);
xor U14220 (N_14220,N_13052,N_13471);
nand U14221 (N_14221,N_13240,N_13896);
xor U14222 (N_14222,N_13833,N_13380);
nand U14223 (N_14223,N_13916,N_13506);
or U14224 (N_14224,N_13304,N_13034);
and U14225 (N_14225,N_13342,N_13687);
and U14226 (N_14226,N_13078,N_13838);
and U14227 (N_14227,N_13463,N_13254);
nor U14228 (N_14228,N_13059,N_13176);
nand U14229 (N_14229,N_13752,N_13410);
xnor U14230 (N_14230,N_13521,N_13354);
or U14231 (N_14231,N_13793,N_13644);
nor U14232 (N_14232,N_13818,N_13343);
and U14233 (N_14233,N_13551,N_13715);
nor U14234 (N_14234,N_13738,N_13847);
and U14235 (N_14235,N_13472,N_13661);
nand U14236 (N_14236,N_13296,N_13298);
nor U14237 (N_14237,N_13718,N_13109);
or U14238 (N_14238,N_13442,N_13800);
xnor U14239 (N_14239,N_13458,N_13888);
nor U14240 (N_14240,N_13131,N_13362);
or U14241 (N_14241,N_13523,N_13428);
or U14242 (N_14242,N_13474,N_13657);
and U14243 (N_14243,N_13531,N_13355);
xor U14244 (N_14244,N_13120,N_13614);
nor U14245 (N_14245,N_13451,N_13264);
nand U14246 (N_14246,N_13184,N_13806);
nor U14247 (N_14247,N_13900,N_13843);
or U14248 (N_14248,N_13241,N_13575);
or U14249 (N_14249,N_13411,N_13673);
nor U14250 (N_14250,N_13111,N_13337);
and U14251 (N_14251,N_13133,N_13127);
nand U14252 (N_14252,N_13597,N_13009);
or U14253 (N_14253,N_13679,N_13199);
and U14254 (N_14254,N_13045,N_13163);
xnor U14255 (N_14255,N_13709,N_13306);
and U14256 (N_14256,N_13748,N_13549);
xor U14257 (N_14257,N_13063,N_13781);
nand U14258 (N_14258,N_13155,N_13443);
nor U14259 (N_14259,N_13867,N_13140);
nand U14260 (N_14260,N_13475,N_13671);
nand U14261 (N_14261,N_13962,N_13347);
nor U14262 (N_14262,N_13948,N_13194);
nand U14263 (N_14263,N_13558,N_13907);
or U14264 (N_14264,N_13775,N_13520);
or U14265 (N_14265,N_13654,N_13588);
and U14266 (N_14266,N_13181,N_13554);
xnor U14267 (N_14267,N_13482,N_13438);
or U14268 (N_14268,N_13352,N_13543);
nor U14269 (N_14269,N_13439,N_13267);
or U14270 (N_14270,N_13810,N_13723);
nor U14271 (N_14271,N_13629,N_13501);
and U14272 (N_14272,N_13790,N_13197);
nand U14273 (N_14273,N_13787,N_13942);
or U14274 (N_14274,N_13168,N_13288);
nand U14275 (N_14275,N_13946,N_13667);
or U14276 (N_14276,N_13457,N_13995);
xor U14277 (N_14277,N_13057,N_13934);
xnor U14278 (N_14278,N_13124,N_13110);
nor U14279 (N_14279,N_13495,N_13326);
or U14280 (N_14280,N_13259,N_13992);
xor U14281 (N_14281,N_13817,N_13681);
or U14282 (N_14282,N_13132,N_13074);
xor U14283 (N_14283,N_13479,N_13512);
or U14284 (N_14284,N_13030,N_13429);
and U14285 (N_14285,N_13915,N_13257);
nor U14286 (N_14286,N_13537,N_13893);
or U14287 (N_14287,N_13371,N_13771);
and U14288 (N_14288,N_13704,N_13522);
and U14289 (N_14289,N_13079,N_13974);
xnor U14290 (N_14290,N_13351,N_13565);
nand U14291 (N_14291,N_13792,N_13786);
and U14292 (N_14292,N_13932,N_13566);
and U14293 (N_14293,N_13011,N_13105);
and U14294 (N_14294,N_13875,N_13073);
xor U14295 (N_14295,N_13641,N_13878);
and U14296 (N_14296,N_13135,N_13437);
or U14297 (N_14297,N_13689,N_13094);
nand U14298 (N_14298,N_13789,N_13130);
nand U14299 (N_14299,N_13751,N_13456);
or U14300 (N_14300,N_13842,N_13119);
or U14301 (N_14301,N_13452,N_13215);
or U14302 (N_14302,N_13801,N_13547);
xnor U14303 (N_14303,N_13845,N_13938);
nand U14304 (N_14304,N_13767,N_13741);
or U14305 (N_14305,N_13552,N_13214);
and U14306 (N_14306,N_13854,N_13139);
or U14307 (N_14307,N_13324,N_13067);
nor U14308 (N_14308,N_13621,N_13121);
and U14309 (N_14309,N_13198,N_13177);
and U14310 (N_14310,N_13877,N_13969);
or U14311 (N_14311,N_13313,N_13364);
and U14312 (N_14312,N_13196,N_13216);
and U14313 (N_14313,N_13726,N_13563);
nor U14314 (N_14314,N_13528,N_13834);
xnor U14315 (N_14315,N_13016,N_13419);
nand U14316 (N_14316,N_13713,N_13293);
or U14317 (N_14317,N_13777,N_13056);
or U14318 (N_14318,N_13497,N_13620);
and U14319 (N_14319,N_13253,N_13676);
xor U14320 (N_14320,N_13169,N_13227);
or U14321 (N_14321,N_13383,N_13491);
nor U14322 (N_14322,N_13396,N_13432);
nand U14323 (N_14323,N_13764,N_13490);
nor U14324 (N_14324,N_13053,N_13076);
nand U14325 (N_14325,N_13084,N_13312);
and U14326 (N_14326,N_13933,N_13095);
nor U14327 (N_14327,N_13980,N_13720);
xor U14328 (N_14328,N_13488,N_13064);
nor U14329 (N_14329,N_13143,N_13421);
nor U14330 (N_14330,N_13508,N_13887);
or U14331 (N_14331,N_13739,N_13024);
nand U14332 (N_14332,N_13556,N_13096);
nand U14333 (N_14333,N_13243,N_13630);
xor U14334 (N_14334,N_13664,N_13917);
nand U14335 (N_14335,N_13256,N_13162);
or U14336 (N_14336,N_13891,N_13949);
and U14337 (N_14337,N_13890,N_13191);
and U14338 (N_14338,N_13659,N_13136);
nor U14339 (N_14339,N_13368,N_13981);
and U14340 (N_14340,N_13517,N_13302);
and U14341 (N_14341,N_13037,N_13595);
xor U14342 (N_14342,N_13811,N_13975);
xor U14343 (N_14343,N_13553,N_13742);
or U14344 (N_14344,N_13964,N_13740);
nor U14345 (N_14345,N_13736,N_13384);
nor U14346 (N_14346,N_13952,N_13378);
xnor U14347 (N_14347,N_13300,N_13206);
nor U14348 (N_14348,N_13779,N_13824);
nand U14349 (N_14349,N_13569,N_13470);
nand U14350 (N_14350,N_13242,N_13100);
nand U14351 (N_14351,N_13208,N_13433);
or U14352 (N_14352,N_13931,N_13601);
and U14353 (N_14353,N_13369,N_13733);
nand U14354 (N_14354,N_13081,N_13538);
nor U14355 (N_14355,N_13379,N_13344);
xnor U14356 (N_14356,N_13529,N_13183);
or U14357 (N_14357,N_13526,N_13481);
xor U14358 (N_14358,N_13593,N_13881);
or U14359 (N_14359,N_13035,N_13971);
xnor U14360 (N_14360,N_13018,N_13768);
or U14361 (N_14361,N_13391,N_13650);
nor U14362 (N_14362,N_13747,N_13393);
xor U14363 (N_14363,N_13578,N_13936);
xor U14364 (N_14364,N_13339,N_13299);
and U14365 (N_14365,N_13912,N_13743);
and U14366 (N_14366,N_13823,N_13232);
and U14367 (N_14367,N_13087,N_13909);
and U14368 (N_14368,N_13640,N_13403);
nand U14369 (N_14369,N_13043,N_13061);
nor U14370 (N_14370,N_13318,N_13572);
xnor U14371 (N_14371,N_13831,N_13498);
and U14372 (N_14372,N_13761,N_13624);
nor U14373 (N_14373,N_13049,N_13603);
nand U14374 (N_14374,N_13866,N_13407);
xor U14375 (N_14375,N_13716,N_13965);
xor U14376 (N_14376,N_13876,N_13334);
or U14377 (N_14377,N_13258,N_13158);
and U14378 (N_14378,N_13335,N_13252);
or U14379 (N_14379,N_13072,N_13085);
nand U14380 (N_14380,N_13058,N_13573);
nor U14381 (N_14381,N_13695,N_13939);
nor U14382 (N_14382,N_13922,N_13570);
nor U14383 (N_14383,N_13755,N_13117);
and U14384 (N_14384,N_13192,N_13653);
or U14385 (N_14385,N_13022,N_13798);
nor U14386 (N_14386,N_13107,N_13023);
or U14387 (N_14387,N_13203,N_13055);
xor U14388 (N_14388,N_13859,N_13157);
and U14389 (N_14389,N_13821,N_13060);
or U14390 (N_14390,N_13505,N_13562);
nor U14391 (N_14391,N_13340,N_13580);
nor U14392 (N_14392,N_13229,N_13998);
and U14393 (N_14393,N_13782,N_13735);
nor U14394 (N_14394,N_13678,N_13927);
nor U14395 (N_14395,N_13808,N_13613);
or U14396 (N_14396,N_13675,N_13530);
or U14397 (N_14397,N_13492,N_13873);
nor U14398 (N_14398,N_13647,N_13564);
nand U14399 (N_14399,N_13886,N_13976);
nor U14400 (N_14400,N_13205,N_13211);
nor U14401 (N_14401,N_13436,N_13104);
and U14402 (N_14402,N_13576,N_13307);
or U14403 (N_14403,N_13799,N_13178);
or U14404 (N_14404,N_13250,N_13928);
or U14405 (N_14405,N_13091,N_13700);
nor U14406 (N_14406,N_13921,N_13559);
nor U14407 (N_14407,N_13469,N_13500);
nor U14408 (N_14408,N_13955,N_13483);
nor U14409 (N_14409,N_13068,N_13174);
xor U14410 (N_14410,N_13765,N_13017);
or U14411 (N_14411,N_13006,N_13099);
nor U14412 (N_14412,N_13172,N_13077);
nor U14413 (N_14413,N_13513,N_13814);
xnor U14414 (N_14414,N_13923,N_13805);
or U14415 (N_14415,N_13905,N_13345);
and U14416 (N_14416,N_13236,N_13348);
and U14417 (N_14417,N_13865,N_13994);
xor U14418 (N_14418,N_13684,N_13769);
or U14419 (N_14419,N_13455,N_13336);
nor U14420 (N_14420,N_13493,N_13555);
or U14421 (N_14421,N_13561,N_13929);
nand U14422 (N_14422,N_13589,N_13682);
or U14423 (N_14423,N_13465,N_13389);
or U14424 (N_14424,N_13218,N_13360);
nand U14425 (N_14425,N_13685,N_13430);
and U14426 (N_14426,N_13453,N_13152);
nor U14427 (N_14427,N_13852,N_13631);
nand U14428 (N_14428,N_13397,N_13602);
nand U14429 (N_14429,N_13728,N_13175);
xor U14430 (N_14430,N_13185,N_13123);
and U14431 (N_14431,N_13062,N_13950);
nand U14432 (N_14432,N_13093,N_13204);
nor U14433 (N_14433,N_13387,N_13841);
or U14434 (N_14434,N_13757,N_13908);
xor U14435 (N_14435,N_13235,N_13289);
or U14436 (N_14436,N_13658,N_13967);
nor U14437 (N_14437,N_13714,N_13514);
or U14438 (N_14438,N_13002,N_13722);
or U14439 (N_14439,N_13646,N_13361);
xor U14440 (N_14440,N_13760,N_13033);
nand U14441 (N_14441,N_13745,N_13050);
nand U14442 (N_14442,N_13262,N_13358);
and U14443 (N_14443,N_13633,N_13270);
nor U14444 (N_14444,N_13125,N_13233);
nor U14445 (N_14445,N_13422,N_13141);
xor U14446 (N_14446,N_13809,N_13273);
nand U14447 (N_14447,N_13772,N_13113);
or U14448 (N_14448,N_13032,N_13285);
and U14449 (N_14449,N_13586,N_13406);
xor U14450 (N_14450,N_13897,N_13012);
nor U14451 (N_14451,N_13000,N_13097);
xor U14452 (N_14452,N_13086,N_13041);
nand U14453 (N_14453,N_13193,N_13382);
or U14454 (N_14454,N_13904,N_13271);
nand U14455 (N_14455,N_13150,N_13164);
nor U14456 (N_14456,N_13323,N_13414);
or U14457 (N_14457,N_13331,N_13753);
nand U14458 (N_14458,N_13245,N_13632);
and U14459 (N_14459,N_13699,N_13116);
xor U14460 (N_14460,N_13219,N_13648);
or U14461 (N_14461,N_13349,N_13311);
nand U14462 (N_14462,N_13763,N_13788);
or U14463 (N_14463,N_13683,N_13287);
nand U14464 (N_14464,N_13548,N_13402);
or U14465 (N_14465,N_13977,N_13696);
and U14466 (N_14466,N_13605,N_13796);
xnor U14467 (N_14467,N_13284,N_13985);
and U14468 (N_14468,N_13265,N_13317);
nor U14469 (N_14469,N_13690,N_13958);
xor U14470 (N_14470,N_13680,N_13898);
nand U14471 (N_14471,N_13794,N_13966);
and U14472 (N_14472,N_13047,N_13960);
xnor U14473 (N_14473,N_13749,N_13773);
nand U14474 (N_14474,N_13724,N_13161);
xor U14475 (N_14475,N_13333,N_13542);
or U14476 (N_14476,N_13188,N_13507);
xor U14477 (N_14477,N_13524,N_13187);
or U14478 (N_14478,N_13122,N_13830);
or U14479 (N_14479,N_13370,N_13294);
and U14480 (N_14480,N_13375,N_13332);
and U14481 (N_14481,N_13691,N_13013);
nor U14482 (N_14482,N_13290,N_13550);
nand U14483 (N_14483,N_13409,N_13982);
xor U14484 (N_14484,N_13545,N_13408);
xor U14485 (N_14485,N_13744,N_13004);
or U14486 (N_14486,N_13171,N_13385);
or U14487 (N_14487,N_13656,N_13727);
nand U14488 (N_14488,N_13230,N_13190);
nor U14489 (N_14489,N_13126,N_13870);
nand U14490 (N_14490,N_13940,N_13567);
and U14491 (N_14491,N_13725,N_13291);
nor U14492 (N_14492,N_13848,N_13101);
xnor U14493 (N_14493,N_13329,N_13462);
nor U14494 (N_14494,N_13478,N_13628);
or U14495 (N_14495,N_13212,N_13473);
nor U14496 (N_14496,N_13527,N_13098);
nor U14497 (N_14497,N_13868,N_13372);
and U14498 (N_14498,N_13712,N_13642);
xnor U14499 (N_14499,N_13019,N_13819);
and U14500 (N_14500,N_13226,N_13786);
nor U14501 (N_14501,N_13913,N_13255);
nor U14502 (N_14502,N_13967,N_13718);
xor U14503 (N_14503,N_13004,N_13669);
nor U14504 (N_14504,N_13763,N_13657);
nand U14505 (N_14505,N_13801,N_13852);
or U14506 (N_14506,N_13769,N_13995);
or U14507 (N_14507,N_13578,N_13260);
nand U14508 (N_14508,N_13102,N_13240);
nand U14509 (N_14509,N_13837,N_13791);
xor U14510 (N_14510,N_13817,N_13452);
and U14511 (N_14511,N_13021,N_13321);
and U14512 (N_14512,N_13243,N_13118);
xor U14513 (N_14513,N_13650,N_13009);
nand U14514 (N_14514,N_13610,N_13374);
xor U14515 (N_14515,N_13690,N_13758);
or U14516 (N_14516,N_13914,N_13417);
nand U14517 (N_14517,N_13225,N_13997);
nand U14518 (N_14518,N_13894,N_13403);
xor U14519 (N_14519,N_13958,N_13938);
nand U14520 (N_14520,N_13091,N_13149);
xnor U14521 (N_14521,N_13428,N_13578);
xnor U14522 (N_14522,N_13952,N_13775);
or U14523 (N_14523,N_13133,N_13280);
and U14524 (N_14524,N_13034,N_13809);
nor U14525 (N_14525,N_13084,N_13025);
nor U14526 (N_14526,N_13659,N_13450);
nor U14527 (N_14527,N_13326,N_13892);
nor U14528 (N_14528,N_13359,N_13270);
nor U14529 (N_14529,N_13673,N_13970);
and U14530 (N_14530,N_13223,N_13357);
nor U14531 (N_14531,N_13194,N_13006);
xor U14532 (N_14532,N_13442,N_13703);
nor U14533 (N_14533,N_13706,N_13138);
or U14534 (N_14534,N_13486,N_13524);
or U14535 (N_14535,N_13442,N_13241);
nand U14536 (N_14536,N_13269,N_13065);
nand U14537 (N_14537,N_13774,N_13961);
xor U14538 (N_14538,N_13934,N_13074);
xor U14539 (N_14539,N_13096,N_13187);
and U14540 (N_14540,N_13822,N_13068);
nand U14541 (N_14541,N_13680,N_13929);
nand U14542 (N_14542,N_13126,N_13910);
and U14543 (N_14543,N_13184,N_13240);
or U14544 (N_14544,N_13219,N_13309);
nor U14545 (N_14545,N_13274,N_13326);
and U14546 (N_14546,N_13447,N_13313);
nand U14547 (N_14547,N_13033,N_13386);
or U14548 (N_14548,N_13039,N_13393);
xor U14549 (N_14549,N_13909,N_13478);
and U14550 (N_14550,N_13854,N_13835);
or U14551 (N_14551,N_13558,N_13626);
or U14552 (N_14552,N_13215,N_13817);
nor U14553 (N_14553,N_13901,N_13744);
nor U14554 (N_14554,N_13462,N_13144);
xor U14555 (N_14555,N_13397,N_13080);
and U14556 (N_14556,N_13851,N_13597);
nor U14557 (N_14557,N_13666,N_13177);
nand U14558 (N_14558,N_13072,N_13027);
nor U14559 (N_14559,N_13945,N_13709);
nand U14560 (N_14560,N_13325,N_13905);
and U14561 (N_14561,N_13809,N_13357);
nor U14562 (N_14562,N_13319,N_13849);
or U14563 (N_14563,N_13286,N_13542);
nand U14564 (N_14564,N_13346,N_13385);
nor U14565 (N_14565,N_13149,N_13362);
xnor U14566 (N_14566,N_13800,N_13313);
or U14567 (N_14567,N_13239,N_13989);
or U14568 (N_14568,N_13178,N_13894);
nor U14569 (N_14569,N_13082,N_13466);
or U14570 (N_14570,N_13973,N_13055);
xnor U14571 (N_14571,N_13088,N_13380);
and U14572 (N_14572,N_13218,N_13511);
xnor U14573 (N_14573,N_13223,N_13124);
and U14574 (N_14574,N_13168,N_13012);
and U14575 (N_14575,N_13459,N_13564);
nand U14576 (N_14576,N_13284,N_13134);
nand U14577 (N_14577,N_13561,N_13133);
or U14578 (N_14578,N_13019,N_13301);
and U14579 (N_14579,N_13960,N_13034);
nor U14580 (N_14580,N_13565,N_13380);
or U14581 (N_14581,N_13240,N_13945);
nor U14582 (N_14582,N_13055,N_13905);
nand U14583 (N_14583,N_13537,N_13393);
nor U14584 (N_14584,N_13834,N_13465);
and U14585 (N_14585,N_13865,N_13016);
nand U14586 (N_14586,N_13859,N_13466);
or U14587 (N_14587,N_13713,N_13697);
and U14588 (N_14588,N_13940,N_13507);
xor U14589 (N_14589,N_13019,N_13743);
nor U14590 (N_14590,N_13550,N_13680);
xnor U14591 (N_14591,N_13451,N_13448);
and U14592 (N_14592,N_13829,N_13568);
or U14593 (N_14593,N_13235,N_13157);
nand U14594 (N_14594,N_13536,N_13938);
and U14595 (N_14595,N_13331,N_13116);
and U14596 (N_14596,N_13733,N_13897);
or U14597 (N_14597,N_13661,N_13174);
xnor U14598 (N_14598,N_13868,N_13869);
or U14599 (N_14599,N_13555,N_13670);
nand U14600 (N_14600,N_13401,N_13202);
and U14601 (N_14601,N_13707,N_13044);
nor U14602 (N_14602,N_13349,N_13785);
and U14603 (N_14603,N_13245,N_13258);
nor U14604 (N_14604,N_13755,N_13747);
nor U14605 (N_14605,N_13836,N_13802);
and U14606 (N_14606,N_13340,N_13327);
nand U14607 (N_14607,N_13230,N_13015);
or U14608 (N_14608,N_13512,N_13228);
and U14609 (N_14609,N_13274,N_13435);
nor U14610 (N_14610,N_13323,N_13190);
nand U14611 (N_14611,N_13256,N_13013);
and U14612 (N_14612,N_13573,N_13685);
nand U14613 (N_14613,N_13375,N_13899);
and U14614 (N_14614,N_13196,N_13504);
or U14615 (N_14615,N_13481,N_13206);
and U14616 (N_14616,N_13724,N_13058);
nor U14617 (N_14617,N_13796,N_13014);
nor U14618 (N_14618,N_13902,N_13930);
or U14619 (N_14619,N_13620,N_13004);
nand U14620 (N_14620,N_13384,N_13864);
or U14621 (N_14621,N_13205,N_13650);
nor U14622 (N_14622,N_13199,N_13951);
nand U14623 (N_14623,N_13996,N_13753);
xnor U14624 (N_14624,N_13662,N_13703);
nor U14625 (N_14625,N_13966,N_13214);
and U14626 (N_14626,N_13032,N_13872);
nor U14627 (N_14627,N_13663,N_13883);
xor U14628 (N_14628,N_13106,N_13647);
nor U14629 (N_14629,N_13995,N_13646);
and U14630 (N_14630,N_13743,N_13717);
nand U14631 (N_14631,N_13966,N_13351);
and U14632 (N_14632,N_13192,N_13585);
or U14633 (N_14633,N_13206,N_13716);
xor U14634 (N_14634,N_13919,N_13215);
nand U14635 (N_14635,N_13407,N_13331);
or U14636 (N_14636,N_13777,N_13662);
nand U14637 (N_14637,N_13370,N_13584);
nand U14638 (N_14638,N_13947,N_13651);
nand U14639 (N_14639,N_13078,N_13640);
or U14640 (N_14640,N_13584,N_13374);
nor U14641 (N_14641,N_13118,N_13211);
or U14642 (N_14642,N_13917,N_13000);
nand U14643 (N_14643,N_13484,N_13242);
and U14644 (N_14644,N_13312,N_13631);
and U14645 (N_14645,N_13273,N_13708);
nor U14646 (N_14646,N_13035,N_13899);
and U14647 (N_14647,N_13569,N_13800);
nor U14648 (N_14648,N_13102,N_13433);
xor U14649 (N_14649,N_13866,N_13780);
nor U14650 (N_14650,N_13138,N_13643);
nand U14651 (N_14651,N_13400,N_13436);
and U14652 (N_14652,N_13917,N_13261);
nor U14653 (N_14653,N_13654,N_13394);
xor U14654 (N_14654,N_13147,N_13885);
or U14655 (N_14655,N_13895,N_13047);
nor U14656 (N_14656,N_13368,N_13375);
or U14657 (N_14657,N_13805,N_13305);
and U14658 (N_14658,N_13943,N_13367);
xor U14659 (N_14659,N_13189,N_13259);
nor U14660 (N_14660,N_13723,N_13560);
nand U14661 (N_14661,N_13042,N_13665);
xor U14662 (N_14662,N_13877,N_13845);
or U14663 (N_14663,N_13589,N_13782);
nand U14664 (N_14664,N_13976,N_13336);
nor U14665 (N_14665,N_13127,N_13583);
nand U14666 (N_14666,N_13075,N_13594);
or U14667 (N_14667,N_13841,N_13737);
nor U14668 (N_14668,N_13885,N_13537);
nor U14669 (N_14669,N_13891,N_13841);
nand U14670 (N_14670,N_13377,N_13576);
nand U14671 (N_14671,N_13955,N_13243);
nand U14672 (N_14672,N_13398,N_13627);
nor U14673 (N_14673,N_13543,N_13786);
nand U14674 (N_14674,N_13169,N_13505);
xor U14675 (N_14675,N_13854,N_13617);
or U14676 (N_14676,N_13318,N_13074);
or U14677 (N_14677,N_13684,N_13304);
xor U14678 (N_14678,N_13137,N_13771);
nand U14679 (N_14679,N_13096,N_13035);
nand U14680 (N_14680,N_13361,N_13025);
xor U14681 (N_14681,N_13941,N_13943);
and U14682 (N_14682,N_13133,N_13251);
nor U14683 (N_14683,N_13457,N_13120);
nor U14684 (N_14684,N_13920,N_13604);
or U14685 (N_14685,N_13170,N_13846);
or U14686 (N_14686,N_13596,N_13434);
nor U14687 (N_14687,N_13451,N_13491);
and U14688 (N_14688,N_13733,N_13964);
nor U14689 (N_14689,N_13861,N_13565);
nor U14690 (N_14690,N_13114,N_13960);
and U14691 (N_14691,N_13618,N_13569);
nand U14692 (N_14692,N_13043,N_13045);
nand U14693 (N_14693,N_13491,N_13942);
nand U14694 (N_14694,N_13878,N_13357);
xnor U14695 (N_14695,N_13406,N_13199);
or U14696 (N_14696,N_13729,N_13857);
nand U14697 (N_14697,N_13983,N_13567);
nor U14698 (N_14698,N_13246,N_13854);
and U14699 (N_14699,N_13465,N_13443);
or U14700 (N_14700,N_13674,N_13503);
nand U14701 (N_14701,N_13173,N_13652);
nor U14702 (N_14702,N_13131,N_13134);
or U14703 (N_14703,N_13107,N_13167);
xnor U14704 (N_14704,N_13088,N_13255);
nor U14705 (N_14705,N_13816,N_13960);
xnor U14706 (N_14706,N_13819,N_13233);
nor U14707 (N_14707,N_13536,N_13837);
xnor U14708 (N_14708,N_13589,N_13260);
nor U14709 (N_14709,N_13746,N_13454);
nor U14710 (N_14710,N_13789,N_13834);
xor U14711 (N_14711,N_13459,N_13543);
xnor U14712 (N_14712,N_13225,N_13684);
xnor U14713 (N_14713,N_13807,N_13866);
or U14714 (N_14714,N_13978,N_13052);
nor U14715 (N_14715,N_13564,N_13576);
xnor U14716 (N_14716,N_13517,N_13278);
nand U14717 (N_14717,N_13498,N_13355);
nand U14718 (N_14718,N_13726,N_13767);
nor U14719 (N_14719,N_13334,N_13611);
nand U14720 (N_14720,N_13821,N_13562);
or U14721 (N_14721,N_13292,N_13075);
nor U14722 (N_14722,N_13177,N_13827);
or U14723 (N_14723,N_13821,N_13995);
nor U14724 (N_14724,N_13054,N_13400);
xnor U14725 (N_14725,N_13977,N_13743);
xor U14726 (N_14726,N_13523,N_13928);
xnor U14727 (N_14727,N_13882,N_13964);
and U14728 (N_14728,N_13177,N_13737);
xor U14729 (N_14729,N_13863,N_13670);
or U14730 (N_14730,N_13404,N_13377);
xor U14731 (N_14731,N_13234,N_13238);
nor U14732 (N_14732,N_13942,N_13259);
and U14733 (N_14733,N_13006,N_13005);
nand U14734 (N_14734,N_13843,N_13171);
xnor U14735 (N_14735,N_13219,N_13255);
nand U14736 (N_14736,N_13721,N_13976);
xnor U14737 (N_14737,N_13816,N_13439);
nand U14738 (N_14738,N_13799,N_13643);
nor U14739 (N_14739,N_13143,N_13293);
nor U14740 (N_14740,N_13967,N_13905);
nand U14741 (N_14741,N_13848,N_13195);
nor U14742 (N_14742,N_13176,N_13752);
nor U14743 (N_14743,N_13118,N_13483);
and U14744 (N_14744,N_13402,N_13651);
xor U14745 (N_14745,N_13658,N_13155);
xor U14746 (N_14746,N_13961,N_13294);
nor U14747 (N_14747,N_13300,N_13998);
and U14748 (N_14748,N_13131,N_13167);
and U14749 (N_14749,N_13263,N_13146);
nand U14750 (N_14750,N_13088,N_13584);
nor U14751 (N_14751,N_13120,N_13534);
and U14752 (N_14752,N_13621,N_13131);
nor U14753 (N_14753,N_13781,N_13169);
nor U14754 (N_14754,N_13430,N_13842);
nand U14755 (N_14755,N_13207,N_13131);
and U14756 (N_14756,N_13034,N_13322);
xnor U14757 (N_14757,N_13917,N_13671);
nand U14758 (N_14758,N_13416,N_13089);
xor U14759 (N_14759,N_13365,N_13759);
nand U14760 (N_14760,N_13023,N_13425);
nand U14761 (N_14761,N_13531,N_13614);
and U14762 (N_14762,N_13319,N_13136);
nand U14763 (N_14763,N_13740,N_13488);
nand U14764 (N_14764,N_13544,N_13449);
xnor U14765 (N_14765,N_13704,N_13218);
nand U14766 (N_14766,N_13321,N_13098);
or U14767 (N_14767,N_13035,N_13252);
and U14768 (N_14768,N_13724,N_13354);
xnor U14769 (N_14769,N_13586,N_13984);
xor U14770 (N_14770,N_13046,N_13158);
or U14771 (N_14771,N_13093,N_13500);
xnor U14772 (N_14772,N_13013,N_13676);
xnor U14773 (N_14773,N_13837,N_13652);
nor U14774 (N_14774,N_13455,N_13289);
and U14775 (N_14775,N_13430,N_13017);
nand U14776 (N_14776,N_13578,N_13037);
or U14777 (N_14777,N_13831,N_13178);
nand U14778 (N_14778,N_13780,N_13694);
nand U14779 (N_14779,N_13384,N_13684);
and U14780 (N_14780,N_13846,N_13476);
nor U14781 (N_14781,N_13687,N_13604);
or U14782 (N_14782,N_13466,N_13761);
or U14783 (N_14783,N_13817,N_13290);
or U14784 (N_14784,N_13690,N_13488);
or U14785 (N_14785,N_13266,N_13161);
and U14786 (N_14786,N_13480,N_13544);
xor U14787 (N_14787,N_13979,N_13297);
or U14788 (N_14788,N_13872,N_13801);
and U14789 (N_14789,N_13354,N_13559);
nand U14790 (N_14790,N_13786,N_13824);
nor U14791 (N_14791,N_13893,N_13593);
and U14792 (N_14792,N_13177,N_13908);
nand U14793 (N_14793,N_13469,N_13205);
nor U14794 (N_14794,N_13623,N_13841);
nand U14795 (N_14795,N_13799,N_13849);
nor U14796 (N_14796,N_13509,N_13677);
xor U14797 (N_14797,N_13922,N_13981);
nor U14798 (N_14798,N_13455,N_13500);
xor U14799 (N_14799,N_13473,N_13918);
or U14800 (N_14800,N_13062,N_13265);
xor U14801 (N_14801,N_13882,N_13640);
or U14802 (N_14802,N_13841,N_13810);
xor U14803 (N_14803,N_13859,N_13048);
or U14804 (N_14804,N_13674,N_13049);
nor U14805 (N_14805,N_13662,N_13737);
and U14806 (N_14806,N_13265,N_13954);
and U14807 (N_14807,N_13825,N_13576);
nand U14808 (N_14808,N_13553,N_13131);
or U14809 (N_14809,N_13737,N_13462);
xor U14810 (N_14810,N_13278,N_13434);
nand U14811 (N_14811,N_13605,N_13753);
nand U14812 (N_14812,N_13711,N_13088);
and U14813 (N_14813,N_13135,N_13423);
nor U14814 (N_14814,N_13699,N_13309);
xor U14815 (N_14815,N_13473,N_13802);
and U14816 (N_14816,N_13846,N_13579);
nor U14817 (N_14817,N_13803,N_13818);
and U14818 (N_14818,N_13980,N_13886);
nand U14819 (N_14819,N_13832,N_13435);
and U14820 (N_14820,N_13582,N_13335);
or U14821 (N_14821,N_13030,N_13665);
or U14822 (N_14822,N_13013,N_13129);
nand U14823 (N_14823,N_13698,N_13240);
or U14824 (N_14824,N_13977,N_13594);
nand U14825 (N_14825,N_13382,N_13347);
or U14826 (N_14826,N_13897,N_13118);
or U14827 (N_14827,N_13587,N_13538);
nand U14828 (N_14828,N_13071,N_13165);
and U14829 (N_14829,N_13320,N_13778);
nand U14830 (N_14830,N_13191,N_13146);
nand U14831 (N_14831,N_13662,N_13467);
xor U14832 (N_14832,N_13748,N_13870);
and U14833 (N_14833,N_13450,N_13437);
xor U14834 (N_14834,N_13486,N_13918);
and U14835 (N_14835,N_13840,N_13367);
xor U14836 (N_14836,N_13874,N_13812);
and U14837 (N_14837,N_13442,N_13492);
xor U14838 (N_14838,N_13687,N_13501);
and U14839 (N_14839,N_13722,N_13425);
and U14840 (N_14840,N_13751,N_13348);
and U14841 (N_14841,N_13023,N_13784);
or U14842 (N_14842,N_13618,N_13424);
nand U14843 (N_14843,N_13567,N_13507);
or U14844 (N_14844,N_13141,N_13625);
xor U14845 (N_14845,N_13345,N_13313);
nand U14846 (N_14846,N_13664,N_13135);
nor U14847 (N_14847,N_13325,N_13377);
nor U14848 (N_14848,N_13455,N_13220);
nand U14849 (N_14849,N_13417,N_13402);
xnor U14850 (N_14850,N_13486,N_13896);
or U14851 (N_14851,N_13768,N_13841);
nand U14852 (N_14852,N_13190,N_13338);
xor U14853 (N_14853,N_13410,N_13517);
and U14854 (N_14854,N_13465,N_13797);
nor U14855 (N_14855,N_13522,N_13386);
nor U14856 (N_14856,N_13912,N_13526);
and U14857 (N_14857,N_13603,N_13531);
nand U14858 (N_14858,N_13024,N_13528);
and U14859 (N_14859,N_13658,N_13956);
or U14860 (N_14860,N_13878,N_13167);
and U14861 (N_14861,N_13104,N_13324);
and U14862 (N_14862,N_13889,N_13919);
nand U14863 (N_14863,N_13263,N_13782);
nand U14864 (N_14864,N_13811,N_13088);
xnor U14865 (N_14865,N_13406,N_13978);
nor U14866 (N_14866,N_13247,N_13518);
xnor U14867 (N_14867,N_13645,N_13624);
nand U14868 (N_14868,N_13936,N_13695);
and U14869 (N_14869,N_13166,N_13049);
or U14870 (N_14870,N_13674,N_13689);
and U14871 (N_14871,N_13845,N_13430);
xnor U14872 (N_14872,N_13000,N_13087);
and U14873 (N_14873,N_13439,N_13070);
nand U14874 (N_14874,N_13117,N_13688);
xnor U14875 (N_14875,N_13293,N_13698);
or U14876 (N_14876,N_13191,N_13704);
xnor U14877 (N_14877,N_13191,N_13017);
nand U14878 (N_14878,N_13361,N_13809);
xnor U14879 (N_14879,N_13761,N_13277);
and U14880 (N_14880,N_13408,N_13318);
xnor U14881 (N_14881,N_13053,N_13228);
nor U14882 (N_14882,N_13801,N_13952);
nand U14883 (N_14883,N_13312,N_13639);
or U14884 (N_14884,N_13277,N_13721);
nor U14885 (N_14885,N_13354,N_13467);
or U14886 (N_14886,N_13294,N_13311);
and U14887 (N_14887,N_13690,N_13098);
and U14888 (N_14888,N_13785,N_13540);
nand U14889 (N_14889,N_13531,N_13749);
nand U14890 (N_14890,N_13378,N_13628);
nor U14891 (N_14891,N_13014,N_13961);
xor U14892 (N_14892,N_13354,N_13473);
nor U14893 (N_14893,N_13835,N_13383);
and U14894 (N_14894,N_13324,N_13028);
and U14895 (N_14895,N_13939,N_13930);
and U14896 (N_14896,N_13669,N_13276);
or U14897 (N_14897,N_13761,N_13172);
nand U14898 (N_14898,N_13496,N_13892);
or U14899 (N_14899,N_13071,N_13414);
and U14900 (N_14900,N_13398,N_13497);
nor U14901 (N_14901,N_13717,N_13017);
nand U14902 (N_14902,N_13532,N_13412);
and U14903 (N_14903,N_13781,N_13161);
and U14904 (N_14904,N_13944,N_13123);
or U14905 (N_14905,N_13798,N_13241);
and U14906 (N_14906,N_13023,N_13969);
or U14907 (N_14907,N_13533,N_13163);
xnor U14908 (N_14908,N_13541,N_13372);
nor U14909 (N_14909,N_13826,N_13086);
nor U14910 (N_14910,N_13533,N_13226);
xnor U14911 (N_14911,N_13614,N_13698);
or U14912 (N_14912,N_13513,N_13481);
and U14913 (N_14913,N_13272,N_13169);
nor U14914 (N_14914,N_13952,N_13120);
nor U14915 (N_14915,N_13993,N_13655);
and U14916 (N_14916,N_13970,N_13846);
nor U14917 (N_14917,N_13422,N_13020);
nand U14918 (N_14918,N_13867,N_13693);
xor U14919 (N_14919,N_13150,N_13617);
xnor U14920 (N_14920,N_13547,N_13105);
nor U14921 (N_14921,N_13072,N_13201);
or U14922 (N_14922,N_13222,N_13738);
or U14923 (N_14923,N_13159,N_13765);
or U14924 (N_14924,N_13815,N_13078);
and U14925 (N_14925,N_13416,N_13582);
xnor U14926 (N_14926,N_13968,N_13627);
and U14927 (N_14927,N_13510,N_13136);
xor U14928 (N_14928,N_13469,N_13544);
xnor U14929 (N_14929,N_13402,N_13515);
and U14930 (N_14930,N_13293,N_13204);
xnor U14931 (N_14931,N_13276,N_13899);
nor U14932 (N_14932,N_13288,N_13381);
nand U14933 (N_14933,N_13144,N_13324);
xnor U14934 (N_14934,N_13125,N_13739);
and U14935 (N_14935,N_13586,N_13778);
nor U14936 (N_14936,N_13921,N_13389);
xnor U14937 (N_14937,N_13894,N_13069);
or U14938 (N_14938,N_13500,N_13578);
xnor U14939 (N_14939,N_13524,N_13994);
xor U14940 (N_14940,N_13341,N_13007);
nor U14941 (N_14941,N_13478,N_13758);
or U14942 (N_14942,N_13775,N_13733);
nand U14943 (N_14943,N_13828,N_13466);
or U14944 (N_14944,N_13536,N_13271);
xnor U14945 (N_14945,N_13573,N_13993);
nand U14946 (N_14946,N_13452,N_13036);
and U14947 (N_14947,N_13919,N_13075);
or U14948 (N_14948,N_13400,N_13514);
xnor U14949 (N_14949,N_13305,N_13596);
nand U14950 (N_14950,N_13113,N_13476);
and U14951 (N_14951,N_13098,N_13065);
or U14952 (N_14952,N_13175,N_13281);
nor U14953 (N_14953,N_13881,N_13358);
and U14954 (N_14954,N_13167,N_13315);
nand U14955 (N_14955,N_13068,N_13745);
xor U14956 (N_14956,N_13803,N_13961);
and U14957 (N_14957,N_13056,N_13769);
and U14958 (N_14958,N_13584,N_13362);
nor U14959 (N_14959,N_13851,N_13983);
nand U14960 (N_14960,N_13121,N_13036);
xor U14961 (N_14961,N_13479,N_13108);
or U14962 (N_14962,N_13290,N_13504);
nand U14963 (N_14963,N_13911,N_13221);
nand U14964 (N_14964,N_13874,N_13064);
nor U14965 (N_14965,N_13086,N_13153);
and U14966 (N_14966,N_13250,N_13545);
nand U14967 (N_14967,N_13237,N_13629);
or U14968 (N_14968,N_13938,N_13763);
xnor U14969 (N_14969,N_13417,N_13528);
and U14970 (N_14970,N_13623,N_13726);
or U14971 (N_14971,N_13244,N_13513);
nand U14972 (N_14972,N_13794,N_13290);
and U14973 (N_14973,N_13887,N_13942);
nand U14974 (N_14974,N_13581,N_13294);
xor U14975 (N_14975,N_13360,N_13402);
xnor U14976 (N_14976,N_13531,N_13124);
or U14977 (N_14977,N_13613,N_13489);
and U14978 (N_14978,N_13256,N_13270);
xnor U14979 (N_14979,N_13016,N_13706);
nor U14980 (N_14980,N_13857,N_13037);
nor U14981 (N_14981,N_13542,N_13871);
xor U14982 (N_14982,N_13140,N_13121);
or U14983 (N_14983,N_13608,N_13387);
or U14984 (N_14984,N_13042,N_13771);
xor U14985 (N_14985,N_13933,N_13693);
nand U14986 (N_14986,N_13317,N_13474);
or U14987 (N_14987,N_13949,N_13321);
nand U14988 (N_14988,N_13210,N_13867);
nand U14989 (N_14989,N_13412,N_13368);
nand U14990 (N_14990,N_13976,N_13497);
and U14991 (N_14991,N_13052,N_13279);
or U14992 (N_14992,N_13798,N_13645);
or U14993 (N_14993,N_13739,N_13597);
and U14994 (N_14994,N_13349,N_13942);
xor U14995 (N_14995,N_13797,N_13731);
and U14996 (N_14996,N_13270,N_13037);
or U14997 (N_14997,N_13161,N_13513);
xnor U14998 (N_14998,N_13954,N_13068);
nand U14999 (N_14999,N_13078,N_13981);
or U15000 (N_15000,N_14233,N_14001);
nand U15001 (N_15001,N_14922,N_14346);
nor U15002 (N_15002,N_14367,N_14109);
nand U15003 (N_15003,N_14643,N_14851);
xnor U15004 (N_15004,N_14297,N_14919);
xnor U15005 (N_15005,N_14280,N_14184);
nand U15006 (N_15006,N_14926,N_14229);
and U15007 (N_15007,N_14528,N_14605);
xor U15008 (N_15008,N_14058,N_14107);
nor U15009 (N_15009,N_14120,N_14847);
nor U15010 (N_15010,N_14440,N_14206);
or U15011 (N_15011,N_14260,N_14086);
nor U15012 (N_15012,N_14145,N_14865);
nand U15013 (N_15013,N_14604,N_14576);
nor U15014 (N_15014,N_14250,N_14942);
nor U15015 (N_15015,N_14842,N_14651);
and U15016 (N_15016,N_14902,N_14007);
xnor U15017 (N_15017,N_14949,N_14684);
nor U15018 (N_15018,N_14728,N_14255);
xor U15019 (N_15019,N_14133,N_14420);
or U15020 (N_15020,N_14337,N_14056);
and U15021 (N_15021,N_14108,N_14426);
nand U15022 (N_15022,N_14670,N_14859);
or U15023 (N_15023,N_14000,N_14144);
or U15024 (N_15024,N_14767,N_14102);
xor U15025 (N_15025,N_14741,N_14492);
nand U15026 (N_15026,N_14074,N_14469);
or U15027 (N_15027,N_14110,N_14873);
and U15028 (N_15028,N_14825,N_14324);
nand U15029 (N_15029,N_14123,N_14616);
and U15030 (N_15030,N_14486,N_14419);
or U15031 (N_15031,N_14603,N_14510);
and U15032 (N_15032,N_14489,N_14882);
and U15033 (N_15033,N_14095,N_14227);
nand U15034 (N_15034,N_14152,N_14397);
or U15035 (N_15035,N_14178,N_14572);
xnor U15036 (N_15036,N_14970,N_14989);
or U15037 (N_15037,N_14965,N_14905);
nor U15038 (N_15038,N_14308,N_14392);
and U15039 (N_15039,N_14092,N_14950);
and U15040 (N_15040,N_14889,N_14550);
xnor U15041 (N_15041,N_14343,N_14774);
xor U15042 (N_15042,N_14691,N_14300);
or U15043 (N_15043,N_14877,N_14017);
xor U15044 (N_15044,N_14656,N_14298);
or U15045 (N_15045,N_14093,N_14739);
and U15046 (N_15046,N_14333,N_14602);
xnor U15047 (N_15047,N_14705,N_14436);
nand U15048 (N_15048,N_14772,N_14499);
nor U15049 (N_15049,N_14228,N_14606);
and U15050 (N_15050,N_14630,N_14833);
nand U15051 (N_15051,N_14968,N_14063);
nor U15052 (N_15052,N_14563,N_14791);
nand U15053 (N_15053,N_14786,N_14209);
xnor U15054 (N_15054,N_14073,N_14854);
nand U15055 (N_15055,N_14004,N_14792);
and U15056 (N_15056,N_14159,N_14773);
and U15057 (N_15057,N_14580,N_14241);
nor U15058 (N_15058,N_14837,N_14646);
nand U15059 (N_15059,N_14676,N_14581);
and U15060 (N_15060,N_14699,N_14849);
xor U15061 (N_15061,N_14824,N_14217);
xor U15062 (N_15062,N_14249,N_14619);
and U15063 (N_15063,N_14078,N_14422);
or U15064 (N_15064,N_14626,N_14655);
or U15065 (N_15065,N_14912,N_14952);
or U15066 (N_15066,N_14679,N_14185);
or U15067 (N_15067,N_14005,N_14597);
and U15068 (N_15068,N_14928,N_14071);
xor U15069 (N_15069,N_14211,N_14666);
nor U15070 (N_15070,N_14946,N_14878);
nor U15071 (N_15071,N_14812,N_14402);
nand U15072 (N_15072,N_14531,N_14053);
xnor U15073 (N_15073,N_14494,N_14041);
nor U15074 (N_15074,N_14628,N_14784);
nor U15075 (N_15075,N_14410,N_14157);
or U15076 (N_15076,N_14521,N_14956);
nor U15077 (N_15077,N_14117,N_14045);
nand U15078 (N_15078,N_14839,N_14681);
or U15079 (N_15079,N_14134,N_14477);
nor U15080 (N_15080,N_14097,N_14051);
or U15081 (N_15081,N_14687,N_14153);
xnor U15082 (N_15082,N_14982,N_14508);
and U15083 (N_15083,N_14328,N_14981);
nor U15084 (N_15084,N_14189,N_14727);
nand U15085 (N_15085,N_14413,N_14932);
nand U15086 (N_15086,N_14316,N_14179);
or U15087 (N_15087,N_14461,N_14176);
or U15088 (N_15088,N_14240,N_14301);
xor U15089 (N_15089,N_14009,N_14829);
or U15090 (N_15090,N_14821,N_14034);
nor U15091 (N_15091,N_14106,N_14718);
xor U15092 (N_15092,N_14857,N_14449);
nand U15093 (N_15093,N_14439,N_14562);
nand U15094 (N_15094,N_14023,N_14969);
or U15095 (N_15095,N_14546,N_14800);
and U15096 (N_15096,N_14814,N_14180);
or U15097 (N_15097,N_14183,N_14174);
and U15098 (N_15098,N_14024,N_14987);
nor U15099 (N_15099,N_14403,N_14822);
and U15100 (N_15100,N_14696,N_14931);
or U15101 (N_15101,N_14043,N_14591);
and U15102 (N_15102,N_14512,N_14471);
nand U15103 (N_15103,N_14277,N_14192);
nand U15104 (N_15104,N_14538,N_14291);
nor U15105 (N_15105,N_14648,N_14458);
and U15106 (N_15106,N_14038,N_14858);
and U15107 (N_15107,N_14483,N_14445);
or U15108 (N_15108,N_14582,N_14526);
or U15109 (N_15109,N_14726,N_14128);
or U15110 (N_15110,N_14985,N_14060);
or U15111 (N_15111,N_14425,N_14997);
nand U15112 (N_15112,N_14374,N_14642);
xnor U15113 (N_15113,N_14904,N_14564);
xor U15114 (N_15114,N_14571,N_14450);
or U15115 (N_15115,N_14763,N_14101);
xnor U15116 (N_15116,N_14488,N_14761);
nand U15117 (N_15117,N_14182,N_14339);
xnor U15118 (N_15118,N_14991,N_14914);
or U15119 (N_15119,N_14811,N_14438);
nand U15120 (N_15120,N_14721,N_14132);
xnor U15121 (N_15121,N_14757,N_14789);
nor U15122 (N_15122,N_14927,N_14378);
xor U15123 (N_15123,N_14365,N_14883);
nor U15124 (N_15124,N_14200,N_14683);
and U15125 (N_15125,N_14527,N_14072);
nor U15126 (N_15126,N_14395,N_14096);
xor U15127 (N_15127,N_14624,N_14223);
nor U15128 (N_15128,N_14370,N_14310);
nand U15129 (N_15129,N_14493,N_14054);
nor U15130 (N_15130,N_14554,N_14972);
or U15131 (N_15131,N_14188,N_14148);
and U15132 (N_15132,N_14411,N_14704);
nor U15133 (N_15133,N_14770,N_14804);
xnor U15134 (N_15134,N_14265,N_14375);
nand U15135 (N_15135,N_14720,N_14087);
xor U15136 (N_15136,N_14371,N_14779);
and U15137 (N_15137,N_14254,N_14639);
and U15138 (N_15138,N_14290,N_14390);
and U15139 (N_15139,N_14487,N_14831);
and U15140 (N_15140,N_14161,N_14372);
nor U15141 (N_15141,N_14934,N_14079);
and U15142 (N_15142,N_14717,N_14544);
and U15143 (N_15143,N_14731,N_14957);
nand U15144 (N_15144,N_14091,N_14121);
and U15145 (N_15145,N_14304,N_14611);
xor U15146 (N_15146,N_14443,N_14677);
xnor U15147 (N_15147,N_14903,N_14273);
xnor U15148 (N_15148,N_14583,N_14215);
nand U15149 (N_15149,N_14797,N_14481);
xnor U15150 (N_15150,N_14142,N_14633);
or U15151 (N_15151,N_14787,N_14203);
or U15152 (N_15152,N_14794,N_14088);
nand U15153 (N_15153,N_14131,N_14612);
or U15154 (N_15154,N_14112,N_14940);
nor U15155 (N_15155,N_14175,N_14678);
or U15156 (N_15156,N_14975,N_14896);
xnor U15157 (N_15157,N_14667,N_14027);
xnor U15158 (N_15158,N_14454,N_14547);
nor U15159 (N_15159,N_14751,N_14744);
and U15160 (N_15160,N_14348,N_14040);
xnor U15161 (N_15161,N_14893,N_14688);
or U15162 (N_15162,N_14524,N_14844);
or U15163 (N_15163,N_14979,N_14194);
nand U15164 (N_15164,N_14160,N_14416);
and U15165 (N_15165,N_14986,N_14959);
xnor U15166 (N_15166,N_14542,N_14430);
xor U15167 (N_15167,N_14801,N_14618);
nand U15168 (N_15168,N_14398,N_14532);
or U15169 (N_15169,N_14270,N_14995);
or U15170 (N_15170,N_14682,N_14266);
or U15171 (N_15171,N_14080,N_14267);
nor U15172 (N_15172,N_14823,N_14468);
nor U15173 (N_15173,N_14881,N_14513);
or U15174 (N_15174,N_14860,N_14460);
or U15175 (N_15175,N_14835,N_14988);
nand U15176 (N_15176,N_14937,N_14709);
or U15177 (N_15177,N_14921,N_14737);
xnor U15178 (N_15178,N_14697,N_14548);
xnor U15179 (N_15179,N_14322,N_14447);
xnor U15180 (N_15180,N_14113,N_14875);
nand U15181 (N_15181,N_14361,N_14129);
or U15182 (N_15182,N_14042,N_14783);
nand U15183 (N_15183,N_14627,N_14652);
nand U15184 (N_15184,N_14295,N_14748);
or U15185 (N_15185,N_14243,N_14190);
xnor U15186 (N_15186,N_14465,N_14664);
nand U15187 (N_15187,N_14708,N_14218);
xor U15188 (N_15188,N_14116,N_14723);
and U15189 (N_15189,N_14738,N_14177);
and U15190 (N_15190,N_14929,N_14930);
nand U15191 (N_15191,N_14125,N_14207);
nand U15192 (N_15192,N_14137,N_14022);
nor U15193 (N_15193,N_14868,N_14455);
nand U15194 (N_15194,N_14050,N_14478);
or U15195 (N_15195,N_14208,N_14334);
nand U15196 (N_15196,N_14408,N_14507);
nand U15197 (N_15197,N_14925,N_14246);
nor U15198 (N_15198,N_14235,N_14703);
or U15199 (N_15199,N_14590,N_14650);
or U15200 (N_15200,N_14514,N_14057);
or U15201 (N_15201,N_14360,N_14615);
nor U15202 (N_15202,N_14622,N_14502);
and U15203 (N_15203,N_14669,N_14695);
xnor U15204 (N_15204,N_14067,N_14342);
nand U15205 (N_15205,N_14003,N_14016);
nand U15206 (N_15206,N_14141,N_14589);
xnor U15207 (N_15207,N_14010,N_14675);
nand U15208 (N_15208,N_14895,N_14911);
and U15209 (N_15209,N_14760,N_14944);
nor U15210 (N_15210,N_14358,N_14242);
and U15211 (N_15211,N_14225,N_14115);
or U15212 (N_15212,N_14463,N_14345);
nor U15213 (N_15213,N_14820,N_14421);
xor U15214 (N_15214,N_14433,N_14165);
nand U15215 (N_15215,N_14853,N_14775);
or U15216 (N_15216,N_14568,N_14424);
nand U15217 (N_15217,N_14848,N_14785);
or U15218 (N_15218,N_14156,N_14248);
xor U15219 (N_15219,N_14015,N_14008);
xor U15220 (N_15220,N_14909,N_14535);
and U15221 (N_15221,N_14168,N_14356);
and U15222 (N_15222,N_14620,N_14898);
and U15223 (N_15223,N_14712,N_14505);
xor U15224 (N_15224,N_14745,N_14490);
xor U15225 (N_15225,N_14352,N_14559);
xor U15226 (N_15226,N_14467,N_14068);
xnor U15227 (N_15227,N_14668,N_14754);
nor U15228 (N_15228,N_14807,N_14466);
xnor U15229 (N_15229,N_14694,N_14158);
nand U15230 (N_15230,N_14018,N_14836);
nand U15231 (N_15231,N_14938,N_14557);
and U15232 (N_15232,N_14543,N_14870);
or U15233 (N_15233,N_14258,N_14186);
xor U15234 (N_15234,N_14777,N_14534);
or U15235 (N_15235,N_14351,N_14588);
nor U15236 (N_15236,N_14778,N_14098);
nand U15237 (N_15237,N_14172,N_14198);
or U15238 (N_15238,N_14173,N_14999);
nor U15239 (N_15239,N_14036,N_14296);
and U15240 (N_15240,N_14220,N_14587);
or U15241 (N_15241,N_14282,N_14974);
or U15242 (N_15242,N_14509,N_14996);
nor U15243 (N_15243,N_14379,N_14948);
and U15244 (N_15244,N_14373,N_14955);
nand U15245 (N_15245,N_14788,N_14625);
nor U15246 (N_15246,N_14124,N_14442);
nand U15247 (N_15247,N_14891,N_14560);
nor U15248 (N_15248,N_14354,N_14039);
and U15249 (N_15249,N_14384,N_14272);
nand U15250 (N_15250,N_14081,N_14756);
nand U15251 (N_15251,N_14685,N_14585);
or U15252 (N_15252,N_14867,N_14653);
or U15253 (N_15253,N_14963,N_14163);
or U15254 (N_15254,N_14269,N_14888);
nand U15255 (N_15255,N_14900,N_14874);
nor U15256 (N_15256,N_14019,N_14719);
or U15257 (N_15257,N_14500,N_14226);
nand U15258 (N_15258,N_14317,N_14511);
nor U15259 (N_15259,N_14923,N_14577);
xnor U15260 (N_15260,N_14575,N_14046);
and U15261 (N_15261,N_14257,N_14863);
nor U15262 (N_15262,N_14998,N_14917);
nand U15263 (N_15263,N_14764,N_14555);
xor U15264 (N_15264,N_14154,N_14473);
nor U15265 (N_15265,N_14933,N_14094);
or U15266 (N_15266,N_14558,N_14879);
or U15267 (N_15267,N_14936,N_14472);
or U15268 (N_15268,N_14232,N_14014);
nand U15269 (N_15269,N_14065,N_14283);
nand U15270 (N_15270,N_14945,N_14307);
xor U15271 (N_15271,N_14796,N_14496);
and U15272 (N_15272,N_14729,N_14143);
nor U15273 (N_15273,N_14150,N_14740);
and U15274 (N_15274,N_14274,N_14195);
nor U15275 (N_15275,N_14059,N_14734);
nor U15276 (N_15276,N_14795,N_14765);
and U15277 (N_15277,N_14993,N_14332);
and U15278 (N_15278,N_14075,N_14918);
or U15279 (N_15279,N_14553,N_14644);
nor U15280 (N_15280,N_14234,N_14032);
xor U15281 (N_15281,N_14052,N_14407);
or U15282 (N_15282,N_14247,N_14686);
or U15283 (N_15283,N_14002,N_14139);
or U15284 (N_15284,N_14813,N_14119);
or U15285 (N_15285,N_14498,N_14400);
nor U15286 (N_15286,N_14111,N_14768);
xnor U15287 (N_15287,N_14805,N_14386);
nand U15288 (N_15288,N_14380,N_14924);
or U15289 (N_15289,N_14654,N_14736);
or U15290 (N_15290,N_14710,N_14536);
xnor U15291 (N_15291,N_14147,N_14711);
or U15292 (N_15292,N_14406,N_14517);
and U15293 (N_15293,N_14169,N_14459);
nor U15294 (N_15294,N_14434,N_14230);
and U15295 (N_15295,N_14122,N_14660);
or U15296 (N_15296,N_14830,N_14127);
or U15297 (N_15297,N_14418,N_14749);
nor U15298 (N_15298,N_14244,N_14105);
or U15299 (N_15299,N_14673,N_14181);
and U15300 (N_15300,N_14816,N_14762);
nand U15301 (N_15301,N_14617,N_14325);
or U15302 (N_15302,N_14966,N_14197);
and U15303 (N_15303,N_14485,N_14961);
nand U15304 (N_15304,N_14608,N_14724);
nand U15305 (N_15305,N_14971,N_14126);
or U15306 (N_15306,N_14025,N_14453);
xor U15307 (N_15307,N_14638,N_14850);
nor U15308 (N_15308,N_14916,N_14278);
xor U15309 (N_15309,N_14140,N_14136);
or U15310 (N_15310,N_14394,N_14412);
xor U15311 (N_15311,N_14569,N_14224);
nand U15312 (N_15312,N_14680,N_14170);
nand U15313 (N_15313,N_14329,N_14798);
nor U15314 (N_15314,N_14263,N_14340);
xnor U15315 (N_15315,N_14947,N_14658);
and U15316 (N_15316,N_14806,N_14722);
or U15317 (N_15317,N_14480,N_14114);
or U15318 (N_15318,N_14201,N_14659);
nor U15319 (N_15319,N_14752,N_14992);
nor U15320 (N_15320,N_14323,N_14594);
nor U15321 (N_15321,N_14279,N_14504);
or U15322 (N_15322,N_14497,N_14423);
nor U15323 (N_15323,N_14167,N_14735);
nand U15324 (N_15324,N_14725,N_14271);
nor U15325 (N_15325,N_14586,N_14556);
xnor U15326 (N_15326,N_14579,N_14908);
xor U15327 (N_15327,N_14070,N_14199);
or U15328 (N_15328,N_14613,N_14803);
and U15329 (N_15329,N_14584,N_14164);
and U15330 (N_15330,N_14529,N_14303);
xnor U15331 (N_15331,N_14817,N_14222);
and U15332 (N_15332,N_14456,N_14960);
and U15333 (N_15333,N_14381,N_14506);
xor U15334 (N_15334,N_14663,N_14312);
nand U15335 (N_15335,N_14565,N_14856);
or U15336 (N_15336,N_14049,N_14026);
nand U15337 (N_15337,N_14753,N_14090);
nand U15338 (N_15338,N_14810,N_14252);
and U15339 (N_15339,N_14256,N_14886);
or U15340 (N_15340,N_14843,N_14368);
nand U15341 (N_15341,N_14064,N_14104);
and U15342 (N_15342,N_14657,N_14780);
nand U15343 (N_15343,N_14976,N_14781);
or U15344 (N_15344,N_14713,N_14501);
xnor U15345 (N_15345,N_14747,N_14238);
nor U15346 (N_15346,N_14689,N_14599);
nand U15347 (N_15347,N_14204,N_14636);
or U15348 (N_15348,N_14006,N_14464);
nand U15349 (N_15349,N_14520,N_14021);
and U15350 (N_15350,N_14245,N_14353);
nor U15351 (N_15351,N_14311,N_14047);
and U15352 (N_15352,N_14645,N_14377);
or U15353 (N_15353,N_14819,N_14714);
or U15354 (N_15354,N_14268,N_14389);
nor U15355 (N_15355,N_14827,N_14399);
xnor U15356 (N_15356,N_14790,N_14845);
xnor U15357 (N_15357,N_14330,N_14069);
and U15358 (N_15358,N_14852,N_14941);
nor U15359 (N_15359,N_14428,N_14013);
nor U15360 (N_15360,N_14077,N_14327);
nand U15361 (N_15361,N_14869,N_14294);
or U15362 (N_15362,N_14808,N_14861);
xnor U15363 (N_15363,N_14503,N_14635);
xor U15364 (N_15364,N_14171,N_14907);
nor U15365 (N_15365,N_14799,N_14028);
and U15366 (N_15366,N_14978,N_14321);
and U15367 (N_15367,N_14693,N_14385);
nor U15368 (N_15368,N_14629,N_14405);
xnor U15369 (N_15369,N_14437,N_14221);
or U15370 (N_15370,N_14884,N_14601);
nand U15371 (N_15371,N_14570,N_14484);
or U15372 (N_15372,N_14314,N_14236);
nand U15373 (N_15373,N_14609,N_14980);
and U15374 (N_15374,N_14326,N_14103);
nor U15375 (N_15375,N_14286,N_14518);
xor U15376 (N_15376,N_14607,N_14030);
and U15377 (N_15377,N_14701,N_14319);
or U15378 (N_15378,N_14637,N_14964);
or U15379 (N_15379,N_14369,N_14495);
nand U15380 (N_15380,N_14876,N_14364);
nand U15381 (N_15381,N_14331,N_14315);
nand U15382 (N_15382,N_14906,N_14541);
or U15383 (N_15383,N_14894,N_14665);
nand U15384 (N_15384,N_14707,N_14076);
nand U15385 (N_15385,N_14519,N_14672);
nor U15386 (N_15386,N_14441,N_14915);
or U15387 (N_15387,N_14427,N_14855);
or U15388 (N_15388,N_14031,N_14193);
xnor U15389 (N_15389,N_14391,N_14187);
and U15390 (N_15390,N_14281,N_14640);
or U15391 (N_15391,N_14264,N_14809);
xor U15392 (N_15392,N_14951,N_14155);
xor U15393 (N_15393,N_14033,N_14162);
or U15394 (N_15394,N_14393,N_14336);
and U15395 (N_15395,N_14404,N_14366);
and U15396 (N_15396,N_14387,N_14973);
xor U15397 (N_15397,N_14470,N_14674);
nor U15398 (N_15398,N_14887,N_14539);
or U15399 (N_15399,N_14089,N_14647);
nor U15400 (N_15400,N_14237,N_14205);
nand U15401 (N_15401,N_14990,N_14259);
xor U15402 (N_15402,N_14771,N_14600);
xor U15403 (N_15403,N_14347,N_14595);
and U15404 (N_15404,N_14292,N_14149);
nand U15405 (N_15405,N_14515,N_14545);
nand U15406 (N_15406,N_14020,N_14516);
nor U15407 (N_15407,N_14135,N_14085);
and U15408 (N_15408,N_14846,N_14567);
nor U15409 (N_15409,N_14885,N_14549);
xor U15410 (N_15410,N_14444,N_14253);
and U15411 (N_15411,N_14920,N_14984);
or U15412 (N_15412,N_14313,N_14084);
and U15413 (N_15413,N_14661,N_14302);
nor U15414 (N_15414,N_14214,N_14448);
nand U15415 (N_15415,N_14341,N_14742);
xor U15416 (N_15416,N_14482,N_14698);
xnor U15417 (N_15417,N_14388,N_14561);
nand U15418 (N_15418,N_14533,N_14362);
and U15419 (N_15419,N_14432,N_14382);
nand U15420 (N_15420,N_14376,N_14261);
or U15421 (N_15421,N_14409,N_14840);
nand U15422 (N_15422,N_14880,N_14954);
xnor U15423 (N_15423,N_14962,N_14901);
or U15424 (N_15424,N_14355,N_14706);
or U15425 (N_15425,N_14598,N_14306);
and U15426 (N_15426,N_14276,N_14415);
nand U15427 (N_15427,N_14750,N_14769);
or U15428 (N_15428,N_14802,N_14083);
nand U15429 (N_15429,N_14530,N_14776);
nor U15430 (N_15430,N_14566,N_14746);
and U15431 (N_15431,N_14320,N_14700);
nand U15432 (N_15432,N_14841,N_14832);
nor U15433 (N_15433,N_14138,N_14864);
nand U15434 (N_15434,N_14755,N_14196);
and U15435 (N_15435,N_14309,N_14793);
or U15436 (N_15436,N_14815,N_14210);
xor U15437 (N_15437,N_14289,N_14151);
xor U15438 (N_15438,N_14596,N_14130);
or U15439 (N_15439,N_14743,N_14318);
xor U15440 (N_15440,N_14216,N_14758);
nand U15441 (N_15441,N_14401,N_14462);
or U15442 (N_15442,N_14476,N_14525);
xnor U15443 (N_15443,N_14055,N_14446);
nor U15444 (N_15444,N_14730,N_14383);
and U15445 (N_15445,N_14732,N_14191);
or U15446 (N_15446,N_14977,N_14452);
or U15447 (N_15447,N_14983,N_14035);
and U15448 (N_15448,N_14491,N_14451);
xor U15449 (N_15449,N_14897,N_14818);
and U15450 (N_15450,N_14118,N_14262);
nand U15451 (N_15451,N_14866,N_14671);
and U15452 (N_15452,N_14435,N_14939);
nor U15453 (N_15453,N_14540,N_14029);
nor U15454 (N_15454,N_14953,N_14166);
or U15455 (N_15455,N_14429,N_14621);
nor U15456 (N_15456,N_14349,N_14457);
or U15457 (N_15457,N_14048,N_14251);
xnor U15458 (N_15458,N_14414,N_14551);
xor U15459 (N_15459,N_14231,N_14632);
nor U15460 (N_15460,N_14288,N_14012);
nor U15461 (N_15461,N_14350,N_14574);
nor U15462 (N_15462,N_14828,N_14061);
nor U15463 (N_15463,N_14522,N_14715);
and U15464 (N_15464,N_14099,N_14287);
or U15465 (N_15465,N_14293,N_14649);
and U15466 (N_15466,N_14641,N_14910);
nor U15467 (N_15467,N_14523,N_14716);
and U15468 (N_15468,N_14593,N_14943);
nand U15469 (N_15469,N_14044,N_14359);
and U15470 (N_15470,N_14396,N_14578);
and U15471 (N_15471,N_14417,N_14935);
xor U15472 (N_15472,N_14537,N_14766);
and U15473 (N_15473,N_14552,N_14066);
nor U15474 (N_15474,N_14826,N_14592);
and U15475 (N_15475,N_14363,N_14913);
and U15476 (N_15476,N_14899,N_14011);
and U15477 (N_15477,N_14475,N_14239);
or U15478 (N_15478,N_14690,N_14474);
xnor U15479 (N_15479,N_14631,N_14692);
and U15480 (N_15480,N_14662,N_14082);
and U15481 (N_15481,N_14702,N_14862);
or U15482 (N_15482,N_14994,N_14305);
nand U15483 (N_15483,N_14357,N_14958);
nand U15484 (N_15484,N_14285,N_14623);
or U15485 (N_15485,N_14213,N_14834);
or U15486 (N_15486,N_14759,N_14838);
nand U15487 (N_15487,N_14871,N_14782);
nor U15488 (N_15488,N_14284,N_14100);
nor U15489 (N_15489,N_14431,N_14146);
or U15490 (N_15490,N_14219,N_14479);
nor U15491 (N_15491,N_14573,N_14614);
xor U15492 (N_15492,N_14338,N_14212);
xor U15493 (N_15493,N_14892,N_14634);
xor U15494 (N_15494,N_14610,N_14872);
nand U15495 (N_15495,N_14062,N_14967);
and U15496 (N_15496,N_14299,N_14202);
and U15497 (N_15497,N_14037,N_14344);
nand U15498 (N_15498,N_14733,N_14275);
or U15499 (N_15499,N_14335,N_14890);
xnor U15500 (N_15500,N_14727,N_14434);
xor U15501 (N_15501,N_14747,N_14094);
nor U15502 (N_15502,N_14430,N_14793);
xor U15503 (N_15503,N_14606,N_14235);
nor U15504 (N_15504,N_14489,N_14985);
or U15505 (N_15505,N_14994,N_14410);
and U15506 (N_15506,N_14730,N_14831);
nor U15507 (N_15507,N_14386,N_14852);
xor U15508 (N_15508,N_14644,N_14655);
or U15509 (N_15509,N_14904,N_14423);
and U15510 (N_15510,N_14785,N_14305);
nand U15511 (N_15511,N_14676,N_14847);
or U15512 (N_15512,N_14792,N_14344);
xnor U15513 (N_15513,N_14008,N_14093);
xnor U15514 (N_15514,N_14241,N_14530);
or U15515 (N_15515,N_14102,N_14789);
and U15516 (N_15516,N_14054,N_14795);
nor U15517 (N_15517,N_14961,N_14126);
nand U15518 (N_15518,N_14970,N_14597);
nor U15519 (N_15519,N_14369,N_14826);
xnor U15520 (N_15520,N_14604,N_14174);
or U15521 (N_15521,N_14570,N_14082);
xor U15522 (N_15522,N_14948,N_14997);
and U15523 (N_15523,N_14515,N_14411);
xor U15524 (N_15524,N_14202,N_14295);
or U15525 (N_15525,N_14602,N_14964);
nor U15526 (N_15526,N_14368,N_14205);
or U15527 (N_15527,N_14541,N_14318);
nor U15528 (N_15528,N_14810,N_14244);
or U15529 (N_15529,N_14263,N_14690);
and U15530 (N_15530,N_14838,N_14588);
xor U15531 (N_15531,N_14142,N_14561);
nor U15532 (N_15532,N_14167,N_14696);
nor U15533 (N_15533,N_14072,N_14829);
or U15534 (N_15534,N_14891,N_14169);
nand U15535 (N_15535,N_14796,N_14939);
nor U15536 (N_15536,N_14395,N_14131);
or U15537 (N_15537,N_14596,N_14309);
xor U15538 (N_15538,N_14348,N_14941);
nand U15539 (N_15539,N_14847,N_14591);
nor U15540 (N_15540,N_14467,N_14459);
nand U15541 (N_15541,N_14471,N_14425);
nor U15542 (N_15542,N_14631,N_14296);
or U15543 (N_15543,N_14256,N_14156);
xor U15544 (N_15544,N_14290,N_14305);
nand U15545 (N_15545,N_14797,N_14117);
or U15546 (N_15546,N_14825,N_14819);
or U15547 (N_15547,N_14244,N_14020);
xnor U15548 (N_15548,N_14856,N_14783);
nor U15549 (N_15549,N_14117,N_14907);
xor U15550 (N_15550,N_14716,N_14126);
nor U15551 (N_15551,N_14217,N_14968);
and U15552 (N_15552,N_14176,N_14840);
nand U15553 (N_15553,N_14194,N_14223);
nor U15554 (N_15554,N_14306,N_14842);
nand U15555 (N_15555,N_14178,N_14971);
or U15556 (N_15556,N_14537,N_14790);
xor U15557 (N_15557,N_14610,N_14311);
nor U15558 (N_15558,N_14896,N_14970);
and U15559 (N_15559,N_14227,N_14631);
or U15560 (N_15560,N_14841,N_14548);
or U15561 (N_15561,N_14575,N_14086);
nand U15562 (N_15562,N_14222,N_14178);
nor U15563 (N_15563,N_14639,N_14154);
nor U15564 (N_15564,N_14670,N_14370);
or U15565 (N_15565,N_14440,N_14356);
nor U15566 (N_15566,N_14756,N_14993);
nand U15567 (N_15567,N_14472,N_14669);
nor U15568 (N_15568,N_14007,N_14034);
and U15569 (N_15569,N_14062,N_14117);
and U15570 (N_15570,N_14989,N_14683);
nand U15571 (N_15571,N_14411,N_14582);
and U15572 (N_15572,N_14104,N_14357);
and U15573 (N_15573,N_14916,N_14160);
and U15574 (N_15574,N_14859,N_14462);
and U15575 (N_15575,N_14637,N_14448);
and U15576 (N_15576,N_14574,N_14738);
and U15577 (N_15577,N_14471,N_14227);
or U15578 (N_15578,N_14321,N_14578);
and U15579 (N_15579,N_14436,N_14682);
and U15580 (N_15580,N_14571,N_14068);
or U15581 (N_15581,N_14847,N_14634);
nand U15582 (N_15582,N_14361,N_14556);
nor U15583 (N_15583,N_14381,N_14745);
nor U15584 (N_15584,N_14333,N_14598);
or U15585 (N_15585,N_14693,N_14400);
and U15586 (N_15586,N_14661,N_14355);
and U15587 (N_15587,N_14660,N_14382);
nor U15588 (N_15588,N_14847,N_14161);
nor U15589 (N_15589,N_14980,N_14495);
nor U15590 (N_15590,N_14419,N_14816);
nor U15591 (N_15591,N_14899,N_14583);
nor U15592 (N_15592,N_14122,N_14963);
nor U15593 (N_15593,N_14612,N_14605);
and U15594 (N_15594,N_14982,N_14889);
nand U15595 (N_15595,N_14208,N_14978);
nor U15596 (N_15596,N_14542,N_14405);
xor U15597 (N_15597,N_14158,N_14592);
nor U15598 (N_15598,N_14209,N_14002);
nor U15599 (N_15599,N_14352,N_14612);
nor U15600 (N_15600,N_14872,N_14228);
and U15601 (N_15601,N_14482,N_14936);
nor U15602 (N_15602,N_14135,N_14809);
nand U15603 (N_15603,N_14028,N_14392);
or U15604 (N_15604,N_14933,N_14342);
or U15605 (N_15605,N_14805,N_14311);
or U15606 (N_15606,N_14118,N_14405);
nand U15607 (N_15607,N_14022,N_14682);
xnor U15608 (N_15608,N_14668,N_14025);
xor U15609 (N_15609,N_14332,N_14104);
and U15610 (N_15610,N_14850,N_14512);
nand U15611 (N_15611,N_14323,N_14658);
xnor U15612 (N_15612,N_14225,N_14770);
and U15613 (N_15613,N_14879,N_14774);
or U15614 (N_15614,N_14032,N_14071);
nor U15615 (N_15615,N_14169,N_14198);
and U15616 (N_15616,N_14351,N_14888);
nor U15617 (N_15617,N_14619,N_14692);
xor U15618 (N_15618,N_14209,N_14704);
or U15619 (N_15619,N_14157,N_14543);
nand U15620 (N_15620,N_14264,N_14061);
xnor U15621 (N_15621,N_14214,N_14690);
or U15622 (N_15622,N_14936,N_14013);
nand U15623 (N_15623,N_14213,N_14669);
nand U15624 (N_15624,N_14309,N_14376);
or U15625 (N_15625,N_14190,N_14785);
xnor U15626 (N_15626,N_14337,N_14836);
nand U15627 (N_15627,N_14520,N_14422);
or U15628 (N_15628,N_14592,N_14665);
and U15629 (N_15629,N_14656,N_14871);
xor U15630 (N_15630,N_14255,N_14906);
nor U15631 (N_15631,N_14809,N_14690);
xor U15632 (N_15632,N_14473,N_14733);
nor U15633 (N_15633,N_14714,N_14044);
nor U15634 (N_15634,N_14313,N_14828);
nor U15635 (N_15635,N_14905,N_14213);
xnor U15636 (N_15636,N_14377,N_14539);
and U15637 (N_15637,N_14927,N_14513);
and U15638 (N_15638,N_14973,N_14934);
or U15639 (N_15639,N_14418,N_14022);
nand U15640 (N_15640,N_14256,N_14181);
xnor U15641 (N_15641,N_14148,N_14520);
xor U15642 (N_15642,N_14335,N_14141);
nand U15643 (N_15643,N_14320,N_14599);
xnor U15644 (N_15644,N_14167,N_14689);
nand U15645 (N_15645,N_14120,N_14414);
or U15646 (N_15646,N_14274,N_14162);
xor U15647 (N_15647,N_14478,N_14108);
and U15648 (N_15648,N_14529,N_14880);
xnor U15649 (N_15649,N_14155,N_14215);
or U15650 (N_15650,N_14386,N_14183);
nor U15651 (N_15651,N_14477,N_14667);
and U15652 (N_15652,N_14009,N_14016);
nor U15653 (N_15653,N_14138,N_14910);
and U15654 (N_15654,N_14450,N_14916);
or U15655 (N_15655,N_14391,N_14143);
nand U15656 (N_15656,N_14713,N_14021);
nor U15657 (N_15657,N_14765,N_14089);
xor U15658 (N_15658,N_14632,N_14930);
and U15659 (N_15659,N_14500,N_14779);
xnor U15660 (N_15660,N_14457,N_14076);
or U15661 (N_15661,N_14267,N_14165);
and U15662 (N_15662,N_14411,N_14185);
and U15663 (N_15663,N_14027,N_14190);
xnor U15664 (N_15664,N_14745,N_14919);
nor U15665 (N_15665,N_14784,N_14941);
nand U15666 (N_15666,N_14302,N_14321);
xnor U15667 (N_15667,N_14546,N_14215);
nand U15668 (N_15668,N_14134,N_14173);
and U15669 (N_15669,N_14269,N_14310);
xnor U15670 (N_15670,N_14663,N_14777);
or U15671 (N_15671,N_14206,N_14790);
nand U15672 (N_15672,N_14427,N_14069);
nand U15673 (N_15673,N_14062,N_14795);
nor U15674 (N_15674,N_14350,N_14218);
xor U15675 (N_15675,N_14666,N_14764);
or U15676 (N_15676,N_14658,N_14102);
nor U15677 (N_15677,N_14130,N_14592);
nor U15678 (N_15678,N_14225,N_14045);
and U15679 (N_15679,N_14660,N_14227);
nor U15680 (N_15680,N_14669,N_14402);
xor U15681 (N_15681,N_14451,N_14788);
xnor U15682 (N_15682,N_14160,N_14866);
and U15683 (N_15683,N_14236,N_14473);
and U15684 (N_15684,N_14031,N_14360);
xor U15685 (N_15685,N_14670,N_14883);
and U15686 (N_15686,N_14170,N_14954);
nand U15687 (N_15687,N_14513,N_14885);
nor U15688 (N_15688,N_14925,N_14774);
and U15689 (N_15689,N_14033,N_14094);
and U15690 (N_15690,N_14976,N_14620);
nor U15691 (N_15691,N_14107,N_14821);
and U15692 (N_15692,N_14677,N_14036);
xnor U15693 (N_15693,N_14376,N_14803);
xnor U15694 (N_15694,N_14072,N_14534);
nand U15695 (N_15695,N_14214,N_14600);
and U15696 (N_15696,N_14970,N_14415);
nand U15697 (N_15697,N_14835,N_14066);
xor U15698 (N_15698,N_14523,N_14634);
or U15699 (N_15699,N_14073,N_14133);
xnor U15700 (N_15700,N_14913,N_14081);
nor U15701 (N_15701,N_14956,N_14291);
xnor U15702 (N_15702,N_14519,N_14916);
nor U15703 (N_15703,N_14625,N_14297);
or U15704 (N_15704,N_14263,N_14169);
and U15705 (N_15705,N_14838,N_14377);
nand U15706 (N_15706,N_14216,N_14221);
xor U15707 (N_15707,N_14154,N_14450);
and U15708 (N_15708,N_14376,N_14762);
nor U15709 (N_15709,N_14519,N_14743);
or U15710 (N_15710,N_14988,N_14743);
nor U15711 (N_15711,N_14830,N_14052);
and U15712 (N_15712,N_14258,N_14562);
nand U15713 (N_15713,N_14514,N_14961);
nand U15714 (N_15714,N_14211,N_14786);
or U15715 (N_15715,N_14978,N_14738);
nand U15716 (N_15716,N_14626,N_14593);
and U15717 (N_15717,N_14566,N_14818);
xnor U15718 (N_15718,N_14910,N_14842);
xor U15719 (N_15719,N_14152,N_14460);
nor U15720 (N_15720,N_14376,N_14057);
and U15721 (N_15721,N_14548,N_14097);
and U15722 (N_15722,N_14127,N_14596);
xor U15723 (N_15723,N_14398,N_14915);
nor U15724 (N_15724,N_14752,N_14519);
xnor U15725 (N_15725,N_14007,N_14272);
xor U15726 (N_15726,N_14274,N_14291);
or U15727 (N_15727,N_14977,N_14584);
nor U15728 (N_15728,N_14599,N_14246);
nand U15729 (N_15729,N_14594,N_14781);
nand U15730 (N_15730,N_14556,N_14654);
and U15731 (N_15731,N_14292,N_14195);
nand U15732 (N_15732,N_14210,N_14043);
and U15733 (N_15733,N_14660,N_14694);
or U15734 (N_15734,N_14776,N_14717);
or U15735 (N_15735,N_14166,N_14884);
xor U15736 (N_15736,N_14966,N_14925);
nand U15737 (N_15737,N_14180,N_14585);
nor U15738 (N_15738,N_14104,N_14116);
nand U15739 (N_15739,N_14623,N_14105);
nand U15740 (N_15740,N_14412,N_14149);
nand U15741 (N_15741,N_14981,N_14545);
and U15742 (N_15742,N_14435,N_14707);
xnor U15743 (N_15743,N_14527,N_14564);
nor U15744 (N_15744,N_14072,N_14229);
nor U15745 (N_15745,N_14261,N_14936);
and U15746 (N_15746,N_14957,N_14100);
nor U15747 (N_15747,N_14720,N_14007);
nand U15748 (N_15748,N_14888,N_14264);
nand U15749 (N_15749,N_14129,N_14908);
xnor U15750 (N_15750,N_14360,N_14280);
xnor U15751 (N_15751,N_14053,N_14002);
nor U15752 (N_15752,N_14202,N_14964);
xor U15753 (N_15753,N_14214,N_14644);
xnor U15754 (N_15754,N_14728,N_14741);
nor U15755 (N_15755,N_14288,N_14942);
nand U15756 (N_15756,N_14742,N_14148);
nand U15757 (N_15757,N_14975,N_14380);
and U15758 (N_15758,N_14471,N_14988);
and U15759 (N_15759,N_14443,N_14335);
or U15760 (N_15760,N_14638,N_14524);
and U15761 (N_15761,N_14919,N_14741);
and U15762 (N_15762,N_14542,N_14088);
nor U15763 (N_15763,N_14651,N_14663);
nor U15764 (N_15764,N_14923,N_14217);
nand U15765 (N_15765,N_14883,N_14003);
or U15766 (N_15766,N_14150,N_14442);
nand U15767 (N_15767,N_14249,N_14400);
nand U15768 (N_15768,N_14308,N_14160);
nor U15769 (N_15769,N_14255,N_14650);
xor U15770 (N_15770,N_14934,N_14118);
nor U15771 (N_15771,N_14444,N_14110);
xor U15772 (N_15772,N_14111,N_14956);
nand U15773 (N_15773,N_14015,N_14672);
and U15774 (N_15774,N_14807,N_14267);
or U15775 (N_15775,N_14713,N_14398);
nor U15776 (N_15776,N_14847,N_14976);
nor U15777 (N_15777,N_14839,N_14587);
xnor U15778 (N_15778,N_14705,N_14384);
nor U15779 (N_15779,N_14617,N_14781);
and U15780 (N_15780,N_14408,N_14975);
nor U15781 (N_15781,N_14829,N_14956);
and U15782 (N_15782,N_14313,N_14285);
xor U15783 (N_15783,N_14497,N_14410);
and U15784 (N_15784,N_14360,N_14771);
nand U15785 (N_15785,N_14059,N_14169);
or U15786 (N_15786,N_14465,N_14157);
nor U15787 (N_15787,N_14631,N_14576);
nand U15788 (N_15788,N_14699,N_14460);
nor U15789 (N_15789,N_14915,N_14821);
and U15790 (N_15790,N_14038,N_14838);
nor U15791 (N_15791,N_14939,N_14650);
nand U15792 (N_15792,N_14661,N_14995);
and U15793 (N_15793,N_14361,N_14996);
or U15794 (N_15794,N_14835,N_14754);
nand U15795 (N_15795,N_14806,N_14308);
nand U15796 (N_15796,N_14924,N_14742);
nand U15797 (N_15797,N_14578,N_14415);
and U15798 (N_15798,N_14811,N_14639);
nor U15799 (N_15799,N_14443,N_14373);
or U15800 (N_15800,N_14408,N_14924);
nor U15801 (N_15801,N_14702,N_14697);
xor U15802 (N_15802,N_14471,N_14859);
nand U15803 (N_15803,N_14887,N_14816);
nor U15804 (N_15804,N_14801,N_14691);
or U15805 (N_15805,N_14832,N_14528);
xnor U15806 (N_15806,N_14877,N_14296);
nand U15807 (N_15807,N_14169,N_14883);
xor U15808 (N_15808,N_14835,N_14060);
and U15809 (N_15809,N_14019,N_14744);
nand U15810 (N_15810,N_14551,N_14954);
and U15811 (N_15811,N_14207,N_14275);
or U15812 (N_15812,N_14452,N_14207);
nor U15813 (N_15813,N_14334,N_14781);
or U15814 (N_15814,N_14772,N_14608);
xor U15815 (N_15815,N_14617,N_14431);
nor U15816 (N_15816,N_14483,N_14571);
or U15817 (N_15817,N_14138,N_14802);
or U15818 (N_15818,N_14545,N_14449);
nor U15819 (N_15819,N_14229,N_14868);
or U15820 (N_15820,N_14691,N_14395);
xor U15821 (N_15821,N_14658,N_14820);
nor U15822 (N_15822,N_14766,N_14553);
xor U15823 (N_15823,N_14099,N_14688);
and U15824 (N_15824,N_14465,N_14546);
or U15825 (N_15825,N_14994,N_14212);
nor U15826 (N_15826,N_14527,N_14434);
and U15827 (N_15827,N_14812,N_14901);
and U15828 (N_15828,N_14423,N_14295);
nor U15829 (N_15829,N_14617,N_14015);
nand U15830 (N_15830,N_14477,N_14877);
nor U15831 (N_15831,N_14214,N_14575);
and U15832 (N_15832,N_14621,N_14258);
and U15833 (N_15833,N_14118,N_14708);
or U15834 (N_15834,N_14596,N_14308);
or U15835 (N_15835,N_14702,N_14252);
nand U15836 (N_15836,N_14764,N_14194);
or U15837 (N_15837,N_14396,N_14032);
xnor U15838 (N_15838,N_14599,N_14995);
xnor U15839 (N_15839,N_14846,N_14042);
nand U15840 (N_15840,N_14058,N_14617);
xor U15841 (N_15841,N_14819,N_14153);
nand U15842 (N_15842,N_14070,N_14840);
or U15843 (N_15843,N_14931,N_14464);
and U15844 (N_15844,N_14937,N_14898);
xnor U15845 (N_15845,N_14265,N_14010);
xor U15846 (N_15846,N_14885,N_14008);
nand U15847 (N_15847,N_14691,N_14818);
and U15848 (N_15848,N_14628,N_14395);
xor U15849 (N_15849,N_14507,N_14375);
nand U15850 (N_15850,N_14638,N_14537);
nand U15851 (N_15851,N_14761,N_14838);
nand U15852 (N_15852,N_14440,N_14773);
nand U15853 (N_15853,N_14497,N_14656);
nand U15854 (N_15854,N_14989,N_14950);
xor U15855 (N_15855,N_14083,N_14492);
or U15856 (N_15856,N_14524,N_14526);
xnor U15857 (N_15857,N_14908,N_14603);
and U15858 (N_15858,N_14318,N_14639);
nor U15859 (N_15859,N_14718,N_14502);
and U15860 (N_15860,N_14838,N_14356);
and U15861 (N_15861,N_14830,N_14439);
xor U15862 (N_15862,N_14742,N_14955);
xnor U15863 (N_15863,N_14736,N_14394);
or U15864 (N_15864,N_14954,N_14299);
or U15865 (N_15865,N_14753,N_14506);
xor U15866 (N_15866,N_14950,N_14622);
xnor U15867 (N_15867,N_14093,N_14393);
and U15868 (N_15868,N_14397,N_14584);
or U15869 (N_15869,N_14461,N_14392);
nor U15870 (N_15870,N_14188,N_14414);
or U15871 (N_15871,N_14692,N_14942);
xor U15872 (N_15872,N_14915,N_14754);
nor U15873 (N_15873,N_14823,N_14504);
nand U15874 (N_15874,N_14578,N_14500);
xnor U15875 (N_15875,N_14067,N_14390);
nor U15876 (N_15876,N_14638,N_14528);
xor U15877 (N_15877,N_14598,N_14227);
nor U15878 (N_15878,N_14559,N_14628);
nor U15879 (N_15879,N_14463,N_14535);
xor U15880 (N_15880,N_14005,N_14289);
nor U15881 (N_15881,N_14714,N_14880);
xnor U15882 (N_15882,N_14620,N_14666);
and U15883 (N_15883,N_14519,N_14910);
and U15884 (N_15884,N_14236,N_14549);
and U15885 (N_15885,N_14355,N_14866);
nor U15886 (N_15886,N_14241,N_14959);
nand U15887 (N_15887,N_14917,N_14984);
xor U15888 (N_15888,N_14511,N_14843);
or U15889 (N_15889,N_14153,N_14462);
and U15890 (N_15890,N_14797,N_14324);
and U15891 (N_15891,N_14851,N_14730);
nor U15892 (N_15892,N_14441,N_14700);
xor U15893 (N_15893,N_14235,N_14531);
nor U15894 (N_15894,N_14536,N_14214);
nor U15895 (N_15895,N_14762,N_14958);
nand U15896 (N_15896,N_14109,N_14251);
and U15897 (N_15897,N_14741,N_14634);
and U15898 (N_15898,N_14212,N_14512);
or U15899 (N_15899,N_14578,N_14350);
xnor U15900 (N_15900,N_14381,N_14372);
nor U15901 (N_15901,N_14177,N_14360);
nor U15902 (N_15902,N_14241,N_14406);
nand U15903 (N_15903,N_14112,N_14349);
or U15904 (N_15904,N_14998,N_14933);
or U15905 (N_15905,N_14277,N_14766);
xor U15906 (N_15906,N_14549,N_14791);
nand U15907 (N_15907,N_14069,N_14816);
xor U15908 (N_15908,N_14503,N_14581);
and U15909 (N_15909,N_14705,N_14883);
or U15910 (N_15910,N_14869,N_14181);
or U15911 (N_15911,N_14344,N_14124);
and U15912 (N_15912,N_14377,N_14549);
nor U15913 (N_15913,N_14316,N_14941);
and U15914 (N_15914,N_14085,N_14677);
xor U15915 (N_15915,N_14145,N_14177);
or U15916 (N_15916,N_14762,N_14171);
nor U15917 (N_15917,N_14959,N_14046);
and U15918 (N_15918,N_14531,N_14372);
nand U15919 (N_15919,N_14836,N_14573);
nand U15920 (N_15920,N_14822,N_14406);
or U15921 (N_15921,N_14165,N_14266);
and U15922 (N_15922,N_14459,N_14241);
xnor U15923 (N_15923,N_14279,N_14790);
xnor U15924 (N_15924,N_14330,N_14299);
xor U15925 (N_15925,N_14787,N_14184);
nor U15926 (N_15926,N_14412,N_14542);
nand U15927 (N_15927,N_14588,N_14788);
xor U15928 (N_15928,N_14229,N_14316);
or U15929 (N_15929,N_14750,N_14634);
or U15930 (N_15930,N_14438,N_14094);
nor U15931 (N_15931,N_14322,N_14417);
nor U15932 (N_15932,N_14458,N_14167);
nand U15933 (N_15933,N_14662,N_14009);
or U15934 (N_15934,N_14644,N_14084);
xnor U15935 (N_15935,N_14706,N_14389);
nand U15936 (N_15936,N_14977,N_14702);
xor U15937 (N_15937,N_14153,N_14798);
nor U15938 (N_15938,N_14560,N_14150);
nand U15939 (N_15939,N_14227,N_14710);
xnor U15940 (N_15940,N_14253,N_14757);
nand U15941 (N_15941,N_14121,N_14863);
nor U15942 (N_15942,N_14867,N_14270);
nand U15943 (N_15943,N_14493,N_14588);
nor U15944 (N_15944,N_14375,N_14555);
nand U15945 (N_15945,N_14494,N_14794);
and U15946 (N_15946,N_14462,N_14822);
and U15947 (N_15947,N_14527,N_14821);
and U15948 (N_15948,N_14620,N_14508);
nand U15949 (N_15949,N_14677,N_14754);
and U15950 (N_15950,N_14819,N_14955);
and U15951 (N_15951,N_14305,N_14125);
nor U15952 (N_15952,N_14017,N_14832);
nand U15953 (N_15953,N_14016,N_14448);
and U15954 (N_15954,N_14652,N_14490);
xor U15955 (N_15955,N_14858,N_14997);
nor U15956 (N_15956,N_14940,N_14623);
xnor U15957 (N_15957,N_14941,N_14397);
and U15958 (N_15958,N_14559,N_14768);
nor U15959 (N_15959,N_14735,N_14892);
or U15960 (N_15960,N_14106,N_14083);
or U15961 (N_15961,N_14725,N_14306);
nor U15962 (N_15962,N_14098,N_14790);
nor U15963 (N_15963,N_14458,N_14608);
or U15964 (N_15964,N_14097,N_14165);
xnor U15965 (N_15965,N_14864,N_14100);
nand U15966 (N_15966,N_14350,N_14720);
xor U15967 (N_15967,N_14045,N_14601);
and U15968 (N_15968,N_14749,N_14012);
and U15969 (N_15969,N_14182,N_14359);
nor U15970 (N_15970,N_14664,N_14922);
xor U15971 (N_15971,N_14559,N_14328);
nand U15972 (N_15972,N_14549,N_14814);
and U15973 (N_15973,N_14701,N_14129);
nand U15974 (N_15974,N_14166,N_14371);
nand U15975 (N_15975,N_14829,N_14762);
or U15976 (N_15976,N_14912,N_14254);
nor U15977 (N_15977,N_14726,N_14037);
nand U15978 (N_15978,N_14926,N_14570);
xnor U15979 (N_15979,N_14760,N_14659);
nor U15980 (N_15980,N_14986,N_14526);
and U15981 (N_15981,N_14168,N_14105);
or U15982 (N_15982,N_14089,N_14477);
xnor U15983 (N_15983,N_14915,N_14148);
nand U15984 (N_15984,N_14388,N_14108);
and U15985 (N_15985,N_14031,N_14339);
or U15986 (N_15986,N_14170,N_14927);
nor U15987 (N_15987,N_14838,N_14942);
xnor U15988 (N_15988,N_14573,N_14306);
or U15989 (N_15989,N_14739,N_14853);
xor U15990 (N_15990,N_14168,N_14832);
xor U15991 (N_15991,N_14343,N_14380);
xnor U15992 (N_15992,N_14181,N_14368);
xnor U15993 (N_15993,N_14907,N_14304);
nand U15994 (N_15994,N_14076,N_14077);
nand U15995 (N_15995,N_14429,N_14583);
nor U15996 (N_15996,N_14421,N_14152);
or U15997 (N_15997,N_14092,N_14130);
or U15998 (N_15998,N_14581,N_14086);
nor U15999 (N_15999,N_14278,N_14997);
or U16000 (N_16000,N_15706,N_15053);
nand U16001 (N_16001,N_15959,N_15962);
and U16002 (N_16002,N_15007,N_15818);
nand U16003 (N_16003,N_15293,N_15665);
nand U16004 (N_16004,N_15064,N_15949);
and U16005 (N_16005,N_15375,N_15082);
or U16006 (N_16006,N_15975,N_15738);
nor U16007 (N_16007,N_15542,N_15645);
nand U16008 (N_16008,N_15809,N_15444);
nand U16009 (N_16009,N_15864,N_15886);
or U16010 (N_16010,N_15572,N_15199);
xor U16011 (N_16011,N_15580,N_15119);
nor U16012 (N_16012,N_15845,N_15495);
and U16013 (N_16013,N_15766,N_15842);
and U16014 (N_16014,N_15807,N_15477);
or U16015 (N_16015,N_15908,N_15009);
nor U16016 (N_16016,N_15750,N_15037);
and U16017 (N_16017,N_15493,N_15203);
or U16018 (N_16018,N_15896,N_15419);
xor U16019 (N_16019,N_15163,N_15618);
nand U16020 (N_16020,N_15800,N_15210);
nand U16021 (N_16021,N_15290,N_15504);
nor U16022 (N_16022,N_15924,N_15660);
and U16023 (N_16023,N_15933,N_15191);
xor U16024 (N_16024,N_15882,N_15992);
nor U16025 (N_16025,N_15252,N_15362);
nor U16026 (N_16026,N_15140,N_15830);
and U16027 (N_16027,N_15793,N_15705);
xnor U16028 (N_16028,N_15556,N_15712);
nand U16029 (N_16029,N_15247,N_15023);
nor U16030 (N_16030,N_15784,N_15781);
or U16031 (N_16031,N_15769,N_15868);
xor U16032 (N_16032,N_15369,N_15161);
or U16033 (N_16033,N_15209,N_15285);
and U16034 (N_16034,N_15219,N_15936);
and U16035 (N_16035,N_15906,N_15520);
and U16036 (N_16036,N_15491,N_15869);
xor U16037 (N_16037,N_15368,N_15325);
xor U16038 (N_16038,N_15694,N_15676);
xnor U16039 (N_16039,N_15630,N_15165);
and U16040 (N_16040,N_15976,N_15576);
nand U16041 (N_16041,N_15981,N_15431);
and U16042 (N_16042,N_15879,N_15217);
or U16043 (N_16043,N_15611,N_15302);
nor U16044 (N_16044,N_15555,N_15841);
or U16045 (N_16045,N_15097,N_15100);
or U16046 (N_16046,N_15207,N_15796);
xor U16047 (N_16047,N_15945,N_15399);
and U16048 (N_16048,N_15497,N_15273);
or U16049 (N_16049,N_15136,N_15022);
xnor U16050 (N_16050,N_15673,N_15454);
nor U16051 (N_16051,N_15755,N_15578);
nand U16052 (N_16052,N_15885,N_15794);
nor U16053 (N_16053,N_15324,N_15288);
nor U16054 (N_16054,N_15175,N_15438);
nor U16055 (N_16055,N_15548,N_15326);
nor U16056 (N_16056,N_15294,N_15249);
and U16057 (N_16057,N_15476,N_15226);
or U16058 (N_16058,N_15122,N_15735);
and U16059 (N_16059,N_15397,N_15066);
nor U16060 (N_16060,N_15982,N_15530);
nor U16061 (N_16061,N_15200,N_15923);
or U16062 (N_16062,N_15212,N_15157);
or U16063 (N_16063,N_15172,N_15246);
and U16064 (N_16064,N_15391,N_15460);
and U16065 (N_16065,N_15029,N_15268);
and U16066 (N_16066,N_15633,N_15357);
xor U16067 (N_16067,N_15797,N_15051);
and U16068 (N_16068,N_15299,N_15147);
xor U16069 (N_16069,N_15545,N_15870);
xnor U16070 (N_16070,N_15899,N_15615);
or U16071 (N_16071,N_15048,N_15472);
xor U16072 (N_16072,N_15732,N_15332);
xor U16073 (N_16073,N_15713,N_15902);
and U16074 (N_16074,N_15060,N_15470);
nand U16075 (N_16075,N_15216,N_15636);
xnor U16076 (N_16076,N_15322,N_15812);
nor U16077 (N_16077,N_15746,N_15271);
xor U16078 (N_16078,N_15792,N_15595);
and U16079 (N_16079,N_15894,N_15608);
and U16080 (N_16080,N_15364,N_15853);
or U16081 (N_16081,N_15654,N_15741);
xnor U16082 (N_16082,N_15878,N_15173);
and U16083 (N_16083,N_15748,N_15671);
nor U16084 (N_16084,N_15047,N_15932);
and U16085 (N_16085,N_15839,N_15604);
nor U16086 (N_16086,N_15838,N_15046);
xor U16087 (N_16087,N_15704,N_15346);
and U16088 (N_16088,N_15774,N_15162);
xor U16089 (N_16089,N_15478,N_15736);
or U16090 (N_16090,N_15450,N_15406);
xor U16091 (N_16091,N_15124,N_15951);
nor U16092 (N_16092,N_15972,N_15335);
xnor U16093 (N_16093,N_15456,N_15843);
nand U16094 (N_16094,N_15502,N_15835);
nor U16095 (N_16095,N_15234,N_15743);
nand U16096 (N_16096,N_15912,N_15967);
nand U16097 (N_16097,N_15319,N_15866);
xnor U16098 (N_16098,N_15170,N_15457);
and U16099 (N_16099,N_15426,N_15400);
nor U16100 (N_16100,N_15821,N_15084);
or U16101 (N_16101,N_15235,N_15928);
xnor U16102 (N_16102,N_15286,N_15516);
xnor U16103 (N_16103,N_15381,N_15907);
and U16104 (N_16104,N_15267,N_15513);
or U16105 (N_16105,N_15336,N_15343);
xor U16106 (N_16106,N_15825,N_15443);
and U16107 (N_16107,N_15767,N_15910);
and U16108 (N_16108,N_15471,N_15638);
nand U16109 (N_16109,N_15881,N_15204);
or U16110 (N_16110,N_15684,N_15939);
and U16111 (N_16111,N_15742,N_15389);
nor U16112 (N_16112,N_15984,N_15639);
and U16113 (N_16113,N_15418,N_15698);
nand U16114 (N_16114,N_15269,N_15806);
nor U16115 (N_16115,N_15832,N_15720);
nor U16116 (N_16116,N_15069,N_15144);
xnor U16117 (N_16117,N_15721,N_15733);
and U16118 (N_16118,N_15768,N_15737);
and U16119 (N_16119,N_15691,N_15863);
and U16120 (N_16120,N_15014,N_15152);
xnor U16121 (N_16121,N_15142,N_15401);
and U16122 (N_16122,N_15801,N_15817);
nor U16123 (N_16123,N_15957,N_15301);
or U16124 (N_16124,N_15120,N_15466);
nor U16125 (N_16125,N_15323,N_15522);
xor U16126 (N_16126,N_15541,N_15651);
or U16127 (N_16127,N_15770,N_15937);
nand U16128 (N_16128,N_15177,N_15820);
and U16129 (N_16129,N_15339,N_15641);
nand U16130 (N_16130,N_15752,N_15396);
nor U16131 (N_16131,N_15888,N_15221);
and U16132 (N_16132,N_15692,N_15222);
xor U16133 (N_16133,N_15554,N_15791);
nand U16134 (N_16134,N_15284,N_15379);
or U16135 (N_16135,N_15535,N_15997);
nand U16136 (N_16136,N_15954,N_15505);
and U16137 (N_16137,N_15617,N_15722);
or U16138 (N_16138,N_15955,N_15042);
nand U16139 (N_16139,N_15340,N_15307);
and U16140 (N_16140,N_15085,N_15151);
nor U16141 (N_16141,N_15353,N_15640);
nor U16142 (N_16142,N_15185,N_15930);
and U16143 (N_16143,N_15697,N_15168);
nor U16144 (N_16144,N_15628,N_15183);
and U16145 (N_16145,N_15537,N_15492);
or U16146 (N_16146,N_15749,N_15433);
or U16147 (N_16147,N_15417,N_15826);
and U16148 (N_16148,N_15484,N_15305);
nand U16149 (N_16149,N_15805,N_15683);
nand U16150 (N_16150,N_15071,N_15757);
nand U16151 (N_16151,N_15412,N_15371);
nand U16152 (N_16152,N_15104,N_15019);
and U16153 (N_16153,N_15459,N_15550);
and U16154 (N_16154,N_15499,N_15708);
or U16155 (N_16155,N_15095,N_15181);
and U16156 (N_16156,N_15099,N_15810);
and U16157 (N_16157,N_15089,N_15624);
and U16158 (N_16158,N_15623,N_15730);
and U16159 (N_16159,N_15897,N_15929);
nand U16160 (N_16160,N_15449,N_15904);
xnor U16161 (N_16161,N_15905,N_15458);
xnor U16162 (N_16162,N_15862,N_15447);
nand U16163 (N_16163,N_15026,N_15110);
nor U16164 (N_16164,N_15509,N_15227);
and U16165 (N_16165,N_15622,N_15822);
xnor U16166 (N_16166,N_15376,N_15446);
xnor U16167 (N_16167,N_15365,N_15875);
and U16168 (N_16168,N_15612,N_15436);
and U16169 (N_16169,N_15424,N_15004);
nor U16170 (N_16170,N_15551,N_15836);
or U16171 (N_16171,N_15614,N_15565);
nor U16172 (N_16172,N_15442,N_15101);
nor U16173 (N_16173,N_15804,N_15359);
nor U16174 (N_16174,N_15036,N_15861);
xnor U16175 (N_16175,N_15880,N_15176);
and U16176 (N_16176,N_15423,N_15489);
and U16177 (N_16177,N_15111,N_15577);
and U16178 (N_16178,N_15616,N_15229);
nor U16179 (N_16179,N_15903,N_15164);
xnor U16180 (N_16180,N_15874,N_15569);
nand U16181 (N_16181,N_15560,N_15663);
and U16182 (N_16182,N_15116,N_15409);
or U16183 (N_16183,N_15010,N_15392);
nor U16184 (N_16184,N_15073,N_15552);
xor U16185 (N_16185,N_15281,N_15236);
nor U16186 (N_16186,N_15374,N_15244);
xor U16187 (N_16187,N_15351,N_15133);
xnor U16188 (N_16188,N_15564,N_15334);
xnor U16189 (N_16189,N_15964,N_15344);
xor U16190 (N_16190,N_15778,N_15581);
or U16191 (N_16191,N_15065,N_15186);
and U16192 (N_16192,N_15402,N_15420);
xor U16193 (N_16193,N_15811,N_15772);
xor U16194 (N_16194,N_15372,N_15202);
nand U16195 (N_16195,N_15734,N_15859);
nor U16196 (N_16196,N_15331,N_15126);
and U16197 (N_16197,N_15263,N_15296);
or U16198 (N_16198,N_15473,N_15919);
or U16199 (N_16199,N_15789,N_15598);
xnor U16200 (N_16200,N_15740,N_15021);
xor U16201 (N_16201,N_15448,N_15974);
and U16202 (N_16202,N_15931,N_15461);
nand U16203 (N_16203,N_15352,N_15309);
nand U16204 (N_16204,N_15096,N_15070);
nand U16205 (N_16205,N_15664,N_15731);
nand U16206 (N_16206,N_15277,N_15189);
nand U16207 (N_16207,N_15264,N_15559);
and U16208 (N_16208,N_15129,N_15206);
and U16209 (N_16209,N_15606,N_15239);
xnor U16210 (N_16210,N_15350,N_15068);
nand U16211 (N_16211,N_15137,N_15819);
and U16212 (N_16212,N_15287,N_15840);
nand U16213 (N_16213,N_15403,N_15873);
nor U16214 (N_16214,N_15190,N_15024);
xor U16215 (N_16215,N_15017,N_15983);
nor U16216 (N_16216,N_15927,N_15251);
nor U16217 (N_16217,N_15751,N_15395);
nand U16218 (N_16218,N_15557,N_15025);
or U16219 (N_16219,N_15970,N_15965);
nand U16220 (N_16220,N_15425,N_15045);
nand U16221 (N_16221,N_15278,N_15103);
xnor U16222 (N_16222,N_15078,N_15107);
nand U16223 (N_16223,N_15649,N_15016);
nand U16224 (N_16224,N_15989,N_15546);
or U16225 (N_16225,N_15451,N_15005);
or U16226 (N_16226,N_15525,N_15867);
xnor U16227 (N_16227,N_15568,N_15410);
and U16228 (N_16228,N_15411,N_15102);
nand U16229 (N_16229,N_15943,N_15058);
nand U16230 (N_16230,N_15166,N_15726);
nand U16231 (N_16231,N_15533,N_15935);
and U16232 (N_16232,N_15098,N_15799);
xnor U16233 (N_16233,N_15637,N_15013);
or U16234 (N_16234,N_15416,N_15709);
or U16235 (N_16235,N_15320,N_15918);
nand U16236 (N_16236,N_15490,N_15231);
and U16237 (N_16237,N_15384,N_15536);
or U16238 (N_16238,N_15380,N_15519);
or U16239 (N_16239,N_15553,N_15215);
xor U16240 (N_16240,N_15475,N_15891);
nor U16241 (N_16241,N_15327,N_15884);
nand U16242 (N_16242,N_15463,N_15600);
nand U16243 (N_16243,N_15871,N_15012);
nor U16244 (N_16244,N_15383,N_15667);
nand U16245 (N_16245,N_15532,N_15243);
xnor U16246 (N_16246,N_15824,N_15790);
nor U16247 (N_16247,N_15890,N_15590);
nand U16248 (N_16248,N_15958,N_15341);
nand U16249 (N_16249,N_15586,N_15682);
xnor U16250 (N_16250,N_15067,N_15218);
xnor U16251 (N_16251,N_15503,N_15828);
nor U16252 (N_16252,N_15934,N_15086);
nor U16253 (N_16253,N_15558,N_15571);
and U16254 (N_16254,N_15583,N_15198);
and U16255 (N_16255,N_15940,N_15224);
xnor U16256 (N_16256,N_15777,N_15501);
nor U16257 (N_16257,N_15312,N_15679);
and U16258 (N_16258,N_15388,N_15213);
and U16259 (N_16259,N_15413,N_15081);
and U16260 (N_16260,N_15776,N_15854);
nor U16261 (N_16261,N_15701,N_15015);
nor U16262 (N_16262,N_15011,N_15494);
nand U16263 (N_16263,N_15926,N_15690);
or U16264 (N_16264,N_15452,N_15193);
xnor U16265 (N_16265,N_15146,N_15963);
and U16266 (N_16266,N_15474,N_15508);
nor U16267 (N_16267,N_15837,N_15169);
and U16268 (N_16268,N_15815,N_15020);
xnor U16269 (N_16269,N_15913,N_15729);
nand U16270 (N_16270,N_15370,N_15232);
and U16271 (N_16271,N_15445,N_15857);
and U16272 (N_16272,N_15160,N_15373);
or U16273 (N_16273,N_15348,N_15059);
or U16274 (N_16274,N_15834,N_15670);
nand U16275 (N_16275,N_15329,N_15194);
or U16276 (N_16276,N_15382,N_15518);
nand U16277 (N_16277,N_15464,N_15969);
xor U16278 (N_16278,N_15192,N_15316);
or U16279 (N_16279,N_15121,N_15597);
nor U16280 (N_16280,N_15892,N_15266);
and U16281 (N_16281,N_15328,N_15174);
xor U16282 (N_16282,N_15582,N_15238);
xnor U16283 (N_16283,N_15860,N_15893);
nor U16284 (N_16284,N_15018,N_15008);
xor U16285 (N_16285,N_15377,N_15703);
and U16286 (N_16286,N_15526,N_15915);
nor U16287 (N_16287,N_15657,N_15487);
nand U16288 (N_16288,N_15063,N_15245);
and U16289 (N_16289,N_15027,N_15753);
nand U16290 (N_16290,N_15167,N_15297);
and U16291 (N_16291,N_15716,N_15944);
nand U16292 (N_16292,N_15437,N_15714);
nand U16293 (N_16293,N_15148,N_15594);
nor U16294 (N_16294,N_15780,N_15242);
xnor U16295 (N_16295,N_15986,N_15061);
xor U16296 (N_16296,N_15515,N_15998);
nor U16297 (N_16297,N_15865,N_15197);
nor U16298 (N_16298,N_15909,N_15523);
nand U16299 (N_16299,N_15653,N_15304);
and U16300 (N_16300,N_15948,N_15076);
nand U16301 (N_16301,N_15872,N_15917);
and U16302 (N_16302,N_15366,N_15338);
xor U16303 (N_16303,N_15440,N_15265);
or U16304 (N_16304,N_15985,N_15488);
and U16305 (N_16305,N_15787,N_15771);
xor U16306 (N_16306,N_15979,N_15681);
and U16307 (N_16307,N_15852,N_15727);
and U16308 (N_16308,N_15123,N_15543);
xor U16309 (N_16309,N_15279,N_15754);
nand U16310 (N_16310,N_15661,N_15428);
nor U16311 (N_16311,N_15938,N_15143);
or U16312 (N_16312,N_15407,N_15056);
xnor U16313 (N_16313,N_15531,N_15625);
and U16314 (N_16314,N_15262,N_15876);
or U16315 (N_16315,N_15851,N_15354);
nand U16316 (N_16316,N_15696,N_15829);
and U16317 (N_16317,N_15626,N_15039);
xnor U16318 (N_16318,N_15850,N_15613);
nor U16319 (N_16319,N_15303,N_15739);
and U16320 (N_16320,N_15674,N_15925);
nand U16321 (N_16321,N_15847,N_15356);
nor U16322 (N_16322,N_15540,N_15980);
and U16323 (N_16323,N_15415,N_15942);
nor U16324 (N_16324,N_15988,N_15486);
nor U16325 (N_16325,N_15744,N_15196);
and U16326 (N_16326,N_15041,N_15241);
nand U16327 (N_16327,N_15155,N_15823);
nand U16328 (N_16328,N_15566,N_15429);
and U16329 (N_16329,N_15666,N_15075);
nand U16330 (N_16330,N_15813,N_15257);
and U16331 (N_16331,N_15035,N_15672);
nand U16332 (N_16332,N_15563,N_15966);
nand U16333 (N_16333,N_15187,N_15139);
xnor U16334 (N_16334,N_15621,N_15977);
and U16335 (N_16335,N_15358,N_15635);
and U16336 (N_16336,N_15877,N_15289);
xor U16337 (N_16337,N_15761,N_15158);
nor U16338 (N_16338,N_15088,N_15816);
nor U16339 (N_16339,N_15117,N_15795);
xor U16340 (N_16340,N_15308,N_15634);
nand U16341 (N_16341,N_15609,N_15511);
and U16342 (N_16342,N_15465,N_15295);
xor U16343 (N_16343,N_15603,N_15469);
nor U16344 (N_16344,N_15788,N_15547);
nand U16345 (N_16345,N_15275,N_15596);
or U16346 (N_16346,N_15507,N_15521);
nor U16347 (N_16347,N_15961,N_15719);
or U16348 (N_16348,N_15171,N_15258);
nand U16349 (N_16349,N_15765,N_15952);
and U16350 (N_16350,N_15724,N_15255);
nand U16351 (N_16351,N_15468,N_15689);
or U16352 (N_16352,N_15481,N_15033);
xnor U16353 (N_16353,N_15145,N_15240);
or U16354 (N_16354,N_15652,N_15747);
xnor U16355 (N_16355,N_15900,N_15404);
and U16356 (N_16356,N_15610,N_15038);
nor U16357 (N_16357,N_15627,N_15055);
or U16358 (N_16358,N_15311,N_15973);
or U16359 (N_16359,N_15785,N_15214);
xnor U16360 (N_16360,N_15659,N_15050);
and U16361 (N_16361,N_15355,N_15180);
or U16362 (N_16362,N_15846,N_15002);
and U16363 (N_16363,N_15802,N_15648);
or U16364 (N_16364,N_15421,N_15363);
xor U16365 (N_16365,N_15321,N_15573);
and U16366 (N_16366,N_15114,N_15602);
nor U16367 (N_16367,N_15688,N_15514);
xor U16368 (N_16368,N_15054,N_15941);
or U16369 (N_16369,N_15220,N_15453);
and U16370 (N_16370,N_15083,N_15298);
or U16371 (N_16371,N_15040,N_15030);
or U16372 (N_16372,N_15074,N_15911);
nand U16373 (N_16373,N_15987,N_15498);
xnor U16374 (N_16374,N_15993,N_15599);
and U16375 (N_16375,N_15080,N_15178);
and U16376 (N_16376,N_15134,N_15978);
nor U16377 (N_16377,N_15028,N_15112);
nor U16378 (N_16378,N_15574,N_15529);
nand U16379 (N_16379,N_15589,N_15131);
nand U16380 (N_16380,N_15629,N_15883);
nor U16381 (N_16381,N_15108,N_15361);
xor U16382 (N_16382,N_15260,N_15662);
and U16383 (N_16383,N_15201,N_15248);
nand U16384 (N_16384,N_15528,N_15125);
xnor U16385 (N_16385,N_15317,N_15642);
xnor U16386 (N_16386,N_15159,N_15585);
xor U16387 (N_16387,N_15314,N_15591);
nand U16388 (N_16388,N_15946,N_15254);
nor U16389 (N_16389,N_15225,N_15632);
nor U16390 (N_16390,N_15833,N_15601);
nand U16391 (N_16391,N_15549,N_15950);
xnor U16392 (N_16392,N_15534,N_15960);
xor U16393 (N_16393,N_15432,N_15130);
nor U16394 (N_16394,N_15898,N_15544);
or U16395 (N_16395,N_15483,N_15077);
xnor U16396 (N_16396,N_15856,N_15711);
nand U16397 (N_16397,N_15539,N_15814);
or U16398 (N_16398,N_15205,N_15844);
nor U16399 (N_16399,N_15282,N_15575);
xnor U16400 (N_16400,N_15827,N_15043);
xor U16401 (N_16401,N_15718,N_15953);
nand U16402 (N_16402,N_15482,N_15091);
nor U16403 (N_16403,N_15693,N_15710);
xor U16404 (N_16404,N_15782,N_15052);
or U16405 (N_16405,N_15687,N_15367);
and U16406 (N_16406,N_15291,N_15745);
or U16407 (N_16407,N_15775,N_15947);
and U16408 (N_16408,N_15485,N_15261);
nor U16409 (N_16409,N_15405,N_15313);
nor U16410 (N_16410,N_15315,N_15562);
or U16411 (N_16411,N_15272,N_15956);
xor U16412 (N_16412,N_15760,N_15803);
nor U16413 (N_16413,N_15996,N_15685);
nand U16414 (N_16414,N_15700,N_15109);
and U16415 (N_16415,N_15593,N_15656);
xor U16416 (N_16416,N_15330,N_15994);
xor U16417 (N_16417,N_15643,N_15524);
and U16418 (N_16418,N_15333,N_15106);
nor U16419 (N_16419,N_15650,N_15274);
or U16420 (N_16420,N_15188,N_15427);
and U16421 (N_16421,N_15049,N_15347);
xor U16422 (N_16422,N_15455,N_15756);
nand U16423 (N_16423,N_15717,N_15414);
xor U16424 (N_16424,N_15233,N_15179);
xnor U16425 (N_16425,N_15631,N_15276);
nand U16426 (N_16426,N_15914,N_15607);
nand U16427 (N_16427,N_15786,N_15115);
and U16428 (N_16428,N_15619,N_15675);
xnor U16429 (N_16429,N_15132,N_15393);
nand U16430 (N_16430,N_15762,N_15360);
nor U16431 (N_16431,N_15763,N_15500);
or U16432 (N_16432,N_15655,N_15150);
xnor U16433 (N_16433,N_15587,N_15093);
and U16434 (N_16434,N_15237,N_15435);
and U16435 (N_16435,N_15995,N_15154);
and U16436 (N_16436,N_15858,N_15434);
or U16437 (N_16437,N_15118,N_15032);
nand U16438 (N_16438,N_15644,N_15773);
nor U16439 (N_16439,N_15678,N_15208);
xor U16440 (N_16440,N_15848,N_15228);
nand U16441 (N_16441,N_15695,N_15467);
and U16442 (N_16442,N_15394,N_15570);
and U16443 (N_16443,N_15079,N_15887);
xnor U16444 (N_16444,N_15156,N_15999);
nand U16445 (N_16445,N_15390,N_15223);
or U16446 (N_16446,N_15280,N_15398);
nand U16447 (N_16447,N_15512,N_15699);
xor U16448 (N_16448,N_15538,N_15044);
xnor U16449 (N_16449,N_15128,N_15031);
nand U16450 (N_16450,N_15001,N_15758);
or U16451 (N_16451,N_15256,N_15916);
nand U16452 (N_16452,N_15759,N_15895);
or U16453 (N_16453,N_15105,N_15310);
nand U16454 (N_16454,N_15971,N_15318);
or U16455 (N_16455,N_15669,N_15345);
xor U16456 (N_16456,N_15991,N_15920);
nand U16457 (N_16457,N_15968,N_15592);
and U16458 (N_16458,N_15658,N_15000);
or U16459 (N_16459,N_15230,N_15408);
xnor U16460 (N_16460,N_15127,N_15422);
nor U16461 (N_16461,N_15462,N_15211);
and U16462 (N_16462,N_15855,N_15300);
nor U16463 (N_16463,N_15003,N_15479);
nor U16464 (N_16464,N_15831,N_15141);
xor U16465 (N_16465,N_15584,N_15527);
nand U16466 (N_16466,N_15728,N_15292);
and U16467 (N_16467,N_15430,N_15349);
and U16468 (N_16468,N_15087,N_15783);
xnor U16469 (N_16469,N_15647,N_15057);
nand U16470 (N_16470,N_15439,N_15725);
xor U16471 (N_16471,N_15496,N_15808);
nand U16472 (N_16472,N_15184,N_15094);
nor U16473 (N_16473,N_15441,N_15378);
or U16474 (N_16474,N_15138,N_15337);
xor U16475 (N_16475,N_15764,N_15510);
nand U16476 (N_16476,N_15605,N_15182);
and U16477 (N_16477,N_15715,N_15561);
nand U16478 (N_16478,N_15385,N_15113);
nor U16479 (N_16479,N_15306,N_15342);
nand U16480 (N_16480,N_15517,N_15889);
xor U16481 (N_16481,N_15779,N_15253);
and U16482 (N_16482,N_15034,N_15072);
nor U16483 (N_16483,N_15990,N_15702);
nor U16484 (N_16484,N_15092,N_15386);
and U16485 (N_16485,N_15270,N_15062);
nand U16486 (N_16486,N_15153,N_15387);
and U16487 (N_16487,N_15668,N_15646);
nand U16488 (N_16488,N_15149,N_15567);
or U16489 (N_16489,N_15283,N_15588);
nand U16490 (N_16490,N_15677,N_15135);
or U16491 (N_16491,N_15006,N_15707);
or U16492 (N_16492,N_15849,N_15259);
nand U16493 (N_16493,N_15723,N_15506);
xnor U16494 (N_16494,N_15620,N_15250);
or U16495 (N_16495,N_15480,N_15090);
or U16496 (N_16496,N_15195,N_15922);
and U16497 (N_16497,N_15579,N_15680);
or U16498 (N_16498,N_15901,N_15921);
xor U16499 (N_16499,N_15798,N_15686);
nand U16500 (N_16500,N_15503,N_15203);
nor U16501 (N_16501,N_15502,N_15636);
and U16502 (N_16502,N_15641,N_15230);
nand U16503 (N_16503,N_15614,N_15646);
or U16504 (N_16504,N_15176,N_15476);
nand U16505 (N_16505,N_15894,N_15662);
or U16506 (N_16506,N_15998,N_15815);
xor U16507 (N_16507,N_15347,N_15737);
nand U16508 (N_16508,N_15424,N_15363);
and U16509 (N_16509,N_15333,N_15080);
nor U16510 (N_16510,N_15658,N_15006);
nor U16511 (N_16511,N_15806,N_15401);
and U16512 (N_16512,N_15348,N_15860);
and U16513 (N_16513,N_15174,N_15028);
nor U16514 (N_16514,N_15454,N_15876);
xor U16515 (N_16515,N_15535,N_15156);
nor U16516 (N_16516,N_15027,N_15456);
xor U16517 (N_16517,N_15427,N_15014);
or U16518 (N_16518,N_15395,N_15999);
or U16519 (N_16519,N_15325,N_15317);
or U16520 (N_16520,N_15752,N_15216);
nor U16521 (N_16521,N_15332,N_15518);
nor U16522 (N_16522,N_15505,N_15120);
and U16523 (N_16523,N_15902,N_15626);
nand U16524 (N_16524,N_15551,N_15697);
or U16525 (N_16525,N_15188,N_15111);
or U16526 (N_16526,N_15724,N_15207);
nand U16527 (N_16527,N_15153,N_15816);
nor U16528 (N_16528,N_15878,N_15022);
nand U16529 (N_16529,N_15546,N_15566);
xor U16530 (N_16530,N_15135,N_15213);
and U16531 (N_16531,N_15467,N_15840);
and U16532 (N_16532,N_15586,N_15431);
nand U16533 (N_16533,N_15570,N_15408);
and U16534 (N_16534,N_15906,N_15401);
or U16535 (N_16535,N_15858,N_15297);
nor U16536 (N_16536,N_15253,N_15096);
and U16537 (N_16537,N_15081,N_15370);
nor U16538 (N_16538,N_15754,N_15363);
nand U16539 (N_16539,N_15624,N_15175);
nor U16540 (N_16540,N_15388,N_15867);
nand U16541 (N_16541,N_15268,N_15574);
and U16542 (N_16542,N_15514,N_15656);
xor U16543 (N_16543,N_15845,N_15132);
nor U16544 (N_16544,N_15195,N_15889);
xor U16545 (N_16545,N_15037,N_15504);
nor U16546 (N_16546,N_15642,N_15957);
nor U16547 (N_16547,N_15947,N_15420);
nand U16548 (N_16548,N_15348,N_15117);
and U16549 (N_16549,N_15462,N_15854);
and U16550 (N_16550,N_15563,N_15324);
nor U16551 (N_16551,N_15036,N_15222);
and U16552 (N_16552,N_15721,N_15574);
and U16553 (N_16553,N_15559,N_15813);
nand U16554 (N_16554,N_15167,N_15168);
and U16555 (N_16555,N_15814,N_15028);
nor U16556 (N_16556,N_15353,N_15958);
and U16557 (N_16557,N_15060,N_15087);
nor U16558 (N_16558,N_15730,N_15359);
nor U16559 (N_16559,N_15950,N_15212);
nand U16560 (N_16560,N_15321,N_15393);
xor U16561 (N_16561,N_15995,N_15310);
nor U16562 (N_16562,N_15991,N_15450);
xnor U16563 (N_16563,N_15078,N_15418);
xor U16564 (N_16564,N_15204,N_15679);
and U16565 (N_16565,N_15510,N_15897);
nand U16566 (N_16566,N_15299,N_15706);
xor U16567 (N_16567,N_15533,N_15300);
and U16568 (N_16568,N_15638,N_15475);
nor U16569 (N_16569,N_15301,N_15105);
nor U16570 (N_16570,N_15992,N_15654);
nand U16571 (N_16571,N_15118,N_15471);
xor U16572 (N_16572,N_15030,N_15339);
and U16573 (N_16573,N_15596,N_15321);
and U16574 (N_16574,N_15283,N_15738);
or U16575 (N_16575,N_15680,N_15931);
nand U16576 (N_16576,N_15188,N_15258);
nor U16577 (N_16577,N_15326,N_15566);
xnor U16578 (N_16578,N_15730,N_15157);
xor U16579 (N_16579,N_15703,N_15277);
xor U16580 (N_16580,N_15971,N_15282);
nand U16581 (N_16581,N_15877,N_15472);
and U16582 (N_16582,N_15278,N_15061);
or U16583 (N_16583,N_15605,N_15676);
nand U16584 (N_16584,N_15823,N_15251);
or U16585 (N_16585,N_15398,N_15896);
and U16586 (N_16586,N_15471,N_15292);
nor U16587 (N_16587,N_15252,N_15395);
nand U16588 (N_16588,N_15957,N_15805);
and U16589 (N_16589,N_15696,N_15565);
xor U16590 (N_16590,N_15286,N_15736);
xnor U16591 (N_16591,N_15822,N_15199);
and U16592 (N_16592,N_15945,N_15282);
nand U16593 (N_16593,N_15042,N_15154);
nor U16594 (N_16594,N_15262,N_15614);
nor U16595 (N_16595,N_15699,N_15348);
xnor U16596 (N_16596,N_15535,N_15131);
or U16597 (N_16597,N_15759,N_15849);
nor U16598 (N_16598,N_15208,N_15025);
and U16599 (N_16599,N_15021,N_15073);
and U16600 (N_16600,N_15840,N_15168);
nand U16601 (N_16601,N_15398,N_15546);
nor U16602 (N_16602,N_15714,N_15904);
and U16603 (N_16603,N_15517,N_15419);
xor U16604 (N_16604,N_15475,N_15368);
or U16605 (N_16605,N_15264,N_15557);
nand U16606 (N_16606,N_15219,N_15745);
xnor U16607 (N_16607,N_15559,N_15296);
and U16608 (N_16608,N_15940,N_15903);
xor U16609 (N_16609,N_15357,N_15242);
xor U16610 (N_16610,N_15487,N_15189);
nand U16611 (N_16611,N_15079,N_15437);
nor U16612 (N_16612,N_15832,N_15650);
and U16613 (N_16613,N_15027,N_15921);
xnor U16614 (N_16614,N_15288,N_15190);
nor U16615 (N_16615,N_15250,N_15454);
or U16616 (N_16616,N_15028,N_15234);
and U16617 (N_16617,N_15459,N_15800);
xnor U16618 (N_16618,N_15424,N_15372);
or U16619 (N_16619,N_15419,N_15538);
xnor U16620 (N_16620,N_15619,N_15118);
nor U16621 (N_16621,N_15376,N_15293);
nor U16622 (N_16622,N_15549,N_15564);
xnor U16623 (N_16623,N_15474,N_15186);
xnor U16624 (N_16624,N_15775,N_15892);
or U16625 (N_16625,N_15284,N_15052);
and U16626 (N_16626,N_15225,N_15234);
nand U16627 (N_16627,N_15740,N_15055);
xor U16628 (N_16628,N_15391,N_15642);
and U16629 (N_16629,N_15257,N_15911);
nand U16630 (N_16630,N_15451,N_15043);
and U16631 (N_16631,N_15028,N_15382);
nor U16632 (N_16632,N_15516,N_15789);
nand U16633 (N_16633,N_15018,N_15907);
and U16634 (N_16634,N_15134,N_15794);
nand U16635 (N_16635,N_15261,N_15302);
or U16636 (N_16636,N_15307,N_15912);
nand U16637 (N_16637,N_15011,N_15853);
and U16638 (N_16638,N_15906,N_15527);
nor U16639 (N_16639,N_15243,N_15278);
nand U16640 (N_16640,N_15091,N_15414);
or U16641 (N_16641,N_15364,N_15078);
or U16642 (N_16642,N_15460,N_15356);
or U16643 (N_16643,N_15865,N_15627);
nand U16644 (N_16644,N_15943,N_15840);
nor U16645 (N_16645,N_15570,N_15521);
xnor U16646 (N_16646,N_15425,N_15106);
and U16647 (N_16647,N_15387,N_15395);
xor U16648 (N_16648,N_15013,N_15863);
and U16649 (N_16649,N_15182,N_15520);
nor U16650 (N_16650,N_15235,N_15948);
and U16651 (N_16651,N_15254,N_15016);
and U16652 (N_16652,N_15975,N_15376);
nor U16653 (N_16653,N_15355,N_15564);
nor U16654 (N_16654,N_15282,N_15782);
xor U16655 (N_16655,N_15541,N_15326);
nand U16656 (N_16656,N_15103,N_15150);
or U16657 (N_16657,N_15653,N_15393);
nand U16658 (N_16658,N_15183,N_15200);
nor U16659 (N_16659,N_15765,N_15720);
and U16660 (N_16660,N_15823,N_15069);
xnor U16661 (N_16661,N_15615,N_15016);
or U16662 (N_16662,N_15649,N_15855);
or U16663 (N_16663,N_15511,N_15526);
nor U16664 (N_16664,N_15517,N_15919);
xor U16665 (N_16665,N_15868,N_15469);
nor U16666 (N_16666,N_15109,N_15679);
or U16667 (N_16667,N_15443,N_15513);
and U16668 (N_16668,N_15196,N_15600);
and U16669 (N_16669,N_15001,N_15259);
xor U16670 (N_16670,N_15905,N_15058);
nand U16671 (N_16671,N_15061,N_15945);
nor U16672 (N_16672,N_15351,N_15457);
nor U16673 (N_16673,N_15619,N_15504);
xnor U16674 (N_16674,N_15848,N_15182);
nand U16675 (N_16675,N_15488,N_15402);
or U16676 (N_16676,N_15908,N_15368);
nor U16677 (N_16677,N_15495,N_15173);
and U16678 (N_16678,N_15956,N_15800);
xnor U16679 (N_16679,N_15174,N_15380);
xor U16680 (N_16680,N_15966,N_15482);
or U16681 (N_16681,N_15778,N_15644);
xor U16682 (N_16682,N_15748,N_15066);
xnor U16683 (N_16683,N_15047,N_15973);
or U16684 (N_16684,N_15651,N_15623);
xnor U16685 (N_16685,N_15284,N_15659);
and U16686 (N_16686,N_15341,N_15083);
nand U16687 (N_16687,N_15965,N_15391);
or U16688 (N_16688,N_15751,N_15016);
nor U16689 (N_16689,N_15455,N_15576);
or U16690 (N_16690,N_15236,N_15274);
nand U16691 (N_16691,N_15312,N_15890);
and U16692 (N_16692,N_15693,N_15914);
nand U16693 (N_16693,N_15478,N_15899);
nor U16694 (N_16694,N_15162,N_15948);
xor U16695 (N_16695,N_15604,N_15315);
nor U16696 (N_16696,N_15240,N_15163);
nand U16697 (N_16697,N_15952,N_15759);
nand U16698 (N_16698,N_15852,N_15222);
nor U16699 (N_16699,N_15352,N_15306);
or U16700 (N_16700,N_15478,N_15734);
nor U16701 (N_16701,N_15066,N_15249);
nor U16702 (N_16702,N_15516,N_15905);
and U16703 (N_16703,N_15964,N_15024);
nor U16704 (N_16704,N_15443,N_15840);
nor U16705 (N_16705,N_15868,N_15910);
nand U16706 (N_16706,N_15886,N_15045);
nor U16707 (N_16707,N_15786,N_15609);
nand U16708 (N_16708,N_15887,N_15652);
xor U16709 (N_16709,N_15884,N_15256);
nor U16710 (N_16710,N_15845,N_15286);
nand U16711 (N_16711,N_15271,N_15544);
and U16712 (N_16712,N_15213,N_15537);
and U16713 (N_16713,N_15987,N_15849);
or U16714 (N_16714,N_15631,N_15454);
or U16715 (N_16715,N_15745,N_15593);
nand U16716 (N_16716,N_15264,N_15556);
or U16717 (N_16717,N_15168,N_15748);
and U16718 (N_16718,N_15959,N_15113);
nor U16719 (N_16719,N_15573,N_15238);
xor U16720 (N_16720,N_15753,N_15425);
nand U16721 (N_16721,N_15421,N_15290);
nand U16722 (N_16722,N_15758,N_15610);
or U16723 (N_16723,N_15960,N_15380);
or U16724 (N_16724,N_15448,N_15768);
xnor U16725 (N_16725,N_15733,N_15913);
nor U16726 (N_16726,N_15126,N_15491);
xor U16727 (N_16727,N_15191,N_15745);
and U16728 (N_16728,N_15077,N_15599);
nand U16729 (N_16729,N_15706,N_15235);
nor U16730 (N_16730,N_15712,N_15661);
and U16731 (N_16731,N_15234,N_15896);
or U16732 (N_16732,N_15542,N_15302);
and U16733 (N_16733,N_15548,N_15493);
and U16734 (N_16734,N_15224,N_15770);
xnor U16735 (N_16735,N_15982,N_15219);
xor U16736 (N_16736,N_15667,N_15871);
nand U16737 (N_16737,N_15735,N_15478);
or U16738 (N_16738,N_15042,N_15288);
xor U16739 (N_16739,N_15105,N_15891);
or U16740 (N_16740,N_15561,N_15231);
xor U16741 (N_16741,N_15188,N_15933);
or U16742 (N_16742,N_15472,N_15234);
or U16743 (N_16743,N_15021,N_15538);
nor U16744 (N_16744,N_15932,N_15234);
or U16745 (N_16745,N_15832,N_15157);
nand U16746 (N_16746,N_15680,N_15752);
xor U16747 (N_16747,N_15738,N_15064);
nor U16748 (N_16748,N_15186,N_15746);
and U16749 (N_16749,N_15964,N_15488);
or U16750 (N_16750,N_15689,N_15742);
nand U16751 (N_16751,N_15282,N_15211);
nor U16752 (N_16752,N_15623,N_15078);
xor U16753 (N_16753,N_15483,N_15953);
nor U16754 (N_16754,N_15735,N_15534);
nor U16755 (N_16755,N_15762,N_15959);
and U16756 (N_16756,N_15472,N_15527);
or U16757 (N_16757,N_15869,N_15637);
nand U16758 (N_16758,N_15446,N_15734);
and U16759 (N_16759,N_15503,N_15807);
nand U16760 (N_16760,N_15018,N_15998);
and U16761 (N_16761,N_15661,N_15966);
nand U16762 (N_16762,N_15591,N_15915);
nand U16763 (N_16763,N_15996,N_15774);
and U16764 (N_16764,N_15627,N_15849);
or U16765 (N_16765,N_15654,N_15114);
nor U16766 (N_16766,N_15122,N_15354);
xor U16767 (N_16767,N_15509,N_15563);
nand U16768 (N_16768,N_15529,N_15855);
xor U16769 (N_16769,N_15865,N_15646);
nand U16770 (N_16770,N_15907,N_15815);
and U16771 (N_16771,N_15135,N_15729);
nor U16772 (N_16772,N_15031,N_15673);
or U16773 (N_16773,N_15449,N_15124);
nor U16774 (N_16774,N_15132,N_15951);
xnor U16775 (N_16775,N_15356,N_15417);
nor U16776 (N_16776,N_15813,N_15953);
xnor U16777 (N_16777,N_15428,N_15796);
and U16778 (N_16778,N_15975,N_15120);
and U16779 (N_16779,N_15098,N_15300);
nand U16780 (N_16780,N_15032,N_15568);
xnor U16781 (N_16781,N_15773,N_15293);
nor U16782 (N_16782,N_15696,N_15909);
nor U16783 (N_16783,N_15466,N_15142);
nor U16784 (N_16784,N_15093,N_15503);
and U16785 (N_16785,N_15211,N_15463);
nor U16786 (N_16786,N_15797,N_15977);
nor U16787 (N_16787,N_15898,N_15448);
nor U16788 (N_16788,N_15895,N_15082);
nor U16789 (N_16789,N_15553,N_15081);
xor U16790 (N_16790,N_15145,N_15707);
xnor U16791 (N_16791,N_15012,N_15171);
xor U16792 (N_16792,N_15780,N_15690);
nand U16793 (N_16793,N_15005,N_15812);
nor U16794 (N_16794,N_15219,N_15696);
xor U16795 (N_16795,N_15286,N_15619);
or U16796 (N_16796,N_15731,N_15138);
nor U16797 (N_16797,N_15582,N_15473);
or U16798 (N_16798,N_15689,N_15273);
and U16799 (N_16799,N_15871,N_15360);
nor U16800 (N_16800,N_15869,N_15875);
xnor U16801 (N_16801,N_15155,N_15800);
nor U16802 (N_16802,N_15320,N_15411);
nor U16803 (N_16803,N_15837,N_15868);
or U16804 (N_16804,N_15225,N_15841);
and U16805 (N_16805,N_15657,N_15974);
nor U16806 (N_16806,N_15993,N_15707);
xnor U16807 (N_16807,N_15843,N_15240);
and U16808 (N_16808,N_15683,N_15136);
xnor U16809 (N_16809,N_15189,N_15922);
or U16810 (N_16810,N_15883,N_15509);
or U16811 (N_16811,N_15749,N_15077);
and U16812 (N_16812,N_15140,N_15305);
nor U16813 (N_16813,N_15598,N_15078);
nand U16814 (N_16814,N_15961,N_15069);
or U16815 (N_16815,N_15944,N_15950);
nand U16816 (N_16816,N_15372,N_15169);
nor U16817 (N_16817,N_15911,N_15303);
nor U16818 (N_16818,N_15897,N_15010);
or U16819 (N_16819,N_15114,N_15069);
nor U16820 (N_16820,N_15635,N_15070);
nor U16821 (N_16821,N_15422,N_15983);
nor U16822 (N_16822,N_15534,N_15514);
nand U16823 (N_16823,N_15248,N_15883);
and U16824 (N_16824,N_15860,N_15750);
nor U16825 (N_16825,N_15417,N_15357);
xnor U16826 (N_16826,N_15821,N_15706);
nor U16827 (N_16827,N_15861,N_15520);
or U16828 (N_16828,N_15810,N_15221);
nand U16829 (N_16829,N_15766,N_15297);
nand U16830 (N_16830,N_15918,N_15459);
nand U16831 (N_16831,N_15616,N_15960);
nor U16832 (N_16832,N_15793,N_15764);
nor U16833 (N_16833,N_15074,N_15924);
and U16834 (N_16834,N_15064,N_15239);
and U16835 (N_16835,N_15747,N_15641);
nor U16836 (N_16836,N_15214,N_15179);
or U16837 (N_16837,N_15332,N_15022);
xnor U16838 (N_16838,N_15026,N_15066);
and U16839 (N_16839,N_15498,N_15695);
and U16840 (N_16840,N_15392,N_15964);
nand U16841 (N_16841,N_15186,N_15677);
or U16842 (N_16842,N_15091,N_15268);
xnor U16843 (N_16843,N_15726,N_15673);
nor U16844 (N_16844,N_15203,N_15033);
nand U16845 (N_16845,N_15523,N_15261);
and U16846 (N_16846,N_15113,N_15365);
or U16847 (N_16847,N_15258,N_15982);
and U16848 (N_16848,N_15510,N_15033);
xnor U16849 (N_16849,N_15312,N_15165);
xor U16850 (N_16850,N_15112,N_15356);
nand U16851 (N_16851,N_15465,N_15960);
nand U16852 (N_16852,N_15104,N_15978);
xor U16853 (N_16853,N_15159,N_15328);
nor U16854 (N_16854,N_15746,N_15893);
xor U16855 (N_16855,N_15907,N_15187);
nor U16856 (N_16856,N_15326,N_15744);
and U16857 (N_16857,N_15698,N_15781);
and U16858 (N_16858,N_15298,N_15892);
nor U16859 (N_16859,N_15144,N_15148);
nor U16860 (N_16860,N_15433,N_15229);
or U16861 (N_16861,N_15769,N_15784);
nor U16862 (N_16862,N_15766,N_15835);
or U16863 (N_16863,N_15417,N_15707);
or U16864 (N_16864,N_15051,N_15835);
nor U16865 (N_16865,N_15850,N_15857);
or U16866 (N_16866,N_15488,N_15194);
xnor U16867 (N_16867,N_15824,N_15451);
xor U16868 (N_16868,N_15206,N_15826);
nand U16869 (N_16869,N_15372,N_15787);
nor U16870 (N_16870,N_15318,N_15525);
or U16871 (N_16871,N_15083,N_15687);
xor U16872 (N_16872,N_15930,N_15877);
or U16873 (N_16873,N_15522,N_15664);
or U16874 (N_16874,N_15358,N_15274);
or U16875 (N_16875,N_15957,N_15546);
and U16876 (N_16876,N_15283,N_15057);
xnor U16877 (N_16877,N_15600,N_15939);
xor U16878 (N_16878,N_15743,N_15302);
nand U16879 (N_16879,N_15898,N_15895);
xor U16880 (N_16880,N_15570,N_15454);
nand U16881 (N_16881,N_15200,N_15570);
nor U16882 (N_16882,N_15691,N_15122);
and U16883 (N_16883,N_15334,N_15697);
or U16884 (N_16884,N_15065,N_15949);
nor U16885 (N_16885,N_15042,N_15092);
nor U16886 (N_16886,N_15253,N_15713);
and U16887 (N_16887,N_15162,N_15508);
or U16888 (N_16888,N_15784,N_15995);
and U16889 (N_16889,N_15376,N_15130);
xor U16890 (N_16890,N_15438,N_15715);
nand U16891 (N_16891,N_15106,N_15066);
nand U16892 (N_16892,N_15719,N_15156);
nor U16893 (N_16893,N_15440,N_15188);
xnor U16894 (N_16894,N_15613,N_15648);
xnor U16895 (N_16895,N_15099,N_15443);
and U16896 (N_16896,N_15466,N_15083);
and U16897 (N_16897,N_15532,N_15774);
or U16898 (N_16898,N_15345,N_15061);
and U16899 (N_16899,N_15558,N_15883);
nand U16900 (N_16900,N_15474,N_15736);
or U16901 (N_16901,N_15763,N_15446);
nor U16902 (N_16902,N_15109,N_15457);
nor U16903 (N_16903,N_15574,N_15771);
xor U16904 (N_16904,N_15945,N_15004);
nand U16905 (N_16905,N_15521,N_15574);
or U16906 (N_16906,N_15557,N_15939);
xnor U16907 (N_16907,N_15500,N_15788);
xnor U16908 (N_16908,N_15182,N_15895);
xor U16909 (N_16909,N_15147,N_15886);
or U16910 (N_16910,N_15247,N_15218);
or U16911 (N_16911,N_15094,N_15096);
xnor U16912 (N_16912,N_15896,N_15071);
xnor U16913 (N_16913,N_15539,N_15700);
nor U16914 (N_16914,N_15283,N_15944);
nor U16915 (N_16915,N_15585,N_15741);
nand U16916 (N_16916,N_15977,N_15778);
nor U16917 (N_16917,N_15103,N_15441);
xor U16918 (N_16918,N_15871,N_15496);
nand U16919 (N_16919,N_15966,N_15455);
nor U16920 (N_16920,N_15291,N_15611);
nand U16921 (N_16921,N_15545,N_15106);
and U16922 (N_16922,N_15705,N_15895);
or U16923 (N_16923,N_15223,N_15546);
and U16924 (N_16924,N_15780,N_15749);
or U16925 (N_16925,N_15482,N_15514);
xor U16926 (N_16926,N_15121,N_15075);
nand U16927 (N_16927,N_15809,N_15308);
or U16928 (N_16928,N_15370,N_15683);
nor U16929 (N_16929,N_15447,N_15838);
or U16930 (N_16930,N_15605,N_15424);
or U16931 (N_16931,N_15478,N_15894);
nand U16932 (N_16932,N_15505,N_15562);
xor U16933 (N_16933,N_15057,N_15689);
nor U16934 (N_16934,N_15916,N_15703);
and U16935 (N_16935,N_15672,N_15909);
xnor U16936 (N_16936,N_15740,N_15511);
or U16937 (N_16937,N_15724,N_15701);
nand U16938 (N_16938,N_15595,N_15361);
nor U16939 (N_16939,N_15195,N_15127);
and U16940 (N_16940,N_15663,N_15895);
or U16941 (N_16941,N_15155,N_15565);
and U16942 (N_16942,N_15967,N_15996);
and U16943 (N_16943,N_15708,N_15517);
and U16944 (N_16944,N_15505,N_15836);
and U16945 (N_16945,N_15651,N_15361);
nand U16946 (N_16946,N_15548,N_15422);
xnor U16947 (N_16947,N_15835,N_15916);
or U16948 (N_16948,N_15262,N_15816);
nand U16949 (N_16949,N_15784,N_15718);
and U16950 (N_16950,N_15119,N_15390);
and U16951 (N_16951,N_15523,N_15995);
or U16952 (N_16952,N_15776,N_15307);
nand U16953 (N_16953,N_15836,N_15266);
and U16954 (N_16954,N_15518,N_15394);
and U16955 (N_16955,N_15980,N_15841);
nor U16956 (N_16956,N_15912,N_15092);
nand U16957 (N_16957,N_15511,N_15813);
nand U16958 (N_16958,N_15678,N_15861);
xnor U16959 (N_16959,N_15959,N_15117);
nor U16960 (N_16960,N_15243,N_15468);
xnor U16961 (N_16961,N_15270,N_15297);
nand U16962 (N_16962,N_15358,N_15696);
and U16963 (N_16963,N_15749,N_15713);
and U16964 (N_16964,N_15369,N_15884);
nor U16965 (N_16965,N_15980,N_15180);
xnor U16966 (N_16966,N_15033,N_15504);
or U16967 (N_16967,N_15113,N_15739);
nand U16968 (N_16968,N_15531,N_15469);
or U16969 (N_16969,N_15782,N_15139);
xnor U16970 (N_16970,N_15753,N_15717);
xor U16971 (N_16971,N_15220,N_15025);
nand U16972 (N_16972,N_15280,N_15307);
nor U16973 (N_16973,N_15709,N_15842);
and U16974 (N_16974,N_15543,N_15296);
nand U16975 (N_16975,N_15562,N_15312);
and U16976 (N_16976,N_15679,N_15061);
and U16977 (N_16977,N_15632,N_15075);
nand U16978 (N_16978,N_15573,N_15552);
nand U16979 (N_16979,N_15570,N_15706);
or U16980 (N_16980,N_15422,N_15211);
xnor U16981 (N_16981,N_15800,N_15400);
or U16982 (N_16982,N_15493,N_15843);
xnor U16983 (N_16983,N_15801,N_15093);
and U16984 (N_16984,N_15454,N_15243);
nor U16985 (N_16985,N_15508,N_15956);
nor U16986 (N_16986,N_15255,N_15396);
nand U16987 (N_16987,N_15185,N_15480);
nor U16988 (N_16988,N_15507,N_15121);
or U16989 (N_16989,N_15763,N_15593);
xnor U16990 (N_16990,N_15745,N_15628);
and U16991 (N_16991,N_15779,N_15499);
or U16992 (N_16992,N_15298,N_15037);
nand U16993 (N_16993,N_15065,N_15989);
and U16994 (N_16994,N_15219,N_15063);
nand U16995 (N_16995,N_15366,N_15486);
nand U16996 (N_16996,N_15585,N_15623);
and U16997 (N_16997,N_15126,N_15864);
nand U16998 (N_16998,N_15082,N_15897);
nand U16999 (N_16999,N_15313,N_15063);
nand U17000 (N_17000,N_16218,N_16204);
or U17001 (N_17001,N_16952,N_16456);
nand U17002 (N_17002,N_16405,N_16416);
nand U17003 (N_17003,N_16347,N_16447);
nand U17004 (N_17004,N_16052,N_16958);
nor U17005 (N_17005,N_16449,N_16384);
or U17006 (N_17006,N_16138,N_16589);
xnor U17007 (N_17007,N_16834,N_16763);
or U17008 (N_17008,N_16974,N_16616);
xnor U17009 (N_17009,N_16503,N_16788);
nor U17010 (N_17010,N_16119,N_16284);
or U17011 (N_17011,N_16376,N_16812);
xnor U17012 (N_17012,N_16082,N_16646);
and U17013 (N_17013,N_16977,N_16723);
nand U17014 (N_17014,N_16028,N_16269);
and U17015 (N_17015,N_16422,N_16427);
nor U17016 (N_17016,N_16051,N_16315);
nand U17017 (N_17017,N_16483,N_16077);
xnor U17018 (N_17018,N_16897,N_16963);
xnor U17019 (N_17019,N_16467,N_16957);
xor U17020 (N_17020,N_16001,N_16608);
or U17021 (N_17021,N_16990,N_16671);
nand U17022 (N_17022,N_16452,N_16828);
or U17023 (N_17023,N_16967,N_16872);
xor U17024 (N_17024,N_16355,N_16264);
or U17025 (N_17025,N_16968,N_16471);
and U17026 (N_17026,N_16124,N_16970);
nor U17027 (N_17027,N_16742,N_16036);
or U17028 (N_17028,N_16078,N_16314);
and U17029 (N_17029,N_16281,N_16691);
or U17030 (N_17030,N_16705,N_16604);
xnor U17031 (N_17031,N_16749,N_16819);
and U17032 (N_17032,N_16121,N_16437);
or U17033 (N_17033,N_16701,N_16510);
and U17034 (N_17034,N_16986,N_16032);
or U17035 (N_17035,N_16876,N_16889);
and U17036 (N_17036,N_16368,N_16141);
and U17037 (N_17037,N_16087,N_16213);
and U17038 (N_17038,N_16855,N_16938);
nand U17039 (N_17039,N_16666,N_16794);
or U17040 (N_17040,N_16267,N_16606);
and U17041 (N_17041,N_16283,N_16319);
nor U17042 (N_17042,N_16707,N_16853);
xnor U17043 (N_17043,N_16445,N_16307);
or U17044 (N_17044,N_16410,N_16475);
and U17045 (N_17045,N_16115,N_16392);
nor U17046 (N_17046,N_16219,N_16557);
and U17047 (N_17047,N_16507,N_16680);
xnor U17048 (N_17048,N_16192,N_16837);
nor U17049 (N_17049,N_16060,N_16620);
xnor U17050 (N_17050,N_16223,N_16665);
xor U17051 (N_17051,N_16401,N_16132);
or U17052 (N_17052,N_16360,N_16173);
or U17053 (N_17053,N_16694,N_16506);
nand U17054 (N_17054,N_16708,N_16029);
xor U17055 (N_17055,N_16913,N_16956);
or U17056 (N_17056,N_16790,N_16209);
or U17057 (N_17057,N_16594,N_16585);
or U17058 (N_17058,N_16830,N_16048);
nor U17059 (N_17059,N_16961,N_16715);
nand U17060 (N_17060,N_16389,N_16193);
xor U17061 (N_17061,N_16260,N_16972);
xor U17062 (N_17062,N_16524,N_16271);
nand U17063 (N_17063,N_16408,N_16817);
nor U17064 (N_17064,N_16917,N_16764);
xor U17065 (N_17065,N_16710,N_16745);
and U17066 (N_17066,N_16272,N_16296);
xnor U17067 (N_17067,N_16748,N_16374);
nor U17068 (N_17068,N_16909,N_16292);
xor U17069 (N_17069,N_16241,N_16380);
and U17070 (N_17070,N_16540,N_16664);
or U17071 (N_17071,N_16020,N_16814);
or U17072 (N_17072,N_16547,N_16933);
or U17073 (N_17073,N_16796,N_16211);
and U17074 (N_17074,N_16751,N_16560);
nand U17075 (N_17075,N_16326,N_16424);
nand U17076 (N_17076,N_16623,N_16139);
or U17077 (N_17077,N_16041,N_16308);
and U17078 (N_17078,N_16976,N_16120);
nand U17079 (N_17079,N_16182,N_16852);
or U17080 (N_17080,N_16572,N_16638);
or U17081 (N_17081,N_16378,N_16239);
xor U17082 (N_17082,N_16780,N_16562);
nor U17083 (N_17083,N_16233,N_16692);
xor U17084 (N_17084,N_16716,N_16131);
or U17085 (N_17085,N_16777,N_16699);
and U17086 (N_17086,N_16720,N_16373);
nor U17087 (N_17087,N_16109,N_16215);
xor U17088 (N_17088,N_16482,N_16366);
nand U17089 (N_17089,N_16655,N_16190);
nand U17090 (N_17090,N_16181,N_16712);
or U17091 (N_17091,N_16058,N_16871);
nand U17092 (N_17092,N_16302,N_16243);
or U17093 (N_17093,N_16300,N_16662);
and U17094 (N_17094,N_16561,N_16174);
and U17095 (N_17095,N_16653,N_16248);
or U17096 (N_17096,N_16912,N_16275);
nor U17097 (N_17097,N_16240,N_16188);
and U17098 (N_17098,N_16153,N_16186);
xor U17099 (N_17099,N_16971,N_16110);
and U17100 (N_17100,N_16929,N_16630);
nor U17101 (N_17101,N_16394,N_16808);
and U17102 (N_17102,N_16914,N_16464);
xor U17103 (N_17103,N_16667,N_16989);
nand U17104 (N_17104,N_16327,N_16840);
nand U17105 (N_17105,N_16943,N_16688);
and U17106 (N_17106,N_16417,N_16455);
or U17107 (N_17107,N_16516,N_16866);
and U17108 (N_17108,N_16448,N_16125);
or U17109 (N_17109,N_16579,N_16799);
or U17110 (N_17110,N_16532,N_16760);
nand U17111 (N_17111,N_16290,N_16045);
or U17112 (N_17112,N_16884,N_16839);
xnor U17113 (N_17113,N_16757,N_16823);
nand U17114 (N_17114,N_16157,N_16461);
and U17115 (N_17115,N_16672,N_16316);
xor U17116 (N_17116,N_16322,N_16928);
and U17117 (N_17117,N_16979,N_16862);
or U17118 (N_17118,N_16249,N_16253);
xnor U17119 (N_17119,N_16856,N_16642);
nor U17120 (N_17120,N_16854,N_16199);
nand U17121 (N_17121,N_16273,N_16194);
nor U17122 (N_17122,N_16878,N_16346);
nand U17123 (N_17123,N_16544,N_16252);
or U17124 (N_17124,N_16183,N_16877);
nor U17125 (N_17125,N_16263,N_16987);
nor U17126 (N_17126,N_16033,N_16896);
or U17127 (N_17127,N_16578,N_16534);
nand U17128 (N_17128,N_16743,N_16729);
nand U17129 (N_17129,N_16126,N_16538);
and U17130 (N_17130,N_16064,N_16010);
or U17131 (N_17131,N_16205,N_16421);
nand U17132 (N_17132,N_16577,N_16221);
nor U17133 (N_17133,N_16166,N_16683);
nand U17134 (N_17134,N_16413,N_16758);
and U17135 (N_17135,N_16053,N_16009);
nand U17136 (N_17136,N_16558,N_16684);
nand U17137 (N_17137,N_16719,N_16093);
xnor U17138 (N_17138,N_16140,N_16744);
xnor U17139 (N_17139,N_16442,N_16108);
and U17140 (N_17140,N_16031,N_16004);
nor U17141 (N_17141,N_16658,N_16288);
nand U17142 (N_17142,N_16874,N_16614);
xor U17143 (N_17143,N_16724,N_16295);
and U17144 (N_17144,N_16945,N_16016);
nor U17145 (N_17145,N_16717,N_16930);
and U17146 (N_17146,N_16737,N_16160);
nor U17147 (N_17147,N_16399,N_16600);
nand U17148 (N_17148,N_16820,N_16918);
nor U17149 (N_17149,N_16202,N_16921);
and U17150 (N_17150,N_16593,N_16795);
and U17151 (N_17151,N_16821,N_16761);
and U17152 (N_17152,N_16244,N_16697);
and U17153 (N_17153,N_16497,N_16505);
nor U17154 (N_17154,N_16739,N_16387);
or U17155 (N_17155,N_16407,N_16008);
xnor U17156 (N_17156,N_16675,N_16881);
or U17157 (N_17157,N_16756,N_16229);
xnor U17158 (N_17158,N_16135,N_16677);
nand U17159 (N_17159,N_16539,N_16640);
and U17160 (N_17160,N_16172,N_16398);
nor U17161 (N_17161,N_16074,N_16321);
nor U17162 (N_17162,N_16887,N_16245);
nor U17163 (N_17163,N_16545,N_16559);
nand U17164 (N_17164,N_16342,N_16338);
xnor U17165 (N_17165,N_16863,N_16364);
xor U17166 (N_17166,N_16668,N_16474);
nand U17167 (N_17167,N_16083,N_16354);
nand U17168 (N_17168,N_16893,N_16792);
nor U17169 (N_17169,N_16353,N_16454);
and U17170 (N_17170,N_16294,N_16673);
or U17171 (N_17171,N_16868,N_16017);
or U17172 (N_17172,N_16280,N_16491);
xor U17173 (N_17173,N_16002,N_16522);
xnor U17174 (N_17174,N_16580,N_16007);
nand U17175 (N_17175,N_16065,N_16509);
nor U17176 (N_17176,N_16303,N_16944);
nor U17177 (N_17177,N_16605,N_16514);
or U17178 (N_17178,N_16627,N_16768);
nor U17179 (N_17179,N_16340,N_16098);
nand U17180 (N_17180,N_16320,N_16328);
xnor U17181 (N_17181,N_16512,N_16428);
and U17182 (N_17182,N_16695,N_16992);
or U17183 (N_17183,N_16994,N_16885);
nor U17184 (N_17184,N_16235,N_16335);
nor U17185 (N_17185,N_16528,N_16836);
nand U17186 (N_17186,N_16966,N_16349);
xnor U17187 (N_17187,N_16311,N_16412);
and U17188 (N_17188,N_16013,N_16494);
or U17189 (N_17189,N_16450,N_16576);
xor U17190 (N_17190,N_16791,N_16116);
nand U17191 (N_17191,N_16479,N_16582);
or U17192 (N_17192,N_16525,N_16753);
nand U17193 (N_17193,N_16624,N_16439);
or U17194 (N_17194,N_16713,N_16693);
or U17195 (N_17195,N_16238,N_16548);
and U17196 (N_17196,N_16750,N_16489);
or U17197 (N_17197,N_16148,N_16037);
and U17198 (N_17198,N_16403,N_16067);
xnor U17199 (N_17199,N_16214,N_16341);
xor U17200 (N_17200,N_16568,N_16983);
xor U17201 (N_17201,N_16434,N_16324);
nand U17202 (N_17202,N_16282,N_16180);
xor U17203 (N_17203,N_16091,N_16021);
nand U17204 (N_17204,N_16325,N_16076);
or U17205 (N_17205,N_16167,N_16459);
nor U17206 (N_17206,N_16847,N_16681);
and U17207 (N_17207,N_16826,N_16833);
and U17208 (N_17208,N_16895,N_16230);
or U17209 (N_17209,N_16487,N_16019);
xnor U17210 (N_17210,N_16152,N_16554);
or U17211 (N_17211,N_16513,N_16099);
nand U17212 (N_17212,N_16102,N_16922);
or U17213 (N_17213,N_16185,N_16546);
and U17214 (N_17214,N_16636,N_16089);
xnor U17215 (N_17215,N_16179,N_16904);
xor U17216 (N_17216,N_16573,N_16363);
or U17217 (N_17217,N_16197,N_16969);
nor U17218 (N_17218,N_16552,N_16553);
nand U17219 (N_17219,N_16344,N_16873);
or U17220 (N_17220,N_16330,N_16187);
nand U17221 (N_17221,N_16414,N_16888);
or U17222 (N_17222,N_16551,N_16998);
nand U17223 (N_17223,N_16923,N_16703);
nand U17224 (N_17224,N_16845,N_16436);
and U17225 (N_17225,N_16476,N_16648);
and U17226 (N_17226,N_16469,N_16163);
xor U17227 (N_17227,N_16372,N_16962);
nand U17228 (N_17228,N_16822,N_16732);
or U17229 (N_17229,N_16784,N_16257);
or U17230 (N_17230,N_16515,N_16440);
and U17231 (N_17231,N_16113,N_16687);
and U17232 (N_17232,N_16850,N_16156);
xnor U17233 (N_17233,N_16619,N_16597);
xor U17234 (N_17234,N_16429,N_16332);
and U17235 (N_17235,N_16674,N_16143);
or U17236 (N_17236,N_16925,N_16468);
nand U17237 (N_17237,N_16523,N_16838);
nand U17238 (N_17238,N_16285,N_16015);
xnor U17239 (N_17239,N_16886,N_16438);
or U17240 (N_17240,N_16189,N_16498);
or U17241 (N_17241,N_16669,N_16988);
and U17242 (N_17242,N_16499,N_16207);
nor U17243 (N_17243,N_16869,N_16406);
nor U17244 (N_17244,N_16607,N_16859);
nand U17245 (N_17245,N_16656,N_16359);
or U17246 (N_17246,N_16396,N_16385);
nor U17247 (N_17247,N_16985,N_16334);
xor U17248 (N_17248,N_16536,N_16256);
nor U17249 (N_17249,N_16261,N_16905);
nand U17250 (N_17250,N_16870,N_16081);
xor U17251 (N_17251,N_16150,N_16789);
and U17252 (N_17252,N_16493,N_16305);
nand U17253 (N_17253,N_16206,N_16208);
or U17254 (N_17254,N_16916,N_16195);
xnor U17255 (N_17255,N_16782,N_16411);
or U17256 (N_17256,N_16637,N_16049);
or U17257 (N_17257,N_16073,N_16776);
or U17258 (N_17258,N_16829,N_16457);
or U17259 (N_17259,N_16220,N_16920);
and U17260 (N_17260,N_16706,N_16430);
nor U17261 (N_17261,N_16178,N_16095);
nor U17262 (N_17262,N_16085,N_16234);
or U17263 (N_17263,N_16331,N_16841);
nor U17264 (N_17264,N_16151,N_16741);
and U17265 (N_17265,N_16170,N_16463);
xor U17266 (N_17266,N_16265,N_16766);
or U17267 (N_17267,N_16798,N_16955);
and U17268 (N_17268,N_16390,N_16993);
or U17269 (N_17269,N_16317,N_16023);
nor U17270 (N_17270,N_16875,N_16114);
and U17271 (N_17271,N_16995,N_16042);
nor U17272 (N_17272,N_16611,N_16891);
nor U17273 (N_17273,N_16415,N_16480);
nor U17274 (N_17274,N_16982,N_16907);
or U17275 (N_17275,N_16954,N_16906);
or U17276 (N_17276,N_16274,N_16803);
nor U17277 (N_17277,N_16084,N_16090);
xnor U17278 (N_17278,N_16569,N_16236);
xnor U17279 (N_17279,N_16381,N_16079);
xor U17280 (N_17280,N_16367,N_16949);
or U17281 (N_17281,N_16043,N_16062);
nor U17282 (N_17282,N_16654,N_16631);
and U17283 (N_17283,N_16472,N_16104);
nor U17284 (N_17284,N_16086,N_16588);
and U17285 (N_17285,N_16386,N_16947);
nor U17286 (N_17286,N_16861,N_16420);
or U17287 (N_17287,N_16289,N_16939);
and U17288 (N_17288,N_16504,N_16329);
and U17289 (N_17289,N_16556,N_16910);
xnor U17290 (N_17290,N_16778,N_16298);
or U17291 (N_17291,N_16807,N_16634);
xnor U17292 (N_17292,N_16809,N_16915);
nor U17293 (N_17293,N_16787,N_16129);
and U17294 (N_17294,N_16158,N_16621);
or U17295 (N_17295,N_16639,N_16232);
or U17296 (N_17296,N_16980,N_16397);
and U17297 (N_17297,N_16356,N_16530);
xnor U17298 (N_17298,N_16747,N_16520);
or U17299 (N_17299,N_16825,N_16867);
nand U17300 (N_17300,N_16304,N_16164);
nor U17301 (N_17301,N_16375,N_16835);
nand U17302 (N_17302,N_16996,N_16728);
nor U17303 (N_17303,N_16286,N_16130);
nand U17304 (N_17304,N_16337,N_16844);
or U17305 (N_17305,N_16709,N_16670);
and U17306 (N_17306,N_16477,N_16950);
xor U17307 (N_17307,N_16254,N_16883);
and U17308 (N_17308,N_16643,N_16924);
or U17309 (N_17309,N_16927,N_16258);
xnor U17310 (N_17310,N_16702,N_16801);
and U17311 (N_17311,N_16860,N_16301);
and U17312 (N_17312,N_16571,N_16134);
or U17313 (N_17313,N_16566,N_16981);
or U17314 (N_17314,N_16740,N_16343);
or U17315 (N_17315,N_16946,N_16024);
nand U17316 (N_17316,N_16805,N_16210);
xnor U17317 (N_17317,N_16765,N_16657);
or U17318 (N_17318,N_16779,N_16583);
xnor U17319 (N_17319,N_16690,N_16849);
nand U17320 (N_17320,N_16492,N_16899);
xnor U17321 (N_17321,N_16435,N_16072);
and U17322 (N_17322,N_16149,N_16632);
nand U17323 (N_17323,N_16775,N_16118);
nor U17324 (N_17324,N_16644,N_16112);
or U17325 (N_17325,N_16615,N_16660);
nand U17326 (N_17326,N_16926,N_16061);
nor U17327 (N_17327,N_16773,N_16419);
nor U17328 (N_17328,N_16537,N_16266);
nor U17329 (N_17329,N_16804,N_16810);
nor U17330 (N_17330,N_16470,N_16942);
or U17331 (N_17331,N_16997,N_16973);
nand U17332 (N_17332,N_16678,N_16940);
or U17333 (N_17333,N_16395,N_16460);
nand U17334 (N_17334,N_16919,N_16984);
xor U17335 (N_17335,N_16858,N_16542);
nor U17336 (N_17336,N_16738,N_16071);
xor U17337 (N_17337,N_16581,N_16184);
or U17338 (N_17338,N_16641,N_16391);
and U17339 (N_17339,N_16313,N_16352);
nor U17340 (N_17340,N_16519,N_16000);
or U17341 (N_17341,N_16857,N_16345);
nand U17342 (N_17342,N_16293,N_16894);
and U17343 (N_17343,N_16793,N_16865);
and U17344 (N_17344,N_16200,N_16890);
or U17345 (N_17345,N_16030,N_16733);
nor U17346 (N_17346,N_16698,N_16441);
nor U17347 (N_17347,N_16934,N_16685);
nand U17348 (N_17348,N_16177,N_16932);
or U17349 (N_17349,N_16370,N_16018);
and U17350 (N_17350,N_16831,N_16903);
xnor U17351 (N_17351,N_16591,N_16953);
or U17352 (N_17352,N_16451,N_16550);
and U17353 (N_17353,N_16046,N_16203);
and U17354 (N_17354,N_16633,N_16222);
nand U17355 (N_17355,N_16570,N_16056);
nor U17356 (N_17356,N_16357,N_16565);
xor U17357 (N_17357,N_16502,N_16650);
nor U17358 (N_17358,N_16549,N_16911);
and U17359 (N_17359,N_16609,N_16055);
xor U17360 (N_17360,N_16689,N_16100);
and U17361 (N_17361,N_16722,N_16726);
or U17362 (N_17362,N_16526,N_16892);
nand U17363 (N_17363,N_16022,N_16225);
nor U17364 (N_17364,N_16059,N_16746);
or U17365 (N_17365,N_16659,N_16767);
nand U17366 (N_17366,N_16312,N_16122);
nor U17367 (N_17367,N_16543,N_16711);
nand U17368 (N_17368,N_16527,N_16882);
nand U17369 (N_17369,N_16161,N_16276);
or U17370 (N_17370,N_16069,N_16299);
nand U17371 (N_17371,N_16661,N_16700);
nand U17372 (N_17372,N_16466,N_16704);
xor U17373 (N_17373,N_16774,N_16811);
nand U17374 (N_17374,N_16409,N_16769);
and U17375 (N_17375,N_16418,N_16369);
nand U17376 (N_17376,N_16402,N_16165);
and U17377 (N_17377,N_16101,N_16517);
nor U17378 (N_17378,N_16226,N_16306);
or U17379 (N_17379,N_16975,N_16171);
and U17380 (N_17380,N_16495,N_16626);
or U17381 (N_17381,N_16142,N_16842);
or U17382 (N_17382,N_16005,N_16908);
xor U17383 (N_17383,N_16679,N_16066);
and U17384 (N_17384,N_16237,N_16951);
or U17385 (N_17385,N_16960,N_16851);
and U17386 (N_17386,N_16377,N_16755);
nand U17387 (N_17387,N_16730,N_16006);
nand U17388 (N_17388,N_16846,N_16880);
and U17389 (N_17389,N_16590,N_16057);
nor U17390 (N_17390,N_16898,N_16270);
nor U17391 (N_17391,N_16106,N_16754);
nor U17392 (N_17392,N_16529,N_16484);
and U17393 (N_17393,N_16040,N_16535);
nor U17394 (N_17394,N_16014,N_16128);
or U17395 (N_17395,N_16478,N_16937);
or U17396 (N_17396,N_16598,N_16848);
and U17397 (N_17397,N_16382,N_16635);
and U17398 (N_17398,N_16843,N_16255);
and U17399 (N_17399,N_16191,N_16063);
or U17400 (N_17400,N_16941,N_16473);
and U17401 (N_17401,N_16278,N_16025);
and U17402 (N_17402,N_16596,N_16433);
and U17403 (N_17403,N_16800,N_16175);
or U17404 (N_17404,N_16383,N_16117);
xor U17405 (N_17405,N_16388,N_16291);
nand U17406 (N_17406,N_16146,N_16080);
nor U17407 (N_17407,N_16511,N_16246);
nor U17408 (N_17408,N_16123,N_16521);
xnor U17409 (N_17409,N_16242,N_16423);
or U17410 (N_17410,N_16196,N_16358);
and U17411 (N_17411,N_16169,N_16771);
nand U17412 (N_17412,N_16462,N_16277);
nor U17413 (N_17413,N_16431,N_16959);
nand U17414 (N_17414,N_16361,N_16797);
xnor U17415 (N_17415,N_16400,N_16617);
nand U17416 (N_17416,N_16287,N_16718);
or U17417 (N_17417,N_16647,N_16147);
nor U17418 (N_17418,N_16518,N_16628);
or U17419 (N_17419,N_16612,N_16268);
xor U17420 (N_17420,N_16759,N_16592);
and U17421 (N_17421,N_16879,N_16154);
nand U17422 (N_17422,N_16563,N_16145);
nand U17423 (N_17423,N_16575,N_16444);
nand U17424 (N_17424,N_16541,N_16336);
nor U17425 (N_17425,N_16155,N_16070);
nor U17426 (N_17426,N_16198,N_16935);
nand U17427 (N_17427,N_16772,N_16649);
or U17428 (N_17428,N_16133,N_16651);
and U17429 (N_17429,N_16603,N_16618);
nand U17430 (N_17430,N_16027,N_16323);
xor U17431 (N_17431,N_16816,N_16054);
nand U17432 (N_17432,N_16490,N_16310);
nor U17433 (N_17433,N_16228,N_16734);
xor U17434 (N_17434,N_16555,N_16813);
and U17435 (N_17435,N_16144,N_16901);
nand U17436 (N_17436,N_16465,N_16224);
nand U17437 (N_17437,N_16047,N_16500);
xnor U17438 (N_17438,N_16786,N_16318);
or U17439 (N_17439,N_16075,N_16103);
or U17440 (N_17440,N_16610,N_16365);
and U17441 (N_17441,N_16625,N_16613);
nor U17442 (N_17442,N_16348,N_16931);
xnor U17443 (N_17443,N_16964,N_16725);
and U17444 (N_17444,N_16567,N_16279);
and U17445 (N_17445,N_16531,N_16574);
or U17446 (N_17446,N_16991,N_16486);
and U17447 (N_17447,N_16035,N_16231);
nor U17448 (N_17448,N_16736,N_16050);
nand U17449 (N_17449,N_16026,N_16379);
nand U17450 (N_17450,N_16251,N_16762);
and U17451 (N_17451,N_16068,N_16508);
xnor U17452 (N_17452,N_16393,N_16136);
and U17453 (N_17453,N_16111,N_16629);
nor U17454 (N_17454,N_16105,N_16351);
xor U17455 (N_17455,N_16092,N_16564);
and U17456 (N_17456,N_16731,N_16501);
nor U17457 (N_17457,N_16696,N_16012);
and U17458 (N_17458,N_16011,N_16587);
nand U17459 (N_17459,N_16770,N_16443);
xor U17460 (N_17460,N_16721,N_16586);
nor U17461 (N_17461,N_16362,N_16802);
and U17462 (N_17462,N_16827,N_16978);
and U17463 (N_17463,N_16965,N_16262);
nand U17464 (N_17464,N_16339,N_16622);
and U17465 (N_17465,N_16727,N_16097);
and U17466 (N_17466,N_16864,N_16247);
nand U17467 (N_17467,N_16815,N_16003);
nand U17468 (N_17468,N_16107,N_16259);
and U17469 (N_17469,N_16039,N_16682);
and U17470 (N_17470,N_16432,N_16663);
and U17471 (N_17471,N_16496,N_16350);
nor U17472 (N_17472,N_16752,N_16137);
and U17473 (N_17473,N_16217,N_16425);
nor U17474 (N_17474,N_16481,N_16212);
and U17475 (N_17475,N_16806,N_16601);
or U17476 (N_17476,N_16088,N_16686);
or U17477 (N_17477,N_16446,N_16948);
and U17478 (N_17478,N_16645,N_16902);
nand U17479 (N_17479,N_16785,N_16584);
or U17480 (N_17480,N_16781,N_16227);
xnor U17481 (N_17481,N_16533,N_16297);
xnor U17482 (N_17482,N_16458,N_16488);
xnor U17483 (N_17483,N_16453,N_16333);
or U17484 (N_17484,N_16832,N_16159);
or U17485 (N_17485,N_16595,N_16096);
nand U17486 (N_17486,N_16714,N_16309);
or U17487 (N_17487,N_16168,N_16602);
nor U17488 (N_17488,N_16676,N_16127);
and U17489 (N_17489,N_16034,N_16824);
or U17490 (N_17490,N_16936,N_16216);
and U17491 (N_17491,N_16094,N_16735);
or U17492 (N_17492,N_16044,N_16652);
or U17493 (N_17493,N_16999,N_16900);
and U17494 (N_17494,N_16250,N_16783);
or U17495 (N_17495,N_16485,N_16162);
xnor U17496 (N_17496,N_16201,N_16426);
nand U17497 (N_17497,N_16404,N_16038);
nand U17498 (N_17498,N_16599,N_16371);
xnor U17499 (N_17499,N_16176,N_16818);
or U17500 (N_17500,N_16046,N_16037);
nor U17501 (N_17501,N_16475,N_16441);
and U17502 (N_17502,N_16121,N_16806);
or U17503 (N_17503,N_16397,N_16744);
and U17504 (N_17504,N_16954,N_16386);
nand U17505 (N_17505,N_16272,N_16946);
nand U17506 (N_17506,N_16440,N_16343);
xor U17507 (N_17507,N_16724,N_16111);
and U17508 (N_17508,N_16653,N_16920);
and U17509 (N_17509,N_16226,N_16389);
nand U17510 (N_17510,N_16356,N_16347);
nor U17511 (N_17511,N_16569,N_16852);
nand U17512 (N_17512,N_16794,N_16089);
nor U17513 (N_17513,N_16194,N_16157);
nor U17514 (N_17514,N_16550,N_16365);
nand U17515 (N_17515,N_16790,N_16237);
nor U17516 (N_17516,N_16914,N_16382);
xor U17517 (N_17517,N_16291,N_16115);
and U17518 (N_17518,N_16999,N_16585);
nor U17519 (N_17519,N_16797,N_16494);
and U17520 (N_17520,N_16470,N_16202);
or U17521 (N_17521,N_16243,N_16331);
xnor U17522 (N_17522,N_16177,N_16027);
nor U17523 (N_17523,N_16677,N_16221);
and U17524 (N_17524,N_16904,N_16892);
and U17525 (N_17525,N_16557,N_16759);
or U17526 (N_17526,N_16045,N_16832);
xor U17527 (N_17527,N_16015,N_16501);
or U17528 (N_17528,N_16053,N_16241);
nand U17529 (N_17529,N_16957,N_16985);
nor U17530 (N_17530,N_16749,N_16585);
nand U17531 (N_17531,N_16240,N_16172);
nor U17532 (N_17532,N_16879,N_16331);
or U17533 (N_17533,N_16618,N_16329);
or U17534 (N_17534,N_16696,N_16663);
or U17535 (N_17535,N_16337,N_16116);
or U17536 (N_17536,N_16272,N_16112);
xnor U17537 (N_17537,N_16182,N_16803);
nor U17538 (N_17538,N_16673,N_16898);
nand U17539 (N_17539,N_16871,N_16360);
xnor U17540 (N_17540,N_16917,N_16980);
or U17541 (N_17541,N_16404,N_16373);
xnor U17542 (N_17542,N_16167,N_16601);
xnor U17543 (N_17543,N_16909,N_16496);
xor U17544 (N_17544,N_16216,N_16928);
nand U17545 (N_17545,N_16134,N_16052);
and U17546 (N_17546,N_16809,N_16001);
and U17547 (N_17547,N_16667,N_16140);
or U17548 (N_17548,N_16075,N_16691);
nor U17549 (N_17549,N_16248,N_16953);
and U17550 (N_17550,N_16367,N_16478);
xor U17551 (N_17551,N_16218,N_16371);
or U17552 (N_17552,N_16182,N_16217);
and U17553 (N_17553,N_16567,N_16873);
and U17554 (N_17554,N_16273,N_16632);
or U17555 (N_17555,N_16007,N_16637);
and U17556 (N_17556,N_16639,N_16641);
and U17557 (N_17557,N_16669,N_16408);
nor U17558 (N_17558,N_16732,N_16555);
or U17559 (N_17559,N_16703,N_16403);
or U17560 (N_17560,N_16485,N_16208);
xnor U17561 (N_17561,N_16101,N_16258);
nor U17562 (N_17562,N_16129,N_16226);
and U17563 (N_17563,N_16335,N_16901);
or U17564 (N_17564,N_16232,N_16924);
and U17565 (N_17565,N_16981,N_16905);
or U17566 (N_17566,N_16696,N_16389);
nand U17567 (N_17567,N_16875,N_16985);
xor U17568 (N_17568,N_16657,N_16649);
nand U17569 (N_17569,N_16275,N_16157);
nor U17570 (N_17570,N_16249,N_16383);
xor U17571 (N_17571,N_16466,N_16788);
nand U17572 (N_17572,N_16148,N_16940);
and U17573 (N_17573,N_16806,N_16781);
or U17574 (N_17574,N_16606,N_16097);
nand U17575 (N_17575,N_16851,N_16162);
xor U17576 (N_17576,N_16810,N_16628);
nand U17577 (N_17577,N_16112,N_16831);
nand U17578 (N_17578,N_16710,N_16307);
and U17579 (N_17579,N_16288,N_16425);
or U17580 (N_17580,N_16987,N_16470);
nor U17581 (N_17581,N_16587,N_16111);
nand U17582 (N_17582,N_16183,N_16623);
xor U17583 (N_17583,N_16288,N_16480);
or U17584 (N_17584,N_16307,N_16098);
nand U17585 (N_17585,N_16403,N_16699);
nor U17586 (N_17586,N_16423,N_16686);
nand U17587 (N_17587,N_16421,N_16166);
and U17588 (N_17588,N_16728,N_16568);
xor U17589 (N_17589,N_16015,N_16355);
and U17590 (N_17590,N_16703,N_16015);
and U17591 (N_17591,N_16727,N_16442);
and U17592 (N_17592,N_16284,N_16718);
or U17593 (N_17593,N_16720,N_16223);
nand U17594 (N_17594,N_16964,N_16928);
nand U17595 (N_17595,N_16832,N_16931);
xnor U17596 (N_17596,N_16299,N_16463);
nor U17597 (N_17597,N_16963,N_16153);
and U17598 (N_17598,N_16752,N_16459);
or U17599 (N_17599,N_16427,N_16005);
nor U17600 (N_17600,N_16934,N_16393);
nand U17601 (N_17601,N_16970,N_16945);
nor U17602 (N_17602,N_16363,N_16219);
and U17603 (N_17603,N_16709,N_16269);
nor U17604 (N_17604,N_16835,N_16590);
and U17605 (N_17605,N_16809,N_16666);
nand U17606 (N_17606,N_16406,N_16970);
xnor U17607 (N_17607,N_16492,N_16545);
xnor U17608 (N_17608,N_16262,N_16120);
or U17609 (N_17609,N_16954,N_16057);
or U17610 (N_17610,N_16872,N_16508);
and U17611 (N_17611,N_16551,N_16710);
xor U17612 (N_17612,N_16598,N_16277);
or U17613 (N_17613,N_16439,N_16852);
and U17614 (N_17614,N_16176,N_16923);
or U17615 (N_17615,N_16757,N_16755);
and U17616 (N_17616,N_16211,N_16941);
nand U17617 (N_17617,N_16570,N_16745);
nand U17618 (N_17618,N_16293,N_16851);
nor U17619 (N_17619,N_16081,N_16985);
nor U17620 (N_17620,N_16801,N_16327);
or U17621 (N_17621,N_16380,N_16775);
nand U17622 (N_17622,N_16019,N_16466);
or U17623 (N_17623,N_16055,N_16762);
and U17624 (N_17624,N_16172,N_16122);
and U17625 (N_17625,N_16890,N_16526);
nor U17626 (N_17626,N_16472,N_16436);
and U17627 (N_17627,N_16997,N_16578);
xor U17628 (N_17628,N_16816,N_16836);
nand U17629 (N_17629,N_16790,N_16823);
xor U17630 (N_17630,N_16039,N_16845);
nand U17631 (N_17631,N_16609,N_16710);
nor U17632 (N_17632,N_16051,N_16879);
xor U17633 (N_17633,N_16847,N_16599);
xnor U17634 (N_17634,N_16061,N_16247);
nand U17635 (N_17635,N_16132,N_16256);
xor U17636 (N_17636,N_16398,N_16592);
or U17637 (N_17637,N_16308,N_16371);
and U17638 (N_17638,N_16601,N_16692);
nor U17639 (N_17639,N_16147,N_16457);
nor U17640 (N_17640,N_16269,N_16516);
nor U17641 (N_17641,N_16949,N_16692);
nand U17642 (N_17642,N_16794,N_16219);
nand U17643 (N_17643,N_16487,N_16592);
or U17644 (N_17644,N_16435,N_16857);
nor U17645 (N_17645,N_16878,N_16253);
nor U17646 (N_17646,N_16796,N_16050);
and U17647 (N_17647,N_16876,N_16619);
nor U17648 (N_17648,N_16298,N_16801);
xor U17649 (N_17649,N_16344,N_16953);
or U17650 (N_17650,N_16048,N_16600);
and U17651 (N_17651,N_16793,N_16638);
and U17652 (N_17652,N_16126,N_16063);
nand U17653 (N_17653,N_16822,N_16883);
xor U17654 (N_17654,N_16591,N_16719);
and U17655 (N_17655,N_16757,N_16548);
xor U17656 (N_17656,N_16077,N_16940);
and U17657 (N_17657,N_16286,N_16929);
xnor U17658 (N_17658,N_16349,N_16046);
or U17659 (N_17659,N_16339,N_16527);
and U17660 (N_17660,N_16873,N_16063);
nand U17661 (N_17661,N_16563,N_16633);
nand U17662 (N_17662,N_16621,N_16104);
and U17663 (N_17663,N_16747,N_16684);
nand U17664 (N_17664,N_16173,N_16998);
or U17665 (N_17665,N_16655,N_16807);
or U17666 (N_17666,N_16348,N_16688);
or U17667 (N_17667,N_16997,N_16901);
and U17668 (N_17668,N_16682,N_16661);
nor U17669 (N_17669,N_16335,N_16669);
nand U17670 (N_17670,N_16711,N_16761);
and U17671 (N_17671,N_16564,N_16324);
xor U17672 (N_17672,N_16622,N_16783);
nor U17673 (N_17673,N_16543,N_16067);
nor U17674 (N_17674,N_16979,N_16704);
nor U17675 (N_17675,N_16543,N_16544);
nand U17676 (N_17676,N_16892,N_16422);
xnor U17677 (N_17677,N_16003,N_16392);
or U17678 (N_17678,N_16087,N_16403);
and U17679 (N_17679,N_16598,N_16599);
or U17680 (N_17680,N_16880,N_16286);
xnor U17681 (N_17681,N_16636,N_16061);
xnor U17682 (N_17682,N_16253,N_16217);
xnor U17683 (N_17683,N_16099,N_16969);
nand U17684 (N_17684,N_16072,N_16748);
or U17685 (N_17685,N_16001,N_16774);
nand U17686 (N_17686,N_16302,N_16241);
nand U17687 (N_17687,N_16320,N_16581);
nand U17688 (N_17688,N_16864,N_16450);
nand U17689 (N_17689,N_16857,N_16996);
nor U17690 (N_17690,N_16694,N_16605);
nor U17691 (N_17691,N_16397,N_16313);
nor U17692 (N_17692,N_16417,N_16837);
and U17693 (N_17693,N_16518,N_16980);
nand U17694 (N_17694,N_16891,N_16321);
nand U17695 (N_17695,N_16383,N_16666);
nor U17696 (N_17696,N_16325,N_16874);
nor U17697 (N_17697,N_16450,N_16194);
nand U17698 (N_17698,N_16865,N_16149);
nand U17699 (N_17699,N_16082,N_16610);
nor U17700 (N_17700,N_16293,N_16811);
and U17701 (N_17701,N_16427,N_16511);
xor U17702 (N_17702,N_16071,N_16862);
nor U17703 (N_17703,N_16317,N_16616);
xnor U17704 (N_17704,N_16627,N_16762);
and U17705 (N_17705,N_16444,N_16118);
and U17706 (N_17706,N_16758,N_16151);
nor U17707 (N_17707,N_16337,N_16327);
or U17708 (N_17708,N_16716,N_16065);
nand U17709 (N_17709,N_16971,N_16505);
xor U17710 (N_17710,N_16347,N_16201);
nor U17711 (N_17711,N_16235,N_16558);
nand U17712 (N_17712,N_16070,N_16897);
nand U17713 (N_17713,N_16430,N_16138);
nor U17714 (N_17714,N_16935,N_16696);
and U17715 (N_17715,N_16660,N_16763);
nand U17716 (N_17716,N_16529,N_16303);
nand U17717 (N_17717,N_16101,N_16835);
xnor U17718 (N_17718,N_16246,N_16765);
or U17719 (N_17719,N_16320,N_16451);
nor U17720 (N_17720,N_16634,N_16112);
nand U17721 (N_17721,N_16413,N_16414);
nand U17722 (N_17722,N_16481,N_16619);
or U17723 (N_17723,N_16166,N_16872);
xor U17724 (N_17724,N_16479,N_16297);
and U17725 (N_17725,N_16697,N_16466);
nand U17726 (N_17726,N_16910,N_16471);
xor U17727 (N_17727,N_16785,N_16028);
nand U17728 (N_17728,N_16281,N_16622);
nand U17729 (N_17729,N_16289,N_16503);
or U17730 (N_17730,N_16110,N_16911);
nor U17731 (N_17731,N_16274,N_16003);
nor U17732 (N_17732,N_16613,N_16970);
nand U17733 (N_17733,N_16268,N_16632);
nor U17734 (N_17734,N_16789,N_16818);
xnor U17735 (N_17735,N_16877,N_16510);
and U17736 (N_17736,N_16274,N_16316);
and U17737 (N_17737,N_16086,N_16903);
xor U17738 (N_17738,N_16996,N_16387);
nor U17739 (N_17739,N_16509,N_16789);
or U17740 (N_17740,N_16503,N_16574);
and U17741 (N_17741,N_16276,N_16600);
and U17742 (N_17742,N_16777,N_16074);
nor U17743 (N_17743,N_16493,N_16085);
and U17744 (N_17744,N_16699,N_16087);
or U17745 (N_17745,N_16950,N_16900);
nand U17746 (N_17746,N_16179,N_16573);
and U17747 (N_17747,N_16808,N_16931);
nor U17748 (N_17748,N_16681,N_16979);
or U17749 (N_17749,N_16554,N_16589);
nand U17750 (N_17750,N_16016,N_16646);
nand U17751 (N_17751,N_16530,N_16975);
or U17752 (N_17752,N_16892,N_16741);
and U17753 (N_17753,N_16956,N_16857);
xnor U17754 (N_17754,N_16371,N_16827);
nand U17755 (N_17755,N_16344,N_16796);
and U17756 (N_17756,N_16480,N_16308);
nor U17757 (N_17757,N_16312,N_16420);
nor U17758 (N_17758,N_16214,N_16903);
and U17759 (N_17759,N_16495,N_16053);
nand U17760 (N_17760,N_16069,N_16791);
nand U17761 (N_17761,N_16007,N_16559);
or U17762 (N_17762,N_16621,N_16823);
nand U17763 (N_17763,N_16161,N_16177);
nand U17764 (N_17764,N_16303,N_16449);
or U17765 (N_17765,N_16317,N_16457);
nand U17766 (N_17766,N_16608,N_16740);
xnor U17767 (N_17767,N_16810,N_16297);
and U17768 (N_17768,N_16492,N_16518);
xor U17769 (N_17769,N_16558,N_16441);
and U17770 (N_17770,N_16562,N_16177);
and U17771 (N_17771,N_16826,N_16636);
nand U17772 (N_17772,N_16800,N_16550);
nand U17773 (N_17773,N_16152,N_16349);
and U17774 (N_17774,N_16342,N_16523);
and U17775 (N_17775,N_16528,N_16293);
and U17776 (N_17776,N_16163,N_16867);
xor U17777 (N_17777,N_16548,N_16715);
nor U17778 (N_17778,N_16248,N_16459);
nor U17779 (N_17779,N_16245,N_16102);
nand U17780 (N_17780,N_16991,N_16057);
xor U17781 (N_17781,N_16573,N_16102);
nand U17782 (N_17782,N_16064,N_16559);
nor U17783 (N_17783,N_16592,N_16660);
nand U17784 (N_17784,N_16241,N_16064);
or U17785 (N_17785,N_16137,N_16278);
or U17786 (N_17786,N_16231,N_16162);
nand U17787 (N_17787,N_16642,N_16959);
nor U17788 (N_17788,N_16454,N_16247);
nand U17789 (N_17789,N_16148,N_16114);
and U17790 (N_17790,N_16008,N_16694);
and U17791 (N_17791,N_16692,N_16290);
or U17792 (N_17792,N_16865,N_16376);
or U17793 (N_17793,N_16192,N_16627);
nand U17794 (N_17794,N_16016,N_16373);
xnor U17795 (N_17795,N_16497,N_16557);
or U17796 (N_17796,N_16361,N_16679);
or U17797 (N_17797,N_16199,N_16644);
nand U17798 (N_17798,N_16343,N_16069);
or U17799 (N_17799,N_16741,N_16838);
or U17800 (N_17800,N_16107,N_16002);
xor U17801 (N_17801,N_16813,N_16967);
nor U17802 (N_17802,N_16503,N_16087);
nor U17803 (N_17803,N_16990,N_16319);
and U17804 (N_17804,N_16836,N_16269);
xor U17805 (N_17805,N_16512,N_16129);
xor U17806 (N_17806,N_16579,N_16958);
nor U17807 (N_17807,N_16921,N_16588);
xnor U17808 (N_17808,N_16858,N_16452);
or U17809 (N_17809,N_16647,N_16374);
xnor U17810 (N_17810,N_16567,N_16363);
xnor U17811 (N_17811,N_16973,N_16062);
and U17812 (N_17812,N_16179,N_16394);
xor U17813 (N_17813,N_16581,N_16982);
or U17814 (N_17814,N_16509,N_16285);
nor U17815 (N_17815,N_16819,N_16451);
xor U17816 (N_17816,N_16912,N_16637);
or U17817 (N_17817,N_16799,N_16305);
or U17818 (N_17818,N_16735,N_16876);
or U17819 (N_17819,N_16596,N_16883);
and U17820 (N_17820,N_16161,N_16837);
nand U17821 (N_17821,N_16231,N_16007);
or U17822 (N_17822,N_16094,N_16967);
nand U17823 (N_17823,N_16804,N_16723);
nand U17824 (N_17824,N_16469,N_16898);
nand U17825 (N_17825,N_16814,N_16033);
xor U17826 (N_17826,N_16169,N_16096);
nor U17827 (N_17827,N_16767,N_16060);
nor U17828 (N_17828,N_16568,N_16460);
or U17829 (N_17829,N_16696,N_16720);
nor U17830 (N_17830,N_16544,N_16296);
and U17831 (N_17831,N_16901,N_16114);
or U17832 (N_17832,N_16036,N_16700);
or U17833 (N_17833,N_16538,N_16090);
or U17834 (N_17834,N_16931,N_16096);
nor U17835 (N_17835,N_16646,N_16840);
or U17836 (N_17836,N_16514,N_16156);
nor U17837 (N_17837,N_16667,N_16710);
nand U17838 (N_17838,N_16653,N_16051);
and U17839 (N_17839,N_16904,N_16650);
or U17840 (N_17840,N_16126,N_16560);
nor U17841 (N_17841,N_16602,N_16543);
xnor U17842 (N_17842,N_16168,N_16049);
and U17843 (N_17843,N_16401,N_16231);
xor U17844 (N_17844,N_16378,N_16572);
nor U17845 (N_17845,N_16492,N_16059);
or U17846 (N_17846,N_16455,N_16082);
or U17847 (N_17847,N_16777,N_16361);
and U17848 (N_17848,N_16818,N_16319);
and U17849 (N_17849,N_16738,N_16176);
nand U17850 (N_17850,N_16184,N_16993);
nand U17851 (N_17851,N_16148,N_16079);
and U17852 (N_17852,N_16314,N_16666);
or U17853 (N_17853,N_16972,N_16509);
and U17854 (N_17854,N_16430,N_16618);
or U17855 (N_17855,N_16645,N_16881);
or U17856 (N_17856,N_16053,N_16146);
nor U17857 (N_17857,N_16957,N_16277);
nor U17858 (N_17858,N_16556,N_16477);
and U17859 (N_17859,N_16490,N_16130);
xor U17860 (N_17860,N_16621,N_16774);
nor U17861 (N_17861,N_16449,N_16171);
nand U17862 (N_17862,N_16153,N_16067);
and U17863 (N_17863,N_16835,N_16980);
xor U17864 (N_17864,N_16204,N_16299);
xnor U17865 (N_17865,N_16337,N_16532);
or U17866 (N_17866,N_16783,N_16782);
nand U17867 (N_17867,N_16579,N_16311);
xnor U17868 (N_17868,N_16132,N_16628);
and U17869 (N_17869,N_16241,N_16106);
or U17870 (N_17870,N_16158,N_16240);
nand U17871 (N_17871,N_16612,N_16607);
xnor U17872 (N_17872,N_16225,N_16016);
or U17873 (N_17873,N_16689,N_16300);
nand U17874 (N_17874,N_16073,N_16230);
and U17875 (N_17875,N_16184,N_16851);
nand U17876 (N_17876,N_16887,N_16019);
and U17877 (N_17877,N_16144,N_16721);
or U17878 (N_17878,N_16601,N_16391);
xor U17879 (N_17879,N_16408,N_16123);
xnor U17880 (N_17880,N_16960,N_16524);
nand U17881 (N_17881,N_16746,N_16834);
nand U17882 (N_17882,N_16001,N_16478);
xnor U17883 (N_17883,N_16621,N_16493);
or U17884 (N_17884,N_16605,N_16317);
nor U17885 (N_17885,N_16784,N_16364);
nand U17886 (N_17886,N_16197,N_16771);
xor U17887 (N_17887,N_16911,N_16817);
xor U17888 (N_17888,N_16006,N_16956);
and U17889 (N_17889,N_16536,N_16534);
nand U17890 (N_17890,N_16961,N_16956);
nor U17891 (N_17891,N_16259,N_16315);
nor U17892 (N_17892,N_16752,N_16821);
or U17893 (N_17893,N_16022,N_16558);
nor U17894 (N_17894,N_16480,N_16321);
and U17895 (N_17895,N_16229,N_16626);
and U17896 (N_17896,N_16918,N_16842);
or U17897 (N_17897,N_16908,N_16563);
xor U17898 (N_17898,N_16319,N_16143);
or U17899 (N_17899,N_16870,N_16572);
or U17900 (N_17900,N_16209,N_16499);
xor U17901 (N_17901,N_16314,N_16882);
nor U17902 (N_17902,N_16217,N_16819);
nor U17903 (N_17903,N_16865,N_16715);
and U17904 (N_17904,N_16327,N_16184);
xnor U17905 (N_17905,N_16480,N_16818);
or U17906 (N_17906,N_16756,N_16725);
nand U17907 (N_17907,N_16609,N_16150);
nand U17908 (N_17908,N_16686,N_16680);
xnor U17909 (N_17909,N_16280,N_16656);
nor U17910 (N_17910,N_16787,N_16989);
nor U17911 (N_17911,N_16273,N_16502);
nor U17912 (N_17912,N_16852,N_16538);
or U17913 (N_17913,N_16285,N_16726);
and U17914 (N_17914,N_16546,N_16807);
nor U17915 (N_17915,N_16335,N_16274);
nand U17916 (N_17916,N_16747,N_16376);
or U17917 (N_17917,N_16189,N_16622);
nand U17918 (N_17918,N_16614,N_16682);
nand U17919 (N_17919,N_16884,N_16802);
and U17920 (N_17920,N_16094,N_16350);
nor U17921 (N_17921,N_16249,N_16445);
xnor U17922 (N_17922,N_16950,N_16220);
or U17923 (N_17923,N_16600,N_16738);
nand U17924 (N_17924,N_16853,N_16471);
nand U17925 (N_17925,N_16569,N_16140);
xor U17926 (N_17926,N_16274,N_16445);
or U17927 (N_17927,N_16636,N_16965);
nand U17928 (N_17928,N_16149,N_16049);
xor U17929 (N_17929,N_16679,N_16974);
and U17930 (N_17930,N_16989,N_16421);
xor U17931 (N_17931,N_16311,N_16969);
xor U17932 (N_17932,N_16292,N_16030);
nand U17933 (N_17933,N_16721,N_16292);
nor U17934 (N_17934,N_16710,N_16008);
nand U17935 (N_17935,N_16465,N_16943);
nand U17936 (N_17936,N_16569,N_16367);
or U17937 (N_17937,N_16361,N_16642);
nand U17938 (N_17938,N_16804,N_16595);
nand U17939 (N_17939,N_16161,N_16031);
or U17940 (N_17940,N_16589,N_16274);
and U17941 (N_17941,N_16822,N_16869);
and U17942 (N_17942,N_16745,N_16418);
and U17943 (N_17943,N_16265,N_16446);
nor U17944 (N_17944,N_16373,N_16669);
xnor U17945 (N_17945,N_16250,N_16204);
xor U17946 (N_17946,N_16847,N_16839);
xnor U17947 (N_17947,N_16117,N_16152);
and U17948 (N_17948,N_16757,N_16734);
or U17949 (N_17949,N_16679,N_16809);
and U17950 (N_17950,N_16273,N_16272);
or U17951 (N_17951,N_16240,N_16757);
and U17952 (N_17952,N_16062,N_16903);
and U17953 (N_17953,N_16291,N_16520);
nor U17954 (N_17954,N_16419,N_16321);
and U17955 (N_17955,N_16800,N_16330);
nor U17956 (N_17956,N_16223,N_16566);
or U17957 (N_17957,N_16340,N_16680);
and U17958 (N_17958,N_16982,N_16349);
and U17959 (N_17959,N_16756,N_16604);
xor U17960 (N_17960,N_16770,N_16301);
and U17961 (N_17961,N_16891,N_16767);
xnor U17962 (N_17962,N_16336,N_16213);
xor U17963 (N_17963,N_16264,N_16854);
and U17964 (N_17964,N_16170,N_16760);
or U17965 (N_17965,N_16448,N_16675);
and U17966 (N_17966,N_16500,N_16715);
nor U17967 (N_17967,N_16712,N_16297);
nand U17968 (N_17968,N_16345,N_16429);
nand U17969 (N_17969,N_16395,N_16711);
xnor U17970 (N_17970,N_16883,N_16832);
or U17971 (N_17971,N_16130,N_16748);
nand U17972 (N_17972,N_16669,N_16330);
nor U17973 (N_17973,N_16900,N_16051);
or U17974 (N_17974,N_16908,N_16157);
or U17975 (N_17975,N_16081,N_16581);
nor U17976 (N_17976,N_16844,N_16849);
and U17977 (N_17977,N_16982,N_16258);
or U17978 (N_17978,N_16361,N_16586);
nand U17979 (N_17979,N_16317,N_16887);
nand U17980 (N_17980,N_16148,N_16718);
nor U17981 (N_17981,N_16048,N_16420);
nand U17982 (N_17982,N_16691,N_16351);
or U17983 (N_17983,N_16035,N_16914);
xor U17984 (N_17984,N_16943,N_16965);
or U17985 (N_17985,N_16006,N_16913);
nor U17986 (N_17986,N_16998,N_16900);
nor U17987 (N_17987,N_16938,N_16914);
or U17988 (N_17988,N_16999,N_16584);
nand U17989 (N_17989,N_16346,N_16506);
and U17990 (N_17990,N_16312,N_16178);
xnor U17991 (N_17991,N_16237,N_16223);
nor U17992 (N_17992,N_16432,N_16181);
xnor U17993 (N_17993,N_16358,N_16673);
xor U17994 (N_17994,N_16733,N_16570);
and U17995 (N_17995,N_16311,N_16987);
and U17996 (N_17996,N_16809,N_16526);
and U17997 (N_17997,N_16336,N_16579);
or U17998 (N_17998,N_16036,N_16853);
xnor U17999 (N_17999,N_16387,N_16597);
xnor U18000 (N_18000,N_17823,N_17968);
xnor U18001 (N_18001,N_17461,N_17716);
nand U18002 (N_18002,N_17237,N_17809);
nand U18003 (N_18003,N_17316,N_17489);
nand U18004 (N_18004,N_17165,N_17057);
nand U18005 (N_18005,N_17937,N_17503);
and U18006 (N_18006,N_17186,N_17211);
nor U18007 (N_18007,N_17976,N_17181);
or U18008 (N_18008,N_17991,N_17178);
nor U18009 (N_18009,N_17870,N_17891);
or U18010 (N_18010,N_17625,N_17312);
or U18011 (N_18011,N_17642,N_17561);
and U18012 (N_18012,N_17566,N_17841);
nor U18013 (N_18013,N_17637,N_17347);
or U18014 (N_18014,N_17224,N_17899);
nand U18015 (N_18015,N_17966,N_17086);
or U18016 (N_18016,N_17518,N_17871);
nand U18017 (N_18017,N_17973,N_17172);
nor U18018 (N_18018,N_17390,N_17905);
nand U18019 (N_18019,N_17038,N_17348);
nor U18020 (N_18020,N_17046,N_17156);
xor U18021 (N_18021,N_17450,N_17840);
and U18022 (N_18022,N_17725,N_17915);
and U18023 (N_18023,N_17689,N_17932);
xor U18024 (N_18024,N_17494,N_17830);
xnor U18025 (N_18025,N_17460,N_17606);
nor U18026 (N_18026,N_17258,N_17677);
or U18027 (N_18027,N_17003,N_17170);
xor U18028 (N_18028,N_17943,N_17977);
nand U18029 (N_18029,N_17836,N_17043);
xor U18030 (N_18030,N_17410,N_17294);
nor U18031 (N_18031,N_17185,N_17713);
nor U18032 (N_18032,N_17240,N_17231);
or U18033 (N_18033,N_17730,N_17884);
xnor U18034 (N_18034,N_17926,N_17555);
nor U18035 (N_18035,N_17184,N_17238);
and U18036 (N_18036,N_17102,N_17493);
or U18037 (N_18037,N_17252,N_17183);
nand U18038 (N_18038,N_17748,N_17417);
nor U18039 (N_18039,N_17299,N_17131);
nor U18040 (N_18040,N_17007,N_17075);
nand U18041 (N_18041,N_17580,N_17717);
xnor U18042 (N_18042,N_17037,N_17249);
or U18043 (N_18043,N_17136,N_17314);
nand U18044 (N_18044,N_17261,N_17601);
xor U18045 (N_18045,N_17922,N_17216);
and U18046 (N_18046,N_17887,N_17711);
and U18047 (N_18047,N_17371,N_17705);
and U18048 (N_18048,N_17066,N_17189);
nand U18049 (N_18049,N_17874,N_17818);
nand U18050 (N_18050,N_17988,N_17635);
nor U18051 (N_18051,N_17069,N_17586);
or U18052 (N_18052,N_17218,N_17276);
nor U18053 (N_18053,N_17033,N_17708);
nand U18054 (N_18054,N_17633,N_17963);
or U18055 (N_18055,N_17659,N_17375);
or U18056 (N_18056,N_17828,N_17403);
or U18057 (N_18057,N_17488,N_17281);
or U18058 (N_18058,N_17023,N_17048);
or U18059 (N_18059,N_17678,N_17885);
nor U18060 (N_18060,N_17663,N_17860);
or U18061 (N_18061,N_17389,N_17453);
and U18062 (N_18062,N_17052,N_17643);
xor U18063 (N_18063,N_17919,N_17970);
and U18064 (N_18064,N_17990,N_17333);
and U18065 (N_18065,N_17498,N_17934);
xnor U18066 (N_18066,N_17569,N_17616);
nand U18067 (N_18067,N_17217,N_17116);
nor U18068 (N_18068,N_17173,N_17564);
and U18069 (N_18069,N_17533,N_17005);
xor U18070 (N_18070,N_17100,N_17902);
nand U18071 (N_18071,N_17826,N_17062);
xor U18072 (N_18072,N_17927,N_17463);
nand U18073 (N_18073,N_17691,N_17767);
and U18074 (N_18074,N_17055,N_17909);
nand U18075 (N_18075,N_17340,N_17827);
or U18076 (N_18076,N_17317,N_17119);
and U18077 (N_18077,N_17148,N_17464);
or U18078 (N_18078,N_17027,N_17204);
or U18079 (N_18079,N_17263,N_17321);
nor U18080 (N_18080,N_17452,N_17802);
xnor U18081 (N_18081,N_17568,N_17829);
or U18082 (N_18082,N_17532,N_17668);
nor U18083 (N_18083,N_17272,N_17866);
xnor U18084 (N_18084,N_17949,N_17089);
nor U18085 (N_18085,N_17168,N_17792);
and U18086 (N_18086,N_17824,N_17160);
or U18087 (N_18087,N_17124,N_17923);
nand U18088 (N_18088,N_17769,N_17481);
and U18089 (N_18089,N_17983,N_17203);
nor U18090 (N_18090,N_17018,N_17227);
xor U18091 (N_18091,N_17239,N_17087);
nand U18092 (N_18092,N_17683,N_17351);
nor U18093 (N_18093,N_17607,N_17125);
nand U18094 (N_18094,N_17992,N_17621);
and U18095 (N_18095,N_17719,N_17507);
nand U18096 (N_18096,N_17393,N_17432);
nand U18097 (N_18097,N_17641,N_17588);
or U18098 (N_18098,N_17422,N_17971);
xnor U18099 (N_18099,N_17442,N_17381);
or U18100 (N_18100,N_17549,N_17735);
and U18101 (N_18101,N_17614,N_17524);
or U18102 (N_18102,N_17650,N_17394);
and U18103 (N_18103,N_17952,N_17400);
and U18104 (N_18104,N_17478,N_17812);
nand U18105 (N_18105,N_17636,N_17806);
and U18106 (N_18106,N_17634,N_17781);
and U18107 (N_18107,N_17080,N_17419);
nand U18108 (N_18108,N_17358,N_17587);
nor U18109 (N_18109,N_17538,N_17001);
and U18110 (N_18110,N_17629,N_17120);
or U18111 (N_18111,N_17554,N_17720);
and U18112 (N_18112,N_17137,N_17512);
nand U18113 (N_18113,N_17330,N_17788);
nand U18114 (N_18114,N_17024,N_17177);
nand U18115 (N_18115,N_17014,N_17448);
xnor U18116 (N_18116,N_17301,N_17756);
nand U18117 (N_18117,N_17245,N_17997);
nand U18118 (N_18118,N_17029,N_17863);
or U18119 (N_18119,N_17598,N_17567);
xnor U18120 (N_18120,N_17685,N_17918);
nand U18121 (N_18121,N_17557,N_17082);
and U18122 (N_18122,N_17912,N_17869);
xnor U18123 (N_18123,N_17940,N_17302);
and U18124 (N_18124,N_17759,N_17962);
or U18125 (N_18125,N_17502,N_17645);
or U18126 (N_18126,N_17010,N_17560);
xnor U18127 (N_18127,N_17382,N_17819);
or U18128 (N_18128,N_17842,N_17545);
nor U18129 (N_18129,N_17061,N_17103);
nand U18130 (N_18130,N_17619,N_17797);
xor U18131 (N_18131,N_17671,N_17473);
xor U18132 (N_18132,N_17993,N_17429);
or U18133 (N_18133,N_17248,N_17449);
and U18134 (N_18134,N_17446,N_17979);
and U18135 (N_18135,N_17649,N_17615);
nor U18136 (N_18136,N_17487,N_17265);
or U18137 (N_18137,N_17126,N_17044);
nor U18138 (N_18138,N_17149,N_17803);
or U18139 (N_18139,N_17627,N_17256);
and U18140 (N_18140,N_17880,N_17304);
and U18141 (N_18141,N_17822,N_17071);
nor U18142 (N_18142,N_17040,N_17195);
nand U18143 (N_18143,N_17867,N_17171);
xor U18144 (N_18144,N_17692,N_17269);
nand U18145 (N_18145,N_17114,N_17270);
and U18146 (N_18146,N_17274,N_17243);
or U18147 (N_18147,N_17201,N_17345);
xor U18148 (N_18148,N_17110,N_17159);
nand U18149 (N_18149,N_17318,N_17698);
xor U18150 (N_18150,N_17710,N_17908);
nor U18151 (N_18151,N_17648,N_17697);
nand U18152 (N_18152,N_17212,N_17540);
xor U18153 (N_18153,N_17776,N_17876);
and U18154 (N_18154,N_17056,N_17839);
nor U18155 (N_18155,N_17613,N_17412);
and U18156 (N_18156,N_17742,N_17222);
or U18157 (N_18157,N_17608,N_17612);
or U18158 (N_18158,N_17680,N_17658);
or U18159 (N_18159,N_17205,N_17595);
and U18160 (N_18160,N_17127,N_17289);
xor U18161 (N_18161,N_17673,N_17196);
nor U18162 (N_18162,N_17435,N_17845);
xnor U18163 (N_18163,N_17959,N_17793);
and U18164 (N_18164,N_17101,N_17581);
nor U18165 (N_18165,N_17287,N_17356);
or U18166 (N_18166,N_17313,N_17399);
and U18167 (N_18167,N_17921,N_17631);
xnor U18168 (N_18168,N_17322,N_17327);
nand U18169 (N_18169,N_17931,N_17406);
nand U18170 (N_18170,N_17379,N_17132);
nand U18171 (N_18171,N_17129,N_17746);
xnor U18172 (N_18172,N_17097,N_17579);
and U18173 (N_18173,N_17938,N_17456);
or U18174 (N_18174,N_17107,N_17404);
nand U18175 (N_18175,N_17833,N_17883);
or U18176 (N_18176,N_17485,N_17143);
nand U18177 (N_18177,N_17197,N_17754);
or U18178 (N_18178,N_17780,N_17760);
nor U18179 (N_18179,N_17571,N_17652);
or U18180 (N_18180,N_17986,N_17431);
and U18181 (N_18181,N_17743,N_17537);
xnor U18182 (N_18182,N_17367,N_17349);
xnor U18183 (N_18183,N_17913,N_17041);
and U18184 (N_18184,N_17147,N_17141);
xor U18185 (N_18185,N_17319,N_17324);
nor U18186 (N_18186,N_17661,N_17961);
and U18187 (N_18187,N_17747,N_17416);
or U18188 (N_18188,N_17994,N_17657);
or U18189 (N_18189,N_17800,N_17213);
nor U18190 (N_18190,N_17734,N_17732);
or U18191 (N_18191,N_17368,N_17343);
and U18192 (N_18192,N_17392,N_17670);
nand U18193 (N_18193,N_17164,N_17896);
and U18194 (N_18194,N_17975,N_17706);
or U18195 (N_18195,N_17329,N_17738);
nand U18196 (N_18196,N_17674,N_17965);
xnor U18197 (N_18197,N_17191,N_17411);
nand U18198 (N_18198,N_17233,N_17690);
nand U18199 (N_18199,N_17548,N_17831);
xnor U18200 (N_18200,N_17401,N_17623);
nor U18201 (N_18201,N_17817,N_17074);
or U18202 (N_18202,N_17235,N_17246);
or U18203 (N_18203,N_17259,N_17445);
xnor U18204 (N_18204,N_17223,N_17072);
xor U18205 (N_18205,N_17112,N_17011);
and U18206 (N_18206,N_17843,N_17577);
or U18207 (N_18207,N_17664,N_17428);
or U18208 (N_18208,N_17958,N_17310);
nand U18209 (N_18209,N_17187,N_17199);
xnor U18210 (N_18210,N_17744,N_17553);
nor U18211 (N_18211,N_17280,N_17834);
nor U18212 (N_18212,N_17541,N_17064);
nor U18213 (N_18213,N_17700,N_17073);
or U18214 (N_18214,N_17391,N_17482);
nor U18215 (N_18215,N_17361,N_17928);
xor U18216 (N_18216,N_17336,N_17153);
or U18217 (N_18217,N_17506,N_17647);
and U18218 (N_18218,N_17207,N_17500);
nor U18219 (N_18219,N_17849,N_17225);
xnor U18220 (N_18220,N_17724,N_17609);
nand U18221 (N_18221,N_17508,N_17474);
nand U18222 (N_18222,N_17167,N_17210);
or U18223 (N_18223,N_17363,N_17941);
nor U18224 (N_18224,N_17437,N_17106);
nor U18225 (N_18225,N_17063,N_17017);
xor U18226 (N_18226,N_17855,N_17282);
nand U18227 (N_18227,N_17531,N_17556);
and U18228 (N_18228,N_17241,N_17140);
nor U18229 (N_18229,N_17472,N_17413);
or U18230 (N_18230,N_17777,N_17542);
nand U18231 (N_18231,N_17479,N_17944);
and U18232 (N_18232,N_17888,N_17602);
and U18233 (N_18233,N_17694,N_17946);
and U18234 (N_18234,N_17315,N_17194);
or U18235 (N_18235,N_17130,N_17501);
and U18236 (N_18236,N_17740,N_17284);
nand U18237 (N_18237,N_17254,N_17513);
and U18238 (N_18238,N_17380,N_17768);
xnor U18239 (N_18239,N_17704,N_17088);
and U18240 (N_18240,N_17104,N_17320);
and U18241 (N_18241,N_17878,N_17520);
nor U18242 (N_18242,N_17296,N_17599);
and U18243 (N_18243,N_17872,N_17665);
xor U18244 (N_18244,N_17045,N_17339);
or U18245 (N_18245,N_17789,N_17752);
nor U18246 (N_18246,N_17105,N_17260);
xor U18247 (N_18247,N_17257,N_17632);
nor U18248 (N_18248,N_17757,N_17536);
nand U18249 (N_18249,N_17681,N_17408);
xnor U18250 (N_18250,N_17832,N_17230);
or U18251 (N_18251,N_17675,N_17605);
nand U18252 (N_18252,N_17696,N_17440);
or U18253 (N_18253,N_17454,N_17215);
xor U18254 (N_18254,N_17590,N_17365);
xnor U18255 (N_18255,N_17525,N_17359);
xnor U18256 (N_18256,N_17558,N_17801);
nand U18257 (N_18257,N_17521,N_17811);
xor U18258 (N_18258,N_17861,N_17355);
or U18259 (N_18259,N_17850,N_17383);
nor U18260 (N_18260,N_17981,N_17157);
nor U18261 (N_18261,N_17423,N_17559);
or U18262 (N_18262,N_17251,N_17267);
and U18263 (N_18263,N_17626,N_17911);
nand U18264 (N_18264,N_17491,N_17220);
and U18265 (N_18265,N_17059,N_17714);
nand U18266 (N_18266,N_17152,N_17236);
nor U18267 (N_18267,N_17639,N_17377);
nand U18268 (N_18268,N_17158,N_17582);
or U18269 (N_18269,N_17480,N_17402);
nand U18270 (N_18270,N_17695,N_17835);
xor U18271 (N_18271,N_17407,N_17718);
nor U18272 (N_18272,N_17139,N_17022);
xor U18273 (N_18273,N_17535,N_17750);
nand U18274 (N_18274,N_17925,N_17775);
xor U18275 (N_18275,N_17755,N_17522);
or U18276 (N_18276,N_17890,N_17622);
nand U18277 (N_18277,N_17729,N_17113);
or U18278 (N_18278,N_17051,N_17892);
nor U18279 (N_18279,N_17050,N_17385);
and U18280 (N_18280,N_17644,N_17462);
xnor U18281 (N_18281,N_17731,N_17285);
and U18282 (N_18282,N_17162,N_17346);
or U18283 (N_18283,N_17728,N_17798);
or U18284 (N_18284,N_17807,N_17444);
and U18285 (N_18285,N_17618,N_17960);
nand U18286 (N_18286,N_17563,N_17693);
nor U18287 (N_18287,N_17956,N_17920);
nor U18288 (N_18288,N_17095,N_17786);
and U18289 (N_18289,N_17858,N_17936);
xor U18290 (N_18290,N_17420,N_17384);
xnor U18291 (N_18291,N_17455,N_17278);
or U18292 (N_18292,N_17596,N_17805);
nor U18293 (N_18293,N_17364,N_17264);
nor U18294 (N_18294,N_17808,N_17109);
and U18295 (N_18295,N_17682,N_17015);
nand U18296 (N_18296,N_17068,N_17311);
nor U18297 (N_18297,N_17935,N_17862);
or U18298 (N_18298,N_17585,N_17369);
and U18299 (N_18299,N_17424,N_17877);
and U18300 (N_18300,N_17477,N_17985);
xnor U18301 (N_18301,N_17758,N_17221);
and U18302 (N_18302,N_17604,N_17060);
or U18303 (N_18303,N_17886,N_17984);
nor U18304 (N_18304,N_17374,N_17111);
nor U18305 (N_18305,N_17950,N_17528);
nand U18306 (N_18306,N_17298,N_17398);
and U18307 (N_18307,N_17900,N_17666);
or U18308 (N_18308,N_17854,N_17293);
or U18309 (N_18309,N_17772,N_17443);
nor U18310 (N_18310,N_17337,N_17360);
nand U18311 (N_18311,N_17593,N_17133);
nand U18312 (N_18312,N_17155,N_17957);
or U18313 (N_18313,N_17209,N_17509);
nor U18314 (N_18314,N_17323,N_17332);
xnor U18315 (N_18315,N_17924,N_17362);
and U18316 (N_18316,N_17433,N_17552);
nand U18317 (N_18317,N_17378,N_17796);
or U18318 (N_18318,N_17669,N_17305);
nor U18319 (N_18319,N_17514,N_17425);
and U18320 (N_18320,N_17467,N_17096);
or U18321 (N_18321,N_17954,N_17034);
or U18322 (N_18322,N_17543,N_17974);
nor U18323 (N_18323,N_17309,N_17002);
nand U18324 (N_18324,N_17978,N_17042);
and U18325 (N_18325,N_17882,N_17953);
xor U18326 (N_18326,N_17815,N_17851);
and U18327 (N_18327,N_17418,N_17415);
xor U18328 (N_18328,N_17942,N_17373);
and U18329 (N_18329,N_17277,N_17099);
or U18330 (N_18330,N_17009,N_17466);
xor U18331 (N_18331,N_17897,N_17290);
or U18332 (N_18332,N_17844,N_17722);
xnor U18333 (N_18333,N_17036,N_17868);
nand U18334 (N_18334,N_17021,N_17334);
nand U18335 (N_18335,N_17510,N_17013);
or U18336 (N_18336,N_17094,N_17570);
nand U18337 (N_18337,N_17436,N_17996);
xnor U18338 (N_18338,N_17138,N_17771);
nor U18339 (N_18339,N_17092,N_17782);
and U18340 (N_18340,N_17065,N_17930);
xor U18341 (N_18341,N_17656,N_17778);
xor U18342 (N_18342,N_17202,N_17039);
xnor U18343 (N_18343,N_17686,N_17576);
xor U18344 (N_18344,N_17047,N_17268);
or U18345 (N_18345,N_17787,N_17497);
xor U18346 (N_18346,N_17654,N_17901);
xnor U18347 (N_18347,N_17012,N_17597);
xnor U18348 (N_18348,N_17486,N_17795);
and U18349 (N_18349,N_17190,N_17286);
nand U18350 (N_18350,N_17594,N_17770);
and U18351 (N_18351,N_17244,N_17085);
xnor U18352 (N_18352,N_17611,N_17784);
nand U18353 (N_18353,N_17762,N_17894);
nand U18354 (N_18354,N_17354,N_17799);
and U18355 (N_18355,N_17853,N_17054);
or U18356 (N_18356,N_17529,N_17283);
nor U18357 (N_18357,N_17458,N_17741);
or U18358 (N_18358,N_17967,N_17300);
or U18359 (N_18359,N_17484,N_17505);
xnor U18360 (N_18360,N_17646,N_17526);
xnor U18361 (N_18361,N_17247,N_17574);
xor U18362 (N_18362,N_17306,N_17206);
nor U18363 (N_18363,N_17721,N_17006);
nor U18364 (N_18364,N_17253,N_17135);
nor U18365 (N_18365,N_17873,N_17297);
or U18366 (N_18366,N_17504,N_17083);
nor U18367 (N_18367,N_17516,N_17551);
or U18368 (N_18368,N_17688,N_17342);
or U18369 (N_18369,N_17192,N_17219);
xor U18370 (N_18370,N_17409,N_17749);
xor U18371 (N_18371,N_17821,N_17288);
and U18372 (N_18372,N_17499,N_17341);
xor U18373 (N_18373,N_17307,N_17651);
nor U18374 (N_18374,N_17955,N_17414);
nor U18375 (N_18375,N_17447,N_17232);
nor U18376 (N_18376,N_17779,N_17350);
or U18377 (N_18377,N_17032,N_17995);
and U18378 (N_18378,N_17530,N_17591);
nor U18379 (N_18379,N_17396,N_17783);
xnor U18380 (N_18380,N_17547,N_17765);
nand U18381 (N_18381,N_17465,N_17081);
nor U18382 (N_18382,N_17434,N_17707);
nand U18383 (N_18383,N_17662,N_17947);
and U18384 (N_18384,N_17791,N_17366);
or U18385 (N_18385,N_17469,N_17929);
xor U18386 (N_18386,N_17904,N_17712);
nor U18387 (N_18387,N_17773,N_17076);
nor U18388 (N_18388,N_17889,N_17910);
and U18389 (N_18389,N_17266,N_17079);
or U18390 (N_18390,N_17134,N_17008);
nor U18391 (N_18391,N_17838,N_17736);
and U18392 (N_18392,N_17331,N_17335);
xor U18393 (N_18393,N_17945,N_17070);
or U18394 (N_18394,N_17603,N_17667);
nand U18395 (N_18395,N_17200,N_17214);
nand U18396 (N_18396,N_17151,N_17439);
nor U18397 (N_18397,N_17163,N_17751);
or U18398 (N_18398,N_17739,N_17262);
or U18399 (N_18399,N_17723,N_17875);
xor U18400 (N_18400,N_17180,N_17895);
nand U18401 (N_18401,N_17078,N_17794);
nor U18402 (N_18402,N_17699,N_17182);
xnor U18403 (N_18403,N_17573,N_17430);
nor U18404 (N_18404,N_17982,N_17630);
nand U18405 (N_18405,N_17701,N_17676);
nand U18406 (N_18406,N_17421,N_17397);
nand U18407 (N_18407,N_17279,N_17546);
xor U18408 (N_18408,N_17933,N_17145);
nor U18409 (N_18409,N_17980,N_17019);
nor U18410 (N_18410,N_17804,N_17492);
or U18411 (N_18411,N_17969,N_17948);
nor U18412 (N_18412,N_17709,N_17405);
nand U18413 (N_18413,N_17534,N_17426);
xor U18414 (N_18414,N_17763,N_17058);
nand U18415 (N_18415,N_17790,N_17441);
and U18416 (N_18416,N_17077,N_17271);
nand U18417 (N_18417,N_17726,N_17624);
and U18418 (N_18418,N_17584,N_17169);
or U18419 (N_18419,N_17628,N_17848);
nand U18420 (N_18420,N_17575,N_17098);
or U18421 (N_18421,N_17091,N_17273);
nand U18422 (N_18422,N_17338,N_17856);
nor U18423 (N_18423,N_17093,N_17496);
nor U18424 (N_18424,N_17292,N_17242);
nor U18425 (N_18425,N_17898,N_17523);
nor U18426 (N_18426,N_17617,N_17030);
nand U18427 (N_18427,N_17176,N_17049);
nor U18428 (N_18428,N_17357,N_17761);
xor U18429 (N_18429,N_17174,N_17972);
or U18430 (N_18430,N_17108,N_17459);
nor U18431 (N_18431,N_17490,N_17325);
nor U18432 (N_18432,N_17703,N_17386);
and U18433 (N_18433,N_17814,N_17353);
and U18434 (N_18434,N_17939,N_17562);
nor U18435 (N_18435,N_17118,N_17825);
or U18436 (N_18436,N_17879,N_17179);
and U18437 (N_18437,N_17951,N_17228);
and U18438 (N_18438,N_17672,N_17640);
and U18439 (N_18439,N_17745,N_17687);
or U18440 (N_18440,N_17090,N_17067);
nand U18441 (N_18441,N_17715,N_17328);
xnor U18442 (N_18442,N_17035,N_17291);
nand U18443 (N_18443,N_17737,N_17837);
or U18444 (N_18444,N_17893,N_17539);
nor U18445 (N_18445,N_17438,N_17679);
xnor U18446 (N_18446,N_17193,N_17517);
xnor U18447 (N_18447,N_17495,N_17122);
nand U18448 (N_18448,N_17903,N_17115);
and U18449 (N_18449,N_17702,N_17150);
nor U18450 (N_18450,N_17527,N_17142);
xor U18451 (N_18451,N_17865,N_17660);
or U18452 (N_18452,N_17727,N_17733);
xor U18453 (N_18453,N_17198,N_17376);
nor U18454 (N_18454,N_17229,N_17188);
xor U18455 (N_18455,N_17226,N_17515);
and U18456 (N_18456,N_17810,N_17764);
nor U18457 (N_18457,N_17550,N_17161);
nor U18458 (N_18458,N_17208,N_17998);
nor U18459 (N_18459,N_17476,N_17544);
nand U18460 (N_18460,N_17020,N_17820);
and U18461 (N_18461,N_17914,N_17511);
and U18462 (N_18462,N_17917,N_17031);
xnor U18463 (N_18463,N_17427,N_17128);
nand U18464 (N_18464,N_17250,N_17370);
nor U18465 (N_18465,N_17589,N_17004);
or U18466 (N_18466,N_17846,N_17000);
xor U18467 (N_18467,N_17620,N_17610);
xnor U18468 (N_18468,N_17016,N_17987);
xor U18469 (N_18469,N_17565,N_17144);
nand U18470 (N_18470,N_17907,N_17388);
nor U18471 (N_18471,N_17470,N_17028);
or U18472 (N_18472,N_17451,N_17352);
nand U18473 (N_18473,N_17852,N_17774);
and U18474 (N_18474,N_17653,N_17753);
and U18475 (N_18475,N_17483,N_17857);
nand U18476 (N_18476,N_17964,N_17084);
nor U18477 (N_18477,N_17457,N_17053);
or U18478 (N_18478,N_17766,N_17117);
or U18479 (N_18479,N_17154,N_17475);
or U18480 (N_18480,N_17468,N_17906);
nand U18481 (N_18481,N_17881,N_17308);
and U18482 (N_18482,N_17638,N_17859);
xnor U18483 (N_18483,N_17592,N_17684);
or U18484 (N_18484,N_17326,N_17303);
and U18485 (N_18485,N_17600,N_17372);
nand U18486 (N_18486,N_17123,N_17025);
xor U18487 (N_18487,N_17816,N_17785);
xnor U18488 (N_18488,N_17175,N_17999);
nor U18489 (N_18489,N_17864,N_17655);
nor U18490 (N_18490,N_17519,N_17578);
nor U18491 (N_18491,N_17387,N_17344);
xnor U18492 (N_18492,N_17847,N_17813);
nor U18493 (N_18493,N_17295,N_17026);
xor U18494 (N_18494,N_17121,N_17234);
xor U18495 (N_18495,N_17583,N_17395);
or U18496 (N_18496,N_17275,N_17146);
xor U18497 (N_18497,N_17471,N_17166);
and U18498 (N_18498,N_17989,N_17255);
nand U18499 (N_18499,N_17916,N_17572);
xor U18500 (N_18500,N_17976,N_17074);
or U18501 (N_18501,N_17270,N_17364);
xor U18502 (N_18502,N_17888,N_17636);
nand U18503 (N_18503,N_17038,N_17362);
xor U18504 (N_18504,N_17938,N_17540);
or U18505 (N_18505,N_17349,N_17477);
or U18506 (N_18506,N_17487,N_17474);
nor U18507 (N_18507,N_17021,N_17856);
nor U18508 (N_18508,N_17759,N_17076);
or U18509 (N_18509,N_17600,N_17654);
nand U18510 (N_18510,N_17919,N_17046);
xor U18511 (N_18511,N_17254,N_17520);
nor U18512 (N_18512,N_17720,N_17853);
xor U18513 (N_18513,N_17153,N_17960);
nand U18514 (N_18514,N_17465,N_17615);
xnor U18515 (N_18515,N_17423,N_17979);
xor U18516 (N_18516,N_17620,N_17405);
and U18517 (N_18517,N_17223,N_17263);
nor U18518 (N_18518,N_17877,N_17879);
or U18519 (N_18519,N_17069,N_17690);
nor U18520 (N_18520,N_17275,N_17642);
nor U18521 (N_18521,N_17915,N_17018);
and U18522 (N_18522,N_17737,N_17946);
nor U18523 (N_18523,N_17826,N_17185);
nand U18524 (N_18524,N_17127,N_17416);
nor U18525 (N_18525,N_17087,N_17921);
or U18526 (N_18526,N_17296,N_17241);
xnor U18527 (N_18527,N_17078,N_17733);
or U18528 (N_18528,N_17388,N_17579);
nand U18529 (N_18529,N_17531,N_17104);
and U18530 (N_18530,N_17834,N_17970);
and U18531 (N_18531,N_17942,N_17559);
and U18532 (N_18532,N_17499,N_17975);
xor U18533 (N_18533,N_17620,N_17591);
nor U18534 (N_18534,N_17373,N_17327);
or U18535 (N_18535,N_17084,N_17126);
or U18536 (N_18536,N_17985,N_17618);
xnor U18537 (N_18537,N_17876,N_17358);
nor U18538 (N_18538,N_17351,N_17420);
and U18539 (N_18539,N_17659,N_17255);
nand U18540 (N_18540,N_17327,N_17467);
nand U18541 (N_18541,N_17788,N_17755);
or U18542 (N_18542,N_17819,N_17471);
xnor U18543 (N_18543,N_17635,N_17719);
and U18544 (N_18544,N_17764,N_17860);
and U18545 (N_18545,N_17812,N_17251);
xnor U18546 (N_18546,N_17946,N_17132);
and U18547 (N_18547,N_17647,N_17975);
xnor U18548 (N_18548,N_17851,N_17036);
nor U18549 (N_18549,N_17869,N_17249);
xnor U18550 (N_18550,N_17316,N_17184);
nand U18551 (N_18551,N_17078,N_17854);
nor U18552 (N_18552,N_17222,N_17447);
or U18553 (N_18553,N_17199,N_17378);
and U18554 (N_18554,N_17704,N_17751);
nor U18555 (N_18555,N_17133,N_17802);
nor U18556 (N_18556,N_17181,N_17598);
xnor U18557 (N_18557,N_17412,N_17745);
and U18558 (N_18558,N_17099,N_17526);
nor U18559 (N_18559,N_17085,N_17200);
nand U18560 (N_18560,N_17686,N_17043);
xnor U18561 (N_18561,N_17007,N_17412);
nand U18562 (N_18562,N_17174,N_17670);
nor U18563 (N_18563,N_17406,N_17758);
and U18564 (N_18564,N_17059,N_17194);
nor U18565 (N_18565,N_17660,N_17186);
and U18566 (N_18566,N_17328,N_17135);
nand U18567 (N_18567,N_17409,N_17362);
nor U18568 (N_18568,N_17277,N_17169);
or U18569 (N_18569,N_17088,N_17925);
nand U18570 (N_18570,N_17257,N_17701);
or U18571 (N_18571,N_17815,N_17358);
or U18572 (N_18572,N_17110,N_17249);
xnor U18573 (N_18573,N_17893,N_17098);
nor U18574 (N_18574,N_17059,N_17765);
and U18575 (N_18575,N_17763,N_17214);
and U18576 (N_18576,N_17818,N_17348);
xor U18577 (N_18577,N_17153,N_17990);
and U18578 (N_18578,N_17795,N_17752);
or U18579 (N_18579,N_17549,N_17346);
or U18580 (N_18580,N_17136,N_17128);
nand U18581 (N_18581,N_17961,N_17072);
nor U18582 (N_18582,N_17814,N_17726);
or U18583 (N_18583,N_17451,N_17933);
xnor U18584 (N_18584,N_17271,N_17736);
or U18585 (N_18585,N_17120,N_17310);
nor U18586 (N_18586,N_17653,N_17013);
or U18587 (N_18587,N_17964,N_17998);
xor U18588 (N_18588,N_17690,N_17266);
and U18589 (N_18589,N_17894,N_17546);
xor U18590 (N_18590,N_17972,N_17838);
nor U18591 (N_18591,N_17967,N_17671);
and U18592 (N_18592,N_17235,N_17170);
nor U18593 (N_18593,N_17052,N_17196);
xnor U18594 (N_18594,N_17733,N_17488);
and U18595 (N_18595,N_17404,N_17679);
nand U18596 (N_18596,N_17979,N_17477);
or U18597 (N_18597,N_17086,N_17928);
or U18598 (N_18598,N_17337,N_17080);
or U18599 (N_18599,N_17412,N_17602);
xor U18600 (N_18600,N_17609,N_17150);
and U18601 (N_18601,N_17328,N_17443);
nand U18602 (N_18602,N_17094,N_17548);
xor U18603 (N_18603,N_17708,N_17645);
and U18604 (N_18604,N_17835,N_17530);
or U18605 (N_18605,N_17798,N_17608);
nand U18606 (N_18606,N_17017,N_17941);
or U18607 (N_18607,N_17570,N_17543);
or U18608 (N_18608,N_17149,N_17877);
and U18609 (N_18609,N_17177,N_17402);
nand U18610 (N_18610,N_17812,N_17656);
nand U18611 (N_18611,N_17273,N_17775);
xnor U18612 (N_18612,N_17874,N_17660);
xnor U18613 (N_18613,N_17501,N_17079);
or U18614 (N_18614,N_17362,N_17594);
or U18615 (N_18615,N_17418,N_17276);
xor U18616 (N_18616,N_17815,N_17512);
nor U18617 (N_18617,N_17059,N_17907);
nand U18618 (N_18618,N_17991,N_17217);
nand U18619 (N_18619,N_17700,N_17094);
or U18620 (N_18620,N_17564,N_17679);
nand U18621 (N_18621,N_17460,N_17778);
xor U18622 (N_18622,N_17367,N_17689);
or U18623 (N_18623,N_17100,N_17519);
nor U18624 (N_18624,N_17862,N_17008);
or U18625 (N_18625,N_17758,N_17555);
or U18626 (N_18626,N_17307,N_17644);
xor U18627 (N_18627,N_17664,N_17854);
or U18628 (N_18628,N_17278,N_17430);
nand U18629 (N_18629,N_17094,N_17044);
nor U18630 (N_18630,N_17578,N_17870);
or U18631 (N_18631,N_17381,N_17913);
xor U18632 (N_18632,N_17368,N_17701);
nor U18633 (N_18633,N_17062,N_17225);
and U18634 (N_18634,N_17775,N_17983);
and U18635 (N_18635,N_17772,N_17816);
or U18636 (N_18636,N_17882,N_17702);
and U18637 (N_18637,N_17519,N_17703);
and U18638 (N_18638,N_17499,N_17072);
xnor U18639 (N_18639,N_17814,N_17937);
and U18640 (N_18640,N_17504,N_17896);
nor U18641 (N_18641,N_17182,N_17619);
xor U18642 (N_18642,N_17565,N_17990);
or U18643 (N_18643,N_17042,N_17470);
nor U18644 (N_18644,N_17177,N_17140);
xnor U18645 (N_18645,N_17588,N_17201);
xor U18646 (N_18646,N_17130,N_17866);
nor U18647 (N_18647,N_17362,N_17340);
or U18648 (N_18648,N_17058,N_17021);
nand U18649 (N_18649,N_17702,N_17799);
nand U18650 (N_18650,N_17155,N_17597);
xnor U18651 (N_18651,N_17066,N_17726);
nand U18652 (N_18652,N_17725,N_17044);
nor U18653 (N_18653,N_17824,N_17419);
nand U18654 (N_18654,N_17137,N_17503);
and U18655 (N_18655,N_17467,N_17606);
and U18656 (N_18656,N_17440,N_17372);
nor U18657 (N_18657,N_17612,N_17662);
and U18658 (N_18658,N_17594,N_17885);
xor U18659 (N_18659,N_17471,N_17583);
xor U18660 (N_18660,N_17743,N_17857);
and U18661 (N_18661,N_17476,N_17087);
nand U18662 (N_18662,N_17047,N_17063);
nand U18663 (N_18663,N_17832,N_17034);
and U18664 (N_18664,N_17068,N_17981);
nor U18665 (N_18665,N_17895,N_17534);
nand U18666 (N_18666,N_17762,N_17876);
nor U18667 (N_18667,N_17223,N_17271);
and U18668 (N_18668,N_17539,N_17371);
and U18669 (N_18669,N_17689,N_17701);
nand U18670 (N_18670,N_17689,N_17497);
xnor U18671 (N_18671,N_17276,N_17387);
nor U18672 (N_18672,N_17418,N_17177);
xor U18673 (N_18673,N_17821,N_17408);
nor U18674 (N_18674,N_17731,N_17893);
xnor U18675 (N_18675,N_17290,N_17039);
nor U18676 (N_18676,N_17496,N_17027);
xor U18677 (N_18677,N_17854,N_17780);
and U18678 (N_18678,N_17365,N_17631);
nand U18679 (N_18679,N_17992,N_17494);
nor U18680 (N_18680,N_17691,N_17746);
nand U18681 (N_18681,N_17733,N_17359);
xnor U18682 (N_18682,N_17695,N_17999);
and U18683 (N_18683,N_17446,N_17525);
or U18684 (N_18684,N_17185,N_17712);
and U18685 (N_18685,N_17078,N_17309);
and U18686 (N_18686,N_17063,N_17761);
and U18687 (N_18687,N_17574,N_17799);
or U18688 (N_18688,N_17892,N_17552);
xnor U18689 (N_18689,N_17239,N_17244);
nand U18690 (N_18690,N_17837,N_17444);
or U18691 (N_18691,N_17301,N_17967);
nor U18692 (N_18692,N_17804,N_17773);
nand U18693 (N_18693,N_17629,N_17710);
nand U18694 (N_18694,N_17360,N_17434);
nand U18695 (N_18695,N_17698,N_17539);
or U18696 (N_18696,N_17273,N_17200);
nor U18697 (N_18697,N_17801,N_17320);
nor U18698 (N_18698,N_17389,N_17154);
or U18699 (N_18699,N_17883,N_17672);
nand U18700 (N_18700,N_17738,N_17281);
or U18701 (N_18701,N_17719,N_17877);
or U18702 (N_18702,N_17216,N_17444);
nor U18703 (N_18703,N_17155,N_17534);
nor U18704 (N_18704,N_17257,N_17995);
or U18705 (N_18705,N_17034,N_17429);
and U18706 (N_18706,N_17585,N_17200);
nor U18707 (N_18707,N_17609,N_17715);
nor U18708 (N_18708,N_17964,N_17187);
nand U18709 (N_18709,N_17666,N_17302);
nand U18710 (N_18710,N_17106,N_17884);
nor U18711 (N_18711,N_17764,N_17026);
nand U18712 (N_18712,N_17682,N_17592);
nor U18713 (N_18713,N_17895,N_17317);
xnor U18714 (N_18714,N_17397,N_17861);
and U18715 (N_18715,N_17549,N_17370);
or U18716 (N_18716,N_17198,N_17139);
nor U18717 (N_18717,N_17069,N_17152);
and U18718 (N_18718,N_17690,N_17763);
and U18719 (N_18719,N_17829,N_17919);
or U18720 (N_18720,N_17173,N_17114);
nor U18721 (N_18721,N_17534,N_17783);
xor U18722 (N_18722,N_17537,N_17949);
xnor U18723 (N_18723,N_17856,N_17900);
xor U18724 (N_18724,N_17564,N_17983);
and U18725 (N_18725,N_17995,N_17114);
or U18726 (N_18726,N_17856,N_17808);
or U18727 (N_18727,N_17600,N_17085);
nand U18728 (N_18728,N_17568,N_17165);
nand U18729 (N_18729,N_17998,N_17121);
nand U18730 (N_18730,N_17501,N_17443);
xor U18731 (N_18731,N_17854,N_17338);
nor U18732 (N_18732,N_17482,N_17689);
nand U18733 (N_18733,N_17805,N_17007);
or U18734 (N_18734,N_17577,N_17124);
nor U18735 (N_18735,N_17995,N_17878);
or U18736 (N_18736,N_17937,N_17695);
and U18737 (N_18737,N_17468,N_17993);
xor U18738 (N_18738,N_17795,N_17822);
or U18739 (N_18739,N_17156,N_17960);
xnor U18740 (N_18740,N_17484,N_17906);
and U18741 (N_18741,N_17334,N_17187);
or U18742 (N_18742,N_17133,N_17869);
or U18743 (N_18743,N_17161,N_17230);
xnor U18744 (N_18744,N_17177,N_17030);
or U18745 (N_18745,N_17377,N_17175);
nand U18746 (N_18746,N_17382,N_17843);
nor U18747 (N_18747,N_17973,N_17951);
and U18748 (N_18748,N_17334,N_17893);
and U18749 (N_18749,N_17093,N_17030);
nor U18750 (N_18750,N_17336,N_17878);
and U18751 (N_18751,N_17440,N_17042);
or U18752 (N_18752,N_17692,N_17956);
or U18753 (N_18753,N_17665,N_17979);
nand U18754 (N_18754,N_17399,N_17920);
xor U18755 (N_18755,N_17214,N_17562);
xor U18756 (N_18756,N_17197,N_17196);
nand U18757 (N_18757,N_17746,N_17895);
or U18758 (N_18758,N_17246,N_17040);
or U18759 (N_18759,N_17369,N_17055);
or U18760 (N_18760,N_17836,N_17266);
or U18761 (N_18761,N_17420,N_17482);
or U18762 (N_18762,N_17533,N_17194);
and U18763 (N_18763,N_17799,N_17601);
nor U18764 (N_18764,N_17211,N_17774);
xor U18765 (N_18765,N_17570,N_17506);
nor U18766 (N_18766,N_17175,N_17621);
xnor U18767 (N_18767,N_17837,N_17592);
and U18768 (N_18768,N_17239,N_17219);
or U18769 (N_18769,N_17979,N_17679);
or U18770 (N_18770,N_17569,N_17754);
xnor U18771 (N_18771,N_17359,N_17207);
and U18772 (N_18772,N_17868,N_17576);
nor U18773 (N_18773,N_17402,N_17183);
nand U18774 (N_18774,N_17238,N_17021);
xnor U18775 (N_18775,N_17920,N_17454);
xnor U18776 (N_18776,N_17578,N_17791);
and U18777 (N_18777,N_17500,N_17351);
nor U18778 (N_18778,N_17243,N_17381);
nor U18779 (N_18779,N_17439,N_17017);
xor U18780 (N_18780,N_17223,N_17040);
xnor U18781 (N_18781,N_17187,N_17457);
or U18782 (N_18782,N_17207,N_17625);
and U18783 (N_18783,N_17415,N_17524);
nor U18784 (N_18784,N_17706,N_17946);
or U18785 (N_18785,N_17171,N_17378);
nor U18786 (N_18786,N_17498,N_17344);
and U18787 (N_18787,N_17242,N_17146);
and U18788 (N_18788,N_17171,N_17410);
nand U18789 (N_18789,N_17891,N_17123);
and U18790 (N_18790,N_17897,N_17690);
or U18791 (N_18791,N_17022,N_17281);
and U18792 (N_18792,N_17918,N_17246);
and U18793 (N_18793,N_17173,N_17775);
or U18794 (N_18794,N_17954,N_17285);
xnor U18795 (N_18795,N_17507,N_17251);
nand U18796 (N_18796,N_17222,N_17982);
and U18797 (N_18797,N_17029,N_17284);
and U18798 (N_18798,N_17396,N_17641);
nand U18799 (N_18799,N_17084,N_17405);
nand U18800 (N_18800,N_17059,N_17759);
nand U18801 (N_18801,N_17626,N_17909);
nand U18802 (N_18802,N_17512,N_17677);
or U18803 (N_18803,N_17924,N_17752);
or U18804 (N_18804,N_17633,N_17229);
or U18805 (N_18805,N_17132,N_17145);
xor U18806 (N_18806,N_17063,N_17167);
and U18807 (N_18807,N_17650,N_17188);
or U18808 (N_18808,N_17091,N_17931);
xor U18809 (N_18809,N_17320,N_17278);
nor U18810 (N_18810,N_17357,N_17160);
and U18811 (N_18811,N_17599,N_17030);
xor U18812 (N_18812,N_17768,N_17975);
xnor U18813 (N_18813,N_17227,N_17425);
and U18814 (N_18814,N_17445,N_17735);
nor U18815 (N_18815,N_17154,N_17495);
and U18816 (N_18816,N_17066,N_17153);
nand U18817 (N_18817,N_17146,N_17853);
and U18818 (N_18818,N_17432,N_17910);
and U18819 (N_18819,N_17432,N_17374);
or U18820 (N_18820,N_17577,N_17840);
xnor U18821 (N_18821,N_17896,N_17464);
nor U18822 (N_18822,N_17162,N_17927);
and U18823 (N_18823,N_17403,N_17802);
nand U18824 (N_18824,N_17949,N_17708);
or U18825 (N_18825,N_17762,N_17757);
xnor U18826 (N_18826,N_17621,N_17671);
nor U18827 (N_18827,N_17160,N_17797);
xnor U18828 (N_18828,N_17825,N_17680);
and U18829 (N_18829,N_17046,N_17796);
xor U18830 (N_18830,N_17048,N_17553);
and U18831 (N_18831,N_17723,N_17624);
nand U18832 (N_18832,N_17077,N_17156);
nor U18833 (N_18833,N_17539,N_17824);
nor U18834 (N_18834,N_17255,N_17857);
xor U18835 (N_18835,N_17799,N_17338);
or U18836 (N_18836,N_17082,N_17808);
nor U18837 (N_18837,N_17295,N_17202);
nand U18838 (N_18838,N_17992,N_17886);
or U18839 (N_18839,N_17095,N_17502);
and U18840 (N_18840,N_17553,N_17387);
xnor U18841 (N_18841,N_17030,N_17778);
nand U18842 (N_18842,N_17086,N_17321);
nor U18843 (N_18843,N_17800,N_17515);
nand U18844 (N_18844,N_17827,N_17886);
nor U18845 (N_18845,N_17980,N_17297);
xnor U18846 (N_18846,N_17038,N_17441);
nand U18847 (N_18847,N_17152,N_17462);
nand U18848 (N_18848,N_17945,N_17874);
nor U18849 (N_18849,N_17751,N_17921);
nand U18850 (N_18850,N_17231,N_17030);
nand U18851 (N_18851,N_17992,N_17010);
and U18852 (N_18852,N_17738,N_17751);
nor U18853 (N_18853,N_17860,N_17458);
or U18854 (N_18854,N_17271,N_17715);
nor U18855 (N_18855,N_17625,N_17482);
nor U18856 (N_18856,N_17427,N_17391);
or U18857 (N_18857,N_17451,N_17997);
and U18858 (N_18858,N_17848,N_17945);
or U18859 (N_18859,N_17980,N_17676);
nor U18860 (N_18860,N_17924,N_17065);
nor U18861 (N_18861,N_17103,N_17404);
and U18862 (N_18862,N_17353,N_17311);
nor U18863 (N_18863,N_17281,N_17380);
nand U18864 (N_18864,N_17295,N_17038);
nor U18865 (N_18865,N_17961,N_17329);
nor U18866 (N_18866,N_17101,N_17029);
nand U18867 (N_18867,N_17461,N_17671);
xnor U18868 (N_18868,N_17247,N_17357);
and U18869 (N_18869,N_17601,N_17393);
nand U18870 (N_18870,N_17291,N_17498);
nand U18871 (N_18871,N_17241,N_17545);
nor U18872 (N_18872,N_17923,N_17667);
or U18873 (N_18873,N_17546,N_17449);
or U18874 (N_18874,N_17077,N_17667);
and U18875 (N_18875,N_17457,N_17888);
or U18876 (N_18876,N_17184,N_17083);
nand U18877 (N_18877,N_17327,N_17864);
and U18878 (N_18878,N_17581,N_17469);
nor U18879 (N_18879,N_17844,N_17598);
nand U18880 (N_18880,N_17088,N_17281);
nand U18881 (N_18881,N_17316,N_17093);
or U18882 (N_18882,N_17036,N_17376);
xnor U18883 (N_18883,N_17801,N_17482);
nand U18884 (N_18884,N_17713,N_17232);
and U18885 (N_18885,N_17024,N_17759);
or U18886 (N_18886,N_17614,N_17454);
nor U18887 (N_18887,N_17278,N_17380);
xnor U18888 (N_18888,N_17280,N_17414);
nor U18889 (N_18889,N_17961,N_17453);
nand U18890 (N_18890,N_17587,N_17406);
nand U18891 (N_18891,N_17384,N_17942);
and U18892 (N_18892,N_17542,N_17478);
xor U18893 (N_18893,N_17614,N_17735);
or U18894 (N_18894,N_17047,N_17459);
or U18895 (N_18895,N_17326,N_17698);
nor U18896 (N_18896,N_17011,N_17665);
xnor U18897 (N_18897,N_17186,N_17231);
and U18898 (N_18898,N_17204,N_17019);
and U18899 (N_18899,N_17297,N_17474);
xnor U18900 (N_18900,N_17315,N_17150);
xor U18901 (N_18901,N_17779,N_17093);
nand U18902 (N_18902,N_17264,N_17973);
xnor U18903 (N_18903,N_17665,N_17805);
nand U18904 (N_18904,N_17636,N_17188);
and U18905 (N_18905,N_17527,N_17826);
and U18906 (N_18906,N_17776,N_17713);
xor U18907 (N_18907,N_17006,N_17480);
or U18908 (N_18908,N_17906,N_17440);
xor U18909 (N_18909,N_17604,N_17236);
and U18910 (N_18910,N_17738,N_17883);
and U18911 (N_18911,N_17238,N_17889);
and U18912 (N_18912,N_17813,N_17806);
or U18913 (N_18913,N_17176,N_17384);
nor U18914 (N_18914,N_17648,N_17123);
xnor U18915 (N_18915,N_17603,N_17957);
or U18916 (N_18916,N_17513,N_17774);
xnor U18917 (N_18917,N_17360,N_17905);
or U18918 (N_18918,N_17094,N_17383);
and U18919 (N_18919,N_17098,N_17947);
xnor U18920 (N_18920,N_17290,N_17106);
and U18921 (N_18921,N_17073,N_17585);
nor U18922 (N_18922,N_17739,N_17218);
nand U18923 (N_18923,N_17647,N_17348);
nor U18924 (N_18924,N_17856,N_17961);
xnor U18925 (N_18925,N_17603,N_17274);
nand U18926 (N_18926,N_17089,N_17760);
nor U18927 (N_18927,N_17968,N_17646);
xnor U18928 (N_18928,N_17145,N_17209);
and U18929 (N_18929,N_17380,N_17745);
or U18930 (N_18930,N_17655,N_17559);
or U18931 (N_18931,N_17194,N_17953);
or U18932 (N_18932,N_17179,N_17470);
and U18933 (N_18933,N_17697,N_17572);
nor U18934 (N_18934,N_17216,N_17185);
and U18935 (N_18935,N_17400,N_17316);
xor U18936 (N_18936,N_17779,N_17709);
nand U18937 (N_18937,N_17110,N_17126);
nand U18938 (N_18938,N_17097,N_17706);
xor U18939 (N_18939,N_17019,N_17396);
nor U18940 (N_18940,N_17041,N_17377);
nor U18941 (N_18941,N_17208,N_17910);
or U18942 (N_18942,N_17344,N_17805);
xnor U18943 (N_18943,N_17654,N_17383);
and U18944 (N_18944,N_17850,N_17035);
xnor U18945 (N_18945,N_17644,N_17104);
xnor U18946 (N_18946,N_17955,N_17997);
and U18947 (N_18947,N_17968,N_17135);
nand U18948 (N_18948,N_17087,N_17652);
xnor U18949 (N_18949,N_17020,N_17164);
or U18950 (N_18950,N_17728,N_17354);
nand U18951 (N_18951,N_17343,N_17102);
nand U18952 (N_18952,N_17224,N_17246);
nor U18953 (N_18953,N_17023,N_17557);
nand U18954 (N_18954,N_17318,N_17777);
nand U18955 (N_18955,N_17273,N_17826);
nor U18956 (N_18956,N_17035,N_17144);
and U18957 (N_18957,N_17945,N_17322);
nand U18958 (N_18958,N_17871,N_17915);
nand U18959 (N_18959,N_17879,N_17898);
nand U18960 (N_18960,N_17765,N_17337);
nand U18961 (N_18961,N_17323,N_17009);
or U18962 (N_18962,N_17405,N_17515);
nor U18963 (N_18963,N_17676,N_17728);
nand U18964 (N_18964,N_17138,N_17654);
or U18965 (N_18965,N_17523,N_17530);
and U18966 (N_18966,N_17857,N_17289);
xnor U18967 (N_18967,N_17093,N_17718);
and U18968 (N_18968,N_17942,N_17480);
and U18969 (N_18969,N_17703,N_17006);
or U18970 (N_18970,N_17421,N_17499);
nand U18971 (N_18971,N_17834,N_17744);
nand U18972 (N_18972,N_17596,N_17084);
or U18973 (N_18973,N_17273,N_17285);
nand U18974 (N_18974,N_17711,N_17281);
nor U18975 (N_18975,N_17789,N_17282);
xor U18976 (N_18976,N_17148,N_17399);
nand U18977 (N_18977,N_17283,N_17606);
or U18978 (N_18978,N_17499,N_17755);
nor U18979 (N_18979,N_17998,N_17444);
nand U18980 (N_18980,N_17058,N_17636);
nand U18981 (N_18981,N_17885,N_17384);
and U18982 (N_18982,N_17157,N_17990);
xnor U18983 (N_18983,N_17830,N_17332);
nand U18984 (N_18984,N_17331,N_17432);
nand U18985 (N_18985,N_17925,N_17706);
nor U18986 (N_18986,N_17657,N_17214);
and U18987 (N_18987,N_17053,N_17743);
or U18988 (N_18988,N_17961,N_17169);
nor U18989 (N_18989,N_17979,N_17802);
or U18990 (N_18990,N_17569,N_17977);
xor U18991 (N_18991,N_17662,N_17753);
and U18992 (N_18992,N_17918,N_17917);
xnor U18993 (N_18993,N_17947,N_17201);
xnor U18994 (N_18994,N_17532,N_17863);
or U18995 (N_18995,N_17014,N_17060);
nor U18996 (N_18996,N_17026,N_17304);
nand U18997 (N_18997,N_17783,N_17029);
and U18998 (N_18998,N_17022,N_17215);
nand U18999 (N_18999,N_17685,N_17646);
xnor U19000 (N_19000,N_18018,N_18969);
nand U19001 (N_19001,N_18378,N_18586);
nor U19002 (N_19002,N_18487,N_18025);
or U19003 (N_19003,N_18235,N_18255);
xnor U19004 (N_19004,N_18281,N_18387);
and U19005 (N_19005,N_18654,N_18540);
nor U19006 (N_19006,N_18841,N_18858);
nor U19007 (N_19007,N_18633,N_18234);
xor U19008 (N_19008,N_18158,N_18127);
and U19009 (N_19009,N_18529,N_18853);
xor U19010 (N_19010,N_18419,N_18137);
nor U19011 (N_19011,N_18100,N_18140);
and U19012 (N_19012,N_18020,N_18056);
or U19013 (N_19013,N_18110,N_18222);
nor U19014 (N_19014,N_18108,N_18711);
or U19015 (N_19015,N_18927,N_18629);
and U19016 (N_19016,N_18545,N_18830);
nor U19017 (N_19017,N_18889,N_18400);
nand U19018 (N_19018,N_18785,N_18036);
or U19019 (N_19019,N_18202,N_18613);
xnor U19020 (N_19020,N_18257,N_18680);
nor U19021 (N_19021,N_18074,N_18526);
nand U19022 (N_19022,N_18209,N_18998);
xnor U19023 (N_19023,N_18031,N_18571);
xnor U19024 (N_19024,N_18005,N_18673);
nand U19025 (N_19025,N_18669,N_18747);
xnor U19026 (N_19026,N_18008,N_18648);
xor U19027 (N_19027,N_18809,N_18489);
xor U19028 (N_19028,N_18563,N_18188);
nor U19029 (N_19029,N_18765,N_18482);
and U19030 (N_19030,N_18694,N_18362);
xnor U19031 (N_19031,N_18186,N_18123);
nor U19032 (N_19032,N_18631,N_18535);
or U19033 (N_19033,N_18312,N_18187);
nand U19034 (N_19034,N_18849,N_18471);
xnor U19035 (N_19035,N_18945,N_18180);
nor U19036 (N_19036,N_18626,N_18182);
and U19037 (N_19037,N_18501,N_18878);
nor U19038 (N_19038,N_18498,N_18951);
nor U19039 (N_19039,N_18383,N_18195);
and U19040 (N_19040,N_18173,N_18065);
and U19041 (N_19041,N_18908,N_18308);
and U19042 (N_19042,N_18178,N_18617);
xnor U19043 (N_19043,N_18455,N_18179);
nor U19044 (N_19044,N_18033,N_18472);
nand U19045 (N_19045,N_18043,N_18363);
or U19046 (N_19046,N_18344,N_18491);
nor U19047 (N_19047,N_18475,N_18875);
nor U19048 (N_19048,N_18652,N_18810);
nand U19049 (N_19049,N_18190,N_18463);
or U19050 (N_19050,N_18721,N_18358);
and U19051 (N_19051,N_18985,N_18439);
or U19052 (N_19052,N_18211,N_18200);
xnor U19053 (N_19053,N_18464,N_18611);
nor U19054 (N_19054,N_18650,N_18960);
nand U19055 (N_19055,N_18585,N_18288);
xnor U19056 (N_19056,N_18414,N_18684);
nor U19057 (N_19057,N_18843,N_18405);
nor U19058 (N_19058,N_18607,N_18800);
and U19059 (N_19059,N_18176,N_18700);
or U19060 (N_19060,N_18445,N_18638);
nor U19061 (N_19061,N_18223,N_18547);
nor U19062 (N_19062,N_18499,N_18208);
and U19063 (N_19063,N_18636,N_18225);
and U19064 (N_19064,N_18032,N_18253);
and U19065 (N_19065,N_18592,N_18321);
and U19066 (N_19066,N_18608,N_18012);
xor U19067 (N_19067,N_18635,N_18512);
nand U19068 (N_19068,N_18041,N_18242);
or U19069 (N_19069,N_18194,N_18888);
or U19070 (N_19070,N_18437,N_18250);
or U19071 (N_19071,N_18885,N_18978);
or U19072 (N_19072,N_18278,N_18566);
xnor U19073 (N_19073,N_18207,N_18319);
or U19074 (N_19074,N_18460,N_18133);
nor U19075 (N_19075,N_18391,N_18569);
and U19076 (N_19076,N_18047,N_18609);
or U19077 (N_19077,N_18593,N_18160);
xor U19078 (N_19078,N_18089,N_18500);
or U19079 (N_19079,N_18000,N_18465);
or U19080 (N_19080,N_18384,N_18456);
or U19081 (N_19081,N_18283,N_18453);
xor U19082 (N_19082,N_18552,N_18597);
xor U19083 (N_19083,N_18594,N_18856);
nand U19084 (N_19084,N_18393,N_18165);
xor U19085 (N_19085,N_18766,N_18351);
nor U19086 (N_19086,N_18360,N_18958);
xnor U19087 (N_19087,N_18861,N_18599);
or U19088 (N_19088,N_18997,N_18651);
nand U19089 (N_19089,N_18873,N_18521);
nor U19090 (N_19090,N_18659,N_18555);
nor U19091 (N_19091,N_18224,N_18893);
or U19092 (N_19092,N_18917,N_18216);
or U19093 (N_19093,N_18963,N_18621);
or U19094 (N_19094,N_18928,N_18476);
xnor U19095 (N_19095,N_18877,N_18930);
nand U19096 (N_19096,N_18117,N_18356);
xnor U19097 (N_19097,N_18315,N_18138);
nand U19098 (N_19098,N_18480,N_18273);
and U19099 (N_19099,N_18851,N_18380);
and U19100 (N_19100,N_18144,N_18115);
and U19101 (N_19101,N_18227,N_18413);
and U19102 (N_19102,N_18107,N_18854);
and U19103 (N_19103,N_18516,N_18935);
or U19104 (N_19104,N_18582,N_18825);
nand U19105 (N_19105,N_18374,N_18554);
nor U19106 (N_19106,N_18090,N_18398);
or U19107 (N_19107,N_18723,N_18757);
or U19108 (N_19108,N_18709,N_18921);
nand U19109 (N_19109,N_18897,N_18708);
nand U19110 (N_19110,N_18579,N_18753);
or U19111 (N_19111,N_18092,N_18277);
nor U19112 (N_19112,N_18578,N_18995);
xor U19113 (N_19113,N_18497,N_18327);
nand U19114 (N_19114,N_18750,N_18191);
and U19115 (N_19115,N_18258,N_18086);
nand U19116 (N_19116,N_18287,N_18731);
nor U19117 (N_19117,N_18937,N_18306);
or U19118 (N_19118,N_18618,N_18347);
and U19119 (N_19119,N_18733,N_18639);
and U19120 (N_19120,N_18063,N_18401);
nand U19121 (N_19121,N_18204,N_18411);
xnor U19122 (N_19122,N_18040,N_18666);
nor U19123 (N_19123,N_18355,N_18271);
nor U19124 (N_19124,N_18403,N_18729);
nor U19125 (N_19125,N_18418,N_18381);
xor U19126 (N_19126,N_18167,N_18519);
xor U19127 (N_19127,N_18890,N_18442);
xor U19128 (N_19128,N_18798,N_18932);
or U19129 (N_19129,N_18506,N_18131);
nand U19130 (N_19130,N_18541,N_18241);
and U19131 (N_19131,N_18598,N_18425);
nand U19132 (N_19132,N_18551,N_18075);
nand U19133 (N_19133,N_18432,N_18857);
nor U19134 (N_19134,N_18793,N_18902);
or U19135 (N_19135,N_18901,N_18938);
or U19136 (N_19136,N_18295,N_18249);
nor U19137 (N_19137,N_18615,N_18048);
and U19138 (N_19138,N_18130,N_18244);
nor U19139 (N_19139,N_18762,N_18256);
nor U19140 (N_19140,N_18574,N_18185);
or U19141 (N_19141,N_18988,N_18286);
or U19142 (N_19142,N_18795,N_18007);
or U19143 (N_19143,N_18697,N_18316);
and U19144 (N_19144,N_18221,N_18368);
nand U19145 (N_19145,N_18270,N_18916);
xor U19146 (N_19146,N_18028,N_18451);
nor U19147 (N_19147,N_18296,N_18324);
and U19148 (N_19148,N_18397,N_18903);
xor U19149 (N_19149,N_18674,N_18198);
and U19150 (N_19150,N_18965,N_18860);
xor U19151 (N_19151,N_18948,N_18070);
xor U19152 (N_19152,N_18575,N_18304);
or U19153 (N_19153,N_18657,N_18494);
nor U19154 (N_19154,N_18004,N_18424);
nor U19155 (N_19155,N_18058,N_18748);
and U19156 (N_19156,N_18534,N_18559);
or U19157 (N_19157,N_18022,N_18136);
nand U19158 (N_19158,N_18490,N_18293);
xnor U19159 (N_19159,N_18911,N_18794);
xor U19160 (N_19160,N_18730,N_18396);
nand U19161 (N_19161,N_18971,N_18077);
nor U19162 (N_19162,N_18299,N_18701);
nor U19163 (N_19163,N_18620,N_18745);
nor U19164 (N_19164,N_18104,N_18996);
xor U19165 (N_19165,N_18936,N_18081);
nor U19166 (N_19166,N_18205,N_18964);
or U19167 (N_19167,N_18514,N_18759);
nand U19168 (N_19168,N_18752,N_18011);
and U19169 (N_19169,N_18504,N_18538);
xnor U19170 (N_19170,N_18703,N_18828);
or U19171 (N_19171,N_18069,N_18778);
nand U19172 (N_19172,N_18436,N_18850);
nand U19173 (N_19173,N_18820,N_18565);
or U19174 (N_19174,N_18839,N_18737);
or U19175 (N_19175,N_18412,N_18163);
nor U19176 (N_19176,N_18807,N_18643);
nand U19177 (N_19177,N_18478,N_18884);
nor U19178 (N_19178,N_18251,N_18789);
and U19179 (N_19179,N_18727,N_18433);
or U19180 (N_19180,N_18966,N_18803);
xor U19181 (N_19181,N_18001,N_18999);
and U19182 (N_19182,N_18226,N_18975);
or U19183 (N_19183,N_18658,N_18972);
or U19184 (N_19184,N_18931,N_18170);
nand U19185 (N_19185,N_18894,N_18738);
nor U19186 (N_19186,N_18863,N_18683);
nor U19187 (N_19187,N_18953,N_18263);
nor U19188 (N_19188,N_18670,N_18819);
or U19189 (N_19189,N_18328,N_18831);
or U19190 (N_19190,N_18905,N_18307);
nor U19191 (N_19191,N_18823,N_18580);
or U19192 (N_19192,N_18764,N_18059);
nand U19193 (N_19193,N_18647,N_18605);
and U19194 (N_19194,N_18103,N_18623);
and U19195 (N_19195,N_18663,N_18015);
nor U19196 (N_19196,N_18461,N_18014);
nor U19197 (N_19197,N_18606,N_18320);
xor U19198 (N_19198,N_18685,N_18749);
xnor U19199 (N_19199,N_18335,N_18238);
xor U19200 (N_19200,N_18044,N_18030);
nand U19201 (N_19201,N_18183,N_18084);
nor U19202 (N_19202,N_18175,N_18950);
xnor U19203 (N_19203,N_18595,N_18724);
xnor U19204 (N_19204,N_18002,N_18681);
or U19205 (N_19205,N_18228,N_18072);
or U19206 (N_19206,N_18024,N_18912);
and U19207 (N_19207,N_18229,N_18062);
nand U19208 (N_19208,N_18247,N_18852);
and U19209 (N_19209,N_18051,N_18172);
nor U19210 (N_19210,N_18054,N_18784);
xnor U19211 (N_19211,N_18233,N_18556);
nor U19212 (N_19212,N_18976,N_18502);
nor U19213 (N_19213,N_18758,N_18267);
xnor U19214 (N_19214,N_18375,N_18243);
nand U19215 (N_19215,N_18067,N_18675);
nor U19216 (N_19216,N_18678,N_18477);
nor U19217 (N_19217,N_18317,N_18768);
and U19218 (N_19218,N_18435,N_18907);
nor U19219 (N_19219,N_18218,N_18632);
xor U19220 (N_19220,N_18408,N_18539);
nand U19221 (N_19221,N_18154,N_18332);
nor U19222 (N_19222,N_18818,N_18874);
or U19223 (N_19223,N_18164,N_18981);
nor U19224 (N_19224,N_18336,N_18867);
nor U19225 (N_19225,N_18899,N_18508);
or U19226 (N_19226,N_18513,N_18676);
or U19227 (N_19227,N_18532,N_18290);
nor U19228 (N_19228,N_18441,N_18664);
nor U19229 (N_19229,N_18704,N_18584);
nor U19230 (N_19230,N_18409,N_18716);
nand U19231 (N_19231,N_18872,N_18956);
and U19232 (N_19232,N_18796,N_18359);
nand U19233 (N_19233,N_18952,N_18904);
and U19234 (N_19234,N_18760,N_18845);
and U19235 (N_19235,N_18630,N_18339);
nor U19236 (N_19236,N_18589,N_18797);
or U19237 (N_19237,N_18248,N_18744);
nor U19238 (N_19238,N_18864,N_18369);
nand U19239 (N_19239,N_18943,N_18832);
nand U19240 (N_19240,N_18771,N_18686);
nor U19241 (N_19241,N_18447,N_18604);
xnor U19242 (N_19242,N_18641,N_18614);
nor U19243 (N_19243,N_18483,N_18155);
or U19244 (N_19244,N_18741,N_18564);
or U19245 (N_19245,N_18919,N_18707);
and U19246 (N_19246,N_18720,N_18364);
and U19247 (N_19247,N_18511,N_18121);
nand U19248 (N_19248,N_18157,N_18990);
and U19249 (N_19249,N_18725,N_18168);
nor U19250 (N_19250,N_18992,N_18993);
nor U19251 (N_19251,N_18891,N_18236);
xor U19252 (N_19252,N_18786,N_18974);
and U19253 (N_19253,N_18496,N_18017);
nor U19254 (N_19254,N_18660,N_18662);
xnor U19255 (N_19255,N_18833,N_18169);
or U19256 (N_19256,N_18029,N_18610);
nor U19257 (N_19257,N_18109,N_18349);
xor U19258 (N_19258,N_18780,N_18634);
nor U19259 (N_19259,N_18313,N_18151);
and U19260 (N_19260,N_18091,N_18791);
xor U19261 (N_19261,N_18314,N_18991);
nor U19262 (N_19262,N_18746,N_18297);
or U19263 (N_19263,N_18543,N_18824);
nor U19264 (N_19264,N_18377,N_18934);
nor U19265 (N_19265,N_18444,N_18423);
xor U19266 (N_19266,N_18944,N_18779);
nor U19267 (N_19267,N_18417,N_18101);
xor U19268 (N_19268,N_18881,N_18060);
nor U19269 (N_19269,N_18019,N_18240);
nand U19270 (N_19270,N_18812,N_18548);
nor U19271 (N_19271,N_18331,N_18612);
nor U19272 (N_19272,N_18021,N_18459);
nand U19273 (N_19273,N_18772,N_18147);
and U19274 (N_19274,N_18879,N_18027);
nand U19275 (N_19275,N_18531,N_18755);
and U19276 (N_19276,N_18341,N_18135);
or U19277 (N_19277,N_18231,N_18206);
xor U19278 (N_19278,N_18484,N_18805);
nand U19279 (N_19279,N_18279,N_18994);
nand U19280 (N_19280,N_18836,N_18695);
xor U19281 (N_19281,N_18064,N_18653);
nand U19282 (N_19282,N_18003,N_18406);
nand U19283 (N_19283,N_18835,N_18602);
nand U19284 (N_19284,N_18149,N_18311);
or U19285 (N_19285,N_18189,N_18310);
xnor U19286 (N_19286,N_18365,N_18237);
and U19287 (N_19287,N_18132,N_18376);
xnor U19288 (N_19288,N_18220,N_18410);
or U19289 (N_19289,N_18567,N_18705);
nor U19290 (N_19290,N_18118,N_18503);
xor U19291 (N_19291,N_18458,N_18714);
nor U19292 (N_19292,N_18688,N_18473);
nand U19293 (N_19293,N_18537,N_18390);
nor U19294 (N_19294,N_18426,N_18192);
nand U19295 (N_19295,N_18949,N_18790);
or U19296 (N_19296,N_18855,N_18718);
nand U19297 (N_19297,N_18918,N_18106);
xnor U19298 (N_19298,N_18834,N_18470);
nor U19299 (N_19299,N_18016,N_18334);
nand U19300 (N_19300,N_18034,N_18361);
xor U19301 (N_19301,N_18507,N_18468);
or U19302 (N_19302,N_18122,N_18479);
or U19303 (N_19303,N_18385,N_18910);
xnor U19304 (N_19304,N_18536,N_18079);
or U19305 (N_19305,N_18126,N_18722);
nor U19306 (N_19306,N_18125,N_18085);
xnor U19307 (N_19307,N_18838,N_18712);
or U19308 (N_19308,N_18914,N_18583);
xor U19309 (N_19309,N_18333,N_18624);
nor U19310 (N_19310,N_18804,N_18906);
xnor U19311 (N_19311,N_18026,N_18230);
or U19312 (N_19312,N_18120,N_18428);
or U19313 (N_19313,N_18525,N_18773);
nor U19314 (N_19314,N_18469,N_18171);
or U19315 (N_19315,N_18862,N_18742);
xnor U19316 (N_19316,N_18869,N_18865);
nand U19317 (N_19317,N_18300,N_18053);
nand U19318 (N_19318,N_18038,N_18429);
and U19319 (N_19319,N_18098,N_18071);
nand U19320 (N_19320,N_18268,N_18119);
nand U19321 (N_19321,N_18808,N_18649);
xnor U19322 (N_19322,N_18156,N_18046);
and U19323 (N_19323,N_18495,N_18099);
and U19324 (N_19324,N_18734,N_18987);
xnor U19325 (N_19325,N_18061,N_18340);
or U19326 (N_19326,N_18751,N_18337);
nand U19327 (N_19327,N_18252,N_18726);
nor U19328 (N_19328,N_18719,N_18967);
nand U19329 (N_19329,N_18811,N_18939);
and U19330 (N_19330,N_18260,N_18350);
nand U19331 (N_19331,N_18285,N_18619);
nand U19332 (N_19332,N_18049,N_18212);
xor U19333 (N_19333,N_18925,N_18407);
nand U19334 (N_19334,N_18097,N_18915);
nor U19335 (N_19335,N_18481,N_18421);
or U19336 (N_19336,N_18754,N_18962);
nor U19337 (N_19337,N_18245,N_18449);
or U19338 (N_19338,N_18146,N_18045);
or U19339 (N_19339,N_18474,N_18422);
or U19340 (N_19340,N_18023,N_18427);
nand U19341 (N_19341,N_18682,N_18148);
xor U19342 (N_19342,N_18774,N_18627);
xnor U19343 (N_19343,N_18710,N_18467);
or U19344 (N_19344,N_18736,N_18094);
and U19345 (N_19345,N_18560,N_18184);
or U19346 (N_19346,N_18886,N_18052);
nor U19347 (N_19347,N_18616,N_18769);
xnor U19348 (N_19348,N_18518,N_18983);
nand U19349 (N_19349,N_18896,N_18326);
nor U19350 (N_19350,N_18039,N_18305);
or U19351 (N_19351,N_18083,N_18799);
nor U19352 (N_19352,N_18761,N_18544);
xnor U19353 (N_19353,N_18706,N_18389);
nand U19354 (N_19354,N_18989,N_18573);
or U19355 (N_19355,N_18438,N_18940);
or U19356 (N_19356,N_18197,N_18876);
nor U19357 (N_19357,N_18542,N_18457);
and U19358 (N_19358,N_18093,N_18066);
xnor U19359 (N_19359,N_18550,N_18371);
xor U19360 (N_19360,N_18837,N_18388);
nor U19361 (N_19361,N_18174,N_18517);
nand U19362 (N_19362,N_18139,N_18450);
or U19363 (N_19363,N_18942,N_18342);
xnor U19364 (N_19364,N_18309,N_18715);
or U19365 (N_19365,N_18303,N_18367);
or U19366 (N_19366,N_18883,N_18984);
and U19367 (N_19367,N_18493,N_18770);
nand U19368 (N_19368,N_18338,N_18096);
nand U19369 (N_19369,N_18203,N_18354);
nand U19370 (N_19370,N_18177,N_18254);
nor U19371 (N_19371,N_18848,N_18275);
or U19372 (N_19372,N_18214,N_18352);
nand U19373 (N_19373,N_18510,N_18166);
or U19374 (N_19374,N_18814,N_18846);
nand U19375 (N_19375,N_18699,N_18870);
nor U19376 (N_19376,N_18829,N_18679);
nor U19377 (N_19377,N_18922,N_18325);
xnor U19378 (N_19378,N_18923,N_18530);
nor U19379 (N_19379,N_18150,N_18392);
xor U19380 (N_19380,N_18454,N_18842);
xnor U19381 (N_19381,N_18581,N_18961);
nand U19382 (N_19382,N_18576,N_18871);
nor U19383 (N_19383,N_18522,N_18929);
and U19384 (N_19384,N_18215,N_18440);
xnor U19385 (N_19385,N_18057,N_18880);
xnor U19386 (N_19386,N_18199,N_18691);
xor U19387 (N_19387,N_18520,N_18196);
xor U19388 (N_19388,N_18161,N_18646);
nor U19389 (N_19389,N_18006,N_18900);
nor U19390 (N_19390,N_18159,N_18667);
nand U19391 (N_19391,N_18739,N_18527);
xor U19392 (N_19392,N_18394,N_18775);
and U19393 (N_19393,N_18515,N_18628);
and U19394 (N_19394,N_18698,N_18524);
xnor U19395 (N_19395,N_18399,N_18859);
nor U19396 (N_19396,N_18078,N_18783);
or U19397 (N_19397,N_18042,N_18372);
nand U19398 (N_19398,N_18558,N_18462);
nor U19399 (N_19399,N_18088,N_18591);
xnor U19400 (N_19400,N_18272,N_18111);
nor U19401 (N_19401,N_18280,N_18213);
nand U19402 (N_19402,N_18767,N_18553);
xor U19403 (N_19403,N_18416,N_18142);
nor U19404 (N_19404,N_18665,N_18112);
and U19405 (N_19405,N_18282,N_18322);
nor U19406 (N_19406,N_18386,N_18348);
or U19407 (N_19407,N_18134,N_18973);
nor U19408 (N_19408,N_18920,N_18289);
and U19409 (N_19409,N_18162,N_18847);
xnor U19410 (N_19410,N_18821,N_18827);
or U19411 (N_19411,N_18264,N_18924);
nor U19412 (N_19412,N_18909,N_18055);
or U19413 (N_19413,N_18080,N_18587);
nand U19414 (N_19414,N_18979,N_18702);
nand U19415 (N_19415,N_18590,N_18370);
nand U19416 (N_19416,N_18181,N_18404);
or U19417 (N_19417,N_18642,N_18588);
nor U19418 (N_19418,N_18068,N_18343);
or U19419 (N_19419,N_18274,N_18728);
nand U19420 (N_19420,N_18672,N_18219);
nor U19421 (N_19421,N_18815,N_18687);
nand U19422 (N_19422,N_18128,N_18986);
and U19423 (N_19423,N_18596,N_18010);
and U19424 (N_19424,N_18941,N_18145);
nor U19425 (N_19425,N_18776,N_18210);
or U19426 (N_19426,N_18265,N_18201);
xor U19427 (N_19427,N_18301,N_18866);
nand U19428 (N_19428,N_18913,N_18382);
nor U19429 (N_19429,N_18129,N_18193);
or U19430 (N_19430,N_18346,N_18671);
or U19431 (N_19431,N_18792,N_18353);
and U19432 (N_19432,N_18577,N_18345);
nand U19433 (N_19433,N_18640,N_18488);
nand U19434 (N_19434,N_18844,N_18806);
and U19435 (N_19435,N_18957,N_18717);
or U19436 (N_19436,N_18082,N_18625);
nor U19437 (N_19437,N_18645,N_18102);
xnor U19438 (N_19438,N_18505,N_18677);
nor U19439 (N_19439,N_18696,N_18466);
or U19440 (N_19440,N_18415,N_18743);
nor U19441 (N_19441,N_18143,N_18968);
or U19442 (N_19442,N_18239,N_18269);
xor U19443 (N_19443,N_18690,N_18492);
xnor U19444 (N_19444,N_18402,N_18732);
or U19445 (N_19445,N_18452,N_18232);
xor U19446 (N_19446,N_18318,N_18561);
or U19447 (N_19447,N_18813,N_18954);
and U19448 (N_19448,N_18114,N_18892);
and U19449 (N_19449,N_18693,N_18259);
or U19450 (N_19450,N_18485,N_18357);
xnor U19451 (N_19451,N_18443,N_18486);
nor U19452 (N_19452,N_18959,N_18735);
nor U19453 (N_19453,N_18970,N_18777);
and U19454 (N_19454,N_18087,N_18124);
or U19455 (N_19455,N_18882,N_18266);
xor U19456 (N_19456,N_18946,N_18509);
nand U19457 (N_19457,N_18528,N_18141);
nand U19458 (N_19458,N_18366,N_18262);
and U19459 (N_19459,N_18373,N_18816);
and U19460 (N_19460,N_18050,N_18603);
nor U19461 (N_19461,N_18546,N_18955);
nor U19462 (N_19462,N_18644,N_18713);
and U19463 (N_19463,N_18787,N_18763);
nand U19464 (N_19464,N_18622,N_18740);
nand U19465 (N_19465,N_18840,N_18073);
or U19466 (N_19466,N_18379,N_18562);
xor U19467 (N_19467,N_18009,N_18298);
xnor U19468 (N_19468,N_18668,N_18898);
xnor U19469 (N_19469,N_18330,N_18116);
nand U19470 (N_19470,N_18568,N_18656);
nand U19471 (N_19471,N_18113,N_18980);
nand U19472 (N_19472,N_18826,N_18933);
and U19473 (N_19473,N_18431,N_18095);
nand U19474 (N_19474,N_18637,N_18801);
nor U19475 (N_19475,N_18261,N_18692);
or U19476 (N_19476,N_18395,N_18868);
nand U19477 (N_19477,N_18788,N_18782);
xnor U19478 (N_19478,N_18802,N_18291);
or U19479 (N_19479,N_18246,N_18781);
nor U19480 (N_19480,N_18977,N_18817);
nand U19481 (N_19481,N_18292,N_18570);
xnor U19482 (N_19482,N_18982,N_18895);
nor U19483 (N_19483,N_18655,N_18523);
nand U19484 (N_19484,N_18600,N_18430);
and U19485 (N_19485,N_18557,N_18329);
nand U19486 (N_19486,N_18035,N_18420);
xor U19487 (N_19487,N_18689,N_18302);
xor U19488 (N_19488,N_18217,N_18037);
or U19489 (N_19489,N_18601,N_18284);
or U19490 (N_19490,N_18887,N_18926);
nand U19491 (N_19491,N_18076,N_18276);
nor U19492 (N_19492,N_18446,N_18152);
nand U19493 (N_19493,N_18323,N_18822);
nor U19494 (N_19494,N_18661,N_18153);
nor U19495 (N_19495,N_18434,N_18549);
or U19496 (N_19496,N_18533,N_18756);
xnor U19497 (N_19497,N_18947,N_18448);
xnor U19498 (N_19498,N_18013,N_18572);
nand U19499 (N_19499,N_18294,N_18105);
or U19500 (N_19500,N_18631,N_18353);
and U19501 (N_19501,N_18333,N_18875);
and U19502 (N_19502,N_18578,N_18582);
nand U19503 (N_19503,N_18417,N_18165);
or U19504 (N_19504,N_18918,N_18538);
or U19505 (N_19505,N_18203,N_18812);
and U19506 (N_19506,N_18933,N_18835);
xnor U19507 (N_19507,N_18991,N_18276);
xor U19508 (N_19508,N_18266,N_18344);
and U19509 (N_19509,N_18403,N_18284);
xor U19510 (N_19510,N_18156,N_18766);
xor U19511 (N_19511,N_18463,N_18777);
and U19512 (N_19512,N_18691,N_18116);
xnor U19513 (N_19513,N_18539,N_18769);
xor U19514 (N_19514,N_18927,N_18604);
nor U19515 (N_19515,N_18274,N_18623);
and U19516 (N_19516,N_18864,N_18791);
nand U19517 (N_19517,N_18256,N_18509);
nand U19518 (N_19518,N_18715,N_18708);
or U19519 (N_19519,N_18338,N_18681);
and U19520 (N_19520,N_18463,N_18548);
nor U19521 (N_19521,N_18848,N_18533);
xnor U19522 (N_19522,N_18775,N_18800);
or U19523 (N_19523,N_18601,N_18260);
or U19524 (N_19524,N_18835,N_18172);
or U19525 (N_19525,N_18220,N_18203);
nor U19526 (N_19526,N_18892,N_18488);
nand U19527 (N_19527,N_18358,N_18735);
nor U19528 (N_19528,N_18323,N_18165);
nor U19529 (N_19529,N_18842,N_18166);
xor U19530 (N_19530,N_18143,N_18541);
xor U19531 (N_19531,N_18425,N_18117);
and U19532 (N_19532,N_18730,N_18776);
and U19533 (N_19533,N_18871,N_18696);
or U19534 (N_19534,N_18373,N_18033);
xor U19535 (N_19535,N_18117,N_18796);
nand U19536 (N_19536,N_18784,N_18762);
or U19537 (N_19537,N_18434,N_18351);
nand U19538 (N_19538,N_18054,N_18802);
and U19539 (N_19539,N_18370,N_18287);
xor U19540 (N_19540,N_18382,N_18619);
and U19541 (N_19541,N_18585,N_18855);
and U19542 (N_19542,N_18631,N_18038);
or U19543 (N_19543,N_18137,N_18464);
nand U19544 (N_19544,N_18258,N_18311);
and U19545 (N_19545,N_18577,N_18885);
nor U19546 (N_19546,N_18656,N_18688);
xor U19547 (N_19547,N_18180,N_18085);
and U19548 (N_19548,N_18653,N_18957);
nand U19549 (N_19549,N_18826,N_18481);
nand U19550 (N_19550,N_18519,N_18210);
nand U19551 (N_19551,N_18649,N_18682);
xnor U19552 (N_19552,N_18440,N_18991);
nand U19553 (N_19553,N_18480,N_18900);
nor U19554 (N_19554,N_18698,N_18334);
and U19555 (N_19555,N_18812,N_18534);
xor U19556 (N_19556,N_18844,N_18269);
nor U19557 (N_19557,N_18063,N_18483);
or U19558 (N_19558,N_18068,N_18783);
nor U19559 (N_19559,N_18610,N_18045);
and U19560 (N_19560,N_18928,N_18955);
or U19561 (N_19561,N_18729,N_18535);
or U19562 (N_19562,N_18634,N_18307);
nor U19563 (N_19563,N_18491,N_18085);
or U19564 (N_19564,N_18760,N_18852);
or U19565 (N_19565,N_18160,N_18224);
xnor U19566 (N_19566,N_18883,N_18746);
xor U19567 (N_19567,N_18962,N_18220);
nor U19568 (N_19568,N_18652,N_18243);
or U19569 (N_19569,N_18201,N_18296);
xor U19570 (N_19570,N_18493,N_18500);
nand U19571 (N_19571,N_18472,N_18942);
nand U19572 (N_19572,N_18676,N_18626);
nand U19573 (N_19573,N_18854,N_18376);
nor U19574 (N_19574,N_18313,N_18913);
nand U19575 (N_19575,N_18443,N_18436);
or U19576 (N_19576,N_18303,N_18547);
and U19577 (N_19577,N_18122,N_18105);
xor U19578 (N_19578,N_18404,N_18445);
xnor U19579 (N_19579,N_18493,N_18786);
or U19580 (N_19580,N_18643,N_18076);
xor U19581 (N_19581,N_18275,N_18214);
nor U19582 (N_19582,N_18027,N_18633);
nand U19583 (N_19583,N_18367,N_18232);
and U19584 (N_19584,N_18430,N_18598);
nor U19585 (N_19585,N_18545,N_18415);
nor U19586 (N_19586,N_18194,N_18120);
and U19587 (N_19587,N_18542,N_18632);
and U19588 (N_19588,N_18493,N_18244);
xor U19589 (N_19589,N_18750,N_18536);
nor U19590 (N_19590,N_18449,N_18683);
xnor U19591 (N_19591,N_18078,N_18253);
xnor U19592 (N_19592,N_18415,N_18560);
or U19593 (N_19593,N_18303,N_18265);
xor U19594 (N_19594,N_18089,N_18176);
or U19595 (N_19595,N_18230,N_18758);
nor U19596 (N_19596,N_18298,N_18672);
or U19597 (N_19597,N_18958,N_18887);
xor U19598 (N_19598,N_18949,N_18396);
or U19599 (N_19599,N_18827,N_18243);
xnor U19600 (N_19600,N_18116,N_18908);
or U19601 (N_19601,N_18928,N_18268);
xnor U19602 (N_19602,N_18074,N_18685);
xor U19603 (N_19603,N_18150,N_18661);
or U19604 (N_19604,N_18844,N_18917);
or U19605 (N_19605,N_18238,N_18443);
nand U19606 (N_19606,N_18982,N_18393);
nor U19607 (N_19607,N_18574,N_18689);
xnor U19608 (N_19608,N_18731,N_18178);
nor U19609 (N_19609,N_18529,N_18081);
nor U19610 (N_19610,N_18298,N_18336);
xor U19611 (N_19611,N_18557,N_18683);
or U19612 (N_19612,N_18422,N_18405);
nor U19613 (N_19613,N_18180,N_18894);
nand U19614 (N_19614,N_18693,N_18231);
xnor U19615 (N_19615,N_18680,N_18669);
or U19616 (N_19616,N_18910,N_18923);
xor U19617 (N_19617,N_18205,N_18464);
or U19618 (N_19618,N_18841,N_18490);
nor U19619 (N_19619,N_18606,N_18904);
nand U19620 (N_19620,N_18571,N_18469);
nor U19621 (N_19621,N_18857,N_18700);
or U19622 (N_19622,N_18298,N_18731);
nand U19623 (N_19623,N_18245,N_18390);
and U19624 (N_19624,N_18252,N_18456);
nor U19625 (N_19625,N_18494,N_18212);
and U19626 (N_19626,N_18326,N_18524);
nor U19627 (N_19627,N_18979,N_18519);
nor U19628 (N_19628,N_18492,N_18208);
and U19629 (N_19629,N_18523,N_18331);
nor U19630 (N_19630,N_18880,N_18526);
nor U19631 (N_19631,N_18316,N_18014);
and U19632 (N_19632,N_18774,N_18250);
and U19633 (N_19633,N_18827,N_18753);
xor U19634 (N_19634,N_18011,N_18196);
nor U19635 (N_19635,N_18778,N_18018);
nand U19636 (N_19636,N_18601,N_18304);
and U19637 (N_19637,N_18310,N_18136);
or U19638 (N_19638,N_18724,N_18203);
and U19639 (N_19639,N_18137,N_18477);
or U19640 (N_19640,N_18956,N_18148);
or U19641 (N_19641,N_18334,N_18247);
or U19642 (N_19642,N_18376,N_18086);
xor U19643 (N_19643,N_18628,N_18924);
and U19644 (N_19644,N_18253,N_18344);
or U19645 (N_19645,N_18813,N_18600);
and U19646 (N_19646,N_18571,N_18351);
nand U19647 (N_19647,N_18398,N_18377);
nand U19648 (N_19648,N_18116,N_18501);
xor U19649 (N_19649,N_18013,N_18356);
nand U19650 (N_19650,N_18406,N_18886);
or U19651 (N_19651,N_18560,N_18706);
or U19652 (N_19652,N_18561,N_18529);
xor U19653 (N_19653,N_18144,N_18795);
nor U19654 (N_19654,N_18839,N_18551);
nand U19655 (N_19655,N_18034,N_18978);
or U19656 (N_19656,N_18144,N_18234);
nor U19657 (N_19657,N_18547,N_18135);
xor U19658 (N_19658,N_18212,N_18752);
nor U19659 (N_19659,N_18723,N_18622);
xnor U19660 (N_19660,N_18035,N_18761);
xnor U19661 (N_19661,N_18316,N_18882);
nor U19662 (N_19662,N_18307,N_18958);
or U19663 (N_19663,N_18147,N_18936);
nand U19664 (N_19664,N_18403,N_18387);
xor U19665 (N_19665,N_18385,N_18489);
or U19666 (N_19666,N_18301,N_18082);
nand U19667 (N_19667,N_18307,N_18565);
xor U19668 (N_19668,N_18008,N_18754);
nand U19669 (N_19669,N_18640,N_18596);
nand U19670 (N_19670,N_18835,N_18207);
nor U19671 (N_19671,N_18791,N_18744);
nand U19672 (N_19672,N_18448,N_18672);
or U19673 (N_19673,N_18211,N_18281);
nor U19674 (N_19674,N_18751,N_18169);
and U19675 (N_19675,N_18828,N_18719);
or U19676 (N_19676,N_18342,N_18849);
and U19677 (N_19677,N_18816,N_18224);
or U19678 (N_19678,N_18507,N_18070);
or U19679 (N_19679,N_18140,N_18654);
nor U19680 (N_19680,N_18012,N_18325);
and U19681 (N_19681,N_18462,N_18864);
nor U19682 (N_19682,N_18915,N_18077);
nand U19683 (N_19683,N_18568,N_18735);
or U19684 (N_19684,N_18356,N_18780);
and U19685 (N_19685,N_18846,N_18161);
xor U19686 (N_19686,N_18850,N_18388);
nand U19687 (N_19687,N_18443,N_18924);
or U19688 (N_19688,N_18448,N_18229);
nand U19689 (N_19689,N_18333,N_18491);
and U19690 (N_19690,N_18809,N_18423);
and U19691 (N_19691,N_18122,N_18882);
xor U19692 (N_19692,N_18815,N_18415);
and U19693 (N_19693,N_18997,N_18673);
nand U19694 (N_19694,N_18057,N_18873);
and U19695 (N_19695,N_18657,N_18759);
xor U19696 (N_19696,N_18960,N_18080);
or U19697 (N_19697,N_18727,N_18529);
nand U19698 (N_19698,N_18000,N_18288);
nand U19699 (N_19699,N_18674,N_18841);
or U19700 (N_19700,N_18201,N_18895);
nor U19701 (N_19701,N_18744,N_18296);
nand U19702 (N_19702,N_18285,N_18932);
xor U19703 (N_19703,N_18641,N_18134);
and U19704 (N_19704,N_18727,N_18371);
nor U19705 (N_19705,N_18788,N_18796);
and U19706 (N_19706,N_18445,N_18956);
nor U19707 (N_19707,N_18925,N_18022);
nand U19708 (N_19708,N_18506,N_18935);
nor U19709 (N_19709,N_18710,N_18679);
nor U19710 (N_19710,N_18582,N_18892);
nor U19711 (N_19711,N_18374,N_18296);
xnor U19712 (N_19712,N_18155,N_18243);
nor U19713 (N_19713,N_18008,N_18440);
nand U19714 (N_19714,N_18836,N_18937);
nand U19715 (N_19715,N_18367,N_18074);
xor U19716 (N_19716,N_18522,N_18820);
and U19717 (N_19717,N_18642,N_18881);
xor U19718 (N_19718,N_18048,N_18685);
xor U19719 (N_19719,N_18780,N_18514);
or U19720 (N_19720,N_18552,N_18342);
and U19721 (N_19721,N_18401,N_18166);
nand U19722 (N_19722,N_18502,N_18312);
nand U19723 (N_19723,N_18132,N_18097);
nand U19724 (N_19724,N_18288,N_18682);
and U19725 (N_19725,N_18591,N_18718);
nor U19726 (N_19726,N_18241,N_18659);
and U19727 (N_19727,N_18185,N_18218);
xnor U19728 (N_19728,N_18919,N_18743);
or U19729 (N_19729,N_18253,N_18769);
nand U19730 (N_19730,N_18636,N_18405);
xor U19731 (N_19731,N_18647,N_18546);
and U19732 (N_19732,N_18796,N_18771);
and U19733 (N_19733,N_18181,N_18325);
nor U19734 (N_19734,N_18299,N_18173);
xor U19735 (N_19735,N_18694,N_18636);
nand U19736 (N_19736,N_18973,N_18414);
and U19737 (N_19737,N_18686,N_18103);
nor U19738 (N_19738,N_18192,N_18962);
xnor U19739 (N_19739,N_18366,N_18405);
or U19740 (N_19740,N_18714,N_18304);
and U19741 (N_19741,N_18121,N_18944);
nand U19742 (N_19742,N_18609,N_18196);
or U19743 (N_19743,N_18639,N_18444);
or U19744 (N_19744,N_18872,N_18772);
and U19745 (N_19745,N_18088,N_18766);
nor U19746 (N_19746,N_18651,N_18750);
nand U19747 (N_19747,N_18656,N_18287);
and U19748 (N_19748,N_18368,N_18876);
nand U19749 (N_19749,N_18866,N_18195);
nand U19750 (N_19750,N_18171,N_18203);
and U19751 (N_19751,N_18216,N_18654);
and U19752 (N_19752,N_18876,N_18352);
xor U19753 (N_19753,N_18080,N_18975);
nor U19754 (N_19754,N_18566,N_18386);
or U19755 (N_19755,N_18452,N_18126);
nand U19756 (N_19756,N_18513,N_18667);
nand U19757 (N_19757,N_18912,N_18940);
nor U19758 (N_19758,N_18087,N_18126);
or U19759 (N_19759,N_18732,N_18569);
or U19760 (N_19760,N_18057,N_18239);
nand U19761 (N_19761,N_18733,N_18473);
or U19762 (N_19762,N_18029,N_18820);
xor U19763 (N_19763,N_18784,N_18468);
and U19764 (N_19764,N_18484,N_18897);
and U19765 (N_19765,N_18697,N_18549);
nor U19766 (N_19766,N_18198,N_18339);
and U19767 (N_19767,N_18029,N_18699);
xor U19768 (N_19768,N_18170,N_18219);
and U19769 (N_19769,N_18127,N_18411);
nor U19770 (N_19770,N_18657,N_18985);
or U19771 (N_19771,N_18194,N_18038);
xnor U19772 (N_19772,N_18782,N_18847);
and U19773 (N_19773,N_18316,N_18826);
nand U19774 (N_19774,N_18760,N_18708);
and U19775 (N_19775,N_18971,N_18177);
and U19776 (N_19776,N_18698,N_18837);
xnor U19777 (N_19777,N_18323,N_18419);
and U19778 (N_19778,N_18894,N_18836);
nor U19779 (N_19779,N_18678,N_18377);
nor U19780 (N_19780,N_18152,N_18783);
nand U19781 (N_19781,N_18038,N_18628);
nor U19782 (N_19782,N_18347,N_18853);
or U19783 (N_19783,N_18992,N_18063);
xor U19784 (N_19784,N_18859,N_18032);
and U19785 (N_19785,N_18673,N_18092);
xor U19786 (N_19786,N_18306,N_18345);
nand U19787 (N_19787,N_18707,N_18660);
nand U19788 (N_19788,N_18703,N_18997);
and U19789 (N_19789,N_18136,N_18820);
or U19790 (N_19790,N_18923,N_18275);
or U19791 (N_19791,N_18827,N_18359);
nor U19792 (N_19792,N_18072,N_18300);
and U19793 (N_19793,N_18452,N_18167);
and U19794 (N_19794,N_18132,N_18017);
or U19795 (N_19795,N_18167,N_18675);
nor U19796 (N_19796,N_18561,N_18446);
or U19797 (N_19797,N_18558,N_18058);
nand U19798 (N_19798,N_18748,N_18541);
or U19799 (N_19799,N_18149,N_18902);
and U19800 (N_19800,N_18043,N_18836);
xnor U19801 (N_19801,N_18225,N_18342);
nor U19802 (N_19802,N_18829,N_18251);
nand U19803 (N_19803,N_18038,N_18570);
nand U19804 (N_19804,N_18599,N_18441);
and U19805 (N_19805,N_18075,N_18852);
nand U19806 (N_19806,N_18468,N_18886);
and U19807 (N_19807,N_18072,N_18638);
or U19808 (N_19808,N_18173,N_18552);
nand U19809 (N_19809,N_18400,N_18678);
or U19810 (N_19810,N_18047,N_18394);
nand U19811 (N_19811,N_18708,N_18748);
and U19812 (N_19812,N_18516,N_18192);
xor U19813 (N_19813,N_18434,N_18170);
nor U19814 (N_19814,N_18700,N_18029);
and U19815 (N_19815,N_18410,N_18011);
nor U19816 (N_19816,N_18070,N_18309);
nor U19817 (N_19817,N_18306,N_18065);
and U19818 (N_19818,N_18098,N_18505);
nand U19819 (N_19819,N_18209,N_18964);
xnor U19820 (N_19820,N_18644,N_18046);
and U19821 (N_19821,N_18870,N_18043);
xnor U19822 (N_19822,N_18240,N_18234);
xor U19823 (N_19823,N_18907,N_18691);
nor U19824 (N_19824,N_18236,N_18084);
nand U19825 (N_19825,N_18654,N_18251);
xor U19826 (N_19826,N_18902,N_18672);
nand U19827 (N_19827,N_18529,N_18583);
and U19828 (N_19828,N_18495,N_18369);
nand U19829 (N_19829,N_18629,N_18944);
or U19830 (N_19830,N_18784,N_18618);
nor U19831 (N_19831,N_18968,N_18951);
or U19832 (N_19832,N_18719,N_18322);
xor U19833 (N_19833,N_18283,N_18520);
nor U19834 (N_19834,N_18752,N_18643);
or U19835 (N_19835,N_18103,N_18375);
or U19836 (N_19836,N_18143,N_18031);
or U19837 (N_19837,N_18918,N_18921);
and U19838 (N_19838,N_18210,N_18345);
and U19839 (N_19839,N_18204,N_18917);
nor U19840 (N_19840,N_18118,N_18341);
nand U19841 (N_19841,N_18208,N_18522);
xor U19842 (N_19842,N_18709,N_18882);
nand U19843 (N_19843,N_18625,N_18361);
nor U19844 (N_19844,N_18189,N_18824);
and U19845 (N_19845,N_18799,N_18745);
and U19846 (N_19846,N_18588,N_18244);
nand U19847 (N_19847,N_18257,N_18130);
or U19848 (N_19848,N_18156,N_18715);
nor U19849 (N_19849,N_18801,N_18836);
and U19850 (N_19850,N_18267,N_18293);
nor U19851 (N_19851,N_18408,N_18121);
nand U19852 (N_19852,N_18757,N_18354);
nand U19853 (N_19853,N_18665,N_18897);
nand U19854 (N_19854,N_18325,N_18330);
nand U19855 (N_19855,N_18718,N_18609);
nor U19856 (N_19856,N_18864,N_18768);
and U19857 (N_19857,N_18668,N_18336);
nand U19858 (N_19858,N_18741,N_18577);
and U19859 (N_19859,N_18540,N_18631);
or U19860 (N_19860,N_18578,N_18588);
nand U19861 (N_19861,N_18497,N_18971);
or U19862 (N_19862,N_18760,N_18467);
xor U19863 (N_19863,N_18313,N_18190);
or U19864 (N_19864,N_18612,N_18228);
nand U19865 (N_19865,N_18705,N_18880);
nand U19866 (N_19866,N_18060,N_18422);
nand U19867 (N_19867,N_18534,N_18781);
xnor U19868 (N_19868,N_18005,N_18901);
and U19869 (N_19869,N_18207,N_18305);
nor U19870 (N_19870,N_18502,N_18103);
xor U19871 (N_19871,N_18143,N_18963);
nor U19872 (N_19872,N_18900,N_18510);
or U19873 (N_19873,N_18930,N_18746);
xor U19874 (N_19874,N_18485,N_18336);
or U19875 (N_19875,N_18668,N_18269);
and U19876 (N_19876,N_18592,N_18005);
and U19877 (N_19877,N_18477,N_18832);
nor U19878 (N_19878,N_18674,N_18946);
or U19879 (N_19879,N_18492,N_18593);
or U19880 (N_19880,N_18364,N_18342);
and U19881 (N_19881,N_18747,N_18513);
and U19882 (N_19882,N_18878,N_18485);
or U19883 (N_19883,N_18280,N_18262);
and U19884 (N_19884,N_18053,N_18827);
nor U19885 (N_19885,N_18461,N_18195);
and U19886 (N_19886,N_18146,N_18831);
nand U19887 (N_19887,N_18922,N_18466);
nand U19888 (N_19888,N_18091,N_18178);
and U19889 (N_19889,N_18720,N_18192);
and U19890 (N_19890,N_18834,N_18000);
or U19891 (N_19891,N_18301,N_18337);
xor U19892 (N_19892,N_18997,N_18717);
or U19893 (N_19893,N_18292,N_18043);
or U19894 (N_19894,N_18622,N_18758);
nand U19895 (N_19895,N_18991,N_18596);
nor U19896 (N_19896,N_18673,N_18874);
nor U19897 (N_19897,N_18356,N_18506);
xor U19898 (N_19898,N_18421,N_18416);
or U19899 (N_19899,N_18992,N_18164);
and U19900 (N_19900,N_18528,N_18364);
nor U19901 (N_19901,N_18887,N_18137);
or U19902 (N_19902,N_18412,N_18759);
or U19903 (N_19903,N_18119,N_18021);
and U19904 (N_19904,N_18546,N_18930);
nand U19905 (N_19905,N_18262,N_18980);
nor U19906 (N_19906,N_18375,N_18011);
xor U19907 (N_19907,N_18669,N_18916);
or U19908 (N_19908,N_18778,N_18876);
nand U19909 (N_19909,N_18572,N_18249);
nand U19910 (N_19910,N_18645,N_18971);
nand U19911 (N_19911,N_18666,N_18669);
nor U19912 (N_19912,N_18070,N_18567);
or U19913 (N_19913,N_18500,N_18564);
nor U19914 (N_19914,N_18276,N_18827);
or U19915 (N_19915,N_18979,N_18193);
and U19916 (N_19916,N_18064,N_18352);
or U19917 (N_19917,N_18257,N_18479);
or U19918 (N_19918,N_18964,N_18672);
xor U19919 (N_19919,N_18308,N_18928);
xor U19920 (N_19920,N_18877,N_18208);
xor U19921 (N_19921,N_18889,N_18792);
nor U19922 (N_19922,N_18622,N_18990);
xor U19923 (N_19923,N_18674,N_18004);
xor U19924 (N_19924,N_18350,N_18459);
and U19925 (N_19925,N_18048,N_18975);
or U19926 (N_19926,N_18349,N_18774);
nand U19927 (N_19927,N_18534,N_18962);
and U19928 (N_19928,N_18548,N_18075);
nand U19929 (N_19929,N_18017,N_18410);
nand U19930 (N_19930,N_18387,N_18682);
and U19931 (N_19931,N_18109,N_18754);
nor U19932 (N_19932,N_18450,N_18806);
nand U19933 (N_19933,N_18116,N_18237);
xor U19934 (N_19934,N_18540,N_18981);
and U19935 (N_19935,N_18822,N_18222);
and U19936 (N_19936,N_18879,N_18608);
nand U19937 (N_19937,N_18850,N_18090);
or U19938 (N_19938,N_18397,N_18489);
nand U19939 (N_19939,N_18755,N_18200);
and U19940 (N_19940,N_18182,N_18438);
and U19941 (N_19941,N_18111,N_18365);
xor U19942 (N_19942,N_18085,N_18087);
xnor U19943 (N_19943,N_18948,N_18108);
and U19944 (N_19944,N_18367,N_18500);
nor U19945 (N_19945,N_18567,N_18099);
and U19946 (N_19946,N_18004,N_18545);
or U19947 (N_19947,N_18820,N_18437);
nor U19948 (N_19948,N_18465,N_18058);
nand U19949 (N_19949,N_18540,N_18848);
xnor U19950 (N_19950,N_18182,N_18391);
or U19951 (N_19951,N_18372,N_18680);
nor U19952 (N_19952,N_18908,N_18699);
and U19953 (N_19953,N_18999,N_18190);
and U19954 (N_19954,N_18885,N_18264);
and U19955 (N_19955,N_18609,N_18394);
nand U19956 (N_19956,N_18009,N_18982);
nand U19957 (N_19957,N_18575,N_18713);
nor U19958 (N_19958,N_18316,N_18913);
and U19959 (N_19959,N_18976,N_18910);
xnor U19960 (N_19960,N_18202,N_18267);
and U19961 (N_19961,N_18192,N_18361);
and U19962 (N_19962,N_18936,N_18194);
nor U19963 (N_19963,N_18207,N_18001);
xor U19964 (N_19964,N_18347,N_18503);
or U19965 (N_19965,N_18227,N_18723);
nand U19966 (N_19966,N_18185,N_18362);
or U19967 (N_19967,N_18946,N_18187);
or U19968 (N_19968,N_18890,N_18025);
xor U19969 (N_19969,N_18803,N_18286);
nand U19970 (N_19970,N_18061,N_18708);
xor U19971 (N_19971,N_18010,N_18762);
nand U19972 (N_19972,N_18178,N_18470);
nand U19973 (N_19973,N_18426,N_18352);
nand U19974 (N_19974,N_18472,N_18575);
nor U19975 (N_19975,N_18981,N_18077);
nand U19976 (N_19976,N_18292,N_18949);
and U19977 (N_19977,N_18035,N_18250);
or U19978 (N_19978,N_18225,N_18604);
and U19979 (N_19979,N_18228,N_18418);
nor U19980 (N_19980,N_18629,N_18929);
or U19981 (N_19981,N_18128,N_18733);
xor U19982 (N_19982,N_18313,N_18845);
or U19983 (N_19983,N_18437,N_18725);
or U19984 (N_19984,N_18492,N_18392);
xnor U19985 (N_19985,N_18216,N_18078);
and U19986 (N_19986,N_18015,N_18031);
and U19987 (N_19987,N_18659,N_18381);
or U19988 (N_19988,N_18655,N_18327);
xnor U19989 (N_19989,N_18007,N_18460);
nand U19990 (N_19990,N_18476,N_18532);
xor U19991 (N_19991,N_18020,N_18617);
and U19992 (N_19992,N_18780,N_18641);
and U19993 (N_19993,N_18995,N_18288);
nor U19994 (N_19994,N_18442,N_18196);
and U19995 (N_19995,N_18250,N_18033);
and U19996 (N_19996,N_18013,N_18680);
nand U19997 (N_19997,N_18755,N_18618);
nor U19998 (N_19998,N_18357,N_18856);
xor U19999 (N_19999,N_18323,N_18608);
nor U20000 (N_20000,N_19601,N_19513);
xor U20001 (N_20001,N_19799,N_19112);
xor U20002 (N_20002,N_19005,N_19454);
nor U20003 (N_20003,N_19812,N_19290);
and U20004 (N_20004,N_19358,N_19853);
and U20005 (N_20005,N_19985,N_19524);
nand U20006 (N_20006,N_19203,N_19456);
and U20007 (N_20007,N_19934,N_19779);
and U20008 (N_20008,N_19202,N_19592);
or U20009 (N_20009,N_19109,N_19478);
nor U20010 (N_20010,N_19229,N_19700);
nor U20011 (N_20011,N_19880,N_19230);
and U20012 (N_20012,N_19283,N_19564);
nand U20013 (N_20013,N_19424,N_19219);
and U20014 (N_20014,N_19741,N_19458);
nand U20015 (N_20015,N_19938,N_19284);
nor U20016 (N_20016,N_19863,N_19923);
nor U20017 (N_20017,N_19655,N_19113);
xor U20018 (N_20018,N_19683,N_19279);
and U20019 (N_20019,N_19169,N_19854);
or U20020 (N_20020,N_19871,N_19015);
xor U20021 (N_20021,N_19050,N_19468);
nor U20022 (N_20022,N_19434,N_19342);
nand U20023 (N_20023,N_19533,N_19632);
or U20024 (N_20024,N_19891,N_19767);
nor U20025 (N_20025,N_19716,N_19411);
or U20026 (N_20026,N_19792,N_19545);
and U20027 (N_20027,N_19364,N_19544);
nor U20028 (N_20028,N_19857,N_19758);
nor U20029 (N_20029,N_19471,N_19894);
nor U20030 (N_20030,N_19173,N_19412);
or U20031 (N_20031,N_19692,N_19377);
nor U20032 (N_20032,N_19776,N_19625);
xor U20033 (N_20033,N_19817,N_19013);
xor U20034 (N_20034,N_19235,N_19046);
nor U20035 (N_20035,N_19795,N_19944);
nand U20036 (N_20036,N_19790,N_19073);
xor U20037 (N_20037,N_19239,N_19218);
and U20038 (N_20038,N_19577,N_19380);
and U20039 (N_20039,N_19905,N_19849);
xor U20040 (N_20040,N_19461,N_19660);
and U20041 (N_20041,N_19262,N_19766);
or U20042 (N_20042,N_19640,N_19269);
nand U20043 (N_20043,N_19039,N_19157);
or U20044 (N_20044,N_19608,N_19910);
nand U20045 (N_20045,N_19907,N_19929);
xnor U20046 (N_20046,N_19549,N_19963);
nor U20047 (N_20047,N_19858,N_19600);
xor U20048 (N_20048,N_19504,N_19052);
and U20049 (N_20049,N_19878,N_19062);
nand U20050 (N_20050,N_19546,N_19210);
or U20051 (N_20051,N_19840,N_19518);
xor U20052 (N_20052,N_19286,N_19401);
nand U20053 (N_20053,N_19724,N_19915);
and U20054 (N_20054,N_19253,N_19676);
nor U20055 (N_20055,N_19069,N_19125);
or U20056 (N_20056,N_19637,N_19502);
nand U20057 (N_20057,N_19605,N_19071);
and U20058 (N_20058,N_19704,N_19460);
nor U20059 (N_20059,N_19523,N_19025);
nand U20060 (N_20060,N_19444,N_19550);
xor U20061 (N_20061,N_19280,N_19031);
or U20062 (N_20062,N_19254,N_19883);
xnor U20063 (N_20063,N_19673,N_19623);
xor U20064 (N_20064,N_19594,N_19833);
and U20065 (N_20065,N_19749,N_19886);
or U20066 (N_20066,N_19788,N_19495);
nand U20067 (N_20067,N_19075,N_19383);
xor U20068 (N_20068,N_19086,N_19787);
nand U20069 (N_20069,N_19011,N_19087);
nand U20070 (N_20070,N_19249,N_19463);
nand U20071 (N_20071,N_19998,N_19535);
nor U20072 (N_20072,N_19597,N_19036);
and U20073 (N_20073,N_19647,N_19346);
nor U20074 (N_20074,N_19861,N_19408);
and U20075 (N_20075,N_19671,N_19498);
and U20076 (N_20076,N_19029,N_19962);
or U20077 (N_20077,N_19128,N_19908);
nor U20078 (N_20078,N_19020,N_19882);
nand U20079 (N_20079,N_19237,N_19761);
xnor U20080 (N_20080,N_19099,N_19734);
xor U20081 (N_20081,N_19226,N_19658);
or U20082 (N_20082,N_19540,N_19974);
and U20083 (N_20083,N_19356,N_19559);
or U20084 (N_20084,N_19924,N_19483);
and U20085 (N_20085,N_19551,N_19063);
or U20086 (N_20086,N_19497,N_19017);
xor U20087 (N_20087,N_19139,N_19289);
and U20088 (N_20088,N_19914,N_19407);
nand U20089 (N_20089,N_19402,N_19182);
or U20090 (N_20090,N_19171,N_19681);
xor U20091 (N_20091,N_19611,N_19663);
xor U20092 (N_20092,N_19141,N_19181);
nand U20093 (N_20093,N_19437,N_19469);
nor U20094 (N_20094,N_19827,N_19371);
and U20095 (N_20095,N_19696,N_19057);
and U20096 (N_20096,N_19599,N_19541);
xnor U20097 (N_20097,N_19505,N_19775);
nor U20098 (N_20098,N_19869,N_19068);
nor U20099 (N_20099,N_19091,N_19324);
xnor U20100 (N_20100,N_19939,N_19482);
or U20101 (N_20101,N_19720,N_19292);
or U20102 (N_20102,N_19521,N_19893);
and U20103 (N_20103,N_19548,N_19555);
xnor U20104 (N_20104,N_19098,N_19170);
and U20105 (N_20105,N_19032,N_19145);
and U20106 (N_20106,N_19064,N_19830);
and U20107 (N_20107,N_19679,N_19423);
nor U20108 (N_20108,N_19193,N_19206);
or U20109 (N_20109,N_19819,N_19890);
nand U20110 (N_20110,N_19185,N_19189);
or U20111 (N_20111,N_19656,N_19430);
nor U20112 (N_20112,N_19682,N_19848);
nor U20113 (N_20113,N_19163,N_19560);
and U20114 (N_20114,N_19887,N_19217);
nand U20115 (N_20115,N_19976,N_19097);
nand U20116 (N_20116,N_19723,N_19855);
nand U20117 (N_20117,N_19657,N_19059);
nor U20118 (N_20118,N_19028,N_19874);
nand U20119 (N_20119,N_19773,N_19768);
nand U20120 (N_20120,N_19680,N_19705);
nor U20121 (N_20121,N_19487,N_19100);
nor U20122 (N_20122,N_19166,N_19715);
or U20123 (N_20123,N_19007,N_19903);
and U20124 (N_20124,N_19542,N_19379);
nor U20125 (N_20125,N_19580,N_19372);
or U20126 (N_20126,N_19575,N_19699);
nor U20127 (N_20127,N_19539,N_19065);
nor U20128 (N_20128,N_19480,N_19162);
or U20129 (N_20129,N_19928,N_19950);
or U20130 (N_20130,N_19376,N_19278);
and U20131 (N_20131,N_19511,N_19186);
and U20132 (N_20132,N_19328,N_19096);
nor U20133 (N_20133,N_19791,N_19631);
xnor U20134 (N_20134,N_19584,N_19969);
or U20135 (N_20135,N_19026,N_19866);
xnor U20136 (N_20136,N_19164,N_19260);
xor U20137 (N_20137,N_19670,N_19778);
and U20138 (N_20138,N_19876,N_19117);
nand U20139 (N_20139,N_19510,N_19582);
or U20140 (N_20140,N_19574,N_19838);
nand U20141 (N_20141,N_19429,N_19390);
nand U20142 (N_20142,N_19256,N_19174);
nand U20143 (N_20143,N_19968,N_19116);
or U20144 (N_20144,N_19947,N_19579);
xor U20145 (N_20145,N_19941,N_19636);
xnor U20146 (N_20146,N_19814,N_19628);
and U20147 (N_20147,N_19588,N_19509);
xnor U20148 (N_20148,N_19561,N_19225);
nand U20149 (N_20149,N_19426,N_19231);
nor U20150 (N_20150,N_19208,N_19406);
and U20151 (N_20151,N_19554,N_19875);
xor U20152 (N_20152,N_19400,N_19422);
nor U20153 (N_20153,N_19095,N_19645);
and U20154 (N_20154,N_19688,N_19476);
nor U20155 (N_20155,N_19034,N_19490);
and U20156 (N_20156,N_19906,N_19785);
xor U20157 (N_20157,N_19023,N_19133);
or U20158 (N_20158,N_19828,N_19911);
nand U20159 (N_20159,N_19439,N_19273);
xor U20160 (N_20160,N_19136,N_19078);
nor U20161 (N_20161,N_19957,N_19357);
xor U20162 (N_20162,N_19194,N_19008);
and U20163 (N_20163,N_19107,N_19144);
xnor U20164 (N_20164,N_19512,N_19578);
nand U20165 (N_20165,N_19634,N_19122);
or U20166 (N_20166,N_19234,N_19367);
xnor U20167 (N_20167,N_19826,N_19298);
and U20168 (N_20168,N_19972,N_19641);
or U20169 (N_20169,N_19806,N_19261);
or U20170 (N_20170,N_19306,N_19151);
nand U20171 (N_20171,N_19121,N_19051);
xnor U20172 (N_20172,N_19088,N_19014);
and U20173 (N_20173,N_19281,N_19248);
nor U20174 (N_20174,N_19000,N_19251);
xnor U20175 (N_20175,N_19530,N_19686);
or U20176 (N_20176,N_19913,N_19102);
and U20177 (N_20177,N_19649,N_19813);
nand U20178 (N_20178,N_19425,N_19103);
and U20179 (N_20179,N_19115,N_19465);
nor U20180 (N_20180,N_19755,N_19847);
or U20181 (N_20181,N_19956,N_19843);
nand U20182 (N_20182,N_19297,N_19945);
and U20183 (N_20183,N_19275,N_19810);
or U20184 (N_20184,N_19515,N_19703);
nand U20185 (N_20185,N_19764,N_19763);
nor U20186 (N_20186,N_19846,N_19149);
xor U20187 (N_20187,N_19481,N_19881);
nor U20188 (N_20188,N_19732,N_19313);
nor U20189 (N_20189,N_19593,N_19517);
nand U20190 (N_20190,N_19360,N_19370);
nor U20191 (N_20191,N_19900,N_19147);
xnor U20192 (N_20192,N_19291,N_19931);
and U20193 (N_20193,N_19339,N_19082);
nand U20194 (N_20194,N_19074,N_19322);
nand U20195 (N_20195,N_19021,N_19815);
nor U20196 (N_20196,N_19693,N_19227);
nor U20197 (N_20197,N_19006,N_19421);
and U20198 (N_20198,N_19943,N_19450);
xor U20199 (N_20199,N_19296,N_19252);
nor U20200 (N_20200,N_19433,N_19503);
or U20201 (N_20201,N_19001,N_19922);
or U20202 (N_20202,N_19624,N_19304);
nor U20203 (N_20203,N_19332,N_19965);
nand U20204 (N_20204,N_19405,N_19056);
and U20205 (N_20205,N_19606,N_19754);
xor U20206 (N_20206,N_19629,N_19678);
nor U20207 (N_20207,N_19753,N_19085);
or U20208 (N_20208,N_19108,N_19730);
nor U20209 (N_20209,N_19491,N_19733);
xor U20210 (N_20210,N_19603,N_19177);
nor U20211 (N_20211,N_19654,N_19436);
and U20212 (N_20212,N_19111,N_19355);
and U20213 (N_20213,N_19816,N_19659);
nor U20214 (N_20214,N_19083,N_19207);
nor U20215 (N_20215,N_19146,N_19867);
nand U20216 (N_20216,N_19630,N_19820);
xor U20217 (N_20217,N_19961,N_19650);
or U20218 (N_20218,N_19419,N_19970);
or U20219 (N_20219,N_19804,N_19598);
or U20220 (N_20220,N_19996,N_19374);
xor U20221 (N_20221,N_19479,N_19079);
and U20222 (N_20222,N_19178,N_19397);
nand U20223 (N_20223,N_19821,N_19836);
xnor U20224 (N_20224,N_19167,N_19721);
nor U20225 (N_20225,N_19457,N_19952);
nand U20226 (N_20226,N_19942,N_19084);
nand U20227 (N_20227,N_19842,N_19038);
and U20228 (N_20228,N_19438,N_19901);
or U20229 (N_20229,N_19839,N_19484);
xnor U20230 (N_20230,N_19211,N_19349);
and U20231 (N_20231,N_19997,N_19470);
xor U20232 (N_20232,N_19199,N_19935);
and U20233 (N_20233,N_19135,N_19807);
xor U20234 (N_20234,N_19667,N_19975);
xnor U20235 (N_20235,N_19652,N_19209);
nand U20236 (N_20236,N_19049,N_19707);
and U20237 (N_20237,N_19414,N_19003);
or U20238 (N_20238,N_19740,N_19337);
and U20239 (N_20239,N_19933,N_19148);
nand U20240 (N_20240,N_19009,N_19562);
nor U20241 (N_20241,N_19916,N_19191);
xor U20242 (N_20242,N_19571,N_19310);
nand U20243 (N_20243,N_19953,N_19303);
and U20244 (N_20244,N_19951,N_19824);
and U20245 (N_20245,N_19832,N_19299);
or U20246 (N_20246,N_19392,N_19973);
or U20247 (N_20247,N_19977,N_19727);
nand U20248 (N_20248,N_19309,N_19835);
or U20249 (N_20249,N_19536,N_19581);
nand U20250 (N_20250,N_19466,N_19662);
and U20251 (N_20251,N_19926,N_19485);
xor U20252 (N_20252,N_19010,N_19442);
xor U20253 (N_20253,N_19311,N_19756);
nor U20254 (N_20254,N_19745,N_19750);
nand U20255 (N_20255,N_19308,N_19198);
or U20256 (N_20256,N_19354,N_19570);
nand U20257 (N_20257,N_19123,N_19999);
or U20258 (N_20258,N_19982,N_19118);
nand U20259 (N_20259,N_19736,N_19387);
nor U20260 (N_20260,N_19132,N_19222);
xor U20261 (N_20261,N_19477,N_19796);
nand U20262 (N_20262,N_19259,N_19447);
nor U20263 (N_20263,N_19563,N_19818);
or U20264 (N_20264,N_19987,N_19738);
and U20265 (N_20265,N_19589,N_19060);
nand U20266 (N_20266,N_19531,N_19687);
and U20267 (N_20267,N_19072,N_19712);
xor U20268 (N_20268,N_19889,N_19615);
or U20269 (N_20269,N_19002,N_19898);
or U20270 (N_20270,N_19917,N_19413);
or U20271 (N_20271,N_19092,N_19389);
nand U20272 (N_20272,N_19844,N_19537);
and U20273 (N_20273,N_19892,N_19744);
or U20274 (N_20274,N_19246,N_19752);
nor U20275 (N_20275,N_19197,N_19446);
nand U20276 (N_20276,N_19475,N_19435);
nand U20277 (N_20277,N_19345,N_19054);
nor U20278 (N_20278,N_19534,N_19702);
nor U20279 (N_20279,N_19607,N_19547);
xor U20280 (N_20280,N_19742,N_19675);
or U20281 (N_20281,N_19264,N_19618);
nor U20282 (N_20282,N_19927,N_19646);
nor U20283 (N_20283,N_19896,N_19385);
nand U20284 (N_20284,N_19321,N_19948);
or U20285 (N_20285,N_19809,N_19301);
and U20286 (N_20286,N_19488,N_19363);
nand U20287 (N_20287,N_19041,N_19232);
xnor U20288 (N_20288,N_19642,N_19610);
xnor U20289 (N_20289,N_19201,N_19271);
xnor U20290 (N_20290,N_19090,N_19165);
or U20291 (N_20291,N_19786,N_19940);
nor U20292 (N_20292,N_19319,N_19860);
and U20293 (N_20293,N_19340,N_19529);
and U20294 (N_20294,N_19765,N_19126);
or U20295 (N_20295,N_19443,N_19305);
nand U20296 (N_20296,N_19771,N_19638);
or U20297 (N_20297,N_19070,N_19983);
xnor U20298 (N_20298,N_19316,N_19845);
nor U20299 (N_20299,N_19930,N_19288);
nand U20300 (N_20300,N_19677,N_19669);
nand U20301 (N_20301,N_19445,N_19396);
nand U20302 (N_20302,N_19022,N_19859);
and U20303 (N_20303,N_19873,N_19595);
nor U20304 (N_20304,N_19293,N_19462);
xor U20305 (N_20305,N_19250,N_19247);
and U20306 (N_20306,N_19501,N_19295);
xor U20307 (N_20307,N_19417,N_19780);
and U20308 (N_20308,N_19770,N_19955);
nor U20309 (N_20309,N_19241,N_19381);
and U20310 (N_20310,N_19464,N_19258);
or U20311 (N_20311,N_19472,N_19048);
nand U20312 (N_20312,N_19664,N_19781);
xnor U20313 (N_20313,N_19691,N_19872);
and U20314 (N_20314,N_19336,N_19195);
xnor U20315 (N_20315,N_19369,N_19661);
or U20316 (N_20316,N_19365,N_19190);
xor U20317 (N_20317,N_19255,N_19666);
nor U20318 (N_20318,N_19850,N_19613);
and U20319 (N_20319,N_19760,N_19089);
nand U20320 (N_20320,N_19585,N_19762);
xor U20321 (N_20321,N_19586,N_19236);
nand U20322 (N_20322,N_19500,N_19263);
nor U20323 (N_20323,N_19382,N_19192);
nand U20324 (N_20324,N_19981,N_19532);
or U20325 (N_20325,N_19708,N_19728);
and U20326 (N_20326,N_19053,N_19617);
and U20327 (N_20327,N_19267,N_19522);
nand U20328 (N_20328,N_19223,N_19757);
or U20329 (N_20329,N_19877,N_19183);
nand U20330 (N_20330,N_19351,N_19706);
or U20331 (N_20331,N_19127,N_19499);
nand U20332 (N_20332,N_19879,N_19731);
nand U20333 (N_20333,N_19489,N_19777);
nand U20334 (N_20334,N_19769,N_19949);
nand U20335 (N_20335,N_19743,N_19416);
and U20336 (N_20336,N_19175,N_19045);
or U20337 (N_20337,N_19394,N_19904);
xnor U20338 (N_20338,N_19044,N_19384);
nor U20339 (N_20339,N_19287,N_19837);
or U20340 (N_20340,N_19018,N_19988);
nand U20341 (N_20341,N_19130,N_19449);
or U20342 (N_20342,N_19516,N_19591);
xor U20343 (N_20343,N_19432,N_19156);
or U20344 (N_20344,N_19320,N_19698);
xnor U20345 (N_20345,N_19954,N_19386);
and U20346 (N_20346,N_19272,N_19153);
or U20347 (N_20347,N_19711,N_19066);
or U20348 (N_20348,N_19134,N_19040);
nand U20349 (N_20349,N_19994,N_19378);
or U20350 (N_20350,N_19282,N_19158);
nor U20351 (N_20351,N_19895,N_19722);
xor U20352 (N_20352,N_19058,N_19967);
or U20353 (N_20353,N_19569,N_19155);
xor U20354 (N_20354,N_19868,N_19725);
and U20355 (N_20355,N_19341,N_19366);
nand U20356 (N_20356,N_19690,N_19841);
xnor U20357 (N_20357,N_19037,N_19635);
or U20358 (N_20358,N_19388,N_19672);
nor U20359 (N_20359,N_19718,N_19215);
xnor U20360 (N_20360,N_19568,N_19979);
xnor U20361 (N_20361,N_19798,N_19142);
nand U20362 (N_20362,N_19077,N_19918);
nand U20363 (N_20363,N_19614,N_19343);
or U20364 (N_20364,N_19205,N_19782);
xor U20365 (N_20365,N_19409,N_19214);
nand U20366 (N_20366,N_19418,N_19265);
nor U20367 (N_20367,N_19325,N_19831);
xnor U20368 (N_20368,N_19101,N_19245);
or U20369 (N_20369,N_19919,N_19984);
and U20370 (N_20370,N_19076,N_19990);
and U20371 (N_20371,N_19131,N_19302);
and U20372 (N_20372,N_19238,N_19344);
nor U20373 (N_20373,N_19800,N_19124);
or U20374 (N_20374,N_19888,N_19701);
or U20375 (N_20375,N_19243,N_19159);
nor U20376 (N_20376,N_19622,N_19335);
nor U20377 (N_20377,N_19627,N_19932);
or U20378 (N_20378,N_19300,N_19644);
or U20379 (N_20379,N_19016,N_19525);
nand U20380 (N_20380,N_19811,N_19403);
xor U20381 (N_20381,N_19616,N_19710);
nand U20382 (N_20382,N_19119,N_19395);
and U20383 (N_20383,N_19494,N_19473);
xor U20384 (N_20384,N_19274,N_19719);
nor U20385 (N_20385,N_19043,N_19067);
nor U20386 (N_20386,N_19240,N_19359);
nand U20387 (N_20387,N_19991,N_19323);
or U20388 (N_20388,N_19404,N_19620);
or U20389 (N_20389,N_19747,N_19114);
nor U20390 (N_20390,N_19714,N_19596);
nor U20391 (N_20391,N_19684,N_19244);
xnor U20392 (N_20392,N_19391,N_19989);
nand U20393 (N_20393,N_19829,N_19856);
and U20394 (N_20394,N_19958,N_19851);
and U20395 (N_20395,N_19285,N_19399);
nand U20396 (N_20396,N_19138,N_19459);
or U20397 (N_20397,N_19980,N_19228);
nor U20398 (N_20398,N_19150,N_19307);
or U20399 (N_20399,N_19154,N_19451);
or U20400 (N_20400,N_19694,N_19587);
xor U20401 (N_20401,N_19266,N_19626);
nand U20402 (N_20402,N_19528,N_19960);
xor U20403 (N_20403,N_19648,N_19793);
and U20404 (N_20404,N_19937,N_19216);
and U20405 (N_20405,N_19713,N_19590);
and U20406 (N_20406,N_19493,N_19350);
or U20407 (N_20407,N_19748,N_19474);
and U20408 (N_20408,N_19353,N_19739);
or U20409 (N_20409,N_19294,N_19326);
nor U20410 (N_20410,N_19276,N_19453);
or U20411 (N_20411,N_19452,N_19496);
and U20412 (N_20412,N_19759,N_19803);
nor U20413 (N_20413,N_19019,N_19899);
or U20414 (N_20414,N_19986,N_19188);
nor U20415 (N_20415,N_19268,N_19212);
or U20416 (N_20416,N_19794,N_19612);
nor U20417 (N_20417,N_19737,N_19331);
nand U20418 (N_20418,N_19870,N_19187);
or U20419 (N_20419,N_19772,N_19129);
xor U20420 (N_20420,N_19427,N_19080);
nor U20421 (N_20421,N_19602,N_19527);
nor U20422 (N_20422,N_19104,N_19746);
xnor U20423 (N_20423,N_19609,N_19106);
xor U20424 (N_20424,N_19318,N_19959);
nor U20425 (N_20425,N_19315,N_19520);
and U20426 (N_20426,N_19514,N_19012);
or U20427 (N_20427,N_19553,N_19619);
or U20428 (N_20428,N_19347,N_19909);
or U20429 (N_20429,N_19964,N_19257);
or U20430 (N_20430,N_19808,N_19506);
nor U20431 (N_20431,N_19140,N_19033);
nand U20432 (N_20432,N_19338,N_19823);
nor U20433 (N_20433,N_19196,N_19558);
nor U20434 (N_20434,N_19172,N_19361);
nor U20435 (N_20435,N_19334,N_19885);
nand U20436 (N_20436,N_19971,N_19572);
nor U20437 (N_20437,N_19176,N_19978);
nor U20438 (N_20438,N_19042,N_19348);
nor U20439 (N_20439,N_19946,N_19161);
nand U20440 (N_20440,N_19695,N_19362);
and U20441 (N_20441,N_19966,N_19864);
nor U20442 (N_20442,N_19801,N_19204);
nand U20443 (N_20443,N_19774,N_19352);
and U20444 (N_20444,N_19884,N_19526);
and U20445 (N_20445,N_19576,N_19538);
nand U20446 (N_20446,N_19508,N_19507);
nand U20447 (N_20447,N_19330,N_19467);
and U20448 (N_20448,N_19789,N_19852);
or U20449 (N_20449,N_19160,N_19519);
xnor U20450 (N_20450,N_19420,N_19668);
xor U20451 (N_20451,N_19865,N_19784);
xor U20452 (N_20452,N_19055,N_19329);
nor U20453 (N_20453,N_19665,N_19375);
and U20454 (N_20454,N_19825,N_19120);
xor U20455 (N_20455,N_19674,N_19902);
xnor U20456 (N_20456,N_19735,N_19543);
xor U20457 (N_20457,N_19729,N_19566);
or U20458 (N_20458,N_19897,N_19992);
and U20459 (N_20459,N_19428,N_19834);
and U20460 (N_20460,N_19557,N_19047);
xnor U20461 (N_20461,N_19448,N_19393);
nor U20462 (N_20462,N_19726,N_19035);
xnor U20463 (N_20463,N_19552,N_19685);
nor U20464 (N_20464,N_19486,N_19621);
and U20465 (N_20465,N_19105,N_19925);
xor U20466 (N_20466,N_19565,N_19368);
nor U20467 (N_20467,N_19143,N_19822);
nor U20468 (N_20468,N_19709,N_19317);
or U20469 (N_20469,N_19921,N_19314);
nor U20470 (N_20470,N_19220,N_19277);
and U20471 (N_20471,N_19213,N_19912);
and U20472 (N_20472,N_19697,N_19556);
xnor U20473 (N_20473,N_19152,N_19567);
nor U20474 (N_20474,N_19200,N_19440);
nor U20475 (N_20475,N_19180,N_19327);
and U20476 (N_20476,N_19604,N_19441);
or U20477 (N_20477,N_19936,N_19633);
and U20478 (N_20478,N_19030,N_19862);
nor U20479 (N_20479,N_19233,N_19653);
xor U20480 (N_20480,N_19179,N_19224);
nor U20481 (N_20481,N_19333,N_19168);
or U20482 (N_20482,N_19027,N_19312);
nand U20483 (N_20483,N_19573,N_19583);
or U20484 (N_20484,N_19993,N_19797);
or U20485 (N_20485,N_19995,N_19270);
nor U20486 (N_20486,N_19717,N_19093);
and U20487 (N_20487,N_19920,N_19802);
and U20488 (N_20488,N_19410,N_19639);
nor U20489 (N_20489,N_19110,N_19004);
or U20490 (N_20490,N_19373,N_19415);
nor U20491 (N_20491,N_19094,N_19061);
xor U20492 (N_20492,N_19751,N_19398);
xnor U20493 (N_20493,N_19242,N_19431);
or U20494 (N_20494,N_19024,N_19184);
nor U20495 (N_20495,N_19805,N_19081);
xnor U20496 (N_20496,N_19221,N_19783);
and U20497 (N_20497,N_19689,N_19492);
nor U20498 (N_20498,N_19455,N_19643);
or U20499 (N_20499,N_19651,N_19137);
or U20500 (N_20500,N_19884,N_19115);
xor U20501 (N_20501,N_19249,N_19250);
nor U20502 (N_20502,N_19552,N_19669);
or U20503 (N_20503,N_19499,N_19092);
nand U20504 (N_20504,N_19613,N_19434);
nand U20505 (N_20505,N_19779,N_19772);
xor U20506 (N_20506,N_19126,N_19419);
or U20507 (N_20507,N_19639,N_19102);
xnor U20508 (N_20508,N_19266,N_19592);
or U20509 (N_20509,N_19554,N_19116);
and U20510 (N_20510,N_19667,N_19537);
and U20511 (N_20511,N_19022,N_19290);
and U20512 (N_20512,N_19663,N_19720);
nand U20513 (N_20513,N_19051,N_19507);
and U20514 (N_20514,N_19340,N_19692);
xnor U20515 (N_20515,N_19120,N_19491);
nand U20516 (N_20516,N_19673,N_19825);
or U20517 (N_20517,N_19965,N_19038);
or U20518 (N_20518,N_19535,N_19464);
nand U20519 (N_20519,N_19630,N_19968);
or U20520 (N_20520,N_19574,N_19554);
or U20521 (N_20521,N_19006,N_19729);
and U20522 (N_20522,N_19648,N_19267);
nor U20523 (N_20523,N_19931,N_19574);
and U20524 (N_20524,N_19748,N_19112);
nor U20525 (N_20525,N_19570,N_19045);
and U20526 (N_20526,N_19698,N_19351);
nand U20527 (N_20527,N_19443,N_19666);
or U20528 (N_20528,N_19765,N_19441);
nand U20529 (N_20529,N_19366,N_19158);
nor U20530 (N_20530,N_19471,N_19278);
xnor U20531 (N_20531,N_19231,N_19680);
nor U20532 (N_20532,N_19318,N_19118);
and U20533 (N_20533,N_19437,N_19845);
and U20534 (N_20534,N_19784,N_19417);
and U20535 (N_20535,N_19266,N_19871);
or U20536 (N_20536,N_19559,N_19589);
xnor U20537 (N_20537,N_19668,N_19435);
or U20538 (N_20538,N_19560,N_19626);
or U20539 (N_20539,N_19779,N_19727);
nand U20540 (N_20540,N_19141,N_19057);
xor U20541 (N_20541,N_19094,N_19129);
and U20542 (N_20542,N_19885,N_19488);
nor U20543 (N_20543,N_19121,N_19894);
and U20544 (N_20544,N_19234,N_19952);
or U20545 (N_20545,N_19652,N_19097);
nand U20546 (N_20546,N_19974,N_19510);
xnor U20547 (N_20547,N_19659,N_19195);
nand U20548 (N_20548,N_19603,N_19766);
xnor U20549 (N_20549,N_19804,N_19829);
nand U20550 (N_20550,N_19117,N_19913);
xor U20551 (N_20551,N_19775,N_19250);
xnor U20552 (N_20552,N_19097,N_19267);
nand U20553 (N_20553,N_19922,N_19595);
nor U20554 (N_20554,N_19868,N_19625);
and U20555 (N_20555,N_19939,N_19181);
xor U20556 (N_20556,N_19620,N_19704);
nor U20557 (N_20557,N_19662,N_19649);
or U20558 (N_20558,N_19041,N_19450);
xnor U20559 (N_20559,N_19150,N_19011);
nand U20560 (N_20560,N_19243,N_19795);
or U20561 (N_20561,N_19650,N_19702);
xnor U20562 (N_20562,N_19209,N_19677);
nand U20563 (N_20563,N_19979,N_19282);
or U20564 (N_20564,N_19500,N_19644);
and U20565 (N_20565,N_19159,N_19759);
nand U20566 (N_20566,N_19784,N_19646);
xnor U20567 (N_20567,N_19834,N_19674);
nor U20568 (N_20568,N_19787,N_19541);
or U20569 (N_20569,N_19274,N_19526);
nand U20570 (N_20570,N_19520,N_19519);
nand U20571 (N_20571,N_19851,N_19859);
xnor U20572 (N_20572,N_19317,N_19196);
or U20573 (N_20573,N_19571,N_19862);
and U20574 (N_20574,N_19697,N_19651);
nor U20575 (N_20575,N_19547,N_19078);
nand U20576 (N_20576,N_19048,N_19541);
nand U20577 (N_20577,N_19849,N_19539);
or U20578 (N_20578,N_19991,N_19794);
and U20579 (N_20579,N_19993,N_19165);
xnor U20580 (N_20580,N_19624,N_19225);
and U20581 (N_20581,N_19168,N_19855);
or U20582 (N_20582,N_19912,N_19333);
and U20583 (N_20583,N_19014,N_19262);
xnor U20584 (N_20584,N_19809,N_19673);
nand U20585 (N_20585,N_19238,N_19803);
and U20586 (N_20586,N_19681,N_19713);
and U20587 (N_20587,N_19436,N_19725);
nor U20588 (N_20588,N_19395,N_19050);
or U20589 (N_20589,N_19157,N_19489);
nor U20590 (N_20590,N_19120,N_19636);
nand U20591 (N_20591,N_19166,N_19609);
nand U20592 (N_20592,N_19817,N_19427);
and U20593 (N_20593,N_19040,N_19054);
and U20594 (N_20594,N_19653,N_19865);
nand U20595 (N_20595,N_19650,N_19170);
or U20596 (N_20596,N_19293,N_19123);
nor U20597 (N_20597,N_19790,N_19262);
and U20598 (N_20598,N_19279,N_19512);
nand U20599 (N_20599,N_19652,N_19627);
nand U20600 (N_20600,N_19777,N_19301);
and U20601 (N_20601,N_19172,N_19842);
nor U20602 (N_20602,N_19583,N_19397);
xor U20603 (N_20603,N_19147,N_19126);
or U20604 (N_20604,N_19455,N_19282);
nand U20605 (N_20605,N_19015,N_19076);
xor U20606 (N_20606,N_19735,N_19797);
or U20607 (N_20607,N_19462,N_19262);
nor U20608 (N_20608,N_19124,N_19819);
nor U20609 (N_20609,N_19619,N_19593);
or U20610 (N_20610,N_19772,N_19951);
nor U20611 (N_20611,N_19105,N_19758);
and U20612 (N_20612,N_19131,N_19246);
nor U20613 (N_20613,N_19530,N_19972);
or U20614 (N_20614,N_19915,N_19201);
nand U20615 (N_20615,N_19117,N_19072);
nand U20616 (N_20616,N_19493,N_19139);
or U20617 (N_20617,N_19880,N_19071);
xnor U20618 (N_20618,N_19153,N_19764);
or U20619 (N_20619,N_19794,N_19313);
xor U20620 (N_20620,N_19485,N_19035);
nand U20621 (N_20621,N_19772,N_19159);
or U20622 (N_20622,N_19854,N_19628);
xnor U20623 (N_20623,N_19608,N_19769);
xor U20624 (N_20624,N_19550,N_19334);
nand U20625 (N_20625,N_19447,N_19403);
nor U20626 (N_20626,N_19916,N_19620);
nand U20627 (N_20627,N_19230,N_19459);
or U20628 (N_20628,N_19868,N_19303);
or U20629 (N_20629,N_19538,N_19414);
or U20630 (N_20630,N_19252,N_19649);
or U20631 (N_20631,N_19931,N_19760);
or U20632 (N_20632,N_19026,N_19923);
nand U20633 (N_20633,N_19064,N_19961);
or U20634 (N_20634,N_19870,N_19090);
or U20635 (N_20635,N_19639,N_19082);
xnor U20636 (N_20636,N_19317,N_19301);
xor U20637 (N_20637,N_19369,N_19913);
xnor U20638 (N_20638,N_19025,N_19695);
or U20639 (N_20639,N_19984,N_19826);
nand U20640 (N_20640,N_19707,N_19143);
nand U20641 (N_20641,N_19968,N_19145);
nand U20642 (N_20642,N_19248,N_19303);
xnor U20643 (N_20643,N_19030,N_19143);
nor U20644 (N_20644,N_19461,N_19413);
nor U20645 (N_20645,N_19575,N_19287);
nor U20646 (N_20646,N_19984,N_19404);
xnor U20647 (N_20647,N_19048,N_19693);
nor U20648 (N_20648,N_19614,N_19970);
nand U20649 (N_20649,N_19735,N_19519);
and U20650 (N_20650,N_19175,N_19430);
or U20651 (N_20651,N_19067,N_19556);
nand U20652 (N_20652,N_19746,N_19322);
nand U20653 (N_20653,N_19898,N_19741);
xnor U20654 (N_20654,N_19837,N_19569);
xnor U20655 (N_20655,N_19965,N_19928);
and U20656 (N_20656,N_19719,N_19888);
and U20657 (N_20657,N_19946,N_19131);
xnor U20658 (N_20658,N_19274,N_19074);
nor U20659 (N_20659,N_19354,N_19164);
xnor U20660 (N_20660,N_19940,N_19467);
nor U20661 (N_20661,N_19486,N_19019);
nor U20662 (N_20662,N_19424,N_19690);
or U20663 (N_20663,N_19618,N_19087);
or U20664 (N_20664,N_19331,N_19827);
xnor U20665 (N_20665,N_19379,N_19548);
or U20666 (N_20666,N_19819,N_19140);
or U20667 (N_20667,N_19626,N_19411);
or U20668 (N_20668,N_19388,N_19568);
or U20669 (N_20669,N_19938,N_19195);
and U20670 (N_20670,N_19389,N_19239);
and U20671 (N_20671,N_19693,N_19471);
or U20672 (N_20672,N_19573,N_19216);
nor U20673 (N_20673,N_19757,N_19358);
or U20674 (N_20674,N_19548,N_19139);
and U20675 (N_20675,N_19043,N_19487);
nand U20676 (N_20676,N_19494,N_19258);
xor U20677 (N_20677,N_19568,N_19461);
and U20678 (N_20678,N_19315,N_19616);
nand U20679 (N_20679,N_19110,N_19977);
and U20680 (N_20680,N_19811,N_19425);
nand U20681 (N_20681,N_19107,N_19156);
nand U20682 (N_20682,N_19189,N_19266);
xnor U20683 (N_20683,N_19787,N_19827);
xnor U20684 (N_20684,N_19574,N_19234);
or U20685 (N_20685,N_19026,N_19307);
xnor U20686 (N_20686,N_19265,N_19969);
and U20687 (N_20687,N_19658,N_19880);
and U20688 (N_20688,N_19067,N_19338);
xnor U20689 (N_20689,N_19037,N_19739);
and U20690 (N_20690,N_19569,N_19197);
or U20691 (N_20691,N_19296,N_19825);
nor U20692 (N_20692,N_19983,N_19597);
xnor U20693 (N_20693,N_19319,N_19875);
and U20694 (N_20694,N_19973,N_19913);
xor U20695 (N_20695,N_19090,N_19756);
and U20696 (N_20696,N_19724,N_19595);
nor U20697 (N_20697,N_19812,N_19749);
nor U20698 (N_20698,N_19837,N_19852);
and U20699 (N_20699,N_19841,N_19641);
or U20700 (N_20700,N_19405,N_19224);
nand U20701 (N_20701,N_19108,N_19838);
nand U20702 (N_20702,N_19957,N_19219);
nand U20703 (N_20703,N_19309,N_19509);
xnor U20704 (N_20704,N_19461,N_19255);
nand U20705 (N_20705,N_19114,N_19074);
nand U20706 (N_20706,N_19033,N_19183);
and U20707 (N_20707,N_19829,N_19218);
or U20708 (N_20708,N_19318,N_19327);
nand U20709 (N_20709,N_19234,N_19838);
xnor U20710 (N_20710,N_19875,N_19469);
xnor U20711 (N_20711,N_19563,N_19843);
and U20712 (N_20712,N_19786,N_19590);
nand U20713 (N_20713,N_19774,N_19482);
and U20714 (N_20714,N_19729,N_19969);
xnor U20715 (N_20715,N_19923,N_19518);
and U20716 (N_20716,N_19714,N_19510);
nand U20717 (N_20717,N_19752,N_19016);
nor U20718 (N_20718,N_19109,N_19917);
or U20719 (N_20719,N_19307,N_19993);
xnor U20720 (N_20720,N_19624,N_19673);
nor U20721 (N_20721,N_19829,N_19177);
or U20722 (N_20722,N_19611,N_19081);
nand U20723 (N_20723,N_19425,N_19001);
or U20724 (N_20724,N_19483,N_19261);
xnor U20725 (N_20725,N_19789,N_19364);
or U20726 (N_20726,N_19040,N_19723);
xor U20727 (N_20727,N_19781,N_19076);
xnor U20728 (N_20728,N_19321,N_19840);
nand U20729 (N_20729,N_19106,N_19802);
or U20730 (N_20730,N_19552,N_19584);
or U20731 (N_20731,N_19375,N_19278);
and U20732 (N_20732,N_19344,N_19757);
xnor U20733 (N_20733,N_19913,N_19847);
nand U20734 (N_20734,N_19552,N_19702);
or U20735 (N_20735,N_19907,N_19460);
xor U20736 (N_20736,N_19403,N_19121);
and U20737 (N_20737,N_19010,N_19992);
xor U20738 (N_20738,N_19877,N_19402);
or U20739 (N_20739,N_19369,N_19960);
xor U20740 (N_20740,N_19641,N_19607);
xnor U20741 (N_20741,N_19931,N_19445);
and U20742 (N_20742,N_19846,N_19555);
nor U20743 (N_20743,N_19398,N_19459);
nor U20744 (N_20744,N_19905,N_19811);
nor U20745 (N_20745,N_19624,N_19801);
xnor U20746 (N_20746,N_19600,N_19476);
nand U20747 (N_20747,N_19557,N_19250);
xor U20748 (N_20748,N_19159,N_19492);
or U20749 (N_20749,N_19116,N_19264);
xor U20750 (N_20750,N_19198,N_19495);
nand U20751 (N_20751,N_19444,N_19385);
or U20752 (N_20752,N_19888,N_19054);
or U20753 (N_20753,N_19475,N_19686);
and U20754 (N_20754,N_19666,N_19154);
nor U20755 (N_20755,N_19429,N_19093);
nor U20756 (N_20756,N_19683,N_19769);
and U20757 (N_20757,N_19951,N_19969);
or U20758 (N_20758,N_19419,N_19242);
nand U20759 (N_20759,N_19858,N_19258);
or U20760 (N_20760,N_19598,N_19870);
nand U20761 (N_20761,N_19736,N_19555);
nand U20762 (N_20762,N_19334,N_19427);
nand U20763 (N_20763,N_19317,N_19192);
nand U20764 (N_20764,N_19685,N_19644);
nor U20765 (N_20765,N_19987,N_19440);
xor U20766 (N_20766,N_19503,N_19138);
and U20767 (N_20767,N_19028,N_19701);
xnor U20768 (N_20768,N_19234,N_19776);
xnor U20769 (N_20769,N_19563,N_19033);
or U20770 (N_20770,N_19813,N_19463);
and U20771 (N_20771,N_19228,N_19022);
and U20772 (N_20772,N_19880,N_19010);
or U20773 (N_20773,N_19494,N_19808);
and U20774 (N_20774,N_19952,N_19475);
and U20775 (N_20775,N_19112,N_19000);
nand U20776 (N_20776,N_19197,N_19532);
nor U20777 (N_20777,N_19967,N_19301);
nand U20778 (N_20778,N_19429,N_19502);
nor U20779 (N_20779,N_19270,N_19517);
or U20780 (N_20780,N_19694,N_19172);
nand U20781 (N_20781,N_19364,N_19760);
and U20782 (N_20782,N_19436,N_19225);
and U20783 (N_20783,N_19134,N_19471);
nand U20784 (N_20784,N_19412,N_19020);
nand U20785 (N_20785,N_19072,N_19550);
xor U20786 (N_20786,N_19250,N_19021);
nor U20787 (N_20787,N_19070,N_19057);
and U20788 (N_20788,N_19379,N_19923);
nand U20789 (N_20789,N_19854,N_19015);
nand U20790 (N_20790,N_19311,N_19253);
xor U20791 (N_20791,N_19283,N_19541);
and U20792 (N_20792,N_19231,N_19768);
nand U20793 (N_20793,N_19779,N_19477);
or U20794 (N_20794,N_19540,N_19639);
nand U20795 (N_20795,N_19890,N_19872);
or U20796 (N_20796,N_19168,N_19598);
and U20797 (N_20797,N_19796,N_19723);
or U20798 (N_20798,N_19620,N_19111);
nand U20799 (N_20799,N_19965,N_19493);
and U20800 (N_20800,N_19459,N_19110);
nor U20801 (N_20801,N_19008,N_19155);
xnor U20802 (N_20802,N_19990,N_19506);
and U20803 (N_20803,N_19863,N_19046);
xor U20804 (N_20804,N_19616,N_19814);
or U20805 (N_20805,N_19380,N_19949);
nor U20806 (N_20806,N_19477,N_19194);
xnor U20807 (N_20807,N_19317,N_19931);
xor U20808 (N_20808,N_19016,N_19413);
or U20809 (N_20809,N_19001,N_19573);
nor U20810 (N_20810,N_19624,N_19144);
xnor U20811 (N_20811,N_19525,N_19554);
nand U20812 (N_20812,N_19495,N_19768);
xnor U20813 (N_20813,N_19216,N_19854);
and U20814 (N_20814,N_19640,N_19417);
or U20815 (N_20815,N_19341,N_19996);
and U20816 (N_20816,N_19901,N_19699);
and U20817 (N_20817,N_19372,N_19327);
xnor U20818 (N_20818,N_19621,N_19680);
xor U20819 (N_20819,N_19570,N_19955);
nor U20820 (N_20820,N_19495,N_19075);
nand U20821 (N_20821,N_19311,N_19738);
nand U20822 (N_20822,N_19517,N_19711);
and U20823 (N_20823,N_19678,N_19875);
nor U20824 (N_20824,N_19803,N_19675);
nand U20825 (N_20825,N_19967,N_19381);
nand U20826 (N_20826,N_19840,N_19824);
xnor U20827 (N_20827,N_19659,N_19995);
or U20828 (N_20828,N_19649,N_19752);
and U20829 (N_20829,N_19448,N_19344);
xor U20830 (N_20830,N_19848,N_19499);
or U20831 (N_20831,N_19215,N_19273);
and U20832 (N_20832,N_19972,N_19102);
xor U20833 (N_20833,N_19064,N_19814);
and U20834 (N_20834,N_19661,N_19334);
or U20835 (N_20835,N_19659,N_19841);
nor U20836 (N_20836,N_19545,N_19469);
xor U20837 (N_20837,N_19886,N_19919);
xnor U20838 (N_20838,N_19783,N_19118);
xor U20839 (N_20839,N_19628,N_19961);
nor U20840 (N_20840,N_19777,N_19856);
and U20841 (N_20841,N_19292,N_19327);
or U20842 (N_20842,N_19929,N_19405);
nor U20843 (N_20843,N_19147,N_19042);
nand U20844 (N_20844,N_19964,N_19835);
nor U20845 (N_20845,N_19478,N_19974);
xor U20846 (N_20846,N_19063,N_19313);
or U20847 (N_20847,N_19858,N_19384);
nor U20848 (N_20848,N_19545,N_19051);
and U20849 (N_20849,N_19323,N_19605);
or U20850 (N_20850,N_19332,N_19584);
xnor U20851 (N_20851,N_19797,N_19172);
xor U20852 (N_20852,N_19568,N_19558);
or U20853 (N_20853,N_19143,N_19587);
or U20854 (N_20854,N_19513,N_19707);
or U20855 (N_20855,N_19344,N_19379);
nor U20856 (N_20856,N_19222,N_19981);
and U20857 (N_20857,N_19674,N_19087);
and U20858 (N_20858,N_19286,N_19440);
nand U20859 (N_20859,N_19654,N_19899);
and U20860 (N_20860,N_19837,N_19041);
nor U20861 (N_20861,N_19197,N_19171);
or U20862 (N_20862,N_19319,N_19601);
xor U20863 (N_20863,N_19924,N_19467);
xor U20864 (N_20864,N_19384,N_19716);
or U20865 (N_20865,N_19866,N_19751);
or U20866 (N_20866,N_19323,N_19661);
or U20867 (N_20867,N_19849,N_19296);
nor U20868 (N_20868,N_19477,N_19031);
and U20869 (N_20869,N_19770,N_19153);
or U20870 (N_20870,N_19511,N_19852);
nor U20871 (N_20871,N_19040,N_19330);
or U20872 (N_20872,N_19599,N_19358);
nor U20873 (N_20873,N_19492,N_19836);
xnor U20874 (N_20874,N_19618,N_19706);
nor U20875 (N_20875,N_19524,N_19650);
xnor U20876 (N_20876,N_19990,N_19577);
or U20877 (N_20877,N_19397,N_19679);
and U20878 (N_20878,N_19694,N_19444);
nor U20879 (N_20879,N_19028,N_19870);
and U20880 (N_20880,N_19847,N_19219);
and U20881 (N_20881,N_19148,N_19824);
nor U20882 (N_20882,N_19778,N_19210);
or U20883 (N_20883,N_19837,N_19746);
xnor U20884 (N_20884,N_19214,N_19851);
and U20885 (N_20885,N_19988,N_19366);
xnor U20886 (N_20886,N_19119,N_19738);
xor U20887 (N_20887,N_19257,N_19901);
nor U20888 (N_20888,N_19310,N_19221);
nor U20889 (N_20889,N_19062,N_19807);
nand U20890 (N_20890,N_19558,N_19882);
and U20891 (N_20891,N_19739,N_19936);
xor U20892 (N_20892,N_19374,N_19958);
nor U20893 (N_20893,N_19709,N_19708);
nand U20894 (N_20894,N_19492,N_19605);
nor U20895 (N_20895,N_19593,N_19012);
xor U20896 (N_20896,N_19095,N_19575);
nand U20897 (N_20897,N_19480,N_19859);
and U20898 (N_20898,N_19333,N_19901);
xor U20899 (N_20899,N_19601,N_19100);
nand U20900 (N_20900,N_19410,N_19533);
nor U20901 (N_20901,N_19115,N_19593);
nor U20902 (N_20902,N_19989,N_19154);
and U20903 (N_20903,N_19616,N_19241);
nor U20904 (N_20904,N_19658,N_19268);
or U20905 (N_20905,N_19052,N_19667);
or U20906 (N_20906,N_19324,N_19479);
nand U20907 (N_20907,N_19611,N_19896);
nand U20908 (N_20908,N_19124,N_19176);
nand U20909 (N_20909,N_19023,N_19086);
nor U20910 (N_20910,N_19095,N_19803);
or U20911 (N_20911,N_19882,N_19058);
or U20912 (N_20912,N_19686,N_19398);
or U20913 (N_20913,N_19614,N_19455);
nor U20914 (N_20914,N_19882,N_19384);
xor U20915 (N_20915,N_19184,N_19675);
or U20916 (N_20916,N_19194,N_19711);
or U20917 (N_20917,N_19947,N_19637);
xnor U20918 (N_20918,N_19203,N_19496);
nor U20919 (N_20919,N_19305,N_19402);
or U20920 (N_20920,N_19093,N_19704);
and U20921 (N_20921,N_19897,N_19049);
nor U20922 (N_20922,N_19988,N_19345);
nor U20923 (N_20923,N_19387,N_19033);
and U20924 (N_20924,N_19236,N_19724);
or U20925 (N_20925,N_19038,N_19503);
xnor U20926 (N_20926,N_19077,N_19907);
xor U20927 (N_20927,N_19711,N_19985);
and U20928 (N_20928,N_19029,N_19314);
nand U20929 (N_20929,N_19071,N_19251);
and U20930 (N_20930,N_19509,N_19001);
xor U20931 (N_20931,N_19165,N_19533);
or U20932 (N_20932,N_19332,N_19313);
and U20933 (N_20933,N_19957,N_19028);
nor U20934 (N_20934,N_19855,N_19301);
and U20935 (N_20935,N_19101,N_19378);
xnor U20936 (N_20936,N_19831,N_19795);
nand U20937 (N_20937,N_19683,N_19198);
nor U20938 (N_20938,N_19985,N_19521);
and U20939 (N_20939,N_19017,N_19256);
or U20940 (N_20940,N_19901,N_19660);
nor U20941 (N_20941,N_19929,N_19067);
and U20942 (N_20942,N_19986,N_19558);
nor U20943 (N_20943,N_19379,N_19063);
xor U20944 (N_20944,N_19717,N_19315);
nor U20945 (N_20945,N_19599,N_19633);
or U20946 (N_20946,N_19661,N_19277);
xor U20947 (N_20947,N_19225,N_19830);
nor U20948 (N_20948,N_19587,N_19130);
nand U20949 (N_20949,N_19019,N_19656);
nor U20950 (N_20950,N_19192,N_19683);
nand U20951 (N_20951,N_19727,N_19815);
nor U20952 (N_20952,N_19142,N_19632);
nor U20953 (N_20953,N_19528,N_19711);
nor U20954 (N_20954,N_19398,N_19832);
nand U20955 (N_20955,N_19097,N_19970);
and U20956 (N_20956,N_19949,N_19521);
xor U20957 (N_20957,N_19948,N_19186);
and U20958 (N_20958,N_19251,N_19751);
nor U20959 (N_20959,N_19376,N_19257);
and U20960 (N_20960,N_19795,N_19834);
and U20961 (N_20961,N_19394,N_19308);
nor U20962 (N_20962,N_19592,N_19494);
xnor U20963 (N_20963,N_19805,N_19145);
nor U20964 (N_20964,N_19853,N_19804);
nand U20965 (N_20965,N_19966,N_19924);
or U20966 (N_20966,N_19660,N_19056);
xor U20967 (N_20967,N_19380,N_19175);
nand U20968 (N_20968,N_19663,N_19555);
and U20969 (N_20969,N_19254,N_19222);
nand U20970 (N_20970,N_19988,N_19404);
nand U20971 (N_20971,N_19014,N_19340);
and U20972 (N_20972,N_19606,N_19325);
xnor U20973 (N_20973,N_19597,N_19543);
and U20974 (N_20974,N_19972,N_19833);
or U20975 (N_20975,N_19339,N_19751);
nand U20976 (N_20976,N_19774,N_19903);
nor U20977 (N_20977,N_19006,N_19410);
nor U20978 (N_20978,N_19481,N_19864);
nor U20979 (N_20979,N_19616,N_19991);
nand U20980 (N_20980,N_19691,N_19662);
nand U20981 (N_20981,N_19615,N_19466);
nand U20982 (N_20982,N_19582,N_19395);
nand U20983 (N_20983,N_19489,N_19132);
nand U20984 (N_20984,N_19484,N_19586);
nand U20985 (N_20985,N_19840,N_19246);
nand U20986 (N_20986,N_19230,N_19945);
nand U20987 (N_20987,N_19160,N_19876);
nand U20988 (N_20988,N_19742,N_19001);
xnor U20989 (N_20989,N_19750,N_19522);
nor U20990 (N_20990,N_19457,N_19260);
nand U20991 (N_20991,N_19846,N_19158);
and U20992 (N_20992,N_19817,N_19103);
xor U20993 (N_20993,N_19933,N_19596);
nor U20994 (N_20994,N_19055,N_19866);
nor U20995 (N_20995,N_19679,N_19550);
or U20996 (N_20996,N_19685,N_19215);
nand U20997 (N_20997,N_19342,N_19934);
nand U20998 (N_20998,N_19690,N_19907);
and U20999 (N_20999,N_19088,N_19498);
and U21000 (N_21000,N_20401,N_20603);
or U21001 (N_21001,N_20069,N_20708);
or U21002 (N_21002,N_20344,N_20205);
or U21003 (N_21003,N_20658,N_20188);
and U21004 (N_21004,N_20670,N_20157);
nand U21005 (N_21005,N_20635,N_20215);
or U21006 (N_21006,N_20546,N_20363);
xnor U21007 (N_21007,N_20046,N_20616);
and U21008 (N_21008,N_20232,N_20963);
or U21009 (N_21009,N_20687,N_20089);
nor U21010 (N_21010,N_20324,N_20633);
nor U21011 (N_21011,N_20896,N_20561);
or U21012 (N_21012,N_20187,N_20384);
nand U21013 (N_21013,N_20202,N_20829);
or U21014 (N_21014,N_20494,N_20101);
nand U21015 (N_21015,N_20349,N_20530);
or U21016 (N_21016,N_20778,N_20292);
and U21017 (N_21017,N_20249,N_20541);
xor U21018 (N_21018,N_20956,N_20775);
and U21019 (N_21019,N_20440,N_20113);
and U21020 (N_21020,N_20964,N_20140);
xor U21021 (N_21021,N_20265,N_20914);
nand U21022 (N_21022,N_20005,N_20293);
xor U21023 (N_21023,N_20343,N_20091);
nand U21024 (N_21024,N_20594,N_20867);
nor U21025 (N_21025,N_20330,N_20998);
and U21026 (N_21026,N_20840,N_20455);
or U21027 (N_21027,N_20507,N_20536);
or U21028 (N_21028,N_20063,N_20605);
or U21029 (N_21029,N_20177,N_20134);
or U21030 (N_21030,N_20675,N_20250);
nand U21031 (N_21031,N_20820,N_20737);
nand U21032 (N_21032,N_20465,N_20464);
and U21033 (N_21033,N_20039,N_20419);
nor U21034 (N_21034,N_20656,N_20805);
nand U21035 (N_21035,N_20035,N_20962);
and U21036 (N_21036,N_20013,N_20207);
nand U21037 (N_21037,N_20789,N_20597);
nor U21038 (N_21038,N_20811,N_20348);
or U21039 (N_21039,N_20787,N_20604);
and U21040 (N_21040,N_20916,N_20154);
nor U21041 (N_21041,N_20759,N_20229);
xor U21042 (N_21042,N_20045,N_20326);
xor U21043 (N_21043,N_20935,N_20717);
nand U21044 (N_21044,N_20946,N_20844);
nand U21045 (N_21045,N_20548,N_20655);
nand U21046 (N_21046,N_20452,N_20160);
nor U21047 (N_21047,N_20025,N_20413);
xor U21048 (N_21048,N_20484,N_20142);
nand U21049 (N_21049,N_20256,N_20321);
and U21050 (N_21050,N_20125,N_20651);
or U21051 (N_21051,N_20190,N_20683);
and U21052 (N_21052,N_20501,N_20569);
and U21053 (N_21053,N_20924,N_20231);
nor U21054 (N_21054,N_20395,N_20736);
xnor U21055 (N_21055,N_20709,N_20741);
and U21056 (N_21056,N_20309,N_20814);
and U21057 (N_21057,N_20317,N_20941);
nand U21058 (N_21058,N_20711,N_20704);
nand U21059 (N_21059,N_20688,N_20463);
and U21060 (N_21060,N_20285,N_20839);
nand U21061 (N_21061,N_20692,N_20532);
and U21062 (N_21062,N_20365,N_20099);
or U21063 (N_21063,N_20334,N_20095);
and U21064 (N_21064,N_20796,N_20166);
or U21065 (N_21065,N_20209,N_20061);
nor U21066 (N_21066,N_20715,N_20499);
nor U21067 (N_21067,N_20891,N_20665);
or U21068 (N_21068,N_20108,N_20346);
nand U21069 (N_21069,N_20980,N_20087);
and U21070 (N_21070,N_20138,N_20024);
xor U21071 (N_21071,N_20011,N_20467);
or U21072 (N_21072,N_20412,N_20892);
nand U21073 (N_21073,N_20340,N_20034);
and U21074 (N_21074,N_20175,N_20682);
or U21075 (N_21075,N_20333,N_20298);
nand U21076 (N_21076,N_20905,N_20247);
xor U21077 (N_21077,N_20018,N_20632);
nor U21078 (N_21078,N_20408,N_20258);
nand U21079 (N_21079,N_20592,N_20766);
nor U21080 (N_21080,N_20922,N_20481);
nor U21081 (N_21081,N_20528,N_20184);
nor U21082 (N_21082,N_20828,N_20391);
or U21083 (N_21083,N_20729,N_20004);
or U21084 (N_21084,N_20386,N_20608);
or U21085 (N_21085,N_20919,N_20264);
or U21086 (N_21086,N_20885,N_20327);
nand U21087 (N_21087,N_20447,N_20826);
xnor U21088 (N_21088,N_20868,N_20429);
nor U21089 (N_21089,N_20007,N_20394);
nand U21090 (N_21090,N_20084,N_20792);
or U21091 (N_21091,N_20162,N_20626);
nor U21092 (N_21092,N_20690,N_20798);
or U21093 (N_21093,N_20918,N_20763);
and U21094 (N_21094,N_20492,N_20705);
nand U21095 (N_21095,N_20571,N_20942);
xnor U21096 (N_21096,N_20299,N_20300);
or U21097 (N_21097,N_20120,N_20197);
and U21098 (N_21098,N_20037,N_20760);
or U21099 (N_21099,N_20017,N_20920);
xor U21100 (N_21100,N_20949,N_20026);
nor U21101 (N_21101,N_20819,N_20927);
and U21102 (N_21102,N_20971,N_20361);
xor U21103 (N_21103,N_20446,N_20168);
xnor U21104 (N_21104,N_20731,N_20029);
or U21105 (N_21105,N_20454,N_20992);
or U21106 (N_21106,N_20518,N_20890);
nor U21107 (N_21107,N_20883,N_20315);
or U21108 (N_21108,N_20156,N_20102);
xor U21109 (N_21109,N_20572,N_20855);
nand U21110 (N_21110,N_20611,N_20195);
or U21111 (N_21111,N_20669,N_20031);
nand U21112 (N_21112,N_20750,N_20444);
nor U21113 (N_21113,N_20448,N_20978);
nand U21114 (N_21114,N_20392,N_20147);
xor U21115 (N_21115,N_20930,N_20472);
nand U21116 (N_21116,N_20505,N_20497);
nand U21117 (N_21117,N_20531,N_20566);
xnor U21118 (N_21118,N_20251,N_20500);
or U21119 (N_21119,N_20100,N_20957);
xnor U21120 (N_21120,N_20359,N_20923);
nand U21121 (N_21121,N_20578,N_20158);
xnor U21122 (N_21122,N_20053,N_20308);
nand U21123 (N_21123,N_20431,N_20771);
or U21124 (N_21124,N_20145,N_20637);
or U21125 (N_21125,N_20442,N_20719);
xnor U21126 (N_21126,N_20904,N_20027);
and U21127 (N_21127,N_20399,N_20712);
nor U21128 (N_21128,N_20153,N_20727);
and U21129 (N_21129,N_20353,N_20527);
nand U21130 (N_21130,N_20289,N_20404);
nand U21131 (N_21131,N_20559,N_20290);
or U21132 (N_21132,N_20791,N_20973);
nand U21133 (N_21133,N_20877,N_20420);
or U21134 (N_21134,N_20021,N_20104);
nand U21135 (N_21135,N_20986,N_20618);
and U21136 (N_21136,N_20533,N_20810);
xor U21137 (N_21137,N_20757,N_20485);
and U21138 (N_21138,N_20538,N_20426);
nor U21139 (N_21139,N_20714,N_20695);
xor U21140 (N_21140,N_20894,N_20549);
nor U21141 (N_21141,N_20267,N_20742);
nand U21142 (N_21142,N_20109,N_20224);
and U21143 (N_21143,N_20641,N_20539);
xor U21144 (N_21144,N_20174,N_20297);
xnor U21145 (N_21145,N_20807,N_20310);
nor U21146 (N_21146,N_20610,N_20774);
or U21147 (N_21147,N_20314,N_20248);
nand U21148 (N_21148,N_20913,N_20523);
nand U21149 (N_21149,N_20364,N_20576);
and U21150 (N_21150,N_20304,N_20457);
and U21151 (N_21151,N_20831,N_20932);
nand U21152 (N_21152,N_20550,N_20002);
and U21153 (N_21153,N_20861,N_20433);
xor U21154 (N_21154,N_20803,N_20794);
nand U21155 (N_21155,N_20048,N_20223);
nor U21156 (N_21156,N_20445,N_20137);
xnor U21157 (N_21157,N_20239,N_20979);
nand U21158 (N_21158,N_20164,N_20598);
nor U21159 (N_21159,N_20403,N_20222);
nor U21160 (N_21160,N_20697,N_20680);
xor U21161 (N_21161,N_20795,N_20133);
nor U21162 (N_21162,N_20393,N_20278);
nand U21163 (N_21163,N_20498,N_20331);
nor U21164 (N_21164,N_20886,N_20458);
xor U21165 (N_21165,N_20483,N_20995);
or U21166 (N_21166,N_20740,N_20191);
xnor U21167 (N_21167,N_20818,N_20000);
xor U21168 (N_21168,N_20303,N_20389);
nor U21169 (N_21169,N_20945,N_20192);
nor U21170 (N_21170,N_20614,N_20336);
nor U21171 (N_21171,N_20534,N_20767);
nor U21172 (N_21172,N_20354,N_20654);
or U21173 (N_21173,N_20241,N_20406);
nor U21174 (N_21174,N_20593,N_20874);
or U21175 (N_21175,N_20123,N_20178);
or U21176 (N_21176,N_20721,N_20753);
xor U21177 (N_21177,N_20277,N_20040);
or U21178 (N_21178,N_20985,N_20043);
xor U21179 (N_21179,N_20119,N_20306);
xor U21180 (N_21180,N_20684,N_20965);
nand U21181 (N_21181,N_20428,N_20764);
and U21182 (N_21182,N_20456,N_20989);
nand U21183 (N_21183,N_20397,N_20228);
and U21184 (N_21184,N_20510,N_20966);
nor U21185 (N_21185,N_20179,N_20718);
xor U21186 (N_21186,N_20014,N_20272);
and U21187 (N_21187,N_20678,N_20269);
or U21188 (N_21188,N_20167,N_20958);
nor U21189 (N_21189,N_20369,N_20136);
or U21190 (N_21190,N_20907,N_20893);
or U21191 (N_21191,N_20469,N_20345);
nor U21192 (N_21192,N_20252,N_20449);
and U21193 (N_21193,N_20490,N_20287);
xnor U21194 (N_21194,N_20944,N_20030);
and U21195 (N_21195,N_20882,N_20852);
xnor U21196 (N_21196,N_20329,N_20881);
and U21197 (N_21197,N_20747,N_20075);
nand U21198 (N_21198,N_20662,N_20400);
and U21199 (N_21199,N_20203,N_20567);
and U21200 (N_21200,N_20439,N_20562);
and U21201 (N_21201,N_20121,N_20044);
nand U21202 (N_21202,N_20902,N_20994);
nor U21203 (N_21203,N_20480,N_20263);
and U21204 (N_21204,N_20198,N_20319);
xnor U21205 (N_21205,N_20067,N_20009);
or U21206 (N_21206,N_20066,N_20612);
nand U21207 (N_21207,N_20887,N_20106);
or U21208 (N_21208,N_20148,N_20423);
nand U21209 (N_21209,N_20129,N_20948);
and U21210 (N_21210,N_20583,N_20540);
xnor U21211 (N_21211,N_20677,N_20783);
xor U21212 (N_21212,N_20318,N_20525);
and U21213 (N_21213,N_20451,N_20859);
nand U21214 (N_21214,N_20707,N_20643);
and U21215 (N_21215,N_20619,N_20652);
xnor U21216 (N_21216,N_20407,N_20065);
nand U21217 (N_21217,N_20720,N_20173);
nand U21218 (N_21218,N_20073,N_20151);
nor U21219 (N_21219,N_20291,N_20591);
or U21220 (N_21220,N_20806,N_20276);
nor U21221 (N_21221,N_20800,N_20915);
nor U21222 (N_21222,N_20357,N_20146);
nand U21223 (N_21223,N_20110,N_20127);
or U21224 (N_21224,N_20246,N_20194);
xor U21225 (N_21225,N_20813,N_20414);
nor U21226 (N_21226,N_20543,N_20496);
nand U21227 (N_21227,N_20097,N_20889);
and U21228 (N_21228,N_20150,N_20060);
xnor U21229 (N_21229,N_20899,N_20878);
nand U21230 (N_21230,N_20186,N_20661);
nand U21231 (N_21231,N_20556,N_20599);
or U21232 (N_21232,N_20141,N_20488);
xor U21233 (N_21233,N_20430,N_20785);
or U21234 (N_21234,N_20696,N_20522);
xor U21235 (N_21235,N_20282,N_20274);
xnor U21236 (N_21236,N_20216,N_20910);
or U21237 (N_21237,N_20520,N_20671);
and U21238 (N_21238,N_20237,N_20159);
or U21239 (N_21239,N_20921,N_20529);
or U21240 (N_21240,N_20926,N_20461);
and U21241 (N_21241,N_20897,N_20863);
or U21242 (N_21242,N_20617,N_20450);
nand U21243 (N_21243,N_20751,N_20879);
nor U21244 (N_21244,N_20375,N_20663);
xnor U21245 (N_21245,N_20460,N_20574);
nor U21246 (N_21246,N_20107,N_20088);
or U21247 (N_21247,N_20041,N_20743);
nand U21248 (N_21248,N_20441,N_20875);
or U21249 (N_21249,N_20575,N_20230);
nor U21250 (N_21250,N_20557,N_20555);
nand U21251 (N_21251,N_20302,N_20581);
and U21252 (N_21252,N_20837,N_20937);
nor U21253 (N_21253,N_20493,N_20316);
or U21254 (N_21254,N_20211,N_20479);
nor U21255 (N_21255,N_20212,N_20952);
nand U21256 (N_21256,N_20733,N_20631);
xnor U21257 (N_21257,N_20755,N_20858);
and U21258 (N_21258,N_20266,N_20325);
and U21259 (N_21259,N_20917,N_20201);
nor U21260 (N_21260,N_20155,N_20967);
xnor U21261 (N_21261,N_20323,N_20782);
nor U21262 (N_21262,N_20240,N_20513);
and U21263 (N_21263,N_20898,N_20925);
xnor U21264 (N_21264,N_20724,N_20681);
xnor U21265 (N_21265,N_20975,N_20242);
and U21266 (N_21266,N_20347,N_20380);
or U21267 (N_21267,N_20078,N_20773);
nor U21268 (N_21268,N_20723,N_20509);
nor U21269 (N_21269,N_20368,N_20587);
xor U21270 (N_21270,N_20243,N_20929);
and U21271 (N_21271,N_20648,N_20585);
and U21272 (N_21272,N_20257,N_20990);
nand U21273 (N_21273,N_20953,N_20884);
nand U21274 (N_21274,N_20294,N_20570);
xnor U21275 (N_21275,N_20385,N_20777);
nand U21276 (N_21276,N_20642,N_20432);
xnor U21277 (N_21277,N_20869,N_20126);
nor U21278 (N_21278,N_20728,N_20114);
xor U21279 (N_21279,N_20906,N_20422);
xor U21280 (N_21280,N_20185,N_20332);
nand U21281 (N_21281,N_20606,N_20558);
and U21282 (N_21282,N_20372,N_20573);
xnor U21283 (N_21283,N_20313,N_20503);
nor U21284 (N_21284,N_20281,N_20674);
nand U21285 (N_21285,N_20815,N_20615);
nor U21286 (N_21286,N_20352,N_20809);
xnor U21287 (N_21287,N_20337,N_20279);
and U21288 (N_21288,N_20780,N_20568);
nor U21289 (N_21289,N_20744,N_20471);
or U21290 (N_21290,N_20105,N_20748);
and U21291 (N_21291,N_20700,N_20416);
or U21292 (N_21292,N_20758,N_20713);
nor U21293 (N_21293,N_20193,N_20703);
xnor U21294 (N_21294,N_20038,N_20475);
xor U21295 (N_21295,N_20183,N_20342);
or U21296 (N_21296,N_20835,N_20676);
nand U21297 (N_21297,N_20981,N_20974);
and U21298 (N_21298,N_20931,N_20554);
or U21299 (N_21299,N_20999,N_20589);
and U21300 (N_21300,N_20311,N_20634);
nor U21301 (N_21301,N_20873,N_20453);
and U21302 (N_21302,N_20094,N_20116);
xnor U21303 (N_21303,N_20478,N_20350);
nor U21304 (N_21304,N_20786,N_20830);
nand U21305 (N_21305,N_20378,N_20756);
or U21306 (N_21306,N_20639,N_20176);
or U21307 (N_21307,N_20398,N_20489);
nor U21308 (N_21308,N_20424,N_20630);
or U21309 (N_21309,N_20977,N_20486);
nor U21310 (N_21310,N_20491,N_20836);
nand U21311 (N_21311,N_20959,N_20772);
or U21312 (N_21312,N_20996,N_20565);
nor U21313 (N_21313,N_20822,N_20117);
and U21314 (N_21314,N_20847,N_20866);
xor U21315 (N_21315,N_20210,N_20693);
and U21316 (N_21316,N_20646,N_20181);
nor U21317 (N_21317,N_20022,N_20411);
xor U21318 (N_21318,N_20801,N_20227);
or U21319 (N_21319,N_20305,N_20495);
nand U21320 (N_21320,N_20664,N_20745);
nor U21321 (N_21321,N_20746,N_20244);
and U21322 (N_21322,N_20936,N_20577);
nand U21323 (N_21323,N_20010,N_20609);
nor U21324 (N_21324,N_20584,N_20901);
nor U21325 (N_21325,N_20221,N_20908);
nor U21326 (N_21326,N_20301,N_20793);
xor U21327 (N_21327,N_20988,N_20508);
or U21328 (N_21328,N_20872,N_20636);
nand U21329 (N_21329,N_20547,N_20003);
or U21330 (N_21330,N_20172,N_20535);
and U21331 (N_21331,N_20976,N_20328);
xnor U21332 (N_21332,N_20895,N_20169);
and U21333 (N_21333,N_20074,N_20388);
nand U21334 (N_21334,N_20351,N_20888);
nor U21335 (N_21335,N_20238,N_20358);
xor U21336 (N_21336,N_20033,N_20443);
or U21337 (N_21337,N_20402,N_20725);
and U21338 (N_21338,N_20832,N_20738);
and U21339 (N_21339,N_20551,N_20233);
or U21340 (N_21340,N_20286,N_20991);
nor U21341 (N_21341,N_20132,N_20544);
and U21342 (N_21342,N_20236,N_20685);
xor U21343 (N_21343,N_20468,N_20812);
nor U21344 (N_21344,N_20752,N_20841);
xnor U21345 (N_21345,N_20607,N_20502);
or U21346 (N_21346,N_20200,N_20434);
and U21347 (N_21347,N_20843,N_20993);
and U21348 (N_21348,N_20362,N_20032);
xnor U21349 (N_21349,N_20161,N_20370);
nand U21350 (N_21350,N_20254,N_20876);
nand U21351 (N_21351,N_20245,N_20042);
nand U21352 (N_21352,N_20784,N_20415);
nor U21353 (N_21353,N_20487,N_20366);
and U21354 (N_21354,N_20821,N_20387);
nor U21355 (N_21355,N_20122,N_20950);
nor U21356 (N_21356,N_20182,N_20081);
or U21357 (N_21357,N_20880,N_20622);
xor U21358 (N_21358,N_20051,N_20058);
or U21359 (N_21359,N_20799,N_20553);
nor U21360 (N_21360,N_20854,N_20059);
and U21361 (N_21361,N_20268,N_20170);
nor U21362 (N_21362,N_20262,N_20580);
xor U21363 (N_21363,N_20943,N_20001);
nand U21364 (N_21364,N_20280,N_20640);
and U21365 (N_21365,N_20694,N_20860);
and U21366 (N_21366,N_20056,N_20912);
or U21367 (N_21367,N_20997,N_20524);
xnor U21368 (N_21368,N_20470,N_20911);
or U21369 (N_21369,N_20410,N_20526);
xor U21370 (N_21370,N_20797,N_20545);
xnor U21371 (N_21371,N_20620,N_20947);
nor U21372 (N_21372,N_20008,N_20706);
xor U21373 (N_21373,N_20335,N_20726);
xor U21374 (N_21374,N_20776,N_20769);
or U21375 (N_21375,N_20217,N_20506);
nor U21376 (N_21376,N_20903,N_20438);
xnor U21377 (N_21377,N_20307,N_20650);
xor U21378 (N_21378,N_20939,N_20668);
nand U21379 (N_21379,N_20851,N_20864);
and U21380 (N_21380,N_20928,N_20761);
nand U21381 (N_21381,N_20749,N_20218);
xnor U21382 (N_21382,N_20339,N_20862);
and U21383 (N_21383,N_20588,N_20982);
nand U21384 (N_21384,N_20940,N_20621);
nor U21385 (N_21385,N_20261,N_20124);
and U21386 (N_21386,N_20020,N_20647);
nor U21387 (N_21387,N_20322,N_20225);
or U21388 (N_21388,N_20199,N_20055);
nand U21389 (N_21389,N_20679,N_20625);
xor U21390 (N_21390,N_20377,N_20425);
xor U21391 (N_21391,N_20077,N_20660);
and U21392 (N_21392,N_20827,N_20673);
nand U21393 (N_21393,N_20131,N_20514);
xor U21394 (N_21394,N_20071,N_20735);
nor U21395 (N_21395,N_20072,N_20015);
nor U21396 (N_21396,N_20984,N_20381);
xor U21397 (N_21397,N_20938,N_20515);
or U21398 (N_21398,N_20054,N_20590);
nor U21399 (N_21399,N_20367,N_20824);
nand U21400 (N_21400,N_20437,N_20698);
and U21401 (N_21401,N_20080,N_20701);
xor U21402 (N_21402,N_20270,N_20466);
xor U21403 (N_21403,N_20716,N_20112);
and U21404 (N_21404,N_20085,N_20057);
xnor U21405 (N_21405,N_20560,N_20103);
nor U21406 (N_21406,N_20070,N_20260);
nand U21407 (N_21407,N_20838,N_20405);
nand U21408 (N_21408,N_20968,N_20552);
or U21409 (N_21409,N_20722,N_20788);
nand U21410 (N_21410,N_20563,N_20804);
nor U21411 (N_21411,N_20208,N_20595);
or U21412 (N_21412,N_20226,N_20739);
or U21413 (N_21413,N_20050,N_20143);
or U21414 (N_21414,N_20064,N_20770);
or U21415 (N_21415,N_20111,N_20295);
nand U21416 (N_21416,N_20600,N_20834);
xor U21417 (N_21417,N_20710,N_20171);
nor U21418 (N_21418,N_20234,N_20355);
nand U21419 (N_21419,N_20283,N_20960);
xor U21420 (N_21420,N_20320,N_20093);
and U21421 (N_21421,N_20833,N_20613);
xnor U21422 (N_21422,N_20667,N_20383);
nor U21423 (N_21423,N_20016,N_20219);
nor U21424 (N_21424,N_20586,N_20052);
and U21425 (N_21425,N_20012,N_20418);
and U21426 (N_21426,N_20645,N_20204);
nand U21427 (N_21427,N_20933,N_20275);
and U21428 (N_21428,N_20427,N_20849);
or U21429 (N_21429,N_20220,N_20396);
xnor U21430 (N_21430,N_20196,N_20983);
xnor U21431 (N_21431,N_20649,N_20781);
or U21432 (N_21432,N_20213,N_20601);
or U21433 (N_21433,N_20163,N_20180);
nor U21434 (N_21434,N_20582,N_20288);
xor U21435 (N_21435,N_20028,N_20462);
or U21436 (N_21436,N_20823,N_20672);
nor U21437 (N_21437,N_20476,N_20596);
or U21438 (N_21438,N_20564,N_20730);
xor U21439 (N_21439,N_20130,N_20699);
and U21440 (N_21440,N_20047,N_20579);
xnor U21441 (N_21441,N_20341,N_20689);
or U21442 (N_21442,N_20623,N_20846);
nand U21443 (N_21443,N_20909,N_20421);
or U21444 (N_21444,N_20006,N_20023);
or U21445 (N_21445,N_20951,N_20284);
or U21446 (N_21446,N_20374,N_20090);
nand U21447 (N_21447,N_20638,N_20371);
or U21448 (N_21448,N_20259,N_20691);
nor U21449 (N_21449,N_20519,N_20086);
xnor U21450 (N_21450,N_20653,N_20845);
and U21451 (N_21451,N_20768,N_20360);
nand U21452 (N_21452,N_20356,N_20082);
nor U21453 (N_21453,N_20808,N_20624);
nor U21454 (N_21454,N_20850,N_20629);
xor U21455 (N_21455,N_20765,N_20144);
nor U21456 (N_21456,N_20762,N_20602);
or U21457 (N_21457,N_20165,N_20790);
nand U21458 (N_21458,N_20235,N_20152);
and U21459 (N_21459,N_20871,N_20214);
xnor U21460 (N_21460,N_20816,N_20754);
xor U21461 (N_21461,N_20273,N_20390);
or U21462 (N_21462,N_20092,N_20537);
nand U21463 (N_21463,N_20036,N_20856);
nand U21464 (N_21464,N_20857,N_20644);
xor U21465 (N_21465,N_20477,N_20068);
or U21466 (N_21466,N_20189,N_20096);
nor U21467 (N_21467,N_20961,N_20296);
or U21468 (N_21468,N_20521,N_20512);
xnor U21469 (N_21469,N_20049,N_20079);
and U21470 (N_21470,N_20865,N_20139);
or U21471 (N_21471,N_20459,N_20409);
or U21472 (N_21472,N_20482,N_20870);
and U21473 (N_21473,N_20842,N_20970);
nand U21474 (N_21474,N_20934,N_20417);
and U21475 (N_21475,N_20376,N_20955);
nor U21476 (N_21476,N_20825,N_20382);
xor U21477 (N_21477,N_20817,N_20734);
nor U21478 (N_21478,N_20373,N_20253);
nor U21479 (N_21479,N_20516,N_20802);
and U21480 (N_21480,N_20019,N_20436);
nor U21481 (N_21481,N_20732,N_20118);
and U21482 (N_21482,N_20628,N_20206);
xnor U21483 (N_21483,N_20083,N_20969);
xnor U21484 (N_21484,N_20473,N_20135);
or U21485 (N_21485,N_20255,N_20987);
and U21486 (N_21486,N_20312,N_20511);
nor U21487 (N_21487,N_20954,N_20659);
xor U21488 (N_21488,N_20338,N_20504);
or U21489 (N_21489,N_20779,N_20076);
nor U21490 (N_21490,N_20271,N_20379);
xor U21491 (N_21491,N_20627,N_20062);
nor U21492 (N_21492,N_20542,N_20853);
and U21493 (N_21493,N_20435,N_20972);
and U21494 (N_21494,N_20517,N_20128);
nand U21495 (N_21495,N_20098,N_20702);
nand U21496 (N_21496,N_20657,N_20474);
xnor U21497 (N_21497,N_20848,N_20686);
or U21498 (N_21498,N_20900,N_20115);
or U21499 (N_21499,N_20149,N_20666);
nand U21500 (N_21500,N_20844,N_20646);
xor U21501 (N_21501,N_20056,N_20939);
nand U21502 (N_21502,N_20824,N_20703);
nand U21503 (N_21503,N_20512,N_20376);
xnor U21504 (N_21504,N_20516,N_20094);
nand U21505 (N_21505,N_20392,N_20073);
nor U21506 (N_21506,N_20576,N_20122);
nor U21507 (N_21507,N_20772,N_20253);
or U21508 (N_21508,N_20460,N_20515);
nor U21509 (N_21509,N_20086,N_20200);
nor U21510 (N_21510,N_20000,N_20945);
nand U21511 (N_21511,N_20386,N_20781);
nor U21512 (N_21512,N_20175,N_20684);
nor U21513 (N_21513,N_20665,N_20376);
nand U21514 (N_21514,N_20639,N_20978);
xor U21515 (N_21515,N_20245,N_20201);
and U21516 (N_21516,N_20926,N_20021);
nor U21517 (N_21517,N_20352,N_20282);
xor U21518 (N_21518,N_20049,N_20921);
xnor U21519 (N_21519,N_20303,N_20867);
nand U21520 (N_21520,N_20473,N_20333);
and U21521 (N_21521,N_20683,N_20498);
and U21522 (N_21522,N_20240,N_20765);
or U21523 (N_21523,N_20328,N_20341);
and U21524 (N_21524,N_20012,N_20597);
nor U21525 (N_21525,N_20738,N_20764);
and U21526 (N_21526,N_20515,N_20313);
nand U21527 (N_21527,N_20609,N_20751);
nor U21528 (N_21528,N_20611,N_20389);
or U21529 (N_21529,N_20514,N_20755);
nor U21530 (N_21530,N_20188,N_20475);
nand U21531 (N_21531,N_20280,N_20705);
xor U21532 (N_21532,N_20871,N_20344);
and U21533 (N_21533,N_20810,N_20187);
xor U21534 (N_21534,N_20782,N_20154);
or U21535 (N_21535,N_20373,N_20608);
xor U21536 (N_21536,N_20245,N_20753);
and U21537 (N_21537,N_20719,N_20830);
xnor U21538 (N_21538,N_20631,N_20395);
nand U21539 (N_21539,N_20087,N_20042);
nor U21540 (N_21540,N_20347,N_20116);
xor U21541 (N_21541,N_20841,N_20965);
nor U21542 (N_21542,N_20935,N_20584);
nor U21543 (N_21543,N_20625,N_20937);
and U21544 (N_21544,N_20569,N_20023);
or U21545 (N_21545,N_20848,N_20031);
and U21546 (N_21546,N_20990,N_20723);
xnor U21547 (N_21547,N_20764,N_20719);
and U21548 (N_21548,N_20021,N_20612);
nand U21549 (N_21549,N_20970,N_20600);
nand U21550 (N_21550,N_20133,N_20843);
xnor U21551 (N_21551,N_20681,N_20390);
and U21552 (N_21552,N_20711,N_20236);
xor U21553 (N_21553,N_20132,N_20009);
or U21554 (N_21554,N_20666,N_20937);
xor U21555 (N_21555,N_20526,N_20776);
and U21556 (N_21556,N_20157,N_20721);
nor U21557 (N_21557,N_20698,N_20408);
or U21558 (N_21558,N_20101,N_20370);
xnor U21559 (N_21559,N_20042,N_20223);
or U21560 (N_21560,N_20133,N_20572);
xnor U21561 (N_21561,N_20000,N_20410);
or U21562 (N_21562,N_20998,N_20187);
nand U21563 (N_21563,N_20617,N_20044);
xnor U21564 (N_21564,N_20254,N_20290);
and U21565 (N_21565,N_20427,N_20236);
xnor U21566 (N_21566,N_20772,N_20224);
and U21567 (N_21567,N_20755,N_20049);
xnor U21568 (N_21568,N_20305,N_20645);
and U21569 (N_21569,N_20275,N_20831);
nor U21570 (N_21570,N_20186,N_20374);
nor U21571 (N_21571,N_20607,N_20796);
xnor U21572 (N_21572,N_20892,N_20349);
nand U21573 (N_21573,N_20631,N_20743);
or U21574 (N_21574,N_20126,N_20345);
or U21575 (N_21575,N_20567,N_20738);
xor U21576 (N_21576,N_20829,N_20651);
nand U21577 (N_21577,N_20714,N_20038);
and U21578 (N_21578,N_20831,N_20407);
and U21579 (N_21579,N_20352,N_20566);
or U21580 (N_21580,N_20212,N_20769);
or U21581 (N_21581,N_20215,N_20525);
or U21582 (N_21582,N_20692,N_20661);
nor U21583 (N_21583,N_20824,N_20712);
nand U21584 (N_21584,N_20209,N_20950);
xor U21585 (N_21585,N_20825,N_20480);
and U21586 (N_21586,N_20541,N_20847);
nor U21587 (N_21587,N_20022,N_20335);
nor U21588 (N_21588,N_20484,N_20711);
or U21589 (N_21589,N_20270,N_20189);
and U21590 (N_21590,N_20747,N_20750);
and U21591 (N_21591,N_20694,N_20164);
or U21592 (N_21592,N_20305,N_20943);
nand U21593 (N_21593,N_20611,N_20433);
xor U21594 (N_21594,N_20621,N_20563);
nor U21595 (N_21595,N_20789,N_20368);
nand U21596 (N_21596,N_20320,N_20088);
nand U21597 (N_21597,N_20161,N_20921);
and U21598 (N_21598,N_20183,N_20326);
nand U21599 (N_21599,N_20914,N_20758);
and U21600 (N_21600,N_20729,N_20564);
or U21601 (N_21601,N_20050,N_20132);
xor U21602 (N_21602,N_20458,N_20062);
and U21603 (N_21603,N_20459,N_20033);
nand U21604 (N_21604,N_20592,N_20073);
nor U21605 (N_21605,N_20425,N_20985);
and U21606 (N_21606,N_20701,N_20351);
or U21607 (N_21607,N_20110,N_20898);
nand U21608 (N_21608,N_20058,N_20094);
and U21609 (N_21609,N_20695,N_20105);
nand U21610 (N_21610,N_20749,N_20797);
nor U21611 (N_21611,N_20148,N_20795);
nor U21612 (N_21612,N_20015,N_20355);
nor U21613 (N_21613,N_20134,N_20291);
xor U21614 (N_21614,N_20653,N_20973);
and U21615 (N_21615,N_20382,N_20456);
or U21616 (N_21616,N_20444,N_20746);
nor U21617 (N_21617,N_20180,N_20406);
xor U21618 (N_21618,N_20980,N_20640);
or U21619 (N_21619,N_20324,N_20893);
xnor U21620 (N_21620,N_20524,N_20617);
or U21621 (N_21621,N_20344,N_20528);
xor U21622 (N_21622,N_20286,N_20129);
xor U21623 (N_21623,N_20989,N_20982);
xor U21624 (N_21624,N_20399,N_20533);
and U21625 (N_21625,N_20038,N_20261);
xnor U21626 (N_21626,N_20780,N_20433);
nand U21627 (N_21627,N_20697,N_20583);
nand U21628 (N_21628,N_20336,N_20807);
nand U21629 (N_21629,N_20384,N_20411);
nor U21630 (N_21630,N_20929,N_20109);
nor U21631 (N_21631,N_20877,N_20607);
xnor U21632 (N_21632,N_20092,N_20157);
nor U21633 (N_21633,N_20995,N_20537);
xor U21634 (N_21634,N_20348,N_20401);
xnor U21635 (N_21635,N_20149,N_20655);
nand U21636 (N_21636,N_20142,N_20176);
and U21637 (N_21637,N_20312,N_20085);
and U21638 (N_21638,N_20659,N_20178);
or U21639 (N_21639,N_20134,N_20053);
nand U21640 (N_21640,N_20456,N_20209);
or U21641 (N_21641,N_20455,N_20937);
nor U21642 (N_21642,N_20377,N_20665);
nand U21643 (N_21643,N_20869,N_20185);
nand U21644 (N_21644,N_20472,N_20680);
or U21645 (N_21645,N_20670,N_20747);
nand U21646 (N_21646,N_20738,N_20151);
or U21647 (N_21647,N_20332,N_20153);
xnor U21648 (N_21648,N_20153,N_20808);
and U21649 (N_21649,N_20124,N_20700);
xor U21650 (N_21650,N_20557,N_20719);
nand U21651 (N_21651,N_20090,N_20517);
xor U21652 (N_21652,N_20906,N_20723);
nand U21653 (N_21653,N_20928,N_20660);
or U21654 (N_21654,N_20595,N_20953);
xor U21655 (N_21655,N_20897,N_20942);
nor U21656 (N_21656,N_20414,N_20534);
xnor U21657 (N_21657,N_20348,N_20058);
xor U21658 (N_21658,N_20411,N_20176);
nor U21659 (N_21659,N_20290,N_20899);
nand U21660 (N_21660,N_20330,N_20758);
nand U21661 (N_21661,N_20827,N_20947);
nand U21662 (N_21662,N_20970,N_20564);
nor U21663 (N_21663,N_20176,N_20841);
and U21664 (N_21664,N_20431,N_20374);
nand U21665 (N_21665,N_20755,N_20656);
nor U21666 (N_21666,N_20778,N_20002);
xor U21667 (N_21667,N_20989,N_20969);
and U21668 (N_21668,N_20036,N_20799);
or U21669 (N_21669,N_20992,N_20980);
nand U21670 (N_21670,N_20990,N_20873);
nand U21671 (N_21671,N_20498,N_20892);
and U21672 (N_21672,N_20467,N_20705);
xnor U21673 (N_21673,N_20576,N_20906);
nand U21674 (N_21674,N_20955,N_20618);
and U21675 (N_21675,N_20380,N_20863);
and U21676 (N_21676,N_20960,N_20817);
xnor U21677 (N_21677,N_20625,N_20405);
nor U21678 (N_21678,N_20316,N_20821);
nor U21679 (N_21679,N_20447,N_20271);
nor U21680 (N_21680,N_20627,N_20999);
and U21681 (N_21681,N_20129,N_20988);
xor U21682 (N_21682,N_20412,N_20825);
nand U21683 (N_21683,N_20519,N_20317);
xnor U21684 (N_21684,N_20817,N_20571);
nor U21685 (N_21685,N_20814,N_20653);
nor U21686 (N_21686,N_20590,N_20061);
nor U21687 (N_21687,N_20683,N_20592);
nand U21688 (N_21688,N_20636,N_20307);
and U21689 (N_21689,N_20818,N_20542);
or U21690 (N_21690,N_20306,N_20309);
nand U21691 (N_21691,N_20427,N_20277);
and U21692 (N_21692,N_20076,N_20717);
and U21693 (N_21693,N_20535,N_20106);
xnor U21694 (N_21694,N_20350,N_20914);
nor U21695 (N_21695,N_20412,N_20329);
nor U21696 (N_21696,N_20185,N_20689);
and U21697 (N_21697,N_20214,N_20195);
or U21698 (N_21698,N_20877,N_20641);
nor U21699 (N_21699,N_20191,N_20785);
or U21700 (N_21700,N_20361,N_20974);
xnor U21701 (N_21701,N_20243,N_20920);
nand U21702 (N_21702,N_20771,N_20740);
xnor U21703 (N_21703,N_20925,N_20776);
xnor U21704 (N_21704,N_20065,N_20694);
and U21705 (N_21705,N_20469,N_20177);
xnor U21706 (N_21706,N_20762,N_20568);
or U21707 (N_21707,N_20883,N_20892);
nor U21708 (N_21708,N_20354,N_20309);
or U21709 (N_21709,N_20640,N_20320);
xnor U21710 (N_21710,N_20556,N_20820);
xor U21711 (N_21711,N_20224,N_20501);
nor U21712 (N_21712,N_20070,N_20561);
nor U21713 (N_21713,N_20105,N_20090);
nand U21714 (N_21714,N_20121,N_20139);
xnor U21715 (N_21715,N_20509,N_20189);
or U21716 (N_21716,N_20721,N_20989);
and U21717 (N_21717,N_20801,N_20970);
nor U21718 (N_21718,N_20492,N_20034);
or U21719 (N_21719,N_20936,N_20449);
xor U21720 (N_21720,N_20148,N_20134);
and U21721 (N_21721,N_20132,N_20612);
and U21722 (N_21722,N_20909,N_20282);
xor U21723 (N_21723,N_20204,N_20018);
nand U21724 (N_21724,N_20060,N_20175);
nor U21725 (N_21725,N_20567,N_20944);
and U21726 (N_21726,N_20902,N_20125);
or U21727 (N_21727,N_20760,N_20851);
xor U21728 (N_21728,N_20873,N_20803);
and U21729 (N_21729,N_20190,N_20935);
xnor U21730 (N_21730,N_20108,N_20265);
xor U21731 (N_21731,N_20275,N_20348);
nand U21732 (N_21732,N_20875,N_20001);
xor U21733 (N_21733,N_20578,N_20418);
xnor U21734 (N_21734,N_20921,N_20915);
and U21735 (N_21735,N_20051,N_20407);
and U21736 (N_21736,N_20311,N_20356);
nand U21737 (N_21737,N_20699,N_20857);
and U21738 (N_21738,N_20811,N_20301);
nand U21739 (N_21739,N_20610,N_20417);
nor U21740 (N_21740,N_20408,N_20315);
or U21741 (N_21741,N_20098,N_20048);
and U21742 (N_21742,N_20303,N_20845);
nand U21743 (N_21743,N_20040,N_20225);
nor U21744 (N_21744,N_20714,N_20361);
nor U21745 (N_21745,N_20446,N_20621);
and U21746 (N_21746,N_20857,N_20753);
and U21747 (N_21747,N_20210,N_20397);
xnor U21748 (N_21748,N_20782,N_20183);
nor U21749 (N_21749,N_20940,N_20240);
or U21750 (N_21750,N_20937,N_20962);
nor U21751 (N_21751,N_20805,N_20673);
and U21752 (N_21752,N_20967,N_20595);
nor U21753 (N_21753,N_20904,N_20862);
xor U21754 (N_21754,N_20972,N_20635);
or U21755 (N_21755,N_20267,N_20151);
nor U21756 (N_21756,N_20096,N_20523);
and U21757 (N_21757,N_20116,N_20863);
xor U21758 (N_21758,N_20329,N_20887);
nor U21759 (N_21759,N_20090,N_20171);
xnor U21760 (N_21760,N_20940,N_20866);
nand U21761 (N_21761,N_20090,N_20646);
nor U21762 (N_21762,N_20869,N_20200);
or U21763 (N_21763,N_20316,N_20611);
xnor U21764 (N_21764,N_20888,N_20322);
or U21765 (N_21765,N_20709,N_20440);
nand U21766 (N_21766,N_20390,N_20641);
xor U21767 (N_21767,N_20176,N_20429);
or U21768 (N_21768,N_20809,N_20691);
or U21769 (N_21769,N_20912,N_20150);
nand U21770 (N_21770,N_20995,N_20265);
xnor U21771 (N_21771,N_20768,N_20172);
and U21772 (N_21772,N_20842,N_20538);
nand U21773 (N_21773,N_20318,N_20773);
nand U21774 (N_21774,N_20690,N_20348);
and U21775 (N_21775,N_20250,N_20555);
or U21776 (N_21776,N_20468,N_20040);
nor U21777 (N_21777,N_20839,N_20995);
or U21778 (N_21778,N_20136,N_20532);
or U21779 (N_21779,N_20406,N_20092);
nand U21780 (N_21780,N_20617,N_20730);
nor U21781 (N_21781,N_20030,N_20655);
xor U21782 (N_21782,N_20735,N_20448);
xnor U21783 (N_21783,N_20166,N_20082);
or U21784 (N_21784,N_20210,N_20267);
and U21785 (N_21785,N_20893,N_20660);
and U21786 (N_21786,N_20487,N_20100);
xnor U21787 (N_21787,N_20863,N_20673);
or U21788 (N_21788,N_20899,N_20747);
xor U21789 (N_21789,N_20249,N_20189);
nor U21790 (N_21790,N_20986,N_20180);
and U21791 (N_21791,N_20343,N_20361);
nand U21792 (N_21792,N_20682,N_20561);
or U21793 (N_21793,N_20521,N_20868);
nand U21794 (N_21794,N_20005,N_20391);
and U21795 (N_21795,N_20647,N_20431);
nor U21796 (N_21796,N_20315,N_20763);
xor U21797 (N_21797,N_20845,N_20529);
nor U21798 (N_21798,N_20557,N_20957);
nand U21799 (N_21799,N_20470,N_20435);
nand U21800 (N_21800,N_20467,N_20164);
and U21801 (N_21801,N_20412,N_20780);
nand U21802 (N_21802,N_20492,N_20413);
nor U21803 (N_21803,N_20750,N_20223);
xor U21804 (N_21804,N_20355,N_20301);
xor U21805 (N_21805,N_20091,N_20990);
nor U21806 (N_21806,N_20448,N_20096);
nor U21807 (N_21807,N_20927,N_20131);
nand U21808 (N_21808,N_20277,N_20324);
and U21809 (N_21809,N_20377,N_20655);
nor U21810 (N_21810,N_20924,N_20003);
nor U21811 (N_21811,N_20280,N_20840);
nor U21812 (N_21812,N_20929,N_20597);
nand U21813 (N_21813,N_20128,N_20592);
xnor U21814 (N_21814,N_20030,N_20649);
xnor U21815 (N_21815,N_20612,N_20218);
and U21816 (N_21816,N_20367,N_20871);
xnor U21817 (N_21817,N_20902,N_20672);
xor U21818 (N_21818,N_20793,N_20697);
nand U21819 (N_21819,N_20466,N_20294);
xor U21820 (N_21820,N_20182,N_20223);
nand U21821 (N_21821,N_20494,N_20871);
nand U21822 (N_21822,N_20635,N_20977);
xor U21823 (N_21823,N_20537,N_20341);
xnor U21824 (N_21824,N_20943,N_20496);
nand U21825 (N_21825,N_20956,N_20110);
and U21826 (N_21826,N_20024,N_20065);
and U21827 (N_21827,N_20714,N_20260);
and U21828 (N_21828,N_20867,N_20640);
xor U21829 (N_21829,N_20662,N_20511);
xnor U21830 (N_21830,N_20301,N_20350);
xnor U21831 (N_21831,N_20951,N_20430);
or U21832 (N_21832,N_20687,N_20689);
nor U21833 (N_21833,N_20626,N_20773);
or U21834 (N_21834,N_20037,N_20334);
nand U21835 (N_21835,N_20131,N_20044);
nand U21836 (N_21836,N_20239,N_20423);
xnor U21837 (N_21837,N_20522,N_20401);
and U21838 (N_21838,N_20615,N_20576);
nand U21839 (N_21839,N_20079,N_20814);
nor U21840 (N_21840,N_20780,N_20505);
xor U21841 (N_21841,N_20745,N_20158);
or U21842 (N_21842,N_20948,N_20532);
and U21843 (N_21843,N_20698,N_20382);
nor U21844 (N_21844,N_20796,N_20997);
nand U21845 (N_21845,N_20119,N_20752);
and U21846 (N_21846,N_20314,N_20517);
nand U21847 (N_21847,N_20713,N_20518);
or U21848 (N_21848,N_20221,N_20549);
and U21849 (N_21849,N_20130,N_20734);
nand U21850 (N_21850,N_20020,N_20063);
nand U21851 (N_21851,N_20180,N_20772);
xor U21852 (N_21852,N_20581,N_20907);
xnor U21853 (N_21853,N_20758,N_20972);
or U21854 (N_21854,N_20327,N_20863);
or U21855 (N_21855,N_20978,N_20256);
nand U21856 (N_21856,N_20912,N_20435);
xor U21857 (N_21857,N_20861,N_20133);
and U21858 (N_21858,N_20471,N_20328);
nor U21859 (N_21859,N_20880,N_20008);
xnor U21860 (N_21860,N_20397,N_20619);
nand U21861 (N_21861,N_20355,N_20058);
nor U21862 (N_21862,N_20552,N_20082);
xor U21863 (N_21863,N_20146,N_20813);
or U21864 (N_21864,N_20681,N_20769);
nor U21865 (N_21865,N_20831,N_20040);
or U21866 (N_21866,N_20490,N_20688);
or U21867 (N_21867,N_20569,N_20101);
and U21868 (N_21868,N_20980,N_20378);
or U21869 (N_21869,N_20110,N_20615);
and U21870 (N_21870,N_20721,N_20190);
and U21871 (N_21871,N_20672,N_20727);
and U21872 (N_21872,N_20066,N_20444);
and U21873 (N_21873,N_20055,N_20599);
and U21874 (N_21874,N_20127,N_20841);
nor U21875 (N_21875,N_20280,N_20621);
and U21876 (N_21876,N_20764,N_20472);
nor U21877 (N_21877,N_20300,N_20365);
nand U21878 (N_21878,N_20994,N_20881);
or U21879 (N_21879,N_20499,N_20579);
and U21880 (N_21880,N_20966,N_20237);
nor U21881 (N_21881,N_20744,N_20903);
nor U21882 (N_21882,N_20715,N_20282);
and U21883 (N_21883,N_20635,N_20541);
nand U21884 (N_21884,N_20968,N_20089);
nor U21885 (N_21885,N_20061,N_20221);
xor U21886 (N_21886,N_20106,N_20223);
nand U21887 (N_21887,N_20014,N_20435);
and U21888 (N_21888,N_20226,N_20915);
and U21889 (N_21889,N_20112,N_20706);
xnor U21890 (N_21890,N_20974,N_20469);
nor U21891 (N_21891,N_20387,N_20524);
xor U21892 (N_21892,N_20950,N_20583);
or U21893 (N_21893,N_20805,N_20382);
and U21894 (N_21894,N_20389,N_20135);
and U21895 (N_21895,N_20962,N_20669);
nor U21896 (N_21896,N_20225,N_20305);
nor U21897 (N_21897,N_20187,N_20801);
or U21898 (N_21898,N_20419,N_20673);
nand U21899 (N_21899,N_20721,N_20364);
or U21900 (N_21900,N_20880,N_20783);
xnor U21901 (N_21901,N_20876,N_20051);
and U21902 (N_21902,N_20213,N_20204);
nor U21903 (N_21903,N_20899,N_20970);
nor U21904 (N_21904,N_20401,N_20634);
nand U21905 (N_21905,N_20919,N_20690);
and U21906 (N_21906,N_20889,N_20012);
xor U21907 (N_21907,N_20644,N_20957);
xor U21908 (N_21908,N_20528,N_20886);
nand U21909 (N_21909,N_20549,N_20601);
nor U21910 (N_21910,N_20653,N_20275);
or U21911 (N_21911,N_20659,N_20935);
nor U21912 (N_21912,N_20849,N_20840);
nand U21913 (N_21913,N_20599,N_20018);
nand U21914 (N_21914,N_20902,N_20839);
xor U21915 (N_21915,N_20128,N_20078);
and U21916 (N_21916,N_20567,N_20322);
or U21917 (N_21917,N_20739,N_20617);
and U21918 (N_21918,N_20019,N_20737);
nor U21919 (N_21919,N_20318,N_20914);
xnor U21920 (N_21920,N_20418,N_20914);
or U21921 (N_21921,N_20851,N_20472);
and U21922 (N_21922,N_20114,N_20197);
nor U21923 (N_21923,N_20118,N_20968);
nor U21924 (N_21924,N_20711,N_20134);
or U21925 (N_21925,N_20928,N_20807);
nand U21926 (N_21926,N_20045,N_20663);
nor U21927 (N_21927,N_20001,N_20426);
and U21928 (N_21928,N_20710,N_20178);
nand U21929 (N_21929,N_20110,N_20601);
xor U21930 (N_21930,N_20343,N_20910);
xor U21931 (N_21931,N_20131,N_20313);
nor U21932 (N_21932,N_20107,N_20522);
nor U21933 (N_21933,N_20091,N_20344);
nor U21934 (N_21934,N_20023,N_20812);
xnor U21935 (N_21935,N_20047,N_20413);
xor U21936 (N_21936,N_20819,N_20095);
nand U21937 (N_21937,N_20337,N_20234);
nand U21938 (N_21938,N_20795,N_20896);
and U21939 (N_21939,N_20933,N_20231);
and U21940 (N_21940,N_20732,N_20402);
or U21941 (N_21941,N_20441,N_20100);
nor U21942 (N_21942,N_20122,N_20720);
or U21943 (N_21943,N_20439,N_20866);
nor U21944 (N_21944,N_20544,N_20614);
nand U21945 (N_21945,N_20912,N_20257);
xnor U21946 (N_21946,N_20690,N_20481);
nand U21947 (N_21947,N_20890,N_20698);
xnor U21948 (N_21948,N_20206,N_20946);
xor U21949 (N_21949,N_20299,N_20723);
nand U21950 (N_21950,N_20184,N_20278);
nand U21951 (N_21951,N_20506,N_20938);
xnor U21952 (N_21952,N_20347,N_20264);
or U21953 (N_21953,N_20935,N_20102);
nor U21954 (N_21954,N_20440,N_20805);
nand U21955 (N_21955,N_20639,N_20735);
xnor U21956 (N_21956,N_20177,N_20267);
nor U21957 (N_21957,N_20324,N_20551);
nand U21958 (N_21958,N_20377,N_20452);
nand U21959 (N_21959,N_20940,N_20725);
or U21960 (N_21960,N_20691,N_20249);
and U21961 (N_21961,N_20564,N_20231);
and U21962 (N_21962,N_20332,N_20479);
nor U21963 (N_21963,N_20212,N_20773);
or U21964 (N_21964,N_20807,N_20506);
and U21965 (N_21965,N_20079,N_20284);
or U21966 (N_21966,N_20983,N_20852);
xnor U21967 (N_21967,N_20738,N_20336);
and U21968 (N_21968,N_20777,N_20357);
nor U21969 (N_21969,N_20244,N_20834);
and U21970 (N_21970,N_20799,N_20981);
nand U21971 (N_21971,N_20041,N_20786);
and U21972 (N_21972,N_20137,N_20862);
and U21973 (N_21973,N_20568,N_20725);
and U21974 (N_21974,N_20860,N_20168);
xor U21975 (N_21975,N_20981,N_20454);
xor U21976 (N_21976,N_20493,N_20231);
nor U21977 (N_21977,N_20977,N_20667);
and U21978 (N_21978,N_20472,N_20738);
and U21979 (N_21979,N_20880,N_20258);
nand U21980 (N_21980,N_20681,N_20353);
and U21981 (N_21981,N_20809,N_20504);
or U21982 (N_21982,N_20169,N_20931);
or U21983 (N_21983,N_20971,N_20451);
and U21984 (N_21984,N_20140,N_20971);
nand U21985 (N_21985,N_20917,N_20035);
nor U21986 (N_21986,N_20739,N_20415);
and U21987 (N_21987,N_20442,N_20081);
or U21988 (N_21988,N_20315,N_20140);
and U21989 (N_21989,N_20061,N_20038);
and U21990 (N_21990,N_20441,N_20899);
xor U21991 (N_21991,N_20985,N_20864);
and U21992 (N_21992,N_20657,N_20565);
xnor U21993 (N_21993,N_20169,N_20708);
nand U21994 (N_21994,N_20017,N_20907);
and U21995 (N_21995,N_20103,N_20192);
and U21996 (N_21996,N_20210,N_20699);
xnor U21997 (N_21997,N_20467,N_20371);
and U21998 (N_21998,N_20218,N_20549);
xnor U21999 (N_21999,N_20204,N_20852);
and U22000 (N_22000,N_21143,N_21388);
xor U22001 (N_22001,N_21080,N_21943);
xnor U22002 (N_22002,N_21269,N_21376);
or U22003 (N_22003,N_21937,N_21239);
xnor U22004 (N_22004,N_21132,N_21825);
nor U22005 (N_22005,N_21791,N_21312);
nand U22006 (N_22006,N_21433,N_21886);
nand U22007 (N_22007,N_21467,N_21168);
nor U22008 (N_22008,N_21698,N_21370);
nor U22009 (N_22009,N_21008,N_21754);
or U22010 (N_22010,N_21578,N_21461);
nor U22011 (N_22011,N_21834,N_21498);
nand U22012 (N_22012,N_21667,N_21592);
xor U22013 (N_22013,N_21776,N_21528);
xnor U22014 (N_22014,N_21518,N_21377);
xor U22015 (N_22015,N_21456,N_21959);
nor U22016 (N_22016,N_21669,N_21551);
or U22017 (N_22017,N_21867,N_21476);
xor U22018 (N_22018,N_21585,N_21733);
xor U22019 (N_22019,N_21182,N_21349);
nand U22020 (N_22020,N_21052,N_21661);
xnor U22021 (N_22021,N_21728,N_21738);
nor U22022 (N_22022,N_21965,N_21473);
nor U22023 (N_22023,N_21193,N_21732);
xnor U22024 (N_22024,N_21119,N_21209);
nor U22025 (N_22025,N_21262,N_21236);
and U22026 (N_22026,N_21093,N_21400);
nor U22027 (N_22027,N_21992,N_21548);
nand U22028 (N_22028,N_21997,N_21336);
nor U22029 (N_22029,N_21729,N_21862);
nand U22030 (N_22030,N_21536,N_21246);
or U22031 (N_22031,N_21833,N_21594);
or U22032 (N_22032,N_21169,N_21748);
and U22033 (N_22033,N_21599,N_21197);
nand U22034 (N_22034,N_21465,N_21383);
xor U22035 (N_22035,N_21247,N_21180);
xnor U22036 (N_22036,N_21295,N_21385);
or U22037 (N_22037,N_21141,N_21437);
nor U22038 (N_22038,N_21410,N_21413);
nor U22039 (N_22039,N_21703,N_21151);
nor U22040 (N_22040,N_21402,N_21251);
nor U22041 (N_22041,N_21106,N_21011);
nand U22042 (N_22042,N_21572,N_21057);
nand U22043 (N_22043,N_21898,N_21082);
or U22044 (N_22044,N_21184,N_21617);
nand U22045 (N_22045,N_21705,N_21042);
or U22046 (N_22046,N_21186,N_21596);
and U22047 (N_22047,N_21475,N_21775);
and U22048 (N_22048,N_21555,N_21190);
xnor U22049 (N_22049,N_21021,N_21665);
xor U22050 (N_22050,N_21774,N_21484);
nor U22051 (N_22051,N_21897,N_21286);
and U22052 (N_22052,N_21065,N_21921);
and U22053 (N_22053,N_21205,N_21519);
xnor U22054 (N_22054,N_21229,N_21894);
and U22055 (N_22055,N_21208,N_21660);
xnor U22056 (N_22056,N_21164,N_21706);
nand U22057 (N_22057,N_21242,N_21238);
and U22058 (N_22058,N_21017,N_21502);
nor U22059 (N_22059,N_21369,N_21772);
nand U22060 (N_22060,N_21367,N_21496);
nand U22061 (N_22061,N_21787,N_21558);
and U22062 (N_22062,N_21541,N_21328);
nor U22063 (N_22063,N_21326,N_21780);
and U22064 (N_22064,N_21167,N_21102);
nand U22065 (N_22065,N_21888,N_21582);
or U22066 (N_22066,N_21575,N_21986);
nand U22067 (N_22067,N_21321,N_21958);
nand U22068 (N_22068,N_21770,N_21796);
and U22069 (N_22069,N_21855,N_21292);
or U22070 (N_22070,N_21671,N_21882);
or U22071 (N_22071,N_21063,N_21913);
nand U22072 (N_22072,N_21195,N_21991);
xnor U22073 (N_22073,N_21023,N_21302);
or U22074 (N_22074,N_21024,N_21391);
xor U22075 (N_22075,N_21490,N_21830);
nand U22076 (N_22076,N_21911,N_21972);
nor U22077 (N_22077,N_21131,N_21634);
or U22078 (N_22078,N_21347,N_21676);
nand U22079 (N_22079,N_21712,N_21944);
xor U22080 (N_22080,N_21068,N_21957);
nor U22081 (N_22081,N_21823,N_21228);
nand U22082 (N_22082,N_21926,N_21115);
nand U22083 (N_22083,N_21511,N_21241);
and U22084 (N_22084,N_21268,N_21222);
nand U22085 (N_22085,N_21560,N_21171);
nor U22086 (N_22086,N_21896,N_21590);
or U22087 (N_22087,N_21727,N_21824);
xnor U22088 (N_22088,N_21666,N_21828);
and U22089 (N_22089,N_21808,N_21633);
nor U22090 (N_22090,N_21346,N_21296);
or U22091 (N_22091,N_21627,N_21015);
xor U22092 (N_22092,N_21371,N_21931);
nor U22093 (N_22093,N_21993,N_21577);
and U22094 (N_22094,N_21084,N_21081);
or U22095 (N_22095,N_21917,N_21569);
xor U22096 (N_22096,N_21799,N_21652);
or U22097 (N_22097,N_21954,N_21053);
xor U22098 (N_22098,N_21146,N_21883);
or U22099 (N_22099,N_21338,N_21134);
and U22100 (N_22100,N_21651,N_21538);
nor U22101 (N_22101,N_21317,N_21275);
xor U22102 (N_22102,N_21087,N_21688);
nand U22103 (N_22103,N_21013,N_21135);
nand U22104 (N_22104,N_21203,N_21805);
nor U22105 (N_22105,N_21500,N_21062);
xor U22106 (N_22106,N_21276,N_21000);
nand U22107 (N_22107,N_21645,N_21263);
nor U22108 (N_22108,N_21429,N_21014);
nand U22109 (N_22109,N_21827,N_21060);
or U22110 (N_22110,N_21010,N_21755);
or U22111 (N_22111,N_21220,N_21891);
xnor U22112 (N_22112,N_21147,N_21604);
and U22113 (N_22113,N_21544,N_21851);
or U22114 (N_22114,N_21339,N_21140);
xor U22115 (N_22115,N_21534,N_21924);
nand U22116 (N_22116,N_21202,N_21985);
xnor U22117 (N_22117,N_21839,N_21743);
nor U22118 (N_22118,N_21201,N_21850);
and U22119 (N_22119,N_21468,N_21477);
and U22120 (N_22120,N_21818,N_21207);
and U22121 (N_22121,N_21393,N_21005);
nand U22122 (N_22122,N_21861,N_21157);
nor U22123 (N_22123,N_21978,N_21411);
nor U22124 (N_22124,N_21460,N_21756);
or U22125 (N_22125,N_21587,N_21749);
and U22126 (N_22126,N_21443,N_21282);
xnor U22127 (N_22127,N_21160,N_21422);
or U22128 (N_22128,N_21724,N_21392);
xnor U22129 (N_22129,N_21952,N_21844);
nand U22130 (N_22130,N_21876,N_21056);
nor U22131 (N_22131,N_21904,N_21387);
nor U22132 (N_22132,N_21407,N_21932);
nor U22133 (N_22133,N_21381,N_21409);
xnor U22134 (N_22134,N_21524,N_21319);
xnor U22135 (N_22135,N_21192,N_21542);
nand U22136 (N_22136,N_21230,N_21900);
nor U22137 (N_22137,N_21880,N_21103);
nor U22138 (N_22138,N_21107,N_21826);
xor U22139 (N_22139,N_21591,N_21557);
and U22140 (N_22140,N_21936,N_21785);
and U22141 (N_22141,N_21117,N_21778);
nor U22142 (N_22142,N_21923,N_21089);
or U22143 (N_22143,N_21514,N_21097);
xnor U22144 (N_22144,N_21974,N_21231);
nand U22145 (N_22145,N_21289,N_21967);
or U22146 (N_22146,N_21664,N_21116);
and U22147 (N_22147,N_21811,N_21970);
nand U22148 (N_22148,N_21311,N_21323);
and U22149 (N_22149,N_21304,N_21104);
or U22150 (N_22150,N_21996,N_21085);
nor U22151 (N_22151,N_21687,N_21139);
nor U22152 (N_22152,N_21836,N_21976);
or U22153 (N_22153,N_21270,N_21709);
nand U22154 (N_22154,N_21865,N_21875);
or U22155 (N_22155,N_21176,N_21330);
and U22156 (N_22156,N_21074,N_21254);
nor U22157 (N_22157,N_21200,N_21797);
and U22158 (N_22158,N_21105,N_21829);
xor U22159 (N_22159,N_21866,N_21945);
and U22160 (N_22160,N_21375,N_21722);
and U22161 (N_22161,N_21148,N_21939);
nor U22162 (N_22162,N_21279,N_21522);
xor U22163 (N_22163,N_21512,N_21988);
nand U22164 (N_22164,N_21055,N_21725);
nor U22165 (N_22165,N_21951,N_21962);
and U22166 (N_22166,N_21320,N_21977);
nand U22167 (N_22167,N_21675,N_21020);
or U22168 (N_22168,N_21981,N_21630);
nor U22169 (N_22169,N_21390,N_21767);
or U22170 (N_22170,N_21837,N_21415);
and U22171 (N_22171,N_21849,N_21601);
and U22172 (N_22172,N_21786,N_21650);
nor U22173 (N_22173,N_21646,N_21002);
or U22174 (N_22174,N_21573,N_21278);
xnor U22175 (N_22175,N_21421,N_21441);
nand U22176 (N_22176,N_21576,N_21354);
nor U22177 (N_22177,N_21293,N_21710);
and U22178 (N_22178,N_21966,N_21812);
or U22179 (N_22179,N_21636,N_21623);
xnor U22180 (N_22180,N_21804,N_21635);
and U22181 (N_22181,N_21740,N_21846);
and U22182 (N_22182,N_21234,N_21004);
nand U22183 (N_22183,N_21048,N_21449);
nand U22184 (N_22184,N_21277,N_21769);
nor U22185 (N_22185,N_21110,N_21533);
xor U22186 (N_22186,N_21737,N_21071);
nand U22187 (N_22187,N_21142,N_21768);
nand U22188 (N_22188,N_21123,N_21436);
xnor U22189 (N_22189,N_21120,N_21610);
xnor U22190 (N_22190,N_21758,N_21657);
and U22191 (N_22191,N_21508,N_21078);
nand U22192 (N_22192,N_21870,N_21424);
xor U22193 (N_22193,N_21495,N_21434);
nor U22194 (N_22194,N_21344,N_21588);
nand U22195 (N_22195,N_21579,N_21948);
nor U22196 (N_22196,N_21677,N_21452);
or U22197 (N_22197,N_21307,N_21294);
nand U22198 (N_22198,N_21674,N_21210);
or U22199 (N_22199,N_21649,N_21418);
nor U22200 (N_22200,N_21189,N_21835);
or U22201 (N_22201,N_21779,N_21406);
or U22202 (N_22202,N_21736,N_21919);
nor U22203 (N_22203,N_21419,N_21156);
nand U22204 (N_22204,N_21540,N_21260);
nand U22205 (N_22205,N_21771,N_21889);
nor U22206 (N_22206,N_21877,N_21154);
xor U22207 (N_22207,N_21290,N_21721);
nor U22208 (N_22208,N_21138,N_21642);
or U22209 (N_22209,N_21751,N_21485);
nor U22210 (N_22210,N_21285,N_21505);
xnor U22211 (N_22211,N_21715,N_21545);
xnor U22212 (N_22212,N_21856,N_21685);
nand U22213 (N_22213,N_21510,N_21194);
nor U22214 (N_22214,N_21953,N_21858);
xnor U22215 (N_22215,N_21343,N_21956);
nor U22216 (N_22216,N_21638,N_21412);
xnor U22217 (N_22217,N_21717,N_21427);
nand U22218 (N_22218,N_21655,N_21987);
nor U22219 (N_22219,N_21621,N_21032);
xor U22220 (N_22220,N_21204,N_21982);
and U22221 (N_22221,N_21380,N_21172);
nand U22222 (N_22222,N_21702,N_21714);
nand U22223 (N_22223,N_21908,N_21860);
nor U22224 (N_22224,N_21525,N_21384);
xor U22225 (N_22225,N_21038,N_21893);
or U22226 (N_22226,N_21240,N_21414);
and U22227 (N_22227,N_21801,N_21611);
xor U22228 (N_22228,N_21223,N_21905);
nor U22229 (N_22229,N_21170,N_21403);
and U22230 (N_22230,N_21352,N_21644);
nor U22231 (N_22231,N_21704,N_21051);
and U22232 (N_22232,N_21798,N_21716);
or U22233 (N_22233,N_21348,N_21752);
nand U22234 (N_22234,N_21399,N_21521);
xor U22235 (N_22235,N_21361,N_21374);
nor U22236 (N_22236,N_21946,N_21784);
or U22237 (N_22237,N_21969,N_21094);
xnor U22238 (N_22238,N_21287,N_21155);
nand U22239 (N_22239,N_21187,N_21554);
xor U22240 (N_22240,N_21373,N_21067);
or U22241 (N_22241,N_21450,N_21859);
nor U22242 (N_22242,N_21464,N_21252);
nor U22243 (N_22243,N_21793,N_21726);
xnor U22244 (N_22244,N_21907,N_21041);
and U22245 (N_22245,N_21095,N_21731);
and U22246 (N_22246,N_21358,N_21746);
xnor U22247 (N_22247,N_21628,N_21637);
nor U22248 (N_22248,N_21513,N_21895);
xor U22249 (N_22249,N_21906,N_21493);
and U22250 (N_22250,N_21274,N_21248);
xnor U22251 (N_22251,N_21090,N_21730);
and U22252 (N_22252,N_21874,N_21890);
and U22253 (N_22253,N_21009,N_21198);
xnor U22254 (N_22254,N_21077,N_21297);
nand U22255 (N_22255,N_21547,N_21757);
xor U22256 (N_22256,N_21149,N_21903);
nor U22257 (N_22257,N_21175,N_21763);
xnor U22258 (N_22258,N_21099,N_21044);
or U22259 (N_22259,N_21446,N_21941);
xor U22260 (N_22260,N_21451,N_21506);
and U22261 (N_22261,N_21947,N_21530);
or U22262 (N_22262,N_21955,N_21114);
xor U22263 (N_22263,N_21625,N_21158);
nand U22264 (N_22264,N_21700,N_21145);
xor U22265 (N_22265,N_21960,N_21491);
nand U22266 (N_22266,N_21631,N_21942);
or U22267 (N_22267,N_21852,N_21012);
xnor U22268 (N_22268,N_21999,N_21092);
xor U22269 (N_22269,N_21574,N_21998);
xor U22270 (N_22270,N_21076,N_21662);
nor U22271 (N_22271,N_21389,N_21790);
nand U22272 (N_22272,N_21603,N_21584);
and U22273 (N_22273,N_21217,N_21764);
xnor U22274 (N_22274,N_21532,N_21641);
nor U22275 (N_22275,N_21161,N_21912);
or U22276 (N_22276,N_21355,N_21118);
nor U22277 (N_22277,N_21291,N_21325);
xor U22278 (N_22278,N_21310,N_21759);
and U22279 (N_22279,N_21100,N_21884);
or U22280 (N_22280,N_21480,N_21341);
and U22281 (N_22281,N_21064,N_21741);
nand U22282 (N_22282,N_21929,N_21214);
and U22283 (N_22283,N_21360,N_21417);
nand U22284 (N_22284,N_21810,N_21892);
or U22285 (N_22285,N_21153,N_21938);
nand U22286 (N_22286,N_21257,N_21624);
nor U22287 (N_22287,N_21455,N_21219);
and U22288 (N_22288,N_21216,N_21045);
nor U22289 (N_22289,N_21620,N_21863);
or U22290 (N_22290,N_21233,N_21463);
nand U22291 (N_22291,N_21968,N_21280);
nand U22292 (N_22292,N_21237,N_21125);
or U22293 (N_22293,N_21487,N_21762);
nand U22294 (N_22294,N_21298,N_21678);
and U22295 (N_22295,N_21553,N_21128);
or U22296 (N_22296,N_21788,N_21813);
or U22297 (N_22297,N_21178,N_21918);
and U22298 (N_22298,N_21447,N_21520);
or U22299 (N_22299,N_21006,N_21211);
nor U22300 (N_22300,N_21322,N_21255);
nand U22301 (N_22301,N_21925,N_21261);
nand U22302 (N_22302,N_21423,N_21070);
nand U22303 (N_22303,N_21227,N_21300);
or U22304 (N_22304,N_21249,N_21781);
and U22305 (N_22305,N_21440,N_21308);
nand U22306 (N_22306,N_21007,N_21398);
or U22307 (N_22307,N_21382,N_21853);
or U22308 (N_22308,N_21137,N_21701);
nand U22309 (N_22309,N_21616,N_21359);
nor U22310 (N_22310,N_21183,N_21822);
nand U22311 (N_22311,N_21018,N_21689);
or U22312 (N_22312,N_21618,N_21609);
and U22313 (N_22313,N_21694,N_21699);
nand U22314 (N_22314,N_21225,N_21843);
and U22315 (N_22315,N_21165,N_21583);
nor U22316 (N_22316,N_21162,N_21831);
nor U22317 (N_22317,N_21035,N_21072);
nor U22318 (N_22318,N_21559,N_21975);
xnor U22319 (N_22319,N_21492,N_21619);
and U22320 (N_22320,N_21878,N_21615);
nor U22321 (N_22321,N_21288,N_21750);
nor U22322 (N_22322,N_21353,N_21306);
nor U22323 (N_22323,N_21848,N_21922);
xnor U22324 (N_22324,N_21656,N_21568);
xor U22325 (N_22325,N_21470,N_21691);
and U22326 (N_22326,N_21144,N_21571);
nand U22327 (N_22327,N_21679,N_21001);
nand U22328 (N_22328,N_21909,N_21163);
xnor U22329 (N_22329,N_21259,N_21486);
nor U22330 (N_22330,N_21901,N_21556);
xor U22331 (N_22331,N_21022,N_21567);
and U22332 (N_22332,N_21019,N_21129);
nor U22333 (N_22333,N_21283,N_21166);
or U22334 (N_22334,N_21562,N_21806);
nor U22335 (N_22335,N_21872,N_21516);
or U22336 (N_22336,N_21586,N_21854);
or U22337 (N_22337,N_21598,N_21819);
xnor U22338 (N_22338,N_21133,N_21504);
nand U22339 (N_22339,N_21364,N_21043);
nor U22340 (N_22340,N_21658,N_21066);
or U22341 (N_22341,N_21789,N_21356);
and U22342 (N_22342,N_21995,N_21916);
xor U22343 (N_22343,N_21408,N_21301);
nand U22344 (N_22344,N_21469,N_21821);
nor U22345 (N_22345,N_21994,N_21272);
nor U22346 (N_22346,N_21483,N_21054);
nor U22347 (N_22347,N_21037,N_21523);
or U22348 (N_22348,N_21466,N_21212);
or U22349 (N_22349,N_21478,N_21593);
or U22350 (N_22350,N_21928,N_21098);
or U22351 (N_22351,N_21159,N_21979);
nor U22352 (N_22352,N_21039,N_21177);
nand U22353 (N_22353,N_21765,N_21462);
or U22354 (N_22354,N_21529,N_21258);
or U22355 (N_22355,N_21885,N_21871);
nand U22356 (N_22356,N_21654,N_21096);
and U22357 (N_22357,N_21425,N_21535);
or U22358 (N_22358,N_21061,N_21807);
or U22359 (N_22359,N_21845,N_21648);
nand U22360 (N_22360,N_21949,N_21564);
and U22361 (N_22361,N_21331,N_21426);
and U22362 (N_22362,N_21842,N_21394);
and U22363 (N_22363,N_21264,N_21050);
or U22364 (N_22364,N_21152,N_21537);
nor U22365 (N_22365,N_21742,N_21397);
nand U22366 (N_22366,N_21179,N_21961);
or U22367 (N_22367,N_21267,N_21899);
nand U22368 (N_22368,N_21783,N_21036);
and U22369 (N_22369,N_21910,N_21747);
nand U22370 (N_22370,N_21494,N_21690);
and U22371 (N_22371,N_21329,N_21795);
xnor U22372 (N_22372,N_21029,N_21950);
and U22373 (N_22373,N_21073,N_21454);
nand U22374 (N_22374,N_21109,N_21570);
nor U22375 (N_22375,N_21471,N_21927);
or U22376 (N_22376,N_21316,N_21059);
xor U22377 (N_22377,N_21033,N_21809);
xnor U22378 (N_22378,N_21915,N_21218);
and U22379 (N_22379,N_21914,N_21430);
or U22380 (N_22380,N_21990,N_21315);
or U22381 (N_22381,N_21457,N_21028);
nor U22382 (N_22382,N_21543,N_21696);
nor U22383 (N_22383,N_21550,N_21711);
or U22384 (N_22384,N_21124,N_21682);
xor U22385 (N_22385,N_21340,N_21964);
nand U22386 (N_22386,N_21058,N_21777);
and U22387 (N_22387,N_21256,N_21265);
nor U22388 (N_22388,N_21047,N_21980);
nor U22389 (N_22389,N_21539,N_21313);
or U22390 (N_22390,N_21351,N_21253);
nor U22391 (N_22391,N_21196,N_21150);
xor U22392 (N_22392,N_21185,N_21920);
xor U22393 (N_22393,N_21489,N_21563);
nor U22394 (N_22394,N_21803,N_21744);
nand U22395 (N_22395,N_21049,N_21439);
xnor U22396 (N_22396,N_21459,N_21357);
xnor U22397 (N_22397,N_21707,N_21940);
nand U22398 (N_22398,N_21453,N_21820);
or U22399 (N_22399,N_21632,N_21111);
or U22400 (N_22400,N_21526,N_21531);
or U22401 (N_22401,N_21509,N_21416);
xor U22402 (N_22402,N_21873,N_21681);
nor U22403 (N_22403,N_21607,N_21552);
nand U22404 (N_22404,N_21378,N_21566);
xor U22405 (N_22405,N_21614,N_21841);
or U22406 (N_22406,N_21224,N_21342);
xnor U22407 (N_22407,N_21445,N_21792);
xor U22408 (N_22408,N_21130,N_21079);
nor U22409 (N_22409,N_21723,N_21363);
nand U22410 (N_22410,N_21814,N_21420);
nor U22411 (N_22411,N_21869,N_21695);
or U22412 (N_22412,N_21431,N_21581);
and U22413 (N_22413,N_21735,N_21602);
nand U22414 (N_22414,N_21622,N_21647);
nor U22415 (N_22415,N_21653,N_21474);
xor U22416 (N_22416,N_21515,N_21713);
and U22417 (N_22417,N_21739,N_21303);
or U22418 (N_22418,N_21503,N_21034);
or U22419 (N_22419,N_21745,N_21507);
nand U22420 (N_22420,N_21639,N_21173);
xnor U22421 (N_22421,N_21501,N_21626);
nor U22422 (N_22422,N_21040,N_21031);
nand U22423 (N_22423,N_21016,N_21395);
nand U22424 (N_22424,N_21472,N_21221);
nor U22425 (N_22425,N_21083,N_21499);
nand U22426 (N_22426,N_21335,N_21663);
xor U22427 (N_22427,N_21815,N_21327);
or U22428 (N_22428,N_21565,N_21840);
xnor U22429 (N_22429,N_21481,N_21332);
or U22430 (N_22430,N_21350,N_21314);
nor U22431 (N_22431,N_21232,N_21984);
nand U22432 (N_22432,N_21113,N_21086);
or U22433 (N_22433,N_21368,N_21324);
xor U22434 (N_22434,N_21435,N_21482);
nand U22435 (N_22435,N_21868,N_21091);
nor U22436 (N_22436,N_21213,N_21405);
or U22437 (N_22437,N_21206,N_21517);
and U22438 (N_22438,N_21718,N_21720);
xor U22439 (N_22439,N_21549,N_21546);
nand U22440 (N_22440,N_21686,N_21273);
or U22441 (N_22441,N_21235,N_21935);
xor U22442 (N_22442,N_21608,N_21643);
or U22443 (N_22443,N_21734,N_21112);
or U22444 (N_22444,N_21847,N_21448);
xor U22445 (N_22445,N_21428,N_21299);
nor U22446 (N_22446,N_21027,N_21127);
or U22447 (N_22447,N_21902,N_21281);
nand U22448 (N_22448,N_21692,N_21345);
xor U22449 (N_22449,N_21773,N_21934);
nor U22450 (N_22450,N_21613,N_21800);
or U22451 (N_22451,N_21881,N_21719);
xor U22452 (N_22452,N_21069,N_21761);
xnor U22453 (N_22453,N_21309,N_21673);
or U22454 (N_22454,N_21003,N_21561);
or U22455 (N_22455,N_21794,N_21226);
nor U22456 (N_22456,N_21030,N_21668);
xnor U22457 (N_22457,N_21753,N_21337);
and U22458 (N_22458,N_21659,N_21136);
nor U22459 (N_22459,N_21181,N_21887);
nand U22460 (N_22460,N_21802,N_21379);
xor U22461 (N_22461,N_21266,N_21488);
xnor U22462 (N_22462,N_21597,N_21075);
nand U22463 (N_22463,N_21188,N_21386);
or U22464 (N_22464,N_21589,N_21693);
nor U22465 (N_22465,N_21672,N_21670);
nand U22466 (N_22466,N_21817,N_21244);
or U22467 (N_22467,N_21963,N_21245);
xor U22468 (N_22468,N_21101,N_21365);
xor U22469 (N_22469,N_21046,N_21989);
nor U22470 (N_22470,N_21971,N_21606);
or U22471 (N_22471,N_21782,N_21527);
nand U22472 (N_22472,N_21366,N_21973);
nor U22473 (N_22473,N_21121,N_21318);
or U22474 (N_22474,N_21930,N_21479);
xnor U22475 (N_22475,N_21983,N_21580);
or U22476 (N_22476,N_21640,N_21088);
xnor U22477 (N_22477,N_21432,N_21497);
nor U22478 (N_22478,N_21444,N_21857);
nand U22479 (N_22479,N_21396,N_21438);
or U22480 (N_22480,N_21215,N_21372);
nor U22481 (N_22481,N_21864,N_21684);
nor U22482 (N_22482,N_21458,N_21174);
and U22483 (N_22483,N_21600,N_21879);
nand U22484 (N_22484,N_21816,N_21442);
nor U22485 (N_22485,N_21612,N_21832);
nor U22486 (N_22486,N_21191,N_21683);
and U22487 (N_22487,N_21025,N_21933);
nor U22488 (N_22488,N_21838,N_21250);
nand U22489 (N_22489,N_21404,N_21305);
nor U22490 (N_22490,N_21697,N_21284);
and U22491 (N_22491,N_21271,N_21333);
xnor U22492 (N_22492,N_21122,N_21605);
xnor U22493 (N_22493,N_21334,N_21766);
and U22494 (N_22494,N_21126,N_21199);
nor U22495 (N_22495,N_21108,N_21401);
and U22496 (N_22496,N_21708,N_21595);
and U22497 (N_22497,N_21680,N_21243);
or U22498 (N_22498,N_21026,N_21629);
nor U22499 (N_22499,N_21760,N_21362);
or U22500 (N_22500,N_21463,N_21989);
and U22501 (N_22501,N_21206,N_21083);
and U22502 (N_22502,N_21735,N_21399);
or U22503 (N_22503,N_21187,N_21178);
nor U22504 (N_22504,N_21113,N_21209);
nor U22505 (N_22505,N_21905,N_21605);
xnor U22506 (N_22506,N_21744,N_21191);
nand U22507 (N_22507,N_21683,N_21344);
nor U22508 (N_22508,N_21990,N_21514);
nor U22509 (N_22509,N_21100,N_21642);
or U22510 (N_22510,N_21945,N_21555);
xnor U22511 (N_22511,N_21849,N_21696);
or U22512 (N_22512,N_21158,N_21775);
and U22513 (N_22513,N_21829,N_21283);
xnor U22514 (N_22514,N_21144,N_21989);
xor U22515 (N_22515,N_21052,N_21709);
nor U22516 (N_22516,N_21517,N_21123);
nor U22517 (N_22517,N_21176,N_21350);
and U22518 (N_22518,N_21080,N_21362);
xnor U22519 (N_22519,N_21081,N_21972);
nor U22520 (N_22520,N_21602,N_21659);
or U22521 (N_22521,N_21386,N_21416);
nand U22522 (N_22522,N_21065,N_21199);
nand U22523 (N_22523,N_21070,N_21322);
nor U22524 (N_22524,N_21374,N_21703);
and U22525 (N_22525,N_21128,N_21954);
xnor U22526 (N_22526,N_21647,N_21630);
or U22527 (N_22527,N_21929,N_21932);
and U22528 (N_22528,N_21240,N_21231);
nor U22529 (N_22529,N_21009,N_21031);
and U22530 (N_22530,N_21209,N_21729);
nand U22531 (N_22531,N_21500,N_21010);
nor U22532 (N_22532,N_21926,N_21785);
and U22533 (N_22533,N_21531,N_21416);
nand U22534 (N_22534,N_21770,N_21435);
and U22535 (N_22535,N_21941,N_21545);
nor U22536 (N_22536,N_21691,N_21616);
and U22537 (N_22537,N_21451,N_21132);
nand U22538 (N_22538,N_21864,N_21253);
and U22539 (N_22539,N_21658,N_21753);
nor U22540 (N_22540,N_21929,N_21060);
or U22541 (N_22541,N_21918,N_21216);
nor U22542 (N_22542,N_21532,N_21197);
and U22543 (N_22543,N_21420,N_21256);
nor U22544 (N_22544,N_21635,N_21791);
and U22545 (N_22545,N_21981,N_21661);
xnor U22546 (N_22546,N_21405,N_21592);
xor U22547 (N_22547,N_21710,N_21307);
nor U22548 (N_22548,N_21401,N_21975);
and U22549 (N_22549,N_21209,N_21761);
xor U22550 (N_22550,N_21077,N_21458);
nor U22551 (N_22551,N_21175,N_21579);
and U22552 (N_22552,N_21762,N_21273);
nor U22553 (N_22553,N_21549,N_21828);
nor U22554 (N_22554,N_21011,N_21785);
nand U22555 (N_22555,N_21087,N_21665);
nor U22556 (N_22556,N_21865,N_21525);
and U22557 (N_22557,N_21489,N_21744);
nor U22558 (N_22558,N_21250,N_21138);
nor U22559 (N_22559,N_21845,N_21393);
xor U22560 (N_22560,N_21622,N_21795);
nand U22561 (N_22561,N_21545,N_21095);
or U22562 (N_22562,N_21920,N_21127);
and U22563 (N_22563,N_21894,N_21756);
and U22564 (N_22564,N_21743,N_21252);
nor U22565 (N_22565,N_21350,N_21686);
nor U22566 (N_22566,N_21828,N_21908);
and U22567 (N_22567,N_21599,N_21630);
or U22568 (N_22568,N_21861,N_21761);
xnor U22569 (N_22569,N_21944,N_21142);
and U22570 (N_22570,N_21140,N_21384);
nand U22571 (N_22571,N_21414,N_21931);
or U22572 (N_22572,N_21888,N_21482);
xnor U22573 (N_22573,N_21657,N_21545);
or U22574 (N_22574,N_21355,N_21838);
nor U22575 (N_22575,N_21979,N_21669);
nor U22576 (N_22576,N_21769,N_21305);
and U22577 (N_22577,N_21808,N_21181);
or U22578 (N_22578,N_21969,N_21016);
or U22579 (N_22579,N_21464,N_21519);
nand U22580 (N_22580,N_21471,N_21233);
or U22581 (N_22581,N_21219,N_21985);
and U22582 (N_22582,N_21499,N_21318);
nor U22583 (N_22583,N_21040,N_21216);
xor U22584 (N_22584,N_21822,N_21037);
nand U22585 (N_22585,N_21929,N_21495);
nand U22586 (N_22586,N_21078,N_21411);
and U22587 (N_22587,N_21225,N_21117);
xor U22588 (N_22588,N_21125,N_21872);
and U22589 (N_22589,N_21761,N_21681);
or U22590 (N_22590,N_21291,N_21840);
nor U22591 (N_22591,N_21920,N_21180);
nor U22592 (N_22592,N_21454,N_21149);
or U22593 (N_22593,N_21053,N_21598);
xnor U22594 (N_22594,N_21788,N_21518);
or U22595 (N_22595,N_21324,N_21818);
and U22596 (N_22596,N_21925,N_21294);
or U22597 (N_22597,N_21676,N_21897);
nand U22598 (N_22598,N_21471,N_21444);
or U22599 (N_22599,N_21406,N_21601);
nand U22600 (N_22600,N_21405,N_21870);
and U22601 (N_22601,N_21909,N_21898);
and U22602 (N_22602,N_21816,N_21175);
or U22603 (N_22603,N_21725,N_21037);
nand U22604 (N_22604,N_21757,N_21187);
xor U22605 (N_22605,N_21826,N_21883);
xor U22606 (N_22606,N_21128,N_21333);
and U22607 (N_22607,N_21942,N_21577);
nor U22608 (N_22608,N_21152,N_21130);
xor U22609 (N_22609,N_21161,N_21926);
nor U22610 (N_22610,N_21192,N_21677);
or U22611 (N_22611,N_21778,N_21688);
xor U22612 (N_22612,N_21170,N_21021);
nor U22613 (N_22613,N_21303,N_21973);
and U22614 (N_22614,N_21071,N_21899);
xnor U22615 (N_22615,N_21552,N_21850);
and U22616 (N_22616,N_21212,N_21326);
nand U22617 (N_22617,N_21019,N_21649);
or U22618 (N_22618,N_21001,N_21044);
and U22619 (N_22619,N_21611,N_21088);
nor U22620 (N_22620,N_21992,N_21970);
nor U22621 (N_22621,N_21753,N_21069);
nand U22622 (N_22622,N_21813,N_21599);
nand U22623 (N_22623,N_21136,N_21290);
xor U22624 (N_22624,N_21663,N_21403);
or U22625 (N_22625,N_21509,N_21719);
nand U22626 (N_22626,N_21899,N_21872);
nand U22627 (N_22627,N_21694,N_21835);
nor U22628 (N_22628,N_21247,N_21422);
or U22629 (N_22629,N_21203,N_21257);
and U22630 (N_22630,N_21710,N_21031);
xor U22631 (N_22631,N_21598,N_21525);
nor U22632 (N_22632,N_21340,N_21874);
nor U22633 (N_22633,N_21578,N_21481);
xnor U22634 (N_22634,N_21192,N_21553);
and U22635 (N_22635,N_21486,N_21374);
and U22636 (N_22636,N_21348,N_21020);
or U22637 (N_22637,N_21795,N_21873);
nor U22638 (N_22638,N_21813,N_21203);
nor U22639 (N_22639,N_21391,N_21249);
and U22640 (N_22640,N_21303,N_21150);
nand U22641 (N_22641,N_21193,N_21097);
and U22642 (N_22642,N_21520,N_21289);
and U22643 (N_22643,N_21761,N_21032);
and U22644 (N_22644,N_21858,N_21451);
nor U22645 (N_22645,N_21659,N_21075);
or U22646 (N_22646,N_21698,N_21431);
nor U22647 (N_22647,N_21071,N_21885);
or U22648 (N_22648,N_21612,N_21280);
and U22649 (N_22649,N_21919,N_21013);
nand U22650 (N_22650,N_21569,N_21850);
nand U22651 (N_22651,N_21047,N_21706);
or U22652 (N_22652,N_21040,N_21079);
xnor U22653 (N_22653,N_21974,N_21018);
nor U22654 (N_22654,N_21653,N_21602);
xor U22655 (N_22655,N_21815,N_21630);
nand U22656 (N_22656,N_21600,N_21073);
nor U22657 (N_22657,N_21124,N_21244);
or U22658 (N_22658,N_21678,N_21564);
or U22659 (N_22659,N_21132,N_21363);
nor U22660 (N_22660,N_21570,N_21210);
nor U22661 (N_22661,N_21100,N_21578);
or U22662 (N_22662,N_21447,N_21795);
nor U22663 (N_22663,N_21615,N_21723);
and U22664 (N_22664,N_21901,N_21649);
and U22665 (N_22665,N_21847,N_21123);
and U22666 (N_22666,N_21274,N_21404);
or U22667 (N_22667,N_21779,N_21987);
xor U22668 (N_22668,N_21937,N_21586);
xnor U22669 (N_22669,N_21762,N_21046);
nor U22670 (N_22670,N_21287,N_21868);
nand U22671 (N_22671,N_21894,N_21131);
nor U22672 (N_22672,N_21903,N_21116);
or U22673 (N_22673,N_21657,N_21757);
nor U22674 (N_22674,N_21238,N_21225);
xor U22675 (N_22675,N_21688,N_21854);
or U22676 (N_22676,N_21924,N_21280);
nand U22677 (N_22677,N_21863,N_21506);
nor U22678 (N_22678,N_21092,N_21715);
nor U22679 (N_22679,N_21046,N_21331);
xnor U22680 (N_22680,N_21606,N_21027);
nand U22681 (N_22681,N_21637,N_21390);
or U22682 (N_22682,N_21265,N_21618);
xnor U22683 (N_22683,N_21127,N_21618);
or U22684 (N_22684,N_21957,N_21496);
and U22685 (N_22685,N_21720,N_21137);
or U22686 (N_22686,N_21723,N_21462);
nor U22687 (N_22687,N_21505,N_21855);
or U22688 (N_22688,N_21640,N_21183);
xor U22689 (N_22689,N_21213,N_21491);
or U22690 (N_22690,N_21531,N_21385);
xor U22691 (N_22691,N_21587,N_21055);
nand U22692 (N_22692,N_21449,N_21076);
nand U22693 (N_22693,N_21118,N_21324);
nand U22694 (N_22694,N_21084,N_21029);
and U22695 (N_22695,N_21023,N_21600);
or U22696 (N_22696,N_21979,N_21682);
nand U22697 (N_22697,N_21794,N_21428);
xor U22698 (N_22698,N_21410,N_21166);
xor U22699 (N_22699,N_21579,N_21913);
and U22700 (N_22700,N_21063,N_21313);
and U22701 (N_22701,N_21098,N_21277);
or U22702 (N_22702,N_21761,N_21956);
xor U22703 (N_22703,N_21693,N_21223);
nor U22704 (N_22704,N_21476,N_21890);
and U22705 (N_22705,N_21142,N_21542);
xnor U22706 (N_22706,N_21683,N_21428);
nor U22707 (N_22707,N_21494,N_21437);
xor U22708 (N_22708,N_21873,N_21156);
xor U22709 (N_22709,N_21983,N_21320);
nor U22710 (N_22710,N_21841,N_21608);
xnor U22711 (N_22711,N_21989,N_21441);
nand U22712 (N_22712,N_21006,N_21922);
or U22713 (N_22713,N_21234,N_21218);
and U22714 (N_22714,N_21500,N_21400);
and U22715 (N_22715,N_21776,N_21995);
xor U22716 (N_22716,N_21494,N_21415);
nand U22717 (N_22717,N_21650,N_21625);
nor U22718 (N_22718,N_21319,N_21454);
xor U22719 (N_22719,N_21658,N_21672);
xnor U22720 (N_22720,N_21592,N_21782);
nand U22721 (N_22721,N_21320,N_21621);
xor U22722 (N_22722,N_21513,N_21342);
and U22723 (N_22723,N_21062,N_21692);
nor U22724 (N_22724,N_21600,N_21434);
and U22725 (N_22725,N_21648,N_21350);
nand U22726 (N_22726,N_21951,N_21028);
xor U22727 (N_22727,N_21537,N_21495);
nor U22728 (N_22728,N_21334,N_21072);
and U22729 (N_22729,N_21872,N_21717);
nor U22730 (N_22730,N_21890,N_21767);
nand U22731 (N_22731,N_21755,N_21322);
or U22732 (N_22732,N_21159,N_21374);
nor U22733 (N_22733,N_21544,N_21885);
and U22734 (N_22734,N_21884,N_21403);
nor U22735 (N_22735,N_21939,N_21157);
xor U22736 (N_22736,N_21003,N_21231);
xor U22737 (N_22737,N_21062,N_21461);
nand U22738 (N_22738,N_21319,N_21114);
xnor U22739 (N_22739,N_21961,N_21934);
nor U22740 (N_22740,N_21595,N_21310);
and U22741 (N_22741,N_21573,N_21087);
nor U22742 (N_22742,N_21163,N_21676);
or U22743 (N_22743,N_21293,N_21956);
nand U22744 (N_22744,N_21545,N_21788);
and U22745 (N_22745,N_21740,N_21419);
and U22746 (N_22746,N_21646,N_21756);
nor U22747 (N_22747,N_21336,N_21610);
xor U22748 (N_22748,N_21067,N_21849);
and U22749 (N_22749,N_21241,N_21751);
or U22750 (N_22750,N_21627,N_21418);
nor U22751 (N_22751,N_21601,N_21326);
xnor U22752 (N_22752,N_21510,N_21448);
nor U22753 (N_22753,N_21223,N_21446);
nand U22754 (N_22754,N_21979,N_21021);
nand U22755 (N_22755,N_21582,N_21529);
nor U22756 (N_22756,N_21944,N_21632);
nor U22757 (N_22757,N_21976,N_21684);
xnor U22758 (N_22758,N_21836,N_21489);
nand U22759 (N_22759,N_21115,N_21451);
or U22760 (N_22760,N_21033,N_21268);
xor U22761 (N_22761,N_21164,N_21865);
nand U22762 (N_22762,N_21208,N_21830);
nor U22763 (N_22763,N_21555,N_21906);
and U22764 (N_22764,N_21151,N_21706);
and U22765 (N_22765,N_21829,N_21217);
and U22766 (N_22766,N_21737,N_21578);
nand U22767 (N_22767,N_21949,N_21170);
nand U22768 (N_22768,N_21153,N_21214);
nor U22769 (N_22769,N_21211,N_21566);
nor U22770 (N_22770,N_21371,N_21112);
nor U22771 (N_22771,N_21443,N_21566);
or U22772 (N_22772,N_21260,N_21672);
nand U22773 (N_22773,N_21455,N_21064);
or U22774 (N_22774,N_21705,N_21826);
or U22775 (N_22775,N_21573,N_21008);
and U22776 (N_22776,N_21275,N_21471);
nor U22777 (N_22777,N_21408,N_21566);
and U22778 (N_22778,N_21374,N_21840);
xnor U22779 (N_22779,N_21334,N_21025);
nor U22780 (N_22780,N_21757,N_21067);
nand U22781 (N_22781,N_21342,N_21732);
nand U22782 (N_22782,N_21556,N_21981);
xor U22783 (N_22783,N_21913,N_21015);
xor U22784 (N_22784,N_21683,N_21698);
and U22785 (N_22785,N_21253,N_21829);
nand U22786 (N_22786,N_21947,N_21936);
xor U22787 (N_22787,N_21023,N_21701);
and U22788 (N_22788,N_21261,N_21219);
and U22789 (N_22789,N_21176,N_21780);
nor U22790 (N_22790,N_21567,N_21644);
nand U22791 (N_22791,N_21874,N_21831);
and U22792 (N_22792,N_21734,N_21993);
and U22793 (N_22793,N_21746,N_21714);
nor U22794 (N_22794,N_21514,N_21411);
and U22795 (N_22795,N_21180,N_21578);
nand U22796 (N_22796,N_21586,N_21912);
nand U22797 (N_22797,N_21365,N_21081);
and U22798 (N_22798,N_21428,N_21365);
xor U22799 (N_22799,N_21289,N_21791);
or U22800 (N_22800,N_21979,N_21378);
nor U22801 (N_22801,N_21082,N_21357);
and U22802 (N_22802,N_21277,N_21802);
nand U22803 (N_22803,N_21752,N_21804);
and U22804 (N_22804,N_21892,N_21817);
nand U22805 (N_22805,N_21252,N_21571);
nand U22806 (N_22806,N_21013,N_21759);
nor U22807 (N_22807,N_21697,N_21902);
xnor U22808 (N_22808,N_21095,N_21483);
and U22809 (N_22809,N_21176,N_21500);
xnor U22810 (N_22810,N_21631,N_21035);
xor U22811 (N_22811,N_21785,N_21579);
xor U22812 (N_22812,N_21191,N_21439);
nor U22813 (N_22813,N_21932,N_21226);
nand U22814 (N_22814,N_21988,N_21963);
nor U22815 (N_22815,N_21297,N_21458);
or U22816 (N_22816,N_21634,N_21020);
nand U22817 (N_22817,N_21866,N_21706);
nor U22818 (N_22818,N_21845,N_21025);
xnor U22819 (N_22819,N_21694,N_21345);
nor U22820 (N_22820,N_21725,N_21353);
and U22821 (N_22821,N_21775,N_21240);
nor U22822 (N_22822,N_21157,N_21752);
or U22823 (N_22823,N_21339,N_21416);
or U22824 (N_22824,N_21173,N_21821);
xor U22825 (N_22825,N_21843,N_21298);
xnor U22826 (N_22826,N_21392,N_21758);
xor U22827 (N_22827,N_21470,N_21457);
and U22828 (N_22828,N_21095,N_21580);
nand U22829 (N_22829,N_21371,N_21594);
or U22830 (N_22830,N_21014,N_21710);
and U22831 (N_22831,N_21733,N_21302);
or U22832 (N_22832,N_21184,N_21770);
nor U22833 (N_22833,N_21460,N_21784);
nor U22834 (N_22834,N_21382,N_21402);
nor U22835 (N_22835,N_21826,N_21422);
nor U22836 (N_22836,N_21102,N_21300);
nor U22837 (N_22837,N_21062,N_21379);
and U22838 (N_22838,N_21875,N_21166);
or U22839 (N_22839,N_21129,N_21626);
and U22840 (N_22840,N_21148,N_21972);
xor U22841 (N_22841,N_21113,N_21434);
nand U22842 (N_22842,N_21592,N_21251);
xnor U22843 (N_22843,N_21796,N_21503);
and U22844 (N_22844,N_21841,N_21920);
and U22845 (N_22845,N_21361,N_21003);
and U22846 (N_22846,N_21551,N_21437);
nand U22847 (N_22847,N_21730,N_21429);
xnor U22848 (N_22848,N_21514,N_21782);
or U22849 (N_22849,N_21490,N_21362);
nand U22850 (N_22850,N_21189,N_21278);
nand U22851 (N_22851,N_21428,N_21728);
or U22852 (N_22852,N_21138,N_21187);
nor U22853 (N_22853,N_21819,N_21558);
or U22854 (N_22854,N_21336,N_21579);
xor U22855 (N_22855,N_21678,N_21855);
nand U22856 (N_22856,N_21516,N_21446);
xnor U22857 (N_22857,N_21324,N_21799);
or U22858 (N_22858,N_21664,N_21726);
and U22859 (N_22859,N_21066,N_21165);
or U22860 (N_22860,N_21018,N_21074);
nor U22861 (N_22861,N_21866,N_21757);
and U22862 (N_22862,N_21133,N_21566);
or U22863 (N_22863,N_21202,N_21299);
xnor U22864 (N_22864,N_21822,N_21134);
xnor U22865 (N_22865,N_21955,N_21671);
nand U22866 (N_22866,N_21662,N_21752);
or U22867 (N_22867,N_21060,N_21151);
or U22868 (N_22868,N_21316,N_21491);
xor U22869 (N_22869,N_21522,N_21558);
or U22870 (N_22870,N_21407,N_21117);
nor U22871 (N_22871,N_21480,N_21828);
xnor U22872 (N_22872,N_21251,N_21097);
or U22873 (N_22873,N_21534,N_21397);
xnor U22874 (N_22874,N_21856,N_21786);
or U22875 (N_22875,N_21997,N_21327);
or U22876 (N_22876,N_21913,N_21094);
xnor U22877 (N_22877,N_21933,N_21722);
or U22878 (N_22878,N_21341,N_21659);
nor U22879 (N_22879,N_21515,N_21403);
nor U22880 (N_22880,N_21559,N_21449);
or U22881 (N_22881,N_21986,N_21593);
xnor U22882 (N_22882,N_21450,N_21539);
xnor U22883 (N_22883,N_21181,N_21474);
nand U22884 (N_22884,N_21240,N_21469);
and U22885 (N_22885,N_21327,N_21262);
nand U22886 (N_22886,N_21543,N_21159);
nor U22887 (N_22887,N_21011,N_21180);
nand U22888 (N_22888,N_21061,N_21996);
xor U22889 (N_22889,N_21043,N_21235);
xnor U22890 (N_22890,N_21267,N_21237);
nand U22891 (N_22891,N_21344,N_21167);
or U22892 (N_22892,N_21460,N_21973);
and U22893 (N_22893,N_21738,N_21355);
or U22894 (N_22894,N_21248,N_21837);
nor U22895 (N_22895,N_21439,N_21409);
xnor U22896 (N_22896,N_21553,N_21314);
xnor U22897 (N_22897,N_21241,N_21093);
xnor U22898 (N_22898,N_21880,N_21156);
nand U22899 (N_22899,N_21863,N_21046);
or U22900 (N_22900,N_21712,N_21389);
and U22901 (N_22901,N_21034,N_21602);
and U22902 (N_22902,N_21529,N_21177);
or U22903 (N_22903,N_21349,N_21620);
xnor U22904 (N_22904,N_21852,N_21266);
and U22905 (N_22905,N_21363,N_21468);
or U22906 (N_22906,N_21868,N_21347);
nand U22907 (N_22907,N_21861,N_21666);
xnor U22908 (N_22908,N_21358,N_21645);
nor U22909 (N_22909,N_21629,N_21624);
xor U22910 (N_22910,N_21146,N_21746);
or U22911 (N_22911,N_21239,N_21505);
nand U22912 (N_22912,N_21373,N_21759);
nor U22913 (N_22913,N_21990,N_21103);
xor U22914 (N_22914,N_21538,N_21070);
xnor U22915 (N_22915,N_21991,N_21389);
xor U22916 (N_22916,N_21692,N_21373);
xor U22917 (N_22917,N_21408,N_21413);
nor U22918 (N_22918,N_21289,N_21519);
nand U22919 (N_22919,N_21767,N_21478);
nor U22920 (N_22920,N_21793,N_21597);
and U22921 (N_22921,N_21107,N_21831);
nor U22922 (N_22922,N_21433,N_21510);
nand U22923 (N_22923,N_21785,N_21389);
and U22924 (N_22924,N_21130,N_21394);
and U22925 (N_22925,N_21389,N_21695);
or U22926 (N_22926,N_21183,N_21981);
nand U22927 (N_22927,N_21042,N_21608);
nand U22928 (N_22928,N_21036,N_21597);
and U22929 (N_22929,N_21537,N_21611);
xor U22930 (N_22930,N_21564,N_21887);
and U22931 (N_22931,N_21702,N_21067);
and U22932 (N_22932,N_21308,N_21564);
xnor U22933 (N_22933,N_21751,N_21418);
and U22934 (N_22934,N_21632,N_21369);
and U22935 (N_22935,N_21421,N_21144);
and U22936 (N_22936,N_21081,N_21022);
xor U22937 (N_22937,N_21905,N_21173);
xnor U22938 (N_22938,N_21112,N_21824);
nand U22939 (N_22939,N_21380,N_21539);
xor U22940 (N_22940,N_21508,N_21971);
nor U22941 (N_22941,N_21128,N_21457);
or U22942 (N_22942,N_21505,N_21829);
nor U22943 (N_22943,N_21049,N_21202);
or U22944 (N_22944,N_21571,N_21315);
and U22945 (N_22945,N_21515,N_21385);
or U22946 (N_22946,N_21662,N_21729);
and U22947 (N_22947,N_21345,N_21101);
or U22948 (N_22948,N_21790,N_21312);
or U22949 (N_22949,N_21751,N_21113);
xor U22950 (N_22950,N_21856,N_21009);
or U22951 (N_22951,N_21650,N_21511);
or U22952 (N_22952,N_21242,N_21198);
xor U22953 (N_22953,N_21912,N_21748);
nor U22954 (N_22954,N_21555,N_21491);
nor U22955 (N_22955,N_21325,N_21122);
nor U22956 (N_22956,N_21606,N_21345);
nand U22957 (N_22957,N_21185,N_21289);
xnor U22958 (N_22958,N_21720,N_21950);
nor U22959 (N_22959,N_21610,N_21570);
or U22960 (N_22960,N_21971,N_21747);
and U22961 (N_22961,N_21780,N_21019);
nor U22962 (N_22962,N_21840,N_21400);
nand U22963 (N_22963,N_21634,N_21990);
xnor U22964 (N_22964,N_21914,N_21350);
nand U22965 (N_22965,N_21869,N_21627);
or U22966 (N_22966,N_21688,N_21050);
xor U22967 (N_22967,N_21340,N_21440);
nor U22968 (N_22968,N_21414,N_21895);
or U22969 (N_22969,N_21598,N_21349);
and U22970 (N_22970,N_21248,N_21005);
xnor U22971 (N_22971,N_21644,N_21417);
xnor U22972 (N_22972,N_21476,N_21079);
nand U22973 (N_22973,N_21379,N_21165);
nand U22974 (N_22974,N_21625,N_21943);
or U22975 (N_22975,N_21097,N_21492);
xor U22976 (N_22976,N_21240,N_21791);
nor U22977 (N_22977,N_21850,N_21083);
or U22978 (N_22978,N_21899,N_21572);
and U22979 (N_22979,N_21632,N_21679);
nand U22980 (N_22980,N_21107,N_21225);
nand U22981 (N_22981,N_21830,N_21673);
nor U22982 (N_22982,N_21107,N_21905);
nand U22983 (N_22983,N_21662,N_21855);
xnor U22984 (N_22984,N_21796,N_21874);
xnor U22985 (N_22985,N_21647,N_21704);
nor U22986 (N_22986,N_21343,N_21213);
or U22987 (N_22987,N_21913,N_21174);
xor U22988 (N_22988,N_21981,N_21953);
or U22989 (N_22989,N_21768,N_21824);
and U22990 (N_22990,N_21489,N_21163);
and U22991 (N_22991,N_21195,N_21839);
and U22992 (N_22992,N_21441,N_21007);
nor U22993 (N_22993,N_21621,N_21967);
and U22994 (N_22994,N_21880,N_21436);
nor U22995 (N_22995,N_21030,N_21545);
nand U22996 (N_22996,N_21475,N_21391);
nor U22997 (N_22997,N_21390,N_21094);
nor U22998 (N_22998,N_21452,N_21208);
xnor U22999 (N_22999,N_21518,N_21497);
nand U23000 (N_23000,N_22196,N_22652);
nor U23001 (N_23001,N_22261,N_22761);
nor U23002 (N_23002,N_22368,N_22880);
nand U23003 (N_23003,N_22699,N_22840);
xnor U23004 (N_23004,N_22144,N_22541);
and U23005 (N_23005,N_22605,N_22602);
or U23006 (N_23006,N_22560,N_22948);
nand U23007 (N_23007,N_22414,N_22298);
or U23008 (N_23008,N_22394,N_22461);
nor U23009 (N_23009,N_22307,N_22143);
or U23010 (N_23010,N_22783,N_22807);
xnor U23011 (N_23011,N_22579,N_22906);
or U23012 (N_23012,N_22964,N_22272);
nand U23013 (N_23013,N_22611,N_22928);
or U23014 (N_23014,N_22572,N_22794);
or U23015 (N_23015,N_22996,N_22773);
and U23016 (N_23016,N_22811,N_22521);
xor U23017 (N_23017,N_22813,N_22289);
and U23018 (N_23018,N_22940,N_22241);
and U23019 (N_23019,N_22525,N_22121);
nand U23020 (N_23020,N_22963,N_22258);
xor U23021 (N_23021,N_22625,N_22573);
or U23022 (N_23022,N_22648,N_22918);
xnor U23023 (N_23023,N_22164,N_22956);
nand U23024 (N_23024,N_22567,N_22270);
nor U23025 (N_23025,N_22505,N_22748);
nand U23026 (N_23026,N_22279,N_22400);
or U23027 (N_23027,N_22549,N_22719);
and U23028 (N_23028,N_22716,N_22062);
nand U23029 (N_23029,N_22054,N_22574);
nand U23030 (N_23030,N_22018,N_22599);
or U23031 (N_23031,N_22077,N_22024);
xnor U23032 (N_23032,N_22836,N_22446);
and U23033 (N_23033,N_22325,N_22514);
or U23034 (N_23034,N_22950,N_22128);
nor U23035 (N_23035,N_22990,N_22337);
nand U23036 (N_23036,N_22027,N_22796);
xnor U23037 (N_23037,N_22684,N_22571);
nand U23038 (N_23038,N_22197,N_22189);
nand U23039 (N_23039,N_22775,N_22386);
nor U23040 (N_23040,N_22905,N_22326);
nor U23041 (N_23041,N_22925,N_22766);
nand U23042 (N_23042,N_22894,N_22510);
or U23043 (N_23043,N_22304,N_22531);
nor U23044 (N_23044,N_22967,N_22667);
nor U23045 (N_23045,N_22344,N_22971);
nand U23046 (N_23046,N_22445,N_22280);
and U23047 (N_23047,N_22937,N_22968);
nor U23048 (N_23048,N_22515,N_22127);
nand U23049 (N_23049,N_22009,N_22483);
xor U23050 (N_23050,N_22601,N_22010);
and U23051 (N_23051,N_22591,N_22491);
and U23052 (N_23052,N_22797,N_22868);
xnor U23053 (N_23053,N_22693,N_22388);
and U23054 (N_23054,N_22767,N_22629);
nor U23055 (N_23055,N_22608,N_22048);
nor U23056 (N_23056,N_22457,N_22268);
nor U23057 (N_23057,N_22607,N_22090);
nor U23058 (N_23058,N_22649,N_22429);
and U23059 (N_23059,N_22901,N_22323);
xor U23060 (N_23060,N_22259,N_22068);
nand U23061 (N_23061,N_22182,N_22743);
and U23062 (N_23062,N_22375,N_22839);
nor U23063 (N_23063,N_22355,N_22481);
or U23064 (N_23064,N_22665,N_22146);
or U23065 (N_23065,N_22785,N_22329);
or U23066 (N_23066,N_22348,N_22092);
and U23067 (N_23067,N_22387,N_22440);
xor U23068 (N_23068,N_22861,N_22660);
xnor U23069 (N_23069,N_22352,N_22626);
nand U23070 (N_23070,N_22857,N_22205);
xnor U23071 (N_23071,N_22341,N_22717);
and U23072 (N_23072,N_22338,N_22398);
xor U23073 (N_23073,N_22154,N_22247);
xnor U23074 (N_23074,N_22472,N_22933);
nand U23075 (N_23075,N_22040,N_22742);
nor U23076 (N_23076,N_22604,N_22022);
nor U23077 (N_23077,N_22673,N_22535);
xnor U23078 (N_23078,N_22911,N_22988);
nor U23079 (N_23079,N_22795,N_22297);
and U23080 (N_23080,N_22319,N_22218);
or U23081 (N_23081,N_22983,N_22370);
nand U23082 (N_23082,N_22830,N_22057);
and U23083 (N_23083,N_22480,N_22529);
or U23084 (N_23084,N_22885,N_22703);
nor U23085 (N_23085,N_22646,N_22255);
or U23086 (N_23086,N_22213,N_22035);
or U23087 (N_23087,N_22697,N_22228);
xnor U23088 (N_23088,N_22706,N_22428);
nor U23089 (N_23089,N_22635,N_22308);
nand U23090 (N_23090,N_22219,N_22876);
xnor U23091 (N_23091,N_22050,N_22680);
nand U23092 (N_23092,N_22416,N_22546);
nor U23093 (N_23093,N_22172,N_22423);
nor U23094 (N_23094,N_22603,N_22454);
nand U23095 (N_23095,N_22942,N_22181);
and U23096 (N_23096,N_22584,N_22257);
nand U23097 (N_23097,N_22818,N_22984);
nand U23098 (N_23098,N_22468,N_22449);
nor U23099 (N_23099,N_22793,N_22837);
nor U23100 (N_23100,N_22670,N_22808);
nand U23101 (N_23101,N_22866,N_22736);
and U23102 (N_23102,N_22185,N_22263);
nand U23103 (N_23103,N_22087,N_22526);
nand U23104 (N_23104,N_22558,N_22696);
nor U23105 (N_23105,N_22539,N_22425);
nand U23106 (N_23106,N_22582,N_22004);
and U23107 (N_23107,N_22506,N_22336);
xnor U23108 (N_23108,N_22407,N_22501);
nor U23109 (N_23109,N_22770,N_22522);
xnor U23110 (N_23110,N_22178,N_22730);
xor U23111 (N_23111,N_22354,N_22755);
nor U23112 (N_23112,N_22628,N_22765);
or U23113 (N_23113,N_22537,N_22170);
nor U23114 (N_23114,N_22473,N_22623);
or U23115 (N_23115,N_22191,N_22071);
xnor U23116 (N_23116,N_22664,N_22909);
nand U23117 (N_23117,N_22915,N_22007);
and U23118 (N_23118,N_22848,N_22311);
or U23119 (N_23119,N_22396,N_22187);
or U23120 (N_23120,N_22508,N_22202);
xor U23121 (N_23121,N_22484,N_22900);
xor U23122 (N_23122,N_22778,N_22944);
and U23123 (N_23123,N_22721,N_22466);
xnor U23124 (N_23124,N_22614,N_22576);
and U23125 (N_23125,N_22391,N_22493);
nand U23126 (N_23126,N_22036,N_22349);
xor U23127 (N_23127,N_22120,N_22681);
nand U23128 (N_23128,N_22978,N_22020);
nor U23129 (N_23129,N_22881,N_22300);
or U23130 (N_23130,N_22215,N_22212);
nor U23131 (N_23131,N_22932,N_22385);
and U23132 (N_23132,N_22923,N_22586);
and U23133 (N_23133,N_22869,N_22162);
or U23134 (N_23134,N_22408,N_22053);
nor U23135 (N_23135,N_22378,N_22816);
or U23136 (N_23136,N_22438,N_22158);
nand U23137 (N_23137,N_22874,N_22554);
nor U23138 (N_23138,N_22331,N_22698);
nor U23139 (N_23139,N_22093,N_22889);
or U23140 (N_23140,N_22126,N_22804);
nor U23141 (N_23141,N_22008,N_22318);
nor U23142 (N_23142,N_22758,N_22516);
or U23143 (N_23143,N_22823,N_22577);
nor U23144 (N_23144,N_22989,N_22662);
nand U23145 (N_23145,N_22015,N_22780);
or U23146 (N_23146,N_22553,N_22565);
nor U23147 (N_23147,N_22108,N_22913);
and U23148 (N_23148,N_22679,N_22924);
and U23149 (N_23149,N_22474,N_22455);
nand U23150 (N_23150,N_22957,N_22676);
nor U23151 (N_23151,N_22895,N_22105);
or U23152 (N_23152,N_22598,N_22262);
xnor U23153 (N_23153,N_22615,N_22760);
or U23154 (N_23154,N_22389,N_22225);
xnor U23155 (N_23155,N_22729,N_22772);
xnor U23156 (N_23156,N_22358,N_22738);
xnor U23157 (N_23157,N_22897,N_22168);
and U23158 (N_23158,N_22347,N_22754);
or U23159 (N_23159,N_22490,N_22283);
or U23160 (N_23160,N_22475,N_22882);
or U23161 (N_23161,N_22627,N_22477);
nor U23162 (N_23162,N_22070,N_22103);
nand U23163 (N_23163,N_22507,N_22829);
nand U23164 (N_23164,N_22444,N_22030);
or U23165 (N_23165,N_22412,N_22981);
nor U23166 (N_23166,N_22091,N_22327);
or U23167 (N_23167,N_22134,N_22700);
or U23168 (N_23168,N_22232,N_22183);
xnor U23169 (N_23169,N_22038,N_22528);
xor U23170 (N_23170,N_22992,N_22124);
nor U23171 (N_23171,N_22192,N_22275);
nor U23172 (N_23172,N_22805,N_22029);
and U23173 (N_23173,N_22421,N_22762);
or U23174 (N_23174,N_22339,N_22759);
or U23175 (N_23175,N_22059,N_22175);
and U23176 (N_23176,N_22860,N_22675);
and U23177 (N_23177,N_22756,N_22116);
and U23178 (N_23178,N_22273,N_22974);
nor U23179 (N_23179,N_22291,N_22418);
nand U23180 (N_23180,N_22141,N_22322);
and U23181 (N_23181,N_22788,N_22687);
and U23182 (N_23182,N_22100,N_22463);
or U23183 (N_23183,N_22089,N_22884);
nand U23184 (N_23184,N_22936,N_22301);
nor U23185 (N_23185,N_22372,N_22176);
and U23186 (N_23186,N_22668,N_22842);
and U23187 (N_23187,N_22306,N_22097);
nand U23188 (N_23188,N_22485,N_22589);
or U23189 (N_23189,N_22246,N_22953);
xnor U23190 (N_23190,N_22216,N_22744);
nand U23191 (N_23191,N_22530,N_22741);
nor U23192 (N_23192,N_22592,N_22982);
xnor U23193 (N_23193,N_22413,N_22986);
or U23194 (N_23194,N_22214,N_22952);
xnor U23195 (N_23195,N_22972,N_22286);
nand U23196 (N_23196,N_22732,N_22640);
nand U23197 (N_23197,N_22637,N_22065);
nand U23198 (N_23198,N_22343,N_22003);
or U23199 (N_23199,N_22624,N_22630);
nor U23200 (N_23200,N_22800,N_22207);
xor U23201 (N_23201,N_22471,N_22056);
and U23202 (N_23202,N_22922,N_22201);
nand U23203 (N_23203,N_22133,N_22271);
xnor U23204 (N_23204,N_22102,N_22538);
xnor U23205 (N_23205,N_22945,N_22487);
or U23206 (N_23206,N_22384,N_22217);
xor U23207 (N_23207,N_22689,N_22821);
xor U23208 (N_23208,N_22227,N_22877);
or U23209 (N_23209,N_22245,N_22991);
and U23210 (N_23210,N_22993,N_22055);
nor U23211 (N_23211,N_22998,N_22790);
or U23212 (N_23212,N_22424,N_22411);
and U23213 (N_23213,N_22317,N_22101);
or U23214 (N_23214,N_22976,N_22135);
and U23215 (N_23215,N_22465,N_22672);
nor U23216 (N_23216,N_22610,N_22067);
and U23217 (N_23217,N_22028,N_22570);
or U23218 (N_23218,N_22132,N_22504);
and U23219 (N_23219,N_22718,N_22557);
nand U23220 (N_23220,N_22432,N_22148);
or U23221 (N_23221,N_22113,N_22524);
or U23222 (N_23222,N_22137,N_22064);
nor U23223 (N_23223,N_22000,N_22498);
xnor U23224 (N_23224,N_22620,N_22791);
nand U23225 (N_23225,N_22237,N_22844);
xnor U23226 (N_23226,N_22859,N_22441);
or U23227 (N_23227,N_22360,N_22099);
nand U23228 (N_23228,N_22095,N_22476);
and U23229 (N_23229,N_22919,N_22434);
nand U23230 (N_23230,N_22583,N_22186);
nor U23231 (N_23231,N_22938,N_22887);
nand U23232 (N_23232,N_22392,N_22140);
nand U23233 (N_23233,N_22786,N_22633);
nor U23234 (N_23234,N_22084,N_22222);
xnor U23235 (N_23235,N_22220,N_22896);
or U23236 (N_23236,N_22208,N_22460);
xor U23237 (N_23237,N_22789,N_22031);
or U23238 (N_23238,N_22117,N_22824);
and U23239 (N_23239,N_22464,N_22403);
xnor U23240 (N_23240,N_22585,N_22858);
nand U23241 (N_23241,N_22488,N_22943);
and U23242 (N_23242,N_22588,N_22929);
and U23243 (N_23243,N_22230,N_22781);
nor U23244 (N_23244,N_22427,N_22578);
and U23245 (N_23245,N_22198,N_22006);
or U23246 (N_23246,N_22569,N_22452);
xor U23247 (N_23247,N_22899,N_22489);
nor U23248 (N_23248,N_22801,N_22155);
nand U23249 (N_23249,N_22890,N_22417);
nand U23250 (N_23250,N_22288,N_22459);
or U23251 (N_23251,N_22683,N_22935);
nor U23252 (N_23252,N_22616,N_22931);
nor U23253 (N_23253,N_22086,N_22921);
and U23254 (N_23254,N_22139,N_22244);
xnor U23255 (N_23255,N_22118,N_22907);
xnor U23256 (N_23256,N_22145,N_22688);
xor U23257 (N_23257,N_22934,N_22277);
nand U23258 (N_23258,N_22657,N_22152);
or U23259 (N_23259,N_22190,N_22013);
or U23260 (N_23260,N_22260,N_22156);
nor U23261 (N_23261,N_22835,N_22253);
nand U23262 (N_23262,N_22725,N_22774);
or U23263 (N_23263,N_22916,N_22194);
and U23264 (N_23264,N_22980,N_22511);
and U23265 (N_23265,N_22044,N_22720);
or U23266 (N_23266,N_22704,N_22771);
nor U23267 (N_23267,N_22871,N_22254);
xnor U23268 (N_23268,N_22757,N_22815);
or U23269 (N_23269,N_22619,N_22638);
or U23270 (N_23270,N_22551,N_22803);
nor U23271 (N_23271,N_22082,N_22290);
nor U23272 (N_23272,N_22238,N_22357);
nor U23273 (N_23273,N_22066,N_22157);
xor U23274 (N_23274,N_22659,N_22052);
nor U23275 (N_23275,N_22617,N_22831);
and U23276 (N_23276,N_22294,N_22677);
or U23277 (N_23277,N_22827,N_22987);
and U23278 (N_23278,N_22714,N_22305);
and U23279 (N_23279,N_22369,N_22872);
or U23280 (N_23280,N_22787,N_22397);
and U23281 (N_23281,N_22379,N_22726);
nand U23282 (N_23282,N_22692,N_22340);
and U23283 (N_23283,N_22431,N_22822);
and U23284 (N_23284,N_22927,N_22946);
nand U23285 (N_23285,N_22740,N_22912);
xor U23286 (N_23286,N_22960,N_22166);
nor U23287 (N_23287,N_22888,N_22041);
and U23288 (N_23288,N_22188,N_22975);
nor U23289 (N_23289,N_22123,N_22776);
nand U23290 (N_23290,N_22083,N_22310);
xnor U23291 (N_23291,N_22856,N_22076);
nor U23292 (N_23292,N_22722,N_22296);
and U23293 (N_23293,N_22845,N_22462);
xnor U23294 (N_23294,N_22406,N_22075);
xnor U23295 (N_23295,N_22647,N_22545);
xnor U23296 (N_23296,N_22174,N_22977);
nand U23297 (N_23297,N_22674,N_22798);
or U23298 (N_23298,N_22954,N_22025);
xor U23299 (N_23299,N_22321,N_22728);
and U23300 (N_23300,N_22994,N_22265);
and U23301 (N_23301,N_22594,N_22711);
nor U23302 (N_23302,N_22658,N_22021);
nor U23303 (N_23303,N_22229,N_22404);
or U23304 (N_23304,N_22512,N_22320);
and U23305 (N_23305,N_22303,N_22540);
nor U23306 (N_23306,N_22820,N_22346);
xnor U23307 (N_23307,N_22639,N_22151);
and U23308 (N_23308,N_22033,N_22383);
and U23309 (N_23309,N_22224,N_22685);
nand U23310 (N_23310,N_22382,N_22707);
or U23311 (N_23311,N_22138,N_22330);
or U23312 (N_23312,N_22597,N_22886);
and U23313 (N_23313,N_22985,N_22299);
xor U23314 (N_23314,N_22002,N_22966);
nor U23315 (N_23315,N_22590,N_22705);
or U23316 (N_23316,N_22892,N_22763);
and U23317 (N_23317,N_22779,N_22492);
xnor U23318 (N_23318,N_22315,N_22017);
or U23319 (N_23319,N_22380,N_22995);
and U23320 (N_23320,N_22542,N_22777);
and U23321 (N_23321,N_22209,N_22903);
xnor U23322 (N_23322,N_22169,N_22547);
or U23323 (N_23323,N_22160,N_22832);
and U23324 (N_23324,N_22879,N_22651);
and U23325 (N_23325,N_22179,N_22532);
xnor U23326 (N_23326,N_22902,N_22834);
nor U23327 (N_23327,N_22023,N_22147);
xor U23328 (N_23328,N_22233,N_22281);
xor U23329 (N_23329,N_22562,N_22032);
xnor U23330 (N_23330,N_22443,N_22250);
xor U23331 (N_23331,N_22069,N_22817);
xnor U23332 (N_23332,N_22731,N_22753);
xor U23333 (N_23333,N_22910,N_22806);
nand U23334 (N_23334,N_22448,N_22661);
or U23335 (N_23335,N_22314,N_22353);
nor U23336 (N_23336,N_22061,N_22851);
nand U23337 (N_23337,N_22415,N_22122);
or U23338 (N_23338,N_22193,N_22366);
or U23339 (N_23339,N_22469,N_22350);
nor U23340 (N_23340,N_22456,N_22478);
and U23341 (N_23341,N_22898,N_22671);
nor U23342 (N_23342,N_22852,N_22701);
nand U23343 (N_23343,N_22575,N_22451);
nand U23344 (N_23344,N_22669,N_22131);
nor U23345 (N_23345,N_22497,N_22447);
nand U23346 (N_23346,N_22768,N_22838);
and U23347 (N_23347,N_22367,N_22655);
xor U23348 (N_23348,N_22482,N_22049);
and U23349 (N_23349,N_22850,N_22606);
xor U23350 (N_23350,N_22163,N_22180);
nand U23351 (N_23351,N_22536,N_22014);
or U23352 (N_23352,N_22746,N_22072);
nor U23353 (N_23353,N_22078,N_22548);
nor U23354 (N_23354,N_22088,N_22034);
xnor U23355 (N_23355,N_22724,N_22285);
or U23356 (N_23356,N_22513,N_22199);
nand U23357 (N_23357,N_22345,N_22011);
and U23358 (N_23358,N_22862,N_22733);
and U23359 (N_23359,N_22080,N_22450);
and U23360 (N_23360,N_22081,N_22110);
and U23361 (N_23361,N_22470,N_22961);
nor U23362 (N_23362,N_22361,N_22500);
xnor U23363 (N_23363,N_22045,N_22248);
nand U23364 (N_23364,N_22282,N_22568);
xnor U23365 (N_23365,N_22737,N_22287);
or U23366 (N_23366,N_22587,N_22833);
and U23367 (N_23367,N_22136,N_22926);
nor U23368 (N_23368,N_22764,N_22709);
nand U23369 (N_23369,N_22373,N_22642);
nor U23370 (N_23370,N_22556,N_22686);
or U23371 (N_23371,N_22694,N_22561);
and U23372 (N_23372,N_22644,N_22249);
or U23373 (N_23373,N_22864,N_22001);
nand U23374 (N_23374,N_22825,N_22891);
or U23375 (N_23375,N_22401,N_22252);
nor U23376 (N_23376,N_22316,N_22437);
xor U23377 (N_23377,N_22409,N_22503);
and U23378 (N_23378,N_22870,N_22734);
or U23379 (N_23379,N_22026,N_22559);
nand U23380 (N_23380,N_22875,N_22377);
nand U23381 (N_23381,N_22841,N_22362);
xnor U23382 (N_23382,N_22405,N_22109);
nor U23383 (N_23383,N_22999,N_22517);
or U23384 (N_23384,N_22073,N_22098);
nand U23385 (N_23385,N_22393,N_22399);
and U23386 (N_23386,N_22613,N_22060);
nand U23387 (N_23387,N_22812,N_22351);
nor U23388 (N_23388,N_22566,N_22552);
xnor U23389 (N_23389,N_22752,N_22802);
nand U23390 (N_23390,N_22678,N_22269);
nor U23391 (N_23391,N_22486,N_22702);
xnor U23392 (N_23392,N_22107,N_22324);
or U23393 (N_23393,N_22969,N_22930);
xnor U23394 (N_23394,N_22826,N_22419);
nor U23395 (N_23395,N_22643,N_22809);
and U23396 (N_23396,N_22631,N_22951);
nand U23397 (N_23397,N_22094,N_22917);
nand U23398 (N_23398,N_22284,N_22792);
and U23399 (N_23399,N_22043,N_22663);
nand U23400 (N_23400,N_22266,N_22063);
nand U23401 (N_23401,N_22328,N_22920);
nor U23402 (N_23402,N_22518,N_22846);
nand U23403 (N_23403,N_22104,N_22267);
nand U23404 (N_23404,N_22959,N_22618);
xnor U23405 (N_23405,N_22593,N_22106);
nor U23406 (N_23406,N_22313,N_22810);
nand U23407 (N_23407,N_22150,N_22226);
xnor U23408 (N_23408,N_22206,N_22690);
nor U23409 (N_23409,N_22161,N_22276);
nand U23410 (N_23410,N_22564,N_22019);
xor U23411 (N_23411,N_22435,N_22111);
and U23412 (N_23412,N_22632,N_22854);
or U23413 (N_23413,N_22200,N_22171);
nor U23414 (N_23414,N_22509,N_22970);
xnor U23415 (N_23415,N_22221,N_22422);
and U23416 (N_23416,N_22374,N_22543);
or U23417 (N_23417,N_22074,N_22236);
nand U23418 (N_23418,N_22533,N_22364);
or U23419 (N_23419,N_22819,N_22550);
nor U23420 (N_23420,N_22112,N_22278);
and U23421 (N_23421,N_22955,N_22342);
nand U23422 (N_23422,N_22853,N_22502);
nand U23423 (N_23423,N_22544,N_22371);
nor U23424 (N_23424,N_22467,N_22843);
nand U23425 (N_23425,N_22799,N_22873);
nand U23426 (N_23426,N_22381,N_22211);
or U23427 (N_23427,N_22695,N_22495);
nor U23428 (N_23428,N_22453,N_22520);
or U23429 (N_23429,N_22653,N_22621);
nor U23430 (N_23430,N_22264,N_22333);
nand U23431 (N_23431,N_22581,N_22650);
and U23432 (N_23432,N_22402,N_22359);
nand U23433 (N_23433,N_22153,N_22251);
nor U23434 (N_23434,N_22363,N_22949);
nor U23435 (N_23435,N_22046,N_22645);
nor U23436 (N_23436,N_22883,N_22365);
nor U23437 (N_23437,N_22274,N_22114);
or U23438 (N_23438,N_22782,N_22234);
nor U23439 (N_23439,N_22079,N_22600);
xor U23440 (N_23440,N_22167,N_22849);
nand U23441 (N_23441,N_22496,N_22312);
nor U23442 (N_23442,N_22893,N_22390);
or U23443 (N_23443,N_22165,N_22527);
nand U23444 (N_23444,N_22047,N_22149);
nor U23445 (N_23445,N_22016,N_22231);
and U23446 (N_23446,N_22979,N_22433);
nand U23447 (N_23447,N_22962,N_22914);
or U23448 (N_23448,N_22939,N_22292);
or U23449 (N_23449,N_22130,N_22295);
nor U23450 (N_23450,N_22376,N_22410);
xnor U23451 (N_23451,N_22177,N_22749);
nand U23452 (N_23452,N_22828,N_22712);
nor U23453 (N_23453,N_22847,N_22534);
xor U23454 (N_23454,N_22739,N_22947);
and U23455 (N_23455,N_22085,N_22420);
or U23456 (N_23456,N_22641,N_22682);
xnor U23457 (N_23457,N_22622,N_22356);
xnor U23458 (N_23458,N_22430,N_22555);
and U23459 (N_23459,N_22210,N_22195);
or U23460 (N_23460,N_22242,N_22612);
or U23461 (N_23461,N_22656,N_22735);
nor U23462 (N_23462,N_22173,N_22908);
and U23463 (N_23463,N_22519,N_22037);
and U23464 (N_23464,N_22609,N_22119);
nor U23465 (N_23465,N_22203,N_22904);
and U23466 (N_23466,N_22595,N_22723);
and U23467 (N_23467,N_22005,N_22727);
and U23468 (N_23468,N_22580,N_22863);
or U23469 (N_23469,N_22256,N_22395);
nand U23470 (N_23470,N_22499,N_22479);
nand U23471 (N_23471,N_22855,N_22634);
or U23472 (N_23472,N_22941,N_22335);
nor U23473 (N_23473,N_22442,N_22997);
xor U23474 (N_23474,N_22309,N_22973);
nand U23475 (N_23475,N_22204,N_22243);
and U23476 (N_23476,N_22750,N_22865);
nand U23477 (N_23477,N_22142,N_22523);
or U23478 (N_23478,N_22039,N_22769);
nand U23479 (N_23479,N_22235,N_22302);
xor U23480 (N_23480,N_22223,N_22184);
xor U23481 (N_23481,N_22965,N_22958);
and U23482 (N_23482,N_22691,N_22426);
or U23483 (N_23483,N_22563,N_22125);
and U23484 (N_23484,N_22051,N_22239);
nand U23485 (N_23485,N_22636,N_22115);
nor U23486 (N_23486,N_22784,N_22293);
or U23487 (N_23487,N_22334,N_22042);
or U23488 (N_23488,N_22159,N_22596);
or U23489 (N_23489,N_22710,N_22240);
and U23490 (N_23490,N_22666,N_22458);
nand U23491 (N_23491,N_22814,N_22129);
nor U23492 (N_23492,N_22436,N_22439);
and U23493 (N_23493,N_22867,N_22494);
or U23494 (N_23494,N_22747,N_22654);
nand U23495 (N_23495,N_22751,N_22713);
or U23496 (N_23496,N_22012,N_22715);
nand U23497 (N_23497,N_22058,N_22332);
and U23498 (N_23498,N_22745,N_22708);
nor U23499 (N_23499,N_22878,N_22096);
or U23500 (N_23500,N_22980,N_22821);
nand U23501 (N_23501,N_22032,N_22233);
and U23502 (N_23502,N_22684,N_22634);
nand U23503 (N_23503,N_22101,N_22273);
nand U23504 (N_23504,N_22456,N_22655);
and U23505 (N_23505,N_22442,N_22122);
or U23506 (N_23506,N_22780,N_22540);
nor U23507 (N_23507,N_22332,N_22600);
or U23508 (N_23508,N_22030,N_22637);
nor U23509 (N_23509,N_22448,N_22056);
or U23510 (N_23510,N_22811,N_22265);
nand U23511 (N_23511,N_22664,N_22303);
nor U23512 (N_23512,N_22467,N_22311);
or U23513 (N_23513,N_22742,N_22602);
nand U23514 (N_23514,N_22953,N_22164);
nand U23515 (N_23515,N_22915,N_22716);
nand U23516 (N_23516,N_22187,N_22205);
xor U23517 (N_23517,N_22197,N_22398);
or U23518 (N_23518,N_22005,N_22242);
or U23519 (N_23519,N_22296,N_22185);
nand U23520 (N_23520,N_22598,N_22892);
xor U23521 (N_23521,N_22468,N_22264);
nor U23522 (N_23522,N_22820,N_22770);
nand U23523 (N_23523,N_22365,N_22962);
nor U23524 (N_23524,N_22028,N_22157);
and U23525 (N_23525,N_22558,N_22047);
nand U23526 (N_23526,N_22570,N_22133);
nor U23527 (N_23527,N_22571,N_22254);
and U23528 (N_23528,N_22271,N_22349);
xnor U23529 (N_23529,N_22944,N_22705);
and U23530 (N_23530,N_22695,N_22971);
and U23531 (N_23531,N_22278,N_22810);
or U23532 (N_23532,N_22548,N_22557);
and U23533 (N_23533,N_22237,N_22426);
nor U23534 (N_23534,N_22046,N_22219);
and U23535 (N_23535,N_22638,N_22915);
nand U23536 (N_23536,N_22309,N_22198);
xnor U23537 (N_23537,N_22227,N_22308);
nor U23538 (N_23538,N_22864,N_22527);
nand U23539 (N_23539,N_22646,N_22410);
or U23540 (N_23540,N_22769,N_22231);
xnor U23541 (N_23541,N_22479,N_22976);
and U23542 (N_23542,N_22018,N_22316);
or U23543 (N_23543,N_22003,N_22762);
or U23544 (N_23544,N_22586,N_22696);
nor U23545 (N_23545,N_22538,N_22571);
nand U23546 (N_23546,N_22102,N_22124);
and U23547 (N_23547,N_22068,N_22563);
or U23548 (N_23548,N_22270,N_22162);
and U23549 (N_23549,N_22911,N_22500);
nor U23550 (N_23550,N_22778,N_22506);
and U23551 (N_23551,N_22321,N_22092);
nor U23552 (N_23552,N_22081,N_22149);
nand U23553 (N_23553,N_22625,N_22198);
xnor U23554 (N_23554,N_22457,N_22492);
nor U23555 (N_23555,N_22591,N_22321);
nor U23556 (N_23556,N_22614,N_22803);
nand U23557 (N_23557,N_22552,N_22108);
and U23558 (N_23558,N_22799,N_22217);
xnor U23559 (N_23559,N_22388,N_22379);
and U23560 (N_23560,N_22962,N_22511);
nand U23561 (N_23561,N_22110,N_22464);
nor U23562 (N_23562,N_22324,N_22893);
nand U23563 (N_23563,N_22900,N_22473);
nand U23564 (N_23564,N_22888,N_22705);
or U23565 (N_23565,N_22157,N_22775);
xnor U23566 (N_23566,N_22689,N_22859);
nor U23567 (N_23567,N_22531,N_22625);
nand U23568 (N_23568,N_22632,N_22934);
xnor U23569 (N_23569,N_22498,N_22608);
or U23570 (N_23570,N_22745,N_22699);
xnor U23571 (N_23571,N_22753,N_22401);
nor U23572 (N_23572,N_22334,N_22229);
xnor U23573 (N_23573,N_22039,N_22027);
nand U23574 (N_23574,N_22307,N_22631);
nor U23575 (N_23575,N_22089,N_22810);
nand U23576 (N_23576,N_22424,N_22912);
and U23577 (N_23577,N_22808,N_22771);
or U23578 (N_23578,N_22903,N_22558);
nor U23579 (N_23579,N_22483,N_22418);
nor U23580 (N_23580,N_22311,N_22645);
xor U23581 (N_23581,N_22925,N_22882);
or U23582 (N_23582,N_22928,N_22310);
nand U23583 (N_23583,N_22403,N_22383);
nor U23584 (N_23584,N_22486,N_22508);
and U23585 (N_23585,N_22240,N_22628);
and U23586 (N_23586,N_22781,N_22904);
nor U23587 (N_23587,N_22520,N_22500);
and U23588 (N_23588,N_22883,N_22295);
xor U23589 (N_23589,N_22660,N_22261);
and U23590 (N_23590,N_22836,N_22776);
or U23591 (N_23591,N_22908,N_22041);
nor U23592 (N_23592,N_22496,N_22989);
xnor U23593 (N_23593,N_22396,N_22147);
nand U23594 (N_23594,N_22122,N_22864);
nor U23595 (N_23595,N_22479,N_22941);
nand U23596 (N_23596,N_22989,N_22068);
or U23597 (N_23597,N_22364,N_22979);
and U23598 (N_23598,N_22024,N_22820);
xnor U23599 (N_23599,N_22818,N_22474);
nand U23600 (N_23600,N_22521,N_22559);
and U23601 (N_23601,N_22048,N_22411);
or U23602 (N_23602,N_22179,N_22671);
xor U23603 (N_23603,N_22347,N_22322);
nor U23604 (N_23604,N_22693,N_22394);
xnor U23605 (N_23605,N_22465,N_22308);
nand U23606 (N_23606,N_22575,N_22019);
and U23607 (N_23607,N_22345,N_22958);
xnor U23608 (N_23608,N_22054,N_22153);
nor U23609 (N_23609,N_22363,N_22052);
or U23610 (N_23610,N_22549,N_22978);
nand U23611 (N_23611,N_22791,N_22217);
nand U23612 (N_23612,N_22933,N_22045);
or U23613 (N_23613,N_22492,N_22742);
nand U23614 (N_23614,N_22984,N_22603);
or U23615 (N_23615,N_22563,N_22444);
nand U23616 (N_23616,N_22910,N_22665);
and U23617 (N_23617,N_22043,N_22332);
xor U23618 (N_23618,N_22423,N_22151);
xnor U23619 (N_23619,N_22113,N_22220);
or U23620 (N_23620,N_22073,N_22211);
nor U23621 (N_23621,N_22576,N_22783);
nor U23622 (N_23622,N_22338,N_22880);
and U23623 (N_23623,N_22721,N_22754);
and U23624 (N_23624,N_22632,N_22438);
or U23625 (N_23625,N_22776,N_22401);
nor U23626 (N_23626,N_22257,N_22054);
nor U23627 (N_23627,N_22395,N_22721);
or U23628 (N_23628,N_22444,N_22196);
or U23629 (N_23629,N_22353,N_22301);
or U23630 (N_23630,N_22984,N_22851);
or U23631 (N_23631,N_22633,N_22454);
nor U23632 (N_23632,N_22117,N_22580);
xor U23633 (N_23633,N_22183,N_22919);
nor U23634 (N_23634,N_22795,N_22294);
nor U23635 (N_23635,N_22512,N_22865);
xor U23636 (N_23636,N_22671,N_22009);
or U23637 (N_23637,N_22387,N_22218);
xnor U23638 (N_23638,N_22469,N_22658);
xor U23639 (N_23639,N_22732,N_22683);
or U23640 (N_23640,N_22103,N_22249);
nand U23641 (N_23641,N_22318,N_22787);
and U23642 (N_23642,N_22832,N_22762);
xnor U23643 (N_23643,N_22735,N_22496);
nand U23644 (N_23644,N_22893,N_22382);
nor U23645 (N_23645,N_22690,N_22647);
nand U23646 (N_23646,N_22114,N_22573);
nor U23647 (N_23647,N_22600,N_22367);
nand U23648 (N_23648,N_22824,N_22619);
nand U23649 (N_23649,N_22922,N_22320);
and U23650 (N_23650,N_22391,N_22623);
nor U23651 (N_23651,N_22771,N_22515);
nand U23652 (N_23652,N_22301,N_22114);
or U23653 (N_23653,N_22613,N_22787);
or U23654 (N_23654,N_22545,N_22775);
nand U23655 (N_23655,N_22845,N_22527);
xor U23656 (N_23656,N_22624,N_22165);
and U23657 (N_23657,N_22369,N_22703);
xor U23658 (N_23658,N_22592,N_22685);
or U23659 (N_23659,N_22803,N_22102);
and U23660 (N_23660,N_22155,N_22224);
nand U23661 (N_23661,N_22800,N_22430);
or U23662 (N_23662,N_22164,N_22277);
nor U23663 (N_23663,N_22107,N_22396);
and U23664 (N_23664,N_22505,N_22057);
or U23665 (N_23665,N_22913,N_22505);
or U23666 (N_23666,N_22330,N_22510);
or U23667 (N_23667,N_22517,N_22939);
nand U23668 (N_23668,N_22697,N_22786);
nor U23669 (N_23669,N_22860,N_22686);
nand U23670 (N_23670,N_22663,N_22040);
or U23671 (N_23671,N_22252,N_22220);
xnor U23672 (N_23672,N_22071,N_22363);
xor U23673 (N_23673,N_22887,N_22976);
or U23674 (N_23674,N_22154,N_22899);
nand U23675 (N_23675,N_22770,N_22061);
or U23676 (N_23676,N_22703,N_22047);
or U23677 (N_23677,N_22249,N_22376);
nor U23678 (N_23678,N_22975,N_22681);
nand U23679 (N_23679,N_22868,N_22543);
nand U23680 (N_23680,N_22147,N_22844);
xnor U23681 (N_23681,N_22949,N_22533);
nand U23682 (N_23682,N_22723,N_22935);
nand U23683 (N_23683,N_22986,N_22548);
nor U23684 (N_23684,N_22024,N_22535);
and U23685 (N_23685,N_22037,N_22752);
and U23686 (N_23686,N_22512,N_22780);
nand U23687 (N_23687,N_22777,N_22001);
and U23688 (N_23688,N_22400,N_22804);
xnor U23689 (N_23689,N_22049,N_22980);
nand U23690 (N_23690,N_22208,N_22272);
nand U23691 (N_23691,N_22638,N_22471);
nand U23692 (N_23692,N_22814,N_22202);
xor U23693 (N_23693,N_22699,N_22959);
or U23694 (N_23694,N_22259,N_22980);
nor U23695 (N_23695,N_22454,N_22742);
nor U23696 (N_23696,N_22489,N_22351);
xor U23697 (N_23697,N_22628,N_22748);
or U23698 (N_23698,N_22926,N_22481);
xnor U23699 (N_23699,N_22559,N_22571);
or U23700 (N_23700,N_22179,N_22584);
and U23701 (N_23701,N_22164,N_22612);
or U23702 (N_23702,N_22908,N_22430);
nand U23703 (N_23703,N_22192,N_22183);
or U23704 (N_23704,N_22418,N_22743);
and U23705 (N_23705,N_22104,N_22734);
nor U23706 (N_23706,N_22674,N_22053);
or U23707 (N_23707,N_22321,N_22173);
or U23708 (N_23708,N_22271,N_22802);
and U23709 (N_23709,N_22554,N_22444);
or U23710 (N_23710,N_22095,N_22790);
and U23711 (N_23711,N_22770,N_22929);
nand U23712 (N_23712,N_22043,N_22558);
nor U23713 (N_23713,N_22697,N_22937);
nor U23714 (N_23714,N_22708,N_22190);
nor U23715 (N_23715,N_22975,N_22017);
xnor U23716 (N_23716,N_22753,N_22607);
nor U23717 (N_23717,N_22788,N_22650);
nand U23718 (N_23718,N_22984,N_22907);
or U23719 (N_23719,N_22264,N_22459);
nand U23720 (N_23720,N_22459,N_22412);
or U23721 (N_23721,N_22063,N_22579);
xnor U23722 (N_23722,N_22765,N_22941);
or U23723 (N_23723,N_22385,N_22989);
and U23724 (N_23724,N_22247,N_22355);
nor U23725 (N_23725,N_22692,N_22252);
xor U23726 (N_23726,N_22844,N_22490);
and U23727 (N_23727,N_22153,N_22529);
and U23728 (N_23728,N_22207,N_22679);
or U23729 (N_23729,N_22638,N_22938);
nand U23730 (N_23730,N_22858,N_22123);
xor U23731 (N_23731,N_22810,N_22470);
nand U23732 (N_23732,N_22937,N_22264);
nand U23733 (N_23733,N_22949,N_22105);
and U23734 (N_23734,N_22952,N_22351);
or U23735 (N_23735,N_22268,N_22174);
or U23736 (N_23736,N_22492,N_22654);
xnor U23737 (N_23737,N_22036,N_22311);
nand U23738 (N_23738,N_22279,N_22860);
and U23739 (N_23739,N_22745,N_22107);
xnor U23740 (N_23740,N_22542,N_22310);
nor U23741 (N_23741,N_22589,N_22933);
nand U23742 (N_23742,N_22879,N_22145);
and U23743 (N_23743,N_22823,N_22890);
or U23744 (N_23744,N_22043,N_22260);
nor U23745 (N_23745,N_22750,N_22684);
nor U23746 (N_23746,N_22610,N_22126);
or U23747 (N_23747,N_22783,N_22360);
or U23748 (N_23748,N_22304,N_22632);
and U23749 (N_23749,N_22499,N_22097);
xor U23750 (N_23750,N_22454,N_22105);
nor U23751 (N_23751,N_22603,N_22058);
nand U23752 (N_23752,N_22823,N_22746);
and U23753 (N_23753,N_22601,N_22678);
xor U23754 (N_23754,N_22932,N_22277);
nand U23755 (N_23755,N_22077,N_22387);
or U23756 (N_23756,N_22511,N_22382);
nand U23757 (N_23757,N_22702,N_22982);
nand U23758 (N_23758,N_22241,N_22487);
or U23759 (N_23759,N_22976,N_22435);
or U23760 (N_23760,N_22357,N_22213);
and U23761 (N_23761,N_22237,N_22572);
xnor U23762 (N_23762,N_22087,N_22158);
xnor U23763 (N_23763,N_22151,N_22822);
and U23764 (N_23764,N_22081,N_22397);
xnor U23765 (N_23765,N_22153,N_22208);
xor U23766 (N_23766,N_22303,N_22831);
nand U23767 (N_23767,N_22752,N_22535);
and U23768 (N_23768,N_22159,N_22308);
xor U23769 (N_23769,N_22485,N_22966);
and U23770 (N_23770,N_22261,N_22431);
nor U23771 (N_23771,N_22543,N_22429);
or U23772 (N_23772,N_22354,N_22537);
nand U23773 (N_23773,N_22748,N_22417);
nor U23774 (N_23774,N_22341,N_22070);
xnor U23775 (N_23775,N_22031,N_22397);
nor U23776 (N_23776,N_22642,N_22654);
and U23777 (N_23777,N_22542,N_22376);
xor U23778 (N_23778,N_22872,N_22549);
xor U23779 (N_23779,N_22246,N_22521);
or U23780 (N_23780,N_22678,N_22850);
nand U23781 (N_23781,N_22468,N_22506);
nand U23782 (N_23782,N_22698,N_22921);
nand U23783 (N_23783,N_22972,N_22795);
and U23784 (N_23784,N_22782,N_22836);
nor U23785 (N_23785,N_22224,N_22438);
nor U23786 (N_23786,N_22304,N_22402);
nor U23787 (N_23787,N_22311,N_22456);
nor U23788 (N_23788,N_22661,N_22892);
xnor U23789 (N_23789,N_22298,N_22799);
nor U23790 (N_23790,N_22217,N_22438);
xnor U23791 (N_23791,N_22386,N_22879);
nor U23792 (N_23792,N_22491,N_22654);
nand U23793 (N_23793,N_22459,N_22617);
xnor U23794 (N_23794,N_22778,N_22865);
or U23795 (N_23795,N_22348,N_22306);
xor U23796 (N_23796,N_22993,N_22393);
and U23797 (N_23797,N_22041,N_22030);
nand U23798 (N_23798,N_22095,N_22568);
nor U23799 (N_23799,N_22729,N_22417);
xnor U23800 (N_23800,N_22737,N_22921);
nor U23801 (N_23801,N_22454,N_22234);
or U23802 (N_23802,N_22632,N_22194);
nand U23803 (N_23803,N_22736,N_22950);
and U23804 (N_23804,N_22229,N_22062);
nor U23805 (N_23805,N_22669,N_22200);
nor U23806 (N_23806,N_22369,N_22217);
nand U23807 (N_23807,N_22722,N_22997);
nor U23808 (N_23808,N_22245,N_22118);
xnor U23809 (N_23809,N_22367,N_22752);
or U23810 (N_23810,N_22028,N_22490);
and U23811 (N_23811,N_22814,N_22444);
and U23812 (N_23812,N_22609,N_22467);
xor U23813 (N_23813,N_22122,N_22895);
nor U23814 (N_23814,N_22278,N_22870);
xnor U23815 (N_23815,N_22194,N_22514);
nand U23816 (N_23816,N_22359,N_22372);
nand U23817 (N_23817,N_22204,N_22132);
xor U23818 (N_23818,N_22457,N_22265);
or U23819 (N_23819,N_22820,N_22747);
nand U23820 (N_23820,N_22748,N_22405);
or U23821 (N_23821,N_22591,N_22349);
nand U23822 (N_23822,N_22104,N_22300);
nand U23823 (N_23823,N_22580,N_22370);
and U23824 (N_23824,N_22364,N_22852);
nor U23825 (N_23825,N_22326,N_22281);
or U23826 (N_23826,N_22881,N_22812);
or U23827 (N_23827,N_22496,N_22017);
xor U23828 (N_23828,N_22044,N_22976);
nor U23829 (N_23829,N_22430,N_22977);
xnor U23830 (N_23830,N_22802,N_22433);
or U23831 (N_23831,N_22245,N_22349);
or U23832 (N_23832,N_22700,N_22807);
nor U23833 (N_23833,N_22103,N_22453);
xnor U23834 (N_23834,N_22586,N_22155);
nand U23835 (N_23835,N_22423,N_22727);
or U23836 (N_23836,N_22000,N_22184);
or U23837 (N_23837,N_22491,N_22083);
nand U23838 (N_23838,N_22820,N_22797);
and U23839 (N_23839,N_22571,N_22109);
and U23840 (N_23840,N_22108,N_22298);
xnor U23841 (N_23841,N_22524,N_22609);
nor U23842 (N_23842,N_22615,N_22193);
and U23843 (N_23843,N_22274,N_22607);
xor U23844 (N_23844,N_22956,N_22098);
and U23845 (N_23845,N_22202,N_22666);
and U23846 (N_23846,N_22587,N_22955);
and U23847 (N_23847,N_22801,N_22267);
or U23848 (N_23848,N_22572,N_22158);
or U23849 (N_23849,N_22566,N_22749);
and U23850 (N_23850,N_22666,N_22220);
and U23851 (N_23851,N_22341,N_22695);
xor U23852 (N_23852,N_22715,N_22181);
nor U23853 (N_23853,N_22231,N_22915);
or U23854 (N_23854,N_22000,N_22023);
or U23855 (N_23855,N_22644,N_22384);
nor U23856 (N_23856,N_22487,N_22141);
nor U23857 (N_23857,N_22861,N_22982);
xor U23858 (N_23858,N_22989,N_22960);
nand U23859 (N_23859,N_22090,N_22407);
nand U23860 (N_23860,N_22718,N_22801);
and U23861 (N_23861,N_22882,N_22454);
or U23862 (N_23862,N_22795,N_22202);
nand U23863 (N_23863,N_22642,N_22756);
or U23864 (N_23864,N_22503,N_22328);
xor U23865 (N_23865,N_22700,N_22535);
or U23866 (N_23866,N_22068,N_22924);
and U23867 (N_23867,N_22174,N_22774);
nor U23868 (N_23868,N_22370,N_22518);
nor U23869 (N_23869,N_22672,N_22961);
nand U23870 (N_23870,N_22309,N_22980);
nand U23871 (N_23871,N_22247,N_22419);
xnor U23872 (N_23872,N_22140,N_22602);
xor U23873 (N_23873,N_22424,N_22009);
nor U23874 (N_23874,N_22157,N_22128);
or U23875 (N_23875,N_22413,N_22306);
nor U23876 (N_23876,N_22849,N_22730);
nand U23877 (N_23877,N_22172,N_22144);
nand U23878 (N_23878,N_22052,N_22465);
or U23879 (N_23879,N_22372,N_22088);
xor U23880 (N_23880,N_22080,N_22576);
and U23881 (N_23881,N_22812,N_22828);
xor U23882 (N_23882,N_22762,N_22021);
nand U23883 (N_23883,N_22322,N_22052);
nor U23884 (N_23884,N_22683,N_22563);
nand U23885 (N_23885,N_22479,N_22518);
nor U23886 (N_23886,N_22176,N_22950);
nor U23887 (N_23887,N_22555,N_22329);
nor U23888 (N_23888,N_22979,N_22292);
xor U23889 (N_23889,N_22768,N_22058);
or U23890 (N_23890,N_22052,N_22306);
nand U23891 (N_23891,N_22422,N_22978);
xor U23892 (N_23892,N_22367,N_22574);
xor U23893 (N_23893,N_22414,N_22775);
nor U23894 (N_23894,N_22892,N_22742);
nand U23895 (N_23895,N_22569,N_22394);
nand U23896 (N_23896,N_22144,N_22382);
nor U23897 (N_23897,N_22446,N_22631);
and U23898 (N_23898,N_22262,N_22609);
nand U23899 (N_23899,N_22341,N_22748);
nor U23900 (N_23900,N_22679,N_22153);
and U23901 (N_23901,N_22714,N_22505);
xor U23902 (N_23902,N_22571,N_22022);
and U23903 (N_23903,N_22267,N_22787);
nand U23904 (N_23904,N_22246,N_22168);
nor U23905 (N_23905,N_22166,N_22812);
nor U23906 (N_23906,N_22750,N_22102);
nand U23907 (N_23907,N_22287,N_22610);
nor U23908 (N_23908,N_22432,N_22191);
nand U23909 (N_23909,N_22174,N_22280);
xor U23910 (N_23910,N_22483,N_22100);
nor U23911 (N_23911,N_22014,N_22242);
nor U23912 (N_23912,N_22621,N_22541);
nand U23913 (N_23913,N_22144,N_22364);
nand U23914 (N_23914,N_22771,N_22697);
and U23915 (N_23915,N_22605,N_22751);
nor U23916 (N_23916,N_22492,N_22841);
nor U23917 (N_23917,N_22256,N_22807);
or U23918 (N_23918,N_22309,N_22502);
or U23919 (N_23919,N_22018,N_22147);
xor U23920 (N_23920,N_22475,N_22450);
nor U23921 (N_23921,N_22739,N_22180);
nor U23922 (N_23922,N_22445,N_22142);
nand U23923 (N_23923,N_22679,N_22149);
nor U23924 (N_23924,N_22759,N_22401);
and U23925 (N_23925,N_22530,N_22317);
xor U23926 (N_23926,N_22190,N_22433);
and U23927 (N_23927,N_22790,N_22807);
xor U23928 (N_23928,N_22228,N_22859);
xnor U23929 (N_23929,N_22220,N_22125);
or U23930 (N_23930,N_22739,N_22075);
nand U23931 (N_23931,N_22463,N_22586);
and U23932 (N_23932,N_22216,N_22383);
nand U23933 (N_23933,N_22364,N_22295);
nand U23934 (N_23934,N_22115,N_22907);
xor U23935 (N_23935,N_22013,N_22676);
nor U23936 (N_23936,N_22752,N_22091);
nand U23937 (N_23937,N_22557,N_22185);
nor U23938 (N_23938,N_22138,N_22924);
or U23939 (N_23939,N_22195,N_22139);
and U23940 (N_23940,N_22058,N_22920);
nor U23941 (N_23941,N_22603,N_22933);
nand U23942 (N_23942,N_22907,N_22889);
nor U23943 (N_23943,N_22232,N_22939);
nor U23944 (N_23944,N_22011,N_22436);
xnor U23945 (N_23945,N_22215,N_22072);
nand U23946 (N_23946,N_22708,N_22959);
and U23947 (N_23947,N_22743,N_22670);
and U23948 (N_23948,N_22181,N_22660);
nor U23949 (N_23949,N_22694,N_22353);
nor U23950 (N_23950,N_22384,N_22365);
nor U23951 (N_23951,N_22998,N_22815);
or U23952 (N_23952,N_22070,N_22393);
xnor U23953 (N_23953,N_22534,N_22341);
and U23954 (N_23954,N_22542,N_22751);
and U23955 (N_23955,N_22187,N_22540);
or U23956 (N_23956,N_22299,N_22027);
or U23957 (N_23957,N_22993,N_22544);
nor U23958 (N_23958,N_22742,N_22342);
and U23959 (N_23959,N_22351,N_22281);
nor U23960 (N_23960,N_22012,N_22193);
nor U23961 (N_23961,N_22442,N_22113);
or U23962 (N_23962,N_22633,N_22577);
and U23963 (N_23963,N_22500,N_22720);
nor U23964 (N_23964,N_22713,N_22891);
or U23965 (N_23965,N_22058,N_22415);
and U23966 (N_23966,N_22320,N_22374);
and U23967 (N_23967,N_22501,N_22681);
and U23968 (N_23968,N_22191,N_22514);
nand U23969 (N_23969,N_22251,N_22671);
and U23970 (N_23970,N_22183,N_22995);
and U23971 (N_23971,N_22815,N_22859);
xor U23972 (N_23972,N_22325,N_22949);
xnor U23973 (N_23973,N_22172,N_22147);
and U23974 (N_23974,N_22302,N_22240);
or U23975 (N_23975,N_22206,N_22156);
nor U23976 (N_23976,N_22987,N_22428);
and U23977 (N_23977,N_22301,N_22434);
and U23978 (N_23978,N_22822,N_22083);
nor U23979 (N_23979,N_22261,N_22588);
xor U23980 (N_23980,N_22701,N_22253);
and U23981 (N_23981,N_22356,N_22315);
nand U23982 (N_23982,N_22412,N_22464);
nand U23983 (N_23983,N_22823,N_22388);
nand U23984 (N_23984,N_22230,N_22515);
or U23985 (N_23985,N_22436,N_22686);
nand U23986 (N_23986,N_22443,N_22332);
nand U23987 (N_23987,N_22774,N_22257);
nor U23988 (N_23988,N_22530,N_22037);
xor U23989 (N_23989,N_22344,N_22956);
and U23990 (N_23990,N_22268,N_22047);
or U23991 (N_23991,N_22273,N_22010);
nor U23992 (N_23992,N_22449,N_22574);
nor U23993 (N_23993,N_22943,N_22461);
and U23994 (N_23994,N_22583,N_22547);
nor U23995 (N_23995,N_22406,N_22968);
or U23996 (N_23996,N_22287,N_22814);
and U23997 (N_23997,N_22930,N_22549);
nand U23998 (N_23998,N_22019,N_22061);
nand U23999 (N_23999,N_22977,N_22954);
or U24000 (N_24000,N_23187,N_23421);
xnor U24001 (N_24001,N_23669,N_23019);
and U24002 (N_24002,N_23442,N_23139);
xor U24003 (N_24003,N_23456,N_23193);
xnor U24004 (N_24004,N_23275,N_23295);
nand U24005 (N_24005,N_23915,N_23099);
nor U24006 (N_24006,N_23638,N_23071);
and U24007 (N_24007,N_23507,N_23986);
and U24008 (N_24008,N_23525,N_23124);
nor U24009 (N_24009,N_23933,N_23870);
or U24010 (N_24010,N_23991,N_23726);
or U24011 (N_24011,N_23311,N_23856);
nand U24012 (N_24012,N_23143,N_23341);
and U24013 (N_24013,N_23619,N_23871);
nor U24014 (N_24014,N_23068,N_23469);
nor U24015 (N_24015,N_23861,N_23766);
xor U24016 (N_24016,N_23715,N_23501);
nand U24017 (N_24017,N_23120,N_23680);
xor U24018 (N_24018,N_23675,N_23605);
nor U24019 (N_24019,N_23452,N_23928);
or U24020 (N_24020,N_23976,N_23502);
nor U24021 (N_24021,N_23086,N_23274);
xor U24022 (N_24022,N_23390,N_23566);
xor U24023 (N_24023,N_23499,N_23495);
nand U24024 (N_24024,N_23937,N_23446);
xor U24025 (N_24025,N_23153,N_23836);
nor U24026 (N_24026,N_23564,N_23169);
nor U24027 (N_24027,N_23480,N_23087);
or U24028 (N_24028,N_23388,N_23303);
and U24029 (N_24029,N_23848,N_23665);
nor U24030 (N_24030,N_23774,N_23326);
nor U24031 (N_24031,N_23111,N_23066);
nor U24032 (N_24032,N_23198,N_23984);
and U24033 (N_24033,N_23339,N_23897);
nor U24034 (N_24034,N_23243,N_23467);
nand U24035 (N_24035,N_23541,N_23651);
nand U24036 (N_24036,N_23258,N_23902);
xor U24037 (N_24037,N_23724,N_23613);
nand U24038 (N_24038,N_23729,N_23385);
or U24039 (N_24039,N_23445,N_23404);
and U24040 (N_24040,N_23573,N_23321);
nand U24041 (N_24041,N_23441,N_23132);
nor U24042 (N_24042,N_23225,N_23824);
or U24043 (N_24043,N_23489,N_23955);
and U24044 (N_24044,N_23759,N_23927);
or U24045 (N_24045,N_23786,N_23118);
or U24046 (N_24046,N_23214,N_23550);
xnor U24047 (N_24047,N_23135,N_23366);
and U24048 (N_24048,N_23438,N_23025);
or U24049 (N_24049,N_23043,N_23455);
xnor U24050 (N_24050,N_23616,N_23355);
and U24051 (N_24051,N_23022,N_23723);
or U24052 (N_24052,N_23805,N_23027);
nor U24053 (N_24053,N_23626,N_23868);
xor U24054 (N_24054,N_23002,N_23867);
or U24055 (N_24055,N_23492,N_23894);
nor U24056 (N_24056,N_23281,N_23748);
nor U24057 (N_24057,N_23136,N_23627);
or U24058 (N_24058,N_23758,N_23182);
and U24059 (N_24059,N_23752,N_23138);
nand U24060 (N_24060,N_23249,N_23858);
and U24061 (N_24061,N_23575,N_23367);
nor U24062 (N_24062,N_23200,N_23743);
nor U24063 (N_24063,N_23907,N_23289);
xnor U24064 (N_24064,N_23211,N_23330);
nand U24065 (N_24065,N_23094,N_23514);
nand U24066 (N_24066,N_23017,N_23375);
nand U24067 (N_24067,N_23213,N_23447);
and U24068 (N_24068,N_23063,N_23217);
or U24069 (N_24069,N_23505,N_23271);
xnor U24070 (N_24070,N_23359,N_23623);
or U24071 (N_24071,N_23992,N_23942);
and U24072 (N_24072,N_23543,N_23049);
and U24073 (N_24073,N_23828,N_23924);
nor U24074 (N_24074,N_23462,N_23067);
or U24075 (N_24075,N_23551,N_23315);
or U24076 (N_24076,N_23686,N_23795);
nand U24077 (N_24077,N_23116,N_23270);
or U24078 (N_24078,N_23678,N_23329);
and U24079 (N_24079,N_23414,N_23978);
or U24080 (N_24080,N_23957,N_23711);
xnor U24081 (N_24081,N_23065,N_23152);
nand U24082 (N_24082,N_23140,N_23659);
nand U24083 (N_24083,N_23267,N_23058);
nand U24084 (N_24084,N_23688,N_23684);
or U24085 (N_24085,N_23356,N_23430);
nor U24086 (N_24086,N_23024,N_23231);
nand U24087 (N_24087,N_23048,N_23674);
and U24088 (N_24088,N_23497,N_23736);
nand U24089 (N_24089,N_23183,N_23996);
nor U24090 (N_24090,N_23685,N_23847);
and U24091 (N_24091,N_23670,N_23000);
xor U24092 (N_24092,N_23888,N_23583);
xnor U24093 (N_24093,N_23005,N_23484);
or U24094 (N_24094,N_23055,N_23895);
and U24095 (N_24095,N_23188,N_23285);
and U24096 (N_24096,N_23589,N_23730);
or U24097 (N_24097,N_23639,N_23648);
or U24098 (N_24098,N_23202,N_23760);
xnor U24099 (N_24099,N_23168,N_23596);
nand U24100 (N_24100,N_23754,N_23052);
nor U24101 (N_24101,N_23150,N_23558);
nand U24102 (N_24102,N_23245,N_23177);
nand U24103 (N_24103,N_23692,N_23379);
nor U24104 (N_24104,N_23069,N_23015);
xnor U24105 (N_24105,N_23640,N_23598);
xor U24106 (N_24106,N_23265,N_23434);
xor U24107 (N_24107,N_23560,N_23905);
nor U24108 (N_24108,N_23632,N_23783);
xor U24109 (N_24109,N_23586,N_23588);
nand U24110 (N_24110,N_23280,N_23221);
and U24111 (N_24111,N_23687,N_23533);
or U24112 (N_24112,N_23407,N_23234);
nand U24113 (N_24113,N_23579,N_23718);
or U24114 (N_24114,N_23468,N_23568);
and U24115 (N_24115,N_23268,N_23037);
or U24116 (N_24116,N_23802,N_23083);
nand U24117 (N_24117,N_23040,N_23879);
and U24118 (N_24118,N_23157,N_23948);
xnor U24119 (N_24119,N_23698,N_23705);
xor U24120 (N_24120,N_23580,N_23765);
and U24121 (N_24121,N_23628,N_23323);
or U24122 (N_24122,N_23018,N_23534);
nand U24123 (N_24123,N_23701,N_23464);
nor U24124 (N_24124,N_23959,N_23725);
nand U24125 (N_24125,N_23056,N_23798);
xnor U24126 (N_24126,N_23463,N_23911);
nor U24127 (N_24127,N_23634,N_23472);
nor U24128 (N_24128,N_23031,N_23232);
xor U24129 (N_24129,N_23522,N_23372);
nor U24130 (N_24130,N_23695,N_23335);
nand U24131 (N_24131,N_23133,N_23337);
or U24132 (N_24132,N_23491,N_23710);
xnor U24133 (N_24133,N_23839,N_23235);
and U24134 (N_24134,N_23382,N_23284);
or U24135 (N_24135,N_23607,N_23935);
and U24136 (N_24136,N_23590,N_23204);
and U24137 (N_24137,N_23361,N_23498);
or U24138 (N_24138,N_23435,N_23961);
xnor U24139 (N_24139,N_23872,N_23577);
nor U24140 (N_24140,N_23841,N_23401);
and U24141 (N_24141,N_23343,N_23413);
and U24142 (N_24142,N_23127,N_23344);
or U24143 (N_24143,N_23768,N_23142);
or U24144 (N_24144,N_23951,N_23047);
xor U24145 (N_24145,N_23950,N_23887);
xor U24146 (N_24146,N_23548,N_23478);
nand U24147 (N_24147,N_23333,N_23418);
and U24148 (N_24148,N_23925,N_23045);
nand U24149 (N_24149,N_23792,N_23220);
nor U24150 (N_24150,N_23131,N_23247);
nand U24151 (N_24151,N_23041,N_23614);
nand U24152 (N_24152,N_23443,N_23500);
nand U24153 (N_24153,N_23091,N_23694);
nor U24154 (N_24154,N_23970,N_23195);
and U24155 (N_24155,N_23165,N_23369);
and U24156 (N_24156,N_23449,N_23511);
nand U24157 (N_24157,N_23877,N_23512);
or U24158 (N_24158,N_23524,N_23529);
nor U24159 (N_24159,N_23601,N_23400);
nand U24160 (N_24160,N_23515,N_23663);
nor U24161 (N_24161,N_23542,N_23676);
xor U24162 (N_24162,N_23237,N_23011);
or U24163 (N_24163,N_23784,N_23318);
nor U24164 (N_24164,N_23657,N_23677);
nand U24165 (N_24165,N_23812,N_23633);
or U24166 (N_24166,N_23395,N_23526);
or U24167 (N_24167,N_23833,N_23277);
and U24168 (N_24168,N_23154,N_23039);
nand U24169 (N_24169,N_23660,N_23399);
xnor U24170 (N_24170,N_23362,N_23749);
and U24171 (N_24171,N_23003,N_23103);
nand U24172 (N_24172,N_23717,N_23163);
nand U24173 (N_24173,N_23365,N_23181);
xor U24174 (N_24174,N_23461,N_23556);
nand U24175 (N_24175,N_23849,N_23020);
and U24176 (N_24176,N_23953,N_23806);
nand U24177 (N_24177,N_23075,N_23900);
xor U24178 (N_24178,N_23174,N_23353);
and U24179 (N_24179,N_23578,N_23458);
nand U24180 (N_24180,N_23819,N_23096);
and U24181 (N_24181,N_23770,N_23913);
and U24182 (N_24182,N_23767,N_23531);
or U24183 (N_24183,N_23779,N_23745);
xnor U24184 (N_24184,N_23538,N_23506);
nor U24185 (N_24185,N_23654,N_23830);
xor U24186 (N_24186,N_23192,N_23123);
and U24187 (N_24187,N_23901,N_23034);
or U24188 (N_24188,N_23916,N_23829);
or U24189 (N_24189,N_23958,N_23302);
or U24190 (N_24190,N_23423,N_23523);
and U24191 (N_24191,N_23797,N_23671);
or U24192 (N_24192,N_23952,N_23304);
nor U24193 (N_24193,N_23473,N_23866);
xor U24194 (N_24194,N_23835,N_23609);
nor U24195 (N_24195,N_23381,N_23788);
and U24196 (N_24196,N_23890,N_23602);
nand U24197 (N_24197,N_23346,N_23403);
nand U24198 (N_24198,N_23763,N_23509);
or U24199 (N_24199,N_23972,N_23929);
xnor U24200 (N_24200,N_23644,N_23857);
xnor U24201 (N_24201,N_23728,N_23439);
nand U24202 (N_24202,N_23023,N_23876);
and U24203 (N_24203,N_23719,N_23371);
nor U24204 (N_24204,N_23918,N_23853);
and U24205 (N_24205,N_23260,N_23079);
and U24206 (N_24206,N_23417,N_23689);
and U24207 (N_24207,N_23815,N_23610);
xor U24208 (N_24208,N_23209,N_23826);
xnor U24209 (N_24209,N_23691,N_23425);
or U24210 (N_24210,N_23300,N_23148);
and U24211 (N_24211,N_23042,N_23149);
xnor U24212 (N_24212,N_23773,N_23386);
or U24213 (N_24213,N_23855,N_23557);
xnor U24214 (N_24214,N_23799,N_23820);
nor U24215 (N_24215,N_23668,N_23842);
xnor U24216 (N_24216,N_23844,N_23097);
nor U24217 (N_24217,N_23158,N_23966);
and U24218 (N_24218,N_23553,N_23062);
and U24219 (N_24219,N_23263,N_23771);
nand U24220 (N_24220,N_23219,N_23721);
or U24221 (N_24221,N_23228,N_23969);
nor U24222 (N_24222,N_23466,N_23903);
nor U24223 (N_24223,N_23248,N_23528);
or U24224 (N_24224,N_23012,N_23536);
or U24225 (N_24225,N_23883,N_23269);
nor U24226 (N_24226,N_23380,N_23622);
nand U24227 (N_24227,N_23089,N_23702);
or U24228 (N_24228,N_23737,N_23394);
nor U24229 (N_24229,N_23882,N_23117);
xor U24230 (N_24230,N_23661,N_23741);
or U24231 (N_24231,N_23134,N_23073);
nor U24232 (N_24232,N_23338,N_23546);
and U24233 (N_24233,N_23794,N_23910);
nor U24234 (N_24234,N_23276,N_23904);
nor U24235 (N_24235,N_23322,N_23813);
or U24236 (N_24236,N_23643,N_23176);
nand U24237 (N_24237,N_23584,N_23532);
nor U24238 (N_24238,N_23823,N_23351);
nor U24239 (N_24239,N_23253,N_23254);
nor U24240 (N_24240,N_23137,N_23530);
and U24241 (N_24241,N_23030,N_23057);
nor U24242 (N_24242,N_23161,N_23947);
xnor U24243 (N_24243,N_23620,N_23215);
nor U24244 (N_24244,N_23283,N_23286);
nor U24245 (N_24245,N_23544,N_23206);
or U24246 (N_24246,N_23964,N_23974);
and U24247 (N_24247,N_23988,N_23255);
xor U24248 (N_24248,N_23510,N_23053);
and U24249 (N_24249,N_23772,N_23340);
and U24250 (N_24250,N_23921,N_23862);
nor U24251 (N_24251,N_23681,N_23860);
nand U24252 (N_24252,N_23886,N_23190);
nor U24253 (N_24253,N_23252,N_23946);
xor U24254 (N_24254,N_23465,N_23873);
and U24255 (N_24255,N_23306,N_23282);
nand U24256 (N_24256,N_23625,N_23426);
or U24257 (N_24257,N_23785,N_23994);
nor U24258 (N_24258,N_23007,N_23384);
and U24259 (N_24259,N_23834,N_23398);
nand U24260 (N_24260,N_23576,N_23451);
nand U24261 (N_24261,N_23299,N_23238);
or U24262 (N_24262,N_23965,N_23405);
or U24263 (N_24263,N_23013,N_23272);
or U24264 (N_24264,N_23880,N_23054);
nand U24265 (N_24265,N_23494,N_23761);
nor U24266 (N_24266,N_23072,N_23803);
and U24267 (N_24267,N_23081,N_23029);
xor U24268 (N_24268,N_23744,N_23008);
or U24269 (N_24269,N_23940,N_23808);
or U24270 (N_24270,N_23036,N_23328);
or U24271 (N_24271,N_23316,N_23664);
nand U24272 (N_24272,N_23453,N_23982);
nor U24273 (N_24273,N_23378,N_23308);
xnor U24274 (N_24274,N_23733,N_23108);
and U24275 (N_24275,N_23391,N_23869);
xnor U24276 (N_24276,N_23076,N_23433);
xnor U24277 (N_24277,N_23571,N_23297);
or U24278 (N_24278,N_23014,N_23679);
xnor U24279 (N_24279,N_23720,N_23327);
and U24280 (N_24280,N_23305,N_23349);
xnor U24281 (N_24281,N_23397,N_23545);
nor U24282 (N_24282,N_23061,N_23840);
and U24283 (N_24283,N_23121,N_23292);
nand U24284 (N_24284,N_23936,N_23059);
or U24285 (N_24285,N_23811,N_23521);
nand U24286 (N_24286,N_23482,N_23508);
nand U24287 (N_24287,N_23113,N_23821);
nand U24288 (N_24288,N_23939,N_23738);
and U24289 (N_24289,N_23769,N_23264);
or U24290 (N_24290,N_23100,N_23776);
xor U24291 (N_24291,N_23889,N_23084);
nor U24292 (N_24292,N_23082,N_23600);
or U24293 (N_24293,N_23156,N_23552);
and U24294 (N_24294,N_23166,N_23230);
nor U24295 (N_24295,N_23934,N_23666);
and U24296 (N_24296,N_23009,N_23621);
nand U24297 (N_24297,N_23406,N_23930);
or U24298 (N_24298,N_23459,N_23298);
or U24299 (N_24299,N_23727,N_23816);
or U24300 (N_24300,N_23440,N_23756);
or U24301 (N_24301,N_23985,N_23878);
and U24302 (N_24302,N_23077,N_23817);
nor U24303 (N_24303,N_23854,N_23350);
nor U24304 (N_24304,N_23962,N_23360);
xor U24305 (N_24305,N_23968,N_23160);
nand U24306 (N_24306,N_23892,N_23408);
and U24307 (N_24307,N_23646,N_23171);
and U24308 (N_24308,N_23092,N_23241);
and U24309 (N_24309,N_23288,N_23064);
or U24310 (N_24310,N_23793,N_23909);
nor U24311 (N_24311,N_23926,N_23611);
xor U24312 (N_24312,N_23266,N_23242);
or U24313 (N_24313,N_23922,N_23098);
nor U24314 (N_24314,N_23262,N_23696);
xnor U24315 (N_24315,N_23863,N_23383);
or U24316 (N_24316,N_23809,N_23419);
xnor U24317 (N_24317,N_23147,N_23368);
and U24318 (N_24318,N_23637,N_23095);
or U24319 (N_24319,N_23592,N_23708);
nand U24320 (N_24320,N_23294,N_23891);
xnor U24321 (N_24321,N_23424,N_23561);
nand U24322 (N_24322,N_23479,N_23212);
and U24323 (N_24323,N_23706,N_23226);
or U24324 (N_24324,N_23975,N_23980);
nor U24325 (N_24325,N_23251,N_23981);
or U24326 (N_24326,N_23093,N_23649);
nor U24327 (N_24327,N_23026,N_23593);
and U24328 (N_24328,N_23070,N_23781);
and U24329 (N_24329,N_23179,N_23700);
nor U24330 (N_24330,N_23631,N_23257);
nor U24331 (N_24331,N_23010,N_23287);
or U24332 (N_24332,N_23410,N_23477);
nand U24333 (N_24333,N_23144,N_23516);
or U24334 (N_24334,N_23218,N_23747);
and U24335 (N_24335,N_23599,N_23309);
nand U24336 (N_24336,N_23085,N_23396);
nand U24337 (N_24337,N_23852,N_23504);
or U24338 (N_24338,N_23683,N_23141);
xor U24339 (N_24339,N_23540,N_23486);
xnor U24340 (N_24340,N_23487,N_23595);
and U24341 (N_24341,N_23581,N_23697);
and U24342 (N_24342,N_23481,N_23606);
or U24343 (N_24343,N_23941,N_23320);
or U24344 (N_24344,N_23537,N_23513);
xnor U24345 (N_24345,N_23313,N_23110);
xor U24346 (N_24346,N_23296,N_23370);
nand U24347 (N_24347,N_23535,N_23427);
nand U24348 (N_24348,N_23731,N_23734);
xnor U24349 (N_24349,N_23347,N_23750);
xor U24350 (N_24350,N_23757,N_23125);
nor U24351 (N_24351,N_23565,N_23653);
nand U24352 (N_24352,N_23570,N_23585);
nor U24353 (N_24353,N_23493,N_23742);
or U24354 (N_24354,N_23210,N_23874);
or U24355 (N_24355,N_23485,N_23859);
or U24356 (N_24356,N_23746,N_23908);
nor U24357 (N_24357,N_23185,N_23810);
xnor U24358 (N_24358,N_23412,N_23105);
or U24359 (N_24359,N_23559,N_23881);
nor U24360 (N_24360,N_23279,N_23652);
and U24361 (N_24361,N_23102,N_23450);
xnor U24362 (N_24362,N_23778,N_23967);
xor U24363 (N_24363,N_23051,N_23216);
or U24364 (N_24364,N_23331,N_23977);
xor U24365 (N_24365,N_23044,N_23028);
nor U24366 (N_24366,N_23196,N_23722);
nor U24367 (N_24367,N_23990,N_23392);
xor U24368 (N_24368,N_23845,N_23751);
or U24369 (N_24369,N_23377,N_23457);
nand U24370 (N_24370,N_23549,N_23246);
nor U24371 (N_24371,N_23864,N_23591);
nor U24372 (N_24372,N_23572,N_23460);
or U24373 (N_24373,N_23923,N_23109);
nor U24374 (N_24374,N_23119,N_23112);
nor U24375 (N_24375,N_23471,N_23709);
and U24376 (N_24376,N_23699,N_23197);
nor U24377 (N_24377,N_23159,N_23920);
and U24378 (N_24378,N_23899,N_23317);
and U24379 (N_24379,N_23470,N_23046);
xor U24380 (N_24380,N_23342,N_23357);
and U24381 (N_24381,N_23334,N_23999);
or U24382 (N_24382,N_23208,N_23199);
or U24383 (N_24383,N_23223,N_23790);
or U24384 (N_24384,N_23129,N_23354);
nor U24385 (N_24385,N_23800,N_23827);
nor U24386 (N_24386,N_23838,N_23431);
nand U24387 (N_24387,N_23567,N_23641);
xor U24388 (N_24388,N_23373,N_23932);
or U24389 (N_24389,N_23618,N_23244);
nor U24390 (N_24390,N_23655,N_23151);
xor U24391 (N_24391,N_23189,N_23594);
or U24392 (N_24392,N_23032,N_23547);
xor U24393 (N_24393,N_23191,N_23325);
or U24394 (N_24394,N_23374,N_23393);
nor U24395 (N_24395,N_23126,N_23569);
xor U24396 (N_24396,N_23250,N_23884);
or U24397 (N_24397,N_23630,N_23520);
nand U24398 (N_24398,N_23496,N_23604);
or U24399 (N_24399,N_23429,N_23703);
or U24400 (N_24400,N_23518,N_23060);
and U24401 (N_24401,N_23409,N_23885);
nor U24402 (N_24402,N_23629,N_23155);
or U24403 (N_24403,N_23850,N_23963);
xnor U24404 (N_24404,N_23420,N_23416);
or U24405 (N_24405,N_23186,N_23352);
xnor U24406 (N_24406,N_23178,N_23814);
and U24407 (N_24407,N_23987,N_23707);
nor U24408 (N_24408,N_23222,N_23006);
and U24409 (N_24409,N_23764,N_23667);
nand U24410 (N_24410,N_23240,N_23114);
xnor U24411 (N_24411,N_23312,N_23791);
nand U24412 (N_24412,N_23837,N_23997);
or U24413 (N_24413,N_23656,N_23818);
or U24414 (N_24414,N_23539,N_23645);
nand U24415 (N_24415,N_23437,N_23693);
nand U24416 (N_24416,N_23832,N_23038);
or U24417 (N_24417,N_23428,N_23115);
xnor U24418 (N_24418,N_23825,N_23517);
and U24419 (N_24419,N_23603,N_23989);
nand U24420 (N_24420,N_23662,N_23104);
and U24421 (N_24421,N_23415,N_23732);
nor U24422 (N_24422,N_23831,N_23033);
and U24423 (N_24423,N_23787,N_23801);
xor U24424 (N_24424,N_23851,N_23650);
xor U24425 (N_24425,N_23107,N_23713);
xnor U24426 (N_24426,N_23804,N_23807);
xnor U24427 (N_24427,N_23363,N_23167);
nand U24428 (N_24428,N_23755,N_23979);
nor U24429 (N_24429,N_23672,N_23448);
nand U24430 (N_24430,N_23389,N_23001);
and U24431 (N_24431,N_23938,N_23130);
or U24432 (N_24432,N_23184,N_23682);
nand U24433 (N_24433,N_23912,N_23919);
nand U24434 (N_24434,N_23615,N_23775);
nor U24435 (N_24435,N_23789,N_23170);
xnor U24436 (N_24436,N_23753,N_23875);
xnor U24437 (N_24437,N_23050,N_23983);
nand U24438 (N_24438,N_23624,N_23612);
nand U24439 (N_24439,N_23436,N_23203);
xnor U24440 (N_24440,N_23822,N_23201);
nand U24441 (N_24441,N_23236,N_23164);
nor U24442 (N_24442,N_23777,N_23843);
nand U24443 (N_24443,N_23454,N_23016);
and U24444 (N_24444,N_23080,N_23293);
or U24445 (N_24445,N_23239,N_23301);
nor U24446 (N_24446,N_23180,N_23324);
xor U24447 (N_24447,N_23233,N_23336);
and U24448 (N_24448,N_23582,N_23960);
or U24449 (N_24449,N_23762,N_23488);
and U24450 (N_24450,N_23555,N_23865);
nor U24451 (N_24451,N_23739,N_23490);
nand U24452 (N_24452,N_23993,N_23358);
nand U24453 (N_24453,N_23714,N_23617);
xor U24454 (N_24454,N_23310,N_23642);
xnor U24455 (N_24455,N_23971,N_23229);
and U24456 (N_24456,N_23782,N_23078);
or U24457 (N_24457,N_23348,N_23291);
and U24458 (N_24458,N_23205,N_23259);
and U24459 (N_24459,N_23345,N_23973);
nor U24460 (N_24460,N_23931,N_23943);
and U24461 (N_24461,N_23307,N_23122);
xor U24462 (N_24462,N_23519,N_23146);
nor U24463 (N_24463,N_23162,N_23290);
and U24464 (N_24464,N_23846,N_23636);
xnor U24465 (N_24465,N_23332,N_23261);
nand U24466 (N_24466,N_23422,N_23173);
nand U24467 (N_24467,N_23194,N_23475);
nand U24468 (N_24468,N_23893,N_23716);
nor U24469 (N_24469,N_23256,N_23945);
and U24470 (N_24470,N_23944,N_23574);
or U24471 (N_24471,N_23949,N_23562);
nand U24472 (N_24472,N_23780,N_23956);
or U24473 (N_24473,N_23319,N_23106);
nor U24474 (N_24474,N_23914,N_23503);
nand U24475 (N_24475,N_23128,N_23917);
or U24476 (N_24476,N_23635,N_23273);
and U24477 (N_24477,N_23796,N_23432);
and U24478 (N_24478,N_23898,N_23740);
or U24479 (N_24479,N_23376,N_23658);
nor U24480 (N_24480,N_23896,N_23444);
nor U24481 (N_24481,N_23004,N_23998);
nor U24482 (N_24482,N_23995,N_23735);
nand U24483 (N_24483,N_23554,N_23387);
nor U24484 (N_24484,N_23364,N_23088);
nand U24485 (N_24485,N_23207,N_23647);
xor U24486 (N_24486,N_23035,N_23527);
nor U24487 (N_24487,N_23954,N_23608);
and U24488 (N_24488,N_23224,N_23563);
nor U24489 (N_24489,N_23402,N_23314);
and U24490 (N_24490,N_23090,N_23278);
and U24491 (N_24491,N_23483,N_23074);
or U24492 (N_24492,N_23476,N_23587);
nand U24493 (N_24493,N_23172,N_23411);
and U24494 (N_24494,N_23145,N_23704);
nand U24495 (N_24495,N_23690,N_23101);
xnor U24496 (N_24496,N_23712,N_23175);
nor U24497 (N_24497,N_23227,N_23673);
or U24498 (N_24498,N_23021,N_23906);
nor U24499 (N_24499,N_23597,N_23474);
nor U24500 (N_24500,N_23349,N_23253);
xnor U24501 (N_24501,N_23844,N_23077);
nor U24502 (N_24502,N_23776,N_23041);
and U24503 (N_24503,N_23963,N_23967);
nand U24504 (N_24504,N_23456,N_23313);
or U24505 (N_24505,N_23301,N_23914);
and U24506 (N_24506,N_23254,N_23152);
nor U24507 (N_24507,N_23697,N_23866);
or U24508 (N_24508,N_23163,N_23015);
nor U24509 (N_24509,N_23153,N_23236);
or U24510 (N_24510,N_23760,N_23710);
and U24511 (N_24511,N_23557,N_23961);
and U24512 (N_24512,N_23023,N_23400);
nor U24513 (N_24513,N_23131,N_23421);
nand U24514 (N_24514,N_23333,N_23078);
or U24515 (N_24515,N_23374,N_23104);
or U24516 (N_24516,N_23909,N_23704);
nor U24517 (N_24517,N_23115,N_23536);
or U24518 (N_24518,N_23230,N_23786);
or U24519 (N_24519,N_23598,N_23625);
xnor U24520 (N_24520,N_23611,N_23974);
nand U24521 (N_24521,N_23894,N_23582);
xor U24522 (N_24522,N_23845,N_23940);
nor U24523 (N_24523,N_23728,N_23351);
nand U24524 (N_24524,N_23134,N_23542);
and U24525 (N_24525,N_23759,N_23721);
or U24526 (N_24526,N_23872,N_23382);
nand U24527 (N_24527,N_23427,N_23209);
nand U24528 (N_24528,N_23981,N_23223);
or U24529 (N_24529,N_23180,N_23593);
nand U24530 (N_24530,N_23028,N_23144);
or U24531 (N_24531,N_23127,N_23116);
and U24532 (N_24532,N_23667,N_23133);
nand U24533 (N_24533,N_23458,N_23280);
or U24534 (N_24534,N_23223,N_23501);
and U24535 (N_24535,N_23611,N_23608);
or U24536 (N_24536,N_23289,N_23598);
and U24537 (N_24537,N_23533,N_23908);
xor U24538 (N_24538,N_23607,N_23775);
and U24539 (N_24539,N_23578,N_23799);
xnor U24540 (N_24540,N_23047,N_23535);
and U24541 (N_24541,N_23658,N_23806);
nor U24542 (N_24542,N_23975,N_23550);
nor U24543 (N_24543,N_23818,N_23012);
or U24544 (N_24544,N_23061,N_23865);
and U24545 (N_24545,N_23045,N_23286);
nor U24546 (N_24546,N_23187,N_23466);
nor U24547 (N_24547,N_23426,N_23266);
nand U24548 (N_24548,N_23514,N_23381);
nor U24549 (N_24549,N_23969,N_23734);
or U24550 (N_24550,N_23576,N_23525);
nor U24551 (N_24551,N_23820,N_23307);
nand U24552 (N_24552,N_23753,N_23181);
nand U24553 (N_24553,N_23329,N_23035);
and U24554 (N_24554,N_23376,N_23565);
xor U24555 (N_24555,N_23025,N_23159);
nand U24556 (N_24556,N_23590,N_23375);
or U24557 (N_24557,N_23453,N_23979);
or U24558 (N_24558,N_23725,N_23415);
or U24559 (N_24559,N_23701,N_23727);
or U24560 (N_24560,N_23728,N_23979);
nor U24561 (N_24561,N_23025,N_23100);
or U24562 (N_24562,N_23560,N_23459);
nor U24563 (N_24563,N_23802,N_23580);
nand U24564 (N_24564,N_23897,N_23553);
nor U24565 (N_24565,N_23239,N_23266);
or U24566 (N_24566,N_23076,N_23883);
nor U24567 (N_24567,N_23096,N_23097);
xor U24568 (N_24568,N_23153,N_23326);
xor U24569 (N_24569,N_23028,N_23981);
or U24570 (N_24570,N_23931,N_23172);
nor U24571 (N_24571,N_23791,N_23187);
xnor U24572 (N_24572,N_23556,N_23930);
or U24573 (N_24573,N_23586,N_23867);
nand U24574 (N_24574,N_23552,N_23449);
and U24575 (N_24575,N_23827,N_23445);
nand U24576 (N_24576,N_23620,N_23812);
and U24577 (N_24577,N_23759,N_23331);
or U24578 (N_24578,N_23768,N_23062);
nand U24579 (N_24579,N_23716,N_23052);
and U24580 (N_24580,N_23752,N_23524);
or U24581 (N_24581,N_23694,N_23389);
and U24582 (N_24582,N_23837,N_23504);
and U24583 (N_24583,N_23424,N_23059);
and U24584 (N_24584,N_23963,N_23323);
or U24585 (N_24585,N_23088,N_23044);
nor U24586 (N_24586,N_23679,N_23643);
nor U24587 (N_24587,N_23872,N_23169);
nand U24588 (N_24588,N_23500,N_23897);
nor U24589 (N_24589,N_23640,N_23763);
and U24590 (N_24590,N_23502,N_23327);
or U24591 (N_24591,N_23302,N_23282);
nor U24592 (N_24592,N_23669,N_23299);
nand U24593 (N_24593,N_23731,N_23159);
nor U24594 (N_24594,N_23029,N_23852);
or U24595 (N_24595,N_23704,N_23710);
xnor U24596 (N_24596,N_23177,N_23738);
nor U24597 (N_24597,N_23987,N_23174);
or U24598 (N_24598,N_23588,N_23666);
and U24599 (N_24599,N_23671,N_23663);
nand U24600 (N_24600,N_23562,N_23907);
and U24601 (N_24601,N_23569,N_23028);
xor U24602 (N_24602,N_23347,N_23671);
nand U24603 (N_24603,N_23330,N_23128);
nor U24604 (N_24604,N_23788,N_23279);
nor U24605 (N_24605,N_23204,N_23870);
nor U24606 (N_24606,N_23702,N_23692);
nand U24607 (N_24607,N_23038,N_23437);
nand U24608 (N_24608,N_23502,N_23401);
nand U24609 (N_24609,N_23339,N_23184);
xnor U24610 (N_24610,N_23780,N_23059);
nor U24611 (N_24611,N_23529,N_23280);
xnor U24612 (N_24612,N_23785,N_23700);
nor U24613 (N_24613,N_23337,N_23972);
nand U24614 (N_24614,N_23450,N_23524);
and U24615 (N_24615,N_23756,N_23717);
or U24616 (N_24616,N_23086,N_23842);
nor U24617 (N_24617,N_23378,N_23538);
and U24618 (N_24618,N_23095,N_23667);
or U24619 (N_24619,N_23288,N_23883);
xnor U24620 (N_24620,N_23145,N_23029);
nor U24621 (N_24621,N_23685,N_23936);
nand U24622 (N_24622,N_23287,N_23914);
nor U24623 (N_24623,N_23380,N_23877);
nor U24624 (N_24624,N_23738,N_23473);
and U24625 (N_24625,N_23092,N_23166);
nand U24626 (N_24626,N_23977,N_23138);
nand U24627 (N_24627,N_23949,N_23417);
xor U24628 (N_24628,N_23253,N_23088);
nand U24629 (N_24629,N_23380,N_23297);
nand U24630 (N_24630,N_23604,N_23800);
nor U24631 (N_24631,N_23813,N_23049);
nor U24632 (N_24632,N_23872,N_23516);
xnor U24633 (N_24633,N_23551,N_23151);
nor U24634 (N_24634,N_23123,N_23256);
nand U24635 (N_24635,N_23252,N_23839);
xnor U24636 (N_24636,N_23973,N_23364);
or U24637 (N_24637,N_23633,N_23258);
or U24638 (N_24638,N_23485,N_23125);
xnor U24639 (N_24639,N_23531,N_23552);
xor U24640 (N_24640,N_23934,N_23552);
nand U24641 (N_24641,N_23914,N_23906);
or U24642 (N_24642,N_23441,N_23963);
or U24643 (N_24643,N_23832,N_23531);
and U24644 (N_24644,N_23430,N_23194);
nor U24645 (N_24645,N_23832,N_23789);
xnor U24646 (N_24646,N_23896,N_23801);
and U24647 (N_24647,N_23476,N_23974);
nor U24648 (N_24648,N_23265,N_23679);
and U24649 (N_24649,N_23288,N_23845);
and U24650 (N_24650,N_23920,N_23544);
nand U24651 (N_24651,N_23121,N_23599);
and U24652 (N_24652,N_23230,N_23091);
xor U24653 (N_24653,N_23735,N_23912);
or U24654 (N_24654,N_23706,N_23099);
and U24655 (N_24655,N_23290,N_23137);
nor U24656 (N_24656,N_23496,N_23682);
or U24657 (N_24657,N_23262,N_23789);
xnor U24658 (N_24658,N_23906,N_23810);
or U24659 (N_24659,N_23053,N_23069);
nand U24660 (N_24660,N_23712,N_23986);
or U24661 (N_24661,N_23144,N_23959);
nand U24662 (N_24662,N_23665,N_23230);
and U24663 (N_24663,N_23053,N_23494);
xor U24664 (N_24664,N_23790,N_23264);
nand U24665 (N_24665,N_23641,N_23880);
nor U24666 (N_24666,N_23295,N_23533);
nor U24667 (N_24667,N_23120,N_23872);
nand U24668 (N_24668,N_23607,N_23783);
nand U24669 (N_24669,N_23950,N_23564);
nor U24670 (N_24670,N_23995,N_23025);
nor U24671 (N_24671,N_23458,N_23386);
and U24672 (N_24672,N_23786,N_23795);
and U24673 (N_24673,N_23652,N_23879);
xor U24674 (N_24674,N_23246,N_23731);
nor U24675 (N_24675,N_23250,N_23262);
or U24676 (N_24676,N_23569,N_23854);
nand U24677 (N_24677,N_23705,N_23794);
and U24678 (N_24678,N_23073,N_23621);
and U24679 (N_24679,N_23420,N_23037);
and U24680 (N_24680,N_23426,N_23371);
or U24681 (N_24681,N_23324,N_23772);
nand U24682 (N_24682,N_23766,N_23675);
nand U24683 (N_24683,N_23622,N_23448);
and U24684 (N_24684,N_23819,N_23330);
and U24685 (N_24685,N_23903,N_23690);
xor U24686 (N_24686,N_23168,N_23340);
and U24687 (N_24687,N_23651,N_23971);
and U24688 (N_24688,N_23220,N_23134);
nor U24689 (N_24689,N_23061,N_23298);
or U24690 (N_24690,N_23287,N_23102);
nor U24691 (N_24691,N_23956,N_23829);
nor U24692 (N_24692,N_23641,N_23699);
and U24693 (N_24693,N_23506,N_23423);
or U24694 (N_24694,N_23357,N_23437);
and U24695 (N_24695,N_23910,N_23450);
or U24696 (N_24696,N_23340,N_23325);
or U24697 (N_24697,N_23625,N_23430);
and U24698 (N_24698,N_23339,N_23213);
and U24699 (N_24699,N_23778,N_23207);
nand U24700 (N_24700,N_23262,N_23718);
xor U24701 (N_24701,N_23970,N_23460);
and U24702 (N_24702,N_23268,N_23790);
xnor U24703 (N_24703,N_23904,N_23706);
and U24704 (N_24704,N_23440,N_23420);
nor U24705 (N_24705,N_23091,N_23697);
nand U24706 (N_24706,N_23048,N_23021);
nand U24707 (N_24707,N_23902,N_23553);
nor U24708 (N_24708,N_23010,N_23358);
xor U24709 (N_24709,N_23308,N_23321);
or U24710 (N_24710,N_23598,N_23680);
nand U24711 (N_24711,N_23070,N_23490);
nor U24712 (N_24712,N_23918,N_23110);
nor U24713 (N_24713,N_23311,N_23659);
or U24714 (N_24714,N_23002,N_23222);
xnor U24715 (N_24715,N_23753,N_23466);
nor U24716 (N_24716,N_23554,N_23983);
or U24717 (N_24717,N_23503,N_23042);
nor U24718 (N_24718,N_23612,N_23408);
or U24719 (N_24719,N_23421,N_23512);
nand U24720 (N_24720,N_23881,N_23783);
or U24721 (N_24721,N_23757,N_23912);
or U24722 (N_24722,N_23128,N_23802);
nand U24723 (N_24723,N_23785,N_23666);
nand U24724 (N_24724,N_23460,N_23160);
and U24725 (N_24725,N_23338,N_23453);
nand U24726 (N_24726,N_23233,N_23519);
and U24727 (N_24727,N_23847,N_23775);
and U24728 (N_24728,N_23144,N_23346);
xor U24729 (N_24729,N_23684,N_23389);
xnor U24730 (N_24730,N_23771,N_23525);
or U24731 (N_24731,N_23510,N_23048);
and U24732 (N_24732,N_23882,N_23096);
nand U24733 (N_24733,N_23583,N_23649);
and U24734 (N_24734,N_23158,N_23280);
or U24735 (N_24735,N_23760,N_23125);
nor U24736 (N_24736,N_23189,N_23862);
or U24737 (N_24737,N_23501,N_23187);
or U24738 (N_24738,N_23420,N_23604);
nor U24739 (N_24739,N_23906,N_23363);
nand U24740 (N_24740,N_23599,N_23719);
and U24741 (N_24741,N_23533,N_23828);
nor U24742 (N_24742,N_23502,N_23573);
xor U24743 (N_24743,N_23762,N_23117);
nor U24744 (N_24744,N_23821,N_23146);
and U24745 (N_24745,N_23460,N_23693);
nor U24746 (N_24746,N_23822,N_23595);
and U24747 (N_24747,N_23992,N_23385);
nand U24748 (N_24748,N_23461,N_23376);
xnor U24749 (N_24749,N_23116,N_23024);
xnor U24750 (N_24750,N_23701,N_23762);
and U24751 (N_24751,N_23838,N_23740);
nand U24752 (N_24752,N_23776,N_23160);
nor U24753 (N_24753,N_23201,N_23807);
nand U24754 (N_24754,N_23400,N_23727);
or U24755 (N_24755,N_23453,N_23362);
or U24756 (N_24756,N_23127,N_23829);
and U24757 (N_24757,N_23711,N_23854);
and U24758 (N_24758,N_23064,N_23469);
and U24759 (N_24759,N_23759,N_23271);
or U24760 (N_24760,N_23255,N_23835);
xnor U24761 (N_24761,N_23557,N_23267);
xor U24762 (N_24762,N_23784,N_23427);
and U24763 (N_24763,N_23113,N_23912);
nand U24764 (N_24764,N_23556,N_23889);
nand U24765 (N_24765,N_23378,N_23963);
or U24766 (N_24766,N_23605,N_23875);
xor U24767 (N_24767,N_23678,N_23430);
xnor U24768 (N_24768,N_23944,N_23966);
xnor U24769 (N_24769,N_23044,N_23167);
xor U24770 (N_24770,N_23038,N_23050);
nand U24771 (N_24771,N_23348,N_23199);
xnor U24772 (N_24772,N_23687,N_23590);
nand U24773 (N_24773,N_23696,N_23935);
nand U24774 (N_24774,N_23152,N_23856);
nand U24775 (N_24775,N_23191,N_23253);
and U24776 (N_24776,N_23973,N_23769);
nand U24777 (N_24777,N_23252,N_23302);
xnor U24778 (N_24778,N_23604,N_23560);
nand U24779 (N_24779,N_23439,N_23690);
nor U24780 (N_24780,N_23134,N_23286);
nand U24781 (N_24781,N_23927,N_23025);
nor U24782 (N_24782,N_23131,N_23357);
or U24783 (N_24783,N_23134,N_23236);
and U24784 (N_24784,N_23881,N_23493);
nor U24785 (N_24785,N_23747,N_23978);
xor U24786 (N_24786,N_23439,N_23383);
or U24787 (N_24787,N_23599,N_23532);
nand U24788 (N_24788,N_23222,N_23715);
xnor U24789 (N_24789,N_23308,N_23208);
nand U24790 (N_24790,N_23519,N_23591);
nor U24791 (N_24791,N_23175,N_23456);
or U24792 (N_24792,N_23187,N_23492);
xnor U24793 (N_24793,N_23876,N_23816);
xnor U24794 (N_24794,N_23181,N_23379);
nor U24795 (N_24795,N_23528,N_23984);
nand U24796 (N_24796,N_23224,N_23596);
nor U24797 (N_24797,N_23866,N_23002);
nand U24798 (N_24798,N_23702,N_23858);
nand U24799 (N_24799,N_23690,N_23766);
or U24800 (N_24800,N_23059,N_23364);
nor U24801 (N_24801,N_23397,N_23548);
nand U24802 (N_24802,N_23030,N_23628);
nand U24803 (N_24803,N_23434,N_23569);
and U24804 (N_24804,N_23536,N_23031);
xor U24805 (N_24805,N_23286,N_23476);
nand U24806 (N_24806,N_23815,N_23582);
xnor U24807 (N_24807,N_23231,N_23314);
and U24808 (N_24808,N_23194,N_23566);
nor U24809 (N_24809,N_23131,N_23132);
xor U24810 (N_24810,N_23256,N_23592);
and U24811 (N_24811,N_23707,N_23102);
nor U24812 (N_24812,N_23303,N_23897);
nor U24813 (N_24813,N_23432,N_23226);
xor U24814 (N_24814,N_23726,N_23946);
or U24815 (N_24815,N_23895,N_23133);
xor U24816 (N_24816,N_23133,N_23785);
nand U24817 (N_24817,N_23671,N_23643);
or U24818 (N_24818,N_23130,N_23893);
xor U24819 (N_24819,N_23443,N_23407);
xnor U24820 (N_24820,N_23618,N_23648);
xor U24821 (N_24821,N_23407,N_23746);
nand U24822 (N_24822,N_23212,N_23342);
and U24823 (N_24823,N_23227,N_23686);
and U24824 (N_24824,N_23493,N_23332);
and U24825 (N_24825,N_23634,N_23969);
nand U24826 (N_24826,N_23592,N_23060);
and U24827 (N_24827,N_23121,N_23301);
xor U24828 (N_24828,N_23149,N_23809);
and U24829 (N_24829,N_23220,N_23468);
nand U24830 (N_24830,N_23751,N_23828);
nand U24831 (N_24831,N_23693,N_23574);
and U24832 (N_24832,N_23501,N_23571);
and U24833 (N_24833,N_23383,N_23077);
nor U24834 (N_24834,N_23316,N_23645);
and U24835 (N_24835,N_23719,N_23137);
nand U24836 (N_24836,N_23916,N_23230);
nor U24837 (N_24837,N_23075,N_23985);
nand U24838 (N_24838,N_23306,N_23148);
xnor U24839 (N_24839,N_23302,N_23670);
or U24840 (N_24840,N_23440,N_23004);
or U24841 (N_24841,N_23292,N_23401);
or U24842 (N_24842,N_23807,N_23338);
and U24843 (N_24843,N_23353,N_23268);
or U24844 (N_24844,N_23741,N_23986);
and U24845 (N_24845,N_23046,N_23845);
or U24846 (N_24846,N_23579,N_23619);
and U24847 (N_24847,N_23646,N_23326);
nand U24848 (N_24848,N_23014,N_23941);
or U24849 (N_24849,N_23785,N_23869);
xor U24850 (N_24850,N_23550,N_23611);
nand U24851 (N_24851,N_23726,N_23448);
or U24852 (N_24852,N_23768,N_23405);
xor U24853 (N_24853,N_23064,N_23870);
nor U24854 (N_24854,N_23636,N_23588);
nand U24855 (N_24855,N_23374,N_23454);
xor U24856 (N_24856,N_23725,N_23914);
nand U24857 (N_24857,N_23086,N_23641);
nor U24858 (N_24858,N_23996,N_23778);
or U24859 (N_24859,N_23737,N_23658);
or U24860 (N_24860,N_23709,N_23410);
and U24861 (N_24861,N_23925,N_23968);
and U24862 (N_24862,N_23683,N_23881);
nand U24863 (N_24863,N_23182,N_23192);
or U24864 (N_24864,N_23325,N_23332);
xnor U24865 (N_24865,N_23529,N_23354);
xor U24866 (N_24866,N_23712,N_23864);
xor U24867 (N_24867,N_23797,N_23371);
and U24868 (N_24868,N_23215,N_23227);
xnor U24869 (N_24869,N_23280,N_23941);
and U24870 (N_24870,N_23311,N_23613);
or U24871 (N_24871,N_23783,N_23798);
nand U24872 (N_24872,N_23968,N_23391);
xor U24873 (N_24873,N_23501,N_23085);
or U24874 (N_24874,N_23073,N_23852);
or U24875 (N_24875,N_23247,N_23201);
and U24876 (N_24876,N_23030,N_23684);
and U24877 (N_24877,N_23500,N_23380);
nor U24878 (N_24878,N_23688,N_23434);
nor U24879 (N_24879,N_23673,N_23656);
nor U24880 (N_24880,N_23161,N_23345);
or U24881 (N_24881,N_23767,N_23837);
nor U24882 (N_24882,N_23159,N_23147);
nand U24883 (N_24883,N_23470,N_23347);
nor U24884 (N_24884,N_23536,N_23468);
nor U24885 (N_24885,N_23170,N_23134);
and U24886 (N_24886,N_23878,N_23511);
or U24887 (N_24887,N_23945,N_23201);
nand U24888 (N_24888,N_23502,N_23653);
xnor U24889 (N_24889,N_23031,N_23118);
nor U24890 (N_24890,N_23442,N_23289);
or U24891 (N_24891,N_23815,N_23553);
or U24892 (N_24892,N_23408,N_23595);
xnor U24893 (N_24893,N_23241,N_23484);
and U24894 (N_24894,N_23134,N_23300);
nor U24895 (N_24895,N_23116,N_23672);
nand U24896 (N_24896,N_23876,N_23005);
nor U24897 (N_24897,N_23364,N_23079);
nand U24898 (N_24898,N_23716,N_23939);
xor U24899 (N_24899,N_23848,N_23315);
and U24900 (N_24900,N_23574,N_23723);
nor U24901 (N_24901,N_23222,N_23614);
or U24902 (N_24902,N_23022,N_23477);
nor U24903 (N_24903,N_23885,N_23538);
nor U24904 (N_24904,N_23550,N_23720);
nand U24905 (N_24905,N_23425,N_23973);
or U24906 (N_24906,N_23380,N_23333);
nand U24907 (N_24907,N_23706,N_23246);
nand U24908 (N_24908,N_23542,N_23923);
nor U24909 (N_24909,N_23942,N_23422);
and U24910 (N_24910,N_23365,N_23349);
and U24911 (N_24911,N_23529,N_23602);
xor U24912 (N_24912,N_23949,N_23902);
and U24913 (N_24913,N_23805,N_23020);
or U24914 (N_24914,N_23228,N_23777);
or U24915 (N_24915,N_23260,N_23961);
nor U24916 (N_24916,N_23936,N_23412);
and U24917 (N_24917,N_23327,N_23680);
nor U24918 (N_24918,N_23002,N_23161);
nor U24919 (N_24919,N_23927,N_23241);
and U24920 (N_24920,N_23701,N_23188);
xnor U24921 (N_24921,N_23578,N_23221);
nand U24922 (N_24922,N_23599,N_23826);
and U24923 (N_24923,N_23738,N_23516);
nor U24924 (N_24924,N_23591,N_23081);
nand U24925 (N_24925,N_23131,N_23986);
xor U24926 (N_24926,N_23841,N_23878);
xnor U24927 (N_24927,N_23777,N_23392);
nor U24928 (N_24928,N_23632,N_23901);
xnor U24929 (N_24929,N_23013,N_23710);
or U24930 (N_24930,N_23247,N_23009);
nor U24931 (N_24931,N_23646,N_23451);
xor U24932 (N_24932,N_23035,N_23008);
nor U24933 (N_24933,N_23068,N_23844);
and U24934 (N_24934,N_23725,N_23578);
or U24935 (N_24935,N_23012,N_23898);
nor U24936 (N_24936,N_23992,N_23048);
nand U24937 (N_24937,N_23259,N_23680);
xor U24938 (N_24938,N_23808,N_23153);
nand U24939 (N_24939,N_23097,N_23090);
xnor U24940 (N_24940,N_23813,N_23084);
nor U24941 (N_24941,N_23798,N_23541);
xnor U24942 (N_24942,N_23862,N_23422);
or U24943 (N_24943,N_23969,N_23257);
or U24944 (N_24944,N_23643,N_23932);
nor U24945 (N_24945,N_23066,N_23365);
nor U24946 (N_24946,N_23712,N_23847);
nor U24947 (N_24947,N_23729,N_23351);
xnor U24948 (N_24948,N_23221,N_23012);
xor U24949 (N_24949,N_23321,N_23201);
xnor U24950 (N_24950,N_23811,N_23545);
nor U24951 (N_24951,N_23799,N_23115);
nand U24952 (N_24952,N_23844,N_23341);
and U24953 (N_24953,N_23342,N_23873);
nand U24954 (N_24954,N_23192,N_23549);
nand U24955 (N_24955,N_23108,N_23365);
nor U24956 (N_24956,N_23075,N_23754);
or U24957 (N_24957,N_23359,N_23309);
or U24958 (N_24958,N_23281,N_23235);
nand U24959 (N_24959,N_23625,N_23668);
and U24960 (N_24960,N_23696,N_23248);
xnor U24961 (N_24961,N_23353,N_23398);
xor U24962 (N_24962,N_23160,N_23175);
nand U24963 (N_24963,N_23407,N_23963);
nor U24964 (N_24964,N_23251,N_23516);
nand U24965 (N_24965,N_23119,N_23207);
or U24966 (N_24966,N_23758,N_23820);
or U24967 (N_24967,N_23593,N_23740);
or U24968 (N_24968,N_23660,N_23262);
nand U24969 (N_24969,N_23052,N_23009);
xnor U24970 (N_24970,N_23044,N_23837);
xor U24971 (N_24971,N_23071,N_23110);
nor U24972 (N_24972,N_23476,N_23149);
xnor U24973 (N_24973,N_23733,N_23429);
nor U24974 (N_24974,N_23339,N_23727);
or U24975 (N_24975,N_23914,N_23865);
nor U24976 (N_24976,N_23090,N_23733);
nand U24977 (N_24977,N_23707,N_23241);
nand U24978 (N_24978,N_23311,N_23798);
nand U24979 (N_24979,N_23403,N_23189);
nand U24980 (N_24980,N_23979,N_23113);
nor U24981 (N_24981,N_23393,N_23356);
xor U24982 (N_24982,N_23421,N_23097);
nor U24983 (N_24983,N_23117,N_23376);
nand U24984 (N_24984,N_23112,N_23109);
nor U24985 (N_24985,N_23929,N_23251);
and U24986 (N_24986,N_23505,N_23952);
or U24987 (N_24987,N_23875,N_23488);
and U24988 (N_24988,N_23128,N_23954);
nor U24989 (N_24989,N_23046,N_23348);
and U24990 (N_24990,N_23316,N_23970);
and U24991 (N_24991,N_23641,N_23342);
nand U24992 (N_24992,N_23246,N_23735);
and U24993 (N_24993,N_23231,N_23012);
or U24994 (N_24994,N_23458,N_23598);
xor U24995 (N_24995,N_23412,N_23000);
or U24996 (N_24996,N_23796,N_23771);
or U24997 (N_24997,N_23396,N_23896);
nor U24998 (N_24998,N_23393,N_23383);
nor U24999 (N_24999,N_23087,N_23393);
nand U25000 (N_25000,N_24802,N_24400);
nor U25001 (N_25001,N_24796,N_24900);
or U25002 (N_25002,N_24511,N_24307);
and U25003 (N_25003,N_24002,N_24493);
xor U25004 (N_25004,N_24490,N_24685);
or U25005 (N_25005,N_24418,N_24079);
xor U25006 (N_25006,N_24394,N_24144);
and U25007 (N_25007,N_24173,N_24043);
and U25008 (N_25008,N_24067,N_24944);
nand U25009 (N_25009,N_24482,N_24617);
and U25010 (N_25010,N_24666,N_24941);
and U25011 (N_25011,N_24724,N_24407);
nand U25012 (N_25012,N_24773,N_24643);
xor U25013 (N_25013,N_24833,N_24164);
or U25014 (N_25014,N_24360,N_24132);
nor U25015 (N_25015,N_24001,N_24426);
and U25016 (N_25016,N_24662,N_24836);
or U25017 (N_25017,N_24105,N_24580);
xor U25018 (N_25018,N_24024,N_24764);
xor U25019 (N_25019,N_24533,N_24838);
xor U25020 (N_25020,N_24985,N_24851);
and U25021 (N_25021,N_24453,N_24992);
nand U25022 (N_25022,N_24478,N_24325);
xnor U25023 (N_25023,N_24709,N_24066);
nand U25024 (N_25024,N_24183,N_24835);
nor U25025 (N_25025,N_24807,N_24540);
nand U25026 (N_25026,N_24410,N_24744);
nand U25027 (N_25027,N_24255,N_24711);
nand U25028 (N_25028,N_24938,N_24800);
and U25029 (N_25029,N_24669,N_24191);
or U25030 (N_25030,N_24266,N_24808);
xnor U25031 (N_25031,N_24752,N_24675);
nand U25032 (N_25032,N_24054,N_24126);
or U25033 (N_25033,N_24009,N_24015);
nor U25034 (N_25034,N_24073,N_24747);
xnor U25035 (N_25035,N_24033,N_24931);
nor U25036 (N_25036,N_24756,N_24981);
xor U25037 (N_25037,N_24775,N_24157);
nand U25038 (N_25038,N_24353,N_24000);
nand U25039 (N_25039,N_24719,N_24821);
nor U25040 (N_25040,N_24894,N_24253);
nor U25041 (N_25041,N_24055,N_24184);
nand U25042 (N_25042,N_24668,N_24012);
and U25043 (N_25043,N_24960,N_24403);
xor U25044 (N_25044,N_24624,N_24117);
or U25045 (N_25045,N_24673,N_24094);
and U25046 (N_25046,N_24522,N_24323);
xnor U25047 (N_25047,N_24832,N_24740);
or U25048 (N_25048,N_24954,N_24893);
xor U25049 (N_25049,N_24371,N_24113);
nand U25050 (N_25050,N_24809,N_24574);
or U25051 (N_25051,N_24721,N_24913);
xnor U25052 (N_25052,N_24141,N_24151);
nor U25053 (N_25053,N_24872,N_24538);
or U25054 (N_25054,N_24163,N_24315);
or U25055 (N_25055,N_24007,N_24275);
nor U25056 (N_25056,N_24571,N_24996);
xnor U25057 (N_25057,N_24652,N_24384);
and U25058 (N_25058,N_24646,N_24119);
xnor U25059 (N_25059,N_24973,N_24774);
xnor U25060 (N_25060,N_24084,N_24260);
xor U25061 (N_25061,N_24081,N_24205);
or U25062 (N_25062,N_24280,N_24468);
nand U25063 (N_25063,N_24306,N_24867);
and U25064 (N_25064,N_24993,N_24458);
nor U25065 (N_25065,N_24381,N_24516);
or U25066 (N_25066,N_24211,N_24063);
or U25067 (N_25067,N_24670,N_24612);
nand U25068 (N_25068,N_24915,N_24050);
and U25069 (N_25069,N_24277,N_24559);
xnor U25070 (N_25070,N_24804,N_24534);
nand U25071 (N_25071,N_24602,N_24189);
nand U25072 (N_25072,N_24147,N_24110);
or U25073 (N_25073,N_24292,N_24090);
xor U25074 (N_25074,N_24447,N_24859);
or U25075 (N_25075,N_24928,N_24671);
nand U25076 (N_25076,N_24723,N_24815);
and U25077 (N_25077,N_24657,N_24272);
nor U25078 (N_25078,N_24146,N_24731);
or U25079 (N_25079,N_24061,N_24582);
xor U25080 (N_25080,N_24914,N_24525);
or U25081 (N_25081,N_24820,N_24978);
nor U25082 (N_25082,N_24647,N_24170);
nor U25083 (N_25083,N_24398,N_24907);
and U25084 (N_25084,N_24549,N_24017);
nand U25085 (N_25085,N_24762,N_24888);
xnor U25086 (N_25086,N_24432,N_24518);
nand U25087 (N_25087,N_24923,N_24310);
nand U25088 (N_25088,N_24885,N_24840);
and U25089 (N_25089,N_24142,N_24854);
nor U25090 (N_25090,N_24233,N_24303);
nand U25091 (N_25091,N_24912,N_24890);
xnor U25092 (N_25092,N_24251,N_24342);
or U25093 (N_25093,N_24868,N_24003);
xor U25094 (N_25094,N_24298,N_24413);
nand U25095 (N_25095,N_24720,N_24145);
xnor U25096 (N_25096,N_24466,N_24738);
and U25097 (N_25097,N_24917,N_24240);
xnor U25098 (N_25098,N_24962,N_24334);
or U25099 (N_25099,N_24417,N_24192);
or U25100 (N_25100,N_24464,N_24062);
or U25101 (N_25101,N_24845,N_24299);
nand U25102 (N_25102,N_24812,N_24335);
and U25103 (N_25103,N_24823,N_24567);
xor U25104 (N_25104,N_24419,N_24361);
xnor U25105 (N_25105,N_24399,N_24691);
nor U25106 (N_25106,N_24193,N_24613);
nand U25107 (N_25107,N_24068,N_24302);
nor U25108 (N_25108,N_24218,N_24182);
nor U25109 (N_25109,N_24169,N_24372);
nor U25110 (N_25110,N_24782,N_24391);
and U25111 (N_25111,N_24052,N_24370);
nand U25112 (N_25112,N_24886,N_24769);
or U25113 (N_25113,N_24224,N_24924);
and U25114 (N_25114,N_24064,N_24958);
or U25115 (N_25115,N_24732,N_24593);
nand U25116 (N_25116,N_24876,N_24311);
and U25117 (N_25117,N_24902,N_24265);
nor U25118 (N_25118,N_24368,N_24392);
or U25119 (N_25119,N_24562,N_24891);
nor U25120 (N_25120,N_24947,N_24942);
xor U25121 (N_25121,N_24159,N_24519);
xnor U25122 (N_25122,N_24550,N_24186);
and U25123 (N_25123,N_24349,N_24795);
and U25124 (N_25124,N_24697,N_24611);
nand U25125 (N_25125,N_24268,N_24354);
nand U25126 (N_25126,N_24860,N_24203);
nor U25127 (N_25127,N_24863,N_24585);
nor U25128 (N_25128,N_24529,N_24247);
or U25129 (N_25129,N_24869,N_24929);
and U25130 (N_25130,N_24554,N_24348);
nand U25131 (N_25131,N_24237,N_24539);
nor U25132 (N_25132,N_24507,N_24693);
nor U25133 (N_25133,N_24058,N_24592);
and U25134 (N_25134,N_24296,N_24285);
nand U25135 (N_25135,N_24664,N_24440);
or U25136 (N_25136,N_24856,N_24014);
nor U25137 (N_25137,N_24805,N_24555);
or U25138 (N_25138,N_24979,N_24242);
nand U25139 (N_25139,N_24025,N_24016);
and U25140 (N_25140,N_24143,N_24627);
or U25141 (N_25141,N_24448,N_24698);
or U25142 (N_25142,N_24716,N_24892);
or U25143 (N_25143,N_24499,N_24160);
xnor U25144 (N_25144,N_24128,N_24314);
nor U25145 (N_25145,N_24462,N_24866);
nor U25146 (N_25146,N_24537,N_24383);
nand U25147 (N_25147,N_24730,N_24616);
xor U25148 (N_25148,N_24523,N_24060);
nor U25149 (N_25149,N_24966,N_24379);
nor U25150 (N_25150,N_24544,N_24974);
xor U25151 (N_25151,N_24236,N_24682);
nand U25152 (N_25152,N_24770,N_24998);
nand U25153 (N_25153,N_24753,N_24229);
or U25154 (N_25154,N_24687,N_24284);
or U25155 (N_25155,N_24729,N_24101);
nand U25156 (N_25156,N_24590,N_24431);
nand U25157 (N_25157,N_24297,N_24583);
nor U25158 (N_25158,N_24615,N_24264);
nand U25159 (N_25159,N_24011,N_24267);
xor U25160 (N_25160,N_24994,N_24148);
xnor U25161 (N_25161,N_24827,N_24965);
nand U25162 (N_25162,N_24526,N_24508);
nand U25163 (N_25163,N_24722,N_24563);
or U25164 (N_25164,N_24925,N_24320);
nor U25165 (N_25165,N_24683,N_24609);
nor U25166 (N_25166,N_24428,N_24341);
and U25167 (N_25167,N_24801,N_24834);
nand U25168 (N_25168,N_24543,N_24376);
nor U25169 (N_25169,N_24136,N_24677);
or U25170 (N_25170,N_24622,N_24112);
or U25171 (N_25171,N_24047,N_24674);
nand U25172 (N_25172,N_24395,N_24256);
and U25173 (N_25173,N_24289,N_24576);
and U25174 (N_25174,N_24776,N_24570);
and U25175 (N_25175,N_24234,N_24109);
nand U25176 (N_25176,N_24547,N_24249);
nor U25177 (N_25177,N_24569,N_24742);
and U25178 (N_25178,N_24129,N_24606);
nand U25179 (N_25179,N_24767,N_24287);
or U25180 (N_25180,N_24991,N_24322);
or U25181 (N_25181,N_24291,N_24489);
and U25182 (N_25182,N_24517,N_24990);
nor U25183 (N_25183,N_24995,N_24887);
xor U25184 (N_25184,N_24989,N_24162);
nand U25185 (N_25185,N_24873,N_24288);
nand U25186 (N_25186,N_24934,N_24704);
and U25187 (N_25187,N_24734,N_24103);
and U25188 (N_25188,N_24380,N_24401);
and U25189 (N_25189,N_24034,N_24588);
or U25190 (N_25190,N_24603,N_24975);
or U25191 (N_25191,N_24138,N_24232);
and U25192 (N_25192,N_24107,N_24181);
nor U25193 (N_25193,N_24423,N_24445);
or U25194 (N_25194,N_24479,N_24935);
nor U25195 (N_25195,N_24751,N_24749);
or U25196 (N_25196,N_24359,N_24207);
and U25197 (N_25197,N_24586,N_24022);
and U25198 (N_25198,N_24118,N_24248);
or U25199 (N_25199,N_24694,N_24654);
nor U25200 (N_25200,N_24195,N_24610);
xor U25201 (N_25201,N_24557,N_24948);
xnor U25202 (N_25202,N_24937,N_24373);
or U25203 (N_25203,N_24279,N_24637);
xor U25204 (N_25204,N_24217,N_24779);
nor U25205 (N_25205,N_24435,N_24601);
xnor U25206 (N_25206,N_24757,N_24235);
and U25207 (N_25207,N_24967,N_24792);
nand U25208 (N_25208,N_24366,N_24220);
nor U25209 (N_25209,N_24505,N_24560);
and U25210 (N_25210,N_24471,N_24127);
or U25211 (N_25211,N_24778,N_24653);
or U25212 (N_25212,N_24347,N_24166);
xor U25213 (N_25213,N_24790,N_24841);
and U25214 (N_25214,N_24338,N_24020);
nand U25215 (N_25215,N_24803,N_24623);
nor U25216 (N_25216,N_24281,N_24871);
and U25217 (N_25217,N_24305,N_24048);
and U25218 (N_25218,N_24125,N_24226);
or U25219 (N_25219,N_24187,N_24553);
nor U25220 (N_25220,N_24436,N_24831);
nor U25221 (N_25221,N_24676,N_24945);
xor U25222 (N_25222,N_24329,N_24660);
nor U25223 (N_25223,N_24438,N_24227);
nand U25224 (N_25224,N_24228,N_24843);
nor U25225 (N_25225,N_24857,N_24918);
nor U25226 (N_25226,N_24520,N_24046);
nor U25227 (N_25227,N_24039,N_24455);
or U25228 (N_25228,N_24093,N_24316);
and U25229 (N_25229,N_24568,N_24758);
nor U25230 (N_25230,N_24686,N_24715);
xor U25231 (N_25231,N_24443,N_24339);
xor U25232 (N_25232,N_24707,N_24225);
nor U25233 (N_25233,N_24761,N_24344);
nand U25234 (N_25234,N_24768,N_24295);
nand U25235 (N_25235,N_24070,N_24969);
or U25236 (N_25236,N_24920,N_24367);
and U25237 (N_25237,N_24254,N_24402);
or U25238 (N_25238,N_24708,N_24065);
nor U25239 (N_25239,N_24754,N_24351);
or U25240 (N_25240,N_24137,N_24575);
and U25241 (N_25241,N_24535,N_24688);
or U25242 (N_25242,N_24263,N_24784);
and U25243 (N_25243,N_24197,N_24352);
or U25244 (N_25244,N_24411,N_24476);
and U25245 (N_25245,N_24806,N_24028);
nor U25246 (N_25246,N_24355,N_24983);
and U25247 (N_25247,N_24030,N_24369);
and U25248 (N_25248,N_24506,N_24317);
nor U25249 (N_25249,N_24706,N_24406);
xnor U25250 (N_25250,N_24513,N_24131);
or U25251 (N_25251,N_24791,N_24389);
nand U25252 (N_25252,N_24171,N_24324);
and U25253 (N_25253,N_24245,N_24986);
nand U25254 (N_25254,N_24971,N_24970);
xnor U25255 (N_25255,N_24442,N_24330);
and U25256 (N_25256,N_24088,N_24420);
nor U25257 (N_25257,N_24899,N_24430);
and U25258 (N_25258,N_24681,N_24656);
nor U25259 (N_25259,N_24083,N_24102);
and U25260 (N_25260,N_24497,N_24626);
xnor U25261 (N_25261,N_24086,N_24564);
or U25262 (N_25262,N_24963,N_24427);
nand U25263 (N_25263,N_24454,N_24469);
or U25264 (N_25264,N_24690,N_24045);
and U25265 (N_25265,N_24422,N_24785);
xor U25266 (N_25266,N_24276,N_24852);
or U25267 (N_25267,N_24745,N_24491);
and U25268 (N_25268,N_24625,N_24908);
nand U25269 (N_25269,N_24922,N_24425);
or U25270 (N_25270,N_24377,N_24964);
or U25271 (N_25271,N_24771,N_24584);
nand U25272 (N_25272,N_24703,N_24955);
nor U25273 (N_25273,N_24056,N_24639);
or U25274 (N_25274,N_24072,N_24269);
xnor U25275 (N_25275,N_24262,N_24541);
nor U25276 (N_25276,N_24274,N_24953);
nor U25277 (N_25277,N_24495,N_24190);
nand U25278 (N_25278,N_24416,N_24665);
or U25279 (N_25279,N_24630,N_24494);
nand U25280 (N_25280,N_24026,N_24177);
nand U25281 (N_25281,N_24139,N_24658);
nand U25282 (N_25282,N_24198,N_24492);
xnor U25283 (N_25283,N_24977,N_24358);
or U25284 (N_25284,N_24772,N_24880);
nor U25285 (N_25285,N_24161,N_24634);
nor U25286 (N_25286,N_24363,N_24608);
and U25287 (N_25287,N_24246,N_24498);
nor U25288 (N_25288,N_24111,N_24879);
nor U25289 (N_25289,N_24984,N_24713);
and U25290 (N_25290,N_24638,N_24441);
xnor U25291 (N_25291,N_24023,N_24799);
or U25292 (N_25292,N_24082,N_24424);
nand U25293 (N_25293,N_24156,N_24035);
and U25294 (N_25294,N_24850,N_24040);
nor U25295 (N_25295,N_24405,N_24365);
or U25296 (N_25296,N_24487,N_24604);
xnor U25297 (N_25297,N_24397,N_24631);
nor U25298 (N_25298,N_24472,N_24106);
nor U25299 (N_25299,N_24629,N_24949);
or U25300 (N_25300,N_24044,N_24847);
nor U25301 (N_25301,N_24244,N_24300);
nand U25302 (N_25302,N_24826,N_24036);
nor U25303 (N_25303,N_24031,N_24504);
or U25304 (N_25304,N_24896,N_24645);
or U25305 (N_25305,N_24474,N_24116);
and U25306 (N_25306,N_24421,N_24210);
xnor U25307 (N_25307,N_24684,N_24952);
xor U25308 (N_25308,N_24940,N_24140);
nand U25309 (N_25309,N_24243,N_24350);
nor U25310 (N_25310,N_24982,N_24294);
or U25311 (N_25311,N_24789,N_24909);
xor U25312 (N_25312,N_24130,N_24844);
and U25313 (N_25313,N_24259,N_24598);
nor U25314 (N_25314,N_24444,N_24378);
xnor U25315 (N_25315,N_24904,N_24393);
or U25316 (N_25316,N_24861,N_24718);
nand U25317 (N_25317,N_24390,N_24746);
and U25318 (N_25318,N_24439,N_24434);
nand U25319 (N_25319,N_24968,N_24502);
and U25320 (N_25320,N_24216,N_24783);
nand U25321 (N_25321,N_24503,N_24018);
nor U25322 (N_25322,N_24816,N_24818);
nor U25323 (N_25323,N_24304,N_24273);
and U25324 (N_25324,N_24500,N_24180);
and U25325 (N_25325,N_24089,N_24680);
nor U25326 (N_25326,N_24855,N_24755);
and U25327 (N_25327,N_24172,N_24095);
nand U25328 (N_25328,N_24230,N_24473);
nand U25329 (N_25329,N_24903,N_24152);
xor U25330 (N_25330,N_24572,N_24409);
nor U25331 (N_25331,N_24010,N_24176);
and U25332 (N_25332,N_24897,N_24278);
and U25333 (N_25333,N_24901,N_24596);
or U25334 (N_25334,N_24336,N_24558);
and U25335 (N_25335,N_24619,N_24270);
nor U25336 (N_25336,N_24614,N_24595);
nand U25337 (N_25337,N_24514,N_24648);
or U25338 (N_25338,N_24710,N_24878);
or U25339 (N_25339,N_24452,N_24607);
nor U25340 (N_25340,N_24741,N_24004);
nand U25341 (N_25341,N_24194,N_24091);
or U25342 (N_25342,N_24512,N_24515);
xnor U25343 (N_25343,N_24882,N_24465);
nand U25344 (N_25344,N_24032,N_24551);
or U25345 (N_25345,N_24702,N_24581);
xor U25346 (N_25346,N_24548,N_24884);
nand U25347 (N_25347,N_24098,N_24362);
and U25348 (N_25348,N_24536,N_24678);
xnor U25349 (N_25349,N_24943,N_24980);
xnor U25350 (N_25350,N_24332,N_24461);
or U25351 (N_25351,N_24810,N_24340);
or U25352 (N_25352,N_24096,N_24739);
nor U25353 (N_25353,N_24618,N_24215);
xor U25354 (N_25354,N_24168,N_24877);
xor U25355 (N_25355,N_24714,N_24124);
and U25356 (N_25356,N_24449,N_24097);
and U25357 (N_25357,N_24100,N_24364);
nand U25358 (N_25358,N_24337,N_24328);
or U25359 (N_25359,N_24178,N_24696);
xor U25360 (N_25360,N_24672,N_24345);
or U25361 (N_25361,N_24864,N_24589);
or U25362 (N_25362,N_24620,N_24038);
nor U25363 (N_25363,N_24532,N_24484);
nor U25364 (N_25364,N_24542,N_24059);
or U25365 (N_25365,N_24241,N_24911);
nand U25366 (N_25366,N_24134,N_24600);
nand U25367 (N_25367,N_24933,N_24735);
nand U25368 (N_25368,N_24837,N_24122);
nor U25369 (N_25369,N_24959,N_24114);
and U25370 (N_25370,N_24293,N_24076);
or U25371 (N_25371,N_24252,N_24926);
nand U25372 (N_25372,N_24830,N_24412);
nand U25373 (N_25373,N_24524,N_24429);
nor U25374 (N_25374,N_24642,N_24635);
and U25375 (N_25375,N_24898,N_24936);
or U25376 (N_25376,N_24357,N_24829);
or U25377 (N_25377,N_24597,N_24573);
nor U25378 (N_25378,N_24385,N_24644);
xnor U25379 (N_25379,N_24486,N_24545);
and U25380 (N_25380,N_24029,N_24636);
or U25381 (N_25381,N_24115,N_24760);
nand U25382 (N_25382,N_24219,N_24318);
xnor U25383 (N_25383,N_24521,N_24951);
xnor U25384 (N_25384,N_24057,N_24080);
and U25385 (N_25385,N_24077,N_24092);
xnor U25386 (N_25386,N_24013,N_24895);
xor U25387 (N_25387,N_24927,N_24049);
xor U25388 (N_25388,N_24813,N_24213);
nor U25389 (N_25389,N_24375,N_24905);
xor U25390 (N_25390,N_24257,N_24087);
nand U25391 (N_25391,N_24460,N_24605);
nand U25392 (N_25392,N_24239,N_24531);
and U25393 (N_25393,N_24717,N_24759);
nor U25394 (N_25394,N_24074,N_24825);
or U25395 (N_25395,N_24599,N_24916);
xnor U25396 (N_25396,N_24777,N_24467);
xnor U25397 (N_25397,N_24733,N_24819);
nor U25398 (N_25398,N_24640,N_24331);
and U25399 (N_25399,N_24972,N_24946);
nor U25400 (N_25400,N_24343,N_24165);
nand U25401 (N_25401,N_24781,N_24655);
xnor U25402 (N_25402,N_24208,N_24488);
or U25403 (N_25403,N_24149,N_24824);
and U25404 (N_25404,N_24204,N_24661);
xor U25405 (N_25405,N_24085,N_24437);
nand U25406 (N_25406,N_24041,N_24578);
and U25407 (N_25407,N_24906,N_24530);
or U25408 (N_25408,N_24150,N_24788);
nand U25409 (N_25409,N_24822,N_24552);
and U25410 (N_25410,N_24123,N_24999);
nor U25411 (N_25411,N_24485,N_24737);
or U25412 (N_25412,N_24201,N_24185);
nand U25413 (N_25413,N_24870,N_24689);
or U25414 (N_25414,N_24797,N_24408);
or U25415 (N_25415,N_24078,N_24120);
nand U25416 (N_25416,N_24765,N_24957);
nand U25417 (N_25417,N_24828,N_24961);
or U25418 (N_25418,N_24939,N_24510);
xor U25419 (N_25419,N_24976,N_24628);
or U25420 (N_25420,N_24459,N_24546);
or U25421 (N_25421,N_24705,N_24480);
nor U25422 (N_25422,N_24667,N_24005);
and U25423 (N_25423,N_24477,N_24135);
and U25424 (N_25424,N_24071,N_24712);
nand U25425 (N_25425,N_24814,N_24651);
nor U25426 (N_25426,N_24496,N_24862);
nor U25427 (N_25427,N_24133,N_24591);
xor U25428 (N_25428,N_24587,N_24457);
nor U25429 (N_25429,N_24238,N_24214);
and U25430 (N_25430,N_24561,N_24209);
and U25431 (N_25431,N_24069,N_24987);
xor U25432 (N_25432,N_24786,N_24725);
xnor U25433 (N_25433,N_24179,N_24396);
or U25434 (N_25434,N_24858,N_24793);
and U25435 (N_25435,N_24679,N_24483);
nor U25436 (N_25436,N_24433,N_24027);
nand U25437 (N_25437,N_24019,N_24556);
and U25438 (N_25438,N_24222,N_24326);
xor U25439 (N_25439,N_24258,N_24921);
xor U25440 (N_25440,N_24632,N_24736);
and U25441 (N_25441,N_24748,N_24261);
and U25442 (N_25442,N_24839,N_24509);
nor U25443 (N_25443,N_24196,N_24283);
xor U25444 (N_25444,N_24728,N_24319);
or U25445 (N_25445,N_24153,N_24692);
or U25446 (N_25446,N_24501,N_24008);
and U25447 (N_25447,N_24650,N_24386);
xnor U25448 (N_25448,N_24356,N_24566);
and U25449 (N_25449,N_24663,N_24271);
xnor U25450 (N_25450,N_24286,N_24099);
nor U25451 (N_25451,N_24881,N_24199);
nand U25452 (N_25452,N_24290,N_24817);
or U25453 (N_25453,N_24053,N_24308);
xnor U25454 (N_25454,N_24700,N_24579);
and U25455 (N_25455,N_24333,N_24798);
xnor U25456 (N_25456,N_24988,N_24950);
nand U25457 (N_25457,N_24212,N_24206);
nor U25458 (N_25458,N_24577,N_24889);
or U25459 (N_25459,N_24301,N_24021);
and U25460 (N_25460,N_24919,N_24463);
nand U25461 (N_25461,N_24794,N_24404);
or U25462 (N_25462,N_24374,N_24188);
xnor U25463 (N_25463,N_24701,N_24167);
nor U25464 (N_25464,N_24415,N_24104);
xor U25465 (N_25465,N_24446,N_24051);
and U25466 (N_25466,N_24649,N_24849);
or U25467 (N_25467,N_24842,N_24388);
nand U25468 (N_25468,N_24699,N_24930);
nand U25469 (N_25469,N_24633,N_24382);
nand U25470 (N_25470,N_24321,N_24451);
nand U25471 (N_25471,N_24621,N_24641);
nand U25472 (N_25472,N_24346,N_24750);
and U25473 (N_25473,N_24202,N_24387);
or U25474 (N_25474,N_24155,N_24456);
nor U25475 (N_25475,N_24811,N_24932);
and U25476 (N_25476,N_24158,N_24475);
nor U25477 (N_25477,N_24743,N_24221);
nand U25478 (N_25478,N_24865,N_24006);
nand U25479 (N_25479,N_24121,N_24875);
and U25480 (N_25480,N_24313,N_24075);
nand U25481 (N_25481,N_24037,N_24594);
nor U25482 (N_25482,N_24787,N_24414);
nor U25483 (N_25483,N_24853,N_24848);
or U25484 (N_25484,N_24883,N_24695);
or U25485 (N_25485,N_24223,N_24282);
xor U25486 (N_25486,N_24108,N_24174);
or U25487 (N_25487,N_24910,N_24780);
nand U25488 (N_25488,N_24450,N_24470);
xor U25489 (N_25489,N_24659,N_24175);
nand U25490 (N_25490,N_24956,N_24327);
or U25491 (N_25491,N_24763,N_24846);
xnor U25492 (N_25492,N_24250,N_24997);
xor U25493 (N_25493,N_24154,N_24527);
nand U25494 (N_25494,N_24766,N_24309);
and U25495 (N_25495,N_24481,N_24312);
and U25496 (N_25496,N_24231,N_24565);
nor U25497 (N_25497,N_24200,N_24726);
and U25498 (N_25498,N_24874,N_24528);
nor U25499 (N_25499,N_24727,N_24042);
nand U25500 (N_25500,N_24410,N_24140);
nor U25501 (N_25501,N_24049,N_24066);
or U25502 (N_25502,N_24407,N_24339);
nor U25503 (N_25503,N_24333,N_24251);
nand U25504 (N_25504,N_24292,N_24769);
nor U25505 (N_25505,N_24516,N_24907);
nor U25506 (N_25506,N_24313,N_24722);
and U25507 (N_25507,N_24056,N_24790);
and U25508 (N_25508,N_24358,N_24728);
nand U25509 (N_25509,N_24613,N_24722);
xor U25510 (N_25510,N_24272,N_24301);
xor U25511 (N_25511,N_24661,N_24659);
nor U25512 (N_25512,N_24994,N_24269);
nand U25513 (N_25513,N_24192,N_24329);
xnor U25514 (N_25514,N_24199,N_24792);
and U25515 (N_25515,N_24016,N_24201);
xor U25516 (N_25516,N_24149,N_24560);
or U25517 (N_25517,N_24103,N_24946);
xor U25518 (N_25518,N_24916,N_24443);
xnor U25519 (N_25519,N_24435,N_24032);
nand U25520 (N_25520,N_24841,N_24119);
nor U25521 (N_25521,N_24694,N_24996);
nor U25522 (N_25522,N_24840,N_24153);
nor U25523 (N_25523,N_24966,N_24768);
and U25524 (N_25524,N_24477,N_24472);
nand U25525 (N_25525,N_24555,N_24652);
and U25526 (N_25526,N_24595,N_24679);
and U25527 (N_25527,N_24794,N_24166);
xor U25528 (N_25528,N_24578,N_24459);
or U25529 (N_25529,N_24370,N_24098);
or U25530 (N_25530,N_24291,N_24939);
and U25531 (N_25531,N_24964,N_24163);
xnor U25532 (N_25532,N_24402,N_24403);
nand U25533 (N_25533,N_24745,N_24311);
xor U25534 (N_25534,N_24031,N_24115);
nor U25535 (N_25535,N_24663,N_24976);
xor U25536 (N_25536,N_24119,N_24347);
xor U25537 (N_25537,N_24489,N_24049);
and U25538 (N_25538,N_24318,N_24981);
or U25539 (N_25539,N_24589,N_24471);
and U25540 (N_25540,N_24098,N_24035);
nand U25541 (N_25541,N_24973,N_24736);
nand U25542 (N_25542,N_24961,N_24749);
nand U25543 (N_25543,N_24424,N_24414);
nor U25544 (N_25544,N_24447,N_24823);
nor U25545 (N_25545,N_24271,N_24978);
and U25546 (N_25546,N_24089,N_24583);
nand U25547 (N_25547,N_24170,N_24849);
nand U25548 (N_25548,N_24145,N_24186);
nand U25549 (N_25549,N_24972,N_24400);
or U25550 (N_25550,N_24422,N_24539);
nor U25551 (N_25551,N_24175,N_24479);
nor U25552 (N_25552,N_24406,N_24887);
nand U25553 (N_25553,N_24715,N_24190);
and U25554 (N_25554,N_24668,N_24085);
nand U25555 (N_25555,N_24063,N_24201);
or U25556 (N_25556,N_24277,N_24534);
and U25557 (N_25557,N_24510,N_24352);
xnor U25558 (N_25558,N_24444,N_24590);
nor U25559 (N_25559,N_24519,N_24243);
xnor U25560 (N_25560,N_24487,N_24348);
nand U25561 (N_25561,N_24685,N_24590);
nor U25562 (N_25562,N_24101,N_24282);
nor U25563 (N_25563,N_24111,N_24741);
nor U25564 (N_25564,N_24332,N_24920);
xnor U25565 (N_25565,N_24484,N_24079);
xnor U25566 (N_25566,N_24605,N_24080);
and U25567 (N_25567,N_24315,N_24941);
and U25568 (N_25568,N_24890,N_24070);
xor U25569 (N_25569,N_24303,N_24934);
and U25570 (N_25570,N_24384,N_24886);
and U25571 (N_25571,N_24134,N_24021);
nand U25572 (N_25572,N_24177,N_24247);
and U25573 (N_25573,N_24304,N_24940);
xnor U25574 (N_25574,N_24975,N_24945);
xor U25575 (N_25575,N_24651,N_24247);
and U25576 (N_25576,N_24189,N_24122);
nand U25577 (N_25577,N_24470,N_24685);
nor U25578 (N_25578,N_24425,N_24864);
nor U25579 (N_25579,N_24703,N_24933);
or U25580 (N_25580,N_24287,N_24713);
and U25581 (N_25581,N_24264,N_24198);
nand U25582 (N_25582,N_24936,N_24079);
nand U25583 (N_25583,N_24280,N_24146);
nand U25584 (N_25584,N_24112,N_24189);
and U25585 (N_25585,N_24250,N_24108);
or U25586 (N_25586,N_24209,N_24768);
xnor U25587 (N_25587,N_24374,N_24937);
nor U25588 (N_25588,N_24815,N_24365);
or U25589 (N_25589,N_24633,N_24356);
nand U25590 (N_25590,N_24021,N_24345);
and U25591 (N_25591,N_24029,N_24358);
nand U25592 (N_25592,N_24015,N_24325);
nand U25593 (N_25593,N_24439,N_24671);
xor U25594 (N_25594,N_24211,N_24757);
nor U25595 (N_25595,N_24512,N_24643);
xnor U25596 (N_25596,N_24146,N_24915);
nand U25597 (N_25597,N_24947,N_24102);
nor U25598 (N_25598,N_24548,N_24812);
xnor U25599 (N_25599,N_24234,N_24267);
or U25600 (N_25600,N_24502,N_24002);
nor U25601 (N_25601,N_24357,N_24546);
nand U25602 (N_25602,N_24375,N_24348);
or U25603 (N_25603,N_24810,N_24270);
xor U25604 (N_25604,N_24128,N_24220);
and U25605 (N_25605,N_24680,N_24279);
nand U25606 (N_25606,N_24425,N_24152);
nor U25607 (N_25607,N_24447,N_24681);
or U25608 (N_25608,N_24823,N_24358);
nand U25609 (N_25609,N_24839,N_24108);
or U25610 (N_25610,N_24482,N_24933);
and U25611 (N_25611,N_24260,N_24285);
or U25612 (N_25612,N_24650,N_24669);
and U25613 (N_25613,N_24573,N_24581);
or U25614 (N_25614,N_24987,N_24211);
and U25615 (N_25615,N_24620,N_24300);
nor U25616 (N_25616,N_24022,N_24653);
or U25617 (N_25617,N_24198,N_24986);
or U25618 (N_25618,N_24308,N_24795);
nor U25619 (N_25619,N_24649,N_24575);
or U25620 (N_25620,N_24805,N_24201);
and U25621 (N_25621,N_24753,N_24100);
and U25622 (N_25622,N_24807,N_24033);
and U25623 (N_25623,N_24283,N_24274);
nand U25624 (N_25624,N_24469,N_24551);
and U25625 (N_25625,N_24733,N_24210);
nand U25626 (N_25626,N_24189,N_24005);
xor U25627 (N_25627,N_24286,N_24282);
or U25628 (N_25628,N_24222,N_24180);
xor U25629 (N_25629,N_24896,N_24249);
and U25630 (N_25630,N_24000,N_24958);
xor U25631 (N_25631,N_24536,N_24375);
or U25632 (N_25632,N_24866,N_24003);
nor U25633 (N_25633,N_24185,N_24371);
or U25634 (N_25634,N_24066,N_24237);
or U25635 (N_25635,N_24951,N_24197);
and U25636 (N_25636,N_24214,N_24930);
nor U25637 (N_25637,N_24598,N_24768);
nand U25638 (N_25638,N_24949,N_24380);
or U25639 (N_25639,N_24085,N_24279);
and U25640 (N_25640,N_24225,N_24750);
or U25641 (N_25641,N_24704,N_24292);
nor U25642 (N_25642,N_24607,N_24155);
and U25643 (N_25643,N_24479,N_24162);
and U25644 (N_25644,N_24672,N_24385);
and U25645 (N_25645,N_24232,N_24306);
nand U25646 (N_25646,N_24612,N_24575);
nand U25647 (N_25647,N_24236,N_24260);
nand U25648 (N_25648,N_24105,N_24478);
xnor U25649 (N_25649,N_24204,N_24777);
xnor U25650 (N_25650,N_24646,N_24038);
and U25651 (N_25651,N_24018,N_24619);
nor U25652 (N_25652,N_24406,N_24563);
nand U25653 (N_25653,N_24092,N_24655);
xor U25654 (N_25654,N_24928,N_24850);
or U25655 (N_25655,N_24934,N_24828);
nor U25656 (N_25656,N_24001,N_24024);
and U25657 (N_25657,N_24294,N_24999);
nor U25658 (N_25658,N_24331,N_24134);
nor U25659 (N_25659,N_24974,N_24869);
nand U25660 (N_25660,N_24440,N_24904);
xor U25661 (N_25661,N_24302,N_24519);
and U25662 (N_25662,N_24515,N_24573);
and U25663 (N_25663,N_24391,N_24477);
nand U25664 (N_25664,N_24280,N_24197);
xnor U25665 (N_25665,N_24693,N_24219);
xnor U25666 (N_25666,N_24047,N_24845);
xnor U25667 (N_25667,N_24341,N_24866);
xor U25668 (N_25668,N_24194,N_24760);
xor U25669 (N_25669,N_24751,N_24573);
nor U25670 (N_25670,N_24216,N_24695);
or U25671 (N_25671,N_24471,N_24911);
or U25672 (N_25672,N_24967,N_24232);
nor U25673 (N_25673,N_24203,N_24143);
nor U25674 (N_25674,N_24843,N_24719);
nor U25675 (N_25675,N_24695,N_24425);
or U25676 (N_25676,N_24393,N_24374);
or U25677 (N_25677,N_24681,N_24082);
nor U25678 (N_25678,N_24688,N_24160);
nand U25679 (N_25679,N_24018,N_24198);
nand U25680 (N_25680,N_24725,N_24421);
or U25681 (N_25681,N_24795,N_24959);
nand U25682 (N_25682,N_24166,N_24942);
or U25683 (N_25683,N_24848,N_24020);
nor U25684 (N_25684,N_24733,N_24116);
xor U25685 (N_25685,N_24726,N_24873);
xnor U25686 (N_25686,N_24070,N_24676);
nor U25687 (N_25687,N_24265,N_24493);
or U25688 (N_25688,N_24748,N_24122);
or U25689 (N_25689,N_24996,N_24804);
nand U25690 (N_25690,N_24884,N_24097);
and U25691 (N_25691,N_24960,N_24546);
nand U25692 (N_25692,N_24852,N_24825);
nand U25693 (N_25693,N_24763,N_24513);
nor U25694 (N_25694,N_24934,N_24332);
and U25695 (N_25695,N_24016,N_24055);
xor U25696 (N_25696,N_24303,N_24357);
xor U25697 (N_25697,N_24739,N_24985);
nor U25698 (N_25698,N_24890,N_24256);
nor U25699 (N_25699,N_24309,N_24707);
nor U25700 (N_25700,N_24201,N_24654);
nand U25701 (N_25701,N_24699,N_24161);
or U25702 (N_25702,N_24680,N_24442);
and U25703 (N_25703,N_24084,N_24555);
xor U25704 (N_25704,N_24126,N_24076);
and U25705 (N_25705,N_24820,N_24464);
and U25706 (N_25706,N_24553,N_24446);
nor U25707 (N_25707,N_24661,N_24857);
nand U25708 (N_25708,N_24866,N_24536);
or U25709 (N_25709,N_24720,N_24939);
and U25710 (N_25710,N_24466,N_24750);
and U25711 (N_25711,N_24942,N_24817);
nor U25712 (N_25712,N_24015,N_24546);
or U25713 (N_25713,N_24082,N_24697);
or U25714 (N_25714,N_24529,N_24712);
or U25715 (N_25715,N_24141,N_24589);
xor U25716 (N_25716,N_24869,N_24518);
and U25717 (N_25717,N_24263,N_24383);
xor U25718 (N_25718,N_24499,N_24776);
xor U25719 (N_25719,N_24835,N_24797);
nand U25720 (N_25720,N_24714,N_24252);
nor U25721 (N_25721,N_24865,N_24454);
and U25722 (N_25722,N_24142,N_24937);
nand U25723 (N_25723,N_24055,N_24286);
nand U25724 (N_25724,N_24282,N_24326);
and U25725 (N_25725,N_24936,N_24998);
nand U25726 (N_25726,N_24734,N_24038);
and U25727 (N_25727,N_24580,N_24958);
xnor U25728 (N_25728,N_24807,N_24803);
xnor U25729 (N_25729,N_24768,N_24837);
nand U25730 (N_25730,N_24244,N_24342);
nand U25731 (N_25731,N_24595,N_24237);
and U25732 (N_25732,N_24469,N_24201);
nor U25733 (N_25733,N_24904,N_24310);
xor U25734 (N_25734,N_24210,N_24458);
and U25735 (N_25735,N_24435,N_24439);
nor U25736 (N_25736,N_24817,N_24906);
nor U25737 (N_25737,N_24684,N_24505);
or U25738 (N_25738,N_24894,N_24672);
or U25739 (N_25739,N_24394,N_24574);
or U25740 (N_25740,N_24999,N_24650);
nor U25741 (N_25741,N_24657,N_24135);
and U25742 (N_25742,N_24169,N_24979);
nor U25743 (N_25743,N_24774,N_24841);
and U25744 (N_25744,N_24797,N_24296);
xnor U25745 (N_25745,N_24192,N_24169);
xnor U25746 (N_25746,N_24169,N_24962);
nand U25747 (N_25747,N_24160,N_24283);
nor U25748 (N_25748,N_24955,N_24486);
nor U25749 (N_25749,N_24974,N_24023);
and U25750 (N_25750,N_24890,N_24860);
xnor U25751 (N_25751,N_24827,N_24992);
and U25752 (N_25752,N_24464,N_24950);
nor U25753 (N_25753,N_24870,N_24621);
and U25754 (N_25754,N_24819,N_24936);
nand U25755 (N_25755,N_24927,N_24270);
nand U25756 (N_25756,N_24844,N_24049);
xnor U25757 (N_25757,N_24072,N_24010);
nor U25758 (N_25758,N_24692,N_24209);
or U25759 (N_25759,N_24972,N_24314);
and U25760 (N_25760,N_24131,N_24737);
or U25761 (N_25761,N_24915,N_24181);
or U25762 (N_25762,N_24012,N_24461);
and U25763 (N_25763,N_24769,N_24207);
or U25764 (N_25764,N_24027,N_24421);
xor U25765 (N_25765,N_24910,N_24725);
nand U25766 (N_25766,N_24977,N_24282);
and U25767 (N_25767,N_24456,N_24988);
nand U25768 (N_25768,N_24406,N_24441);
nor U25769 (N_25769,N_24174,N_24804);
and U25770 (N_25770,N_24695,N_24679);
and U25771 (N_25771,N_24389,N_24862);
nand U25772 (N_25772,N_24788,N_24583);
nor U25773 (N_25773,N_24865,N_24392);
nand U25774 (N_25774,N_24782,N_24143);
xor U25775 (N_25775,N_24963,N_24120);
nand U25776 (N_25776,N_24836,N_24631);
nand U25777 (N_25777,N_24352,N_24301);
nand U25778 (N_25778,N_24294,N_24800);
or U25779 (N_25779,N_24943,N_24601);
or U25780 (N_25780,N_24638,N_24780);
or U25781 (N_25781,N_24116,N_24143);
nor U25782 (N_25782,N_24107,N_24589);
nor U25783 (N_25783,N_24200,N_24792);
or U25784 (N_25784,N_24154,N_24776);
and U25785 (N_25785,N_24429,N_24170);
xnor U25786 (N_25786,N_24832,N_24230);
or U25787 (N_25787,N_24473,N_24058);
nand U25788 (N_25788,N_24873,N_24130);
nand U25789 (N_25789,N_24830,N_24403);
and U25790 (N_25790,N_24089,N_24799);
xnor U25791 (N_25791,N_24102,N_24848);
nor U25792 (N_25792,N_24253,N_24453);
xor U25793 (N_25793,N_24356,N_24270);
and U25794 (N_25794,N_24795,N_24511);
xor U25795 (N_25795,N_24119,N_24647);
and U25796 (N_25796,N_24047,N_24739);
and U25797 (N_25797,N_24778,N_24975);
nor U25798 (N_25798,N_24616,N_24245);
xor U25799 (N_25799,N_24172,N_24130);
nor U25800 (N_25800,N_24681,N_24915);
or U25801 (N_25801,N_24600,N_24806);
nand U25802 (N_25802,N_24598,N_24161);
or U25803 (N_25803,N_24474,N_24732);
and U25804 (N_25804,N_24633,N_24319);
or U25805 (N_25805,N_24742,N_24389);
nand U25806 (N_25806,N_24854,N_24369);
xnor U25807 (N_25807,N_24143,N_24576);
nand U25808 (N_25808,N_24889,N_24890);
and U25809 (N_25809,N_24218,N_24011);
and U25810 (N_25810,N_24290,N_24567);
or U25811 (N_25811,N_24786,N_24679);
nand U25812 (N_25812,N_24003,N_24152);
nor U25813 (N_25813,N_24715,N_24090);
nand U25814 (N_25814,N_24684,N_24487);
and U25815 (N_25815,N_24984,N_24204);
or U25816 (N_25816,N_24738,N_24513);
nand U25817 (N_25817,N_24613,N_24607);
or U25818 (N_25818,N_24142,N_24422);
and U25819 (N_25819,N_24086,N_24543);
xnor U25820 (N_25820,N_24214,N_24479);
nand U25821 (N_25821,N_24786,N_24389);
nor U25822 (N_25822,N_24083,N_24011);
and U25823 (N_25823,N_24766,N_24365);
and U25824 (N_25824,N_24573,N_24755);
and U25825 (N_25825,N_24562,N_24213);
xor U25826 (N_25826,N_24213,N_24504);
xor U25827 (N_25827,N_24989,N_24044);
nand U25828 (N_25828,N_24276,N_24820);
nor U25829 (N_25829,N_24773,N_24020);
and U25830 (N_25830,N_24705,N_24022);
and U25831 (N_25831,N_24356,N_24955);
nand U25832 (N_25832,N_24090,N_24518);
nand U25833 (N_25833,N_24599,N_24870);
or U25834 (N_25834,N_24427,N_24409);
nor U25835 (N_25835,N_24205,N_24328);
and U25836 (N_25836,N_24800,N_24426);
nor U25837 (N_25837,N_24174,N_24164);
or U25838 (N_25838,N_24458,N_24659);
or U25839 (N_25839,N_24918,N_24492);
nor U25840 (N_25840,N_24693,N_24441);
or U25841 (N_25841,N_24151,N_24656);
nor U25842 (N_25842,N_24010,N_24145);
nand U25843 (N_25843,N_24073,N_24357);
xnor U25844 (N_25844,N_24596,N_24989);
and U25845 (N_25845,N_24109,N_24714);
and U25846 (N_25846,N_24906,N_24112);
nand U25847 (N_25847,N_24943,N_24933);
nand U25848 (N_25848,N_24449,N_24011);
or U25849 (N_25849,N_24010,N_24754);
or U25850 (N_25850,N_24887,N_24429);
or U25851 (N_25851,N_24175,N_24716);
xnor U25852 (N_25852,N_24155,N_24515);
nor U25853 (N_25853,N_24474,N_24963);
xor U25854 (N_25854,N_24661,N_24614);
and U25855 (N_25855,N_24724,N_24922);
or U25856 (N_25856,N_24718,N_24899);
and U25857 (N_25857,N_24043,N_24275);
nand U25858 (N_25858,N_24262,N_24219);
nor U25859 (N_25859,N_24468,N_24339);
nand U25860 (N_25860,N_24826,N_24839);
and U25861 (N_25861,N_24957,N_24905);
nor U25862 (N_25862,N_24634,N_24758);
nor U25863 (N_25863,N_24552,N_24043);
nand U25864 (N_25864,N_24204,N_24227);
nand U25865 (N_25865,N_24105,N_24692);
xor U25866 (N_25866,N_24986,N_24304);
xnor U25867 (N_25867,N_24875,N_24763);
nand U25868 (N_25868,N_24525,N_24581);
or U25869 (N_25869,N_24539,N_24636);
xor U25870 (N_25870,N_24499,N_24432);
nand U25871 (N_25871,N_24664,N_24705);
xor U25872 (N_25872,N_24283,N_24824);
nor U25873 (N_25873,N_24575,N_24559);
or U25874 (N_25874,N_24108,N_24887);
and U25875 (N_25875,N_24925,N_24917);
xor U25876 (N_25876,N_24962,N_24441);
and U25877 (N_25877,N_24867,N_24838);
nand U25878 (N_25878,N_24738,N_24215);
xnor U25879 (N_25879,N_24059,N_24972);
or U25880 (N_25880,N_24038,N_24471);
nor U25881 (N_25881,N_24176,N_24328);
xor U25882 (N_25882,N_24288,N_24393);
nand U25883 (N_25883,N_24492,N_24485);
xnor U25884 (N_25884,N_24315,N_24855);
nor U25885 (N_25885,N_24767,N_24447);
nand U25886 (N_25886,N_24250,N_24422);
and U25887 (N_25887,N_24020,N_24013);
nand U25888 (N_25888,N_24228,N_24250);
nand U25889 (N_25889,N_24082,N_24803);
nand U25890 (N_25890,N_24756,N_24934);
and U25891 (N_25891,N_24995,N_24870);
nor U25892 (N_25892,N_24501,N_24196);
nand U25893 (N_25893,N_24604,N_24144);
and U25894 (N_25894,N_24351,N_24879);
nand U25895 (N_25895,N_24514,N_24121);
and U25896 (N_25896,N_24039,N_24307);
nand U25897 (N_25897,N_24037,N_24786);
and U25898 (N_25898,N_24126,N_24924);
or U25899 (N_25899,N_24882,N_24476);
xor U25900 (N_25900,N_24851,N_24142);
and U25901 (N_25901,N_24124,N_24654);
nand U25902 (N_25902,N_24431,N_24675);
or U25903 (N_25903,N_24799,N_24560);
nand U25904 (N_25904,N_24626,N_24280);
nor U25905 (N_25905,N_24014,N_24971);
and U25906 (N_25906,N_24339,N_24706);
and U25907 (N_25907,N_24486,N_24146);
and U25908 (N_25908,N_24318,N_24879);
xnor U25909 (N_25909,N_24861,N_24140);
nand U25910 (N_25910,N_24694,N_24137);
and U25911 (N_25911,N_24113,N_24089);
nand U25912 (N_25912,N_24122,N_24982);
nand U25913 (N_25913,N_24088,N_24553);
or U25914 (N_25914,N_24091,N_24154);
xor U25915 (N_25915,N_24746,N_24948);
or U25916 (N_25916,N_24165,N_24125);
xnor U25917 (N_25917,N_24902,N_24379);
or U25918 (N_25918,N_24819,N_24219);
xnor U25919 (N_25919,N_24304,N_24719);
or U25920 (N_25920,N_24752,N_24701);
nand U25921 (N_25921,N_24314,N_24403);
and U25922 (N_25922,N_24199,N_24159);
nand U25923 (N_25923,N_24744,N_24074);
nand U25924 (N_25924,N_24009,N_24819);
or U25925 (N_25925,N_24305,N_24880);
xnor U25926 (N_25926,N_24253,N_24374);
or U25927 (N_25927,N_24154,N_24452);
nand U25928 (N_25928,N_24853,N_24602);
nor U25929 (N_25929,N_24661,N_24618);
nand U25930 (N_25930,N_24296,N_24872);
nor U25931 (N_25931,N_24729,N_24826);
nand U25932 (N_25932,N_24114,N_24954);
nor U25933 (N_25933,N_24613,N_24465);
xnor U25934 (N_25934,N_24547,N_24712);
or U25935 (N_25935,N_24639,N_24456);
or U25936 (N_25936,N_24786,N_24348);
nand U25937 (N_25937,N_24128,N_24647);
nand U25938 (N_25938,N_24381,N_24662);
nor U25939 (N_25939,N_24223,N_24032);
and U25940 (N_25940,N_24960,N_24799);
xor U25941 (N_25941,N_24346,N_24988);
nand U25942 (N_25942,N_24314,N_24186);
or U25943 (N_25943,N_24806,N_24156);
and U25944 (N_25944,N_24651,N_24337);
nor U25945 (N_25945,N_24294,N_24332);
and U25946 (N_25946,N_24000,N_24684);
nor U25947 (N_25947,N_24636,N_24950);
xor U25948 (N_25948,N_24283,N_24362);
nand U25949 (N_25949,N_24540,N_24182);
or U25950 (N_25950,N_24905,N_24201);
or U25951 (N_25951,N_24342,N_24518);
and U25952 (N_25952,N_24764,N_24767);
nand U25953 (N_25953,N_24893,N_24508);
xnor U25954 (N_25954,N_24595,N_24722);
and U25955 (N_25955,N_24931,N_24550);
and U25956 (N_25956,N_24203,N_24377);
xor U25957 (N_25957,N_24958,N_24564);
xnor U25958 (N_25958,N_24829,N_24438);
xnor U25959 (N_25959,N_24096,N_24398);
nor U25960 (N_25960,N_24232,N_24830);
xor U25961 (N_25961,N_24073,N_24661);
or U25962 (N_25962,N_24203,N_24053);
xor U25963 (N_25963,N_24983,N_24029);
nor U25964 (N_25964,N_24647,N_24876);
nand U25965 (N_25965,N_24570,N_24932);
xor U25966 (N_25966,N_24026,N_24216);
nor U25967 (N_25967,N_24341,N_24713);
or U25968 (N_25968,N_24325,N_24742);
xnor U25969 (N_25969,N_24971,N_24688);
xnor U25970 (N_25970,N_24869,N_24961);
nor U25971 (N_25971,N_24640,N_24146);
or U25972 (N_25972,N_24470,N_24701);
and U25973 (N_25973,N_24191,N_24529);
nand U25974 (N_25974,N_24036,N_24635);
or U25975 (N_25975,N_24558,N_24165);
nand U25976 (N_25976,N_24297,N_24355);
and U25977 (N_25977,N_24822,N_24946);
xnor U25978 (N_25978,N_24219,N_24292);
nor U25979 (N_25979,N_24736,N_24966);
xor U25980 (N_25980,N_24297,N_24602);
nand U25981 (N_25981,N_24484,N_24109);
and U25982 (N_25982,N_24480,N_24649);
nand U25983 (N_25983,N_24158,N_24465);
or U25984 (N_25984,N_24958,N_24261);
xnor U25985 (N_25985,N_24238,N_24018);
or U25986 (N_25986,N_24212,N_24541);
nor U25987 (N_25987,N_24300,N_24948);
xor U25988 (N_25988,N_24119,N_24790);
and U25989 (N_25989,N_24064,N_24197);
nor U25990 (N_25990,N_24566,N_24795);
nor U25991 (N_25991,N_24991,N_24186);
and U25992 (N_25992,N_24344,N_24099);
nor U25993 (N_25993,N_24122,N_24248);
nand U25994 (N_25994,N_24560,N_24287);
nand U25995 (N_25995,N_24051,N_24491);
and U25996 (N_25996,N_24046,N_24352);
nand U25997 (N_25997,N_24046,N_24828);
or U25998 (N_25998,N_24581,N_24277);
nand U25999 (N_25999,N_24258,N_24293);
nand U26000 (N_26000,N_25367,N_25225);
and U26001 (N_26001,N_25251,N_25463);
or U26002 (N_26002,N_25525,N_25204);
or U26003 (N_26003,N_25377,N_25779);
nor U26004 (N_26004,N_25338,N_25383);
and U26005 (N_26005,N_25630,N_25471);
and U26006 (N_26006,N_25864,N_25918);
xor U26007 (N_26007,N_25831,N_25589);
nor U26008 (N_26008,N_25060,N_25640);
or U26009 (N_26009,N_25873,N_25303);
or U26010 (N_26010,N_25897,N_25657);
and U26011 (N_26011,N_25645,N_25175);
and U26012 (N_26012,N_25600,N_25389);
nand U26013 (N_26013,N_25989,N_25635);
nor U26014 (N_26014,N_25050,N_25135);
or U26015 (N_26015,N_25540,N_25947);
or U26016 (N_26016,N_25654,N_25242);
nand U26017 (N_26017,N_25777,N_25130);
or U26018 (N_26018,N_25797,N_25223);
xnor U26019 (N_26019,N_25519,N_25205);
xnor U26020 (N_26020,N_25104,N_25454);
or U26021 (N_26021,N_25033,N_25821);
xor U26022 (N_26022,N_25714,N_25169);
nand U26023 (N_26023,N_25070,N_25928);
xor U26024 (N_26024,N_25841,N_25909);
xnor U26025 (N_26025,N_25839,N_25751);
nand U26026 (N_26026,N_25164,N_25951);
nand U26027 (N_26027,N_25412,N_25224);
or U26028 (N_26028,N_25510,N_25384);
and U26029 (N_26029,N_25980,N_25792);
or U26030 (N_26030,N_25903,N_25261);
and U26031 (N_26031,N_25983,N_25585);
and U26032 (N_26032,N_25647,N_25019);
nor U26033 (N_26033,N_25183,N_25290);
nand U26034 (N_26034,N_25730,N_25310);
and U26035 (N_26035,N_25020,N_25313);
nand U26036 (N_26036,N_25505,N_25443);
nand U26037 (N_26037,N_25087,N_25532);
nand U26038 (N_26038,N_25473,N_25031);
or U26039 (N_26039,N_25602,N_25518);
xor U26040 (N_26040,N_25770,N_25355);
nand U26041 (N_26041,N_25101,N_25123);
xnor U26042 (N_26042,N_25764,N_25206);
xor U26043 (N_26043,N_25984,N_25273);
nor U26044 (N_26044,N_25590,N_25131);
nand U26045 (N_26045,N_25682,N_25535);
and U26046 (N_26046,N_25154,N_25812);
xor U26047 (N_26047,N_25361,N_25650);
and U26048 (N_26048,N_25920,N_25360);
and U26049 (N_26049,N_25567,N_25392);
xnor U26050 (N_26050,N_25830,N_25969);
xnor U26051 (N_26051,N_25304,N_25450);
nand U26052 (N_26052,N_25874,N_25807);
or U26053 (N_26053,N_25343,N_25368);
and U26054 (N_26054,N_25055,N_25100);
nand U26055 (N_26055,N_25374,N_25965);
and U26056 (N_26056,N_25817,N_25744);
xor U26057 (N_26057,N_25769,N_25964);
nor U26058 (N_26058,N_25165,N_25021);
xnor U26059 (N_26059,N_25347,N_25746);
or U26060 (N_26060,N_25911,N_25943);
nand U26061 (N_26061,N_25599,N_25474);
nand U26062 (N_26062,N_25760,N_25973);
xor U26063 (N_26063,N_25143,N_25122);
nand U26064 (N_26064,N_25722,N_25944);
xor U26065 (N_26065,N_25125,N_25774);
and U26066 (N_26066,N_25315,N_25761);
xnor U26067 (N_26067,N_25234,N_25278);
and U26068 (N_26068,N_25913,N_25128);
nand U26069 (N_26069,N_25924,N_25086);
or U26070 (N_26070,N_25322,N_25621);
nand U26071 (N_26071,N_25255,N_25741);
nand U26072 (N_26072,N_25869,N_25414);
and U26073 (N_26073,N_25340,N_25112);
or U26074 (N_26074,N_25974,N_25546);
or U26075 (N_26075,N_25045,N_25954);
or U26076 (N_26076,N_25925,N_25399);
nand U26077 (N_26077,N_25622,N_25228);
nand U26078 (N_26078,N_25179,N_25010);
and U26079 (N_26079,N_25369,N_25079);
nor U26080 (N_26080,N_25678,N_25308);
xor U26081 (N_26081,N_25213,N_25407);
nor U26082 (N_26082,N_25092,N_25140);
nand U26083 (N_26083,N_25476,N_25642);
or U26084 (N_26084,N_25419,N_25398);
xor U26085 (N_26085,N_25811,N_25819);
xnor U26086 (N_26086,N_25966,N_25058);
and U26087 (N_26087,N_25043,N_25095);
nand U26088 (N_26088,N_25544,N_25272);
and U26089 (N_26089,N_25366,N_25145);
and U26090 (N_26090,N_25653,N_25666);
nor U26091 (N_26091,N_25047,N_25523);
and U26092 (N_26092,N_25007,N_25513);
nor U26093 (N_26093,N_25017,N_25591);
nor U26094 (N_26094,N_25006,N_25296);
nor U26095 (N_26095,N_25960,N_25431);
nand U26096 (N_26096,N_25117,N_25511);
and U26097 (N_26097,N_25910,N_25293);
or U26098 (N_26098,N_25916,N_25302);
nand U26099 (N_26099,N_25765,N_25762);
nor U26100 (N_26100,N_25702,N_25468);
nor U26101 (N_26101,N_25306,N_25766);
or U26102 (N_26102,N_25705,N_25294);
nor U26103 (N_26103,N_25784,N_25876);
nor U26104 (N_26104,N_25351,N_25096);
nand U26105 (N_26105,N_25814,N_25161);
and U26106 (N_26106,N_25957,N_25276);
nor U26107 (N_26107,N_25708,N_25977);
or U26108 (N_26108,N_25402,N_25053);
nand U26109 (N_26109,N_25978,N_25815);
xor U26110 (N_26110,N_25598,N_25734);
xnor U26111 (N_26111,N_25756,N_25805);
nor U26112 (N_26112,N_25328,N_25502);
or U26113 (N_26113,N_25512,N_25250);
nand U26114 (N_26114,N_25386,N_25063);
xor U26115 (N_26115,N_25936,N_25156);
nor U26116 (N_26116,N_25789,N_25067);
xnor U26117 (N_26117,N_25847,N_25845);
and U26118 (N_26118,N_25241,N_25478);
xor U26119 (N_26119,N_25046,N_25271);
and U26120 (N_26120,N_25329,N_25556);
nand U26121 (N_26121,N_25015,N_25578);
xnor U26122 (N_26122,N_25754,N_25301);
xor U26123 (N_26123,N_25324,N_25417);
xor U26124 (N_26124,N_25504,N_25549);
and U26125 (N_26125,N_25515,N_25090);
nand U26126 (N_26126,N_25452,N_25687);
nand U26127 (N_26127,N_25037,N_25217);
nand U26128 (N_26128,N_25371,N_25268);
or U26129 (N_26129,N_25231,N_25061);
xor U26130 (N_26130,N_25976,N_25636);
nor U26131 (N_26131,N_25758,N_25029);
or U26132 (N_26132,N_25114,N_25262);
and U26133 (N_26133,N_25042,N_25562);
xnor U26134 (N_26134,N_25962,N_25877);
nor U26135 (N_26135,N_25575,N_25625);
nand U26136 (N_26136,N_25923,N_25227);
nand U26137 (N_26137,N_25721,N_25307);
xor U26138 (N_26138,N_25970,N_25616);
nand U26139 (N_26139,N_25782,N_25023);
or U26140 (N_26140,N_25768,N_25898);
and U26141 (N_26141,N_25305,N_25545);
nor U26142 (N_26142,N_25285,N_25215);
nor U26143 (N_26143,N_25894,N_25693);
and U26144 (N_26144,N_25345,N_25813);
and U26145 (N_26145,N_25915,N_25009);
nor U26146 (N_26146,N_25427,N_25646);
or U26147 (N_26147,N_25449,N_25159);
or U26148 (N_26148,N_25181,N_25890);
and U26149 (N_26149,N_25150,N_25025);
nand U26150 (N_26150,N_25882,N_25445);
xor U26151 (N_26151,N_25275,N_25036);
xnor U26152 (N_26152,N_25942,N_25363);
nand U26153 (N_26153,N_25553,N_25319);
or U26154 (N_26154,N_25587,N_25052);
xnor U26155 (N_26155,N_25379,N_25073);
and U26156 (N_26156,N_25593,N_25182);
and U26157 (N_26157,N_25953,N_25012);
xnor U26158 (N_26158,N_25677,N_25628);
and U26159 (N_26159,N_25480,N_25212);
or U26160 (N_26160,N_25277,N_25866);
xnor U26161 (N_26161,N_25479,N_25317);
nand U26162 (N_26162,N_25800,N_25733);
nor U26163 (N_26163,N_25415,N_25499);
nor U26164 (N_26164,N_25465,N_25517);
nor U26165 (N_26165,N_25728,N_25103);
xor U26166 (N_26166,N_25078,N_25134);
and U26167 (N_26167,N_25786,N_25219);
and U26168 (N_26168,N_25948,N_25421);
or U26169 (N_26169,N_25259,N_25679);
and U26170 (N_26170,N_25372,N_25249);
or U26171 (N_26171,N_25854,N_25993);
and U26172 (N_26172,N_25424,N_25002);
nor U26173 (N_26173,N_25542,N_25240);
xor U26174 (N_26174,N_25879,N_25837);
nand U26175 (N_26175,N_25526,N_25281);
nand U26176 (N_26176,N_25149,N_25945);
or U26177 (N_26177,N_25522,N_25501);
and U26178 (N_26178,N_25193,N_25083);
nand U26179 (N_26179,N_25573,N_25039);
xnor U26180 (N_26180,N_25218,N_25245);
nor U26181 (N_26181,N_25472,N_25334);
and U26182 (N_26182,N_25483,N_25005);
xnor U26183 (N_26183,N_25516,N_25855);
nand U26184 (N_26184,N_25497,N_25539);
nor U26185 (N_26185,N_25489,N_25146);
nor U26186 (N_26186,N_25208,N_25180);
or U26187 (N_26187,N_25342,N_25672);
and U26188 (N_26188,N_25878,N_25138);
and U26189 (N_26189,N_25385,N_25094);
or U26190 (N_26190,N_25986,N_25394);
or U26191 (N_26191,N_25325,N_25946);
or U26192 (N_26192,N_25441,N_25331);
and U26193 (N_26193,N_25393,N_25258);
nand U26194 (N_26194,N_25641,N_25108);
nor U26195 (N_26195,N_25530,N_25004);
nand U26196 (N_26196,N_25011,N_25111);
or U26197 (N_26197,N_25742,N_25314);
nor U26198 (N_26198,N_25166,N_25247);
xor U26199 (N_26199,N_25596,N_25288);
nand U26200 (N_26200,N_25403,N_25353);
or U26201 (N_26201,N_25507,N_25740);
xor U26202 (N_26202,N_25605,N_25905);
nand U26203 (N_26203,N_25209,N_25375);
nor U26204 (N_26204,N_25110,N_25274);
nor U26205 (N_26205,N_25893,N_25610);
xnor U26206 (N_26206,N_25026,N_25833);
xnor U26207 (N_26207,N_25664,N_25935);
and U26208 (N_26208,N_25674,N_25267);
xor U26209 (N_26209,N_25199,N_25703);
or U26210 (N_26210,N_25109,N_25597);
xnor U26211 (N_26211,N_25853,N_25624);
nand U26212 (N_26212,N_25257,N_25686);
or U26213 (N_26213,N_25886,N_25142);
nand U26214 (N_26214,N_25099,N_25634);
and U26215 (N_26215,N_25858,N_25827);
or U26216 (N_26216,N_25048,N_25115);
and U26217 (N_26217,N_25357,N_25279);
nor U26218 (N_26218,N_25401,N_25192);
nand U26219 (N_26219,N_25373,N_25027);
xor U26220 (N_26220,N_25406,N_25840);
or U26221 (N_26221,N_25732,N_25333);
nor U26222 (N_26222,N_25466,N_25222);
or U26223 (N_26223,N_25896,N_25119);
and U26224 (N_26224,N_25299,N_25171);
nor U26225 (N_26225,N_25459,N_25365);
nand U26226 (N_26226,N_25902,N_25711);
and U26227 (N_26227,N_25804,N_25237);
xor U26228 (N_26228,N_25660,N_25084);
nand U26229 (N_26229,N_25844,N_25330);
xnor U26230 (N_26230,N_25062,N_25432);
nor U26231 (N_26231,N_25337,N_25147);
nor U26232 (N_26232,N_25808,N_25609);
nor U26233 (N_26233,N_25775,N_25176);
and U26234 (N_26234,N_25536,N_25210);
nor U26235 (N_26235,N_25555,N_25152);
nor U26236 (N_26236,N_25057,N_25269);
or U26237 (N_26237,N_25888,N_25576);
and U26238 (N_26238,N_25998,N_25030);
or U26239 (N_26239,N_25196,N_25081);
or U26240 (N_26240,N_25243,N_25638);
xor U26241 (N_26241,N_25126,N_25753);
nand U26242 (N_26242,N_25991,N_25318);
or U26243 (N_26243,N_25089,N_25380);
or U26244 (N_26244,N_25627,N_25836);
nor U26245 (N_26245,N_25038,N_25848);
and U26246 (N_26246,N_25717,N_25469);
nand U26247 (N_26247,N_25433,N_25743);
nand U26248 (N_26248,N_25851,N_25491);
or U26249 (N_26249,N_25695,N_25698);
nand U26250 (N_26250,N_25603,N_25327);
or U26251 (N_26251,N_25551,N_25798);
nand U26252 (N_26252,N_25785,N_25534);
nor U26253 (N_26253,N_25106,N_25051);
and U26254 (N_26254,N_25736,N_25323);
nand U26255 (N_26255,N_25554,N_25120);
xor U26256 (N_26256,N_25064,N_25035);
nor U26257 (N_26257,N_25552,N_25133);
nand U26258 (N_26258,N_25835,N_25632);
or U26259 (N_26259,N_25887,N_25320);
nor U26260 (N_26260,N_25436,N_25619);
xnor U26261 (N_26261,N_25757,N_25999);
nor U26262 (N_26262,N_25395,N_25767);
nand U26263 (N_26263,N_25940,N_25477);
and U26264 (N_26264,N_25694,N_25097);
nand U26265 (N_26265,N_25282,N_25527);
or U26266 (N_26266,N_25652,N_25435);
and U26267 (N_26267,N_25790,N_25700);
and U26268 (N_26268,N_25952,N_25076);
or U26269 (N_26269,N_25644,N_25912);
or U26270 (N_26270,N_25701,N_25872);
nand U26271 (N_26271,N_25994,N_25580);
nand U26272 (N_26272,N_25794,N_25195);
and U26273 (N_26273,N_25132,N_25773);
nor U26274 (N_26274,N_25982,N_25167);
and U26275 (N_26275,N_25229,N_25929);
nor U26276 (N_26276,N_25256,N_25214);
and U26277 (N_26277,N_25157,N_25633);
nand U26278 (N_26278,N_25085,N_25688);
xnor U26279 (N_26279,N_25447,N_25559);
or U26280 (N_26280,N_25783,N_25174);
nand U26281 (N_26281,N_25316,N_25704);
nor U26282 (N_26282,N_25715,N_25930);
or U26283 (N_26283,N_25088,N_25617);
nor U26284 (N_26284,N_25608,N_25709);
nor U26285 (N_26285,N_25828,N_25014);
or U26286 (N_26286,N_25297,N_25173);
or U26287 (N_26287,N_25865,N_25482);
nand U26288 (N_26288,N_25665,N_25669);
xor U26289 (N_26289,N_25113,N_25458);
nor U26290 (N_26290,N_25791,N_25668);
xnor U26291 (N_26291,N_25016,N_25129);
nand U26292 (N_26292,N_25822,N_25226);
xor U26293 (N_26293,N_25404,N_25056);
or U26294 (N_26294,N_25074,N_25356);
nor U26295 (N_26295,N_25799,N_25985);
and U26296 (N_26296,N_25579,N_25455);
nor U26297 (N_26297,N_25091,N_25620);
or U26298 (N_26298,N_25658,N_25931);
xor U26299 (N_26299,N_25809,N_25298);
nor U26300 (N_26300,N_25781,N_25891);
or U26301 (N_26301,N_25136,N_25068);
and U26302 (N_26302,N_25233,N_25253);
nand U26303 (N_26303,N_25460,N_25198);
xor U26304 (N_26304,N_25601,N_25321);
and U26305 (N_26305,N_25852,N_25571);
or U26306 (N_26306,N_25494,N_25283);
and U26307 (N_26307,N_25719,N_25706);
nand U26308 (N_26308,N_25300,N_25186);
and U26309 (N_26309,N_25244,N_25266);
nand U26310 (N_26310,N_25659,N_25163);
nor U26311 (N_26311,N_25082,N_25586);
or U26312 (N_26312,N_25656,N_25000);
and U26313 (N_26313,N_25971,N_25560);
and U26314 (N_26314,N_25892,N_25376);
and U26315 (N_26315,N_25710,N_25054);
and U26316 (N_26316,N_25759,N_25739);
nand U26317 (N_26317,N_25956,N_25034);
nand U26318 (N_26318,N_25881,N_25661);
xor U26319 (N_26319,N_25286,N_25606);
nor U26320 (N_26320,N_25618,N_25335);
or U26321 (N_26321,N_25843,N_25558);
and U26322 (N_26322,N_25748,N_25572);
nand U26323 (N_26323,N_25184,N_25349);
xor U26324 (N_26324,N_25197,N_25919);
and U26325 (N_26325,N_25292,N_25487);
nand U26326 (N_26326,N_25118,N_25422);
nor U26327 (N_26327,N_25981,N_25236);
nor U26328 (N_26328,N_25252,N_25533);
and U26329 (N_26329,N_25990,N_25071);
and U26330 (N_26330,N_25339,N_25448);
nand U26331 (N_26331,N_25639,N_25311);
or U26332 (N_26332,N_25676,N_25577);
and U26333 (N_26333,N_25581,N_25416);
or U26334 (N_26334,N_25028,N_25202);
and U26335 (N_26335,N_25690,N_25801);
xnor U26336 (N_26336,N_25537,N_25364);
and U26337 (N_26337,N_25270,N_25796);
nand U26338 (N_26338,N_25370,N_25408);
or U26339 (N_26339,N_25655,N_25749);
nor U26340 (N_26340,N_25889,N_25397);
nor U26341 (N_26341,N_25806,N_25003);
or U26342 (N_26342,N_25795,N_25570);
xnor U26343 (N_26343,N_25098,N_25699);
and U26344 (N_26344,N_25032,N_25295);
and U26345 (N_26345,N_25220,N_25508);
or U26346 (N_26346,N_25938,N_25939);
or U26347 (N_26347,N_25780,N_25863);
xnor U26348 (N_26348,N_25541,N_25914);
and U26349 (N_26349,N_25388,N_25191);
or U26350 (N_26350,N_25072,N_25158);
nor U26351 (N_26351,N_25595,N_25456);
or U26352 (N_26352,N_25439,N_25901);
nand U26353 (N_26353,N_25834,N_25643);
xnor U26354 (N_26354,N_25883,N_25613);
or U26355 (N_26355,N_25662,N_25899);
xor U26356 (N_26356,N_25437,N_25684);
or U26357 (N_26357,N_25462,N_25438);
or U26358 (N_26358,N_25420,N_25260);
xor U26359 (N_26359,N_25937,N_25850);
nand U26360 (N_26360,N_25856,N_25391);
nand U26361 (N_26361,N_25490,N_25309);
nor U26362 (N_26362,N_25712,N_25583);
nor U26363 (N_26363,N_25453,N_25442);
nand U26364 (N_26364,N_25521,N_25148);
xor U26365 (N_26365,N_25689,N_25188);
nand U26366 (N_26366,N_25354,N_25200);
xor U26367 (N_26367,N_25488,N_25102);
xnor U26368 (N_26368,N_25629,N_25972);
and U26369 (N_26369,N_25254,N_25168);
nor U26370 (N_26370,N_25211,N_25673);
or U26371 (N_26371,N_25531,N_25607);
and U26372 (N_26372,N_25409,N_25506);
xnor U26373 (N_26373,N_25547,N_25838);
or U26374 (N_26374,N_25958,N_25248);
and U26375 (N_26375,N_25857,N_25289);
nand U26376 (N_26376,N_25348,N_25190);
xnor U26377 (N_26377,N_25153,N_25604);
xor U26378 (N_26378,N_25961,N_25968);
nor U26379 (N_26379,N_25829,N_25492);
xor U26380 (N_26380,N_25235,N_25413);
nand U26381 (N_26381,N_25750,N_25423);
nor U26382 (N_26382,N_25917,N_25975);
nor U26383 (N_26383,N_25387,N_25246);
and U26384 (N_26384,N_25995,N_25378);
or U26385 (N_26385,N_25824,N_25735);
xnor U26386 (N_26386,N_25172,N_25680);
nor U26387 (N_26387,N_25194,N_25692);
xor U26388 (N_26388,N_25691,N_25651);
nand U26389 (N_26389,N_25696,N_25429);
nor U26390 (N_26390,N_25729,N_25093);
nor U26391 (N_26391,N_25862,N_25685);
or U26392 (N_26392,N_25987,N_25265);
nand U26393 (N_26393,N_25950,N_25457);
or U26394 (N_26394,N_25486,N_25359);
nor U26395 (N_26395,N_25671,N_25529);
and U26396 (N_26396,N_25959,N_25921);
or U26397 (N_26397,N_25904,N_25121);
nor U26398 (N_26398,N_25232,N_25470);
or U26399 (N_26399,N_25069,N_25430);
or U26400 (N_26400,N_25411,N_25612);
and U26401 (N_26401,N_25885,N_25967);
nand U26402 (N_26402,N_25823,N_25683);
or U26403 (N_26403,N_25563,N_25346);
xnor U26404 (N_26404,N_25207,N_25718);
and U26405 (N_26405,N_25820,N_25726);
and U26406 (N_26406,N_25239,N_25336);
and U26407 (N_26407,N_25933,N_25065);
and U26408 (N_26408,N_25538,N_25731);
or U26409 (N_26409,N_25810,N_25842);
and U26410 (N_26410,N_25264,N_25344);
nor U26411 (N_26411,N_25880,N_25428);
nand U26412 (N_26412,N_25631,N_25475);
and U26413 (N_26413,N_25001,N_25802);
and U26414 (N_26414,N_25396,N_25594);
and U26415 (N_26415,N_25160,N_25155);
and U26416 (N_26416,N_25040,N_25481);
and U26417 (N_26417,N_25932,N_25564);
nor U26418 (N_26418,N_25776,N_25162);
nand U26419 (N_26419,N_25187,N_25362);
and U26420 (N_26420,N_25611,N_25390);
or U26421 (N_26421,N_25500,N_25941);
nor U26422 (N_26422,N_25495,N_25907);
xnor U26423 (N_26423,N_25528,N_25569);
or U26424 (N_26424,N_25752,N_25178);
and U26425 (N_26425,N_25787,N_25713);
or U26426 (N_26426,N_25151,N_25332);
and U26427 (N_26427,N_25681,N_25992);
and U26428 (N_26428,N_25008,N_25574);
nor U26429 (N_26429,N_25464,N_25926);
and U26430 (N_26430,N_25350,N_25818);
nor U26431 (N_26431,N_25238,N_25170);
xnor U26432 (N_26432,N_25216,N_25745);
nor U26433 (N_26433,N_25584,N_25788);
or U26434 (N_26434,N_25352,N_25024);
nand U26435 (N_26435,N_25358,N_25410);
and U26436 (N_26436,N_25623,N_25870);
or U26437 (N_26437,N_25550,N_25906);
nor U26438 (N_26438,N_25141,N_25565);
xor U26439 (N_26439,N_25013,N_25738);
xnor U26440 (N_26440,N_25520,N_25484);
nand U26441 (N_26441,N_25440,N_25697);
nand U26442 (N_26442,N_25626,N_25418);
nand U26443 (N_26443,N_25044,N_25588);
nand U26444 (N_26444,N_25041,N_25514);
nand U26445 (N_26445,N_25022,N_25291);
nand U26446 (N_26446,N_25018,N_25615);
or U26447 (N_26447,N_25663,N_25825);
nor U26448 (N_26448,N_25871,N_25934);
xor U26449 (N_26449,N_25868,N_25614);
xor U26450 (N_26450,N_25201,N_25949);
nand U26451 (N_26451,N_25816,N_25080);
and U26452 (N_26452,N_25723,N_25716);
or U26453 (N_26453,N_25077,N_25105);
and U26454 (N_26454,N_25493,N_25509);
or U26455 (N_26455,N_25724,N_25426);
and U26456 (N_26456,N_25312,N_25116);
and U26457 (N_26457,N_25737,N_25059);
nor U26458 (N_26458,N_25524,N_25400);
or U26459 (N_26459,N_25221,N_25280);
xnor U26460 (N_26460,N_25875,N_25772);
nand U26461 (N_26461,N_25832,N_25496);
nand U26462 (N_26462,N_25049,N_25867);
xor U26463 (N_26463,N_25997,N_25467);
xor U26464 (N_26464,N_25955,N_25287);
and U26465 (N_26465,N_25725,N_25263);
and U26466 (N_26466,N_25763,N_25861);
and U26467 (N_26467,N_25434,N_25230);
and U26468 (N_26468,N_25498,N_25637);
and U26469 (N_26469,N_25503,N_25127);
or U26470 (N_26470,N_25381,N_25075);
and U26471 (N_26471,N_25543,N_25203);
xor U26472 (N_26472,N_25727,N_25988);
or U26473 (N_26473,N_25284,N_25326);
nor U26474 (N_26474,N_25405,N_25649);
and U26475 (N_26475,N_25922,N_25648);
nand U26476 (N_26476,N_25548,N_25979);
nand U26477 (N_26477,N_25582,N_25675);
or U26478 (N_26478,N_25557,N_25747);
nand U26479 (N_26479,N_25124,N_25860);
and U26480 (N_26480,N_25859,N_25568);
xor U26481 (N_26481,N_25849,N_25139);
xnor U26482 (N_26482,N_25803,N_25066);
nand U26483 (N_26483,N_25341,N_25707);
and U26484 (N_26484,N_25451,N_25566);
xnor U26485 (N_26485,N_25137,N_25778);
nand U26486 (N_26486,N_25461,N_25189);
nand U26487 (N_26487,N_25895,N_25561);
nand U26488 (N_26488,N_25755,N_25177);
and U26489 (N_26489,N_25884,N_25771);
and U26490 (N_26490,N_25720,N_25446);
and U26491 (N_26491,N_25425,N_25485);
nor U26492 (N_26492,N_25444,N_25382);
or U26493 (N_26493,N_25793,N_25927);
nand U26494 (N_26494,N_25846,N_25667);
nand U26495 (N_26495,N_25144,N_25908);
nand U26496 (N_26496,N_25107,N_25996);
xnor U26497 (N_26497,N_25592,N_25185);
nor U26498 (N_26498,N_25900,N_25963);
nor U26499 (N_26499,N_25826,N_25670);
and U26500 (N_26500,N_25810,N_25519);
nor U26501 (N_26501,N_25808,N_25519);
and U26502 (N_26502,N_25850,N_25523);
and U26503 (N_26503,N_25738,N_25230);
and U26504 (N_26504,N_25430,N_25908);
nand U26505 (N_26505,N_25125,N_25647);
or U26506 (N_26506,N_25959,N_25376);
and U26507 (N_26507,N_25775,N_25223);
nand U26508 (N_26508,N_25694,N_25655);
or U26509 (N_26509,N_25159,N_25584);
xor U26510 (N_26510,N_25170,N_25718);
and U26511 (N_26511,N_25341,N_25811);
xor U26512 (N_26512,N_25385,N_25340);
nor U26513 (N_26513,N_25655,N_25503);
nor U26514 (N_26514,N_25512,N_25853);
nor U26515 (N_26515,N_25037,N_25741);
or U26516 (N_26516,N_25633,N_25963);
and U26517 (N_26517,N_25340,N_25037);
or U26518 (N_26518,N_25948,N_25290);
or U26519 (N_26519,N_25449,N_25258);
nand U26520 (N_26520,N_25660,N_25461);
nor U26521 (N_26521,N_25556,N_25728);
nand U26522 (N_26522,N_25237,N_25252);
nor U26523 (N_26523,N_25659,N_25083);
nand U26524 (N_26524,N_25733,N_25603);
xor U26525 (N_26525,N_25724,N_25258);
and U26526 (N_26526,N_25649,N_25420);
nor U26527 (N_26527,N_25316,N_25416);
or U26528 (N_26528,N_25895,N_25823);
xor U26529 (N_26529,N_25340,N_25976);
xor U26530 (N_26530,N_25275,N_25256);
or U26531 (N_26531,N_25300,N_25014);
and U26532 (N_26532,N_25354,N_25459);
xor U26533 (N_26533,N_25389,N_25143);
and U26534 (N_26534,N_25232,N_25714);
nor U26535 (N_26535,N_25475,N_25702);
nor U26536 (N_26536,N_25231,N_25170);
nand U26537 (N_26537,N_25869,N_25830);
nor U26538 (N_26538,N_25979,N_25403);
xnor U26539 (N_26539,N_25563,N_25793);
or U26540 (N_26540,N_25674,N_25915);
nor U26541 (N_26541,N_25597,N_25066);
xnor U26542 (N_26542,N_25185,N_25508);
xnor U26543 (N_26543,N_25449,N_25925);
nor U26544 (N_26544,N_25215,N_25287);
nand U26545 (N_26545,N_25046,N_25382);
or U26546 (N_26546,N_25341,N_25663);
and U26547 (N_26547,N_25651,N_25183);
or U26548 (N_26548,N_25811,N_25613);
nand U26549 (N_26549,N_25720,N_25759);
xor U26550 (N_26550,N_25424,N_25789);
nand U26551 (N_26551,N_25547,N_25992);
nor U26552 (N_26552,N_25081,N_25019);
nand U26553 (N_26553,N_25521,N_25265);
or U26554 (N_26554,N_25992,N_25389);
nor U26555 (N_26555,N_25368,N_25504);
xor U26556 (N_26556,N_25652,N_25543);
nor U26557 (N_26557,N_25088,N_25866);
nor U26558 (N_26558,N_25072,N_25569);
nand U26559 (N_26559,N_25318,N_25136);
nor U26560 (N_26560,N_25757,N_25218);
nor U26561 (N_26561,N_25487,N_25020);
or U26562 (N_26562,N_25710,N_25137);
nor U26563 (N_26563,N_25360,N_25994);
nor U26564 (N_26564,N_25590,N_25698);
and U26565 (N_26565,N_25508,N_25663);
nand U26566 (N_26566,N_25715,N_25234);
or U26567 (N_26567,N_25630,N_25331);
and U26568 (N_26568,N_25283,N_25657);
nand U26569 (N_26569,N_25510,N_25985);
nand U26570 (N_26570,N_25316,N_25563);
xor U26571 (N_26571,N_25220,N_25655);
nor U26572 (N_26572,N_25604,N_25365);
nor U26573 (N_26573,N_25999,N_25851);
and U26574 (N_26574,N_25307,N_25561);
or U26575 (N_26575,N_25337,N_25115);
nor U26576 (N_26576,N_25937,N_25051);
nand U26577 (N_26577,N_25764,N_25670);
nand U26578 (N_26578,N_25990,N_25548);
nor U26579 (N_26579,N_25792,N_25848);
or U26580 (N_26580,N_25998,N_25259);
nor U26581 (N_26581,N_25797,N_25752);
and U26582 (N_26582,N_25944,N_25769);
nand U26583 (N_26583,N_25729,N_25217);
nor U26584 (N_26584,N_25136,N_25185);
nor U26585 (N_26585,N_25314,N_25083);
nor U26586 (N_26586,N_25270,N_25753);
or U26587 (N_26587,N_25843,N_25972);
and U26588 (N_26588,N_25980,N_25881);
and U26589 (N_26589,N_25479,N_25979);
xor U26590 (N_26590,N_25431,N_25444);
xnor U26591 (N_26591,N_25329,N_25130);
or U26592 (N_26592,N_25189,N_25944);
nor U26593 (N_26593,N_25872,N_25561);
nor U26594 (N_26594,N_25091,N_25038);
nand U26595 (N_26595,N_25873,N_25677);
or U26596 (N_26596,N_25368,N_25178);
nor U26597 (N_26597,N_25849,N_25766);
or U26598 (N_26598,N_25771,N_25313);
xnor U26599 (N_26599,N_25022,N_25451);
xor U26600 (N_26600,N_25271,N_25226);
nor U26601 (N_26601,N_25197,N_25978);
nand U26602 (N_26602,N_25947,N_25417);
nor U26603 (N_26603,N_25981,N_25173);
and U26604 (N_26604,N_25620,N_25762);
nand U26605 (N_26605,N_25940,N_25194);
and U26606 (N_26606,N_25559,N_25021);
xnor U26607 (N_26607,N_25912,N_25330);
nand U26608 (N_26608,N_25223,N_25030);
xor U26609 (N_26609,N_25150,N_25914);
nand U26610 (N_26610,N_25839,N_25494);
or U26611 (N_26611,N_25597,N_25790);
nor U26612 (N_26612,N_25274,N_25414);
nor U26613 (N_26613,N_25975,N_25524);
xor U26614 (N_26614,N_25697,N_25438);
nand U26615 (N_26615,N_25974,N_25915);
and U26616 (N_26616,N_25013,N_25539);
nand U26617 (N_26617,N_25231,N_25466);
nor U26618 (N_26618,N_25761,N_25138);
or U26619 (N_26619,N_25212,N_25592);
nand U26620 (N_26620,N_25873,N_25250);
or U26621 (N_26621,N_25432,N_25179);
nand U26622 (N_26622,N_25232,N_25158);
and U26623 (N_26623,N_25807,N_25395);
or U26624 (N_26624,N_25755,N_25393);
or U26625 (N_26625,N_25564,N_25017);
nand U26626 (N_26626,N_25109,N_25419);
xor U26627 (N_26627,N_25029,N_25760);
nand U26628 (N_26628,N_25983,N_25111);
nor U26629 (N_26629,N_25964,N_25678);
nor U26630 (N_26630,N_25353,N_25882);
or U26631 (N_26631,N_25483,N_25880);
and U26632 (N_26632,N_25183,N_25137);
or U26633 (N_26633,N_25717,N_25570);
or U26634 (N_26634,N_25948,N_25893);
xor U26635 (N_26635,N_25078,N_25057);
nor U26636 (N_26636,N_25835,N_25272);
xor U26637 (N_26637,N_25178,N_25069);
nand U26638 (N_26638,N_25922,N_25264);
xnor U26639 (N_26639,N_25945,N_25385);
nand U26640 (N_26640,N_25410,N_25097);
and U26641 (N_26641,N_25774,N_25718);
or U26642 (N_26642,N_25754,N_25835);
xor U26643 (N_26643,N_25262,N_25311);
nand U26644 (N_26644,N_25784,N_25364);
nand U26645 (N_26645,N_25961,N_25882);
or U26646 (N_26646,N_25881,N_25153);
xnor U26647 (N_26647,N_25701,N_25670);
nor U26648 (N_26648,N_25133,N_25260);
nand U26649 (N_26649,N_25428,N_25329);
and U26650 (N_26650,N_25112,N_25379);
or U26651 (N_26651,N_25720,N_25590);
nor U26652 (N_26652,N_25889,N_25842);
xnor U26653 (N_26653,N_25253,N_25611);
nor U26654 (N_26654,N_25889,N_25876);
nor U26655 (N_26655,N_25526,N_25802);
nand U26656 (N_26656,N_25090,N_25736);
nand U26657 (N_26657,N_25903,N_25156);
nand U26658 (N_26658,N_25380,N_25963);
nand U26659 (N_26659,N_25040,N_25049);
nand U26660 (N_26660,N_25846,N_25687);
and U26661 (N_26661,N_25963,N_25472);
nand U26662 (N_26662,N_25402,N_25083);
or U26663 (N_26663,N_25934,N_25150);
nand U26664 (N_26664,N_25806,N_25674);
nand U26665 (N_26665,N_25242,N_25089);
or U26666 (N_26666,N_25715,N_25782);
nand U26667 (N_26667,N_25014,N_25938);
nand U26668 (N_26668,N_25311,N_25738);
or U26669 (N_26669,N_25405,N_25938);
or U26670 (N_26670,N_25921,N_25665);
xor U26671 (N_26671,N_25918,N_25939);
or U26672 (N_26672,N_25560,N_25784);
nor U26673 (N_26673,N_25843,N_25049);
nor U26674 (N_26674,N_25676,N_25354);
nor U26675 (N_26675,N_25967,N_25102);
or U26676 (N_26676,N_25174,N_25085);
nand U26677 (N_26677,N_25471,N_25945);
xnor U26678 (N_26678,N_25778,N_25479);
nor U26679 (N_26679,N_25181,N_25766);
nor U26680 (N_26680,N_25909,N_25791);
nor U26681 (N_26681,N_25042,N_25682);
nor U26682 (N_26682,N_25991,N_25044);
xnor U26683 (N_26683,N_25073,N_25238);
nand U26684 (N_26684,N_25364,N_25724);
or U26685 (N_26685,N_25264,N_25622);
xnor U26686 (N_26686,N_25744,N_25500);
and U26687 (N_26687,N_25375,N_25153);
nor U26688 (N_26688,N_25224,N_25887);
and U26689 (N_26689,N_25476,N_25542);
xnor U26690 (N_26690,N_25074,N_25613);
or U26691 (N_26691,N_25500,N_25487);
or U26692 (N_26692,N_25279,N_25364);
or U26693 (N_26693,N_25847,N_25907);
or U26694 (N_26694,N_25503,N_25536);
and U26695 (N_26695,N_25787,N_25717);
or U26696 (N_26696,N_25857,N_25299);
xor U26697 (N_26697,N_25172,N_25299);
and U26698 (N_26698,N_25870,N_25625);
xnor U26699 (N_26699,N_25019,N_25180);
nand U26700 (N_26700,N_25668,N_25834);
and U26701 (N_26701,N_25996,N_25474);
xor U26702 (N_26702,N_25688,N_25161);
nor U26703 (N_26703,N_25263,N_25601);
nor U26704 (N_26704,N_25145,N_25010);
nand U26705 (N_26705,N_25839,N_25766);
nor U26706 (N_26706,N_25137,N_25919);
nor U26707 (N_26707,N_25364,N_25672);
nand U26708 (N_26708,N_25014,N_25843);
and U26709 (N_26709,N_25438,N_25130);
nand U26710 (N_26710,N_25118,N_25190);
and U26711 (N_26711,N_25310,N_25773);
xor U26712 (N_26712,N_25061,N_25023);
nand U26713 (N_26713,N_25147,N_25778);
nand U26714 (N_26714,N_25474,N_25600);
and U26715 (N_26715,N_25507,N_25196);
xor U26716 (N_26716,N_25353,N_25110);
nor U26717 (N_26717,N_25586,N_25649);
nand U26718 (N_26718,N_25014,N_25957);
xor U26719 (N_26719,N_25054,N_25248);
or U26720 (N_26720,N_25272,N_25418);
nor U26721 (N_26721,N_25307,N_25930);
and U26722 (N_26722,N_25918,N_25399);
xor U26723 (N_26723,N_25346,N_25384);
and U26724 (N_26724,N_25333,N_25738);
nand U26725 (N_26725,N_25368,N_25947);
nand U26726 (N_26726,N_25873,N_25864);
and U26727 (N_26727,N_25410,N_25420);
nor U26728 (N_26728,N_25096,N_25105);
and U26729 (N_26729,N_25756,N_25790);
or U26730 (N_26730,N_25621,N_25819);
nand U26731 (N_26731,N_25320,N_25909);
or U26732 (N_26732,N_25699,N_25134);
nor U26733 (N_26733,N_25067,N_25381);
xnor U26734 (N_26734,N_25126,N_25997);
and U26735 (N_26735,N_25745,N_25593);
and U26736 (N_26736,N_25855,N_25395);
and U26737 (N_26737,N_25880,N_25977);
nor U26738 (N_26738,N_25219,N_25050);
nor U26739 (N_26739,N_25520,N_25418);
xor U26740 (N_26740,N_25843,N_25664);
nand U26741 (N_26741,N_25541,N_25368);
xor U26742 (N_26742,N_25008,N_25898);
or U26743 (N_26743,N_25400,N_25692);
and U26744 (N_26744,N_25513,N_25672);
xor U26745 (N_26745,N_25365,N_25949);
or U26746 (N_26746,N_25438,N_25428);
and U26747 (N_26747,N_25472,N_25344);
nand U26748 (N_26748,N_25771,N_25503);
xor U26749 (N_26749,N_25846,N_25478);
nor U26750 (N_26750,N_25759,N_25329);
and U26751 (N_26751,N_25100,N_25085);
nand U26752 (N_26752,N_25789,N_25347);
nand U26753 (N_26753,N_25380,N_25343);
xnor U26754 (N_26754,N_25854,N_25655);
and U26755 (N_26755,N_25081,N_25172);
xnor U26756 (N_26756,N_25801,N_25513);
xor U26757 (N_26757,N_25186,N_25321);
xor U26758 (N_26758,N_25000,N_25478);
or U26759 (N_26759,N_25580,N_25973);
nor U26760 (N_26760,N_25837,N_25495);
and U26761 (N_26761,N_25995,N_25262);
nand U26762 (N_26762,N_25922,N_25445);
nor U26763 (N_26763,N_25356,N_25669);
nand U26764 (N_26764,N_25443,N_25858);
and U26765 (N_26765,N_25358,N_25178);
or U26766 (N_26766,N_25236,N_25650);
nor U26767 (N_26767,N_25985,N_25638);
and U26768 (N_26768,N_25825,N_25840);
and U26769 (N_26769,N_25847,N_25927);
xor U26770 (N_26770,N_25965,N_25959);
and U26771 (N_26771,N_25435,N_25331);
or U26772 (N_26772,N_25135,N_25924);
nand U26773 (N_26773,N_25568,N_25165);
nand U26774 (N_26774,N_25335,N_25403);
xor U26775 (N_26775,N_25742,N_25462);
nand U26776 (N_26776,N_25328,N_25629);
or U26777 (N_26777,N_25962,N_25224);
or U26778 (N_26778,N_25729,N_25121);
nand U26779 (N_26779,N_25109,N_25773);
or U26780 (N_26780,N_25244,N_25471);
nand U26781 (N_26781,N_25490,N_25974);
nor U26782 (N_26782,N_25076,N_25871);
xor U26783 (N_26783,N_25376,N_25499);
or U26784 (N_26784,N_25908,N_25739);
xnor U26785 (N_26785,N_25166,N_25151);
and U26786 (N_26786,N_25868,N_25391);
or U26787 (N_26787,N_25892,N_25016);
or U26788 (N_26788,N_25205,N_25485);
or U26789 (N_26789,N_25345,N_25586);
or U26790 (N_26790,N_25437,N_25150);
or U26791 (N_26791,N_25575,N_25904);
nor U26792 (N_26792,N_25770,N_25675);
or U26793 (N_26793,N_25246,N_25315);
nor U26794 (N_26794,N_25068,N_25668);
nor U26795 (N_26795,N_25951,N_25089);
nor U26796 (N_26796,N_25259,N_25757);
nand U26797 (N_26797,N_25777,N_25830);
or U26798 (N_26798,N_25904,N_25328);
nand U26799 (N_26799,N_25555,N_25118);
nor U26800 (N_26800,N_25211,N_25844);
nand U26801 (N_26801,N_25271,N_25332);
nor U26802 (N_26802,N_25486,N_25983);
and U26803 (N_26803,N_25260,N_25331);
or U26804 (N_26804,N_25419,N_25040);
and U26805 (N_26805,N_25164,N_25159);
and U26806 (N_26806,N_25663,N_25013);
xnor U26807 (N_26807,N_25786,N_25768);
and U26808 (N_26808,N_25427,N_25445);
or U26809 (N_26809,N_25727,N_25385);
nor U26810 (N_26810,N_25755,N_25193);
and U26811 (N_26811,N_25270,N_25488);
and U26812 (N_26812,N_25040,N_25483);
xnor U26813 (N_26813,N_25044,N_25150);
xnor U26814 (N_26814,N_25996,N_25105);
nor U26815 (N_26815,N_25546,N_25326);
nand U26816 (N_26816,N_25050,N_25294);
nor U26817 (N_26817,N_25789,N_25003);
xnor U26818 (N_26818,N_25483,N_25970);
nor U26819 (N_26819,N_25642,N_25439);
nand U26820 (N_26820,N_25870,N_25088);
and U26821 (N_26821,N_25715,N_25468);
xnor U26822 (N_26822,N_25137,N_25177);
nor U26823 (N_26823,N_25444,N_25455);
xor U26824 (N_26824,N_25088,N_25618);
or U26825 (N_26825,N_25394,N_25785);
xnor U26826 (N_26826,N_25326,N_25483);
nor U26827 (N_26827,N_25397,N_25137);
or U26828 (N_26828,N_25499,N_25925);
and U26829 (N_26829,N_25418,N_25138);
and U26830 (N_26830,N_25594,N_25986);
nor U26831 (N_26831,N_25730,N_25006);
xnor U26832 (N_26832,N_25462,N_25653);
and U26833 (N_26833,N_25651,N_25177);
nor U26834 (N_26834,N_25135,N_25638);
and U26835 (N_26835,N_25740,N_25378);
or U26836 (N_26836,N_25041,N_25844);
xor U26837 (N_26837,N_25110,N_25686);
nor U26838 (N_26838,N_25148,N_25771);
and U26839 (N_26839,N_25197,N_25448);
and U26840 (N_26840,N_25626,N_25020);
or U26841 (N_26841,N_25248,N_25134);
nand U26842 (N_26842,N_25559,N_25173);
xnor U26843 (N_26843,N_25704,N_25946);
nand U26844 (N_26844,N_25009,N_25698);
nand U26845 (N_26845,N_25816,N_25510);
nor U26846 (N_26846,N_25012,N_25857);
nor U26847 (N_26847,N_25436,N_25615);
xnor U26848 (N_26848,N_25859,N_25693);
or U26849 (N_26849,N_25982,N_25595);
and U26850 (N_26850,N_25862,N_25369);
nand U26851 (N_26851,N_25351,N_25162);
and U26852 (N_26852,N_25791,N_25953);
nor U26853 (N_26853,N_25901,N_25678);
or U26854 (N_26854,N_25372,N_25511);
nor U26855 (N_26855,N_25791,N_25048);
and U26856 (N_26856,N_25422,N_25031);
nand U26857 (N_26857,N_25984,N_25034);
or U26858 (N_26858,N_25947,N_25245);
or U26859 (N_26859,N_25182,N_25099);
nand U26860 (N_26860,N_25259,N_25795);
xor U26861 (N_26861,N_25836,N_25773);
and U26862 (N_26862,N_25077,N_25303);
nor U26863 (N_26863,N_25577,N_25759);
nand U26864 (N_26864,N_25154,N_25843);
nor U26865 (N_26865,N_25758,N_25349);
nor U26866 (N_26866,N_25997,N_25100);
or U26867 (N_26867,N_25250,N_25016);
nor U26868 (N_26868,N_25474,N_25025);
xor U26869 (N_26869,N_25478,N_25815);
or U26870 (N_26870,N_25089,N_25903);
nor U26871 (N_26871,N_25058,N_25561);
and U26872 (N_26872,N_25003,N_25907);
or U26873 (N_26873,N_25517,N_25811);
and U26874 (N_26874,N_25678,N_25618);
xnor U26875 (N_26875,N_25624,N_25662);
or U26876 (N_26876,N_25354,N_25654);
xnor U26877 (N_26877,N_25553,N_25408);
or U26878 (N_26878,N_25439,N_25372);
xor U26879 (N_26879,N_25800,N_25840);
or U26880 (N_26880,N_25817,N_25048);
or U26881 (N_26881,N_25549,N_25626);
or U26882 (N_26882,N_25188,N_25348);
or U26883 (N_26883,N_25908,N_25355);
xnor U26884 (N_26884,N_25997,N_25998);
and U26885 (N_26885,N_25526,N_25183);
or U26886 (N_26886,N_25679,N_25206);
nand U26887 (N_26887,N_25042,N_25689);
and U26888 (N_26888,N_25891,N_25882);
xnor U26889 (N_26889,N_25497,N_25223);
nand U26890 (N_26890,N_25645,N_25497);
or U26891 (N_26891,N_25146,N_25388);
or U26892 (N_26892,N_25737,N_25553);
or U26893 (N_26893,N_25404,N_25934);
nand U26894 (N_26894,N_25625,N_25229);
nor U26895 (N_26895,N_25894,N_25395);
xor U26896 (N_26896,N_25228,N_25472);
xor U26897 (N_26897,N_25402,N_25233);
and U26898 (N_26898,N_25753,N_25622);
and U26899 (N_26899,N_25813,N_25641);
xnor U26900 (N_26900,N_25674,N_25602);
or U26901 (N_26901,N_25267,N_25436);
nand U26902 (N_26902,N_25150,N_25251);
nor U26903 (N_26903,N_25139,N_25144);
xnor U26904 (N_26904,N_25686,N_25979);
nor U26905 (N_26905,N_25681,N_25978);
and U26906 (N_26906,N_25478,N_25627);
nand U26907 (N_26907,N_25528,N_25346);
or U26908 (N_26908,N_25146,N_25295);
and U26909 (N_26909,N_25767,N_25829);
and U26910 (N_26910,N_25614,N_25058);
and U26911 (N_26911,N_25898,N_25886);
nand U26912 (N_26912,N_25285,N_25605);
and U26913 (N_26913,N_25140,N_25531);
and U26914 (N_26914,N_25706,N_25083);
nand U26915 (N_26915,N_25217,N_25889);
or U26916 (N_26916,N_25005,N_25573);
xnor U26917 (N_26917,N_25145,N_25489);
and U26918 (N_26918,N_25548,N_25196);
nand U26919 (N_26919,N_25792,N_25300);
or U26920 (N_26920,N_25543,N_25404);
nor U26921 (N_26921,N_25608,N_25770);
or U26922 (N_26922,N_25865,N_25840);
nor U26923 (N_26923,N_25366,N_25227);
nand U26924 (N_26924,N_25301,N_25762);
nor U26925 (N_26925,N_25599,N_25976);
and U26926 (N_26926,N_25679,N_25997);
nor U26927 (N_26927,N_25738,N_25547);
or U26928 (N_26928,N_25467,N_25551);
xor U26929 (N_26929,N_25688,N_25274);
or U26930 (N_26930,N_25030,N_25555);
nor U26931 (N_26931,N_25743,N_25331);
nor U26932 (N_26932,N_25496,N_25431);
nand U26933 (N_26933,N_25140,N_25651);
or U26934 (N_26934,N_25911,N_25228);
nor U26935 (N_26935,N_25984,N_25832);
nor U26936 (N_26936,N_25810,N_25176);
nand U26937 (N_26937,N_25419,N_25967);
or U26938 (N_26938,N_25285,N_25415);
xor U26939 (N_26939,N_25748,N_25230);
xnor U26940 (N_26940,N_25148,N_25570);
and U26941 (N_26941,N_25628,N_25244);
xor U26942 (N_26942,N_25319,N_25727);
xnor U26943 (N_26943,N_25467,N_25035);
nand U26944 (N_26944,N_25358,N_25585);
xor U26945 (N_26945,N_25472,N_25908);
and U26946 (N_26946,N_25754,N_25856);
and U26947 (N_26947,N_25022,N_25879);
nor U26948 (N_26948,N_25231,N_25367);
and U26949 (N_26949,N_25000,N_25262);
xor U26950 (N_26950,N_25416,N_25095);
or U26951 (N_26951,N_25234,N_25777);
nand U26952 (N_26952,N_25414,N_25527);
xnor U26953 (N_26953,N_25752,N_25048);
nor U26954 (N_26954,N_25831,N_25567);
or U26955 (N_26955,N_25255,N_25270);
xor U26956 (N_26956,N_25079,N_25790);
nor U26957 (N_26957,N_25493,N_25888);
and U26958 (N_26958,N_25044,N_25637);
and U26959 (N_26959,N_25931,N_25572);
xnor U26960 (N_26960,N_25404,N_25751);
nand U26961 (N_26961,N_25661,N_25356);
or U26962 (N_26962,N_25853,N_25646);
nand U26963 (N_26963,N_25475,N_25296);
xor U26964 (N_26964,N_25792,N_25680);
xor U26965 (N_26965,N_25568,N_25896);
nor U26966 (N_26966,N_25082,N_25452);
nand U26967 (N_26967,N_25319,N_25102);
xor U26968 (N_26968,N_25521,N_25031);
and U26969 (N_26969,N_25420,N_25730);
xor U26970 (N_26970,N_25355,N_25353);
and U26971 (N_26971,N_25019,N_25490);
or U26972 (N_26972,N_25988,N_25821);
and U26973 (N_26973,N_25648,N_25737);
nor U26974 (N_26974,N_25201,N_25189);
nand U26975 (N_26975,N_25307,N_25253);
nand U26976 (N_26976,N_25283,N_25239);
and U26977 (N_26977,N_25147,N_25053);
and U26978 (N_26978,N_25257,N_25165);
or U26979 (N_26979,N_25607,N_25800);
and U26980 (N_26980,N_25072,N_25615);
or U26981 (N_26981,N_25092,N_25601);
and U26982 (N_26982,N_25458,N_25512);
nor U26983 (N_26983,N_25387,N_25043);
or U26984 (N_26984,N_25695,N_25269);
xnor U26985 (N_26985,N_25124,N_25757);
nor U26986 (N_26986,N_25026,N_25864);
or U26987 (N_26987,N_25821,N_25625);
or U26988 (N_26988,N_25398,N_25118);
or U26989 (N_26989,N_25224,N_25035);
nor U26990 (N_26990,N_25431,N_25571);
nor U26991 (N_26991,N_25191,N_25265);
nand U26992 (N_26992,N_25434,N_25588);
xor U26993 (N_26993,N_25664,N_25944);
nand U26994 (N_26994,N_25251,N_25587);
or U26995 (N_26995,N_25224,N_25516);
nand U26996 (N_26996,N_25444,N_25174);
nand U26997 (N_26997,N_25544,N_25916);
and U26998 (N_26998,N_25874,N_25521);
and U26999 (N_26999,N_25183,N_25799);
or U27000 (N_27000,N_26960,N_26196);
xnor U27001 (N_27001,N_26727,N_26414);
or U27002 (N_27002,N_26470,N_26895);
nor U27003 (N_27003,N_26569,N_26233);
and U27004 (N_27004,N_26086,N_26862);
nor U27005 (N_27005,N_26833,N_26326);
nand U27006 (N_27006,N_26530,N_26402);
and U27007 (N_27007,N_26867,N_26579);
or U27008 (N_27008,N_26774,N_26445);
nor U27009 (N_27009,N_26949,N_26693);
xnor U27010 (N_27010,N_26410,N_26267);
and U27011 (N_27011,N_26930,N_26487);
or U27012 (N_27012,N_26108,N_26708);
or U27013 (N_27013,N_26134,N_26559);
nand U27014 (N_27014,N_26151,N_26453);
xor U27015 (N_27015,N_26551,N_26713);
xnor U27016 (N_27016,N_26666,N_26981);
or U27017 (N_27017,N_26678,N_26244);
or U27018 (N_27018,N_26316,N_26481);
and U27019 (N_27019,N_26679,N_26576);
or U27020 (N_27020,N_26815,N_26088);
xnor U27021 (N_27021,N_26804,N_26103);
nand U27022 (N_27022,N_26923,N_26442);
nand U27023 (N_27023,N_26548,N_26312);
and U27024 (N_27024,N_26615,N_26726);
nor U27025 (N_27025,N_26252,N_26148);
xnor U27026 (N_27026,N_26078,N_26992);
and U27027 (N_27027,N_26536,N_26502);
nor U27028 (N_27028,N_26877,N_26075);
nand U27029 (N_27029,N_26011,N_26879);
or U27030 (N_27030,N_26717,N_26213);
or U27031 (N_27031,N_26076,N_26753);
nor U27032 (N_27032,N_26800,N_26786);
and U27033 (N_27033,N_26578,N_26712);
nor U27034 (N_27034,N_26023,N_26262);
or U27035 (N_27035,N_26232,N_26953);
xnor U27036 (N_27036,N_26157,N_26235);
nor U27037 (N_27037,N_26639,N_26967);
nor U27038 (N_27038,N_26869,N_26614);
nor U27039 (N_27039,N_26117,N_26513);
or U27040 (N_27040,N_26896,N_26126);
nor U27041 (N_27041,N_26831,N_26253);
xnor U27042 (N_27042,N_26610,N_26936);
xor U27043 (N_27043,N_26849,N_26847);
or U27044 (N_27044,N_26689,N_26227);
xnor U27045 (N_27045,N_26258,N_26566);
and U27046 (N_27046,N_26655,N_26072);
and U27047 (N_27047,N_26411,N_26390);
nor U27048 (N_27048,N_26926,N_26854);
nor U27049 (N_27049,N_26781,N_26618);
xnor U27050 (N_27050,N_26684,N_26856);
nor U27051 (N_27051,N_26860,N_26226);
xor U27052 (N_27052,N_26797,N_26394);
nor U27053 (N_27053,N_26575,N_26826);
nor U27054 (N_27054,N_26754,N_26527);
and U27055 (N_27055,N_26208,N_26845);
xor U27056 (N_27056,N_26902,N_26698);
nor U27057 (N_27057,N_26083,N_26526);
or U27058 (N_27058,N_26280,N_26700);
nand U27059 (N_27059,N_26249,N_26324);
nor U27060 (N_27060,N_26870,N_26829);
or U27061 (N_27061,N_26626,N_26984);
or U27062 (N_27062,N_26522,N_26447);
xor U27063 (N_27063,N_26756,N_26416);
or U27064 (N_27064,N_26941,N_26118);
nand U27065 (N_27065,N_26670,N_26517);
or U27066 (N_27066,N_26971,N_26676);
and U27067 (N_27067,N_26285,N_26003);
xor U27068 (N_27068,N_26444,N_26738);
nand U27069 (N_27069,N_26799,N_26934);
or U27070 (N_27070,N_26143,N_26054);
or U27071 (N_27071,N_26940,N_26180);
xnor U27072 (N_27072,N_26729,N_26682);
nor U27073 (N_27073,N_26466,N_26939);
or U27074 (N_27074,N_26874,N_26749);
xor U27075 (N_27075,N_26292,N_26459);
and U27076 (N_27076,N_26355,N_26909);
nor U27077 (N_27077,N_26040,N_26777);
or U27078 (N_27078,N_26281,N_26325);
nand U27079 (N_27079,N_26454,N_26150);
xnor U27080 (N_27080,N_26509,N_26376);
or U27081 (N_27081,N_26375,N_26135);
nor U27082 (N_27082,N_26813,N_26979);
xor U27083 (N_27083,N_26773,N_26601);
nand U27084 (N_27084,N_26987,N_26273);
xnor U27085 (N_27085,N_26049,N_26499);
or U27086 (N_27086,N_26819,N_26635);
and U27087 (N_27087,N_26767,N_26825);
or U27088 (N_27088,N_26776,N_26131);
nand U27089 (N_27089,N_26065,N_26858);
and U27090 (N_27090,N_26769,N_26332);
or U27091 (N_27091,N_26866,N_26068);
and U27092 (N_27092,N_26495,N_26932);
or U27093 (N_27093,N_26945,N_26897);
nor U27094 (N_27094,N_26133,N_26523);
and U27095 (N_27095,N_26525,N_26090);
and U27096 (N_27096,N_26784,N_26184);
or U27097 (N_27097,N_26174,N_26837);
xor U27098 (N_27098,N_26384,N_26374);
nor U27099 (N_27099,N_26972,N_26101);
and U27100 (N_27100,N_26515,N_26623);
nand U27101 (N_27101,N_26082,N_26707);
or U27102 (N_27102,N_26508,N_26467);
and U27103 (N_27103,N_26603,N_26853);
or U27104 (N_27104,N_26295,N_26588);
xnor U27105 (N_27105,N_26261,N_26658);
or U27106 (N_27106,N_26356,N_26197);
and U27107 (N_27107,N_26287,N_26921);
nor U27108 (N_27108,N_26299,N_26427);
or U27109 (N_27109,N_26516,N_26889);
and U27110 (N_27110,N_26032,N_26608);
nor U27111 (N_27111,N_26757,N_26391);
nor U27112 (N_27112,N_26051,N_26720);
and U27113 (N_27113,N_26547,N_26912);
or U27114 (N_27114,N_26152,N_26824);
nand U27115 (N_27115,N_26549,N_26340);
nor U27116 (N_27116,N_26600,N_26059);
nand U27117 (N_27117,N_26359,N_26307);
xnor U27118 (N_27118,N_26571,N_26794);
nand U27119 (N_27119,N_26604,N_26611);
nor U27120 (N_27120,N_26802,N_26367);
nor U27121 (N_27121,N_26048,N_26296);
or U27122 (N_27122,N_26890,N_26851);
nand U27123 (N_27123,N_26675,N_26449);
and U27124 (N_27124,N_26621,N_26345);
and U27125 (N_27125,N_26104,N_26424);
or U27126 (N_27126,N_26452,N_26216);
nand U27127 (N_27127,N_26472,N_26099);
and U27128 (N_27128,N_26153,N_26801);
nor U27129 (N_27129,N_26683,N_26925);
xor U27130 (N_27130,N_26938,N_26422);
nor U27131 (N_27131,N_26719,N_26328);
xnor U27132 (N_27132,N_26861,N_26412);
or U27133 (N_27133,N_26415,N_26451);
and U27134 (N_27134,N_26263,N_26742);
and U27135 (N_27135,N_26583,N_26961);
nand U27136 (N_27136,N_26311,N_26545);
nand U27137 (N_27137,N_26033,N_26916);
nor U27138 (N_27138,N_26266,N_26024);
nand U27139 (N_27139,N_26620,N_26834);
xnor U27140 (N_27140,N_26747,N_26306);
nand U27141 (N_27141,N_26910,N_26218);
or U27142 (N_27142,N_26012,N_26725);
nor U27143 (N_27143,N_26373,N_26816);
nand U27144 (N_27144,N_26061,N_26294);
or U27145 (N_27145,N_26095,N_26277);
nor U27146 (N_27146,N_26970,N_26085);
xnor U27147 (N_27147,N_26031,N_26360);
nand U27148 (N_27148,N_26577,N_26602);
nor U27149 (N_27149,N_26900,N_26557);
and U27150 (N_27150,N_26385,N_26714);
xnor U27151 (N_27151,N_26546,N_26388);
or U27152 (N_27152,N_26805,N_26279);
nor U27153 (N_27153,N_26366,N_26172);
nand U27154 (N_27154,N_26187,N_26543);
nand U27155 (N_27155,N_26195,N_26885);
or U27156 (N_27156,N_26063,N_26671);
nor U27157 (N_27157,N_26413,N_26111);
xnor U27158 (N_27158,N_26149,N_26673);
nor U27159 (N_27159,N_26944,N_26840);
nor U27160 (N_27160,N_26483,N_26990);
xnor U27161 (N_27161,N_26759,N_26034);
and U27162 (N_27162,N_26486,N_26175);
nand U27163 (N_27163,N_26370,N_26962);
or U27164 (N_27164,N_26915,N_26511);
nand U27165 (N_27165,N_26162,N_26798);
nand U27166 (N_27166,N_26762,N_26336);
xor U27167 (N_27167,N_26419,N_26275);
nor U27168 (N_27168,N_26692,N_26768);
or U27169 (N_27169,N_26737,N_26230);
xnor U27170 (N_27170,N_26349,N_26124);
nor U27171 (N_27171,N_26521,N_26329);
xor U27172 (N_27172,N_26144,N_26044);
nand U27173 (N_27173,N_26497,N_26734);
and U27174 (N_27174,N_26901,N_26562);
xor U27175 (N_27175,N_26080,N_26793);
nand U27176 (N_27176,N_26787,N_26116);
and U27177 (N_27177,N_26919,N_26455);
nor U27178 (N_27178,N_26421,N_26544);
and U27179 (N_27179,N_26141,N_26705);
nand U27180 (N_27180,N_26745,N_26221);
or U27181 (N_27181,N_26430,N_26036);
nor U27182 (N_27182,N_26037,N_26047);
and U27183 (N_27183,N_26672,N_26848);
and U27184 (N_27184,N_26920,N_26386);
nand U27185 (N_27185,N_26129,N_26617);
nor U27186 (N_27186,N_26701,N_26400);
nand U27187 (N_27187,N_26631,N_26137);
nor U27188 (N_27188,N_26492,N_26409);
nor U27189 (N_27189,N_26441,N_26660);
nand U27190 (N_27190,N_26105,N_26718);
nand U27191 (N_27191,N_26022,N_26166);
or U27192 (N_27192,N_26758,N_26641);
nor U27193 (N_27193,N_26209,N_26790);
nor U27194 (N_27194,N_26703,N_26810);
or U27195 (N_27195,N_26573,N_26835);
or U27196 (N_27196,N_26322,N_26590);
xnor U27197 (N_27197,N_26724,N_26035);
and U27198 (N_27198,N_26778,N_26956);
or U27199 (N_27199,N_26943,N_26711);
and U27200 (N_27200,N_26403,N_26320);
nor U27201 (N_27201,N_26928,N_26659);
nand U27202 (N_27202,N_26731,N_26688);
and U27203 (N_27203,N_26250,N_26857);
nor U27204 (N_27204,N_26437,N_26062);
nand U27205 (N_27205,N_26598,N_26438);
xnor U27206 (N_27206,N_26461,N_26982);
xor U27207 (N_27207,N_26665,N_26709);
xor U27208 (N_27208,N_26908,N_26529);
xnor U27209 (N_27209,N_26130,N_26746);
or U27210 (N_27210,N_26818,N_26382);
and U27211 (N_27211,N_26796,N_26690);
nand U27212 (N_27212,N_26236,N_26334);
and U27213 (N_27213,N_26188,N_26779);
or U27214 (N_27214,N_26782,N_26428);
and U27215 (N_27215,N_26788,N_26343);
and U27216 (N_27216,N_26183,N_26630);
nand U27217 (N_27217,N_26891,N_26272);
nand U27218 (N_27218,N_26638,N_26323);
nand U27219 (N_27219,N_26850,N_26182);
nor U27220 (N_27220,N_26247,N_26558);
or U27221 (N_27221,N_26740,N_26138);
xor U27222 (N_27222,N_26168,N_26446);
xnor U27223 (N_27223,N_26214,N_26278);
xor U27224 (N_27224,N_26844,N_26217);
nor U27225 (N_27225,N_26222,N_26286);
and U27226 (N_27226,N_26114,N_26715);
or U27227 (N_27227,N_26219,N_26903);
nor U27228 (N_27228,N_26026,N_26479);
and U27229 (N_27229,N_26491,N_26297);
xor U27230 (N_27230,N_26827,N_26643);
nand U27231 (N_27231,N_26674,N_26518);
or U27232 (N_27232,N_26496,N_26539);
xnor U27233 (N_27233,N_26636,N_26234);
nor U27234 (N_27234,N_26308,N_26426);
xor U27235 (N_27235,N_26785,N_26974);
nor U27236 (N_27236,N_26282,N_26046);
and U27237 (N_27237,N_26755,N_26770);
xnor U27238 (N_27238,N_26434,N_26021);
xnor U27239 (N_27239,N_26121,N_26339);
nand U27240 (N_27240,N_26716,N_26884);
or U27241 (N_27241,N_26830,N_26586);
xor U27242 (N_27242,N_26224,N_26730);
nor U27243 (N_27243,N_26791,N_26161);
nand U27244 (N_27244,N_26506,N_26504);
or U27245 (N_27245,N_26457,N_26667);
and U27246 (N_27246,N_26493,N_26302);
nor U27247 (N_27247,N_26880,N_26211);
nor U27248 (N_27248,N_26288,N_26741);
nor U27249 (N_27249,N_26728,N_26927);
nor U27250 (N_27250,N_26190,N_26119);
or U27251 (N_27251,N_26071,N_26397);
xnor U27252 (N_27252,N_26165,N_26110);
or U27253 (N_27253,N_26352,N_26680);
nor U27254 (N_27254,N_26193,N_26488);
and U27255 (N_27255,N_26098,N_26220);
xor U27256 (N_27256,N_26045,N_26875);
or U27257 (N_27257,N_26652,N_26647);
and U27258 (N_27258,N_26351,N_26396);
nor U27259 (N_27259,N_26186,N_26806);
and U27260 (N_27260,N_26561,N_26425);
and U27261 (N_27261,N_26589,N_26337);
nor U27262 (N_27262,N_26079,N_26534);
or U27263 (N_27263,N_26836,N_26661);
xnor U27264 (N_27264,N_26871,N_26644);
nand U27265 (N_27265,N_26330,N_26669);
xnor U27266 (N_27266,N_26887,N_26807);
nor U27267 (N_27267,N_26008,N_26494);
nand U27268 (N_27268,N_26191,N_26176);
nor U27269 (N_27269,N_26533,N_26448);
xnor U27270 (N_27270,N_26238,N_26087);
or U27271 (N_27271,N_26399,N_26556);
nand U27272 (N_27272,N_26993,N_26899);
or U27273 (N_27273,N_26542,N_26505);
nand U27274 (N_27274,N_26568,N_26260);
nor U27275 (N_27275,N_26458,N_26321);
nor U27276 (N_27276,N_26996,N_26812);
nand U27277 (N_27277,N_26911,N_26274);
and U27278 (N_27278,N_26301,N_26520);
or U27279 (N_27279,N_26398,N_26538);
xnor U27280 (N_27280,N_26364,N_26016);
or U27281 (N_27281,N_26064,N_26607);
xnor U27282 (N_27282,N_26907,N_26464);
nor U27283 (N_27283,N_26942,N_26735);
xnor U27284 (N_27284,N_26239,N_26156);
and U27285 (N_27285,N_26648,N_26145);
xor U27286 (N_27286,N_26937,N_26991);
and U27287 (N_27287,N_26084,N_26803);
or U27288 (N_27288,N_26846,N_26722);
or U27289 (N_27289,N_26317,N_26436);
xor U27290 (N_27290,N_26952,N_26342);
nor U27291 (N_27291,N_26820,N_26013);
or U27292 (N_27292,N_26363,N_26456);
xor U27293 (N_27293,N_26954,N_26231);
and U27294 (N_27294,N_26946,N_26264);
nand U27295 (N_27295,N_26839,N_26592);
xnor U27296 (N_27296,N_26924,N_26178);
nand U27297 (N_27297,N_26642,N_26204);
xor U27298 (N_27298,N_26248,N_26093);
xnor U27299 (N_27299,N_26255,N_26706);
nand U27300 (N_27300,N_26290,N_26914);
or U27301 (N_27301,N_26254,N_26055);
nor U27302 (N_27302,N_26744,N_26609);
xor U27303 (N_27303,N_26507,N_26002);
nand U27304 (N_27304,N_26973,N_26750);
or U27305 (N_27305,N_26335,N_26443);
nor U27306 (N_27306,N_26469,N_26057);
nor U27307 (N_27307,N_26268,N_26009);
and U27308 (N_27308,N_26185,N_26637);
or U27309 (N_27309,N_26593,N_26663);
nand U27310 (N_27310,N_26313,N_26969);
or U27311 (N_27311,N_26276,N_26649);
nor U27312 (N_27312,N_26001,N_26344);
or U27313 (N_27313,N_26347,N_26179);
or U27314 (N_27314,N_26739,N_26843);
and U27315 (N_27315,N_26181,N_26624);
nand U27316 (N_27316,N_26348,N_26664);
nand U27317 (N_27317,N_26687,N_26256);
and U27318 (N_27318,N_26811,N_26951);
or U27319 (N_27319,N_26107,N_26512);
and U27320 (N_27320,N_26167,N_26580);
nand U27321 (N_27321,N_26976,N_26056);
xnor U27322 (N_27322,N_26291,N_26476);
xor U27323 (N_27323,N_26381,N_26431);
nand U27324 (N_27324,N_26929,N_26237);
nand U27325 (N_27325,N_26077,N_26977);
nand U27326 (N_27326,N_26950,N_26694);
nand U27327 (N_27327,N_26817,N_26058);
or U27328 (N_27328,N_26863,N_26898);
or U27329 (N_27329,N_26695,N_26986);
or U27330 (N_27330,N_26066,N_26265);
and U27331 (N_27331,N_26112,N_26710);
or U27332 (N_27332,N_26948,N_26379);
and U27333 (N_27333,N_26524,N_26407);
nor U27334 (N_27334,N_26203,N_26155);
nand U27335 (N_27335,N_26091,N_26599);
and U27336 (N_27336,N_26240,N_26319);
nand U27337 (N_27337,N_26365,N_26070);
xnor U27338 (N_27338,N_26957,N_26743);
xor U27339 (N_27339,N_26293,N_26284);
nor U27340 (N_27340,N_26215,N_26489);
xnor U27341 (N_27341,N_26270,N_26341);
or U27342 (N_27342,N_26395,N_26535);
and U27343 (N_27343,N_26014,N_26894);
nor U27344 (N_27344,N_26189,N_26732);
nand U27345 (N_27345,N_26020,N_26918);
or U27346 (N_27346,N_26913,N_26677);
nor U27347 (N_27347,N_26823,N_26122);
nand U27348 (N_27348,N_26300,N_26873);
nor U27349 (N_27349,N_26500,N_26094);
nand U27350 (N_27350,N_26625,N_26229);
nand U27351 (N_27351,N_26372,N_26338);
xnor U27352 (N_27352,N_26978,N_26567);
nor U27353 (N_27353,N_26000,N_26471);
or U27354 (N_27354,N_26005,N_26763);
nor U27355 (N_27355,N_26947,N_26792);
nor U27356 (N_27356,N_26042,N_26243);
xnor U27357 (N_27357,N_26283,N_26140);
or U27358 (N_27358,N_26893,N_26985);
nand U27359 (N_27359,N_26766,N_26052);
and U27360 (N_27360,N_26404,N_26752);
nand U27361 (N_27361,N_26751,N_26654);
or U27362 (N_27362,N_26584,N_26205);
xor U27363 (N_27363,N_26640,N_26565);
nor U27364 (N_27364,N_26519,N_26115);
or U27365 (N_27365,N_26783,N_26852);
nor U27366 (N_27366,N_26723,N_26532);
nor U27367 (N_27367,N_26808,N_26865);
and U27368 (N_27368,N_26074,N_26257);
nor U27369 (N_27369,N_26369,N_26092);
xnor U27370 (N_27370,N_26147,N_26616);
and U27371 (N_27371,N_26132,N_26761);
and U27372 (N_27372,N_26420,N_26681);
nand U27373 (N_27373,N_26435,N_26780);
and U27374 (N_27374,N_26160,N_26510);
xor U27375 (N_27375,N_26628,N_26906);
and U27376 (N_27376,N_26069,N_26886);
or U27377 (N_27377,N_26027,N_26622);
nor U27378 (N_27378,N_26772,N_26795);
or U27379 (N_27379,N_26246,N_26159);
and U27380 (N_27380,N_26966,N_26832);
xor U27381 (N_27381,N_26463,N_26192);
nor U27382 (N_27382,N_26067,N_26004);
nand U27383 (N_27383,N_26019,N_26841);
nand U27384 (N_27384,N_26392,N_26223);
nand U27385 (N_27385,N_26922,N_26540);
nor U27386 (N_27386,N_26881,N_26771);
or U27387 (N_27387,N_26838,N_26963);
and U27388 (N_27388,N_26553,N_26965);
and U27389 (N_27389,N_26146,N_26439);
or U27390 (N_27390,N_26025,N_26199);
xnor U27391 (N_27391,N_26634,N_26251);
and U27392 (N_27392,N_26582,N_26473);
xor U27393 (N_27393,N_26998,N_26177);
or U27394 (N_27394,N_26989,N_26096);
or U27395 (N_27395,N_26354,N_26310);
and U27396 (N_27396,N_26968,N_26959);
xnor U27397 (N_27397,N_26170,N_26868);
nand U27398 (N_27398,N_26298,N_26498);
xnor U27399 (N_27399,N_26657,N_26645);
or U27400 (N_27400,N_26163,N_26194);
and U27401 (N_27401,N_26490,N_26828);
or U27402 (N_27402,N_26478,N_26935);
or U27403 (N_27403,N_26387,N_26888);
nor U27404 (N_27404,N_26474,N_26315);
nand U27405 (N_27405,N_26405,N_26173);
and U27406 (N_27406,N_26017,N_26555);
or U27407 (N_27407,N_26465,N_26883);
xnor U27408 (N_27408,N_26039,N_26225);
or U27409 (N_27409,N_26429,N_26169);
xnor U27410 (N_27410,N_26503,N_26632);
and U27411 (N_27411,N_26650,N_26595);
and U27412 (N_27412,N_26380,N_26988);
xnor U27413 (N_27413,N_26574,N_26029);
or U27414 (N_27414,N_26864,N_26477);
and U27415 (N_27415,N_26353,N_26605);
or U27416 (N_27416,N_26433,N_26855);
xnor U27417 (N_27417,N_26905,N_26955);
nand U27418 (N_27418,N_26089,N_26537);
and U27419 (N_27419,N_26333,N_26748);
nor U27420 (N_27420,N_26564,N_26814);
nand U27421 (N_27421,N_26872,N_26668);
and U27422 (N_27422,N_26450,N_26822);
and U27423 (N_27423,N_26171,N_26721);
nor U27424 (N_27424,N_26999,N_26983);
nand U27425 (N_27425,N_26462,N_26309);
or U27426 (N_27426,N_26200,N_26485);
or U27427 (N_27427,N_26050,N_26010);
xnor U27428 (N_27428,N_26653,N_26358);
xnor U27429 (N_27429,N_26081,N_26073);
nor U27430 (N_27430,N_26475,N_26550);
nor U27431 (N_27431,N_26245,N_26514);
or U27432 (N_27432,N_26030,N_26201);
or U27433 (N_27433,N_26389,N_26606);
xor U27434 (N_27434,N_26371,N_26007);
xnor U27435 (N_27435,N_26859,N_26305);
nor U27436 (N_27436,N_26041,N_26393);
and U27437 (N_27437,N_26612,N_26136);
or U27438 (N_27438,N_26289,N_26560);
or U27439 (N_27439,N_26269,N_26125);
xor U27440 (N_27440,N_26202,N_26699);
or U27441 (N_27441,N_26646,N_26346);
nand U27442 (N_27442,N_26383,N_26331);
nand U27443 (N_27443,N_26357,N_26878);
and U27444 (N_27444,N_26362,N_26933);
xor U27445 (N_27445,N_26997,N_26350);
nor U27446 (N_27446,N_26563,N_26406);
nand U27447 (N_27447,N_26212,N_26480);
nor U27448 (N_27448,N_26760,N_26418);
xnor U27449 (N_27449,N_26691,N_26206);
or U27450 (N_27450,N_26432,N_26043);
xnor U27451 (N_27451,N_26685,N_26789);
xnor U27452 (N_27452,N_26882,N_26736);
nor U27453 (N_27453,N_26127,N_26733);
and U27454 (N_27454,N_26765,N_26596);
nor U27455 (N_27455,N_26975,N_26629);
nor U27456 (N_27456,N_26656,N_26100);
nand U27457 (N_27457,N_26028,N_26876);
nor U27458 (N_27458,N_26633,N_26980);
nor U27459 (N_27459,N_26139,N_26271);
xor U27460 (N_27460,N_26821,N_26142);
nand U27461 (N_27461,N_26303,N_26917);
or U27462 (N_27462,N_26587,N_26460);
xor U27463 (N_27463,N_26619,N_26210);
and U27464 (N_27464,N_26697,N_26995);
nand U27465 (N_27465,N_26482,N_26408);
xnor U27466 (N_27466,N_26994,N_26120);
and U27467 (N_27467,N_26097,N_26304);
nor U27468 (N_27468,N_26164,N_26241);
or U27469 (N_27469,N_26892,N_26597);
xor U27470 (N_27470,N_26006,N_26613);
nand U27471 (N_27471,N_26327,N_26686);
nor U27472 (N_27472,N_26554,N_26552);
nor U27473 (N_27473,N_26377,N_26207);
xnor U27474 (N_27474,N_26704,N_26158);
nor U27475 (N_27475,N_26113,N_26228);
and U27476 (N_27476,N_26662,N_26696);
xnor U27477 (N_27477,N_26053,N_26242);
nand U27478 (N_27478,N_26531,N_26038);
and U27479 (N_27479,N_26594,N_26585);
or U27480 (N_27480,N_26102,N_26106);
and U27481 (N_27481,N_26581,N_26809);
or U27482 (N_27482,N_26591,N_26468);
and U27483 (N_27483,N_26259,N_26318);
and U27484 (N_27484,N_26423,N_26123);
nand U27485 (N_27485,N_26484,N_26015);
nor U27486 (N_27486,N_26931,N_26775);
or U27487 (N_27487,N_26501,N_26964);
xor U27488 (N_27488,N_26361,N_26541);
nand U27489 (N_27489,N_26570,N_26368);
or U27490 (N_27490,N_26314,N_26764);
nor U27491 (N_27491,N_26627,N_26128);
nand U27492 (N_27492,N_26958,N_26378);
nand U27493 (N_27493,N_26904,N_26154);
nand U27494 (N_27494,N_26401,N_26060);
and U27495 (N_27495,N_26528,N_26417);
or U27496 (N_27496,N_26109,N_26018);
nand U27497 (N_27497,N_26702,N_26572);
xnor U27498 (N_27498,N_26651,N_26198);
and U27499 (N_27499,N_26440,N_26842);
xnor U27500 (N_27500,N_26027,N_26801);
nand U27501 (N_27501,N_26891,N_26621);
and U27502 (N_27502,N_26099,N_26105);
nand U27503 (N_27503,N_26513,N_26086);
and U27504 (N_27504,N_26061,N_26068);
xnor U27505 (N_27505,N_26114,N_26345);
xor U27506 (N_27506,N_26731,N_26326);
or U27507 (N_27507,N_26941,N_26777);
or U27508 (N_27508,N_26836,N_26046);
and U27509 (N_27509,N_26656,N_26454);
nor U27510 (N_27510,N_26126,N_26438);
xnor U27511 (N_27511,N_26684,N_26362);
nand U27512 (N_27512,N_26912,N_26477);
nor U27513 (N_27513,N_26151,N_26080);
nor U27514 (N_27514,N_26782,N_26024);
and U27515 (N_27515,N_26179,N_26319);
nand U27516 (N_27516,N_26196,N_26892);
xor U27517 (N_27517,N_26465,N_26133);
nor U27518 (N_27518,N_26350,N_26951);
or U27519 (N_27519,N_26473,N_26642);
nor U27520 (N_27520,N_26268,N_26956);
and U27521 (N_27521,N_26444,N_26153);
xor U27522 (N_27522,N_26969,N_26248);
nor U27523 (N_27523,N_26477,N_26960);
nor U27524 (N_27524,N_26868,N_26096);
and U27525 (N_27525,N_26401,N_26892);
nor U27526 (N_27526,N_26516,N_26428);
nor U27527 (N_27527,N_26325,N_26260);
xnor U27528 (N_27528,N_26184,N_26832);
and U27529 (N_27529,N_26206,N_26756);
xor U27530 (N_27530,N_26475,N_26835);
nor U27531 (N_27531,N_26272,N_26456);
and U27532 (N_27532,N_26921,N_26559);
and U27533 (N_27533,N_26015,N_26721);
or U27534 (N_27534,N_26884,N_26974);
nand U27535 (N_27535,N_26965,N_26504);
or U27536 (N_27536,N_26544,N_26864);
nor U27537 (N_27537,N_26828,N_26189);
xnor U27538 (N_27538,N_26528,N_26291);
nor U27539 (N_27539,N_26488,N_26744);
xnor U27540 (N_27540,N_26076,N_26428);
nor U27541 (N_27541,N_26445,N_26734);
nor U27542 (N_27542,N_26447,N_26276);
nor U27543 (N_27543,N_26836,N_26344);
and U27544 (N_27544,N_26054,N_26883);
and U27545 (N_27545,N_26785,N_26397);
nor U27546 (N_27546,N_26587,N_26615);
nor U27547 (N_27547,N_26187,N_26666);
and U27548 (N_27548,N_26750,N_26305);
and U27549 (N_27549,N_26657,N_26721);
nor U27550 (N_27550,N_26081,N_26823);
nand U27551 (N_27551,N_26620,N_26325);
nand U27552 (N_27552,N_26120,N_26658);
xnor U27553 (N_27553,N_26840,N_26747);
nand U27554 (N_27554,N_26869,N_26213);
xnor U27555 (N_27555,N_26122,N_26294);
and U27556 (N_27556,N_26438,N_26198);
nor U27557 (N_27557,N_26761,N_26976);
or U27558 (N_27558,N_26718,N_26260);
nand U27559 (N_27559,N_26308,N_26555);
and U27560 (N_27560,N_26641,N_26215);
or U27561 (N_27561,N_26952,N_26949);
and U27562 (N_27562,N_26119,N_26319);
or U27563 (N_27563,N_26278,N_26866);
and U27564 (N_27564,N_26174,N_26293);
and U27565 (N_27565,N_26176,N_26322);
and U27566 (N_27566,N_26981,N_26776);
and U27567 (N_27567,N_26399,N_26100);
or U27568 (N_27568,N_26343,N_26910);
nor U27569 (N_27569,N_26205,N_26932);
xnor U27570 (N_27570,N_26151,N_26673);
xor U27571 (N_27571,N_26615,N_26307);
xnor U27572 (N_27572,N_26506,N_26336);
xnor U27573 (N_27573,N_26052,N_26583);
or U27574 (N_27574,N_26080,N_26563);
xnor U27575 (N_27575,N_26443,N_26091);
xor U27576 (N_27576,N_26785,N_26839);
and U27577 (N_27577,N_26428,N_26705);
nor U27578 (N_27578,N_26048,N_26361);
or U27579 (N_27579,N_26747,N_26777);
nor U27580 (N_27580,N_26133,N_26134);
or U27581 (N_27581,N_26921,N_26302);
or U27582 (N_27582,N_26678,N_26422);
nand U27583 (N_27583,N_26133,N_26532);
nor U27584 (N_27584,N_26834,N_26545);
xor U27585 (N_27585,N_26545,N_26739);
xor U27586 (N_27586,N_26536,N_26369);
nand U27587 (N_27587,N_26316,N_26883);
or U27588 (N_27588,N_26894,N_26118);
xnor U27589 (N_27589,N_26429,N_26625);
nand U27590 (N_27590,N_26636,N_26702);
nand U27591 (N_27591,N_26606,N_26328);
and U27592 (N_27592,N_26889,N_26640);
nand U27593 (N_27593,N_26932,N_26040);
nor U27594 (N_27594,N_26760,N_26464);
nand U27595 (N_27595,N_26468,N_26832);
or U27596 (N_27596,N_26257,N_26346);
and U27597 (N_27597,N_26941,N_26799);
or U27598 (N_27598,N_26268,N_26208);
xor U27599 (N_27599,N_26699,N_26305);
nand U27600 (N_27600,N_26518,N_26383);
or U27601 (N_27601,N_26860,N_26240);
and U27602 (N_27602,N_26684,N_26511);
xor U27603 (N_27603,N_26098,N_26751);
and U27604 (N_27604,N_26801,N_26432);
or U27605 (N_27605,N_26592,N_26352);
nand U27606 (N_27606,N_26578,N_26970);
nand U27607 (N_27607,N_26261,N_26673);
xnor U27608 (N_27608,N_26908,N_26110);
and U27609 (N_27609,N_26060,N_26191);
nor U27610 (N_27610,N_26927,N_26909);
xnor U27611 (N_27611,N_26668,N_26304);
and U27612 (N_27612,N_26316,N_26319);
nor U27613 (N_27613,N_26389,N_26051);
and U27614 (N_27614,N_26561,N_26050);
and U27615 (N_27615,N_26468,N_26529);
nand U27616 (N_27616,N_26259,N_26468);
xor U27617 (N_27617,N_26221,N_26461);
nand U27618 (N_27618,N_26418,N_26072);
and U27619 (N_27619,N_26559,N_26609);
xor U27620 (N_27620,N_26043,N_26472);
nor U27621 (N_27621,N_26842,N_26818);
nand U27622 (N_27622,N_26919,N_26809);
or U27623 (N_27623,N_26285,N_26616);
nor U27624 (N_27624,N_26077,N_26664);
or U27625 (N_27625,N_26031,N_26098);
xnor U27626 (N_27626,N_26168,N_26457);
nand U27627 (N_27627,N_26444,N_26389);
or U27628 (N_27628,N_26168,N_26122);
nor U27629 (N_27629,N_26412,N_26373);
or U27630 (N_27630,N_26573,N_26374);
and U27631 (N_27631,N_26691,N_26396);
nand U27632 (N_27632,N_26773,N_26945);
and U27633 (N_27633,N_26238,N_26636);
xnor U27634 (N_27634,N_26005,N_26093);
nor U27635 (N_27635,N_26109,N_26305);
nand U27636 (N_27636,N_26480,N_26405);
and U27637 (N_27637,N_26294,N_26171);
or U27638 (N_27638,N_26688,N_26914);
and U27639 (N_27639,N_26462,N_26709);
xor U27640 (N_27640,N_26764,N_26568);
nor U27641 (N_27641,N_26111,N_26096);
nor U27642 (N_27642,N_26466,N_26716);
nand U27643 (N_27643,N_26545,N_26338);
xor U27644 (N_27644,N_26591,N_26747);
or U27645 (N_27645,N_26483,N_26715);
nand U27646 (N_27646,N_26543,N_26917);
nor U27647 (N_27647,N_26580,N_26269);
or U27648 (N_27648,N_26704,N_26986);
nand U27649 (N_27649,N_26034,N_26332);
nand U27650 (N_27650,N_26334,N_26557);
nand U27651 (N_27651,N_26425,N_26916);
xnor U27652 (N_27652,N_26929,N_26290);
nand U27653 (N_27653,N_26007,N_26270);
or U27654 (N_27654,N_26142,N_26555);
nor U27655 (N_27655,N_26926,N_26295);
nor U27656 (N_27656,N_26987,N_26802);
or U27657 (N_27657,N_26606,N_26625);
xnor U27658 (N_27658,N_26908,N_26959);
and U27659 (N_27659,N_26776,N_26873);
xnor U27660 (N_27660,N_26436,N_26073);
and U27661 (N_27661,N_26760,N_26923);
or U27662 (N_27662,N_26640,N_26804);
nor U27663 (N_27663,N_26777,N_26543);
or U27664 (N_27664,N_26833,N_26066);
or U27665 (N_27665,N_26021,N_26088);
and U27666 (N_27666,N_26921,N_26936);
nor U27667 (N_27667,N_26703,N_26756);
and U27668 (N_27668,N_26951,N_26613);
nand U27669 (N_27669,N_26501,N_26215);
and U27670 (N_27670,N_26744,N_26822);
or U27671 (N_27671,N_26455,N_26254);
xor U27672 (N_27672,N_26325,N_26106);
nor U27673 (N_27673,N_26111,N_26836);
xnor U27674 (N_27674,N_26168,N_26146);
or U27675 (N_27675,N_26428,N_26054);
and U27676 (N_27676,N_26101,N_26665);
nor U27677 (N_27677,N_26790,N_26996);
or U27678 (N_27678,N_26281,N_26156);
nand U27679 (N_27679,N_26230,N_26574);
or U27680 (N_27680,N_26339,N_26751);
nand U27681 (N_27681,N_26828,N_26534);
and U27682 (N_27682,N_26658,N_26054);
nor U27683 (N_27683,N_26756,N_26205);
nor U27684 (N_27684,N_26529,N_26733);
nand U27685 (N_27685,N_26913,N_26776);
nor U27686 (N_27686,N_26389,N_26995);
xor U27687 (N_27687,N_26262,N_26780);
nor U27688 (N_27688,N_26943,N_26831);
or U27689 (N_27689,N_26465,N_26807);
nand U27690 (N_27690,N_26481,N_26657);
or U27691 (N_27691,N_26417,N_26803);
nand U27692 (N_27692,N_26207,N_26976);
nor U27693 (N_27693,N_26290,N_26835);
nor U27694 (N_27694,N_26040,N_26214);
xor U27695 (N_27695,N_26033,N_26498);
nor U27696 (N_27696,N_26693,N_26720);
xnor U27697 (N_27697,N_26277,N_26387);
or U27698 (N_27698,N_26814,N_26932);
and U27699 (N_27699,N_26544,N_26267);
and U27700 (N_27700,N_26226,N_26137);
xnor U27701 (N_27701,N_26802,N_26836);
and U27702 (N_27702,N_26804,N_26405);
xor U27703 (N_27703,N_26581,N_26973);
and U27704 (N_27704,N_26943,N_26644);
xnor U27705 (N_27705,N_26303,N_26650);
or U27706 (N_27706,N_26115,N_26764);
nor U27707 (N_27707,N_26200,N_26830);
nor U27708 (N_27708,N_26352,N_26170);
xor U27709 (N_27709,N_26946,N_26427);
nor U27710 (N_27710,N_26004,N_26462);
and U27711 (N_27711,N_26359,N_26205);
xor U27712 (N_27712,N_26862,N_26916);
or U27713 (N_27713,N_26155,N_26227);
or U27714 (N_27714,N_26039,N_26785);
xnor U27715 (N_27715,N_26510,N_26688);
xnor U27716 (N_27716,N_26283,N_26385);
or U27717 (N_27717,N_26672,N_26806);
nand U27718 (N_27718,N_26447,N_26167);
and U27719 (N_27719,N_26331,N_26895);
xnor U27720 (N_27720,N_26862,N_26511);
and U27721 (N_27721,N_26295,N_26860);
or U27722 (N_27722,N_26680,N_26775);
nor U27723 (N_27723,N_26630,N_26097);
or U27724 (N_27724,N_26548,N_26951);
nor U27725 (N_27725,N_26829,N_26195);
nand U27726 (N_27726,N_26415,N_26887);
and U27727 (N_27727,N_26151,N_26498);
nand U27728 (N_27728,N_26110,N_26448);
or U27729 (N_27729,N_26923,N_26114);
nand U27730 (N_27730,N_26117,N_26404);
xor U27731 (N_27731,N_26717,N_26852);
nor U27732 (N_27732,N_26268,N_26720);
or U27733 (N_27733,N_26395,N_26427);
and U27734 (N_27734,N_26181,N_26625);
nor U27735 (N_27735,N_26993,N_26902);
nor U27736 (N_27736,N_26572,N_26251);
and U27737 (N_27737,N_26922,N_26805);
nor U27738 (N_27738,N_26633,N_26409);
nand U27739 (N_27739,N_26485,N_26693);
nand U27740 (N_27740,N_26780,N_26840);
nor U27741 (N_27741,N_26095,N_26700);
xor U27742 (N_27742,N_26386,N_26432);
nand U27743 (N_27743,N_26780,N_26286);
xnor U27744 (N_27744,N_26054,N_26342);
and U27745 (N_27745,N_26840,N_26922);
xnor U27746 (N_27746,N_26682,N_26745);
or U27747 (N_27747,N_26847,N_26778);
and U27748 (N_27748,N_26996,N_26046);
nor U27749 (N_27749,N_26285,N_26489);
and U27750 (N_27750,N_26536,N_26734);
nor U27751 (N_27751,N_26349,N_26477);
and U27752 (N_27752,N_26897,N_26996);
nand U27753 (N_27753,N_26907,N_26357);
nor U27754 (N_27754,N_26576,N_26318);
and U27755 (N_27755,N_26059,N_26029);
nand U27756 (N_27756,N_26716,N_26441);
xor U27757 (N_27757,N_26913,N_26143);
nor U27758 (N_27758,N_26606,N_26654);
nand U27759 (N_27759,N_26809,N_26326);
nand U27760 (N_27760,N_26484,N_26512);
and U27761 (N_27761,N_26279,N_26344);
nor U27762 (N_27762,N_26847,N_26564);
xnor U27763 (N_27763,N_26811,N_26557);
nand U27764 (N_27764,N_26088,N_26873);
nand U27765 (N_27765,N_26594,N_26560);
nand U27766 (N_27766,N_26593,N_26408);
and U27767 (N_27767,N_26768,N_26266);
or U27768 (N_27768,N_26208,N_26467);
and U27769 (N_27769,N_26126,N_26018);
or U27770 (N_27770,N_26688,N_26669);
nand U27771 (N_27771,N_26131,N_26592);
or U27772 (N_27772,N_26427,N_26093);
nand U27773 (N_27773,N_26104,N_26145);
or U27774 (N_27774,N_26412,N_26680);
or U27775 (N_27775,N_26092,N_26599);
nor U27776 (N_27776,N_26622,N_26303);
or U27777 (N_27777,N_26628,N_26619);
nor U27778 (N_27778,N_26785,N_26530);
nand U27779 (N_27779,N_26430,N_26534);
nor U27780 (N_27780,N_26858,N_26520);
nor U27781 (N_27781,N_26658,N_26684);
and U27782 (N_27782,N_26488,N_26923);
nor U27783 (N_27783,N_26125,N_26590);
xor U27784 (N_27784,N_26774,N_26972);
nor U27785 (N_27785,N_26443,N_26472);
or U27786 (N_27786,N_26191,N_26253);
nand U27787 (N_27787,N_26330,N_26886);
nand U27788 (N_27788,N_26071,N_26286);
or U27789 (N_27789,N_26926,N_26708);
nor U27790 (N_27790,N_26390,N_26047);
nand U27791 (N_27791,N_26344,N_26921);
and U27792 (N_27792,N_26570,N_26739);
xor U27793 (N_27793,N_26514,N_26799);
xnor U27794 (N_27794,N_26010,N_26647);
and U27795 (N_27795,N_26021,N_26026);
or U27796 (N_27796,N_26403,N_26134);
and U27797 (N_27797,N_26180,N_26479);
nand U27798 (N_27798,N_26997,N_26151);
xnor U27799 (N_27799,N_26592,N_26400);
or U27800 (N_27800,N_26161,N_26617);
or U27801 (N_27801,N_26821,N_26736);
nand U27802 (N_27802,N_26319,N_26293);
xnor U27803 (N_27803,N_26530,N_26104);
nor U27804 (N_27804,N_26472,N_26384);
and U27805 (N_27805,N_26279,N_26894);
nor U27806 (N_27806,N_26237,N_26204);
xor U27807 (N_27807,N_26939,N_26705);
or U27808 (N_27808,N_26976,N_26544);
or U27809 (N_27809,N_26018,N_26048);
nand U27810 (N_27810,N_26536,N_26166);
nor U27811 (N_27811,N_26845,N_26141);
nor U27812 (N_27812,N_26052,N_26130);
or U27813 (N_27813,N_26109,N_26006);
or U27814 (N_27814,N_26624,N_26473);
or U27815 (N_27815,N_26943,N_26435);
and U27816 (N_27816,N_26646,N_26816);
nand U27817 (N_27817,N_26018,N_26419);
xnor U27818 (N_27818,N_26557,N_26780);
and U27819 (N_27819,N_26110,N_26351);
nand U27820 (N_27820,N_26965,N_26968);
nand U27821 (N_27821,N_26910,N_26421);
xor U27822 (N_27822,N_26218,N_26075);
nand U27823 (N_27823,N_26204,N_26180);
nor U27824 (N_27824,N_26288,N_26877);
nand U27825 (N_27825,N_26001,N_26736);
nand U27826 (N_27826,N_26654,N_26071);
nor U27827 (N_27827,N_26003,N_26383);
and U27828 (N_27828,N_26994,N_26043);
and U27829 (N_27829,N_26860,N_26422);
and U27830 (N_27830,N_26795,N_26943);
xor U27831 (N_27831,N_26334,N_26544);
or U27832 (N_27832,N_26632,N_26775);
nand U27833 (N_27833,N_26833,N_26291);
and U27834 (N_27834,N_26289,N_26116);
and U27835 (N_27835,N_26488,N_26646);
nand U27836 (N_27836,N_26044,N_26186);
nand U27837 (N_27837,N_26158,N_26272);
xnor U27838 (N_27838,N_26736,N_26680);
nand U27839 (N_27839,N_26168,N_26243);
or U27840 (N_27840,N_26840,N_26610);
nand U27841 (N_27841,N_26635,N_26380);
or U27842 (N_27842,N_26843,N_26058);
nand U27843 (N_27843,N_26026,N_26981);
and U27844 (N_27844,N_26962,N_26239);
or U27845 (N_27845,N_26361,N_26831);
xor U27846 (N_27846,N_26647,N_26054);
nand U27847 (N_27847,N_26320,N_26402);
or U27848 (N_27848,N_26181,N_26088);
xnor U27849 (N_27849,N_26005,N_26909);
nor U27850 (N_27850,N_26583,N_26741);
or U27851 (N_27851,N_26780,N_26475);
nand U27852 (N_27852,N_26714,N_26479);
xnor U27853 (N_27853,N_26297,N_26601);
nor U27854 (N_27854,N_26617,N_26411);
or U27855 (N_27855,N_26233,N_26134);
nand U27856 (N_27856,N_26672,N_26212);
nand U27857 (N_27857,N_26568,N_26496);
and U27858 (N_27858,N_26013,N_26145);
or U27859 (N_27859,N_26264,N_26758);
or U27860 (N_27860,N_26957,N_26145);
or U27861 (N_27861,N_26202,N_26372);
or U27862 (N_27862,N_26967,N_26041);
and U27863 (N_27863,N_26072,N_26100);
nand U27864 (N_27864,N_26876,N_26166);
and U27865 (N_27865,N_26839,N_26850);
xnor U27866 (N_27866,N_26334,N_26124);
nor U27867 (N_27867,N_26352,N_26165);
nand U27868 (N_27868,N_26272,N_26145);
nand U27869 (N_27869,N_26515,N_26031);
nand U27870 (N_27870,N_26375,N_26986);
nand U27871 (N_27871,N_26236,N_26186);
xnor U27872 (N_27872,N_26191,N_26694);
and U27873 (N_27873,N_26866,N_26586);
and U27874 (N_27874,N_26194,N_26804);
xor U27875 (N_27875,N_26960,N_26819);
xor U27876 (N_27876,N_26998,N_26599);
and U27877 (N_27877,N_26175,N_26163);
nand U27878 (N_27878,N_26186,N_26656);
nor U27879 (N_27879,N_26096,N_26474);
and U27880 (N_27880,N_26367,N_26702);
nor U27881 (N_27881,N_26193,N_26817);
or U27882 (N_27882,N_26336,N_26825);
and U27883 (N_27883,N_26997,N_26847);
xor U27884 (N_27884,N_26528,N_26855);
and U27885 (N_27885,N_26581,N_26610);
or U27886 (N_27886,N_26485,N_26964);
nand U27887 (N_27887,N_26429,N_26308);
xnor U27888 (N_27888,N_26425,N_26686);
xnor U27889 (N_27889,N_26934,N_26408);
or U27890 (N_27890,N_26654,N_26509);
nand U27891 (N_27891,N_26949,N_26882);
or U27892 (N_27892,N_26147,N_26447);
and U27893 (N_27893,N_26701,N_26900);
xnor U27894 (N_27894,N_26101,N_26439);
or U27895 (N_27895,N_26704,N_26685);
or U27896 (N_27896,N_26554,N_26524);
nor U27897 (N_27897,N_26646,N_26854);
nor U27898 (N_27898,N_26860,N_26276);
xnor U27899 (N_27899,N_26038,N_26609);
nor U27900 (N_27900,N_26285,N_26173);
nand U27901 (N_27901,N_26942,N_26126);
nand U27902 (N_27902,N_26508,N_26433);
nor U27903 (N_27903,N_26491,N_26446);
xor U27904 (N_27904,N_26521,N_26727);
nor U27905 (N_27905,N_26741,N_26027);
nand U27906 (N_27906,N_26837,N_26714);
or U27907 (N_27907,N_26869,N_26849);
and U27908 (N_27908,N_26072,N_26201);
and U27909 (N_27909,N_26450,N_26732);
nand U27910 (N_27910,N_26128,N_26579);
and U27911 (N_27911,N_26934,N_26123);
and U27912 (N_27912,N_26703,N_26731);
nand U27913 (N_27913,N_26534,N_26977);
nor U27914 (N_27914,N_26583,N_26306);
or U27915 (N_27915,N_26117,N_26218);
and U27916 (N_27916,N_26996,N_26952);
nor U27917 (N_27917,N_26703,N_26867);
or U27918 (N_27918,N_26863,N_26916);
nor U27919 (N_27919,N_26743,N_26523);
nand U27920 (N_27920,N_26043,N_26947);
or U27921 (N_27921,N_26765,N_26146);
xnor U27922 (N_27922,N_26840,N_26469);
xnor U27923 (N_27923,N_26252,N_26632);
or U27924 (N_27924,N_26623,N_26666);
xor U27925 (N_27925,N_26701,N_26213);
xor U27926 (N_27926,N_26392,N_26921);
nand U27927 (N_27927,N_26494,N_26435);
or U27928 (N_27928,N_26536,N_26419);
and U27929 (N_27929,N_26548,N_26048);
and U27930 (N_27930,N_26141,N_26258);
xnor U27931 (N_27931,N_26087,N_26260);
xor U27932 (N_27932,N_26618,N_26922);
nand U27933 (N_27933,N_26506,N_26069);
or U27934 (N_27934,N_26357,N_26375);
nand U27935 (N_27935,N_26470,N_26310);
nor U27936 (N_27936,N_26421,N_26822);
xnor U27937 (N_27937,N_26823,N_26020);
nand U27938 (N_27938,N_26319,N_26752);
nor U27939 (N_27939,N_26225,N_26859);
nand U27940 (N_27940,N_26965,N_26888);
xor U27941 (N_27941,N_26507,N_26966);
xor U27942 (N_27942,N_26563,N_26581);
xnor U27943 (N_27943,N_26201,N_26813);
and U27944 (N_27944,N_26170,N_26543);
nor U27945 (N_27945,N_26158,N_26727);
and U27946 (N_27946,N_26794,N_26098);
xnor U27947 (N_27947,N_26053,N_26137);
nand U27948 (N_27948,N_26212,N_26275);
nor U27949 (N_27949,N_26507,N_26175);
xnor U27950 (N_27950,N_26234,N_26380);
xnor U27951 (N_27951,N_26824,N_26036);
and U27952 (N_27952,N_26191,N_26669);
nand U27953 (N_27953,N_26669,N_26893);
xor U27954 (N_27954,N_26007,N_26436);
xnor U27955 (N_27955,N_26177,N_26334);
or U27956 (N_27956,N_26546,N_26847);
xnor U27957 (N_27957,N_26864,N_26068);
nand U27958 (N_27958,N_26960,N_26588);
nand U27959 (N_27959,N_26012,N_26573);
xnor U27960 (N_27960,N_26771,N_26009);
and U27961 (N_27961,N_26925,N_26461);
and U27962 (N_27962,N_26953,N_26140);
or U27963 (N_27963,N_26656,N_26677);
xor U27964 (N_27964,N_26499,N_26017);
xor U27965 (N_27965,N_26091,N_26491);
or U27966 (N_27966,N_26808,N_26298);
nand U27967 (N_27967,N_26310,N_26921);
and U27968 (N_27968,N_26971,N_26823);
and U27969 (N_27969,N_26000,N_26460);
or U27970 (N_27970,N_26095,N_26276);
xor U27971 (N_27971,N_26692,N_26394);
nor U27972 (N_27972,N_26723,N_26068);
nand U27973 (N_27973,N_26299,N_26442);
and U27974 (N_27974,N_26905,N_26244);
nand U27975 (N_27975,N_26713,N_26430);
nor U27976 (N_27976,N_26796,N_26555);
or U27977 (N_27977,N_26621,N_26115);
and U27978 (N_27978,N_26557,N_26256);
or U27979 (N_27979,N_26984,N_26318);
and U27980 (N_27980,N_26916,N_26387);
nor U27981 (N_27981,N_26428,N_26121);
and U27982 (N_27982,N_26351,N_26349);
nand U27983 (N_27983,N_26970,N_26131);
nand U27984 (N_27984,N_26155,N_26949);
and U27985 (N_27985,N_26709,N_26681);
nor U27986 (N_27986,N_26121,N_26578);
or U27987 (N_27987,N_26528,N_26699);
and U27988 (N_27988,N_26283,N_26603);
nor U27989 (N_27989,N_26548,N_26931);
and U27990 (N_27990,N_26699,N_26135);
nand U27991 (N_27991,N_26685,N_26697);
xor U27992 (N_27992,N_26143,N_26191);
nor U27993 (N_27993,N_26953,N_26018);
nor U27994 (N_27994,N_26646,N_26381);
or U27995 (N_27995,N_26001,N_26097);
and U27996 (N_27996,N_26873,N_26236);
nor U27997 (N_27997,N_26926,N_26662);
nand U27998 (N_27998,N_26473,N_26579);
or U27999 (N_27999,N_26444,N_26359);
xor U28000 (N_28000,N_27632,N_27831);
and U28001 (N_28001,N_27160,N_27413);
xor U28002 (N_28002,N_27166,N_27326);
xnor U28003 (N_28003,N_27492,N_27955);
nor U28004 (N_28004,N_27587,N_27571);
or U28005 (N_28005,N_27266,N_27081);
nor U28006 (N_28006,N_27287,N_27162);
nor U28007 (N_28007,N_27380,N_27531);
or U28008 (N_28008,N_27916,N_27150);
xnor U28009 (N_28009,N_27611,N_27251);
xnor U28010 (N_28010,N_27829,N_27414);
and U28011 (N_28011,N_27276,N_27067);
nor U28012 (N_28012,N_27727,N_27941);
or U28013 (N_28013,N_27917,N_27176);
nor U28014 (N_28014,N_27205,N_27719);
nor U28015 (N_28015,N_27455,N_27991);
nor U28016 (N_28016,N_27456,N_27695);
xor U28017 (N_28017,N_27522,N_27648);
and U28018 (N_28018,N_27878,N_27045);
and U28019 (N_28019,N_27093,N_27604);
or U28020 (N_28020,N_27370,N_27161);
nand U28021 (N_28021,N_27404,N_27507);
nand U28022 (N_28022,N_27841,N_27471);
nand U28023 (N_28023,N_27810,N_27749);
nor U28024 (N_28024,N_27072,N_27567);
or U28025 (N_28025,N_27011,N_27464);
nand U28026 (N_28026,N_27508,N_27994);
xnor U28027 (N_28027,N_27257,N_27446);
xor U28028 (N_28028,N_27865,N_27859);
nor U28029 (N_28029,N_27636,N_27718);
nand U28030 (N_28030,N_27599,N_27964);
or U28031 (N_28031,N_27324,N_27408);
nand U28032 (N_28032,N_27225,N_27772);
nand U28033 (N_28033,N_27348,N_27521);
nand U28034 (N_28034,N_27275,N_27237);
nor U28035 (N_28035,N_27042,N_27304);
or U28036 (N_28036,N_27364,N_27959);
nand U28037 (N_28037,N_27863,N_27181);
nand U28038 (N_28038,N_27242,N_27790);
nor U28039 (N_28039,N_27976,N_27137);
nand U28040 (N_28040,N_27342,N_27579);
or U28041 (N_28041,N_27131,N_27103);
nand U28042 (N_28042,N_27548,N_27821);
nand U28043 (N_28043,N_27180,N_27393);
xnor U28044 (N_28044,N_27639,N_27154);
or U28045 (N_28045,N_27842,N_27862);
or U28046 (N_28046,N_27539,N_27637);
or U28047 (N_28047,N_27889,N_27236);
nand U28048 (N_28048,N_27728,N_27776);
nand U28049 (N_28049,N_27215,N_27660);
xnor U28050 (N_28050,N_27759,N_27851);
xor U28051 (N_28051,N_27712,N_27801);
and U28052 (N_28052,N_27947,N_27778);
and U28053 (N_28053,N_27808,N_27077);
and U28054 (N_28054,N_27744,N_27904);
xnor U28055 (N_28055,N_27902,N_27460);
xor U28056 (N_28056,N_27788,N_27058);
xnor U28057 (N_28057,N_27490,N_27111);
nand U28058 (N_28058,N_27543,N_27930);
nand U28059 (N_28059,N_27331,N_27577);
nor U28060 (N_28060,N_27975,N_27729);
xor U28061 (N_28061,N_27377,N_27189);
nand U28062 (N_28062,N_27957,N_27797);
nand U28063 (N_28063,N_27389,N_27062);
nor U28064 (N_28064,N_27200,N_27277);
and U28065 (N_28065,N_27164,N_27444);
xor U28066 (N_28066,N_27676,N_27417);
nor U28067 (N_28067,N_27913,N_27855);
and U28068 (N_28068,N_27282,N_27666);
and U28069 (N_28069,N_27985,N_27982);
nand U28070 (N_28070,N_27918,N_27177);
xnor U28071 (N_28071,N_27149,N_27448);
nand U28072 (N_28072,N_27032,N_27584);
nand U28073 (N_28073,N_27600,N_27512);
and U28074 (N_28074,N_27929,N_27523);
nand U28075 (N_28075,N_27601,N_27306);
nand U28076 (N_28076,N_27899,N_27950);
nor U28077 (N_28077,N_27938,N_27562);
and U28078 (N_28078,N_27933,N_27877);
or U28079 (N_28079,N_27707,N_27777);
or U28080 (N_28080,N_27989,N_27514);
and U28081 (N_28081,N_27317,N_27720);
nor U28082 (N_28082,N_27027,N_27315);
nor U28083 (N_28083,N_27307,N_27977);
or U28084 (N_28084,N_27844,N_27942);
and U28085 (N_28085,N_27618,N_27968);
nor U28086 (N_28086,N_27170,N_27084);
and U28087 (N_28087,N_27468,N_27643);
xnor U28088 (N_28088,N_27121,N_27965);
xor U28089 (N_28089,N_27352,N_27954);
or U28090 (N_28090,N_27185,N_27421);
and U28091 (N_28091,N_27222,N_27376);
nand U28092 (N_28092,N_27211,N_27586);
nand U28093 (N_28093,N_27010,N_27650);
nor U28094 (N_28094,N_27798,N_27802);
or U28095 (N_28095,N_27167,N_27133);
nor U28096 (N_28096,N_27241,N_27921);
and U28097 (N_28097,N_27480,N_27756);
and U28098 (N_28098,N_27203,N_27207);
and U28099 (N_28099,N_27974,N_27429);
nor U28100 (N_28100,N_27519,N_27119);
xor U28101 (N_28101,N_27725,N_27513);
and U28102 (N_28102,N_27581,N_27983);
nor U28103 (N_28103,N_27425,N_27270);
nand U28104 (N_28104,N_27678,N_27803);
or U28105 (N_28105,N_27849,N_27388);
xor U28106 (N_28106,N_27229,N_27196);
nor U28107 (N_28107,N_27644,N_27765);
or U28108 (N_28108,N_27091,N_27190);
nand U28109 (N_28109,N_27269,N_27467);
nor U28110 (N_28110,N_27335,N_27589);
and U28111 (N_28111,N_27854,N_27520);
or U28112 (N_28112,N_27195,N_27732);
or U28113 (N_28113,N_27297,N_27073);
or U28114 (N_28114,N_27006,N_27069);
nor U28115 (N_28115,N_27793,N_27993);
or U28116 (N_28116,N_27527,N_27786);
or U28117 (N_28117,N_27961,N_27049);
nor U28118 (N_28118,N_27807,N_27485);
xor U28119 (N_28119,N_27595,N_27828);
xor U28120 (N_28120,N_27063,N_27186);
and U28121 (N_28121,N_27920,N_27140);
nand U28122 (N_28122,N_27670,N_27748);
xor U28123 (N_28123,N_27112,N_27281);
and U28124 (N_28124,N_27116,N_27845);
xnor U28125 (N_28125,N_27784,N_27505);
or U28126 (N_28126,N_27083,N_27375);
and U28127 (N_28127,N_27476,N_27419);
nand U28128 (N_28128,N_27592,N_27056);
nand U28129 (N_28129,N_27440,N_27191);
nand U28130 (N_28130,N_27672,N_27610);
or U28131 (N_28131,N_27293,N_27546);
and U28132 (N_28132,N_27373,N_27538);
nand U28133 (N_28133,N_27614,N_27343);
nor U28134 (N_28134,N_27198,N_27247);
and U28135 (N_28135,N_27840,N_27602);
nand U28136 (N_28136,N_27000,N_27396);
xor U28137 (N_28137,N_27858,N_27060);
nor U28138 (N_28138,N_27358,N_27780);
nand U28139 (N_28139,N_27911,N_27469);
and U28140 (N_28140,N_27213,N_27526);
xor U28141 (N_28141,N_27675,N_27145);
xnor U28142 (N_28142,N_27769,N_27381);
or U28143 (N_28143,N_27059,N_27474);
and U28144 (N_28144,N_27262,N_27924);
and U28145 (N_28145,N_27028,N_27700);
and U28146 (N_28146,N_27830,N_27135);
nor U28147 (N_28147,N_27972,N_27463);
or U28148 (N_28148,N_27124,N_27254);
or U28149 (N_28149,N_27591,N_27894);
nor U28150 (N_28150,N_27228,N_27015);
xnor U28151 (N_28151,N_27753,N_27770);
or U28152 (N_28152,N_27184,N_27263);
and U28153 (N_28153,N_27239,N_27635);
and U28154 (N_28154,N_27470,N_27547);
or U28155 (N_28155,N_27433,N_27187);
nand U28156 (N_28156,N_27664,N_27412);
or U28157 (N_28157,N_27407,N_27019);
or U28158 (N_28158,N_27880,N_27369);
and U28159 (N_28159,N_27716,N_27768);
xnor U28160 (N_28160,N_27745,N_27178);
or U28161 (N_28161,N_27402,N_27397);
xor U28162 (N_28162,N_27787,N_27026);
nand U28163 (N_28163,N_27937,N_27336);
xor U28164 (N_28164,N_27742,N_27202);
and U28165 (N_28165,N_27816,N_27979);
nor U28166 (N_28166,N_27504,N_27090);
nand U28167 (N_28167,N_27152,N_27428);
nand U28168 (N_28168,N_27450,N_27025);
xnor U28169 (N_28169,N_27697,N_27875);
and U28170 (N_28170,N_27836,N_27515);
xnor U28171 (N_28171,N_27677,N_27289);
or U28172 (N_28172,N_27936,N_27750);
nand U28173 (N_28173,N_27743,N_27147);
nor U28174 (N_28174,N_27308,N_27018);
or U28175 (N_28175,N_27426,N_27616);
and U28176 (N_28176,N_27169,N_27327);
nor U28177 (N_28177,N_27290,N_27949);
or U28178 (N_28178,N_27762,N_27051);
or U28179 (N_28179,N_27273,N_27879);
nor U28180 (N_28180,N_27477,N_27940);
xor U28181 (N_28181,N_27657,N_27052);
nor U28182 (N_28182,N_27895,N_27540);
and U28183 (N_28183,N_27640,N_27785);
or U28184 (N_28184,N_27303,N_27127);
nand U28185 (N_28185,N_27582,N_27245);
nor U28186 (N_28186,N_27710,N_27734);
nor U28187 (N_28187,N_27883,N_27510);
xnor U28188 (N_28188,N_27654,N_27298);
xnor U28189 (N_28189,N_27781,N_27261);
nor U28190 (N_28190,N_27679,N_27909);
nor U28191 (N_28191,N_27322,N_27128);
nand U28192 (N_28192,N_27900,N_27009);
or U28193 (N_28193,N_27486,N_27299);
xnor U28194 (N_28194,N_27035,N_27300);
and U28195 (N_28195,N_27148,N_27649);
xor U28196 (N_28196,N_27773,N_27366);
xnor U28197 (N_28197,N_27627,N_27212);
or U28198 (N_28198,N_27175,N_27182);
xnor U28199 (N_28199,N_27819,N_27096);
nand U28200 (N_28200,N_27055,N_27848);
nor U28201 (N_28201,N_27356,N_27100);
nand U28202 (N_28202,N_27061,N_27956);
nor U28203 (N_28203,N_27489,N_27488);
xor U28204 (N_28204,N_27250,N_27893);
or U28205 (N_28205,N_27665,N_27885);
or U28206 (N_28206,N_27039,N_27487);
or U28207 (N_28207,N_27570,N_27853);
nor U28208 (N_28208,N_27881,N_27509);
xor U28209 (N_28209,N_27107,N_27503);
xor U28210 (N_28210,N_27812,N_27832);
and U28211 (N_28211,N_27876,N_27701);
and U28212 (N_28212,N_27799,N_27106);
or U28213 (N_28213,N_27607,N_27496);
or U28214 (N_28214,N_27108,N_27458);
or U28215 (N_28215,N_27687,N_27925);
or U28216 (N_28216,N_27197,N_27260);
and U28217 (N_28217,N_27283,N_27048);
xor U28218 (N_28218,N_27690,N_27984);
nor U28219 (N_28219,N_27398,N_27651);
and U28220 (N_28220,N_27274,N_27033);
xnor U28221 (N_28221,N_27967,N_27951);
or U28222 (N_28222,N_27201,N_27642);
and U28223 (N_28223,N_27715,N_27453);
xor U28224 (N_28224,N_27806,N_27410);
and U28225 (N_28225,N_27384,N_27479);
nor U28226 (N_28226,N_27958,N_27826);
or U28227 (N_28227,N_27374,N_27530);
nor U28228 (N_28228,N_27981,N_27866);
nand U28229 (N_28229,N_27367,N_27932);
or U28230 (N_28230,N_27804,N_27795);
nand U28231 (N_28231,N_27430,N_27887);
or U28232 (N_28232,N_27462,N_27691);
nor U28233 (N_28233,N_27406,N_27811);
or U28234 (N_28234,N_27118,N_27020);
xnor U28235 (N_28235,N_27003,N_27126);
and U28236 (N_28236,N_27673,N_27559);
or U28237 (N_28237,N_27316,N_27647);
xnor U28238 (N_28238,N_27761,N_27763);
nand U28239 (N_28239,N_27054,N_27272);
xor U28240 (N_28240,N_27002,N_27192);
or U28241 (N_28241,N_27731,N_27330);
nor U28242 (N_28242,N_27927,N_27861);
nand U28243 (N_28243,N_27739,N_27117);
xor U28244 (N_28244,N_27130,N_27325);
nand U28245 (N_28245,N_27037,N_27846);
and U28246 (N_28246,N_27199,N_27357);
and U28247 (N_28247,N_27168,N_27905);
nand U28248 (N_28248,N_27053,N_27593);
xnor U28249 (N_28249,N_27231,N_27386);
nor U28250 (N_28250,N_27442,N_27767);
nor U28251 (N_28251,N_27655,N_27012);
xnor U28252 (N_28252,N_27724,N_27722);
and U28253 (N_28253,N_27232,N_27246);
xor U28254 (N_28254,N_27334,N_27087);
nor U28255 (N_28255,N_27301,N_27822);
and U28256 (N_28256,N_27646,N_27706);
xor U28257 (N_28257,N_27850,N_27963);
xnor U28258 (N_28258,N_27594,N_27741);
xor U28259 (N_28259,N_27572,N_27392);
or U28260 (N_28260,N_27014,N_27075);
and U28261 (N_28261,N_27556,N_27500);
xor U28262 (N_28262,N_27279,N_27590);
or U28263 (N_28263,N_27516,N_27353);
nand U28264 (N_28264,N_27578,N_27612);
and U28265 (N_28265,N_27007,N_27216);
nand U28266 (N_28266,N_27792,N_27259);
xnor U28267 (N_28267,N_27005,N_27016);
nor U28268 (N_28268,N_27023,N_27079);
and U28269 (N_28269,N_27074,N_27472);
and U28270 (N_28270,N_27436,N_27387);
and U28271 (N_28271,N_27104,N_27481);
xnor U28272 (N_28272,N_27783,N_27814);
or U28273 (N_28273,N_27194,N_27493);
and U28274 (N_28274,N_27333,N_27606);
nand U28275 (N_28275,N_27217,N_27692);
nand U28276 (N_28276,N_27340,N_27620);
xor U28277 (N_28277,N_27943,N_27319);
and U28278 (N_28278,N_27910,N_27337);
or U28279 (N_28279,N_27449,N_27835);
xor U28280 (N_28280,N_27574,N_27615);
nand U28281 (N_28281,N_27721,N_27362);
or U28282 (N_28282,N_27805,N_27013);
nand U28283 (N_28283,N_27702,N_27796);
nand U28284 (N_28284,N_27457,N_27043);
and U28285 (N_28285,N_27667,N_27758);
nor U28286 (N_28286,N_27057,N_27939);
nor U28287 (N_28287,N_27536,N_27372);
and U28288 (N_28288,N_27545,N_27995);
or U28289 (N_28289,N_27136,N_27782);
nand U28290 (N_28290,N_27794,N_27903);
nor U28291 (N_28291,N_27554,N_27529);
xnor U28292 (N_28292,N_27847,N_27423);
nand U28293 (N_28293,N_27537,N_27681);
nor U28294 (N_28294,N_27209,N_27354);
nand U28295 (N_28295,N_27435,N_27931);
xor U28296 (N_28296,N_27230,N_27638);
nor U28297 (N_28297,N_27224,N_27935);
and U28298 (N_28298,N_27142,N_27411);
xor U28299 (N_28299,N_27159,N_27709);
nor U28300 (N_28300,N_27608,N_27094);
nor U28301 (N_28301,N_27820,N_27065);
or U28302 (N_28302,N_27004,N_27800);
and U28303 (N_28303,N_27465,N_27248);
nand U28304 (N_28304,N_27233,N_27328);
nand U28305 (N_28305,N_27001,N_27506);
and U28306 (N_28306,N_27313,N_27815);
and U28307 (N_28307,N_27869,N_27349);
nand U28308 (N_28308,N_27310,N_27757);
or U28309 (N_28309,N_27332,N_27641);
xor U28310 (N_28310,N_27078,N_27155);
nor U28311 (N_28311,N_27365,N_27249);
and U28312 (N_28312,N_27491,N_27923);
or U28313 (N_28313,N_27305,N_27309);
xnor U28314 (N_28314,N_27441,N_27494);
nor U28315 (N_28315,N_27361,N_27834);
nor U28316 (N_28316,N_27320,N_27158);
and U28317 (N_28317,N_27422,N_27669);
nand U28318 (N_28318,N_27466,N_27824);
nor U28319 (N_28319,N_27041,N_27418);
xor U28320 (N_28320,N_27318,N_27971);
xor U28321 (N_28321,N_27478,N_27017);
and U28322 (N_28322,N_27717,N_27125);
nand U28323 (N_28323,N_27141,N_27906);
xor U28324 (N_28324,N_27383,N_27622);
xor U28325 (N_28325,N_27898,N_27652);
nor U28326 (N_28326,N_27143,N_27292);
nand U28327 (N_28327,N_27626,N_27870);
nor U28328 (N_28328,N_27220,N_27359);
nor U28329 (N_28329,N_27427,N_27511);
or U28330 (N_28330,N_27922,N_27431);
nor U28331 (N_28331,N_27825,N_27240);
or U28332 (N_28332,N_27085,N_27071);
xnor U28333 (N_28333,N_27437,N_27817);
xor U28334 (N_28334,N_27134,N_27944);
nor U28335 (N_28335,N_27597,N_27771);
nand U28336 (N_28336,N_27542,N_27401);
and U28337 (N_28337,N_27110,N_27311);
and U28338 (N_28338,N_27347,N_27703);
nand U28339 (N_28339,N_27746,N_27268);
or U28340 (N_28340,N_27945,N_27996);
nand U28341 (N_28341,N_27568,N_27897);
nor U28342 (N_28342,N_27482,N_27843);
and U28343 (N_28343,N_27583,N_27022);
nand U28344 (N_28344,N_27029,N_27760);
xnor U28345 (N_28345,N_27928,N_27399);
nor U28346 (N_28346,N_27223,N_27946);
xor U28347 (N_28347,N_27838,N_27775);
nor U28348 (N_28348,N_27686,N_27696);
xnor U28349 (N_28349,N_27129,N_27882);
xnor U28350 (N_28350,N_27288,N_27258);
xnor U28351 (N_28351,N_27573,N_27827);
or U28352 (N_28352,N_27339,N_27234);
nor U28353 (N_28353,N_27378,N_27535);
xnor U28354 (N_28354,N_27066,N_27541);
nand U28355 (N_28355,N_27653,N_27497);
and U28356 (N_28356,N_27285,N_27892);
nor U28357 (N_28357,N_27525,N_27857);
or U28358 (N_28358,N_27114,N_27867);
nor U28359 (N_28359,N_27912,N_27235);
nor U28360 (N_28360,N_27031,N_27238);
nand U28361 (N_28361,N_27082,N_27962);
or U28362 (N_28362,N_27046,N_27210);
nand U28363 (N_28363,N_27024,N_27395);
nor U28364 (N_28364,N_27736,N_27558);
and U28365 (N_28365,N_27550,N_27755);
and U28366 (N_28366,N_27064,N_27524);
or U28367 (N_28367,N_27873,N_27621);
nor U28368 (N_28368,N_27454,N_27532);
or U28369 (N_28369,N_27113,N_27534);
and U28370 (N_28370,N_27791,N_27628);
xor U28371 (N_28371,N_27747,N_27382);
nor U28372 (N_28372,N_27405,N_27634);
or U28373 (N_28373,N_27713,N_27751);
and U28374 (N_28374,N_27021,N_27998);
nand U28375 (N_28375,N_27969,N_27360);
or U28376 (N_28376,N_27907,N_27557);
and U28377 (N_28377,N_27163,N_27735);
and U28378 (N_28378,N_27551,N_27438);
or U28379 (N_28379,N_27092,N_27295);
nand U28380 (N_28380,N_27415,N_27999);
or U28381 (N_28381,N_27122,N_27475);
nor U28382 (N_28382,N_27645,N_27050);
nand U28383 (N_28383,N_27101,N_27265);
and U28384 (N_28384,N_27901,N_27864);
nor U28385 (N_28385,N_27227,N_27852);
nand U28386 (N_28386,N_27682,N_27099);
or U28387 (N_28387,N_27986,N_27139);
nor U28388 (N_28388,N_27656,N_27344);
nand U28389 (N_28389,N_27208,N_27764);
or U28390 (N_28390,N_27294,N_27754);
or U28391 (N_28391,N_27445,N_27416);
xnor U28392 (N_28392,N_27264,N_27284);
and U28393 (N_28393,N_27886,N_27598);
or U28394 (N_28394,N_27561,N_27605);
nor U28395 (N_28395,N_27323,N_27329);
and U28396 (N_28396,N_27693,N_27179);
nor U28397 (N_28397,N_27068,N_27278);
xnor U28398 (N_28398,N_27633,N_27156);
and U28399 (N_28399,N_27625,N_27576);
xnor U28400 (N_28400,N_27371,N_27047);
and U28401 (N_28401,N_27214,N_27566);
xor U28402 (N_28402,N_27174,N_27823);
nor U28403 (N_28403,N_27555,N_27560);
or U28404 (N_28404,N_27874,N_27439);
nand U28405 (N_28405,N_27960,N_27188);
or U28406 (N_28406,N_27390,N_27603);
nand U28407 (N_28407,N_27517,N_27694);
or U28408 (N_28408,N_27171,N_27280);
xnor U28409 (N_28409,N_27987,N_27711);
xor U28410 (N_28410,N_27157,N_27256);
nor U28411 (N_28411,N_27394,N_27990);
nor U28412 (N_28412,N_27350,N_27818);
nor U28413 (N_28413,N_27120,N_27351);
nand U28414 (N_28414,N_27473,N_27105);
nor U28415 (N_28415,N_27684,N_27890);
and U28416 (N_28416,N_27860,N_27363);
xor U28417 (N_28417,N_27988,N_27226);
and U28418 (N_28418,N_27737,N_27443);
and U28419 (N_28419,N_27345,N_27856);
and U28420 (N_28420,N_27766,N_27498);
or U28421 (N_28421,N_27206,N_27914);
nand U28422 (N_28422,N_27564,N_27165);
or U28423 (N_28423,N_27888,N_27617);
nand U28424 (N_28424,N_27321,N_27668);
or U28425 (N_28425,N_27837,N_27553);
or U28426 (N_28426,N_27080,N_27919);
and U28427 (N_28427,N_27252,N_27659);
xor U28428 (N_28428,N_27596,N_27338);
nor U28429 (N_28429,N_27738,N_27008);
or U28430 (N_28430,N_27451,N_27569);
nor U28431 (N_28431,N_27183,N_27495);
nand U28432 (N_28432,N_27624,N_27774);
xor U28433 (N_28433,N_27253,N_27671);
or U28434 (N_28434,N_27588,N_27502);
xnor U28435 (N_28435,N_27544,N_27044);
nand U28436 (N_28436,N_27219,N_27459);
and U28437 (N_28437,N_27575,N_27699);
xor U28438 (N_28438,N_27565,N_27296);
xor U28439 (N_28439,N_27086,N_27221);
nand U28440 (N_28440,N_27533,N_27409);
xnor U28441 (N_28441,N_27661,N_27115);
nand U28442 (N_28442,N_27173,N_27978);
and U28443 (N_28443,N_27952,N_27740);
xnor U28444 (N_28444,N_27076,N_27461);
xor U28445 (N_28445,N_27726,N_27244);
nand U28446 (N_28446,N_27549,N_27663);
or U28447 (N_28447,N_27123,N_27619);
and U28448 (N_28448,N_27030,N_27286);
or U28449 (N_28449,N_27193,N_27585);
nor U28450 (N_28450,N_27391,N_27089);
nor U28451 (N_28451,N_27915,N_27403);
nand U28452 (N_28452,N_27151,N_27243);
or U28453 (N_28453,N_27434,N_27698);
nor U28454 (N_28454,N_27779,N_27501);
nand U28455 (N_28455,N_27379,N_27872);
nor U28456 (N_28456,N_27662,N_27036);
nor U28457 (N_28457,N_27034,N_27683);
xor U28458 (N_28458,N_27789,N_27631);
and U28459 (N_28459,N_27097,N_27271);
and U28460 (N_28460,N_27095,N_27708);
nand U28461 (N_28461,N_27132,N_27973);
xnor U28462 (N_28462,N_27432,N_27884);
nand U28463 (N_28463,N_27813,N_27302);
xor U28464 (N_28464,N_27891,N_27680);
xor U28465 (N_28465,N_27146,N_27658);
nor U28466 (N_28466,N_27070,N_27934);
nor U28467 (N_28467,N_27752,N_27704);
xnor U28468 (N_28468,N_27970,N_27630);
xor U28469 (N_28469,N_27144,N_27953);
nand U28470 (N_28470,N_27314,N_27714);
nor U28471 (N_28471,N_27153,N_27580);
nor U28472 (N_28472,N_27267,N_27420);
or U28473 (N_28473,N_27552,N_27839);
and U28474 (N_28474,N_27674,N_27966);
nor U28475 (N_28475,N_27896,N_27871);
nor U28476 (N_28476,N_27355,N_27908);
and U28477 (N_28477,N_27484,N_27629);
nand U28478 (N_28478,N_27980,N_27038);
nor U28479 (N_28479,N_27613,N_27346);
xnor U28480 (N_28480,N_27623,N_27609);
or U28481 (N_28481,N_27688,N_27518);
or U28482 (N_28482,N_27992,N_27926);
nand U28483 (N_28483,N_27528,N_27723);
and U28484 (N_28484,N_27424,N_27689);
nor U28485 (N_28485,N_27368,N_27685);
nor U28486 (N_28486,N_27948,N_27138);
and U28487 (N_28487,N_27705,N_27102);
nand U28488 (N_28488,N_27809,N_27088);
and U28489 (N_28489,N_27563,N_27204);
nand U28490 (N_28490,N_27109,N_27499);
nor U28491 (N_28491,N_27730,N_27452);
nand U28492 (N_28492,N_27098,N_27172);
nor U28493 (N_28493,N_27447,N_27483);
nand U28494 (N_28494,N_27868,N_27385);
and U28495 (N_28495,N_27733,N_27291);
or U28496 (N_28496,N_27218,N_27997);
and U28497 (N_28497,N_27400,N_27341);
and U28498 (N_28498,N_27255,N_27312);
nand U28499 (N_28499,N_27040,N_27833);
or U28500 (N_28500,N_27509,N_27245);
and U28501 (N_28501,N_27955,N_27319);
xnor U28502 (N_28502,N_27212,N_27663);
nor U28503 (N_28503,N_27924,N_27085);
and U28504 (N_28504,N_27509,N_27694);
nor U28505 (N_28505,N_27814,N_27742);
xor U28506 (N_28506,N_27385,N_27744);
and U28507 (N_28507,N_27151,N_27029);
or U28508 (N_28508,N_27045,N_27896);
xor U28509 (N_28509,N_27495,N_27787);
and U28510 (N_28510,N_27485,N_27114);
or U28511 (N_28511,N_27424,N_27216);
nand U28512 (N_28512,N_27436,N_27792);
and U28513 (N_28513,N_27569,N_27227);
nor U28514 (N_28514,N_27544,N_27879);
xor U28515 (N_28515,N_27574,N_27090);
or U28516 (N_28516,N_27462,N_27209);
nor U28517 (N_28517,N_27409,N_27509);
and U28518 (N_28518,N_27604,N_27770);
nor U28519 (N_28519,N_27603,N_27322);
and U28520 (N_28520,N_27217,N_27424);
and U28521 (N_28521,N_27368,N_27588);
or U28522 (N_28522,N_27282,N_27386);
nor U28523 (N_28523,N_27263,N_27110);
nor U28524 (N_28524,N_27184,N_27245);
nand U28525 (N_28525,N_27121,N_27791);
nand U28526 (N_28526,N_27273,N_27915);
and U28527 (N_28527,N_27719,N_27717);
nand U28528 (N_28528,N_27636,N_27189);
xor U28529 (N_28529,N_27971,N_27109);
and U28530 (N_28530,N_27350,N_27403);
nor U28531 (N_28531,N_27035,N_27145);
and U28532 (N_28532,N_27615,N_27422);
or U28533 (N_28533,N_27185,N_27379);
nor U28534 (N_28534,N_27626,N_27988);
nor U28535 (N_28535,N_27101,N_27537);
and U28536 (N_28536,N_27976,N_27969);
and U28537 (N_28537,N_27339,N_27002);
or U28538 (N_28538,N_27931,N_27982);
and U28539 (N_28539,N_27141,N_27914);
xnor U28540 (N_28540,N_27615,N_27222);
nor U28541 (N_28541,N_27062,N_27775);
xor U28542 (N_28542,N_27726,N_27509);
and U28543 (N_28543,N_27097,N_27678);
or U28544 (N_28544,N_27294,N_27215);
and U28545 (N_28545,N_27260,N_27589);
or U28546 (N_28546,N_27507,N_27475);
nor U28547 (N_28547,N_27275,N_27231);
and U28548 (N_28548,N_27758,N_27121);
nor U28549 (N_28549,N_27301,N_27228);
xnor U28550 (N_28550,N_27920,N_27103);
nand U28551 (N_28551,N_27404,N_27333);
or U28552 (N_28552,N_27367,N_27907);
or U28553 (N_28553,N_27399,N_27809);
nor U28554 (N_28554,N_27872,N_27659);
nand U28555 (N_28555,N_27994,N_27839);
and U28556 (N_28556,N_27796,N_27581);
xnor U28557 (N_28557,N_27694,N_27002);
nor U28558 (N_28558,N_27617,N_27021);
nor U28559 (N_28559,N_27697,N_27773);
nand U28560 (N_28560,N_27117,N_27169);
xnor U28561 (N_28561,N_27249,N_27291);
or U28562 (N_28562,N_27760,N_27228);
nor U28563 (N_28563,N_27103,N_27983);
or U28564 (N_28564,N_27588,N_27761);
nand U28565 (N_28565,N_27315,N_27174);
or U28566 (N_28566,N_27269,N_27911);
and U28567 (N_28567,N_27409,N_27901);
or U28568 (N_28568,N_27740,N_27095);
and U28569 (N_28569,N_27318,N_27624);
nor U28570 (N_28570,N_27988,N_27536);
or U28571 (N_28571,N_27519,N_27934);
nor U28572 (N_28572,N_27758,N_27509);
xor U28573 (N_28573,N_27662,N_27997);
xor U28574 (N_28574,N_27808,N_27339);
nand U28575 (N_28575,N_27798,N_27269);
or U28576 (N_28576,N_27434,N_27292);
or U28577 (N_28577,N_27782,N_27152);
nand U28578 (N_28578,N_27617,N_27044);
nand U28579 (N_28579,N_27735,N_27243);
xor U28580 (N_28580,N_27802,N_27184);
nand U28581 (N_28581,N_27386,N_27321);
xor U28582 (N_28582,N_27400,N_27595);
xor U28583 (N_28583,N_27791,N_27574);
xnor U28584 (N_28584,N_27677,N_27302);
nand U28585 (N_28585,N_27222,N_27005);
or U28586 (N_28586,N_27327,N_27234);
and U28587 (N_28587,N_27058,N_27969);
nand U28588 (N_28588,N_27130,N_27818);
and U28589 (N_28589,N_27774,N_27943);
nor U28590 (N_28590,N_27620,N_27561);
nor U28591 (N_28591,N_27231,N_27037);
xor U28592 (N_28592,N_27936,N_27557);
or U28593 (N_28593,N_27494,N_27311);
nor U28594 (N_28594,N_27017,N_27364);
nand U28595 (N_28595,N_27484,N_27789);
nor U28596 (N_28596,N_27667,N_27613);
xnor U28597 (N_28597,N_27638,N_27291);
or U28598 (N_28598,N_27354,N_27457);
or U28599 (N_28599,N_27918,N_27619);
nor U28600 (N_28600,N_27381,N_27190);
nor U28601 (N_28601,N_27707,N_27812);
nor U28602 (N_28602,N_27322,N_27725);
nand U28603 (N_28603,N_27955,N_27642);
xnor U28604 (N_28604,N_27460,N_27360);
nand U28605 (N_28605,N_27241,N_27612);
nand U28606 (N_28606,N_27578,N_27203);
and U28607 (N_28607,N_27717,N_27971);
nor U28608 (N_28608,N_27476,N_27477);
nand U28609 (N_28609,N_27528,N_27736);
nor U28610 (N_28610,N_27025,N_27320);
and U28611 (N_28611,N_27340,N_27585);
or U28612 (N_28612,N_27754,N_27695);
xnor U28613 (N_28613,N_27083,N_27064);
and U28614 (N_28614,N_27591,N_27138);
nand U28615 (N_28615,N_27026,N_27904);
nor U28616 (N_28616,N_27499,N_27578);
xor U28617 (N_28617,N_27032,N_27418);
xnor U28618 (N_28618,N_27419,N_27274);
or U28619 (N_28619,N_27970,N_27781);
nand U28620 (N_28620,N_27938,N_27244);
nor U28621 (N_28621,N_27817,N_27324);
and U28622 (N_28622,N_27591,N_27606);
xnor U28623 (N_28623,N_27491,N_27953);
xor U28624 (N_28624,N_27586,N_27548);
nor U28625 (N_28625,N_27504,N_27640);
and U28626 (N_28626,N_27330,N_27177);
xor U28627 (N_28627,N_27710,N_27251);
nand U28628 (N_28628,N_27682,N_27718);
and U28629 (N_28629,N_27284,N_27926);
nand U28630 (N_28630,N_27471,N_27347);
or U28631 (N_28631,N_27689,N_27041);
and U28632 (N_28632,N_27811,N_27927);
nor U28633 (N_28633,N_27492,N_27091);
or U28634 (N_28634,N_27570,N_27086);
nor U28635 (N_28635,N_27655,N_27267);
nor U28636 (N_28636,N_27639,N_27614);
and U28637 (N_28637,N_27967,N_27446);
xnor U28638 (N_28638,N_27258,N_27380);
or U28639 (N_28639,N_27713,N_27507);
xor U28640 (N_28640,N_27804,N_27214);
nand U28641 (N_28641,N_27385,N_27457);
or U28642 (N_28642,N_27539,N_27331);
nor U28643 (N_28643,N_27578,N_27857);
nand U28644 (N_28644,N_27263,N_27064);
nand U28645 (N_28645,N_27715,N_27677);
or U28646 (N_28646,N_27907,N_27683);
xnor U28647 (N_28647,N_27808,N_27723);
xor U28648 (N_28648,N_27231,N_27235);
or U28649 (N_28649,N_27116,N_27604);
nand U28650 (N_28650,N_27844,N_27397);
nand U28651 (N_28651,N_27460,N_27013);
nor U28652 (N_28652,N_27483,N_27479);
xnor U28653 (N_28653,N_27802,N_27253);
nand U28654 (N_28654,N_27955,N_27227);
or U28655 (N_28655,N_27422,N_27969);
nand U28656 (N_28656,N_27221,N_27686);
nor U28657 (N_28657,N_27138,N_27091);
xor U28658 (N_28658,N_27910,N_27503);
xnor U28659 (N_28659,N_27576,N_27628);
xnor U28660 (N_28660,N_27026,N_27101);
nor U28661 (N_28661,N_27368,N_27192);
and U28662 (N_28662,N_27857,N_27029);
nor U28663 (N_28663,N_27654,N_27690);
xor U28664 (N_28664,N_27289,N_27058);
nor U28665 (N_28665,N_27108,N_27834);
or U28666 (N_28666,N_27486,N_27062);
nor U28667 (N_28667,N_27349,N_27227);
xnor U28668 (N_28668,N_27436,N_27279);
xnor U28669 (N_28669,N_27914,N_27757);
and U28670 (N_28670,N_27896,N_27695);
or U28671 (N_28671,N_27265,N_27018);
nor U28672 (N_28672,N_27646,N_27943);
xor U28673 (N_28673,N_27933,N_27776);
xnor U28674 (N_28674,N_27641,N_27064);
nor U28675 (N_28675,N_27721,N_27799);
nor U28676 (N_28676,N_27193,N_27783);
nor U28677 (N_28677,N_27871,N_27732);
xor U28678 (N_28678,N_27064,N_27037);
or U28679 (N_28679,N_27545,N_27323);
and U28680 (N_28680,N_27592,N_27436);
or U28681 (N_28681,N_27750,N_27013);
xnor U28682 (N_28682,N_27593,N_27257);
and U28683 (N_28683,N_27419,N_27248);
nor U28684 (N_28684,N_27902,N_27883);
xnor U28685 (N_28685,N_27881,N_27971);
nor U28686 (N_28686,N_27965,N_27946);
xor U28687 (N_28687,N_27029,N_27929);
or U28688 (N_28688,N_27888,N_27909);
nand U28689 (N_28689,N_27134,N_27623);
nor U28690 (N_28690,N_27331,N_27013);
or U28691 (N_28691,N_27731,N_27244);
xor U28692 (N_28692,N_27227,N_27739);
nor U28693 (N_28693,N_27673,N_27560);
and U28694 (N_28694,N_27504,N_27630);
nand U28695 (N_28695,N_27502,N_27824);
or U28696 (N_28696,N_27915,N_27866);
and U28697 (N_28697,N_27407,N_27168);
and U28698 (N_28698,N_27510,N_27930);
and U28699 (N_28699,N_27522,N_27749);
xor U28700 (N_28700,N_27063,N_27577);
nand U28701 (N_28701,N_27727,N_27764);
or U28702 (N_28702,N_27291,N_27059);
xnor U28703 (N_28703,N_27780,N_27401);
nand U28704 (N_28704,N_27439,N_27099);
and U28705 (N_28705,N_27450,N_27633);
or U28706 (N_28706,N_27557,N_27381);
xnor U28707 (N_28707,N_27408,N_27522);
nor U28708 (N_28708,N_27354,N_27778);
nand U28709 (N_28709,N_27840,N_27779);
nor U28710 (N_28710,N_27171,N_27955);
nand U28711 (N_28711,N_27078,N_27558);
or U28712 (N_28712,N_27798,N_27176);
nand U28713 (N_28713,N_27292,N_27088);
nor U28714 (N_28714,N_27904,N_27110);
xor U28715 (N_28715,N_27214,N_27588);
or U28716 (N_28716,N_27580,N_27576);
nor U28717 (N_28717,N_27397,N_27137);
and U28718 (N_28718,N_27158,N_27187);
or U28719 (N_28719,N_27944,N_27530);
and U28720 (N_28720,N_27961,N_27809);
xor U28721 (N_28721,N_27534,N_27799);
and U28722 (N_28722,N_27132,N_27408);
nor U28723 (N_28723,N_27861,N_27122);
nand U28724 (N_28724,N_27971,N_27996);
nand U28725 (N_28725,N_27231,N_27887);
and U28726 (N_28726,N_27227,N_27245);
xor U28727 (N_28727,N_27326,N_27009);
or U28728 (N_28728,N_27303,N_27829);
nand U28729 (N_28729,N_27359,N_27974);
nand U28730 (N_28730,N_27717,N_27817);
and U28731 (N_28731,N_27056,N_27709);
or U28732 (N_28732,N_27287,N_27062);
xor U28733 (N_28733,N_27342,N_27059);
nor U28734 (N_28734,N_27133,N_27602);
nand U28735 (N_28735,N_27170,N_27858);
nor U28736 (N_28736,N_27141,N_27736);
or U28737 (N_28737,N_27975,N_27175);
xor U28738 (N_28738,N_27952,N_27407);
xor U28739 (N_28739,N_27093,N_27885);
and U28740 (N_28740,N_27935,N_27332);
or U28741 (N_28741,N_27442,N_27320);
and U28742 (N_28742,N_27710,N_27848);
xor U28743 (N_28743,N_27462,N_27153);
nand U28744 (N_28744,N_27809,N_27674);
and U28745 (N_28745,N_27246,N_27077);
xnor U28746 (N_28746,N_27794,N_27575);
nor U28747 (N_28747,N_27247,N_27538);
xor U28748 (N_28748,N_27932,N_27693);
and U28749 (N_28749,N_27968,N_27625);
nor U28750 (N_28750,N_27390,N_27226);
nor U28751 (N_28751,N_27867,N_27041);
nor U28752 (N_28752,N_27319,N_27564);
nand U28753 (N_28753,N_27283,N_27300);
nand U28754 (N_28754,N_27684,N_27141);
or U28755 (N_28755,N_27390,N_27141);
nor U28756 (N_28756,N_27622,N_27962);
nor U28757 (N_28757,N_27475,N_27518);
nor U28758 (N_28758,N_27514,N_27091);
nor U28759 (N_28759,N_27187,N_27671);
nor U28760 (N_28760,N_27471,N_27009);
xor U28761 (N_28761,N_27314,N_27294);
and U28762 (N_28762,N_27860,N_27826);
or U28763 (N_28763,N_27490,N_27159);
and U28764 (N_28764,N_27924,N_27997);
and U28765 (N_28765,N_27199,N_27792);
or U28766 (N_28766,N_27703,N_27097);
nand U28767 (N_28767,N_27579,N_27319);
nand U28768 (N_28768,N_27451,N_27143);
xor U28769 (N_28769,N_27969,N_27751);
nand U28770 (N_28770,N_27753,N_27529);
or U28771 (N_28771,N_27089,N_27675);
or U28772 (N_28772,N_27375,N_27596);
xor U28773 (N_28773,N_27275,N_27795);
nand U28774 (N_28774,N_27706,N_27428);
xor U28775 (N_28775,N_27685,N_27364);
nand U28776 (N_28776,N_27677,N_27511);
nand U28777 (N_28777,N_27641,N_27730);
nor U28778 (N_28778,N_27499,N_27156);
nor U28779 (N_28779,N_27656,N_27242);
nor U28780 (N_28780,N_27309,N_27951);
xor U28781 (N_28781,N_27737,N_27947);
or U28782 (N_28782,N_27930,N_27345);
nor U28783 (N_28783,N_27908,N_27361);
and U28784 (N_28784,N_27562,N_27912);
nand U28785 (N_28785,N_27613,N_27049);
and U28786 (N_28786,N_27079,N_27270);
and U28787 (N_28787,N_27653,N_27724);
nor U28788 (N_28788,N_27831,N_27879);
nor U28789 (N_28789,N_27880,N_27045);
or U28790 (N_28790,N_27250,N_27341);
xor U28791 (N_28791,N_27241,N_27679);
and U28792 (N_28792,N_27270,N_27173);
xor U28793 (N_28793,N_27546,N_27562);
nor U28794 (N_28794,N_27190,N_27135);
and U28795 (N_28795,N_27488,N_27467);
and U28796 (N_28796,N_27389,N_27745);
and U28797 (N_28797,N_27383,N_27020);
and U28798 (N_28798,N_27135,N_27594);
and U28799 (N_28799,N_27603,N_27213);
nand U28800 (N_28800,N_27004,N_27494);
and U28801 (N_28801,N_27311,N_27348);
nor U28802 (N_28802,N_27400,N_27045);
or U28803 (N_28803,N_27700,N_27108);
xor U28804 (N_28804,N_27911,N_27196);
nand U28805 (N_28805,N_27866,N_27612);
and U28806 (N_28806,N_27979,N_27679);
and U28807 (N_28807,N_27842,N_27419);
and U28808 (N_28808,N_27157,N_27216);
xnor U28809 (N_28809,N_27441,N_27776);
and U28810 (N_28810,N_27611,N_27332);
xnor U28811 (N_28811,N_27193,N_27042);
or U28812 (N_28812,N_27336,N_27296);
or U28813 (N_28813,N_27530,N_27606);
and U28814 (N_28814,N_27831,N_27971);
nor U28815 (N_28815,N_27168,N_27990);
or U28816 (N_28816,N_27673,N_27891);
nand U28817 (N_28817,N_27379,N_27430);
and U28818 (N_28818,N_27942,N_27884);
nand U28819 (N_28819,N_27106,N_27617);
nor U28820 (N_28820,N_27692,N_27152);
or U28821 (N_28821,N_27756,N_27840);
xnor U28822 (N_28822,N_27952,N_27371);
or U28823 (N_28823,N_27859,N_27262);
or U28824 (N_28824,N_27143,N_27621);
nand U28825 (N_28825,N_27246,N_27414);
nor U28826 (N_28826,N_27559,N_27365);
or U28827 (N_28827,N_27011,N_27514);
and U28828 (N_28828,N_27509,N_27007);
and U28829 (N_28829,N_27200,N_27081);
xor U28830 (N_28830,N_27910,N_27954);
or U28831 (N_28831,N_27097,N_27923);
or U28832 (N_28832,N_27349,N_27640);
nand U28833 (N_28833,N_27703,N_27763);
nand U28834 (N_28834,N_27134,N_27520);
or U28835 (N_28835,N_27716,N_27335);
or U28836 (N_28836,N_27100,N_27575);
and U28837 (N_28837,N_27488,N_27125);
and U28838 (N_28838,N_27899,N_27651);
and U28839 (N_28839,N_27323,N_27941);
nor U28840 (N_28840,N_27263,N_27819);
and U28841 (N_28841,N_27563,N_27306);
or U28842 (N_28842,N_27399,N_27461);
nand U28843 (N_28843,N_27010,N_27448);
and U28844 (N_28844,N_27954,N_27044);
nand U28845 (N_28845,N_27370,N_27955);
or U28846 (N_28846,N_27010,N_27238);
or U28847 (N_28847,N_27055,N_27697);
nor U28848 (N_28848,N_27658,N_27443);
or U28849 (N_28849,N_27721,N_27965);
xor U28850 (N_28850,N_27488,N_27722);
xnor U28851 (N_28851,N_27448,N_27497);
xnor U28852 (N_28852,N_27270,N_27061);
nor U28853 (N_28853,N_27338,N_27825);
or U28854 (N_28854,N_27720,N_27854);
nor U28855 (N_28855,N_27055,N_27129);
nor U28856 (N_28856,N_27225,N_27031);
or U28857 (N_28857,N_27436,N_27750);
or U28858 (N_28858,N_27007,N_27663);
nor U28859 (N_28859,N_27132,N_27537);
nor U28860 (N_28860,N_27330,N_27860);
nand U28861 (N_28861,N_27536,N_27090);
nor U28862 (N_28862,N_27563,N_27915);
and U28863 (N_28863,N_27156,N_27760);
and U28864 (N_28864,N_27579,N_27308);
nor U28865 (N_28865,N_27848,N_27782);
or U28866 (N_28866,N_27943,N_27007);
nand U28867 (N_28867,N_27999,N_27309);
xnor U28868 (N_28868,N_27696,N_27382);
or U28869 (N_28869,N_27212,N_27263);
xor U28870 (N_28870,N_27801,N_27524);
or U28871 (N_28871,N_27581,N_27479);
nor U28872 (N_28872,N_27872,N_27440);
xor U28873 (N_28873,N_27748,N_27190);
xnor U28874 (N_28874,N_27524,N_27477);
or U28875 (N_28875,N_27905,N_27736);
or U28876 (N_28876,N_27039,N_27260);
xor U28877 (N_28877,N_27682,N_27298);
and U28878 (N_28878,N_27248,N_27483);
nor U28879 (N_28879,N_27556,N_27481);
and U28880 (N_28880,N_27300,N_27809);
nor U28881 (N_28881,N_27950,N_27578);
nand U28882 (N_28882,N_27539,N_27315);
or U28883 (N_28883,N_27613,N_27692);
or U28884 (N_28884,N_27572,N_27577);
nand U28885 (N_28885,N_27300,N_27213);
nor U28886 (N_28886,N_27545,N_27917);
or U28887 (N_28887,N_27735,N_27671);
xnor U28888 (N_28888,N_27095,N_27204);
nand U28889 (N_28889,N_27923,N_27990);
and U28890 (N_28890,N_27277,N_27811);
nand U28891 (N_28891,N_27748,N_27510);
nand U28892 (N_28892,N_27111,N_27164);
and U28893 (N_28893,N_27091,N_27119);
nand U28894 (N_28894,N_27555,N_27577);
or U28895 (N_28895,N_27918,N_27032);
nor U28896 (N_28896,N_27488,N_27170);
nor U28897 (N_28897,N_27584,N_27940);
and U28898 (N_28898,N_27564,N_27253);
or U28899 (N_28899,N_27557,N_27275);
nand U28900 (N_28900,N_27695,N_27863);
nor U28901 (N_28901,N_27870,N_27855);
nand U28902 (N_28902,N_27939,N_27872);
and U28903 (N_28903,N_27458,N_27440);
nor U28904 (N_28904,N_27491,N_27145);
and U28905 (N_28905,N_27399,N_27717);
nor U28906 (N_28906,N_27251,N_27931);
nor U28907 (N_28907,N_27597,N_27399);
or U28908 (N_28908,N_27419,N_27834);
nand U28909 (N_28909,N_27904,N_27215);
xnor U28910 (N_28910,N_27571,N_27364);
nand U28911 (N_28911,N_27775,N_27677);
nor U28912 (N_28912,N_27982,N_27979);
or U28913 (N_28913,N_27754,N_27245);
and U28914 (N_28914,N_27097,N_27949);
xor U28915 (N_28915,N_27564,N_27481);
and U28916 (N_28916,N_27685,N_27051);
xor U28917 (N_28917,N_27925,N_27816);
or U28918 (N_28918,N_27065,N_27180);
nor U28919 (N_28919,N_27756,N_27564);
xnor U28920 (N_28920,N_27459,N_27461);
nand U28921 (N_28921,N_27733,N_27937);
or U28922 (N_28922,N_27582,N_27845);
nor U28923 (N_28923,N_27738,N_27150);
xor U28924 (N_28924,N_27360,N_27455);
nor U28925 (N_28925,N_27215,N_27298);
nor U28926 (N_28926,N_27748,N_27437);
nand U28927 (N_28927,N_27656,N_27941);
and U28928 (N_28928,N_27487,N_27387);
and U28929 (N_28929,N_27059,N_27896);
nor U28930 (N_28930,N_27204,N_27177);
nor U28931 (N_28931,N_27418,N_27033);
xor U28932 (N_28932,N_27747,N_27255);
nor U28933 (N_28933,N_27630,N_27239);
or U28934 (N_28934,N_27900,N_27641);
xnor U28935 (N_28935,N_27693,N_27038);
or U28936 (N_28936,N_27692,N_27390);
and U28937 (N_28937,N_27776,N_27532);
xor U28938 (N_28938,N_27820,N_27774);
or U28939 (N_28939,N_27174,N_27572);
xor U28940 (N_28940,N_27820,N_27157);
nand U28941 (N_28941,N_27940,N_27089);
nor U28942 (N_28942,N_27494,N_27458);
nand U28943 (N_28943,N_27386,N_27484);
nor U28944 (N_28944,N_27141,N_27450);
xor U28945 (N_28945,N_27091,N_27701);
xnor U28946 (N_28946,N_27035,N_27262);
nor U28947 (N_28947,N_27305,N_27731);
nor U28948 (N_28948,N_27305,N_27199);
or U28949 (N_28949,N_27601,N_27021);
xnor U28950 (N_28950,N_27778,N_27116);
or U28951 (N_28951,N_27470,N_27111);
xor U28952 (N_28952,N_27225,N_27214);
nor U28953 (N_28953,N_27231,N_27599);
nand U28954 (N_28954,N_27103,N_27820);
or U28955 (N_28955,N_27649,N_27730);
nor U28956 (N_28956,N_27563,N_27205);
and U28957 (N_28957,N_27333,N_27749);
nor U28958 (N_28958,N_27061,N_27058);
nand U28959 (N_28959,N_27133,N_27766);
nor U28960 (N_28960,N_27093,N_27688);
nor U28961 (N_28961,N_27421,N_27473);
and U28962 (N_28962,N_27794,N_27594);
nor U28963 (N_28963,N_27461,N_27523);
xnor U28964 (N_28964,N_27199,N_27665);
nand U28965 (N_28965,N_27788,N_27387);
and U28966 (N_28966,N_27192,N_27522);
nand U28967 (N_28967,N_27052,N_27620);
nand U28968 (N_28968,N_27769,N_27931);
or U28969 (N_28969,N_27972,N_27851);
and U28970 (N_28970,N_27541,N_27385);
nor U28971 (N_28971,N_27554,N_27782);
nand U28972 (N_28972,N_27474,N_27717);
nor U28973 (N_28973,N_27349,N_27852);
nor U28974 (N_28974,N_27669,N_27007);
or U28975 (N_28975,N_27013,N_27325);
nor U28976 (N_28976,N_27189,N_27403);
nand U28977 (N_28977,N_27654,N_27305);
xnor U28978 (N_28978,N_27872,N_27130);
xnor U28979 (N_28979,N_27616,N_27473);
and U28980 (N_28980,N_27653,N_27169);
nand U28981 (N_28981,N_27441,N_27334);
nor U28982 (N_28982,N_27194,N_27570);
or U28983 (N_28983,N_27995,N_27289);
or U28984 (N_28984,N_27297,N_27557);
nand U28985 (N_28985,N_27705,N_27661);
and U28986 (N_28986,N_27117,N_27282);
nor U28987 (N_28987,N_27380,N_27548);
nor U28988 (N_28988,N_27613,N_27822);
or U28989 (N_28989,N_27326,N_27389);
xor U28990 (N_28990,N_27880,N_27767);
xor U28991 (N_28991,N_27146,N_27949);
nor U28992 (N_28992,N_27871,N_27550);
nand U28993 (N_28993,N_27689,N_27742);
xor U28994 (N_28994,N_27884,N_27385);
nor U28995 (N_28995,N_27659,N_27170);
nand U28996 (N_28996,N_27386,N_27350);
nand U28997 (N_28997,N_27901,N_27078);
xor U28998 (N_28998,N_27256,N_27794);
or U28999 (N_28999,N_27396,N_27398);
nand U29000 (N_29000,N_28843,N_28178);
nor U29001 (N_29001,N_28722,N_28236);
xor U29002 (N_29002,N_28195,N_28642);
nand U29003 (N_29003,N_28384,N_28139);
or U29004 (N_29004,N_28047,N_28716);
and U29005 (N_29005,N_28957,N_28652);
or U29006 (N_29006,N_28787,N_28617);
nor U29007 (N_29007,N_28588,N_28737);
nor U29008 (N_29008,N_28590,N_28846);
and U29009 (N_29009,N_28181,N_28557);
nand U29010 (N_29010,N_28503,N_28426);
or U29011 (N_29011,N_28659,N_28314);
nand U29012 (N_29012,N_28976,N_28167);
xor U29013 (N_29013,N_28979,N_28430);
nand U29014 (N_29014,N_28261,N_28033);
nand U29015 (N_29015,N_28940,N_28337);
or U29016 (N_29016,N_28247,N_28687);
nand U29017 (N_29017,N_28072,N_28855);
nand U29018 (N_29018,N_28292,N_28810);
nand U29019 (N_29019,N_28028,N_28419);
and U29020 (N_29020,N_28446,N_28582);
or U29021 (N_29021,N_28852,N_28682);
nor U29022 (N_29022,N_28772,N_28739);
nor U29023 (N_29023,N_28137,N_28632);
or U29024 (N_29024,N_28147,N_28003);
nand U29025 (N_29025,N_28796,N_28129);
or U29026 (N_29026,N_28297,N_28081);
and U29027 (N_29027,N_28216,N_28126);
and U29028 (N_29028,N_28197,N_28117);
nand U29029 (N_29029,N_28420,N_28404);
or U29030 (N_29030,N_28945,N_28403);
or U29031 (N_29031,N_28581,N_28202);
nand U29032 (N_29032,N_28781,N_28671);
nand U29033 (N_29033,N_28115,N_28792);
and U29034 (N_29034,N_28230,N_28738);
xnor U29035 (N_29035,N_28618,N_28941);
and U29036 (N_29036,N_28333,N_28146);
nand U29037 (N_29037,N_28828,N_28470);
and U29038 (N_29038,N_28054,N_28969);
nor U29039 (N_29039,N_28250,N_28519);
nand U29040 (N_29040,N_28764,N_28258);
xnor U29041 (N_29041,N_28901,N_28030);
xnor U29042 (N_29042,N_28443,N_28460);
nand U29043 (N_29043,N_28244,N_28599);
and U29044 (N_29044,N_28587,N_28410);
xor U29045 (N_29045,N_28449,N_28809);
xnor U29046 (N_29046,N_28733,N_28063);
and U29047 (N_29047,N_28748,N_28909);
xnor U29048 (N_29048,N_28508,N_28658);
nand U29049 (N_29049,N_28817,N_28741);
xnor U29050 (N_29050,N_28433,N_28592);
xnor U29051 (N_29051,N_28758,N_28083);
nand U29052 (N_29052,N_28098,N_28059);
and U29053 (N_29053,N_28623,N_28136);
or U29054 (N_29054,N_28660,N_28260);
nand U29055 (N_29055,N_28627,N_28832);
or U29056 (N_29056,N_28051,N_28637);
xor U29057 (N_29057,N_28208,N_28156);
xor U29058 (N_29058,N_28389,N_28283);
nand U29059 (N_29059,N_28994,N_28756);
and U29060 (N_29060,N_28308,N_28972);
nor U29061 (N_29061,N_28376,N_28076);
nor U29062 (N_29062,N_28541,N_28417);
nor U29063 (N_29063,N_28330,N_28980);
or U29064 (N_29064,N_28124,N_28094);
nand U29065 (N_29065,N_28844,N_28624);
xnor U29066 (N_29066,N_28188,N_28499);
and U29067 (N_29067,N_28513,N_28847);
nor U29068 (N_29068,N_28085,N_28349);
nand U29069 (N_29069,N_28301,N_28755);
nand U29070 (N_29070,N_28375,N_28552);
and U29071 (N_29071,N_28488,N_28401);
or U29072 (N_29072,N_28480,N_28039);
nor U29073 (N_29073,N_28769,N_28043);
xor U29074 (N_29074,N_28239,N_28092);
xnor U29075 (N_29075,N_28911,N_28254);
and U29076 (N_29076,N_28300,N_28062);
or U29077 (N_29077,N_28485,N_28171);
xnor U29078 (N_29078,N_28251,N_28646);
nand U29079 (N_29079,N_28439,N_28436);
nand U29080 (N_29080,N_28850,N_28892);
nand U29081 (N_29081,N_28670,N_28610);
nor U29082 (N_29082,N_28386,N_28021);
or U29083 (N_29083,N_28912,N_28935);
nand U29084 (N_29084,N_28408,N_28151);
or U29085 (N_29085,N_28473,N_28827);
nand U29086 (N_29086,N_28255,N_28857);
nand U29087 (N_29087,N_28790,N_28365);
nand U29088 (N_29088,N_28342,N_28999);
nor U29089 (N_29089,N_28992,N_28531);
and U29090 (N_29090,N_28876,N_28701);
and U29091 (N_29091,N_28037,N_28016);
nand U29092 (N_29092,N_28483,N_28138);
nor U29093 (N_29093,N_28690,N_28931);
xnor U29094 (N_29094,N_28593,N_28150);
nor U29095 (N_29095,N_28715,N_28162);
nand U29096 (N_29096,N_28311,N_28639);
nand U29097 (N_29097,N_28668,N_28416);
or U29098 (N_29098,N_28681,N_28411);
nand U29099 (N_29099,N_28257,N_28661);
or U29100 (N_29100,N_28740,N_28600);
nand U29101 (N_29101,N_28949,N_28108);
nor U29102 (N_29102,N_28077,N_28669);
xnor U29103 (N_29103,N_28192,N_28506);
nand U29104 (N_29104,N_28517,N_28774);
and U29105 (N_29105,N_28793,N_28641);
nand U29106 (N_29106,N_28112,N_28749);
and U29107 (N_29107,N_28042,N_28221);
xnor U29108 (N_29108,N_28731,N_28331);
and U29109 (N_29109,N_28630,N_28163);
nand U29110 (N_29110,N_28858,N_28607);
xnor U29111 (N_29111,N_28183,N_28169);
nand U29112 (N_29112,N_28194,N_28390);
and U29113 (N_29113,N_28626,N_28328);
or U29114 (N_29114,N_28206,N_28629);
nand U29115 (N_29115,N_28084,N_28451);
xor U29116 (N_29116,N_28939,N_28145);
nand U29117 (N_29117,N_28981,N_28152);
nand U29118 (N_29118,N_28921,N_28176);
nor U29119 (N_29119,N_28380,N_28482);
nand U29120 (N_29120,N_28636,N_28110);
nor U29121 (N_29121,N_28776,N_28611);
nor U29122 (N_29122,N_28805,N_28825);
nand U29123 (N_29123,N_28354,N_28452);
xor U29124 (N_29124,N_28780,N_28881);
nor U29125 (N_29125,N_28966,N_28768);
nand U29126 (N_29126,N_28823,N_28116);
and U29127 (N_29127,N_28276,N_28707);
nor U29128 (N_29128,N_28395,N_28179);
and U29129 (N_29129,N_28565,N_28511);
xor U29130 (N_29130,N_28227,N_28364);
or U29131 (N_29131,N_28559,N_28536);
and U29132 (N_29132,N_28685,N_28053);
xnor U29133 (N_29133,N_28154,N_28734);
and U29134 (N_29134,N_28427,N_28412);
nand U29135 (N_29135,N_28543,N_28019);
nor U29136 (N_29136,N_28873,N_28877);
and U29137 (N_29137,N_28664,N_28104);
or U29138 (N_29138,N_28710,N_28732);
or U29139 (N_29139,N_28878,N_28026);
nand U29140 (N_29140,N_28578,N_28907);
nand U29141 (N_29141,N_28281,N_28683);
nand U29142 (N_29142,N_28714,N_28285);
nor U29143 (N_29143,N_28533,N_28615);
or U29144 (N_29144,N_28951,N_28510);
xor U29145 (N_29145,N_28554,N_28555);
or U29146 (N_29146,N_28289,N_28985);
nand U29147 (N_29147,N_28340,N_28566);
or U29148 (N_29148,N_28421,N_28341);
nor U29149 (N_29149,N_28649,N_28445);
nand U29150 (N_29150,N_28943,N_28932);
xor U29151 (N_29151,N_28325,N_28620);
or U29152 (N_29152,N_28310,N_28351);
nor U29153 (N_29153,N_28274,N_28747);
and U29154 (N_29154,N_28381,N_28675);
and U29155 (N_29155,N_28879,N_28212);
nor U29156 (N_29156,N_28491,N_28672);
and U29157 (N_29157,N_28204,N_28135);
nand U29158 (N_29158,N_28918,N_28101);
and U29159 (N_29159,N_28215,N_28462);
or U29160 (N_29160,N_28391,N_28459);
nor U29161 (N_29161,N_28471,N_28968);
xnor U29162 (N_29162,N_28222,N_28867);
or U29163 (N_29163,N_28423,N_28914);
xor U29164 (N_29164,N_28840,N_28754);
nor U29165 (N_29165,N_28926,N_28928);
and U29166 (N_29166,N_28534,N_28561);
nand U29167 (N_29167,N_28367,N_28338);
and U29168 (N_29168,N_28686,N_28679);
or U29169 (N_29169,N_28699,N_28144);
and U29170 (N_29170,N_28930,N_28476);
nand U29171 (N_29171,N_28794,N_28698);
nand U29172 (N_29172,N_28778,N_28605);
nor U29173 (N_29173,N_28818,N_28291);
or U29174 (N_29174,N_28119,N_28157);
or U29175 (N_29175,N_28174,N_28882);
nor U29176 (N_29176,N_28429,N_28132);
and U29177 (N_29177,N_28345,N_28111);
and U29178 (N_29178,N_28424,N_28363);
or U29179 (N_29179,N_28551,N_28093);
or U29180 (N_29180,N_28650,N_28467);
and U29181 (N_29181,N_28086,N_28266);
and U29182 (N_29182,N_28315,N_28942);
and U29183 (N_29183,N_28529,N_28464);
and U29184 (N_29184,N_28572,N_28834);
or U29185 (N_29185,N_28967,N_28091);
nand U29186 (N_29186,N_28589,N_28223);
or U29187 (N_29187,N_28232,N_28360);
nor U29188 (N_29188,N_28773,N_28763);
nor U29189 (N_29189,N_28229,N_28512);
and U29190 (N_29190,N_28567,N_28068);
nor U29191 (N_29191,N_28456,N_28087);
and U29192 (N_29192,N_28305,N_28546);
or U29193 (N_29193,N_28831,N_28186);
xor U29194 (N_29194,N_28856,N_28450);
or U29195 (N_29195,N_28910,N_28346);
and U29196 (N_29196,N_28560,N_28288);
and U29197 (N_29197,N_28538,N_28321);
and U29198 (N_29198,N_28454,N_28388);
xor U29199 (N_29199,N_28872,N_28984);
or U29200 (N_29200,N_28184,N_28891);
and U29201 (N_29201,N_28307,N_28118);
and U29202 (N_29202,N_28044,N_28997);
nor U29203 (N_29203,N_28603,N_28596);
xnor U29204 (N_29204,N_28213,N_28908);
xor U29205 (N_29205,N_28676,N_28007);
and U29206 (N_29206,N_28893,N_28697);
xnor U29207 (N_29207,N_28720,N_28050);
and U29208 (N_29208,N_28556,N_28962);
nor U29209 (N_29209,N_28319,N_28457);
nand U29210 (N_29210,N_28800,N_28568);
or U29211 (N_29211,N_28000,N_28440);
or U29212 (N_29212,N_28718,N_28399);
and U29213 (N_29213,N_28861,N_28868);
or U29214 (N_29214,N_28608,N_28493);
xnor U29215 (N_29215,N_28514,N_28998);
xnor U29216 (N_29216,N_28383,N_28466);
xor U29217 (N_29217,N_28677,N_28955);
or U29218 (N_29218,N_28954,N_28574);
xnor U29219 (N_29219,N_28849,N_28622);
and U29220 (N_29220,N_28487,N_28518);
xnor U29221 (N_29221,N_28235,N_28965);
or U29222 (N_29222,N_28895,N_28760);
and U29223 (N_29223,N_28294,N_28695);
nor U29224 (N_29224,N_28278,N_28329);
and U29225 (N_29225,N_28180,N_28474);
and U29226 (N_29226,N_28708,N_28766);
xnor U29227 (N_29227,N_28521,N_28189);
and U29228 (N_29228,N_28128,N_28058);
and U29229 (N_29229,N_28437,N_28153);
nor U29230 (N_29230,N_28495,N_28634);
and U29231 (N_29231,N_28327,N_28286);
xor U29232 (N_29232,N_28075,N_28564);
xor U29233 (N_29233,N_28576,N_28114);
or U29234 (N_29234,N_28067,N_28752);
and U29235 (N_29235,N_28066,N_28570);
or U29236 (N_29236,N_28692,N_28079);
nand U29237 (N_29237,N_28366,N_28334);
and U29238 (N_29238,N_28964,N_28501);
nand U29239 (N_29239,N_28854,N_28220);
xor U29240 (N_29240,N_28869,N_28712);
or U29241 (N_29241,N_28548,N_28614);
and U29242 (N_29242,N_28020,N_28516);
nand U29243 (N_29243,N_28379,N_28061);
xnor U29244 (N_29244,N_28277,N_28502);
nand U29245 (N_29245,N_28666,N_28830);
nand U29246 (N_29246,N_28191,N_28326);
nand U29247 (N_29247,N_28874,N_28655);
nand U29248 (N_29248,N_28728,N_28762);
xnor U29249 (N_29249,N_28298,N_28963);
and U29250 (N_29250,N_28397,N_28371);
xnor U29251 (N_29251,N_28350,N_28819);
or U29252 (N_29252,N_28688,N_28958);
xor U29253 (N_29253,N_28448,N_28727);
or U29254 (N_29254,N_28761,N_28082);
and U29255 (N_29255,N_28526,N_28591);
nand U29256 (N_29256,N_28392,N_28583);
nand U29257 (N_29257,N_28065,N_28961);
and U29258 (N_29258,N_28324,N_28496);
nor U29259 (N_29259,N_28127,N_28296);
and U29260 (N_29260,N_28432,N_28977);
nor U29261 (N_29261,N_28268,N_28662);
nand U29262 (N_29262,N_28657,N_28807);
and U29263 (N_29263,N_28262,N_28175);
nand U29264 (N_29264,N_28120,N_28264);
nand U29265 (N_29265,N_28700,N_28396);
and U29266 (N_29266,N_28166,N_28031);
and U29267 (N_29267,N_28711,N_28725);
nand U29268 (N_29268,N_28249,N_28394);
or U29269 (N_29269,N_28929,N_28099);
nand U29270 (N_29270,N_28860,N_28187);
nor U29271 (N_29271,N_28055,N_28170);
nor U29272 (N_29272,N_28225,N_28013);
xnor U29273 (N_29273,N_28975,N_28263);
or U29274 (N_29274,N_28275,N_28241);
and U29275 (N_29275,N_28923,N_28060);
nor U29276 (N_29276,N_28418,N_28090);
xnor U29277 (N_29277,N_28505,N_28484);
nand U29278 (N_29278,N_28052,N_28024);
nor U29279 (N_29279,N_28034,N_28751);
and U29280 (N_29280,N_28829,N_28562);
and U29281 (N_29281,N_28045,N_28903);
and U29282 (N_29282,N_28097,N_28302);
and U29283 (N_29283,N_28804,N_28214);
xnor U29284 (N_29284,N_28571,N_28736);
or U29285 (N_29285,N_28211,N_28133);
xor U29286 (N_29286,N_28049,N_28207);
and U29287 (N_29287,N_28594,N_28073);
nor U29288 (N_29288,N_28273,N_28004);
and U29289 (N_29289,N_28015,N_28573);
nor U29290 (N_29290,N_28479,N_28469);
nand U29291 (N_29291,N_28237,N_28005);
nand U29292 (N_29292,N_28777,N_28633);
or U29293 (N_29293,N_28372,N_28332);
and U29294 (N_29294,N_28936,N_28841);
and U29295 (N_29295,N_28987,N_28447);
nor U29296 (N_29296,N_28231,N_28387);
nor U29297 (N_29297,N_28358,N_28883);
and U29298 (N_29298,N_28674,N_28498);
and U29299 (N_29299,N_28988,N_28284);
and U29300 (N_29300,N_28497,N_28706);
xor U29301 (N_29301,N_28402,N_28547);
and U29302 (N_29302,N_28875,N_28680);
xnor U29303 (N_29303,N_28933,N_28569);
xor U29304 (N_29304,N_28989,N_28287);
nor U29305 (N_29305,N_28735,N_28312);
and U29306 (N_29306,N_28259,N_28103);
nand U29307 (N_29307,N_28362,N_28201);
nor U29308 (N_29308,N_28651,N_28406);
or U29309 (N_29309,N_28673,N_28927);
nor U29310 (N_29310,N_28890,N_28463);
xor U29311 (N_29311,N_28172,N_28703);
and U29312 (N_29312,N_28504,N_28096);
nor U29313 (N_29313,N_28123,N_28228);
nand U29314 (N_29314,N_28509,N_28920);
nor U29315 (N_29315,N_28602,N_28960);
xnor U29316 (N_29316,N_28656,N_28647);
and U29317 (N_29317,N_28088,N_28267);
xor U29318 (N_29318,N_28377,N_28532);
nor U29319 (N_29319,N_28871,N_28667);
and U29320 (N_29320,N_28035,N_28428);
nor U29321 (N_29321,N_28434,N_28265);
xor U29322 (N_29322,N_28799,N_28782);
nand U29323 (N_29323,N_28057,N_28431);
and U29324 (N_29324,N_28545,N_28866);
xor U29325 (N_29325,N_28523,N_28226);
and U29326 (N_29326,N_28970,N_28356);
or U29327 (N_29327,N_28029,N_28444);
xnor U29328 (N_29328,N_28894,N_28640);
or U29329 (N_29329,N_28125,N_28313);
or U29330 (N_29330,N_28385,N_28937);
xnor U29331 (N_29331,N_28798,N_28036);
xnor U29332 (N_29332,N_28619,N_28813);
nand U29333 (N_29333,N_28783,N_28865);
nand U29334 (N_29334,N_28887,N_28134);
or U29335 (N_29335,N_28713,N_28643);
nand U29336 (N_29336,N_28767,N_28316);
xor U29337 (N_29337,N_28078,N_28986);
nand U29338 (N_29338,N_28048,N_28442);
or U29339 (N_29339,N_28527,N_28357);
or U29340 (N_29340,N_28374,N_28142);
nor U29341 (N_29341,N_28746,N_28595);
xnor U29342 (N_29342,N_28950,N_28904);
nor U29343 (N_29343,N_28757,N_28468);
xor U29344 (N_29344,N_28486,N_28859);
or U29345 (N_29345,N_28461,N_28352);
nand U29346 (N_29346,N_28753,N_28654);
xor U29347 (N_29347,N_28826,N_28884);
nor U29348 (N_29348,N_28665,N_28797);
nor U29349 (N_29349,N_28791,N_28190);
or U29350 (N_29350,N_28477,N_28899);
and U29351 (N_29351,N_28919,N_28472);
nand U29352 (N_29352,N_28822,N_28653);
xor U29353 (N_29353,N_28323,N_28322);
nand U29354 (N_29354,N_28347,N_28107);
nor U29355 (N_29355,N_28290,N_28027);
nor U29356 (N_29356,N_28272,N_28946);
nor U29357 (N_29357,N_28293,N_28824);
nor U29358 (N_29358,N_28056,N_28304);
and U29359 (N_29359,N_28801,N_28696);
and U29360 (N_29360,N_28438,N_28784);
xnor U29361 (N_29361,N_28648,N_28719);
or U29362 (N_29362,N_28282,N_28148);
nand U29363 (N_29363,N_28925,N_28540);
nor U29364 (N_29364,N_28168,N_28494);
nand U29365 (N_29365,N_28750,N_28130);
nor U29366 (N_29366,N_28730,N_28563);
nand U29367 (N_29367,N_28597,N_28956);
nor U29368 (N_29368,N_28089,N_28023);
nor U29369 (N_29369,N_28744,N_28638);
or U29370 (N_29370,N_28694,N_28795);
xnor U29371 (N_29371,N_28609,N_28100);
nor U29372 (N_29372,N_28205,N_28422);
or U29373 (N_29373,N_28368,N_28723);
nor U29374 (N_29374,N_28001,N_28539);
xor U29375 (N_29375,N_28243,N_28270);
nor U29376 (N_29376,N_28644,N_28253);
and U29377 (N_29377,N_28947,N_28425);
or U29378 (N_29378,N_28269,N_28726);
or U29379 (N_29379,N_28771,N_28155);
and U29380 (N_29380,N_28944,N_28811);
xnor U29381 (N_29381,N_28833,N_28271);
nor U29382 (N_29382,N_28398,N_28663);
nor U29383 (N_29383,N_28575,N_28765);
or U29384 (N_29384,N_28177,N_28924);
nand U29385 (N_29385,N_28369,N_28848);
or U29386 (N_29386,N_28990,N_28080);
or U29387 (N_29387,N_28458,N_28584);
nor U29388 (N_29388,N_28400,N_28018);
nand U29389 (N_29389,N_28631,N_28040);
xor U29390 (N_29390,N_28948,N_28789);
nor U29391 (N_29391,N_28489,N_28343);
and U29392 (N_29392,N_28318,N_28336);
and U29393 (N_29393,N_28069,N_28173);
nand U29394 (N_29394,N_28478,N_28074);
or U29395 (N_29395,N_28218,N_28759);
xor U29396 (N_29396,N_28806,N_28842);
nor U29397 (N_29397,N_28182,N_28185);
nor U29398 (N_29398,N_28544,N_28612);
nand U29399 (N_29399,N_28971,N_28689);
or U29400 (N_29400,N_28373,N_28886);
nor U29401 (N_29401,N_28993,N_28317);
or U29402 (N_29402,N_28070,N_28530);
nand U29403 (N_29403,N_28121,N_28558);
xnor U29404 (N_29404,N_28845,N_28238);
xnor U29405 (N_29405,N_28002,N_28779);
xnor U29406 (N_29406,N_28528,N_28233);
xnor U29407 (N_29407,N_28898,N_28978);
or U29408 (N_29408,N_28210,N_28645);
and U29409 (N_29409,N_28586,N_28815);
nand U29410 (N_29410,N_28934,N_28577);
or U29411 (N_29411,N_28678,N_28009);
nor U29412 (N_29412,N_28515,N_28014);
nor U29413 (N_29413,N_28888,N_28775);
nor U29414 (N_29414,N_28995,N_28837);
and U29415 (N_29415,N_28820,N_28729);
nor U29416 (N_29416,N_28038,N_28585);
xnor U29417 (N_29417,N_28006,N_28525);
nor U29418 (N_29418,N_28982,N_28938);
and U29419 (N_29419,N_28196,N_28522);
nor U29420 (N_29420,N_28628,N_28348);
nand U29421 (N_29421,N_28952,N_28041);
nand U29422 (N_29422,N_28724,N_28198);
and U29423 (N_29423,N_28248,N_28745);
and U29424 (N_29424,N_28953,N_28974);
nand U29425 (N_29425,N_28915,N_28008);
nor U29426 (N_29426,N_28973,N_28102);
xnor U29427 (N_29427,N_28355,N_28786);
nand U29428 (N_29428,N_28393,N_28335);
nand U29429 (N_29429,N_28299,N_28122);
xor U29430 (N_29430,N_28160,N_28245);
nand U29431 (N_29431,N_28621,N_28802);
nor U29432 (N_29432,N_28507,N_28481);
nand U29433 (N_29433,N_28158,N_28808);
and U29434 (N_29434,N_28240,N_28816);
nor U29435 (N_29435,N_28550,N_28885);
and U29436 (N_29436,N_28702,N_28870);
nand U29437 (N_29437,N_28704,N_28922);
and U29438 (N_29438,N_28071,N_28113);
or U29439 (N_29439,N_28475,N_28017);
or U29440 (N_29440,N_28022,N_28252);
xnor U29441 (N_29441,N_28361,N_28896);
nor U29442 (N_29442,N_28106,N_28897);
or U29443 (N_29443,N_28542,N_28520);
nor U29444 (N_29444,N_28200,N_28905);
xnor U29445 (N_29445,N_28131,N_28785);
nor U29446 (N_29446,N_28219,N_28812);
and U29447 (N_29447,N_28105,N_28579);
xnor U29448 (N_29448,N_28959,N_28500);
or U29449 (N_29449,N_28203,N_28889);
or U29450 (N_29450,N_28853,N_28295);
nor U29451 (N_29451,N_28705,N_28109);
and U29452 (N_29452,N_28902,N_28234);
or U29453 (N_29453,N_28161,N_28339);
nor U29454 (N_29454,N_28838,N_28164);
or U29455 (N_29455,N_28344,N_28917);
nor U29456 (N_29456,N_28435,N_28409);
nor U29457 (N_29457,N_28012,N_28246);
nor U29458 (N_29458,N_28625,N_28717);
or U29459 (N_29459,N_28580,N_28770);
nor U29460 (N_29460,N_28839,N_28309);
xor U29461 (N_29461,N_28613,N_28413);
xnor U29462 (N_29462,N_28835,N_28149);
nand U29463 (N_29463,N_28306,N_28721);
nor U29464 (N_29464,N_28535,N_28256);
and U29465 (N_29465,N_28320,N_28991);
nand U29466 (N_29466,N_28996,N_28370);
xor U29467 (N_29467,N_28913,N_28814);
nor U29468 (N_29468,N_28441,N_28906);
and U29469 (N_29469,N_28378,N_28635);
xnor U29470 (N_29470,N_28742,N_28916);
nand U29471 (N_29471,N_28803,N_28025);
or U29472 (N_29472,N_28046,N_28303);
xor U29473 (N_29473,N_28524,N_28095);
nor U29474 (N_29474,N_28863,N_28616);
or U29475 (N_29475,N_28064,N_28553);
xnor U29476 (N_29476,N_28143,N_28140);
nand U29477 (N_29477,N_28141,N_28193);
xnor U29478 (N_29478,N_28405,N_28490);
or U29479 (N_29479,N_28165,N_28862);
or U29480 (N_29480,N_28453,N_28414);
nand U29481 (N_29481,N_28159,N_28601);
nor U29482 (N_29482,N_28864,N_28851);
nor U29483 (N_29483,N_28604,N_28821);
and U29484 (N_29484,N_28382,N_28465);
nor U29485 (N_29485,N_28836,N_28549);
and U29486 (N_29486,N_28032,N_28691);
and U29487 (N_29487,N_28455,N_28010);
xnor U29488 (N_29488,N_28199,N_28415);
xor U29489 (N_29489,N_28224,N_28280);
or U29490 (N_29490,N_28684,N_28598);
or U29491 (N_29491,N_28880,N_28492);
nor U29492 (N_29492,N_28242,N_28743);
xor U29493 (N_29493,N_28353,N_28709);
nand U29494 (N_29494,N_28359,N_28983);
nand U29495 (N_29495,N_28693,N_28209);
and U29496 (N_29496,N_28011,N_28217);
or U29497 (N_29497,N_28407,N_28606);
nor U29498 (N_29498,N_28788,N_28279);
nand U29499 (N_29499,N_28537,N_28900);
and U29500 (N_29500,N_28892,N_28931);
or U29501 (N_29501,N_28283,N_28061);
nor U29502 (N_29502,N_28988,N_28755);
and U29503 (N_29503,N_28025,N_28510);
or U29504 (N_29504,N_28282,N_28984);
nor U29505 (N_29505,N_28843,N_28636);
nor U29506 (N_29506,N_28934,N_28122);
nand U29507 (N_29507,N_28112,N_28212);
xor U29508 (N_29508,N_28650,N_28795);
nor U29509 (N_29509,N_28885,N_28290);
or U29510 (N_29510,N_28659,N_28718);
nor U29511 (N_29511,N_28899,N_28985);
or U29512 (N_29512,N_28835,N_28011);
xnor U29513 (N_29513,N_28106,N_28020);
xor U29514 (N_29514,N_28147,N_28677);
nor U29515 (N_29515,N_28427,N_28544);
nand U29516 (N_29516,N_28057,N_28804);
and U29517 (N_29517,N_28786,N_28742);
xor U29518 (N_29518,N_28666,N_28257);
nor U29519 (N_29519,N_28069,N_28001);
and U29520 (N_29520,N_28965,N_28279);
nor U29521 (N_29521,N_28719,N_28098);
and U29522 (N_29522,N_28993,N_28667);
nor U29523 (N_29523,N_28584,N_28384);
xnor U29524 (N_29524,N_28073,N_28602);
or U29525 (N_29525,N_28945,N_28043);
xor U29526 (N_29526,N_28040,N_28455);
or U29527 (N_29527,N_28422,N_28901);
and U29528 (N_29528,N_28277,N_28194);
nor U29529 (N_29529,N_28259,N_28283);
or U29530 (N_29530,N_28650,N_28938);
xor U29531 (N_29531,N_28146,N_28747);
xnor U29532 (N_29532,N_28645,N_28398);
or U29533 (N_29533,N_28489,N_28327);
nor U29534 (N_29534,N_28391,N_28214);
xnor U29535 (N_29535,N_28155,N_28996);
xor U29536 (N_29536,N_28197,N_28082);
nand U29537 (N_29537,N_28889,N_28927);
nand U29538 (N_29538,N_28662,N_28168);
or U29539 (N_29539,N_28699,N_28169);
or U29540 (N_29540,N_28649,N_28003);
nor U29541 (N_29541,N_28794,N_28126);
nor U29542 (N_29542,N_28057,N_28476);
nand U29543 (N_29543,N_28468,N_28664);
xnor U29544 (N_29544,N_28779,N_28602);
nand U29545 (N_29545,N_28536,N_28411);
or U29546 (N_29546,N_28539,N_28167);
xnor U29547 (N_29547,N_28493,N_28416);
xnor U29548 (N_29548,N_28798,N_28243);
nor U29549 (N_29549,N_28818,N_28565);
or U29550 (N_29550,N_28944,N_28837);
nor U29551 (N_29551,N_28507,N_28679);
and U29552 (N_29552,N_28508,N_28114);
nand U29553 (N_29553,N_28387,N_28945);
and U29554 (N_29554,N_28724,N_28892);
nand U29555 (N_29555,N_28160,N_28503);
nor U29556 (N_29556,N_28785,N_28811);
nand U29557 (N_29557,N_28641,N_28438);
nand U29558 (N_29558,N_28448,N_28056);
and U29559 (N_29559,N_28720,N_28475);
nand U29560 (N_29560,N_28808,N_28743);
nand U29561 (N_29561,N_28917,N_28421);
or U29562 (N_29562,N_28458,N_28520);
or U29563 (N_29563,N_28576,N_28049);
nor U29564 (N_29564,N_28773,N_28741);
nor U29565 (N_29565,N_28139,N_28766);
and U29566 (N_29566,N_28648,N_28205);
xnor U29567 (N_29567,N_28994,N_28105);
nand U29568 (N_29568,N_28068,N_28862);
nand U29569 (N_29569,N_28920,N_28047);
or U29570 (N_29570,N_28012,N_28167);
or U29571 (N_29571,N_28467,N_28866);
nand U29572 (N_29572,N_28784,N_28511);
nor U29573 (N_29573,N_28247,N_28919);
nand U29574 (N_29574,N_28754,N_28665);
or U29575 (N_29575,N_28821,N_28150);
or U29576 (N_29576,N_28523,N_28035);
nand U29577 (N_29577,N_28909,N_28218);
xnor U29578 (N_29578,N_28727,N_28141);
nand U29579 (N_29579,N_28732,N_28172);
and U29580 (N_29580,N_28870,N_28297);
nand U29581 (N_29581,N_28396,N_28535);
nand U29582 (N_29582,N_28887,N_28524);
and U29583 (N_29583,N_28142,N_28322);
and U29584 (N_29584,N_28405,N_28996);
or U29585 (N_29585,N_28775,N_28124);
xnor U29586 (N_29586,N_28903,N_28188);
nand U29587 (N_29587,N_28881,N_28999);
nor U29588 (N_29588,N_28651,N_28454);
nor U29589 (N_29589,N_28115,N_28950);
nand U29590 (N_29590,N_28359,N_28757);
nor U29591 (N_29591,N_28395,N_28814);
xor U29592 (N_29592,N_28496,N_28258);
or U29593 (N_29593,N_28940,N_28385);
nand U29594 (N_29594,N_28035,N_28450);
nand U29595 (N_29595,N_28788,N_28135);
nor U29596 (N_29596,N_28121,N_28156);
or U29597 (N_29597,N_28292,N_28378);
and U29598 (N_29598,N_28292,N_28821);
and U29599 (N_29599,N_28114,N_28187);
xor U29600 (N_29600,N_28266,N_28059);
nand U29601 (N_29601,N_28192,N_28562);
and U29602 (N_29602,N_28591,N_28482);
nor U29603 (N_29603,N_28082,N_28456);
nand U29604 (N_29604,N_28288,N_28712);
and U29605 (N_29605,N_28813,N_28820);
nand U29606 (N_29606,N_28159,N_28539);
nor U29607 (N_29607,N_28666,N_28988);
nand U29608 (N_29608,N_28613,N_28553);
or U29609 (N_29609,N_28022,N_28863);
nand U29610 (N_29610,N_28401,N_28835);
and U29611 (N_29611,N_28522,N_28417);
or U29612 (N_29612,N_28848,N_28505);
and U29613 (N_29613,N_28607,N_28165);
nor U29614 (N_29614,N_28362,N_28638);
nand U29615 (N_29615,N_28669,N_28373);
xnor U29616 (N_29616,N_28371,N_28987);
xor U29617 (N_29617,N_28568,N_28282);
and U29618 (N_29618,N_28181,N_28568);
nand U29619 (N_29619,N_28973,N_28532);
nand U29620 (N_29620,N_28374,N_28426);
nor U29621 (N_29621,N_28742,N_28534);
nand U29622 (N_29622,N_28600,N_28677);
or U29623 (N_29623,N_28053,N_28170);
xnor U29624 (N_29624,N_28989,N_28820);
xnor U29625 (N_29625,N_28256,N_28997);
xnor U29626 (N_29626,N_28241,N_28682);
nand U29627 (N_29627,N_28766,N_28627);
xnor U29628 (N_29628,N_28607,N_28849);
nor U29629 (N_29629,N_28741,N_28121);
xnor U29630 (N_29630,N_28992,N_28058);
or U29631 (N_29631,N_28397,N_28664);
xnor U29632 (N_29632,N_28038,N_28099);
and U29633 (N_29633,N_28179,N_28929);
xnor U29634 (N_29634,N_28575,N_28147);
nor U29635 (N_29635,N_28363,N_28598);
xnor U29636 (N_29636,N_28168,N_28611);
and U29637 (N_29637,N_28473,N_28238);
nor U29638 (N_29638,N_28889,N_28989);
or U29639 (N_29639,N_28546,N_28562);
nor U29640 (N_29640,N_28466,N_28902);
and U29641 (N_29641,N_28113,N_28967);
or U29642 (N_29642,N_28165,N_28307);
or U29643 (N_29643,N_28242,N_28561);
nor U29644 (N_29644,N_28474,N_28129);
and U29645 (N_29645,N_28986,N_28403);
or U29646 (N_29646,N_28089,N_28549);
xnor U29647 (N_29647,N_28549,N_28160);
nor U29648 (N_29648,N_28576,N_28669);
nand U29649 (N_29649,N_28820,N_28120);
xor U29650 (N_29650,N_28060,N_28770);
xnor U29651 (N_29651,N_28478,N_28754);
nor U29652 (N_29652,N_28350,N_28780);
or U29653 (N_29653,N_28810,N_28613);
and U29654 (N_29654,N_28294,N_28833);
nor U29655 (N_29655,N_28168,N_28626);
xnor U29656 (N_29656,N_28169,N_28488);
nand U29657 (N_29657,N_28267,N_28274);
xor U29658 (N_29658,N_28731,N_28468);
or U29659 (N_29659,N_28886,N_28610);
nand U29660 (N_29660,N_28211,N_28742);
or U29661 (N_29661,N_28599,N_28495);
and U29662 (N_29662,N_28147,N_28930);
nand U29663 (N_29663,N_28022,N_28462);
and U29664 (N_29664,N_28079,N_28417);
nor U29665 (N_29665,N_28381,N_28761);
nand U29666 (N_29666,N_28677,N_28936);
nand U29667 (N_29667,N_28308,N_28287);
nor U29668 (N_29668,N_28852,N_28046);
xnor U29669 (N_29669,N_28807,N_28027);
nand U29670 (N_29670,N_28419,N_28159);
xor U29671 (N_29671,N_28053,N_28161);
nand U29672 (N_29672,N_28253,N_28500);
and U29673 (N_29673,N_28689,N_28256);
nor U29674 (N_29674,N_28740,N_28918);
xor U29675 (N_29675,N_28856,N_28717);
or U29676 (N_29676,N_28556,N_28593);
xor U29677 (N_29677,N_28832,N_28915);
or U29678 (N_29678,N_28203,N_28851);
nand U29679 (N_29679,N_28611,N_28585);
nand U29680 (N_29680,N_28452,N_28468);
and U29681 (N_29681,N_28402,N_28859);
or U29682 (N_29682,N_28295,N_28244);
or U29683 (N_29683,N_28976,N_28623);
or U29684 (N_29684,N_28445,N_28105);
nor U29685 (N_29685,N_28503,N_28806);
nor U29686 (N_29686,N_28241,N_28692);
and U29687 (N_29687,N_28376,N_28809);
xor U29688 (N_29688,N_28425,N_28179);
or U29689 (N_29689,N_28030,N_28103);
nand U29690 (N_29690,N_28534,N_28180);
nor U29691 (N_29691,N_28584,N_28706);
and U29692 (N_29692,N_28528,N_28457);
or U29693 (N_29693,N_28628,N_28985);
nand U29694 (N_29694,N_28410,N_28084);
nor U29695 (N_29695,N_28036,N_28517);
nand U29696 (N_29696,N_28612,N_28310);
or U29697 (N_29697,N_28238,N_28326);
nand U29698 (N_29698,N_28946,N_28963);
and U29699 (N_29699,N_28738,N_28724);
and U29700 (N_29700,N_28726,N_28625);
nand U29701 (N_29701,N_28503,N_28841);
or U29702 (N_29702,N_28578,N_28217);
and U29703 (N_29703,N_28318,N_28643);
and U29704 (N_29704,N_28747,N_28703);
xnor U29705 (N_29705,N_28707,N_28095);
or U29706 (N_29706,N_28822,N_28278);
nand U29707 (N_29707,N_28783,N_28739);
xnor U29708 (N_29708,N_28400,N_28095);
and U29709 (N_29709,N_28576,N_28622);
nor U29710 (N_29710,N_28958,N_28620);
xnor U29711 (N_29711,N_28211,N_28072);
or U29712 (N_29712,N_28840,N_28974);
nand U29713 (N_29713,N_28952,N_28977);
nor U29714 (N_29714,N_28148,N_28864);
nor U29715 (N_29715,N_28857,N_28681);
nand U29716 (N_29716,N_28034,N_28950);
and U29717 (N_29717,N_28164,N_28109);
and U29718 (N_29718,N_28789,N_28753);
or U29719 (N_29719,N_28252,N_28670);
nand U29720 (N_29720,N_28812,N_28404);
or U29721 (N_29721,N_28249,N_28737);
nor U29722 (N_29722,N_28942,N_28101);
xor U29723 (N_29723,N_28461,N_28887);
xnor U29724 (N_29724,N_28080,N_28237);
xnor U29725 (N_29725,N_28826,N_28241);
xor U29726 (N_29726,N_28583,N_28047);
and U29727 (N_29727,N_28386,N_28330);
xnor U29728 (N_29728,N_28136,N_28361);
xnor U29729 (N_29729,N_28995,N_28808);
and U29730 (N_29730,N_28538,N_28227);
nand U29731 (N_29731,N_28275,N_28301);
or U29732 (N_29732,N_28715,N_28765);
nand U29733 (N_29733,N_28077,N_28855);
nand U29734 (N_29734,N_28117,N_28881);
or U29735 (N_29735,N_28484,N_28661);
xor U29736 (N_29736,N_28379,N_28009);
nand U29737 (N_29737,N_28949,N_28670);
or U29738 (N_29738,N_28285,N_28090);
nand U29739 (N_29739,N_28059,N_28388);
xor U29740 (N_29740,N_28689,N_28633);
and U29741 (N_29741,N_28794,N_28246);
nand U29742 (N_29742,N_28286,N_28060);
nor U29743 (N_29743,N_28972,N_28661);
xor U29744 (N_29744,N_28381,N_28966);
nor U29745 (N_29745,N_28756,N_28925);
nand U29746 (N_29746,N_28918,N_28495);
and U29747 (N_29747,N_28200,N_28152);
nor U29748 (N_29748,N_28717,N_28872);
nor U29749 (N_29749,N_28033,N_28227);
xor U29750 (N_29750,N_28825,N_28146);
xor U29751 (N_29751,N_28994,N_28484);
nand U29752 (N_29752,N_28042,N_28149);
and U29753 (N_29753,N_28202,N_28459);
nor U29754 (N_29754,N_28511,N_28826);
xor U29755 (N_29755,N_28806,N_28520);
or U29756 (N_29756,N_28821,N_28459);
nor U29757 (N_29757,N_28344,N_28157);
and U29758 (N_29758,N_28951,N_28542);
xor U29759 (N_29759,N_28046,N_28883);
nand U29760 (N_29760,N_28575,N_28502);
and U29761 (N_29761,N_28716,N_28428);
and U29762 (N_29762,N_28815,N_28712);
nor U29763 (N_29763,N_28463,N_28953);
xnor U29764 (N_29764,N_28810,N_28415);
nand U29765 (N_29765,N_28914,N_28560);
xor U29766 (N_29766,N_28164,N_28726);
nand U29767 (N_29767,N_28436,N_28487);
nor U29768 (N_29768,N_28144,N_28943);
and U29769 (N_29769,N_28250,N_28255);
nor U29770 (N_29770,N_28159,N_28567);
xnor U29771 (N_29771,N_28079,N_28613);
and U29772 (N_29772,N_28409,N_28821);
nand U29773 (N_29773,N_28506,N_28709);
nand U29774 (N_29774,N_28267,N_28401);
xnor U29775 (N_29775,N_28361,N_28334);
and U29776 (N_29776,N_28982,N_28564);
nor U29777 (N_29777,N_28514,N_28251);
nor U29778 (N_29778,N_28332,N_28278);
and U29779 (N_29779,N_28956,N_28725);
nand U29780 (N_29780,N_28548,N_28437);
xor U29781 (N_29781,N_28083,N_28275);
xor U29782 (N_29782,N_28353,N_28916);
or U29783 (N_29783,N_28892,N_28096);
nor U29784 (N_29784,N_28707,N_28522);
or U29785 (N_29785,N_28680,N_28786);
and U29786 (N_29786,N_28059,N_28503);
xor U29787 (N_29787,N_28690,N_28491);
xnor U29788 (N_29788,N_28452,N_28277);
nor U29789 (N_29789,N_28204,N_28854);
nand U29790 (N_29790,N_28419,N_28725);
xor U29791 (N_29791,N_28304,N_28209);
nor U29792 (N_29792,N_28953,N_28354);
or U29793 (N_29793,N_28757,N_28911);
or U29794 (N_29794,N_28893,N_28569);
or U29795 (N_29795,N_28024,N_28669);
nor U29796 (N_29796,N_28549,N_28120);
or U29797 (N_29797,N_28011,N_28059);
nand U29798 (N_29798,N_28494,N_28913);
and U29799 (N_29799,N_28588,N_28318);
and U29800 (N_29800,N_28945,N_28338);
xor U29801 (N_29801,N_28093,N_28812);
and U29802 (N_29802,N_28697,N_28861);
and U29803 (N_29803,N_28671,N_28661);
nor U29804 (N_29804,N_28076,N_28288);
or U29805 (N_29805,N_28584,N_28518);
xor U29806 (N_29806,N_28956,N_28975);
nor U29807 (N_29807,N_28466,N_28071);
or U29808 (N_29808,N_28070,N_28574);
nand U29809 (N_29809,N_28016,N_28643);
nor U29810 (N_29810,N_28901,N_28185);
nor U29811 (N_29811,N_28907,N_28213);
and U29812 (N_29812,N_28268,N_28226);
nand U29813 (N_29813,N_28259,N_28211);
or U29814 (N_29814,N_28632,N_28493);
xor U29815 (N_29815,N_28523,N_28806);
and U29816 (N_29816,N_28804,N_28756);
nor U29817 (N_29817,N_28219,N_28652);
nand U29818 (N_29818,N_28506,N_28261);
or U29819 (N_29819,N_28092,N_28189);
nor U29820 (N_29820,N_28929,N_28734);
and U29821 (N_29821,N_28801,N_28231);
nand U29822 (N_29822,N_28406,N_28890);
and U29823 (N_29823,N_28922,N_28888);
and U29824 (N_29824,N_28643,N_28873);
xnor U29825 (N_29825,N_28021,N_28602);
or U29826 (N_29826,N_28826,N_28975);
or U29827 (N_29827,N_28450,N_28481);
or U29828 (N_29828,N_28168,N_28613);
xor U29829 (N_29829,N_28471,N_28969);
nor U29830 (N_29830,N_28679,N_28727);
and U29831 (N_29831,N_28799,N_28016);
xor U29832 (N_29832,N_28979,N_28363);
and U29833 (N_29833,N_28784,N_28162);
xor U29834 (N_29834,N_28473,N_28550);
xnor U29835 (N_29835,N_28357,N_28734);
xor U29836 (N_29836,N_28075,N_28143);
or U29837 (N_29837,N_28763,N_28067);
nor U29838 (N_29838,N_28526,N_28954);
xor U29839 (N_29839,N_28281,N_28225);
xor U29840 (N_29840,N_28360,N_28110);
or U29841 (N_29841,N_28838,N_28858);
nor U29842 (N_29842,N_28270,N_28823);
nand U29843 (N_29843,N_28431,N_28165);
nor U29844 (N_29844,N_28585,N_28370);
xor U29845 (N_29845,N_28303,N_28185);
nor U29846 (N_29846,N_28602,N_28422);
nand U29847 (N_29847,N_28132,N_28434);
xnor U29848 (N_29848,N_28240,N_28744);
nand U29849 (N_29849,N_28092,N_28369);
nor U29850 (N_29850,N_28083,N_28415);
or U29851 (N_29851,N_28562,N_28868);
nand U29852 (N_29852,N_28236,N_28940);
or U29853 (N_29853,N_28981,N_28835);
or U29854 (N_29854,N_28995,N_28597);
xor U29855 (N_29855,N_28218,N_28401);
and U29856 (N_29856,N_28919,N_28392);
nor U29857 (N_29857,N_28888,N_28497);
or U29858 (N_29858,N_28078,N_28043);
xnor U29859 (N_29859,N_28717,N_28051);
nor U29860 (N_29860,N_28970,N_28977);
and U29861 (N_29861,N_28890,N_28743);
or U29862 (N_29862,N_28998,N_28922);
or U29863 (N_29863,N_28394,N_28742);
or U29864 (N_29864,N_28415,N_28745);
nand U29865 (N_29865,N_28592,N_28752);
nand U29866 (N_29866,N_28056,N_28405);
nor U29867 (N_29867,N_28221,N_28520);
nand U29868 (N_29868,N_28036,N_28429);
nor U29869 (N_29869,N_28093,N_28221);
nand U29870 (N_29870,N_28623,N_28862);
or U29871 (N_29871,N_28237,N_28732);
nand U29872 (N_29872,N_28200,N_28735);
xnor U29873 (N_29873,N_28589,N_28072);
nand U29874 (N_29874,N_28780,N_28742);
nor U29875 (N_29875,N_28463,N_28970);
or U29876 (N_29876,N_28255,N_28244);
xnor U29877 (N_29877,N_28937,N_28172);
nand U29878 (N_29878,N_28732,N_28163);
and U29879 (N_29879,N_28132,N_28977);
nor U29880 (N_29880,N_28923,N_28389);
nand U29881 (N_29881,N_28191,N_28911);
xnor U29882 (N_29882,N_28984,N_28243);
nand U29883 (N_29883,N_28963,N_28538);
and U29884 (N_29884,N_28024,N_28099);
nand U29885 (N_29885,N_28963,N_28781);
xor U29886 (N_29886,N_28847,N_28202);
and U29887 (N_29887,N_28621,N_28807);
and U29888 (N_29888,N_28815,N_28441);
and U29889 (N_29889,N_28034,N_28910);
nand U29890 (N_29890,N_28978,N_28101);
xor U29891 (N_29891,N_28990,N_28973);
xnor U29892 (N_29892,N_28611,N_28985);
xnor U29893 (N_29893,N_28143,N_28125);
nor U29894 (N_29894,N_28608,N_28786);
nand U29895 (N_29895,N_28246,N_28745);
or U29896 (N_29896,N_28648,N_28217);
or U29897 (N_29897,N_28082,N_28053);
xor U29898 (N_29898,N_28109,N_28036);
nand U29899 (N_29899,N_28127,N_28187);
xnor U29900 (N_29900,N_28460,N_28473);
nand U29901 (N_29901,N_28739,N_28491);
nor U29902 (N_29902,N_28087,N_28761);
and U29903 (N_29903,N_28691,N_28200);
nand U29904 (N_29904,N_28590,N_28851);
nor U29905 (N_29905,N_28270,N_28414);
nand U29906 (N_29906,N_28880,N_28098);
nand U29907 (N_29907,N_28012,N_28850);
nand U29908 (N_29908,N_28345,N_28998);
nor U29909 (N_29909,N_28883,N_28645);
or U29910 (N_29910,N_28028,N_28942);
nand U29911 (N_29911,N_28679,N_28040);
xnor U29912 (N_29912,N_28003,N_28496);
and U29913 (N_29913,N_28359,N_28801);
nand U29914 (N_29914,N_28552,N_28173);
nand U29915 (N_29915,N_28055,N_28441);
nor U29916 (N_29916,N_28347,N_28106);
xor U29917 (N_29917,N_28316,N_28918);
and U29918 (N_29918,N_28205,N_28288);
nor U29919 (N_29919,N_28100,N_28627);
or U29920 (N_29920,N_28311,N_28169);
or U29921 (N_29921,N_28989,N_28355);
xnor U29922 (N_29922,N_28356,N_28119);
nor U29923 (N_29923,N_28863,N_28732);
xor U29924 (N_29924,N_28585,N_28033);
nor U29925 (N_29925,N_28126,N_28976);
xor U29926 (N_29926,N_28871,N_28535);
and U29927 (N_29927,N_28844,N_28383);
and U29928 (N_29928,N_28780,N_28107);
and U29929 (N_29929,N_28100,N_28853);
and U29930 (N_29930,N_28839,N_28658);
or U29931 (N_29931,N_28102,N_28846);
or U29932 (N_29932,N_28842,N_28180);
and U29933 (N_29933,N_28767,N_28274);
nand U29934 (N_29934,N_28965,N_28381);
or U29935 (N_29935,N_28494,N_28923);
and U29936 (N_29936,N_28724,N_28700);
and U29937 (N_29937,N_28692,N_28019);
or U29938 (N_29938,N_28086,N_28866);
nor U29939 (N_29939,N_28558,N_28832);
xnor U29940 (N_29940,N_28013,N_28124);
xor U29941 (N_29941,N_28317,N_28899);
nor U29942 (N_29942,N_28125,N_28843);
nand U29943 (N_29943,N_28208,N_28535);
xor U29944 (N_29944,N_28254,N_28773);
and U29945 (N_29945,N_28514,N_28264);
and U29946 (N_29946,N_28585,N_28754);
or U29947 (N_29947,N_28467,N_28769);
xor U29948 (N_29948,N_28507,N_28944);
or U29949 (N_29949,N_28665,N_28545);
nand U29950 (N_29950,N_28760,N_28649);
nand U29951 (N_29951,N_28629,N_28771);
or U29952 (N_29952,N_28583,N_28237);
nand U29953 (N_29953,N_28893,N_28641);
nor U29954 (N_29954,N_28993,N_28966);
or U29955 (N_29955,N_28326,N_28537);
xor U29956 (N_29956,N_28630,N_28549);
and U29957 (N_29957,N_28662,N_28462);
xor U29958 (N_29958,N_28153,N_28134);
nand U29959 (N_29959,N_28668,N_28106);
xnor U29960 (N_29960,N_28071,N_28024);
and U29961 (N_29961,N_28135,N_28213);
nor U29962 (N_29962,N_28941,N_28734);
or U29963 (N_29963,N_28005,N_28851);
nand U29964 (N_29964,N_28269,N_28080);
nor U29965 (N_29965,N_28089,N_28610);
or U29966 (N_29966,N_28863,N_28832);
nand U29967 (N_29967,N_28163,N_28019);
and U29968 (N_29968,N_28098,N_28599);
nor U29969 (N_29969,N_28802,N_28456);
xor U29970 (N_29970,N_28633,N_28940);
xor U29971 (N_29971,N_28286,N_28953);
xor U29972 (N_29972,N_28525,N_28385);
xor U29973 (N_29973,N_28670,N_28018);
and U29974 (N_29974,N_28036,N_28762);
and U29975 (N_29975,N_28800,N_28464);
nand U29976 (N_29976,N_28427,N_28319);
nor U29977 (N_29977,N_28236,N_28844);
xor U29978 (N_29978,N_28673,N_28282);
and U29979 (N_29979,N_28706,N_28872);
xor U29980 (N_29980,N_28628,N_28794);
nor U29981 (N_29981,N_28329,N_28726);
nor U29982 (N_29982,N_28578,N_28868);
nor U29983 (N_29983,N_28216,N_28309);
nor U29984 (N_29984,N_28366,N_28202);
and U29985 (N_29985,N_28440,N_28324);
xor U29986 (N_29986,N_28727,N_28501);
xnor U29987 (N_29987,N_28658,N_28087);
nor U29988 (N_29988,N_28192,N_28182);
or U29989 (N_29989,N_28004,N_28821);
or U29990 (N_29990,N_28999,N_28495);
and U29991 (N_29991,N_28781,N_28995);
or U29992 (N_29992,N_28861,N_28986);
nor U29993 (N_29993,N_28422,N_28958);
or U29994 (N_29994,N_28358,N_28660);
xor U29995 (N_29995,N_28066,N_28103);
nor U29996 (N_29996,N_28159,N_28016);
and U29997 (N_29997,N_28838,N_28034);
nor U29998 (N_29998,N_28036,N_28651);
nand U29999 (N_29999,N_28573,N_28443);
and U30000 (N_30000,N_29087,N_29635);
and U30001 (N_30001,N_29423,N_29319);
or U30002 (N_30002,N_29771,N_29745);
xnor U30003 (N_30003,N_29311,N_29980);
nor U30004 (N_30004,N_29967,N_29168);
nor U30005 (N_30005,N_29075,N_29554);
nor U30006 (N_30006,N_29058,N_29751);
nor U30007 (N_30007,N_29563,N_29203);
nand U30008 (N_30008,N_29723,N_29436);
or U30009 (N_30009,N_29976,N_29930);
and U30010 (N_30010,N_29792,N_29542);
xor U30011 (N_30011,N_29935,N_29505);
nor U30012 (N_30012,N_29199,N_29948);
nor U30013 (N_30013,N_29756,N_29581);
nand U30014 (N_30014,N_29130,N_29177);
nor U30015 (N_30015,N_29000,N_29790);
and U30016 (N_30016,N_29955,N_29021);
nor U30017 (N_30017,N_29424,N_29922);
xor U30018 (N_30018,N_29874,N_29913);
and U30019 (N_30019,N_29559,N_29172);
or U30020 (N_30020,N_29103,N_29896);
xnor U30021 (N_30021,N_29959,N_29812);
xor U30022 (N_30022,N_29093,N_29176);
nor U30023 (N_30023,N_29739,N_29750);
xnor U30024 (N_30024,N_29866,N_29523);
and U30025 (N_30025,N_29947,N_29125);
and U30026 (N_30026,N_29462,N_29032);
and U30027 (N_30027,N_29919,N_29720);
nand U30028 (N_30028,N_29736,N_29583);
or U30029 (N_30029,N_29134,N_29915);
xnor U30030 (N_30030,N_29666,N_29208);
xor U30031 (N_30031,N_29492,N_29634);
nor U30032 (N_30032,N_29908,N_29502);
xor U30033 (N_30033,N_29050,N_29419);
nor U30034 (N_30034,N_29317,N_29326);
xnor U30035 (N_30035,N_29167,N_29937);
or U30036 (N_30036,N_29119,N_29071);
nor U30037 (N_30037,N_29705,N_29840);
nor U30038 (N_30038,N_29104,N_29612);
xor U30039 (N_30039,N_29073,N_29615);
and U30040 (N_30040,N_29527,N_29604);
or U30041 (N_30041,N_29096,N_29216);
nor U30042 (N_30042,N_29137,N_29392);
xnor U30043 (N_30043,N_29290,N_29831);
nor U30044 (N_30044,N_29782,N_29701);
nand U30045 (N_30045,N_29297,N_29191);
xor U30046 (N_30046,N_29507,N_29257);
nand U30047 (N_30047,N_29360,N_29886);
nor U30048 (N_30048,N_29764,N_29689);
or U30049 (N_30049,N_29625,N_29522);
or U30050 (N_30050,N_29649,N_29135);
nand U30051 (N_30051,N_29642,N_29110);
xor U30052 (N_30052,N_29025,N_29999);
nand U30053 (N_30053,N_29275,N_29148);
xnor U30054 (N_30054,N_29893,N_29152);
nor U30055 (N_30055,N_29925,N_29306);
or U30056 (N_30056,N_29802,N_29828);
or U30057 (N_30057,N_29882,N_29579);
nor U30058 (N_30058,N_29232,N_29270);
xor U30059 (N_30059,N_29658,N_29222);
xor U30060 (N_30060,N_29267,N_29427);
or U30061 (N_30061,N_29993,N_29433);
and U30062 (N_30062,N_29911,N_29713);
nor U30063 (N_30063,N_29706,N_29430);
or U30064 (N_30064,N_29968,N_29154);
nor U30065 (N_30065,N_29160,N_29421);
and U30066 (N_30066,N_29344,N_29243);
nand U30067 (N_30067,N_29046,N_29490);
nor U30068 (N_30068,N_29962,N_29384);
and U30069 (N_30069,N_29719,N_29459);
nand U30070 (N_30070,N_29084,N_29241);
nor U30071 (N_30071,N_29928,N_29970);
or U30072 (N_30072,N_29905,N_29389);
nand U30073 (N_30073,N_29985,N_29182);
and U30074 (N_30074,N_29259,N_29287);
nor U30075 (N_30075,N_29582,N_29906);
and U30076 (N_30076,N_29858,N_29795);
and U30077 (N_30077,N_29853,N_29048);
and U30078 (N_30078,N_29310,N_29730);
and U30079 (N_30079,N_29499,N_29686);
or U30080 (N_30080,N_29741,N_29616);
or U30081 (N_30081,N_29005,N_29098);
nand U30082 (N_30082,N_29877,N_29388);
or U30083 (N_30083,N_29255,N_29367);
and U30084 (N_30084,N_29153,N_29619);
nor U30085 (N_30085,N_29480,N_29406);
nor U30086 (N_30086,N_29489,N_29724);
nand U30087 (N_30087,N_29975,N_29843);
and U30088 (N_30088,N_29218,N_29230);
xnor U30089 (N_30089,N_29195,N_29054);
or U30090 (N_30090,N_29322,N_29260);
nand U30091 (N_30091,N_29456,N_29451);
and U30092 (N_30092,N_29690,N_29747);
nor U30093 (N_30093,N_29857,N_29276);
and U30094 (N_30094,N_29385,N_29114);
nor U30095 (N_30095,N_29233,N_29161);
nand U30096 (N_30096,N_29892,N_29921);
and U30097 (N_30097,N_29258,N_29691);
nand U30098 (N_30098,N_29425,N_29571);
and U30099 (N_30099,N_29386,N_29431);
and U30100 (N_30100,N_29924,N_29065);
xnor U30101 (N_30101,N_29128,N_29136);
xor U30102 (N_30102,N_29219,N_29851);
and U30103 (N_30103,N_29943,N_29081);
nand U30104 (N_30104,N_29361,N_29336);
nand U30105 (N_30105,N_29051,N_29530);
and U30106 (N_30106,N_29078,N_29210);
xor U30107 (N_30107,N_29618,N_29282);
nand U30108 (N_30108,N_29163,N_29052);
or U30109 (N_30109,N_29272,N_29638);
and U30110 (N_30110,N_29965,N_29503);
and U30111 (N_30111,N_29300,N_29209);
nand U30112 (N_30112,N_29022,N_29623);
xnor U30113 (N_30113,N_29823,N_29335);
nand U30114 (N_30114,N_29028,N_29568);
or U30115 (N_30115,N_29510,N_29446);
or U30116 (N_30116,N_29034,N_29629);
nand U30117 (N_30117,N_29438,N_29536);
and U30118 (N_30118,N_29403,N_29268);
or U30119 (N_30119,N_29998,N_29767);
nand U30120 (N_30120,N_29670,N_29907);
xor U30121 (N_30121,N_29526,N_29483);
nor U30122 (N_30122,N_29097,N_29914);
xor U30123 (N_30123,N_29090,N_29320);
nand U30124 (N_30124,N_29504,N_29945);
nand U30125 (N_30125,N_29017,N_29498);
or U30126 (N_30126,N_29997,N_29733);
xnor U30127 (N_30127,N_29067,N_29363);
nor U30128 (N_30128,N_29331,N_29482);
nand U30129 (N_30129,N_29340,N_29165);
xor U30130 (N_30130,N_29584,N_29781);
and U30131 (N_30131,N_29121,N_29334);
nor U30132 (N_30132,N_29951,N_29819);
nand U30133 (N_30133,N_29752,N_29465);
and U30134 (N_30134,N_29697,N_29683);
nor U30135 (N_30135,N_29029,N_29227);
and U30136 (N_30136,N_29555,N_29605);
nor U30137 (N_30137,N_29133,N_29197);
and U30138 (N_30138,N_29547,N_29417);
or U30139 (N_30139,N_29007,N_29570);
nand U30140 (N_30140,N_29718,N_29765);
or U30141 (N_30141,N_29606,N_29013);
or U30142 (N_30142,N_29657,N_29693);
and U30143 (N_30143,N_29211,N_29374);
nor U30144 (N_30144,N_29445,N_29743);
or U30145 (N_30145,N_29788,N_29901);
and U30146 (N_30146,N_29162,N_29453);
nor U30147 (N_30147,N_29545,N_29904);
nor U30148 (N_30148,N_29236,N_29252);
xnor U30149 (N_30149,N_29215,N_29711);
or U30150 (N_30150,N_29867,N_29042);
and U30151 (N_30151,N_29049,N_29958);
nand U30152 (N_30152,N_29237,N_29738);
xnor U30153 (N_30153,N_29246,N_29721);
and U30154 (N_30154,N_29910,N_29969);
nor U30155 (N_30155,N_29577,N_29652);
xor U30156 (N_30156,N_29437,N_29755);
or U30157 (N_30157,N_29595,N_29318);
nor U30158 (N_30158,N_29550,N_29366);
nand U30159 (N_30159,N_29289,N_29481);
or U30160 (N_30160,N_29776,N_29725);
or U30161 (N_30161,N_29086,N_29146);
or U30162 (N_30162,N_29355,N_29938);
xnor U30163 (N_30163,N_29871,N_29405);
nand U30164 (N_30164,N_29607,N_29833);
xor U30165 (N_30165,N_29974,N_29578);
nor U30166 (N_30166,N_29728,N_29884);
or U30167 (N_30167,N_29784,N_29617);
nand U30168 (N_30168,N_29744,N_29348);
or U30169 (N_30169,N_29012,N_29622);
or U30170 (N_30170,N_29979,N_29856);
nand U30171 (N_30171,N_29680,N_29519);
and U30172 (N_30172,N_29056,N_29118);
nand U30173 (N_30173,N_29292,N_29284);
xor U30174 (N_30174,N_29589,N_29357);
or U30175 (N_30175,N_29105,N_29917);
or U30176 (N_30176,N_29316,N_29957);
nand U30177 (N_30177,N_29407,N_29122);
nand U30178 (N_30178,N_29889,N_29663);
nor U30179 (N_30179,N_29301,N_29574);
or U30180 (N_30180,N_29832,N_29457);
nor U30181 (N_30181,N_29512,N_29712);
or U30182 (N_30182,N_29224,N_29019);
or U30183 (N_30183,N_29429,N_29314);
and U30184 (N_30184,N_29143,N_29181);
xor U30185 (N_30185,N_29089,N_29973);
nand U30186 (N_30186,N_29740,N_29517);
xnor U30187 (N_30187,N_29796,N_29278);
nand U30188 (N_30188,N_29754,N_29834);
and U30189 (N_30189,N_29003,N_29347);
or U30190 (N_30190,N_29702,N_29426);
or U30191 (N_30191,N_29971,N_29375);
nand U30192 (N_30192,N_29806,N_29651);
nand U30193 (N_30193,N_29699,N_29008);
and U30194 (N_30194,N_29018,N_29359);
nand U30195 (N_30195,N_29047,N_29532);
xor U30196 (N_30196,N_29835,N_29212);
and U30197 (N_30197,N_29854,N_29986);
or U30198 (N_30198,N_29830,N_29801);
xnor U30199 (N_30199,N_29870,N_29035);
and U30200 (N_30200,N_29593,N_29171);
nand U30201 (N_30201,N_29369,N_29178);
nor U30202 (N_30202,N_29434,N_29598);
and U30203 (N_30203,N_29920,N_29285);
nor U30204 (N_30204,N_29271,N_29394);
and U30205 (N_30205,N_29679,N_29961);
nand U30206 (N_30206,N_29956,N_29729);
xnor U30207 (N_30207,N_29513,N_29362);
nor U30208 (N_30208,N_29274,N_29586);
nor U30209 (N_30209,N_29132,N_29671);
xor U30210 (N_30210,N_29769,N_29041);
xnor U30211 (N_30211,N_29416,N_29471);
or U30212 (N_30212,N_29989,N_29912);
nand U30213 (N_30213,N_29040,N_29647);
nor U30214 (N_30214,N_29820,N_29378);
and U30215 (N_30215,N_29383,N_29539);
nor U30216 (N_30216,N_29213,N_29524);
nand U30217 (N_30217,N_29592,N_29414);
nor U30218 (N_30218,N_29780,N_29330);
or U30219 (N_30219,N_29692,N_29847);
xnor U30220 (N_30220,N_29468,N_29109);
or U30221 (N_30221,N_29332,N_29328);
xor U30222 (N_30222,N_29562,N_29564);
nor U30223 (N_30223,N_29390,N_29115);
and U30224 (N_30224,N_29011,N_29194);
xnor U30225 (N_30225,N_29777,N_29124);
and U30226 (N_30226,N_29266,N_29558);
or U30227 (N_30227,N_29014,N_29805);
and U30228 (N_30228,N_29145,N_29566);
nor U30229 (N_30229,N_29544,N_29159);
and U30230 (N_30230,N_29814,N_29783);
and U30231 (N_30231,N_29599,N_29594);
nand U30232 (N_30232,N_29472,N_29324);
nor U30233 (N_30233,N_29992,N_29428);
xor U30234 (N_30234,N_29063,N_29715);
nor U30235 (N_30235,N_29408,N_29894);
nor U30236 (N_30236,N_29960,N_29688);
nand U30237 (N_30237,N_29600,N_29393);
and U30238 (N_30238,N_29214,N_29295);
or U30239 (N_30239,N_29256,N_29313);
xnor U30240 (N_30240,N_29076,N_29624);
and U30241 (N_30241,N_29639,N_29188);
and U30242 (N_30242,N_29952,N_29682);
xor U30243 (N_30243,N_29726,N_29356);
or U30244 (N_30244,N_29420,N_29338);
nor U30245 (N_30245,N_29043,N_29070);
nor U30246 (N_30246,N_29966,N_29633);
xnor U30247 (N_30247,N_29838,N_29778);
nand U30248 (N_30248,N_29198,N_29373);
xnor U30249 (N_30249,N_29753,N_29376);
xnor U30250 (N_30250,N_29698,N_29452);
and U30251 (N_30251,N_29441,N_29916);
nor U30252 (N_30252,N_29850,N_29824);
nand U30253 (N_30253,N_29166,N_29826);
nor U30254 (N_30254,N_29281,N_29339);
and U30255 (N_30255,N_29120,N_29897);
or U30256 (N_30256,N_29501,N_29238);
and U30257 (N_30257,N_29982,N_29775);
xor U30258 (N_30258,N_29485,N_29247);
or U30259 (N_30259,N_29662,N_29793);
and U30260 (N_30260,N_29466,N_29737);
or U30261 (N_30261,N_29092,N_29944);
nand U30262 (N_30262,N_29573,N_29987);
or U30263 (N_30263,N_29529,N_29469);
and U30264 (N_30264,N_29508,N_29677);
and U30265 (N_30265,N_29064,N_29898);
nor U30266 (N_30266,N_29343,N_29187);
nand U30267 (N_30267,N_29139,N_29493);
or U30268 (N_30268,N_29949,N_29878);
nand U30269 (N_30269,N_29060,N_29800);
nand U30270 (N_30270,N_29500,N_29848);
xor U30271 (N_30271,N_29669,N_29066);
or U30272 (N_30272,N_29413,N_29749);
or U30273 (N_30273,N_29239,N_29888);
xor U30274 (N_30274,N_29415,N_29354);
and U30275 (N_30275,N_29789,N_29100);
xor U30276 (N_30276,N_29742,N_29026);
nand U30277 (N_30277,N_29827,N_29156);
nor U30278 (N_30278,N_29387,N_29668);
nor U30279 (N_30279,N_29370,N_29575);
and U30280 (N_30280,N_29309,N_29127);
nand U30281 (N_30281,N_29641,N_29205);
or U30282 (N_30282,N_29646,N_29791);
or U30283 (N_30283,N_29077,N_29708);
nor U30284 (N_30284,N_29841,N_29759);
and U30285 (N_30285,N_29621,N_29116);
xnor U30286 (N_30286,N_29150,N_29020);
nand U30287 (N_30287,N_29861,N_29653);
nand U30288 (N_30288,N_29447,N_29506);
and U30289 (N_30289,N_29352,N_29321);
or U30290 (N_30290,N_29543,N_29106);
or U30291 (N_30291,N_29817,N_29179);
or U30292 (N_30292,N_29746,N_29440);
nor U30293 (N_30293,N_29511,N_29248);
and U30294 (N_30294,N_29443,N_29102);
nor U30295 (N_30295,N_29580,N_29868);
nand U30296 (N_30296,N_29186,N_29852);
or U30297 (N_30297,N_29637,N_29804);
and U30298 (N_30298,N_29184,N_29023);
xor U30299 (N_30299,N_29264,N_29860);
nand U30300 (N_30300,N_29496,N_29602);
nor U30301 (N_30301,N_29061,N_29872);
xor U30302 (N_30302,N_29811,N_29470);
nor U30303 (N_30303,N_29091,N_29033);
or U30304 (N_30304,N_29463,N_29398);
or U30305 (N_30305,N_29918,N_29876);
nor U30306 (N_30306,N_29196,N_29346);
or U30307 (N_30307,N_29059,N_29454);
nor U30308 (N_30308,N_29044,N_29809);
xor U30309 (N_30309,N_29620,N_29164);
or U30310 (N_30310,N_29991,N_29984);
nor U30311 (N_30311,N_29821,N_29661);
xnor U30312 (N_30312,N_29467,N_29151);
nand U30313 (N_30313,N_29085,N_29036);
nand U30314 (N_30314,N_29977,N_29631);
nor U30315 (N_30315,N_29941,N_29461);
nand U30316 (N_30316,N_29030,N_29681);
nor U30317 (N_30317,N_29829,N_29189);
and U30318 (N_30318,N_29365,N_29228);
and U30319 (N_30319,N_29099,N_29766);
xor U30320 (N_30320,N_29418,N_29280);
nand U30321 (N_30321,N_29138,N_29567);
or U30322 (N_30322,N_29614,N_29027);
nor U30323 (N_30323,N_29350,N_29541);
xor U30324 (N_30324,N_29455,N_29869);
and U30325 (N_30325,N_29644,N_29895);
xnor U30326 (N_30326,N_29972,N_29836);
xor U30327 (N_30327,N_29927,N_29822);
xnor U30328 (N_30328,N_29813,N_29149);
or U30329 (N_30329,N_29696,N_29588);
nand U30330 (N_30330,N_29379,N_29074);
xor U30331 (N_30331,N_29283,N_29714);
nor U30332 (N_30332,N_29364,N_29533);
nor U30333 (N_30333,N_29942,N_29899);
or U30334 (N_30334,N_29286,N_29807);
nor U30335 (N_30335,N_29204,N_29113);
nand U30336 (N_30336,N_29068,N_29643);
and U30337 (N_30337,N_29879,N_29207);
nor U30338 (N_30338,N_29610,N_29760);
nor U30339 (N_30339,N_29703,N_29534);
and U30340 (N_30340,N_29694,N_29173);
and U30341 (N_30341,N_29865,N_29630);
nor U30342 (N_30342,N_29439,N_29678);
nor U30343 (N_30343,N_29299,N_29716);
nor U30344 (N_30344,N_29101,N_29603);
and U30345 (N_30345,N_29402,N_29734);
nor U30346 (N_30346,N_29180,N_29082);
xor U30347 (N_30347,N_29185,N_29996);
nand U30348 (N_30348,N_29475,N_29978);
and U30349 (N_30349,N_29799,N_29002);
and U30350 (N_30350,N_29169,N_29548);
or U30351 (N_30351,N_29983,N_29351);
and U30352 (N_30352,N_29518,N_29887);
xnor U30353 (N_30353,N_29923,N_29514);
or U30354 (N_30354,N_29262,N_29004);
xor U30355 (N_30355,N_29794,N_29072);
xor U30356 (N_30356,N_29774,N_29862);
and U30357 (N_30357,N_29001,N_29234);
nor U30358 (N_30358,N_29265,N_29994);
xnor U30359 (N_30359,N_29601,N_29660);
nor U30360 (N_30360,N_29240,N_29039);
or U30361 (N_30361,N_29561,N_29810);
nand U30362 (N_30362,N_29797,N_29397);
and U30363 (N_30363,N_29825,N_29371);
and U30364 (N_30364,N_29037,N_29141);
nor U30365 (N_30365,N_29302,N_29242);
xnor U30366 (N_30366,N_29412,N_29655);
nand U30367 (N_30367,N_29656,N_29231);
or U30368 (N_30368,N_29549,N_29704);
nor U30369 (N_30369,N_29131,N_29142);
or U30370 (N_30370,N_29223,N_29845);
nor U30371 (N_30371,N_29377,N_29525);
or U30372 (N_30372,N_29628,N_29476);
or U30373 (N_30373,N_29748,N_29900);
xnor U30374 (N_30374,N_29395,N_29486);
nand U30375 (N_30375,N_29675,N_29565);
nand U30376 (N_30376,N_29842,N_29226);
nor U30377 (N_30377,N_29244,N_29569);
and U30378 (N_30378,N_29659,N_29399);
and U30379 (N_30379,N_29645,N_29926);
or U30380 (N_30380,N_29590,N_29873);
nand U30381 (N_30381,N_29846,N_29787);
nand U30382 (N_30382,N_29932,N_29798);
and U30383 (N_30383,N_29909,N_29844);
nor U30384 (N_30384,N_29855,N_29016);
and U30385 (N_30385,N_29859,N_29988);
and U30386 (N_30386,N_29722,N_29864);
nor U30387 (N_30387,N_29665,N_29261);
nor U30388 (N_30388,N_29667,N_29818);
and U30389 (N_30389,N_29024,N_29516);
or U30390 (N_30390,N_29293,N_29038);
xnor U30391 (N_30391,N_29596,N_29839);
nor U30392 (N_30392,N_29478,N_29731);
and U30393 (N_30393,N_29934,N_29990);
and U30394 (N_30394,N_29816,N_29903);
xnor U30395 (N_30395,N_29556,N_29477);
and U30396 (N_30396,N_29576,N_29939);
nand U30397 (N_30397,N_29815,N_29785);
and U30398 (N_30398,N_29158,N_29382);
and U30399 (N_30399,N_29627,N_29931);
xnor U30400 (N_30400,N_29225,N_29540);
or U30401 (N_30401,N_29053,N_29304);
nor U30402 (N_30402,N_29953,N_29732);
nand U30403 (N_30403,N_29981,N_29535);
nand U30404 (N_30404,N_29672,N_29757);
nand U30405 (N_30405,N_29009,N_29464);
nand U30406 (N_30406,N_29080,N_29863);
and U30407 (N_30407,N_29254,N_29770);
and U30408 (N_30408,N_29391,N_29761);
xor U30409 (N_30409,N_29123,N_29307);
nand U30410 (N_30410,N_29277,N_29432);
nand U30411 (N_30411,N_29632,N_29717);
xor U30412 (N_30412,N_29312,N_29676);
nand U30413 (N_30413,N_29358,N_29636);
nor U30414 (N_30414,N_29409,N_29111);
xor U30415 (N_30415,N_29079,N_29709);
nand U30416 (N_30416,N_29201,N_29411);
xnor U30417 (N_30417,N_29837,N_29294);
xor U30418 (N_30418,N_29484,N_29758);
or U30419 (N_30419,N_29479,N_29587);
nand U30420 (N_30420,N_29245,N_29560);
nor U30421 (N_30421,N_29305,N_29083);
nand U30422 (N_30422,N_29140,N_29626);
xor U30423 (N_30423,N_29515,N_29929);
nor U30424 (N_30424,N_29250,N_29448);
and U30425 (N_30425,N_29057,N_29553);
or U30426 (N_30426,N_29674,N_29885);
nand U30427 (N_30427,N_29337,N_29372);
or U30428 (N_30428,N_29727,N_29269);
and U30429 (N_30429,N_29458,N_29401);
or U30430 (N_30430,N_29006,N_29298);
and U30431 (N_30431,N_29045,N_29572);
xnor U30432 (N_30432,N_29353,N_29380);
or U30433 (N_30433,N_29654,N_29202);
nor U30434 (N_30434,N_29803,N_29497);
xnor U30435 (N_30435,N_29235,N_29273);
xnor U30436 (N_30436,N_29183,N_29954);
nand U30437 (N_30437,N_29495,N_29609);
nor U30438 (N_30438,N_29538,N_29494);
nor U30439 (N_30439,N_29221,N_29253);
or U30440 (N_30440,N_29329,N_29591);
and U30441 (N_30441,N_29460,N_29875);
nor U30442 (N_30442,N_29710,N_29531);
nand U30443 (N_30443,N_29808,N_29220);
and U30444 (N_30444,N_29308,N_29673);
nor U30445 (N_30445,N_29650,N_29107);
and U30446 (N_30446,N_29763,N_29608);
nor U30447 (N_30447,N_29206,N_29528);
and U30448 (N_30448,N_29664,N_29786);
xor U30449 (N_30449,N_29450,N_29112);
nand U30450 (N_30450,N_29117,N_29963);
nand U30451 (N_30451,N_29700,N_29950);
or U30452 (N_30452,N_29341,N_29200);
and U30453 (N_30453,N_29031,N_29279);
and U30454 (N_30454,N_29249,N_29296);
and U30455 (N_30455,N_29291,N_29229);
nor U30456 (N_30456,N_29521,N_29147);
nor U30457 (N_30457,N_29449,N_29193);
xnor U30458 (N_30458,N_29155,N_29883);
xnor U30459 (N_30459,N_29933,N_29404);
nand U30460 (N_30460,N_29773,N_29488);
and U30461 (N_30461,N_29687,N_29400);
nand U30462 (N_30462,N_29349,N_29520);
nor U30463 (N_30463,N_29735,N_29217);
or U30464 (N_30464,N_29946,N_29435);
or U30465 (N_30465,N_29546,N_29487);
xnor U30466 (N_30466,N_29902,N_29126);
nor U30467 (N_30467,N_29345,N_29323);
nor U30468 (N_30468,N_29613,N_29964);
nand U30469 (N_30469,N_29940,N_29880);
or U30470 (N_30470,N_29890,N_29442);
xor U30471 (N_30471,N_29768,N_29263);
or U30472 (N_30472,N_29288,N_29170);
nand U30473 (N_30473,N_29422,N_29585);
nand U30474 (N_30474,N_29995,N_29333);
and U30475 (N_30475,N_29144,N_29410);
nand U30476 (N_30476,N_29551,N_29685);
or U30477 (N_30477,N_29695,N_29327);
xor U30478 (N_30478,N_29192,N_29491);
nor U30479 (N_30479,N_29891,N_29396);
nor U30480 (N_30480,N_29779,N_29174);
and U30481 (N_30481,N_29509,N_29552);
and U30482 (N_30482,N_29684,N_29640);
nand U30483 (N_30483,N_29055,N_29015);
and U30484 (N_30484,N_29368,N_29325);
nor U30485 (N_30485,N_29010,N_29936);
nor U30486 (N_30486,N_29095,N_29088);
or U30487 (N_30487,N_29315,N_29381);
nor U30488 (N_30488,N_29597,N_29648);
nand U30489 (N_30489,N_29444,N_29094);
nor U30490 (N_30490,N_29557,N_29537);
nor U30491 (N_30491,N_29611,N_29190);
xnor U30492 (N_30492,N_29303,N_29849);
or U30493 (N_30493,N_29157,N_29881);
and U30494 (N_30494,N_29342,N_29473);
xor U30495 (N_30495,N_29069,N_29062);
nand U30496 (N_30496,N_29707,N_29772);
xor U30497 (N_30497,N_29762,N_29474);
nor U30498 (N_30498,N_29129,N_29175);
nor U30499 (N_30499,N_29251,N_29108);
or U30500 (N_30500,N_29511,N_29551);
and U30501 (N_30501,N_29904,N_29054);
nor U30502 (N_30502,N_29479,N_29988);
or U30503 (N_30503,N_29998,N_29499);
and U30504 (N_30504,N_29845,N_29026);
and U30505 (N_30505,N_29177,N_29194);
and U30506 (N_30506,N_29751,N_29422);
nand U30507 (N_30507,N_29323,N_29895);
nand U30508 (N_30508,N_29264,N_29507);
and U30509 (N_30509,N_29601,N_29985);
or U30510 (N_30510,N_29718,N_29831);
and U30511 (N_30511,N_29546,N_29548);
and U30512 (N_30512,N_29031,N_29058);
or U30513 (N_30513,N_29546,N_29957);
or U30514 (N_30514,N_29481,N_29489);
nor U30515 (N_30515,N_29724,N_29739);
xor U30516 (N_30516,N_29584,N_29807);
or U30517 (N_30517,N_29093,N_29829);
nor U30518 (N_30518,N_29076,N_29083);
nand U30519 (N_30519,N_29170,N_29191);
and U30520 (N_30520,N_29766,N_29312);
and U30521 (N_30521,N_29126,N_29465);
xnor U30522 (N_30522,N_29093,N_29644);
nand U30523 (N_30523,N_29066,N_29940);
nor U30524 (N_30524,N_29797,N_29127);
nor U30525 (N_30525,N_29082,N_29010);
nand U30526 (N_30526,N_29652,N_29545);
nor U30527 (N_30527,N_29483,N_29947);
and U30528 (N_30528,N_29176,N_29701);
and U30529 (N_30529,N_29475,N_29191);
and U30530 (N_30530,N_29907,N_29598);
nor U30531 (N_30531,N_29321,N_29517);
xor U30532 (N_30532,N_29100,N_29256);
and U30533 (N_30533,N_29015,N_29038);
xor U30534 (N_30534,N_29112,N_29683);
and U30535 (N_30535,N_29648,N_29201);
nand U30536 (N_30536,N_29998,N_29957);
xnor U30537 (N_30537,N_29453,N_29452);
xor U30538 (N_30538,N_29690,N_29478);
and U30539 (N_30539,N_29604,N_29751);
nor U30540 (N_30540,N_29947,N_29808);
nand U30541 (N_30541,N_29146,N_29650);
or U30542 (N_30542,N_29145,N_29906);
or U30543 (N_30543,N_29794,N_29892);
nand U30544 (N_30544,N_29270,N_29719);
xor U30545 (N_30545,N_29646,N_29608);
xnor U30546 (N_30546,N_29716,N_29723);
xor U30547 (N_30547,N_29092,N_29662);
nor U30548 (N_30548,N_29854,N_29816);
xnor U30549 (N_30549,N_29590,N_29312);
nand U30550 (N_30550,N_29582,N_29353);
xor U30551 (N_30551,N_29032,N_29466);
xor U30552 (N_30552,N_29729,N_29467);
xor U30553 (N_30553,N_29039,N_29168);
xor U30554 (N_30554,N_29291,N_29347);
xor U30555 (N_30555,N_29578,N_29744);
xor U30556 (N_30556,N_29646,N_29581);
or U30557 (N_30557,N_29154,N_29873);
or U30558 (N_30558,N_29968,N_29533);
or U30559 (N_30559,N_29653,N_29583);
and U30560 (N_30560,N_29190,N_29254);
or U30561 (N_30561,N_29334,N_29153);
nor U30562 (N_30562,N_29005,N_29701);
or U30563 (N_30563,N_29824,N_29887);
xor U30564 (N_30564,N_29203,N_29525);
and U30565 (N_30565,N_29799,N_29409);
nand U30566 (N_30566,N_29528,N_29637);
nor U30567 (N_30567,N_29853,N_29540);
nand U30568 (N_30568,N_29221,N_29812);
or U30569 (N_30569,N_29656,N_29901);
and U30570 (N_30570,N_29017,N_29900);
nor U30571 (N_30571,N_29182,N_29514);
nor U30572 (N_30572,N_29965,N_29253);
nand U30573 (N_30573,N_29615,N_29541);
nand U30574 (N_30574,N_29813,N_29439);
and U30575 (N_30575,N_29889,N_29333);
nor U30576 (N_30576,N_29594,N_29870);
or U30577 (N_30577,N_29663,N_29871);
nand U30578 (N_30578,N_29463,N_29537);
and U30579 (N_30579,N_29053,N_29174);
xor U30580 (N_30580,N_29546,N_29381);
xor U30581 (N_30581,N_29071,N_29228);
or U30582 (N_30582,N_29205,N_29708);
and U30583 (N_30583,N_29201,N_29125);
nand U30584 (N_30584,N_29165,N_29740);
xnor U30585 (N_30585,N_29456,N_29722);
nand U30586 (N_30586,N_29454,N_29989);
and U30587 (N_30587,N_29692,N_29389);
and U30588 (N_30588,N_29865,N_29519);
nand U30589 (N_30589,N_29293,N_29689);
or U30590 (N_30590,N_29099,N_29320);
and U30591 (N_30591,N_29037,N_29410);
nand U30592 (N_30592,N_29796,N_29190);
nand U30593 (N_30593,N_29128,N_29478);
xor U30594 (N_30594,N_29644,N_29075);
and U30595 (N_30595,N_29563,N_29797);
xor U30596 (N_30596,N_29390,N_29262);
xnor U30597 (N_30597,N_29708,N_29255);
xor U30598 (N_30598,N_29433,N_29448);
and U30599 (N_30599,N_29424,N_29384);
or U30600 (N_30600,N_29723,N_29112);
nor U30601 (N_30601,N_29081,N_29006);
nor U30602 (N_30602,N_29386,N_29502);
xor U30603 (N_30603,N_29657,N_29827);
and U30604 (N_30604,N_29001,N_29050);
xor U30605 (N_30605,N_29833,N_29823);
or U30606 (N_30606,N_29247,N_29550);
xnor U30607 (N_30607,N_29012,N_29875);
xnor U30608 (N_30608,N_29055,N_29609);
nand U30609 (N_30609,N_29296,N_29960);
or U30610 (N_30610,N_29490,N_29008);
nor U30611 (N_30611,N_29988,N_29231);
or U30612 (N_30612,N_29720,N_29652);
xnor U30613 (N_30613,N_29215,N_29536);
and U30614 (N_30614,N_29464,N_29245);
or U30615 (N_30615,N_29343,N_29275);
xnor U30616 (N_30616,N_29592,N_29470);
nand U30617 (N_30617,N_29545,N_29601);
xor U30618 (N_30618,N_29873,N_29736);
or U30619 (N_30619,N_29388,N_29601);
nand U30620 (N_30620,N_29405,N_29991);
nand U30621 (N_30621,N_29575,N_29548);
xnor U30622 (N_30622,N_29126,N_29021);
nor U30623 (N_30623,N_29613,N_29825);
nand U30624 (N_30624,N_29165,N_29043);
nor U30625 (N_30625,N_29598,N_29027);
nor U30626 (N_30626,N_29709,N_29897);
or U30627 (N_30627,N_29617,N_29190);
or U30628 (N_30628,N_29747,N_29209);
or U30629 (N_30629,N_29526,N_29531);
or U30630 (N_30630,N_29042,N_29333);
nand U30631 (N_30631,N_29967,N_29333);
nor U30632 (N_30632,N_29700,N_29874);
nand U30633 (N_30633,N_29940,N_29155);
or U30634 (N_30634,N_29351,N_29196);
nor U30635 (N_30635,N_29877,N_29516);
xor U30636 (N_30636,N_29295,N_29243);
xor U30637 (N_30637,N_29641,N_29819);
or U30638 (N_30638,N_29006,N_29532);
nor U30639 (N_30639,N_29996,N_29512);
xnor U30640 (N_30640,N_29591,N_29653);
xnor U30641 (N_30641,N_29199,N_29147);
xnor U30642 (N_30642,N_29454,N_29406);
nand U30643 (N_30643,N_29171,N_29875);
nor U30644 (N_30644,N_29088,N_29453);
and U30645 (N_30645,N_29703,N_29652);
xnor U30646 (N_30646,N_29664,N_29862);
nand U30647 (N_30647,N_29933,N_29709);
nand U30648 (N_30648,N_29009,N_29394);
and U30649 (N_30649,N_29616,N_29035);
nand U30650 (N_30650,N_29465,N_29491);
nor U30651 (N_30651,N_29951,N_29990);
nor U30652 (N_30652,N_29377,N_29159);
and U30653 (N_30653,N_29054,N_29062);
nor U30654 (N_30654,N_29250,N_29212);
or U30655 (N_30655,N_29813,N_29756);
and U30656 (N_30656,N_29069,N_29765);
xor U30657 (N_30657,N_29953,N_29550);
nand U30658 (N_30658,N_29586,N_29105);
nand U30659 (N_30659,N_29207,N_29752);
nand U30660 (N_30660,N_29618,N_29302);
and U30661 (N_30661,N_29028,N_29201);
nor U30662 (N_30662,N_29946,N_29350);
and U30663 (N_30663,N_29753,N_29523);
or U30664 (N_30664,N_29868,N_29648);
or U30665 (N_30665,N_29676,N_29077);
xnor U30666 (N_30666,N_29124,N_29009);
nand U30667 (N_30667,N_29344,N_29234);
xor U30668 (N_30668,N_29700,N_29650);
nand U30669 (N_30669,N_29878,N_29863);
or U30670 (N_30670,N_29363,N_29792);
nand U30671 (N_30671,N_29103,N_29306);
and U30672 (N_30672,N_29063,N_29156);
and U30673 (N_30673,N_29096,N_29052);
nor U30674 (N_30674,N_29290,N_29134);
and U30675 (N_30675,N_29237,N_29618);
xnor U30676 (N_30676,N_29656,N_29314);
nand U30677 (N_30677,N_29710,N_29297);
and U30678 (N_30678,N_29519,N_29672);
nand U30679 (N_30679,N_29914,N_29880);
or U30680 (N_30680,N_29235,N_29251);
or U30681 (N_30681,N_29563,N_29306);
xor U30682 (N_30682,N_29153,N_29123);
and U30683 (N_30683,N_29931,N_29281);
xnor U30684 (N_30684,N_29768,N_29182);
nand U30685 (N_30685,N_29343,N_29045);
and U30686 (N_30686,N_29065,N_29932);
and U30687 (N_30687,N_29448,N_29505);
nor U30688 (N_30688,N_29227,N_29921);
and U30689 (N_30689,N_29881,N_29523);
and U30690 (N_30690,N_29724,N_29861);
or U30691 (N_30691,N_29836,N_29502);
nor U30692 (N_30692,N_29503,N_29012);
or U30693 (N_30693,N_29364,N_29556);
xnor U30694 (N_30694,N_29029,N_29343);
nand U30695 (N_30695,N_29613,N_29131);
nor U30696 (N_30696,N_29445,N_29959);
nand U30697 (N_30697,N_29082,N_29009);
nand U30698 (N_30698,N_29253,N_29296);
nand U30699 (N_30699,N_29700,N_29431);
and U30700 (N_30700,N_29872,N_29305);
xor U30701 (N_30701,N_29689,N_29183);
and U30702 (N_30702,N_29002,N_29591);
nand U30703 (N_30703,N_29887,N_29163);
or U30704 (N_30704,N_29436,N_29126);
and U30705 (N_30705,N_29761,N_29859);
nand U30706 (N_30706,N_29560,N_29108);
and U30707 (N_30707,N_29504,N_29992);
nand U30708 (N_30708,N_29082,N_29307);
nor U30709 (N_30709,N_29639,N_29262);
xor U30710 (N_30710,N_29423,N_29662);
and U30711 (N_30711,N_29395,N_29682);
nand U30712 (N_30712,N_29126,N_29206);
nand U30713 (N_30713,N_29083,N_29775);
xnor U30714 (N_30714,N_29237,N_29542);
xor U30715 (N_30715,N_29864,N_29672);
and U30716 (N_30716,N_29032,N_29374);
xnor U30717 (N_30717,N_29413,N_29420);
and U30718 (N_30718,N_29885,N_29364);
or U30719 (N_30719,N_29157,N_29780);
and U30720 (N_30720,N_29468,N_29215);
or U30721 (N_30721,N_29221,N_29226);
nand U30722 (N_30722,N_29674,N_29490);
xor U30723 (N_30723,N_29240,N_29996);
xor U30724 (N_30724,N_29259,N_29680);
xnor U30725 (N_30725,N_29758,N_29972);
xnor U30726 (N_30726,N_29687,N_29568);
xnor U30727 (N_30727,N_29254,N_29866);
or U30728 (N_30728,N_29850,N_29483);
xor U30729 (N_30729,N_29337,N_29672);
or U30730 (N_30730,N_29270,N_29371);
and U30731 (N_30731,N_29525,N_29354);
nand U30732 (N_30732,N_29176,N_29082);
and U30733 (N_30733,N_29725,N_29112);
xor U30734 (N_30734,N_29827,N_29539);
nor U30735 (N_30735,N_29668,N_29804);
or U30736 (N_30736,N_29705,N_29345);
and U30737 (N_30737,N_29086,N_29936);
nor U30738 (N_30738,N_29229,N_29018);
nor U30739 (N_30739,N_29430,N_29892);
xnor U30740 (N_30740,N_29270,N_29705);
or U30741 (N_30741,N_29141,N_29370);
nor U30742 (N_30742,N_29509,N_29926);
nor U30743 (N_30743,N_29918,N_29986);
or U30744 (N_30744,N_29342,N_29952);
nand U30745 (N_30745,N_29331,N_29762);
nor U30746 (N_30746,N_29458,N_29476);
or U30747 (N_30747,N_29057,N_29490);
xnor U30748 (N_30748,N_29707,N_29703);
and U30749 (N_30749,N_29028,N_29278);
xor U30750 (N_30750,N_29550,N_29138);
and U30751 (N_30751,N_29759,N_29717);
xnor U30752 (N_30752,N_29665,N_29313);
xnor U30753 (N_30753,N_29382,N_29600);
and U30754 (N_30754,N_29065,N_29714);
and U30755 (N_30755,N_29234,N_29961);
and U30756 (N_30756,N_29919,N_29546);
and U30757 (N_30757,N_29055,N_29291);
or U30758 (N_30758,N_29966,N_29888);
xnor U30759 (N_30759,N_29672,N_29952);
nor U30760 (N_30760,N_29035,N_29957);
xnor U30761 (N_30761,N_29105,N_29357);
xor U30762 (N_30762,N_29154,N_29256);
and U30763 (N_30763,N_29259,N_29520);
nor U30764 (N_30764,N_29032,N_29744);
and U30765 (N_30765,N_29354,N_29141);
nand U30766 (N_30766,N_29675,N_29161);
nand U30767 (N_30767,N_29895,N_29819);
and U30768 (N_30768,N_29552,N_29201);
xor U30769 (N_30769,N_29815,N_29704);
nand U30770 (N_30770,N_29306,N_29060);
or U30771 (N_30771,N_29805,N_29222);
and U30772 (N_30772,N_29560,N_29750);
nor U30773 (N_30773,N_29136,N_29908);
nand U30774 (N_30774,N_29673,N_29378);
nor U30775 (N_30775,N_29609,N_29700);
and U30776 (N_30776,N_29509,N_29630);
nand U30777 (N_30777,N_29992,N_29650);
xor U30778 (N_30778,N_29576,N_29681);
or U30779 (N_30779,N_29976,N_29182);
or U30780 (N_30780,N_29483,N_29274);
nand U30781 (N_30781,N_29276,N_29367);
and U30782 (N_30782,N_29967,N_29727);
nand U30783 (N_30783,N_29102,N_29681);
xnor U30784 (N_30784,N_29519,N_29536);
nor U30785 (N_30785,N_29791,N_29483);
xor U30786 (N_30786,N_29886,N_29999);
nand U30787 (N_30787,N_29326,N_29561);
and U30788 (N_30788,N_29207,N_29608);
or U30789 (N_30789,N_29748,N_29461);
or U30790 (N_30790,N_29901,N_29095);
or U30791 (N_30791,N_29040,N_29393);
or U30792 (N_30792,N_29522,N_29670);
and U30793 (N_30793,N_29034,N_29903);
xnor U30794 (N_30794,N_29763,N_29559);
nor U30795 (N_30795,N_29699,N_29737);
nand U30796 (N_30796,N_29430,N_29765);
and U30797 (N_30797,N_29932,N_29259);
and U30798 (N_30798,N_29116,N_29220);
nor U30799 (N_30799,N_29495,N_29840);
nand U30800 (N_30800,N_29032,N_29378);
xor U30801 (N_30801,N_29197,N_29723);
xnor U30802 (N_30802,N_29187,N_29426);
nand U30803 (N_30803,N_29984,N_29955);
nand U30804 (N_30804,N_29010,N_29738);
nand U30805 (N_30805,N_29167,N_29784);
nand U30806 (N_30806,N_29963,N_29745);
nor U30807 (N_30807,N_29587,N_29631);
nand U30808 (N_30808,N_29307,N_29731);
xnor U30809 (N_30809,N_29400,N_29444);
nand U30810 (N_30810,N_29163,N_29238);
nor U30811 (N_30811,N_29686,N_29012);
nor U30812 (N_30812,N_29267,N_29796);
nor U30813 (N_30813,N_29120,N_29798);
xnor U30814 (N_30814,N_29549,N_29280);
nand U30815 (N_30815,N_29303,N_29483);
or U30816 (N_30816,N_29354,N_29223);
nand U30817 (N_30817,N_29828,N_29305);
and U30818 (N_30818,N_29808,N_29702);
nor U30819 (N_30819,N_29017,N_29876);
or U30820 (N_30820,N_29939,N_29556);
nor U30821 (N_30821,N_29707,N_29869);
or U30822 (N_30822,N_29835,N_29884);
or U30823 (N_30823,N_29291,N_29001);
or U30824 (N_30824,N_29535,N_29901);
xor U30825 (N_30825,N_29209,N_29811);
nor U30826 (N_30826,N_29546,N_29315);
or U30827 (N_30827,N_29951,N_29418);
nand U30828 (N_30828,N_29176,N_29549);
and U30829 (N_30829,N_29771,N_29002);
nor U30830 (N_30830,N_29774,N_29262);
and U30831 (N_30831,N_29816,N_29118);
or U30832 (N_30832,N_29207,N_29378);
xnor U30833 (N_30833,N_29828,N_29976);
nor U30834 (N_30834,N_29146,N_29177);
or U30835 (N_30835,N_29745,N_29641);
xor U30836 (N_30836,N_29286,N_29096);
and U30837 (N_30837,N_29987,N_29484);
nand U30838 (N_30838,N_29543,N_29398);
nor U30839 (N_30839,N_29097,N_29180);
and U30840 (N_30840,N_29352,N_29377);
and U30841 (N_30841,N_29801,N_29982);
xor U30842 (N_30842,N_29424,N_29723);
and U30843 (N_30843,N_29523,N_29086);
nor U30844 (N_30844,N_29167,N_29753);
or U30845 (N_30845,N_29580,N_29442);
and U30846 (N_30846,N_29982,N_29731);
xnor U30847 (N_30847,N_29760,N_29303);
and U30848 (N_30848,N_29787,N_29411);
nor U30849 (N_30849,N_29907,N_29950);
nand U30850 (N_30850,N_29926,N_29861);
and U30851 (N_30851,N_29506,N_29642);
or U30852 (N_30852,N_29452,N_29290);
and U30853 (N_30853,N_29077,N_29555);
xnor U30854 (N_30854,N_29154,N_29916);
nand U30855 (N_30855,N_29063,N_29223);
nor U30856 (N_30856,N_29705,N_29053);
xor U30857 (N_30857,N_29272,N_29739);
xor U30858 (N_30858,N_29073,N_29209);
nor U30859 (N_30859,N_29762,N_29168);
and U30860 (N_30860,N_29724,N_29781);
and U30861 (N_30861,N_29048,N_29252);
nor U30862 (N_30862,N_29339,N_29721);
nand U30863 (N_30863,N_29790,N_29511);
nor U30864 (N_30864,N_29850,N_29544);
xnor U30865 (N_30865,N_29914,N_29665);
or U30866 (N_30866,N_29440,N_29284);
and U30867 (N_30867,N_29300,N_29007);
and U30868 (N_30868,N_29469,N_29020);
nor U30869 (N_30869,N_29338,N_29762);
nor U30870 (N_30870,N_29031,N_29677);
and U30871 (N_30871,N_29260,N_29718);
nor U30872 (N_30872,N_29296,N_29301);
xnor U30873 (N_30873,N_29497,N_29728);
xnor U30874 (N_30874,N_29338,N_29939);
nand U30875 (N_30875,N_29704,N_29244);
or U30876 (N_30876,N_29795,N_29850);
nand U30877 (N_30877,N_29207,N_29124);
nor U30878 (N_30878,N_29700,N_29361);
xnor U30879 (N_30879,N_29293,N_29452);
nand U30880 (N_30880,N_29477,N_29671);
xor U30881 (N_30881,N_29882,N_29732);
nor U30882 (N_30882,N_29732,N_29147);
and U30883 (N_30883,N_29486,N_29961);
nor U30884 (N_30884,N_29564,N_29934);
and U30885 (N_30885,N_29179,N_29134);
nor U30886 (N_30886,N_29439,N_29004);
nor U30887 (N_30887,N_29800,N_29283);
or U30888 (N_30888,N_29225,N_29452);
xnor U30889 (N_30889,N_29524,N_29897);
and U30890 (N_30890,N_29786,N_29231);
and U30891 (N_30891,N_29924,N_29326);
or U30892 (N_30892,N_29668,N_29136);
and U30893 (N_30893,N_29358,N_29073);
nand U30894 (N_30894,N_29988,N_29159);
and U30895 (N_30895,N_29154,N_29422);
and U30896 (N_30896,N_29217,N_29280);
and U30897 (N_30897,N_29815,N_29003);
or U30898 (N_30898,N_29698,N_29767);
nor U30899 (N_30899,N_29060,N_29256);
nor U30900 (N_30900,N_29161,N_29766);
nor U30901 (N_30901,N_29294,N_29770);
xnor U30902 (N_30902,N_29547,N_29356);
or U30903 (N_30903,N_29593,N_29039);
and U30904 (N_30904,N_29181,N_29735);
nand U30905 (N_30905,N_29443,N_29066);
nor U30906 (N_30906,N_29346,N_29870);
or U30907 (N_30907,N_29823,N_29520);
xnor U30908 (N_30908,N_29696,N_29402);
nand U30909 (N_30909,N_29547,N_29511);
and U30910 (N_30910,N_29530,N_29642);
nor U30911 (N_30911,N_29275,N_29873);
xor U30912 (N_30912,N_29287,N_29107);
nand U30913 (N_30913,N_29168,N_29736);
nand U30914 (N_30914,N_29822,N_29071);
xnor U30915 (N_30915,N_29967,N_29342);
xnor U30916 (N_30916,N_29056,N_29140);
and U30917 (N_30917,N_29147,N_29394);
xor U30918 (N_30918,N_29530,N_29594);
nand U30919 (N_30919,N_29205,N_29499);
nand U30920 (N_30920,N_29517,N_29273);
or U30921 (N_30921,N_29388,N_29448);
xnor U30922 (N_30922,N_29416,N_29899);
xnor U30923 (N_30923,N_29167,N_29840);
or U30924 (N_30924,N_29112,N_29166);
and U30925 (N_30925,N_29060,N_29666);
and U30926 (N_30926,N_29578,N_29018);
nand U30927 (N_30927,N_29767,N_29978);
nor U30928 (N_30928,N_29375,N_29523);
nor U30929 (N_30929,N_29302,N_29995);
nor U30930 (N_30930,N_29072,N_29068);
nor U30931 (N_30931,N_29690,N_29842);
nand U30932 (N_30932,N_29906,N_29987);
or U30933 (N_30933,N_29990,N_29340);
and U30934 (N_30934,N_29348,N_29564);
xor U30935 (N_30935,N_29918,N_29256);
or U30936 (N_30936,N_29666,N_29112);
or U30937 (N_30937,N_29826,N_29141);
xnor U30938 (N_30938,N_29526,N_29330);
or U30939 (N_30939,N_29747,N_29178);
or U30940 (N_30940,N_29073,N_29425);
xnor U30941 (N_30941,N_29665,N_29252);
and U30942 (N_30942,N_29547,N_29683);
xnor U30943 (N_30943,N_29035,N_29796);
nand U30944 (N_30944,N_29872,N_29594);
xor U30945 (N_30945,N_29164,N_29666);
and U30946 (N_30946,N_29841,N_29458);
xor U30947 (N_30947,N_29839,N_29921);
and U30948 (N_30948,N_29668,N_29722);
nor U30949 (N_30949,N_29744,N_29390);
or U30950 (N_30950,N_29718,N_29664);
or U30951 (N_30951,N_29036,N_29698);
xnor U30952 (N_30952,N_29379,N_29715);
nor U30953 (N_30953,N_29365,N_29225);
or U30954 (N_30954,N_29976,N_29985);
nand U30955 (N_30955,N_29945,N_29953);
nor U30956 (N_30956,N_29397,N_29766);
and U30957 (N_30957,N_29941,N_29352);
xnor U30958 (N_30958,N_29881,N_29573);
xor U30959 (N_30959,N_29561,N_29122);
or U30960 (N_30960,N_29700,N_29738);
xnor U30961 (N_30961,N_29469,N_29948);
or U30962 (N_30962,N_29530,N_29317);
and U30963 (N_30963,N_29702,N_29911);
and U30964 (N_30964,N_29125,N_29485);
nand U30965 (N_30965,N_29953,N_29770);
xnor U30966 (N_30966,N_29352,N_29375);
or U30967 (N_30967,N_29289,N_29926);
nand U30968 (N_30968,N_29776,N_29889);
and U30969 (N_30969,N_29873,N_29989);
and U30970 (N_30970,N_29721,N_29564);
and U30971 (N_30971,N_29420,N_29836);
xor U30972 (N_30972,N_29549,N_29354);
or U30973 (N_30973,N_29917,N_29223);
nor U30974 (N_30974,N_29796,N_29034);
nand U30975 (N_30975,N_29831,N_29916);
nor U30976 (N_30976,N_29067,N_29208);
nand U30977 (N_30977,N_29935,N_29757);
nor U30978 (N_30978,N_29963,N_29494);
xnor U30979 (N_30979,N_29557,N_29067);
xnor U30980 (N_30980,N_29250,N_29836);
xnor U30981 (N_30981,N_29846,N_29143);
nand U30982 (N_30982,N_29456,N_29036);
xor U30983 (N_30983,N_29878,N_29966);
and U30984 (N_30984,N_29179,N_29191);
xnor U30985 (N_30985,N_29104,N_29697);
nand U30986 (N_30986,N_29664,N_29060);
or U30987 (N_30987,N_29627,N_29811);
nor U30988 (N_30988,N_29029,N_29153);
and U30989 (N_30989,N_29322,N_29112);
nor U30990 (N_30990,N_29868,N_29554);
nand U30991 (N_30991,N_29816,N_29838);
and U30992 (N_30992,N_29859,N_29937);
and U30993 (N_30993,N_29069,N_29143);
or U30994 (N_30994,N_29913,N_29329);
xor U30995 (N_30995,N_29191,N_29496);
xor U30996 (N_30996,N_29918,N_29872);
nor U30997 (N_30997,N_29735,N_29463);
xor U30998 (N_30998,N_29748,N_29612);
and U30999 (N_30999,N_29208,N_29678);
or U31000 (N_31000,N_30041,N_30835);
and U31001 (N_31001,N_30534,N_30833);
nand U31002 (N_31002,N_30321,N_30425);
xor U31003 (N_31003,N_30402,N_30516);
and U31004 (N_31004,N_30865,N_30649);
or U31005 (N_31005,N_30351,N_30793);
nand U31006 (N_31006,N_30597,N_30130);
nand U31007 (N_31007,N_30613,N_30347);
or U31008 (N_31008,N_30274,N_30573);
nor U31009 (N_31009,N_30326,N_30030);
xnor U31010 (N_31010,N_30114,N_30561);
nor U31011 (N_31011,N_30890,N_30188);
nand U31012 (N_31012,N_30633,N_30583);
or U31013 (N_31013,N_30420,N_30788);
or U31014 (N_31014,N_30626,N_30636);
or U31015 (N_31015,N_30140,N_30127);
xor U31016 (N_31016,N_30875,N_30574);
nor U31017 (N_31017,N_30932,N_30846);
and U31018 (N_31018,N_30060,N_30172);
and U31019 (N_31019,N_30906,N_30553);
or U31020 (N_31020,N_30520,N_30285);
xnor U31021 (N_31021,N_30779,N_30888);
xnor U31022 (N_31022,N_30017,N_30822);
xor U31023 (N_31023,N_30388,N_30912);
xnor U31024 (N_31024,N_30809,N_30955);
or U31025 (N_31025,N_30526,N_30176);
and U31026 (N_31026,N_30338,N_30086);
nand U31027 (N_31027,N_30400,N_30264);
or U31028 (N_31028,N_30319,N_30929);
xnor U31029 (N_31029,N_30591,N_30052);
and U31030 (N_31030,N_30128,N_30480);
and U31031 (N_31031,N_30614,N_30366);
or U31032 (N_31032,N_30358,N_30839);
nand U31033 (N_31033,N_30403,N_30313);
nand U31034 (N_31034,N_30456,N_30005);
xnor U31035 (N_31035,N_30826,N_30728);
nand U31036 (N_31036,N_30872,N_30923);
nand U31037 (N_31037,N_30930,N_30717);
xnor U31038 (N_31038,N_30429,N_30075);
nor U31039 (N_31039,N_30265,N_30397);
xor U31040 (N_31040,N_30020,N_30853);
or U31041 (N_31041,N_30723,N_30604);
or U31042 (N_31042,N_30705,N_30279);
or U31043 (N_31043,N_30451,N_30972);
nor U31044 (N_31044,N_30902,N_30297);
or U31045 (N_31045,N_30161,N_30982);
nand U31046 (N_31046,N_30242,N_30071);
or U31047 (N_31047,N_30448,N_30565);
xor U31048 (N_31048,N_30744,N_30605);
nand U31049 (N_31049,N_30981,N_30523);
nand U31050 (N_31050,N_30371,N_30631);
and U31051 (N_31051,N_30382,N_30829);
or U31052 (N_31052,N_30192,N_30948);
and U31053 (N_31053,N_30707,N_30150);
or U31054 (N_31054,N_30396,N_30812);
and U31055 (N_31055,N_30083,N_30200);
or U31056 (N_31056,N_30231,N_30337);
or U31057 (N_31057,N_30891,N_30806);
nand U31058 (N_31058,N_30484,N_30349);
and U31059 (N_31059,N_30627,N_30008);
xor U31060 (N_31060,N_30327,N_30276);
xor U31061 (N_31061,N_30610,N_30792);
and U31062 (N_31062,N_30584,N_30973);
or U31063 (N_31063,N_30260,N_30203);
and U31064 (N_31064,N_30715,N_30009);
nor U31065 (N_31065,N_30594,N_30196);
and U31066 (N_31066,N_30046,N_30849);
or U31067 (N_31067,N_30765,N_30845);
and U31068 (N_31068,N_30097,N_30034);
xor U31069 (N_31069,N_30881,N_30947);
nor U31070 (N_31070,N_30813,N_30716);
xor U31071 (N_31071,N_30840,N_30921);
and U31072 (N_31072,N_30990,N_30160);
and U31073 (N_31073,N_30832,N_30299);
or U31074 (N_31074,N_30064,N_30453);
nand U31075 (N_31075,N_30886,N_30143);
and U31076 (N_31076,N_30080,N_30772);
or U31077 (N_31077,N_30378,N_30072);
nand U31078 (N_31078,N_30157,N_30039);
nand U31079 (N_31079,N_30364,N_30615);
xnor U31080 (N_31080,N_30758,N_30939);
and U31081 (N_31081,N_30712,N_30133);
nand U31082 (N_31082,N_30827,N_30010);
and U31083 (N_31083,N_30908,N_30136);
xor U31084 (N_31084,N_30748,N_30962);
nor U31085 (N_31085,N_30113,N_30243);
or U31086 (N_31086,N_30729,N_30632);
and U31087 (N_31087,N_30467,N_30894);
xnor U31088 (N_31088,N_30170,N_30089);
or U31089 (N_31089,N_30624,N_30958);
xor U31090 (N_31090,N_30205,N_30530);
and U31091 (N_31091,N_30258,N_30752);
or U31092 (N_31092,N_30213,N_30401);
or U31093 (N_31093,N_30183,N_30120);
and U31094 (N_31094,N_30013,N_30036);
or U31095 (N_31095,N_30685,N_30166);
nand U31096 (N_31096,N_30146,N_30117);
and U31097 (N_31097,N_30244,N_30411);
or U31098 (N_31098,N_30447,N_30278);
nor U31099 (N_31099,N_30029,N_30375);
nor U31100 (N_31100,N_30759,N_30771);
nor U31101 (N_31101,N_30018,N_30253);
or U31102 (N_31102,N_30836,N_30045);
nor U31103 (N_31103,N_30545,N_30619);
and U31104 (N_31104,N_30111,N_30734);
or U31105 (N_31105,N_30525,N_30303);
or U31106 (N_31106,N_30907,N_30625);
or U31107 (N_31107,N_30171,N_30206);
nand U31108 (N_31108,N_30343,N_30065);
or U31109 (N_31109,N_30595,N_30365);
and U31110 (N_31110,N_30547,N_30082);
nor U31111 (N_31111,N_30803,N_30811);
xor U31112 (N_31112,N_30404,N_30847);
or U31113 (N_31113,N_30468,N_30515);
and U31114 (N_31114,N_30441,N_30786);
nand U31115 (N_31115,N_30926,N_30164);
or U31116 (N_31116,N_30011,N_30155);
and U31117 (N_31117,N_30068,N_30897);
xor U31118 (N_31118,N_30738,N_30254);
and U31119 (N_31119,N_30061,N_30344);
nor U31120 (N_31120,N_30913,N_30693);
xnor U31121 (N_31121,N_30450,N_30147);
xor U31122 (N_31122,N_30678,N_30755);
xor U31123 (N_31123,N_30399,N_30014);
xnor U31124 (N_31124,N_30630,N_30587);
xnor U31125 (N_31125,N_30554,N_30996);
or U31126 (N_31126,N_30684,N_30848);
and U31127 (N_31127,N_30257,N_30925);
nand U31128 (N_31128,N_30575,N_30690);
nand U31129 (N_31129,N_30680,N_30866);
nor U31130 (N_31130,N_30979,N_30413);
nand U31131 (N_31131,N_30519,N_30670);
nor U31132 (N_31132,N_30514,N_30437);
nand U31133 (N_31133,N_30863,N_30556);
nand U31134 (N_31134,N_30681,N_30641);
nand U31135 (N_31135,N_30935,N_30659);
nor U31136 (N_31136,N_30392,N_30379);
nor U31137 (N_31137,N_30090,N_30645);
and U31138 (N_31138,N_30601,N_30699);
and U31139 (N_31139,N_30223,N_30198);
and U31140 (N_31140,N_30696,N_30263);
xor U31141 (N_31141,N_30126,N_30138);
nand U31142 (N_31142,N_30739,N_30362);
xnor U31143 (N_31143,N_30042,N_30747);
nand U31144 (N_31144,N_30528,N_30741);
and U31145 (N_31145,N_30828,N_30774);
and U31146 (N_31146,N_30189,N_30478);
and U31147 (N_31147,N_30533,N_30750);
and U31148 (N_31148,N_30778,N_30997);
nor U31149 (N_31149,N_30989,N_30733);
nor U31150 (N_31150,N_30799,N_30286);
nor U31151 (N_31151,N_30674,N_30977);
nor U31152 (N_31152,N_30269,N_30855);
nand U31153 (N_31153,N_30621,N_30354);
nand U31154 (N_31154,N_30336,N_30586);
nor U31155 (N_31155,N_30821,N_30050);
and U31156 (N_31156,N_30284,N_30592);
or U31157 (N_31157,N_30510,N_30654);
nand U31158 (N_31158,N_30296,N_30049);
or U31159 (N_31159,N_30145,N_30518);
nand U31160 (N_31160,N_30817,N_30187);
nor U31161 (N_31161,N_30311,N_30389);
xor U31162 (N_31162,N_30834,N_30410);
or U31163 (N_31163,N_30234,N_30230);
xor U31164 (N_31164,N_30949,N_30629);
xnor U31165 (N_31165,N_30119,N_30802);
nor U31166 (N_31166,N_30212,N_30787);
and U31167 (N_31167,N_30608,N_30668);
nor U31168 (N_31168,N_30324,N_30361);
nor U31169 (N_31169,N_30181,N_30919);
xnor U31170 (N_31170,N_30495,N_30325);
xnor U31171 (N_31171,N_30679,N_30044);
nand U31172 (N_31172,N_30353,N_30616);
nand U31173 (N_31173,N_30665,N_30452);
or U31174 (N_31174,N_30442,N_30222);
xnor U31175 (N_31175,N_30277,N_30531);
and U31176 (N_31176,N_30557,N_30314);
nor U31177 (N_31177,N_30298,N_30571);
nor U31178 (N_31178,N_30194,N_30129);
xor U31179 (N_31179,N_30386,N_30843);
nand U31180 (N_31180,N_30304,N_30537);
or U31181 (N_31181,N_30569,N_30596);
nand U31182 (N_31182,N_30905,N_30577);
or U31183 (N_31183,N_30652,N_30706);
xnor U31184 (N_31184,N_30966,N_30922);
nor U31185 (N_31185,N_30004,N_30639);
and U31186 (N_31186,N_30965,N_30995);
nor U31187 (N_31187,N_30543,N_30179);
nand U31188 (N_31188,N_30106,N_30238);
nand U31189 (N_31189,N_30944,N_30567);
nand U31190 (N_31190,N_30991,N_30988);
or U31191 (N_31191,N_30920,N_30975);
nand U31192 (N_31192,N_30439,N_30663);
or U31193 (N_31193,N_30418,N_30262);
or U31194 (N_31194,N_30945,N_30882);
and U31195 (N_31195,N_30256,N_30770);
nand U31196 (N_31196,N_30315,N_30193);
nor U31197 (N_31197,N_30391,N_30667);
nand U31198 (N_31198,N_30635,N_30491);
or U31199 (N_31199,N_30539,N_30967);
nand U31200 (N_31200,N_30927,N_30585);
nor U31201 (N_31201,N_30000,N_30310);
and U31202 (N_31202,N_30019,N_30178);
nor U31203 (N_31203,N_30012,N_30470);
nand U31204 (N_31204,N_30898,N_30640);
xor U31205 (N_31205,N_30085,N_30251);
and U31206 (N_31206,N_30938,N_30713);
nor U31207 (N_31207,N_30318,N_30186);
nor U31208 (N_31208,N_30736,N_30015);
nand U31209 (N_31209,N_30850,N_30031);
and U31210 (N_31210,N_30791,N_30762);
xor U31211 (N_31211,N_30730,N_30942);
or U31212 (N_31212,N_30182,N_30798);
nand U31213 (N_31213,N_30440,N_30214);
and U31214 (N_31214,N_30245,N_30634);
nor U31215 (N_31215,N_30721,N_30007);
xor U31216 (N_31216,N_30941,N_30499);
nor U31217 (N_31217,N_30316,N_30374);
xnor U31218 (N_31218,N_30043,N_30094);
or U31219 (N_31219,N_30151,N_30227);
nor U31220 (N_31220,N_30153,N_30454);
xor U31221 (N_31221,N_30954,N_30312);
nor U31222 (N_31222,N_30578,N_30618);
xnor U31223 (N_31223,N_30077,N_30795);
or U31224 (N_31224,N_30003,N_30204);
nor U31225 (N_31225,N_30141,N_30419);
and U31226 (N_31226,N_30661,N_30394);
or U31227 (N_31227,N_30504,N_30356);
nand U31228 (N_31228,N_30173,N_30348);
and U31229 (N_31229,N_30588,N_30651);
nor U31230 (N_31230,N_30858,N_30436);
and U31231 (N_31231,N_30956,N_30305);
or U31232 (N_31232,N_30880,N_30560);
or U31233 (N_31233,N_30497,N_30438);
or U31234 (N_31234,N_30293,N_30745);
and U31235 (N_31235,N_30078,N_30766);
nand U31236 (N_31236,N_30102,N_30682);
and U31237 (N_31237,N_30067,N_30953);
nor U31238 (N_31238,N_30423,N_30329);
nand U31239 (N_31239,N_30884,N_30564);
xnor U31240 (N_31240,N_30503,N_30540);
nor U31241 (N_31241,N_30426,N_30070);
xnor U31242 (N_31242,N_30159,N_30226);
or U31243 (N_31243,N_30820,N_30790);
and U31244 (N_31244,N_30870,N_30333);
nor U31245 (N_31245,N_30727,N_30692);
xnor U31246 (N_31246,N_30506,N_30091);
and U31247 (N_31247,N_30248,N_30058);
xor U31248 (N_31248,N_30720,N_30993);
nand U31249 (N_31249,N_30202,N_30032);
nor U31250 (N_31250,N_30725,N_30458);
or U31251 (N_31251,N_30037,N_30864);
nor U31252 (N_31252,N_30465,N_30963);
and U31253 (N_31253,N_30461,N_30658);
xnor U31254 (N_31254,N_30152,N_30675);
and U31255 (N_31255,N_30676,N_30341);
nor U31256 (N_31256,N_30580,N_30646);
xnor U31257 (N_31257,N_30856,N_30877);
nor U31258 (N_31258,N_30924,N_30191);
nand U31259 (N_31259,N_30377,N_30475);
xor U31260 (N_31260,N_30529,N_30370);
nand U31261 (N_31261,N_30550,N_30084);
nand U31262 (N_31262,N_30096,N_30271);
nor U31263 (N_31263,N_30026,N_30022);
xnor U31264 (N_31264,N_30054,N_30782);
nand U31265 (N_31265,N_30910,N_30381);
nor U31266 (N_31266,N_30757,N_30511);
or U31267 (N_31267,N_30095,N_30622);
xnor U31268 (N_31268,N_30208,N_30422);
or U31269 (N_31269,N_30224,N_30322);
or U31270 (N_31270,N_30479,N_30273);
xor U31271 (N_31271,N_30346,N_30777);
and U31272 (N_31272,N_30323,N_30968);
or U31273 (N_31273,N_30776,N_30753);
and U31274 (N_31274,N_30027,N_30309);
nor U31275 (N_31275,N_30088,N_30240);
nand U31276 (N_31276,N_30746,N_30301);
and U31277 (N_31277,N_30185,N_30548);
or U31278 (N_31278,N_30644,N_30726);
or U31279 (N_31279,N_30142,N_30637);
xor U31280 (N_31280,N_30001,N_30446);
nand U31281 (N_31281,N_30909,N_30517);
and U31282 (N_31282,N_30369,N_30066);
or U31283 (N_31283,N_30781,N_30538);
xnor U31284 (N_31284,N_30950,N_30814);
nor U31285 (N_31285,N_30959,N_30047);
and U31286 (N_31286,N_30252,N_30562);
or U31287 (N_31287,N_30883,N_30215);
or U31288 (N_31288,N_30756,N_30300);
xor U31289 (N_31289,N_30267,N_30057);
nand U31290 (N_31290,N_30098,N_30940);
nand U31291 (N_31291,N_30686,N_30104);
or U31292 (N_31292,N_30334,N_30784);
xnor U31293 (N_31293,N_30816,N_30718);
or U31294 (N_31294,N_30689,N_30474);
nor U31295 (N_31295,N_30476,N_30559);
nand U31296 (N_31296,N_30421,N_30081);
nand U31297 (N_31297,N_30546,N_30195);
and U31298 (N_31298,N_30570,N_30177);
and U31299 (N_31299,N_30342,N_30241);
and U31300 (N_31300,N_30638,N_30536);
nand U31301 (N_31301,N_30180,N_30035);
nor U31302 (N_31302,N_30357,N_30016);
and U31303 (N_31303,N_30331,N_30563);
nand U31304 (N_31304,N_30040,N_30021);
nand U31305 (N_31305,N_30598,N_30719);
nor U31306 (N_31306,N_30387,N_30308);
nor U31307 (N_31307,N_30869,N_30703);
xor U31308 (N_31308,N_30092,N_30099);
nor U31309 (N_31309,N_30783,N_30249);
and U31310 (N_31310,N_30167,N_30861);
nor U31311 (N_31311,N_30647,N_30607);
nor U31312 (N_31312,N_30210,N_30220);
or U31313 (N_31313,N_30449,N_30033);
nor U31314 (N_31314,N_30428,N_30320);
and U31315 (N_31315,N_30288,N_30289);
and U31316 (N_31316,N_30255,N_30122);
and U31317 (N_31317,N_30431,N_30576);
nand U31318 (N_31318,N_30500,N_30871);
and U31319 (N_31319,N_30443,N_30768);
and U31320 (N_31320,N_30860,N_30079);
nor U31321 (N_31321,N_30937,N_30841);
nand U31322 (N_31322,N_30487,N_30737);
nand U31323 (N_31323,N_30648,N_30144);
and U31324 (N_31324,N_30852,N_30272);
nand U31325 (N_31325,N_30568,N_30606);
nor U31326 (N_31326,N_30100,N_30581);
nand U31327 (N_31327,N_30112,N_30134);
xor U31328 (N_31328,N_30551,N_30994);
and U31329 (N_31329,N_30427,N_30281);
and U31330 (N_31330,N_30804,N_30911);
and U31331 (N_31331,N_30970,N_30800);
and U31332 (N_31332,N_30899,N_30494);
and U31333 (N_31333,N_30290,N_30496);
nor U31334 (N_31334,N_30268,N_30857);
and U31335 (N_31335,N_30282,N_30775);
nor U31336 (N_31336,N_30270,N_30350);
and U31337 (N_31337,N_30459,N_30915);
and U31338 (N_31338,N_30471,N_30724);
xor U31339 (N_31339,N_30711,N_30885);
xor U31340 (N_31340,N_30405,N_30390);
xnor U31341 (N_31341,N_30612,N_30359);
and U31342 (N_31342,N_30132,N_30190);
and U31343 (N_31343,N_30708,N_30895);
and U31344 (N_31344,N_30823,N_30876);
xnor U31345 (N_31345,N_30769,N_30261);
nor U31346 (N_31346,N_30412,N_30710);
nor U31347 (N_31347,N_30946,N_30229);
xor U31348 (N_31348,N_30507,N_30055);
or U31349 (N_31349,N_30928,N_30671);
nor U31350 (N_31350,N_30808,N_30797);
or U31351 (N_31351,N_30367,N_30743);
xnor U31352 (N_31352,N_30302,N_30677);
nand U31353 (N_31353,N_30483,N_30105);
and U31354 (N_31354,N_30666,N_30878);
nor U31355 (N_31355,N_30063,N_30056);
and U31356 (N_31356,N_30542,N_30283);
and U31357 (N_31357,N_30059,N_30662);
xor U31358 (N_31358,N_30751,N_30053);
nand U31359 (N_31359,N_30702,N_30363);
and U31360 (N_31360,N_30385,N_30493);
nor U31361 (N_31361,N_30498,N_30722);
or U31362 (N_31362,N_30051,N_30867);
or U31363 (N_31363,N_30603,N_30672);
nor U31364 (N_31364,N_30239,N_30742);
and U31365 (N_31365,N_30714,N_30512);
and U31366 (N_31366,N_30028,N_30393);
or U31367 (N_31367,N_30069,N_30424);
nor U31368 (N_31368,N_30462,N_30687);
nand U31369 (N_31369,N_30006,N_30048);
nand U31370 (N_31370,N_30532,N_30445);
nor U31371 (N_31371,N_30986,N_30232);
nand U31372 (N_31372,N_30825,N_30103);
nor U31373 (N_31373,N_30199,N_30740);
nand U31374 (N_31374,N_30628,N_30339);
nor U31375 (N_31375,N_30280,N_30754);
nor U31376 (N_31376,N_30892,N_30887);
xor U31377 (N_31377,N_30544,N_30969);
and U31378 (N_31378,N_30233,N_30934);
xor U31379 (N_31379,N_30101,N_30455);
nor U31380 (N_31380,N_30373,N_30398);
xnor U31381 (N_31381,N_30810,N_30169);
nand U31382 (N_31382,N_30785,N_30992);
xor U31383 (N_31383,N_30960,N_30156);
or U31384 (N_31384,N_30330,N_30062);
nand U31385 (N_31385,N_30815,N_30837);
or U31386 (N_31386,N_30221,N_30914);
nor U31387 (N_31387,N_30549,N_30552);
and U31388 (N_31388,N_30695,N_30216);
nand U31389 (N_31389,N_30209,N_30521);
xnor U31390 (N_31390,N_30558,N_30831);
xnor U31391 (N_31391,N_30168,N_30481);
xnor U31392 (N_31392,N_30137,N_30023);
nand U31393 (N_31393,N_30295,N_30900);
or U31394 (N_31394,N_30207,N_30780);
nor U31395 (N_31395,N_30109,N_30355);
nor U31396 (N_31396,N_30660,N_30599);
and U31397 (N_31397,N_30492,N_30961);
nand U31398 (N_31398,N_30998,N_30287);
xnor U31399 (N_31399,N_30317,N_30918);
and U31400 (N_31400,N_30175,N_30118);
nand U31401 (N_31401,N_30964,N_30896);
nand U31402 (N_31402,N_30698,N_30201);
nand U31403 (N_31403,N_30760,N_30482);
nor U31404 (N_31404,N_30236,N_30225);
nand U31405 (N_31405,N_30976,N_30688);
nand U31406 (N_31406,N_30978,N_30415);
xnor U31407 (N_31407,N_30974,N_30408);
nor U31408 (N_31408,N_30555,N_30444);
nor U31409 (N_31409,N_30859,N_30368);
xnor U31410 (N_31410,N_30228,N_30306);
and U31411 (N_31411,N_30524,N_30952);
nor U31412 (N_31412,N_30844,N_30767);
and U31413 (N_31413,N_30488,N_30076);
and U31414 (N_31414,N_30162,N_30664);
and U31415 (N_31415,N_30395,N_30824);
nor U31416 (N_31416,N_30773,N_30148);
nand U31417 (N_31417,N_30380,N_30352);
xor U31418 (N_31418,N_30197,N_30617);
and U31419 (N_31419,N_30165,N_30893);
and U31420 (N_31420,N_30149,N_30219);
xnor U31421 (N_31421,N_30259,N_30691);
or U31422 (N_31422,N_30983,N_30464);
xor U31423 (N_31423,N_30805,N_30139);
xor U31424 (N_31424,N_30217,N_30602);
and U31425 (N_31425,N_30116,N_30406);
or U31426 (N_31426,N_30211,N_30943);
nor U31427 (N_31427,N_30332,N_30435);
and U31428 (N_31428,N_30763,N_30620);
or U31429 (N_31429,N_30237,N_30527);
or U31430 (N_31430,N_30460,N_30854);
xor U31431 (N_31431,N_30246,N_30623);
nand U31432 (N_31432,N_30489,N_30345);
nor U31433 (N_31433,N_30184,N_30414);
xor U31434 (N_31434,N_30903,N_30490);
or U31435 (N_31435,N_30694,N_30294);
nand U31436 (N_31436,N_30335,N_30174);
and U31437 (N_31437,N_30879,N_30818);
nor U31438 (N_31438,N_30582,N_30761);
xnor U31439 (N_31439,N_30472,N_30291);
and U31440 (N_31440,N_30384,N_30505);
or U31441 (N_31441,N_30541,N_30794);
and U31442 (N_31442,N_30074,N_30700);
or U31443 (N_31443,N_30110,N_30469);
xnor U31444 (N_31444,N_30509,N_30764);
xnor U31445 (N_31445,N_30247,N_30121);
or U31446 (N_31446,N_30002,N_30951);
xor U31447 (N_31447,N_30838,N_30579);
and U31448 (N_31448,N_30124,N_30466);
nor U31449 (N_31449,N_30789,N_30038);
and U31450 (N_31450,N_30154,N_30611);
nor U31451 (N_31451,N_30340,N_30501);
xnor U31452 (N_31452,N_30407,N_30731);
or U31453 (N_31453,N_30709,N_30508);
xnor U31454 (N_31454,N_30590,N_30250);
nand U31455 (N_31455,N_30643,N_30916);
and U31456 (N_31456,N_30372,N_30486);
nor U31457 (N_31457,N_30999,N_30673);
nand U31458 (N_31458,N_30819,N_30093);
or U31459 (N_31459,N_30656,N_30980);
xor U31460 (N_31460,N_30901,N_30704);
xnor U31461 (N_31461,N_30125,N_30383);
or U31462 (N_31462,N_30697,N_30936);
xor U31463 (N_31463,N_30107,N_30522);
nor U31464 (N_31464,N_30158,N_30433);
nand U31465 (N_31465,N_30931,N_30430);
xor U31466 (N_31466,N_30434,N_30328);
and U31467 (N_31467,N_30796,N_30108);
nand U31468 (N_31468,N_30123,N_30485);
and U31469 (N_31469,N_30873,N_30463);
or U31470 (N_31470,N_30701,N_30749);
or U31471 (N_31471,N_30566,N_30409);
and U31472 (N_31472,N_30417,N_30874);
xnor U31473 (N_31473,N_30657,N_30732);
and U31474 (N_31474,N_30917,N_30513);
xnor U31475 (N_31475,N_30457,N_30642);
and U31476 (N_31476,N_30163,N_30218);
xor U31477 (N_31477,N_30376,N_30024);
and U31478 (N_31478,N_30131,N_30985);
nand U31479 (N_31479,N_30987,N_30572);
xnor U31480 (N_31480,N_30653,N_30984);
and U31481 (N_31481,N_30589,N_30235);
or U31482 (N_31482,N_30266,N_30868);
and U31483 (N_31483,N_30933,N_30957);
and U31484 (N_31484,N_30416,N_30655);
nor U31485 (N_31485,N_30432,N_30593);
nor U31486 (N_31486,N_30862,N_30683);
or U31487 (N_31487,N_30477,N_30473);
nand U31488 (N_31488,N_30135,N_30842);
xnor U31489 (N_31489,N_30535,N_30115);
xnor U31490 (N_31490,N_30830,N_30851);
nor U31491 (N_31491,N_30889,N_30807);
nand U31492 (N_31492,N_30600,N_30307);
and U31493 (N_31493,N_30502,N_30609);
xor U31494 (N_31494,N_30025,N_30801);
or U31495 (N_31495,N_30087,N_30275);
nor U31496 (N_31496,N_30360,N_30073);
nor U31497 (N_31497,N_30904,N_30971);
nor U31498 (N_31498,N_30650,N_30735);
and U31499 (N_31499,N_30292,N_30669);
nor U31500 (N_31500,N_30239,N_30209);
nor U31501 (N_31501,N_30180,N_30646);
nand U31502 (N_31502,N_30229,N_30844);
nor U31503 (N_31503,N_30312,N_30902);
xor U31504 (N_31504,N_30747,N_30551);
or U31505 (N_31505,N_30261,N_30999);
xor U31506 (N_31506,N_30166,N_30044);
and U31507 (N_31507,N_30220,N_30238);
and U31508 (N_31508,N_30756,N_30587);
nor U31509 (N_31509,N_30668,N_30020);
nor U31510 (N_31510,N_30881,N_30894);
and U31511 (N_31511,N_30098,N_30301);
and U31512 (N_31512,N_30625,N_30956);
or U31513 (N_31513,N_30225,N_30478);
xnor U31514 (N_31514,N_30178,N_30516);
nor U31515 (N_31515,N_30112,N_30072);
or U31516 (N_31516,N_30595,N_30633);
xnor U31517 (N_31517,N_30750,N_30703);
nand U31518 (N_31518,N_30690,N_30199);
nor U31519 (N_31519,N_30735,N_30371);
or U31520 (N_31520,N_30348,N_30996);
or U31521 (N_31521,N_30929,N_30893);
and U31522 (N_31522,N_30845,N_30511);
and U31523 (N_31523,N_30274,N_30272);
xor U31524 (N_31524,N_30452,N_30299);
xnor U31525 (N_31525,N_30242,N_30222);
nor U31526 (N_31526,N_30196,N_30874);
nand U31527 (N_31527,N_30112,N_30532);
and U31528 (N_31528,N_30095,N_30311);
and U31529 (N_31529,N_30300,N_30601);
xor U31530 (N_31530,N_30263,N_30887);
nor U31531 (N_31531,N_30785,N_30540);
xnor U31532 (N_31532,N_30440,N_30236);
or U31533 (N_31533,N_30031,N_30468);
or U31534 (N_31534,N_30568,N_30404);
nor U31535 (N_31535,N_30622,N_30769);
and U31536 (N_31536,N_30943,N_30454);
nor U31537 (N_31537,N_30787,N_30591);
and U31538 (N_31538,N_30719,N_30128);
nor U31539 (N_31539,N_30793,N_30872);
xnor U31540 (N_31540,N_30767,N_30253);
or U31541 (N_31541,N_30607,N_30114);
and U31542 (N_31542,N_30288,N_30933);
xor U31543 (N_31543,N_30968,N_30076);
xor U31544 (N_31544,N_30583,N_30162);
or U31545 (N_31545,N_30603,N_30835);
or U31546 (N_31546,N_30485,N_30586);
xnor U31547 (N_31547,N_30358,N_30641);
nand U31548 (N_31548,N_30071,N_30066);
and U31549 (N_31549,N_30145,N_30372);
nand U31550 (N_31550,N_30514,N_30922);
xor U31551 (N_31551,N_30418,N_30861);
or U31552 (N_31552,N_30716,N_30573);
nor U31553 (N_31553,N_30546,N_30132);
and U31554 (N_31554,N_30537,N_30820);
xnor U31555 (N_31555,N_30153,N_30107);
or U31556 (N_31556,N_30641,N_30412);
nand U31557 (N_31557,N_30161,N_30780);
and U31558 (N_31558,N_30159,N_30057);
and U31559 (N_31559,N_30864,N_30839);
nand U31560 (N_31560,N_30081,N_30199);
xnor U31561 (N_31561,N_30030,N_30958);
or U31562 (N_31562,N_30501,N_30474);
and U31563 (N_31563,N_30246,N_30746);
nor U31564 (N_31564,N_30942,N_30983);
and U31565 (N_31565,N_30188,N_30709);
nor U31566 (N_31566,N_30034,N_30642);
nand U31567 (N_31567,N_30386,N_30115);
or U31568 (N_31568,N_30195,N_30191);
nand U31569 (N_31569,N_30028,N_30372);
nand U31570 (N_31570,N_30976,N_30761);
nor U31571 (N_31571,N_30524,N_30651);
or U31572 (N_31572,N_30963,N_30617);
nor U31573 (N_31573,N_30617,N_30109);
nor U31574 (N_31574,N_30590,N_30550);
nor U31575 (N_31575,N_30349,N_30961);
or U31576 (N_31576,N_30747,N_30408);
nand U31577 (N_31577,N_30522,N_30601);
nand U31578 (N_31578,N_30063,N_30183);
xnor U31579 (N_31579,N_30060,N_30173);
or U31580 (N_31580,N_30961,N_30019);
nor U31581 (N_31581,N_30574,N_30525);
and U31582 (N_31582,N_30085,N_30545);
xnor U31583 (N_31583,N_30297,N_30977);
nand U31584 (N_31584,N_30165,N_30021);
or U31585 (N_31585,N_30981,N_30618);
nor U31586 (N_31586,N_30764,N_30820);
nor U31587 (N_31587,N_30730,N_30547);
xor U31588 (N_31588,N_30717,N_30072);
xnor U31589 (N_31589,N_30721,N_30388);
or U31590 (N_31590,N_30853,N_30474);
nor U31591 (N_31591,N_30813,N_30826);
and U31592 (N_31592,N_30731,N_30072);
nor U31593 (N_31593,N_30405,N_30091);
xor U31594 (N_31594,N_30477,N_30077);
nor U31595 (N_31595,N_30856,N_30272);
and U31596 (N_31596,N_30202,N_30088);
nand U31597 (N_31597,N_30612,N_30278);
nor U31598 (N_31598,N_30583,N_30593);
nor U31599 (N_31599,N_30784,N_30881);
or U31600 (N_31600,N_30476,N_30919);
and U31601 (N_31601,N_30151,N_30153);
xnor U31602 (N_31602,N_30960,N_30127);
and U31603 (N_31603,N_30759,N_30342);
xor U31604 (N_31604,N_30671,N_30444);
xnor U31605 (N_31605,N_30651,N_30846);
and U31606 (N_31606,N_30432,N_30210);
xor U31607 (N_31607,N_30026,N_30501);
or U31608 (N_31608,N_30334,N_30775);
and U31609 (N_31609,N_30966,N_30133);
or U31610 (N_31610,N_30344,N_30723);
xor U31611 (N_31611,N_30305,N_30701);
xor U31612 (N_31612,N_30759,N_30787);
and U31613 (N_31613,N_30969,N_30600);
nand U31614 (N_31614,N_30703,N_30575);
and U31615 (N_31615,N_30173,N_30466);
xor U31616 (N_31616,N_30239,N_30998);
xnor U31617 (N_31617,N_30419,N_30600);
nand U31618 (N_31618,N_30616,N_30659);
nor U31619 (N_31619,N_30499,N_30101);
or U31620 (N_31620,N_30057,N_30918);
nor U31621 (N_31621,N_30847,N_30987);
nor U31622 (N_31622,N_30815,N_30816);
xnor U31623 (N_31623,N_30339,N_30704);
and U31624 (N_31624,N_30526,N_30214);
and U31625 (N_31625,N_30265,N_30622);
xor U31626 (N_31626,N_30883,N_30515);
xor U31627 (N_31627,N_30493,N_30343);
and U31628 (N_31628,N_30252,N_30105);
xnor U31629 (N_31629,N_30459,N_30181);
or U31630 (N_31630,N_30466,N_30534);
nor U31631 (N_31631,N_30275,N_30892);
or U31632 (N_31632,N_30860,N_30065);
nor U31633 (N_31633,N_30297,N_30464);
nand U31634 (N_31634,N_30932,N_30237);
or U31635 (N_31635,N_30572,N_30396);
nand U31636 (N_31636,N_30885,N_30880);
nor U31637 (N_31637,N_30881,N_30096);
xnor U31638 (N_31638,N_30633,N_30791);
nand U31639 (N_31639,N_30099,N_30465);
and U31640 (N_31640,N_30971,N_30110);
nand U31641 (N_31641,N_30853,N_30437);
or U31642 (N_31642,N_30514,N_30586);
xnor U31643 (N_31643,N_30934,N_30814);
nor U31644 (N_31644,N_30606,N_30540);
nand U31645 (N_31645,N_30244,N_30084);
and U31646 (N_31646,N_30690,N_30842);
xnor U31647 (N_31647,N_30852,N_30949);
and U31648 (N_31648,N_30035,N_30692);
or U31649 (N_31649,N_30104,N_30316);
nor U31650 (N_31650,N_30132,N_30900);
or U31651 (N_31651,N_30850,N_30161);
or U31652 (N_31652,N_30549,N_30389);
xor U31653 (N_31653,N_30394,N_30430);
nand U31654 (N_31654,N_30806,N_30002);
or U31655 (N_31655,N_30324,N_30283);
or U31656 (N_31656,N_30022,N_30124);
nor U31657 (N_31657,N_30056,N_30652);
and U31658 (N_31658,N_30293,N_30287);
and U31659 (N_31659,N_30553,N_30613);
nor U31660 (N_31660,N_30466,N_30778);
xnor U31661 (N_31661,N_30952,N_30884);
nand U31662 (N_31662,N_30749,N_30723);
or U31663 (N_31663,N_30570,N_30094);
nor U31664 (N_31664,N_30316,N_30973);
xor U31665 (N_31665,N_30122,N_30439);
or U31666 (N_31666,N_30924,N_30703);
nand U31667 (N_31667,N_30046,N_30043);
and U31668 (N_31668,N_30311,N_30149);
nand U31669 (N_31669,N_30528,N_30037);
nand U31670 (N_31670,N_30144,N_30199);
nand U31671 (N_31671,N_30467,N_30045);
nand U31672 (N_31672,N_30763,N_30523);
and U31673 (N_31673,N_30551,N_30252);
or U31674 (N_31674,N_30880,N_30210);
nand U31675 (N_31675,N_30286,N_30644);
or U31676 (N_31676,N_30152,N_30954);
xnor U31677 (N_31677,N_30917,N_30126);
nor U31678 (N_31678,N_30643,N_30988);
and U31679 (N_31679,N_30401,N_30001);
xor U31680 (N_31680,N_30555,N_30512);
nand U31681 (N_31681,N_30311,N_30336);
nor U31682 (N_31682,N_30723,N_30178);
or U31683 (N_31683,N_30344,N_30816);
xnor U31684 (N_31684,N_30258,N_30953);
or U31685 (N_31685,N_30628,N_30277);
or U31686 (N_31686,N_30272,N_30443);
xor U31687 (N_31687,N_30791,N_30458);
nor U31688 (N_31688,N_30676,N_30107);
and U31689 (N_31689,N_30500,N_30574);
nor U31690 (N_31690,N_30465,N_30948);
xor U31691 (N_31691,N_30170,N_30909);
nor U31692 (N_31692,N_30952,N_30821);
xor U31693 (N_31693,N_30886,N_30082);
nor U31694 (N_31694,N_30350,N_30465);
nand U31695 (N_31695,N_30522,N_30566);
and U31696 (N_31696,N_30681,N_30905);
and U31697 (N_31697,N_30291,N_30953);
nor U31698 (N_31698,N_30588,N_30620);
xor U31699 (N_31699,N_30826,N_30162);
xor U31700 (N_31700,N_30401,N_30610);
xor U31701 (N_31701,N_30614,N_30862);
nand U31702 (N_31702,N_30819,N_30994);
and U31703 (N_31703,N_30321,N_30332);
nor U31704 (N_31704,N_30170,N_30640);
xor U31705 (N_31705,N_30156,N_30341);
nor U31706 (N_31706,N_30032,N_30913);
or U31707 (N_31707,N_30583,N_30032);
and U31708 (N_31708,N_30049,N_30294);
nor U31709 (N_31709,N_30980,N_30962);
nor U31710 (N_31710,N_30056,N_30060);
xor U31711 (N_31711,N_30355,N_30155);
or U31712 (N_31712,N_30276,N_30795);
and U31713 (N_31713,N_30265,N_30608);
nand U31714 (N_31714,N_30156,N_30775);
nand U31715 (N_31715,N_30564,N_30451);
or U31716 (N_31716,N_30379,N_30300);
nand U31717 (N_31717,N_30126,N_30732);
xor U31718 (N_31718,N_30330,N_30507);
or U31719 (N_31719,N_30995,N_30797);
nand U31720 (N_31720,N_30977,N_30012);
nand U31721 (N_31721,N_30355,N_30694);
nor U31722 (N_31722,N_30866,N_30101);
and U31723 (N_31723,N_30578,N_30462);
and U31724 (N_31724,N_30683,N_30993);
nand U31725 (N_31725,N_30438,N_30062);
xnor U31726 (N_31726,N_30433,N_30384);
or U31727 (N_31727,N_30402,N_30378);
xor U31728 (N_31728,N_30842,N_30523);
or U31729 (N_31729,N_30994,N_30645);
and U31730 (N_31730,N_30274,N_30974);
and U31731 (N_31731,N_30351,N_30520);
and U31732 (N_31732,N_30153,N_30161);
or U31733 (N_31733,N_30917,N_30056);
and U31734 (N_31734,N_30338,N_30528);
and U31735 (N_31735,N_30416,N_30304);
or U31736 (N_31736,N_30587,N_30320);
or U31737 (N_31737,N_30124,N_30074);
nand U31738 (N_31738,N_30468,N_30308);
or U31739 (N_31739,N_30052,N_30764);
nor U31740 (N_31740,N_30419,N_30692);
and U31741 (N_31741,N_30392,N_30929);
or U31742 (N_31742,N_30858,N_30760);
and U31743 (N_31743,N_30971,N_30441);
or U31744 (N_31744,N_30979,N_30626);
and U31745 (N_31745,N_30530,N_30871);
and U31746 (N_31746,N_30019,N_30293);
or U31747 (N_31747,N_30274,N_30572);
nand U31748 (N_31748,N_30725,N_30960);
xnor U31749 (N_31749,N_30605,N_30772);
or U31750 (N_31750,N_30024,N_30759);
nor U31751 (N_31751,N_30975,N_30364);
nor U31752 (N_31752,N_30124,N_30587);
nand U31753 (N_31753,N_30943,N_30792);
or U31754 (N_31754,N_30454,N_30251);
xnor U31755 (N_31755,N_30460,N_30937);
nor U31756 (N_31756,N_30211,N_30656);
xnor U31757 (N_31757,N_30605,N_30756);
and U31758 (N_31758,N_30563,N_30062);
xor U31759 (N_31759,N_30225,N_30128);
and U31760 (N_31760,N_30687,N_30409);
nand U31761 (N_31761,N_30956,N_30543);
or U31762 (N_31762,N_30250,N_30628);
nand U31763 (N_31763,N_30445,N_30987);
nor U31764 (N_31764,N_30706,N_30734);
xnor U31765 (N_31765,N_30801,N_30883);
and U31766 (N_31766,N_30900,N_30542);
nand U31767 (N_31767,N_30182,N_30721);
and U31768 (N_31768,N_30453,N_30172);
nor U31769 (N_31769,N_30265,N_30858);
nand U31770 (N_31770,N_30683,N_30424);
nand U31771 (N_31771,N_30342,N_30405);
or U31772 (N_31772,N_30280,N_30885);
nand U31773 (N_31773,N_30842,N_30206);
nand U31774 (N_31774,N_30971,N_30895);
nor U31775 (N_31775,N_30717,N_30236);
nand U31776 (N_31776,N_30198,N_30293);
nor U31777 (N_31777,N_30951,N_30518);
nand U31778 (N_31778,N_30379,N_30080);
nor U31779 (N_31779,N_30360,N_30852);
nor U31780 (N_31780,N_30574,N_30932);
nor U31781 (N_31781,N_30968,N_30617);
and U31782 (N_31782,N_30704,N_30608);
xor U31783 (N_31783,N_30783,N_30729);
xnor U31784 (N_31784,N_30406,N_30732);
nand U31785 (N_31785,N_30545,N_30380);
or U31786 (N_31786,N_30196,N_30974);
nand U31787 (N_31787,N_30500,N_30266);
nand U31788 (N_31788,N_30034,N_30937);
nor U31789 (N_31789,N_30674,N_30009);
and U31790 (N_31790,N_30124,N_30160);
xor U31791 (N_31791,N_30299,N_30838);
nand U31792 (N_31792,N_30752,N_30964);
nand U31793 (N_31793,N_30476,N_30802);
or U31794 (N_31794,N_30309,N_30467);
xnor U31795 (N_31795,N_30730,N_30921);
xnor U31796 (N_31796,N_30364,N_30818);
and U31797 (N_31797,N_30136,N_30239);
and U31798 (N_31798,N_30114,N_30699);
nand U31799 (N_31799,N_30327,N_30945);
nand U31800 (N_31800,N_30405,N_30176);
or U31801 (N_31801,N_30138,N_30035);
or U31802 (N_31802,N_30400,N_30988);
nand U31803 (N_31803,N_30222,N_30354);
nand U31804 (N_31804,N_30709,N_30211);
nand U31805 (N_31805,N_30325,N_30413);
xor U31806 (N_31806,N_30191,N_30021);
and U31807 (N_31807,N_30504,N_30704);
and U31808 (N_31808,N_30824,N_30896);
or U31809 (N_31809,N_30554,N_30838);
nand U31810 (N_31810,N_30648,N_30914);
nand U31811 (N_31811,N_30911,N_30318);
nand U31812 (N_31812,N_30626,N_30596);
nor U31813 (N_31813,N_30324,N_30695);
nand U31814 (N_31814,N_30429,N_30143);
or U31815 (N_31815,N_30969,N_30492);
nand U31816 (N_31816,N_30232,N_30565);
nand U31817 (N_31817,N_30387,N_30104);
or U31818 (N_31818,N_30646,N_30016);
nand U31819 (N_31819,N_30627,N_30943);
or U31820 (N_31820,N_30670,N_30711);
nand U31821 (N_31821,N_30841,N_30159);
and U31822 (N_31822,N_30688,N_30336);
nand U31823 (N_31823,N_30246,N_30052);
or U31824 (N_31824,N_30562,N_30331);
nor U31825 (N_31825,N_30674,N_30288);
and U31826 (N_31826,N_30649,N_30291);
and U31827 (N_31827,N_30332,N_30991);
and U31828 (N_31828,N_30675,N_30206);
nand U31829 (N_31829,N_30270,N_30536);
nor U31830 (N_31830,N_30921,N_30051);
or U31831 (N_31831,N_30958,N_30303);
nand U31832 (N_31832,N_30874,N_30552);
nor U31833 (N_31833,N_30152,N_30736);
or U31834 (N_31834,N_30181,N_30315);
nor U31835 (N_31835,N_30851,N_30490);
nor U31836 (N_31836,N_30208,N_30412);
nor U31837 (N_31837,N_30661,N_30751);
nor U31838 (N_31838,N_30269,N_30456);
xnor U31839 (N_31839,N_30527,N_30714);
or U31840 (N_31840,N_30940,N_30900);
nand U31841 (N_31841,N_30878,N_30248);
and U31842 (N_31842,N_30594,N_30134);
or U31843 (N_31843,N_30151,N_30609);
nor U31844 (N_31844,N_30365,N_30443);
nor U31845 (N_31845,N_30861,N_30120);
nor U31846 (N_31846,N_30216,N_30174);
or U31847 (N_31847,N_30774,N_30102);
nand U31848 (N_31848,N_30508,N_30813);
nand U31849 (N_31849,N_30888,N_30477);
nor U31850 (N_31850,N_30568,N_30378);
and U31851 (N_31851,N_30717,N_30803);
or U31852 (N_31852,N_30261,N_30869);
and U31853 (N_31853,N_30985,N_30027);
or U31854 (N_31854,N_30091,N_30186);
xnor U31855 (N_31855,N_30175,N_30416);
and U31856 (N_31856,N_30022,N_30013);
or U31857 (N_31857,N_30311,N_30928);
nand U31858 (N_31858,N_30085,N_30039);
xnor U31859 (N_31859,N_30267,N_30977);
xor U31860 (N_31860,N_30230,N_30072);
and U31861 (N_31861,N_30276,N_30671);
nand U31862 (N_31862,N_30993,N_30724);
nor U31863 (N_31863,N_30885,N_30962);
and U31864 (N_31864,N_30722,N_30520);
and U31865 (N_31865,N_30236,N_30704);
nor U31866 (N_31866,N_30329,N_30866);
nand U31867 (N_31867,N_30162,N_30832);
nor U31868 (N_31868,N_30981,N_30875);
and U31869 (N_31869,N_30750,N_30717);
nand U31870 (N_31870,N_30680,N_30474);
xor U31871 (N_31871,N_30954,N_30989);
xnor U31872 (N_31872,N_30142,N_30566);
and U31873 (N_31873,N_30415,N_30158);
nor U31874 (N_31874,N_30492,N_30433);
and U31875 (N_31875,N_30876,N_30127);
nand U31876 (N_31876,N_30030,N_30050);
and U31877 (N_31877,N_30893,N_30453);
and U31878 (N_31878,N_30145,N_30982);
and U31879 (N_31879,N_30816,N_30918);
or U31880 (N_31880,N_30505,N_30302);
nor U31881 (N_31881,N_30676,N_30914);
nand U31882 (N_31882,N_30981,N_30358);
nand U31883 (N_31883,N_30273,N_30931);
and U31884 (N_31884,N_30986,N_30096);
xnor U31885 (N_31885,N_30833,N_30425);
nand U31886 (N_31886,N_30827,N_30088);
and U31887 (N_31887,N_30103,N_30795);
nor U31888 (N_31888,N_30238,N_30039);
xor U31889 (N_31889,N_30713,N_30542);
nor U31890 (N_31890,N_30165,N_30133);
and U31891 (N_31891,N_30822,N_30021);
and U31892 (N_31892,N_30234,N_30472);
nand U31893 (N_31893,N_30516,N_30446);
xor U31894 (N_31894,N_30765,N_30799);
nand U31895 (N_31895,N_30023,N_30354);
nor U31896 (N_31896,N_30663,N_30067);
nor U31897 (N_31897,N_30147,N_30018);
and U31898 (N_31898,N_30272,N_30034);
and U31899 (N_31899,N_30937,N_30531);
and U31900 (N_31900,N_30279,N_30111);
or U31901 (N_31901,N_30645,N_30244);
xor U31902 (N_31902,N_30949,N_30642);
xnor U31903 (N_31903,N_30752,N_30154);
xor U31904 (N_31904,N_30657,N_30007);
nor U31905 (N_31905,N_30686,N_30308);
nor U31906 (N_31906,N_30274,N_30835);
xnor U31907 (N_31907,N_30786,N_30105);
nand U31908 (N_31908,N_30518,N_30650);
or U31909 (N_31909,N_30768,N_30737);
nor U31910 (N_31910,N_30271,N_30147);
nor U31911 (N_31911,N_30399,N_30940);
xnor U31912 (N_31912,N_30147,N_30998);
nor U31913 (N_31913,N_30628,N_30321);
nand U31914 (N_31914,N_30743,N_30423);
and U31915 (N_31915,N_30895,N_30436);
and U31916 (N_31916,N_30403,N_30962);
nand U31917 (N_31917,N_30501,N_30419);
xor U31918 (N_31918,N_30061,N_30871);
nand U31919 (N_31919,N_30727,N_30444);
xnor U31920 (N_31920,N_30889,N_30070);
or U31921 (N_31921,N_30039,N_30059);
nor U31922 (N_31922,N_30831,N_30921);
and U31923 (N_31923,N_30047,N_30434);
nor U31924 (N_31924,N_30196,N_30835);
or U31925 (N_31925,N_30966,N_30231);
or U31926 (N_31926,N_30214,N_30815);
or U31927 (N_31927,N_30568,N_30428);
nand U31928 (N_31928,N_30591,N_30980);
xor U31929 (N_31929,N_30306,N_30753);
or U31930 (N_31930,N_30950,N_30441);
xor U31931 (N_31931,N_30221,N_30391);
nor U31932 (N_31932,N_30612,N_30543);
xor U31933 (N_31933,N_30425,N_30408);
nor U31934 (N_31934,N_30858,N_30068);
xnor U31935 (N_31935,N_30438,N_30372);
or U31936 (N_31936,N_30414,N_30987);
nand U31937 (N_31937,N_30537,N_30159);
nand U31938 (N_31938,N_30564,N_30056);
xor U31939 (N_31939,N_30002,N_30802);
nand U31940 (N_31940,N_30365,N_30700);
xnor U31941 (N_31941,N_30331,N_30636);
nand U31942 (N_31942,N_30320,N_30743);
or U31943 (N_31943,N_30428,N_30397);
xor U31944 (N_31944,N_30752,N_30669);
or U31945 (N_31945,N_30185,N_30516);
nand U31946 (N_31946,N_30860,N_30746);
nor U31947 (N_31947,N_30776,N_30677);
nand U31948 (N_31948,N_30320,N_30381);
xor U31949 (N_31949,N_30296,N_30982);
xor U31950 (N_31950,N_30991,N_30100);
xor U31951 (N_31951,N_30929,N_30846);
or U31952 (N_31952,N_30828,N_30740);
nor U31953 (N_31953,N_30172,N_30522);
nand U31954 (N_31954,N_30516,N_30801);
nor U31955 (N_31955,N_30304,N_30013);
or U31956 (N_31956,N_30447,N_30402);
nand U31957 (N_31957,N_30990,N_30521);
xor U31958 (N_31958,N_30737,N_30228);
or U31959 (N_31959,N_30584,N_30164);
or U31960 (N_31960,N_30904,N_30947);
or U31961 (N_31961,N_30066,N_30476);
nand U31962 (N_31962,N_30271,N_30912);
and U31963 (N_31963,N_30268,N_30415);
or U31964 (N_31964,N_30396,N_30076);
nand U31965 (N_31965,N_30283,N_30284);
nor U31966 (N_31966,N_30444,N_30959);
or U31967 (N_31967,N_30800,N_30460);
xor U31968 (N_31968,N_30136,N_30630);
nor U31969 (N_31969,N_30938,N_30297);
nor U31970 (N_31970,N_30527,N_30764);
nand U31971 (N_31971,N_30763,N_30402);
xor U31972 (N_31972,N_30178,N_30598);
nand U31973 (N_31973,N_30753,N_30923);
xor U31974 (N_31974,N_30614,N_30761);
or U31975 (N_31975,N_30710,N_30399);
nand U31976 (N_31976,N_30674,N_30866);
xor U31977 (N_31977,N_30246,N_30810);
or U31978 (N_31978,N_30679,N_30004);
or U31979 (N_31979,N_30345,N_30226);
and U31980 (N_31980,N_30421,N_30211);
nor U31981 (N_31981,N_30921,N_30013);
or U31982 (N_31982,N_30051,N_30125);
xnor U31983 (N_31983,N_30948,N_30448);
xnor U31984 (N_31984,N_30263,N_30908);
xnor U31985 (N_31985,N_30971,N_30729);
nand U31986 (N_31986,N_30017,N_30211);
or U31987 (N_31987,N_30901,N_30978);
nor U31988 (N_31988,N_30279,N_30059);
and U31989 (N_31989,N_30261,N_30448);
xnor U31990 (N_31990,N_30923,N_30551);
nand U31991 (N_31991,N_30515,N_30849);
nor U31992 (N_31992,N_30101,N_30131);
nor U31993 (N_31993,N_30335,N_30005);
nand U31994 (N_31994,N_30243,N_30152);
nor U31995 (N_31995,N_30953,N_30723);
nand U31996 (N_31996,N_30421,N_30382);
nor U31997 (N_31997,N_30947,N_30554);
nor U31998 (N_31998,N_30275,N_30838);
xor U31999 (N_31999,N_30553,N_30070);
nor U32000 (N_32000,N_31836,N_31810);
and U32001 (N_32001,N_31672,N_31545);
or U32002 (N_32002,N_31544,N_31042);
xor U32003 (N_32003,N_31803,N_31126);
and U32004 (N_32004,N_31727,N_31409);
xnor U32005 (N_32005,N_31040,N_31826);
or U32006 (N_32006,N_31453,N_31934);
or U32007 (N_32007,N_31654,N_31266);
or U32008 (N_32008,N_31228,N_31804);
nand U32009 (N_32009,N_31820,N_31536);
or U32010 (N_32010,N_31895,N_31915);
or U32011 (N_32011,N_31220,N_31921);
nor U32012 (N_32012,N_31087,N_31842);
and U32013 (N_32013,N_31492,N_31817);
nor U32014 (N_32014,N_31923,N_31933);
and U32015 (N_32015,N_31257,N_31355);
or U32016 (N_32016,N_31527,N_31186);
xnor U32017 (N_32017,N_31778,N_31936);
xnor U32018 (N_32018,N_31956,N_31005);
nand U32019 (N_32019,N_31127,N_31128);
xor U32020 (N_32020,N_31738,N_31427);
or U32021 (N_32021,N_31911,N_31219);
and U32022 (N_32022,N_31213,N_31236);
nand U32023 (N_32023,N_31590,N_31606);
or U32024 (N_32024,N_31607,N_31084);
nor U32025 (N_32025,N_31295,N_31207);
or U32026 (N_32026,N_31902,N_31748);
xor U32027 (N_32027,N_31206,N_31857);
or U32028 (N_32028,N_31404,N_31178);
nor U32029 (N_32029,N_31106,N_31929);
xor U32030 (N_32030,N_31979,N_31839);
nor U32031 (N_32031,N_31208,N_31927);
and U32032 (N_32032,N_31299,N_31007);
nand U32033 (N_32033,N_31950,N_31639);
and U32034 (N_32034,N_31449,N_31474);
and U32035 (N_32035,N_31098,N_31522);
xor U32036 (N_32036,N_31035,N_31258);
nor U32037 (N_32037,N_31465,N_31766);
and U32038 (N_32038,N_31070,N_31452);
xnor U32039 (N_32039,N_31556,N_31702);
and U32040 (N_32040,N_31381,N_31942);
xor U32041 (N_32041,N_31245,N_31154);
and U32042 (N_32042,N_31442,N_31670);
xnor U32043 (N_32043,N_31759,N_31172);
and U32044 (N_32044,N_31359,N_31507);
and U32045 (N_32045,N_31510,N_31113);
nor U32046 (N_32046,N_31852,N_31109);
nand U32047 (N_32047,N_31749,N_31982);
xor U32048 (N_32048,N_31953,N_31612);
and U32049 (N_32049,N_31231,N_31755);
nor U32050 (N_32050,N_31275,N_31673);
nor U32051 (N_32051,N_31320,N_31588);
xor U32052 (N_32052,N_31387,N_31580);
xor U32053 (N_32053,N_31402,N_31559);
nand U32054 (N_32054,N_31989,N_31488);
nor U32055 (N_32055,N_31124,N_31284);
nand U32056 (N_32056,N_31045,N_31781);
nand U32057 (N_32057,N_31656,N_31578);
and U32058 (N_32058,N_31615,N_31688);
or U32059 (N_32059,N_31288,N_31726);
and U32060 (N_32060,N_31375,N_31062);
xor U32061 (N_32061,N_31369,N_31036);
and U32062 (N_32062,N_31379,N_31205);
nand U32063 (N_32063,N_31175,N_31669);
and U32064 (N_32064,N_31912,N_31383);
nor U32065 (N_32065,N_31489,N_31156);
xor U32066 (N_32066,N_31159,N_31714);
nor U32067 (N_32067,N_31535,N_31328);
nand U32068 (N_32068,N_31451,N_31722);
xnor U32069 (N_32069,N_31708,N_31573);
xnor U32070 (N_32070,N_31102,N_31283);
nand U32071 (N_32071,N_31420,N_31300);
or U32072 (N_32072,N_31905,N_31017);
nand U32073 (N_32073,N_31813,N_31278);
and U32074 (N_32074,N_31783,N_31909);
nor U32075 (N_32075,N_31082,N_31080);
and U32076 (N_32076,N_31692,N_31318);
nor U32077 (N_32077,N_31408,N_31282);
nor U32078 (N_32078,N_31610,N_31091);
or U32079 (N_32079,N_31486,N_31724);
or U32080 (N_32080,N_31533,N_31313);
and U32081 (N_32081,N_31711,N_31097);
xor U32082 (N_32082,N_31104,N_31643);
and U32083 (N_32083,N_31890,N_31757);
nor U32084 (N_32084,N_31083,N_31562);
nor U32085 (N_32085,N_31150,N_31806);
or U32086 (N_32086,N_31189,N_31210);
nand U32087 (N_32087,N_31763,N_31505);
nand U32088 (N_32088,N_31430,N_31553);
or U32089 (N_32089,N_31253,N_31149);
or U32090 (N_32090,N_31233,N_31260);
xor U32091 (N_32091,N_31495,N_31770);
or U32092 (N_32092,N_31021,N_31595);
and U32093 (N_32093,N_31437,N_31309);
nand U32094 (N_32094,N_31114,N_31237);
or U32095 (N_32095,N_31779,N_31843);
and U32096 (N_32096,N_31286,N_31006);
xnor U32097 (N_32097,N_31012,N_31315);
and U32098 (N_32098,N_31107,N_31191);
nand U32099 (N_32099,N_31686,N_31725);
and U32100 (N_32100,N_31969,N_31509);
xor U32101 (N_32101,N_31223,N_31135);
nor U32102 (N_32102,N_31877,N_31690);
and U32103 (N_32103,N_31424,N_31745);
nor U32104 (N_32104,N_31517,N_31940);
nor U32105 (N_32105,N_31646,N_31202);
nor U32106 (N_32106,N_31808,N_31963);
nand U32107 (N_32107,N_31425,N_31576);
and U32108 (N_32108,N_31732,N_31209);
nand U32109 (N_32109,N_31119,N_31914);
and U32110 (N_32110,N_31976,N_31805);
nand U32111 (N_32111,N_31644,N_31992);
xnor U32112 (N_32112,N_31086,N_31957);
nor U32113 (N_32113,N_31141,N_31234);
or U32114 (N_32114,N_31008,N_31990);
or U32115 (N_32115,N_31397,N_31329);
nor U32116 (N_32116,N_31037,N_31818);
or U32117 (N_32117,N_31991,N_31735);
or U32118 (N_32118,N_31377,N_31652);
xor U32119 (N_32119,N_31853,N_31750);
or U32120 (N_32120,N_31078,N_31326);
or U32121 (N_32121,N_31807,N_31193);
nor U32122 (N_32122,N_31985,N_31226);
nor U32123 (N_32123,N_31015,N_31687);
xnor U32124 (N_32124,N_31565,N_31602);
xnor U32125 (N_32125,N_31401,N_31906);
nand U32126 (N_32126,N_31204,N_31583);
and U32127 (N_32127,N_31541,N_31621);
nor U32128 (N_32128,N_31334,N_31613);
xnor U32129 (N_32129,N_31285,N_31540);
nand U32130 (N_32130,N_31648,N_31306);
nand U32131 (N_32131,N_31019,N_31052);
xnor U32132 (N_32132,N_31693,N_31589);
xnor U32133 (N_32133,N_31461,N_31919);
nor U32134 (N_32134,N_31938,N_31790);
and U32135 (N_32135,N_31605,N_31626);
nor U32136 (N_32136,N_31993,N_31865);
or U32137 (N_32137,N_31782,N_31618);
xor U32138 (N_32138,N_31887,N_31632);
nor U32139 (N_32139,N_31834,N_31366);
nand U32140 (N_32140,N_31094,N_31571);
and U32141 (N_32141,N_31352,N_31166);
nor U32142 (N_32142,N_31473,N_31570);
xnor U32143 (N_32143,N_31214,N_31970);
xnor U32144 (N_32144,N_31707,N_31044);
nand U32145 (N_32145,N_31450,N_31415);
or U32146 (N_32146,N_31279,N_31767);
and U32147 (N_32147,N_31534,N_31860);
nor U32148 (N_32148,N_31439,N_31247);
nand U32149 (N_32149,N_31876,N_31203);
xnor U32150 (N_32150,N_31825,N_31764);
and U32151 (N_32151,N_31793,N_31162);
nand U32152 (N_32152,N_31350,N_31551);
nor U32153 (N_32153,N_31868,N_31068);
nor U32154 (N_32154,N_31248,N_31229);
nand U32155 (N_32155,N_31034,N_31685);
and U32156 (N_32156,N_31875,N_31776);
or U32157 (N_32157,N_31682,N_31872);
xor U32158 (N_32158,N_31343,N_31252);
nand U32159 (N_32159,N_31182,N_31059);
or U32160 (N_32160,N_31634,N_31038);
and U32161 (N_32161,N_31893,N_31396);
nand U32162 (N_32162,N_31294,N_31411);
xnor U32163 (N_32163,N_31557,N_31768);
nand U32164 (N_32164,N_31760,N_31600);
nand U32165 (N_32165,N_31471,N_31357);
nor U32166 (N_32166,N_31703,N_31910);
or U32167 (N_32167,N_31122,N_31538);
nand U32168 (N_32168,N_31809,N_31271);
xor U32169 (N_32169,N_31561,N_31997);
nor U32170 (N_32170,N_31093,N_31001);
or U32171 (N_32171,N_31624,N_31617);
nor U32172 (N_32172,N_31130,N_31849);
xnor U32173 (N_32173,N_31095,N_31668);
xnor U32174 (N_32174,N_31847,N_31344);
xnor U32175 (N_32175,N_31874,N_31892);
or U32176 (N_32176,N_31597,N_31330);
or U32177 (N_32177,N_31577,N_31242);
or U32178 (N_32178,N_31593,N_31504);
nand U32179 (N_32179,N_31143,N_31096);
and U32180 (N_32180,N_31569,N_31072);
nor U32181 (N_32181,N_31903,N_31477);
and U32182 (N_32182,N_31647,N_31697);
and U32183 (N_32183,N_31947,N_31394);
nand U32184 (N_32184,N_31199,N_31152);
nand U32185 (N_32185,N_31188,N_31981);
or U32186 (N_32186,N_31163,N_31446);
or U32187 (N_32187,N_31462,N_31429);
and U32188 (N_32188,N_31850,N_31838);
or U32189 (N_32189,N_31515,N_31512);
and U32190 (N_32190,N_31530,N_31131);
or U32191 (N_32191,N_31251,N_31389);
xor U32192 (N_32192,N_31321,N_31388);
nor U32193 (N_32193,N_31314,N_31476);
or U32194 (N_32194,N_31882,N_31201);
nand U32195 (N_32195,N_31901,N_31419);
nand U32196 (N_32196,N_31448,N_31659);
nor U32197 (N_32197,N_31625,N_31884);
nand U32198 (N_32198,N_31564,N_31787);
or U32199 (N_32199,N_31351,N_31599);
and U32200 (N_32200,N_31434,N_31926);
and U32201 (N_32201,N_31000,N_31758);
nand U32202 (N_32202,N_31835,N_31339);
xor U32203 (N_32203,N_31123,N_31115);
xor U32204 (N_32204,N_31291,N_31497);
or U32205 (N_32205,N_31814,N_31939);
nand U32206 (N_32206,N_31460,N_31503);
nor U32207 (N_32207,N_31470,N_31658);
nor U32208 (N_32208,N_31443,N_31650);
and U32209 (N_32209,N_31145,N_31620);
nor U32210 (N_32210,N_31418,N_31752);
or U32211 (N_32211,N_31792,N_31338);
xor U32212 (N_32212,N_31341,N_31480);
nand U32213 (N_32213,N_31550,N_31681);
nor U32214 (N_32214,N_31880,N_31706);
and U32215 (N_32215,N_31274,N_31181);
xnor U32216 (N_32216,N_31454,N_31636);
xnor U32217 (N_32217,N_31928,N_31340);
nor U32218 (N_32218,N_31160,N_31854);
or U32219 (N_32219,N_31523,N_31904);
or U32220 (N_32220,N_31064,N_31691);
and U32221 (N_32221,N_31728,N_31346);
nor U32222 (N_32222,N_31500,N_31406);
or U32223 (N_32223,N_31116,N_31709);
and U32224 (N_32224,N_31185,N_31302);
and U32225 (N_32225,N_31713,N_31718);
nor U32226 (N_32226,N_31134,N_31312);
xnor U32227 (N_32227,N_31563,N_31864);
xnor U32228 (N_32228,N_31305,N_31103);
and U32229 (N_32229,N_31676,N_31241);
or U32230 (N_32230,N_31878,N_31308);
nor U32231 (N_32231,N_31074,N_31655);
nand U32232 (N_32232,N_31705,N_31018);
nor U32233 (N_32233,N_31458,N_31235);
xor U32234 (N_32234,N_31296,N_31378);
or U32235 (N_32235,N_31791,N_31053);
nor U32236 (N_32236,N_31431,N_31977);
xor U32237 (N_32237,N_31002,N_31494);
nand U32238 (N_32238,N_31325,N_31367);
and U32239 (N_32239,N_31348,N_31974);
nand U32240 (N_32240,N_31873,N_31537);
nor U32241 (N_32241,N_31054,N_31171);
or U32242 (N_32242,N_31372,N_31640);
and U32243 (N_32243,N_31319,N_31555);
xnor U32244 (N_32244,N_31572,N_31829);
and U32245 (N_32245,N_31591,N_31525);
nor U32246 (N_32246,N_31031,N_31332);
and U32247 (N_32247,N_31586,N_31773);
nand U32248 (N_32248,N_31333,N_31469);
and U32249 (N_32249,N_31496,N_31222);
xnor U32250 (N_32250,N_31400,N_31949);
and U32251 (N_32251,N_31975,N_31121);
xnor U32252 (N_32252,N_31310,N_31117);
xor U32253 (N_32253,N_31441,N_31033);
and U32254 (N_32254,N_31678,N_31444);
nand U32255 (N_32255,N_31243,N_31614);
nor U32256 (N_32256,N_31290,N_31794);
and U32257 (N_32257,N_31965,N_31240);
xor U32258 (N_32258,N_31393,N_31174);
nand U32259 (N_32259,N_31165,N_31177);
nand U32260 (N_32260,N_31812,N_31558);
nor U32261 (N_32261,N_31828,N_31280);
and U32262 (N_32262,N_31049,N_31730);
nand U32263 (N_32263,N_31513,N_31567);
nand U32264 (N_32264,N_31399,N_31827);
and U32265 (N_32265,N_31548,N_31866);
and U32266 (N_32266,N_31298,N_31520);
or U32267 (N_32267,N_31373,N_31638);
or U32268 (N_32268,N_31039,N_31137);
or U32269 (N_32269,N_31841,N_31467);
nor U32270 (N_32270,N_31629,N_31978);
xor U32271 (N_32271,N_31907,N_31362);
and U32272 (N_32272,N_31491,N_31741);
xor U32273 (N_32273,N_31365,N_31061);
and U32274 (N_32274,N_31777,N_31475);
and U32275 (N_32275,N_31047,N_31723);
or U32276 (N_32276,N_31657,N_31742);
xor U32277 (N_32277,N_31932,N_31604);
nand U32278 (N_32278,N_31347,N_31376);
and U32279 (N_32279,N_31317,N_31584);
nor U32280 (N_32280,N_31153,N_31746);
xor U32281 (N_32281,N_31633,N_31421);
or U32282 (N_32282,N_31016,N_31164);
xor U32283 (N_32283,N_31830,N_31661);
nor U32284 (N_32284,N_31870,N_31984);
nand U32285 (N_32285,N_31816,N_31631);
and U32286 (N_32286,N_31058,N_31958);
and U32287 (N_32287,N_31345,N_31844);
xnor U32288 (N_32288,N_31771,N_31071);
nor U32289 (N_32289,N_31144,N_31526);
or U32290 (N_32290,N_31195,N_31256);
nand U32291 (N_32291,N_31414,N_31867);
nand U32292 (N_32292,N_31024,N_31224);
xor U32293 (N_32293,N_31753,N_31802);
or U32294 (N_32294,N_31221,N_31772);
or U32295 (N_32295,N_31013,N_31342);
or U32296 (N_32296,N_31955,N_31148);
nor U32297 (N_32297,N_31754,N_31821);
nor U32298 (N_32298,N_31079,N_31798);
or U32299 (N_32299,N_31920,N_31667);
or U32300 (N_32300,N_31898,N_31761);
nand U32301 (N_32301,N_31239,N_31729);
xnor U32302 (N_32302,N_31531,N_31627);
nor U32303 (N_32303,N_31133,N_31010);
and U32304 (N_32304,N_31931,N_31412);
nand U32305 (N_32305,N_31370,N_31263);
xor U32306 (N_32306,N_31216,N_31717);
nand U32307 (N_32307,N_31304,N_31581);
or U32308 (N_32308,N_31695,N_31698);
and U32309 (N_32309,N_31436,N_31869);
and U32310 (N_32310,N_31384,N_31398);
and U32311 (N_32311,N_31960,N_31076);
nor U32312 (N_32312,N_31392,N_31215);
nand U32313 (N_32313,N_31894,N_31200);
nand U32314 (N_32314,N_31679,N_31478);
nor U32315 (N_32315,N_31785,N_31187);
xor U32316 (N_32316,N_31170,N_31996);
and U32317 (N_32317,N_31311,N_31479);
and U32318 (N_32318,N_31316,N_31273);
and U32319 (N_32319,N_31374,N_31218);
xor U32320 (N_32320,N_31270,N_31100);
xor U32321 (N_32321,N_31542,N_31025);
nor U32322 (N_32322,N_31050,N_31246);
and U32323 (N_32323,N_31155,N_31579);
nand U32324 (N_32324,N_31999,N_31323);
xor U32325 (N_32325,N_31788,N_31023);
and U32326 (N_32326,N_31734,N_31712);
xnor U32327 (N_32327,N_31307,N_31603);
and U32328 (N_32328,N_31566,N_31995);
or U32329 (N_32329,N_31660,N_31490);
nor U32330 (N_32330,N_31032,N_31716);
nor U32331 (N_32331,N_31699,N_31554);
nor U32332 (N_32332,N_31980,N_31780);
xnor U32333 (N_32333,N_31353,N_31549);
nand U32334 (N_32334,N_31769,N_31674);
and U32335 (N_32335,N_31371,N_31719);
and U32336 (N_32336,N_31030,N_31085);
xnor U32337 (N_32337,N_31710,N_31261);
nand U32338 (N_32338,N_31067,N_31184);
nand U32339 (N_32339,N_31951,N_31514);
or U32340 (N_32340,N_31484,N_31594);
nand U32341 (N_32341,N_31922,N_31403);
or U32342 (N_32342,N_31180,N_31823);
nor U32343 (N_32343,N_31861,N_31731);
xor U32344 (N_32344,N_31238,N_31740);
and U32345 (N_32345,N_31879,N_31945);
nand U32346 (N_32346,N_31651,N_31060);
nand U32347 (N_32347,N_31268,N_31161);
or U32348 (N_32348,N_31988,N_31587);
nor U32349 (N_32349,N_31151,N_31846);
and U32350 (N_32350,N_31608,N_31382);
nor U32351 (N_32351,N_31158,N_31671);
nor U32352 (N_32352,N_31715,N_31575);
and U32353 (N_32353,N_31292,N_31508);
nand U32354 (N_32354,N_31831,N_31635);
xor U32355 (N_32355,N_31386,N_31139);
nand U32356 (N_32356,N_31485,N_31499);
nand U32357 (N_32357,N_31455,N_31466);
nor U32358 (N_32358,N_31972,N_31363);
and U32359 (N_32359,N_31147,N_31211);
nor U32360 (N_32360,N_31385,N_31028);
xor U32361 (N_32361,N_31637,N_31413);
or U32362 (N_32362,N_31003,N_31129);
and U32363 (N_32363,N_31183,N_31254);
nand U32364 (N_32364,N_31649,N_31360);
xnor U32365 (N_32365,N_31736,N_31743);
and U32366 (N_32366,N_31789,N_31796);
or U32367 (N_32367,N_31354,N_31361);
nand U32368 (N_32368,N_31026,N_31293);
nor U32369 (N_32369,N_31250,N_31459);
nor U32370 (N_32370,N_31837,N_31800);
xor U32371 (N_32371,N_31848,N_31368);
nor U32372 (N_32372,N_31675,N_31851);
xnor U32373 (N_32373,N_31666,N_31762);
xnor U32374 (N_32374,N_31998,N_31009);
and U32375 (N_32375,N_31108,N_31198);
nand U32376 (N_32376,N_31582,N_31801);
nor U32377 (N_32377,N_31063,N_31983);
or U32378 (N_32378,N_31498,N_31324);
nor U32379 (N_32379,N_31696,N_31822);
and U32380 (N_32380,N_31964,N_31303);
nor U32381 (N_32381,N_31881,N_31701);
or U32382 (N_32382,N_31179,N_31733);
nand U32383 (N_32383,N_31653,N_31774);
or U32384 (N_32384,N_31546,N_31528);
xnor U32385 (N_32385,N_31410,N_31616);
nor U32386 (N_32386,N_31112,N_31663);
nor U32387 (N_32387,N_31721,N_31069);
and U32388 (N_32388,N_31259,N_31986);
nand U32389 (N_32389,N_31518,N_31751);
and U32390 (N_32390,N_31720,N_31176);
and U32391 (N_32391,N_31468,N_31694);
and U32392 (N_32392,N_31547,N_31786);
or U32393 (N_32393,N_31457,N_31739);
nor U32394 (N_32394,N_31322,N_31066);
nor U32395 (N_32395,N_31856,N_31407);
xor U32396 (N_32396,N_31105,N_31700);
xnor U32397 (N_32397,N_31232,N_31438);
nor U32398 (N_32398,N_31568,N_31560);
or U32399 (N_32399,N_31088,N_31432);
and U32400 (N_32400,N_31433,N_31885);
nand U32401 (N_32401,N_31775,N_31090);
xnor U32402 (N_32402,N_31611,N_31335);
nand U32403 (N_32403,N_31125,N_31886);
nor U32404 (N_32404,N_31994,N_31004);
nor U32405 (N_32405,N_31048,N_31011);
and U32406 (N_32406,N_31987,N_31765);
nand U32407 (N_32407,N_31623,N_31840);
nor U32408 (N_32408,N_31502,N_31287);
and U32409 (N_32409,N_31930,N_31337);
and U32410 (N_32410,N_31422,N_31811);
nor U32411 (N_32411,N_31883,N_31684);
xnor U32412 (N_32412,N_31301,N_31795);
nor U32413 (N_32413,N_31642,N_31140);
xnor U32414 (N_32414,N_31440,N_31941);
xor U32415 (N_32415,N_31390,N_31022);
nand U32416 (N_32416,N_31281,N_31543);
and U32417 (N_32417,N_31967,N_31212);
nand U32418 (N_32418,N_31269,N_31845);
nor U32419 (N_32419,N_31099,N_31092);
nor U32420 (N_32420,N_31364,N_31395);
or U32421 (N_32421,N_31046,N_31483);
xor U32422 (N_32422,N_31255,N_31120);
or U32423 (N_32423,N_31959,N_31824);
nor U32424 (N_32424,N_31924,N_31056);
nand U32425 (N_32425,N_31157,N_31417);
or U32426 (N_32426,N_31689,N_31871);
xnor U32427 (N_32427,N_31973,N_31908);
xnor U32428 (N_32428,N_31797,N_31356);
nand U32429 (N_32429,N_31196,N_31426);
nor U32430 (N_32430,N_31968,N_31487);
nand U32431 (N_32431,N_31336,N_31173);
nor U32432 (N_32432,N_31622,N_31267);
nand U32433 (N_32433,N_31598,N_31948);
xor U32434 (N_32434,N_31516,N_31896);
or U32435 (N_32435,N_31832,N_31416);
nor U32436 (N_32436,N_31925,N_31574);
nor U32437 (N_32437,N_31227,N_31506);
nor U32438 (N_32438,N_31815,N_31020);
nor U32439 (N_32439,N_31737,N_31552);
xor U32440 (N_32440,N_31971,N_31349);
nor U32441 (N_32441,N_31065,N_31075);
nand U32442 (N_32442,N_31858,N_31862);
nand U32443 (N_32443,N_31521,N_31327);
xor U32444 (N_32444,N_31665,N_31511);
or U32445 (N_32445,N_31519,N_31194);
xor U32446 (N_32446,N_31619,N_31423);
and U32447 (N_32447,N_31073,N_31089);
nor U32448 (N_32448,N_31081,N_31916);
or U32449 (N_32449,N_31833,N_31380);
xor U32450 (N_32450,N_31331,N_31532);
nor U32451 (N_32451,N_31954,N_31913);
and U32452 (N_32452,N_31272,N_31799);
and U32453 (N_32453,N_31677,N_31704);
xnor U32454 (N_32454,N_31146,N_31900);
and U32455 (N_32455,N_31592,N_31944);
nor U32456 (N_32456,N_31961,N_31264);
or U32457 (N_32457,N_31277,N_31217);
and U32458 (N_32458,N_31493,N_31641);
xnor U32459 (N_32459,N_31077,N_31230);
nand U32460 (N_32460,N_31888,N_31169);
nor U32461 (N_32461,N_31680,N_31585);
nand U32462 (N_32462,N_31265,N_31014);
and U32463 (N_32463,N_31276,N_31167);
or U32464 (N_32464,N_31168,N_31744);
or U32465 (N_32465,N_31055,N_31859);
xnor U32466 (N_32466,N_31897,N_31937);
nand U32467 (N_32467,N_31043,N_31952);
nand U32468 (N_32468,N_31962,N_31110);
xnor U32469 (N_32469,N_31192,N_31917);
or U32470 (N_32470,N_31784,N_31136);
nor U32471 (N_32471,N_31946,N_31118);
xnor U32472 (N_32472,N_31297,N_31628);
nand U32473 (N_32473,N_31456,N_31111);
nand U32474 (N_32474,N_31662,N_31445);
and U32475 (N_32475,N_31041,N_31630);
or U32476 (N_32476,N_31539,N_31464);
or U32477 (N_32477,N_31482,N_31027);
nand U32478 (N_32478,N_31943,N_31889);
nand U32479 (N_32479,N_31132,N_31601);
xnor U32480 (N_32480,N_31501,N_31596);
nor U32481 (N_32481,N_31249,N_31244);
or U32482 (N_32482,N_31529,N_31190);
or U32483 (N_32483,N_31664,N_31899);
nand U32484 (N_32484,N_31855,N_31029);
nand U32485 (N_32485,N_31472,N_31966);
and U32486 (N_32486,N_31358,N_31463);
nand U32487 (N_32487,N_31262,N_31428);
nand U32488 (N_32488,N_31863,N_31101);
nor U32489 (N_32489,N_31683,N_31057);
and U32490 (N_32490,N_31142,N_31524);
nor U32491 (N_32491,N_31391,N_31609);
and U32492 (N_32492,N_31645,N_31891);
nor U32493 (N_32493,N_31447,N_31747);
and U32494 (N_32494,N_31935,N_31481);
and U32495 (N_32495,N_31289,N_31197);
nand U32496 (N_32496,N_31756,N_31819);
nor U32497 (N_32497,N_31051,N_31918);
nor U32498 (N_32498,N_31225,N_31435);
xor U32499 (N_32499,N_31405,N_31138);
nand U32500 (N_32500,N_31995,N_31741);
xor U32501 (N_32501,N_31121,N_31055);
or U32502 (N_32502,N_31648,N_31275);
nand U32503 (N_32503,N_31896,N_31036);
nand U32504 (N_32504,N_31300,N_31839);
xnor U32505 (N_32505,N_31137,N_31512);
nor U32506 (N_32506,N_31620,N_31421);
or U32507 (N_32507,N_31751,N_31136);
nor U32508 (N_32508,N_31907,N_31707);
nor U32509 (N_32509,N_31047,N_31427);
nand U32510 (N_32510,N_31248,N_31473);
nor U32511 (N_32511,N_31561,N_31152);
or U32512 (N_32512,N_31550,N_31828);
or U32513 (N_32513,N_31076,N_31730);
and U32514 (N_32514,N_31758,N_31031);
nor U32515 (N_32515,N_31578,N_31597);
nor U32516 (N_32516,N_31955,N_31871);
and U32517 (N_32517,N_31499,N_31833);
nor U32518 (N_32518,N_31926,N_31276);
xnor U32519 (N_32519,N_31957,N_31583);
xor U32520 (N_32520,N_31977,N_31198);
xnor U32521 (N_32521,N_31290,N_31997);
or U32522 (N_32522,N_31936,N_31137);
xor U32523 (N_32523,N_31220,N_31659);
or U32524 (N_32524,N_31595,N_31144);
nand U32525 (N_32525,N_31913,N_31369);
nor U32526 (N_32526,N_31392,N_31999);
or U32527 (N_32527,N_31894,N_31992);
nand U32528 (N_32528,N_31272,N_31402);
and U32529 (N_32529,N_31921,N_31967);
nand U32530 (N_32530,N_31984,N_31288);
nor U32531 (N_32531,N_31600,N_31627);
nor U32532 (N_32532,N_31502,N_31300);
nand U32533 (N_32533,N_31155,N_31535);
nand U32534 (N_32534,N_31745,N_31121);
nor U32535 (N_32535,N_31716,N_31031);
nor U32536 (N_32536,N_31901,N_31171);
and U32537 (N_32537,N_31795,N_31012);
or U32538 (N_32538,N_31988,N_31001);
nor U32539 (N_32539,N_31070,N_31516);
xor U32540 (N_32540,N_31385,N_31726);
nand U32541 (N_32541,N_31318,N_31133);
or U32542 (N_32542,N_31117,N_31263);
xor U32543 (N_32543,N_31390,N_31773);
or U32544 (N_32544,N_31461,N_31800);
xnor U32545 (N_32545,N_31501,N_31241);
or U32546 (N_32546,N_31520,N_31971);
nor U32547 (N_32547,N_31476,N_31015);
and U32548 (N_32548,N_31646,N_31025);
xor U32549 (N_32549,N_31390,N_31451);
xnor U32550 (N_32550,N_31709,N_31704);
xor U32551 (N_32551,N_31071,N_31050);
or U32552 (N_32552,N_31551,N_31198);
and U32553 (N_32553,N_31153,N_31816);
nor U32554 (N_32554,N_31429,N_31177);
nand U32555 (N_32555,N_31457,N_31254);
or U32556 (N_32556,N_31764,N_31259);
xor U32557 (N_32557,N_31040,N_31171);
xnor U32558 (N_32558,N_31466,N_31133);
xor U32559 (N_32559,N_31852,N_31417);
nand U32560 (N_32560,N_31677,N_31155);
and U32561 (N_32561,N_31363,N_31824);
and U32562 (N_32562,N_31597,N_31475);
nand U32563 (N_32563,N_31007,N_31654);
xnor U32564 (N_32564,N_31867,N_31098);
and U32565 (N_32565,N_31197,N_31469);
nand U32566 (N_32566,N_31241,N_31121);
nand U32567 (N_32567,N_31699,N_31497);
xor U32568 (N_32568,N_31695,N_31610);
nand U32569 (N_32569,N_31304,N_31604);
nand U32570 (N_32570,N_31868,N_31698);
nor U32571 (N_32571,N_31013,N_31675);
nand U32572 (N_32572,N_31096,N_31487);
nand U32573 (N_32573,N_31437,N_31570);
xnor U32574 (N_32574,N_31391,N_31828);
nor U32575 (N_32575,N_31577,N_31403);
nand U32576 (N_32576,N_31887,N_31608);
nand U32577 (N_32577,N_31837,N_31491);
or U32578 (N_32578,N_31252,N_31988);
nor U32579 (N_32579,N_31566,N_31627);
nand U32580 (N_32580,N_31044,N_31367);
and U32581 (N_32581,N_31125,N_31554);
nand U32582 (N_32582,N_31974,N_31337);
nor U32583 (N_32583,N_31702,N_31490);
nand U32584 (N_32584,N_31067,N_31249);
xor U32585 (N_32585,N_31003,N_31670);
or U32586 (N_32586,N_31829,N_31234);
xor U32587 (N_32587,N_31838,N_31581);
xnor U32588 (N_32588,N_31583,N_31673);
and U32589 (N_32589,N_31474,N_31447);
xnor U32590 (N_32590,N_31322,N_31925);
or U32591 (N_32591,N_31990,N_31197);
and U32592 (N_32592,N_31876,N_31129);
and U32593 (N_32593,N_31996,N_31027);
nand U32594 (N_32594,N_31649,N_31630);
nor U32595 (N_32595,N_31344,N_31747);
nor U32596 (N_32596,N_31022,N_31110);
xor U32597 (N_32597,N_31013,N_31938);
nor U32598 (N_32598,N_31686,N_31391);
or U32599 (N_32599,N_31919,N_31753);
and U32600 (N_32600,N_31763,N_31591);
and U32601 (N_32601,N_31086,N_31696);
nor U32602 (N_32602,N_31648,N_31809);
or U32603 (N_32603,N_31434,N_31799);
and U32604 (N_32604,N_31499,N_31599);
nor U32605 (N_32605,N_31555,N_31490);
xnor U32606 (N_32606,N_31448,N_31658);
or U32607 (N_32607,N_31863,N_31457);
nor U32608 (N_32608,N_31671,N_31016);
xnor U32609 (N_32609,N_31192,N_31898);
nand U32610 (N_32610,N_31565,N_31738);
or U32611 (N_32611,N_31238,N_31866);
nor U32612 (N_32612,N_31765,N_31806);
xor U32613 (N_32613,N_31595,N_31305);
nor U32614 (N_32614,N_31410,N_31861);
nand U32615 (N_32615,N_31617,N_31059);
nor U32616 (N_32616,N_31943,N_31248);
nor U32617 (N_32617,N_31842,N_31395);
xnor U32618 (N_32618,N_31024,N_31204);
nand U32619 (N_32619,N_31615,N_31915);
xor U32620 (N_32620,N_31793,N_31020);
nand U32621 (N_32621,N_31385,N_31164);
nor U32622 (N_32622,N_31964,N_31054);
nand U32623 (N_32623,N_31670,N_31049);
nor U32624 (N_32624,N_31529,N_31625);
nand U32625 (N_32625,N_31052,N_31508);
nand U32626 (N_32626,N_31294,N_31738);
and U32627 (N_32627,N_31630,N_31835);
xor U32628 (N_32628,N_31853,N_31246);
and U32629 (N_32629,N_31691,N_31093);
and U32630 (N_32630,N_31990,N_31403);
nor U32631 (N_32631,N_31853,N_31898);
nor U32632 (N_32632,N_31944,N_31453);
nand U32633 (N_32633,N_31378,N_31434);
nand U32634 (N_32634,N_31970,N_31673);
and U32635 (N_32635,N_31336,N_31932);
and U32636 (N_32636,N_31919,N_31376);
and U32637 (N_32637,N_31562,N_31036);
and U32638 (N_32638,N_31636,N_31577);
nor U32639 (N_32639,N_31329,N_31913);
or U32640 (N_32640,N_31055,N_31845);
or U32641 (N_32641,N_31123,N_31392);
nor U32642 (N_32642,N_31114,N_31540);
nand U32643 (N_32643,N_31787,N_31304);
xor U32644 (N_32644,N_31508,N_31507);
xnor U32645 (N_32645,N_31308,N_31523);
xnor U32646 (N_32646,N_31562,N_31459);
nand U32647 (N_32647,N_31275,N_31618);
and U32648 (N_32648,N_31299,N_31135);
and U32649 (N_32649,N_31002,N_31117);
nor U32650 (N_32650,N_31801,N_31655);
or U32651 (N_32651,N_31521,N_31623);
xnor U32652 (N_32652,N_31991,N_31318);
or U32653 (N_32653,N_31242,N_31930);
or U32654 (N_32654,N_31052,N_31253);
xnor U32655 (N_32655,N_31796,N_31494);
nand U32656 (N_32656,N_31252,N_31966);
nand U32657 (N_32657,N_31320,N_31407);
and U32658 (N_32658,N_31728,N_31611);
and U32659 (N_32659,N_31177,N_31702);
nand U32660 (N_32660,N_31878,N_31417);
nor U32661 (N_32661,N_31913,N_31014);
nor U32662 (N_32662,N_31050,N_31826);
and U32663 (N_32663,N_31967,N_31334);
nand U32664 (N_32664,N_31065,N_31598);
xnor U32665 (N_32665,N_31547,N_31608);
xor U32666 (N_32666,N_31610,N_31981);
nand U32667 (N_32667,N_31041,N_31856);
or U32668 (N_32668,N_31021,N_31222);
xnor U32669 (N_32669,N_31560,N_31700);
xnor U32670 (N_32670,N_31185,N_31927);
and U32671 (N_32671,N_31949,N_31907);
nor U32672 (N_32672,N_31092,N_31811);
or U32673 (N_32673,N_31821,N_31152);
or U32674 (N_32674,N_31565,N_31008);
and U32675 (N_32675,N_31197,N_31815);
nand U32676 (N_32676,N_31126,N_31621);
nor U32677 (N_32677,N_31420,N_31438);
nand U32678 (N_32678,N_31477,N_31408);
nor U32679 (N_32679,N_31783,N_31491);
and U32680 (N_32680,N_31462,N_31189);
xnor U32681 (N_32681,N_31305,N_31406);
xor U32682 (N_32682,N_31546,N_31583);
or U32683 (N_32683,N_31059,N_31194);
or U32684 (N_32684,N_31074,N_31625);
nor U32685 (N_32685,N_31440,N_31334);
nand U32686 (N_32686,N_31729,N_31563);
nand U32687 (N_32687,N_31222,N_31659);
nand U32688 (N_32688,N_31098,N_31120);
and U32689 (N_32689,N_31445,N_31572);
xor U32690 (N_32690,N_31147,N_31827);
and U32691 (N_32691,N_31467,N_31812);
nand U32692 (N_32692,N_31903,N_31737);
or U32693 (N_32693,N_31828,N_31754);
or U32694 (N_32694,N_31680,N_31270);
nand U32695 (N_32695,N_31014,N_31354);
or U32696 (N_32696,N_31228,N_31067);
xnor U32697 (N_32697,N_31575,N_31172);
or U32698 (N_32698,N_31176,N_31113);
nand U32699 (N_32699,N_31591,N_31168);
or U32700 (N_32700,N_31244,N_31870);
or U32701 (N_32701,N_31846,N_31510);
nor U32702 (N_32702,N_31244,N_31306);
nor U32703 (N_32703,N_31134,N_31256);
xor U32704 (N_32704,N_31580,N_31763);
and U32705 (N_32705,N_31011,N_31928);
nand U32706 (N_32706,N_31616,N_31300);
nand U32707 (N_32707,N_31302,N_31353);
and U32708 (N_32708,N_31597,N_31096);
and U32709 (N_32709,N_31248,N_31004);
and U32710 (N_32710,N_31193,N_31096);
nor U32711 (N_32711,N_31627,N_31625);
nor U32712 (N_32712,N_31603,N_31322);
and U32713 (N_32713,N_31317,N_31697);
nand U32714 (N_32714,N_31312,N_31589);
nor U32715 (N_32715,N_31714,N_31653);
or U32716 (N_32716,N_31074,N_31874);
xor U32717 (N_32717,N_31301,N_31785);
nor U32718 (N_32718,N_31889,N_31873);
xnor U32719 (N_32719,N_31666,N_31618);
nor U32720 (N_32720,N_31144,N_31754);
and U32721 (N_32721,N_31058,N_31312);
or U32722 (N_32722,N_31449,N_31256);
or U32723 (N_32723,N_31342,N_31645);
nand U32724 (N_32724,N_31136,N_31313);
and U32725 (N_32725,N_31469,N_31170);
xor U32726 (N_32726,N_31048,N_31597);
xnor U32727 (N_32727,N_31178,N_31319);
nor U32728 (N_32728,N_31896,N_31747);
nor U32729 (N_32729,N_31325,N_31407);
and U32730 (N_32730,N_31003,N_31827);
nand U32731 (N_32731,N_31099,N_31633);
and U32732 (N_32732,N_31112,N_31881);
or U32733 (N_32733,N_31189,N_31387);
or U32734 (N_32734,N_31864,N_31397);
xnor U32735 (N_32735,N_31289,N_31917);
nor U32736 (N_32736,N_31713,N_31013);
xnor U32737 (N_32737,N_31836,N_31750);
or U32738 (N_32738,N_31642,N_31794);
nor U32739 (N_32739,N_31052,N_31070);
and U32740 (N_32740,N_31260,N_31695);
and U32741 (N_32741,N_31721,N_31220);
xor U32742 (N_32742,N_31095,N_31827);
nand U32743 (N_32743,N_31602,N_31161);
and U32744 (N_32744,N_31545,N_31869);
xnor U32745 (N_32745,N_31450,N_31568);
nor U32746 (N_32746,N_31412,N_31648);
nor U32747 (N_32747,N_31861,N_31437);
nand U32748 (N_32748,N_31801,N_31908);
xor U32749 (N_32749,N_31897,N_31697);
or U32750 (N_32750,N_31945,N_31119);
nand U32751 (N_32751,N_31383,N_31266);
nand U32752 (N_32752,N_31047,N_31846);
nor U32753 (N_32753,N_31124,N_31462);
xnor U32754 (N_32754,N_31419,N_31346);
nand U32755 (N_32755,N_31456,N_31933);
or U32756 (N_32756,N_31276,N_31588);
xor U32757 (N_32757,N_31032,N_31282);
nand U32758 (N_32758,N_31094,N_31779);
nor U32759 (N_32759,N_31448,N_31003);
and U32760 (N_32760,N_31222,N_31132);
xnor U32761 (N_32761,N_31872,N_31306);
nand U32762 (N_32762,N_31672,N_31296);
nor U32763 (N_32763,N_31927,N_31655);
nand U32764 (N_32764,N_31790,N_31670);
and U32765 (N_32765,N_31853,N_31419);
or U32766 (N_32766,N_31680,N_31376);
and U32767 (N_32767,N_31173,N_31653);
nand U32768 (N_32768,N_31571,N_31265);
and U32769 (N_32769,N_31288,N_31273);
xor U32770 (N_32770,N_31351,N_31010);
nand U32771 (N_32771,N_31939,N_31740);
and U32772 (N_32772,N_31832,N_31814);
xor U32773 (N_32773,N_31382,N_31777);
nor U32774 (N_32774,N_31336,N_31913);
nor U32775 (N_32775,N_31224,N_31263);
and U32776 (N_32776,N_31504,N_31679);
and U32777 (N_32777,N_31169,N_31589);
nand U32778 (N_32778,N_31709,N_31804);
or U32779 (N_32779,N_31391,N_31647);
and U32780 (N_32780,N_31174,N_31111);
nor U32781 (N_32781,N_31881,N_31521);
nand U32782 (N_32782,N_31220,N_31032);
xnor U32783 (N_32783,N_31237,N_31571);
xnor U32784 (N_32784,N_31420,N_31025);
and U32785 (N_32785,N_31688,N_31138);
and U32786 (N_32786,N_31715,N_31546);
nor U32787 (N_32787,N_31062,N_31286);
xor U32788 (N_32788,N_31841,N_31557);
and U32789 (N_32789,N_31569,N_31330);
or U32790 (N_32790,N_31055,N_31101);
xor U32791 (N_32791,N_31481,N_31383);
and U32792 (N_32792,N_31268,N_31142);
and U32793 (N_32793,N_31450,N_31576);
or U32794 (N_32794,N_31420,N_31550);
and U32795 (N_32795,N_31975,N_31941);
xor U32796 (N_32796,N_31856,N_31817);
xnor U32797 (N_32797,N_31742,N_31781);
nand U32798 (N_32798,N_31994,N_31394);
or U32799 (N_32799,N_31517,N_31983);
nand U32800 (N_32800,N_31170,N_31834);
nand U32801 (N_32801,N_31336,N_31217);
xor U32802 (N_32802,N_31949,N_31737);
xnor U32803 (N_32803,N_31089,N_31675);
or U32804 (N_32804,N_31140,N_31045);
or U32805 (N_32805,N_31592,N_31965);
nand U32806 (N_32806,N_31641,N_31559);
or U32807 (N_32807,N_31159,N_31326);
or U32808 (N_32808,N_31118,N_31564);
xor U32809 (N_32809,N_31331,N_31492);
nor U32810 (N_32810,N_31537,N_31847);
nand U32811 (N_32811,N_31337,N_31239);
and U32812 (N_32812,N_31225,N_31374);
nand U32813 (N_32813,N_31614,N_31130);
or U32814 (N_32814,N_31135,N_31644);
or U32815 (N_32815,N_31047,N_31141);
or U32816 (N_32816,N_31778,N_31743);
nor U32817 (N_32817,N_31965,N_31237);
or U32818 (N_32818,N_31524,N_31365);
or U32819 (N_32819,N_31542,N_31847);
nand U32820 (N_32820,N_31696,N_31716);
nand U32821 (N_32821,N_31766,N_31526);
or U32822 (N_32822,N_31654,N_31106);
xnor U32823 (N_32823,N_31318,N_31118);
xor U32824 (N_32824,N_31459,N_31384);
nor U32825 (N_32825,N_31004,N_31543);
or U32826 (N_32826,N_31226,N_31305);
nor U32827 (N_32827,N_31484,N_31589);
and U32828 (N_32828,N_31879,N_31917);
or U32829 (N_32829,N_31079,N_31917);
and U32830 (N_32830,N_31826,N_31970);
and U32831 (N_32831,N_31563,N_31413);
and U32832 (N_32832,N_31473,N_31738);
nand U32833 (N_32833,N_31715,N_31796);
xnor U32834 (N_32834,N_31673,N_31299);
nand U32835 (N_32835,N_31134,N_31099);
and U32836 (N_32836,N_31025,N_31935);
and U32837 (N_32837,N_31024,N_31096);
nand U32838 (N_32838,N_31170,N_31643);
nand U32839 (N_32839,N_31133,N_31991);
and U32840 (N_32840,N_31531,N_31179);
nand U32841 (N_32841,N_31870,N_31691);
and U32842 (N_32842,N_31257,N_31307);
nor U32843 (N_32843,N_31183,N_31507);
or U32844 (N_32844,N_31058,N_31635);
or U32845 (N_32845,N_31389,N_31286);
and U32846 (N_32846,N_31071,N_31297);
nand U32847 (N_32847,N_31714,N_31434);
xnor U32848 (N_32848,N_31600,N_31526);
or U32849 (N_32849,N_31487,N_31592);
nor U32850 (N_32850,N_31795,N_31582);
or U32851 (N_32851,N_31269,N_31139);
nand U32852 (N_32852,N_31780,N_31064);
and U32853 (N_32853,N_31428,N_31842);
nand U32854 (N_32854,N_31679,N_31768);
nand U32855 (N_32855,N_31785,N_31509);
and U32856 (N_32856,N_31912,N_31072);
xor U32857 (N_32857,N_31614,N_31930);
nor U32858 (N_32858,N_31848,N_31637);
or U32859 (N_32859,N_31051,N_31389);
xor U32860 (N_32860,N_31522,N_31877);
nand U32861 (N_32861,N_31229,N_31629);
and U32862 (N_32862,N_31275,N_31933);
or U32863 (N_32863,N_31219,N_31469);
or U32864 (N_32864,N_31314,N_31514);
nor U32865 (N_32865,N_31809,N_31013);
or U32866 (N_32866,N_31272,N_31596);
nor U32867 (N_32867,N_31532,N_31904);
xor U32868 (N_32868,N_31652,N_31011);
or U32869 (N_32869,N_31141,N_31796);
nor U32870 (N_32870,N_31686,N_31752);
or U32871 (N_32871,N_31847,N_31582);
or U32872 (N_32872,N_31800,N_31181);
and U32873 (N_32873,N_31524,N_31367);
nand U32874 (N_32874,N_31293,N_31782);
nor U32875 (N_32875,N_31178,N_31974);
nand U32876 (N_32876,N_31051,N_31990);
nand U32877 (N_32877,N_31752,N_31657);
xor U32878 (N_32878,N_31637,N_31639);
nand U32879 (N_32879,N_31575,N_31438);
nor U32880 (N_32880,N_31428,N_31865);
or U32881 (N_32881,N_31251,N_31310);
xnor U32882 (N_32882,N_31501,N_31153);
xnor U32883 (N_32883,N_31551,N_31179);
xnor U32884 (N_32884,N_31036,N_31935);
xor U32885 (N_32885,N_31626,N_31863);
nor U32886 (N_32886,N_31940,N_31884);
nand U32887 (N_32887,N_31661,N_31621);
nand U32888 (N_32888,N_31921,N_31664);
or U32889 (N_32889,N_31628,N_31680);
nor U32890 (N_32890,N_31748,N_31320);
nand U32891 (N_32891,N_31652,N_31528);
or U32892 (N_32892,N_31601,N_31793);
or U32893 (N_32893,N_31317,N_31517);
nor U32894 (N_32894,N_31208,N_31763);
or U32895 (N_32895,N_31185,N_31073);
and U32896 (N_32896,N_31734,N_31523);
and U32897 (N_32897,N_31994,N_31336);
xor U32898 (N_32898,N_31249,N_31602);
xnor U32899 (N_32899,N_31663,N_31742);
or U32900 (N_32900,N_31926,N_31478);
and U32901 (N_32901,N_31604,N_31351);
xnor U32902 (N_32902,N_31401,N_31188);
nand U32903 (N_32903,N_31613,N_31232);
or U32904 (N_32904,N_31049,N_31169);
or U32905 (N_32905,N_31477,N_31555);
nor U32906 (N_32906,N_31798,N_31926);
nor U32907 (N_32907,N_31203,N_31303);
or U32908 (N_32908,N_31202,N_31603);
or U32909 (N_32909,N_31779,N_31107);
xor U32910 (N_32910,N_31328,N_31311);
nand U32911 (N_32911,N_31285,N_31296);
nor U32912 (N_32912,N_31440,N_31739);
or U32913 (N_32913,N_31219,N_31488);
or U32914 (N_32914,N_31726,N_31890);
nor U32915 (N_32915,N_31481,N_31531);
or U32916 (N_32916,N_31409,N_31403);
and U32917 (N_32917,N_31098,N_31864);
nand U32918 (N_32918,N_31274,N_31430);
or U32919 (N_32919,N_31089,N_31898);
or U32920 (N_32920,N_31383,N_31425);
and U32921 (N_32921,N_31964,N_31832);
xor U32922 (N_32922,N_31817,N_31018);
xor U32923 (N_32923,N_31617,N_31408);
xor U32924 (N_32924,N_31199,N_31067);
xnor U32925 (N_32925,N_31445,N_31523);
nor U32926 (N_32926,N_31715,N_31862);
or U32927 (N_32927,N_31611,N_31675);
nand U32928 (N_32928,N_31479,N_31338);
nand U32929 (N_32929,N_31409,N_31582);
nand U32930 (N_32930,N_31604,N_31812);
or U32931 (N_32931,N_31545,N_31492);
nor U32932 (N_32932,N_31906,N_31688);
nand U32933 (N_32933,N_31212,N_31614);
nor U32934 (N_32934,N_31146,N_31919);
or U32935 (N_32935,N_31538,N_31610);
or U32936 (N_32936,N_31105,N_31290);
nor U32937 (N_32937,N_31213,N_31372);
nor U32938 (N_32938,N_31516,N_31125);
xor U32939 (N_32939,N_31497,N_31838);
xnor U32940 (N_32940,N_31446,N_31402);
nor U32941 (N_32941,N_31404,N_31014);
or U32942 (N_32942,N_31748,N_31570);
xor U32943 (N_32943,N_31595,N_31176);
and U32944 (N_32944,N_31305,N_31432);
and U32945 (N_32945,N_31424,N_31748);
or U32946 (N_32946,N_31073,N_31075);
xor U32947 (N_32947,N_31480,N_31115);
nand U32948 (N_32948,N_31630,N_31878);
or U32949 (N_32949,N_31589,N_31915);
and U32950 (N_32950,N_31440,N_31237);
and U32951 (N_32951,N_31207,N_31545);
nand U32952 (N_32952,N_31613,N_31452);
nor U32953 (N_32953,N_31074,N_31189);
nand U32954 (N_32954,N_31700,N_31578);
and U32955 (N_32955,N_31680,N_31911);
or U32956 (N_32956,N_31820,N_31859);
xor U32957 (N_32957,N_31910,N_31654);
and U32958 (N_32958,N_31131,N_31232);
nor U32959 (N_32959,N_31800,N_31149);
xnor U32960 (N_32960,N_31632,N_31558);
nor U32961 (N_32961,N_31113,N_31227);
or U32962 (N_32962,N_31008,N_31218);
or U32963 (N_32963,N_31087,N_31552);
and U32964 (N_32964,N_31439,N_31179);
xor U32965 (N_32965,N_31433,N_31640);
and U32966 (N_32966,N_31063,N_31194);
nor U32967 (N_32967,N_31933,N_31617);
and U32968 (N_32968,N_31679,N_31335);
and U32969 (N_32969,N_31255,N_31830);
nor U32970 (N_32970,N_31914,N_31915);
xor U32971 (N_32971,N_31769,N_31040);
xor U32972 (N_32972,N_31484,N_31363);
and U32973 (N_32973,N_31495,N_31668);
and U32974 (N_32974,N_31390,N_31739);
nand U32975 (N_32975,N_31430,N_31143);
xor U32976 (N_32976,N_31362,N_31165);
nor U32977 (N_32977,N_31652,N_31273);
nand U32978 (N_32978,N_31457,N_31636);
nor U32979 (N_32979,N_31338,N_31744);
xnor U32980 (N_32980,N_31360,N_31601);
nand U32981 (N_32981,N_31662,N_31751);
or U32982 (N_32982,N_31050,N_31347);
or U32983 (N_32983,N_31215,N_31892);
or U32984 (N_32984,N_31360,N_31180);
or U32985 (N_32985,N_31607,N_31140);
and U32986 (N_32986,N_31463,N_31231);
nor U32987 (N_32987,N_31114,N_31041);
or U32988 (N_32988,N_31915,N_31177);
nor U32989 (N_32989,N_31884,N_31497);
xnor U32990 (N_32990,N_31950,N_31968);
nor U32991 (N_32991,N_31335,N_31233);
nor U32992 (N_32992,N_31045,N_31808);
or U32993 (N_32993,N_31568,N_31660);
nor U32994 (N_32994,N_31825,N_31108);
and U32995 (N_32995,N_31870,N_31410);
and U32996 (N_32996,N_31140,N_31294);
nand U32997 (N_32997,N_31270,N_31945);
or U32998 (N_32998,N_31170,N_31646);
or U32999 (N_32999,N_31665,N_31640);
xnor U33000 (N_33000,N_32097,N_32863);
nor U33001 (N_33001,N_32968,N_32534);
xnor U33002 (N_33002,N_32342,N_32159);
and U33003 (N_33003,N_32796,N_32565);
nand U33004 (N_33004,N_32024,N_32588);
nand U33005 (N_33005,N_32561,N_32013);
or U33006 (N_33006,N_32734,N_32022);
xor U33007 (N_33007,N_32877,N_32261);
nor U33008 (N_33008,N_32800,N_32209);
nand U33009 (N_33009,N_32300,N_32569);
and U33010 (N_33010,N_32179,N_32089);
nor U33011 (N_33011,N_32496,N_32702);
nor U33012 (N_33012,N_32416,N_32350);
nand U33013 (N_33013,N_32180,N_32079);
nor U33014 (N_33014,N_32033,N_32436);
and U33015 (N_33015,N_32012,N_32239);
xnor U33016 (N_33016,N_32622,N_32509);
or U33017 (N_33017,N_32462,N_32156);
or U33018 (N_33018,N_32113,N_32754);
nor U33019 (N_33019,N_32882,N_32065);
xor U33020 (N_33020,N_32211,N_32521);
and U33021 (N_33021,N_32658,N_32711);
and U33022 (N_33022,N_32267,N_32452);
nand U33023 (N_33023,N_32178,N_32590);
or U33024 (N_33024,N_32422,N_32653);
nor U33025 (N_33025,N_32373,N_32834);
and U33026 (N_33026,N_32652,N_32666);
nand U33027 (N_33027,N_32369,N_32963);
xnor U33028 (N_33028,N_32837,N_32070);
or U33029 (N_33029,N_32096,N_32895);
or U33030 (N_33030,N_32778,N_32101);
nand U33031 (N_33031,N_32829,N_32680);
nand U33032 (N_33032,N_32134,N_32400);
nand U33033 (N_33033,N_32655,N_32981);
nand U33034 (N_33034,N_32913,N_32689);
nor U33035 (N_33035,N_32579,N_32757);
or U33036 (N_33036,N_32459,N_32606);
nor U33037 (N_33037,N_32930,N_32463);
or U33038 (N_33038,N_32679,N_32911);
and U33039 (N_33039,N_32885,N_32811);
or U33040 (N_33040,N_32087,N_32292);
or U33041 (N_33041,N_32784,N_32036);
nor U33042 (N_33042,N_32944,N_32009);
nand U33043 (N_33043,N_32061,N_32765);
xor U33044 (N_33044,N_32493,N_32368);
or U33045 (N_33045,N_32248,N_32171);
xnor U33046 (N_33046,N_32219,N_32257);
nor U33047 (N_33047,N_32490,N_32827);
and U33048 (N_33048,N_32527,N_32254);
xor U33049 (N_33049,N_32978,N_32724);
nor U33050 (N_33050,N_32224,N_32010);
or U33051 (N_33051,N_32716,N_32105);
nor U33052 (N_33052,N_32767,N_32624);
nand U33053 (N_33053,N_32130,N_32423);
xnor U33054 (N_33054,N_32327,N_32318);
and U33055 (N_33055,N_32456,N_32903);
nand U33056 (N_33056,N_32603,N_32011);
nand U33057 (N_33057,N_32642,N_32235);
and U33058 (N_33058,N_32104,N_32917);
xor U33059 (N_33059,N_32667,N_32578);
or U33060 (N_33060,N_32934,N_32390);
or U33061 (N_33061,N_32382,N_32234);
and U33062 (N_33062,N_32512,N_32501);
nor U33063 (N_33063,N_32779,N_32646);
xnor U33064 (N_33064,N_32564,N_32393);
nor U33065 (N_33065,N_32976,N_32277);
nand U33066 (N_33066,N_32682,N_32684);
or U33067 (N_33067,N_32537,N_32006);
nand U33068 (N_33068,N_32676,N_32242);
nor U33069 (N_33069,N_32320,N_32799);
nor U33070 (N_33070,N_32983,N_32957);
nor U33071 (N_33071,N_32357,N_32835);
nand U33072 (N_33072,N_32214,N_32019);
nand U33073 (N_33073,N_32819,N_32973);
and U33074 (N_33074,N_32795,N_32056);
nand U33075 (N_33075,N_32952,N_32084);
and U33076 (N_33076,N_32741,N_32344);
xnor U33077 (N_33077,N_32748,N_32516);
or U33078 (N_33078,N_32420,N_32632);
or U33079 (N_33079,N_32558,N_32458);
xor U33080 (N_33080,N_32678,N_32181);
nand U33081 (N_33081,N_32455,N_32439);
xnor U33082 (N_33082,N_32683,N_32886);
xnor U33083 (N_33083,N_32897,N_32773);
or U33084 (N_33084,N_32151,N_32189);
and U33085 (N_33085,N_32645,N_32958);
or U33086 (N_33086,N_32876,N_32383);
xnor U33087 (N_33087,N_32836,N_32172);
or U33088 (N_33088,N_32777,N_32494);
and U33089 (N_33089,N_32208,N_32807);
nor U33090 (N_33090,N_32194,N_32585);
nor U33091 (N_33091,N_32291,N_32128);
xnor U33092 (N_33092,N_32062,N_32788);
and U33093 (N_33093,N_32607,N_32285);
or U33094 (N_33094,N_32020,N_32939);
nand U33095 (N_33095,N_32095,N_32129);
nor U33096 (N_33096,N_32117,N_32007);
nor U33097 (N_33097,N_32774,N_32551);
nand U33098 (N_33098,N_32058,N_32999);
or U33099 (N_33099,N_32449,N_32766);
or U33100 (N_33100,N_32805,N_32677);
nor U33101 (N_33101,N_32060,N_32814);
and U33102 (N_33102,N_32281,N_32563);
or U33103 (N_33103,N_32043,N_32136);
xor U33104 (N_33104,N_32916,N_32441);
xnor U33105 (N_33105,N_32987,N_32661);
nand U33106 (N_33106,N_32681,N_32207);
or U33107 (N_33107,N_32522,N_32185);
and U33108 (N_33108,N_32241,N_32370);
or U33109 (N_33109,N_32355,N_32953);
or U33110 (N_33110,N_32424,N_32586);
xnor U33111 (N_33111,N_32502,N_32665);
xnor U33112 (N_33112,N_32478,N_32099);
and U33113 (N_33113,N_32240,N_32595);
or U33114 (N_33114,N_32432,N_32845);
nor U33115 (N_33115,N_32638,N_32164);
or U33116 (N_33116,N_32121,N_32387);
xor U33117 (N_33117,N_32946,N_32896);
and U33118 (N_33118,N_32379,N_32830);
and U33119 (N_33119,N_32428,N_32206);
and U33120 (N_33120,N_32451,N_32878);
or U33121 (N_33121,N_32037,N_32046);
xnor U33122 (N_33122,N_32700,N_32321);
and U33123 (N_33123,N_32941,N_32336);
nor U33124 (N_33124,N_32995,N_32443);
and U33125 (N_33125,N_32786,N_32378);
nand U33126 (N_33126,N_32985,N_32950);
nor U33127 (N_33127,N_32054,N_32531);
and U33128 (N_33128,N_32940,N_32562);
and U33129 (N_33129,N_32278,N_32457);
xnor U33130 (N_33130,N_32971,N_32881);
nand U33131 (N_33131,N_32589,N_32312);
and U33132 (N_33132,N_32377,N_32488);
nor U33133 (N_33133,N_32334,N_32236);
xor U33134 (N_33134,N_32005,N_32102);
nor U33135 (N_33135,N_32801,N_32523);
xnor U33136 (N_33136,N_32053,N_32608);
nand U33137 (N_33137,N_32560,N_32447);
xor U33138 (N_33138,N_32686,N_32550);
nor U33139 (N_33139,N_32055,N_32988);
or U33140 (N_33140,N_32764,N_32044);
nor U33141 (N_33141,N_32962,N_32391);
xnor U33142 (N_33142,N_32574,N_32848);
nor U33143 (N_33143,N_32816,N_32361);
or U33144 (N_33144,N_32915,N_32631);
or U33145 (N_33145,N_32268,N_32310);
nand U33146 (N_33146,N_32229,N_32205);
nand U33147 (N_33147,N_32535,N_32749);
nor U33148 (N_33148,N_32854,N_32536);
or U33149 (N_33149,N_32402,N_32161);
nand U33150 (N_33150,N_32825,N_32354);
and U33151 (N_33151,N_32826,N_32228);
or U33152 (N_33152,N_32050,N_32620);
or U33153 (N_33153,N_32345,N_32153);
and U33154 (N_33154,N_32328,N_32704);
and U33155 (N_33155,N_32860,N_32448);
and U33156 (N_33156,N_32910,N_32954);
and U33157 (N_33157,N_32813,N_32601);
nor U33158 (N_33158,N_32571,N_32468);
nor U33159 (N_33159,N_32500,N_32162);
and U33160 (N_33160,N_32831,N_32873);
nor U33161 (N_33161,N_32026,N_32945);
nand U33162 (N_33162,N_32559,N_32049);
xor U33163 (N_33163,N_32371,N_32525);
or U33164 (N_33164,N_32635,N_32810);
nand U33165 (N_33165,N_32844,N_32906);
nand U33166 (N_33166,N_32992,N_32284);
nand U33167 (N_33167,N_32331,N_32028);
nand U33168 (N_33168,N_32489,N_32143);
nand U33169 (N_33169,N_32313,N_32991);
nand U33170 (N_33170,N_32637,N_32583);
and U33171 (N_33171,N_32904,N_32260);
and U33172 (N_33172,N_32444,N_32597);
or U33173 (N_33173,N_32707,N_32972);
nor U33174 (N_33174,N_32204,N_32727);
nor U33175 (N_33175,N_32141,N_32119);
and U33176 (N_33176,N_32406,N_32002);
xnor U33177 (N_33177,N_32004,N_32614);
and U33178 (N_33178,N_32879,N_32990);
nand U33179 (N_33179,N_32532,N_32581);
nor U33180 (N_33180,N_32710,N_32309);
nand U33181 (N_33181,N_32880,N_32446);
or U33182 (N_33182,N_32431,N_32644);
or U33183 (N_33183,N_32869,N_32437);
nor U33184 (N_33184,N_32576,N_32623);
or U33185 (N_33185,N_32027,N_32201);
nand U33186 (N_33186,N_32169,N_32127);
nor U33187 (N_33187,N_32744,N_32418);
xnor U33188 (N_33188,N_32762,N_32360);
nor U33189 (N_33189,N_32809,N_32388);
nand U33190 (N_33190,N_32654,N_32783);
xnor U33191 (N_33191,N_32469,N_32543);
or U33192 (N_33192,N_32615,N_32649);
and U33193 (N_33193,N_32158,N_32514);
or U33194 (N_33194,N_32289,N_32769);
nor U33195 (N_33195,N_32883,N_32346);
nand U33196 (N_33196,N_32924,N_32401);
nand U33197 (N_33197,N_32761,N_32376);
xnor U33198 (N_33198,N_32487,N_32131);
and U33199 (N_33199,N_32951,N_32326);
and U33200 (N_33200,N_32894,N_32605);
or U33201 (N_33201,N_32865,N_32887);
xnor U33202 (N_33202,N_32567,N_32392);
nand U33203 (N_33203,N_32789,N_32850);
nor U33204 (N_33204,N_32698,N_32071);
xnor U33205 (N_33205,N_32187,N_32621);
xor U33206 (N_33206,N_32948,N_32304);
nand U33207 (N_33207,N_32454,N_32057);
and U33208 (N_33208,N_32639,N_32465);
or U33209 (N_33209,N_32955,N_32301);
nor U33210 (N_33210,N_32529,N_32083);
xor U33211 (N_33211,N_32986,N_32513);
nand U33212 (N_33212,N_32023,N_32249);
and U33213 (N_33213,N_32902,N_32703);
nor U33214 (N_33214,N_32085,N_32504);
nand U33215 (N_33215,N_32855,N_32929);
nor U33216 (N_33216,N_32453,N_32045);
xor U33217 (N_33217,N_32386,N_32602);
or U33218 (N_33218,N_32627,N_32317);
and U33219 (N_33219,N_32619,N_32506);
xor U33220 (N_33220,N_32935,N_32440);
nor U33221 (N_33221,N_32450,N_32616);
nor U33222 (N_33222,N_32338,N_32419);
or U33223 (N_33223,N_32518,N_32195);
and U33224 (N_33224,N_32231,N_32372);
or U33225 (N_33225,N_32780,N_32862);
and U33226 (N_33226,N_32015,N_32146);
nor U33227 (N_33227,N_32928,N_32977);
and U33228 (N_33228,N_32110,N_32163);
nand U33229 (N_33229,N_32251,N_32899);
xnor U33230 (N_33230,N_32192,N_32688);
nand U33231 (N_33231,N_32442,N_32908);
xor U33232 (N_33232,N_32712,N_32395);
or U33233 (N_33233,N_32617,N_32174);
nor U33234 (N_33234,N_32706,N_32225);
or U33235 (N_33235,N_32467,N_32319);
nand U33236 (N_33236,N_32031,N_32429);
nor U33237 (N_33237,N_32167,N_32647);
and U33238 (N_33238,N_32330,N_32996);
nand U33239 (N_33239,N_32694,N_32259);
and U33240 (N_33240,N_32316,N_32651);
nand U33241 (N_33241,N_32549,N_32733);
xnor U33242 (N_33242,N_32818,N_32542);
or U33243 (N_33243,N_32598,N_32247);
and U33244 (N_33244,N_32152,N_32526);
and U33245 (N_33245,N_32286,N_32273);
or U33246 (N_33246,N_32112,N_32464);
xor U33247 (N_33247,N_32931,N_32255);
nand U33248 (N_33248,N_32979,N_32824);
nand U33249 (N_33249,N_32275,N_32108);
nor U33250 (N_33250,N_32220,N_32575);
nor U33251 (N_33251,N_32604,N_32756);
and U33252 (N_33252,N_32849,N_32507);
or U33253 (N_33253,N_32258,N_32466);
nor U33254 (N_33254,N_32923,N_32905);
or U33255 (N_33255,N_32040,N_32557);
or U33256 (N_33256,N_32287,N_32280);
nor U33257 (N_33257,N_32909,N_32546);
and U33258 (N_33258,N_32636,N_32611);
or U33259 (N_33259,N_32937,N_32759);
and U33260 (N_33260,N_32133,N_32864);
or U33261 (N_33261,N_32018,N_32785);
and U33262 (N_33262,N_32517,N_32212);
and U33263 (N_33263,N_32302,N_32486);
nand U33264 (N_33264,N_32182,N_32374);
xor U33265 (N_33265,N_32114,N_32891);
xnor U33266 (N_33266,N_32052,N_32751);
and U33267 (N_33267,N_32218,N_32592);
nand U33268 (N_33268,N_32365,N_32256);
and U33269 (N_33269,N_32746,N_32539);
xnor U33270 (N_33270,N_32723,N_32394);
and U33271 (N_33271,N_32520,N_32792);
nor U33272 (N_33272,N_32874,N_32403);
or U33273 (N_33273,N_32696,N_32599);
and U33274 (N_33274,N_32411,N_32397);
or U33275 (N_33275,N_32843,N_32772);
nor U33276 (N_33276,N_32970,N_32262);
and U33277 (N_33277,N_32483,N_32966);
nor U33278 (N_33278,N_32471,N_32687);
or U33279 (N_33279,N_32787,N_32884);
or U33280 (N_33280,N_32349,N_32739);
or U33281 (N_33281,N_32547,N_32352);
or U33282 (N_33282,N_32705,N_32719);
nand U33283 (N_33283,N_32570,N_32122);
and U33284 (N_33284,N_32125,N_32190);
and U33285 (N_33285,N_32495,N_32307);
xor U33286 (N_33286,N_32918,N_32137);
or U33287 (N_33287,N_32685,N_32842);
or U33288 (N_33288,N_32306,N_32035);
xnor U33289 (N_33289,N_32184,N_32409);
and U33290 (N_33290,N_32960,N_32399);
nor U33291 (N_33291,N_32069,N_32077);
or U33292 (N_33292,N_32794,N_32132);
xor U33293 (N_33293,N_32697,N_32771);
xor U33294 (N_33294,N_32237,N_32160);
nor U33295 (N_33295,N_32362,N_32434);
xnor U33296 (N_33296,N_32538,N_32690);
nand U33297 (N_33297,N_32491,N_32846);
and U33298 (N_33298,N_32124,N_32870);
or U33299 (N_33299,N_32815,N_32732);
xnor U33300 (N_33300,N_32822,N_32802);
nor U33301 (N_33301,N_32123,N_32485);
nand U33302 (N_33302,N_32294,N_32656);
xnor U33303 (N_33303,N_32691,N_32866);
xor U33304 (N_33304,N_32210,N_32149);
xnor U33305 (N_33305,N_32039,N_32295);
or U33306 (N_33306,N_32343,N_32366);
or U33307 (N_33307,N_32577,N_32817);
xnor U33308 (N_33308,N_32725,N_32568);
nor U33309 (N_33309,N_32367,N_32790);
nand U33310 (N_33310,N_32166,N_32282);
nand U33311 (N_33311,N_32092,N_32859);
xnor U33312 (N_33312,N_32750,N_32852);
nor U33313 (N_33313,N_32919,N_32139);
nand U33314 (N_33314,N_32264,N_32051);
and U33315 (N_33315,N_32969,N_32003);
nand U33316 (N_33316,N_32708,N_32072);
or U33317 (N_33317,N_32186,N_32821);
or U33318 (N_33318,N_32175,N_32322);
and U33319 (N_33319,N_32359,N_32250);
xor U33320 (N_33320,N_32662,N_32901);
nand U33321 (N_33321,N_32290,N_32329);
and U33322 (N_33322,N_32148,N_32157);
nor U33323 (N_33323,N_32276,N_32106);
nand U33324 (N_33324,N_32781,N_32417);
nand U33325 (N_33325,N_32433,N_32659);
nand U33326 (N_33326,N_32713,N_32073);
nand U33327 (N_33327,N_32410,N_32797);
or U33328 (N_33328,N_32385,N_32356);
and U33329 (N_33329,N_32857,N_32925);
nor U33330 (N_33330,N_32470,N_32090);
nor U33331 (N_33331,N_32657,N_32841);
nor U33332 (N_33332,N_32271,N_32381);
or U33333 (N_33333,N_32861,N_32492);
or U33334 (N_33334,N_32947,N_32580);
or U33335 (N_33335,N_32274,N_32311);
nor U33336 (N_33336,N_32519,N_32147);
or U33337 (N_33337,N_32279,N_32412);
nand U33338 (N_33338,N_32715,N_32445);
or U33339 (N_33339,N_32475,N_32804);
and U33340 (N_33340,N_32042,N_32135);
nand U33341 (N_33341,N_32803,N_32335);
and U33342 (N_33342,N_32303,N_32067);
and U33343 (N_33343,N_32872,N_32384);
or U33344 (N_33344,N_32484,N_32230);
nor U33345 (N_33345,N_32552,N_32118);
nand U33346 (N_33346,N_32650,N_32047);
nand U33347 (N_33347,N_32351,N_32100);
nand U33348 (N_33348,N_32223,N_32720);
or U33349 (N_33349,N_32183,N_32625);
and U33350 (N_33350,N_32613,N_32348);
nand U33351 (N_33351,N_32017,N_32964);
nand U33352 (N_33352,N_32956,N_32413);
or U33353 (N_33353,N_32408,N_32337);
and U33354 (N_33354,N_32503,N_32693);
nor U33355 (N_33355,N_32064,N_32730);
nor U33356 (N_33356,N_32221,N_32168);
or U33357 (N_33357,N_32188,N_32499);
and U33358 (N_33358,N_32907,N_32758);
nand U33359 (N_33359,N_32942,N_32669);
nand U33360 (N_33360,N_32847,N_32226);
nand U33361 (N_33361,N_32202,N_32199);
or U33362 (N_33362,N_32116,N_32460);
nand U33363 (N_33363,N_32528,N_32692);
and U33364 (N_33364,N_32200,N_32333);
nand U33365 (N_33365,N_32075,N_32269);
nor U33366 (N_33366,N_32890,N_32791);
nor U33367 (N_33367,N_32041,N_32480);
nor U33368 (N_33368,N_32497,N_32438);
nor U33369 (N_33369,N_32213,N_32640);
nand U33370 (N_33370,N_32283,N_32325);
nand U33371 (N_33371,N_32555,N_32430);
and U33372 (N_33372,N_32533,N_32670);
nand U33373 (N_33373,N_32612,N_32752);
xnor U33374 (N_33374,N_32427,N_32076);
and U33375 (N_33375,N_32556,N_32729);
or U33376 (N_33376,N_32980,N_32252);
and U33377 (N_33377,N_32144,N_32566);
and U33378 (N_33378,N_32341,N_32375);
xor U33379 (N_33379,N_32066,N_32093);
nor U33380 (N_33380,N_32435,N_32288);
or U33381 (N_33381,N_32296,N_32196);
nor U33382 (N_33382,N_32120,N_32695);
xnor U33383 (N_33383,N_32404,N_32782);
xor U33384 (N_33384,N_32000,N_32699);
or U33385 (N_33385,N_32554,N_32738);
nor U33386 (N_33386,N_32984,N_32889);
nand U33387 (N_33387,N_32634,N_32227);
xnor U33388 (N_33388,N_32912,N_32339);
xor U33389 (N_33389,N_32340,N_32898);
nor U33390 (N_33390,N_32840,N_32347);
xnor U33391 (N_33391,N_32609,N_32511);
nand U33392 (N_33392,N_32851,N_32820);
xnor U33393 (N_33393,N_32177,N_32936);
and U33394 (N_33394,N_32203,N_32736);
xor U33395 (N_33395,N_32993,N_32150);
nor U33396 (N_33396,N_32823,N_32610);
nand U33397 (N_33397,N_32932,N_32740);
and U33398 (N_33398,N_32743,N_32414);
or U33399 (N_33399,N_32776,N_32098);
xnor U33400 (N_33400,N_32775,N_32660);
nor U33401 (N_33401,N_32107,N_32596);
xnor U33402 (N_33402,N_32246,N_32505);
nor U33403 (N_33403,N_32173,N_32461);
nor U33404 (N_33404,N_32943,N_32998);
nand U33405 (N_33405,N_32474,N_32838);
nand U33406 (N_33406,N_32920,N_32216);
nand U33407 (N_33407,N_32008,N_32630);
xor U33408 (N_33408,N_32832,N_32308);
nor U33409 (N_33409,N_32938,N_32671);
or U33410 (N_33410,N_32191,N_32358);
nand U33411 (N_33411,N_32103,N_32197);
xnor U33412 (N_33412,N_32892,N_32868);
or U33413 (N_33413,N_32109,N_32270);
or U33414 (N_33414,N_32875,N_32315);
nor U33415 (N_33415,N_32591,N_32722);
and U33416 (N_33416,N_32798,N_32245);
nand U33417 (N_33417,N_32389,N_32297);
nor U33418 (N_33418,N_32324,N_32138);
nand U33419 (N_33419,N_32217,N_32545);
nor U33420 (N_33420,N_32298,N_32111);
or U33421 (N_33421,N_32553,N_32243);
nor U33422 (N_33422,N_32063,N_32673);
and U33423 (N_33423,N_32668,N_32415);
or U33424 (N_33424,N_32548,N_32232);
and U33425 (N_33425,N_32476,N_32222);
and U33426 (N_33426,N_32030,N_32082);
nor U33427 (N_33427,N_32305,N_32714);
and U33428 (N_33428,N_32155,N_32473);
and U33429 (N_33429,N_32426,N_32735);
xnor U33430 (N_33430,N_32094,N_32126);
nor U33431 (N_33431,N_32747,N_32989);
and U33432 (N_33432,N_32048,N_32994);
nor U33433 (N_33433,N_32115,N_32266);
nand U33434 (N_33434,N_32293,N_32481);
nor U33435 (N_33435,N_32643,N_32793);
and U33436 (N_33436,N_32663,N_32633);
nand U33437 (N_33437,N_32768,N_32080);
nor U33438 (N_33438,N_32353,N_32091);
xnor U33439 (N_33439,N_32038,N_32721);
and U33440 (N_33440,N_32472,N_32629);
or U33441 (N_33441,N_32997,N_32672);
xor U33442 (N_33442,N_32479,N_32407);
nor U33443 (N_33443,N_32701,N_32364);
nand U33444 (N_33444,N_32933,N_32573);
and U33445 (N_33445,N_32016,N_32626);
and U33446 (N_33446,N_32059,N_32272);
nor U33447 (N_33447,N_32215,N_32728);
or U33448 (N_33448,N_32021,N_32641);
nor U33449 (N_33449,N_32893,N_32584);
nand U33450 (N_33450,N_32165,N_32856);
and U33451 (N_33451,N_32753,N_32709);
or U33452 (N_33452,N_32198,N_32675);
xnor U33453 (N_33453,N_32142,N_32323);
nor U33454 (N_33454,N_32405,N_32806);
nand U33455 (N_33455,N_32032,N_32808);
and U33456 (N_33456,N_32025,N_32363);
and U33457 (N_33457,N_32594,N_32398);
nor U33458 (N_33458,N_32927,N_32648);
nor U33459 (N_33459,N_32593,N_32858);
and U33460 (N_33460,N_32068,N_32628);
and U33461 (N_33461,N_32541,N_32078);
nand U33462 (N_33462,N_32425,N_32742);
or U33463 (N_33463,N_32853,N_32745);
nor U33464 (N_33464,N_32034,N_32029);
nor U33465 (N_33465,N_32396,N_32014);
or U33466 (N_33466,N_32193,N_32074);
xnor U33467 (N_33467,N_32572,N_32828);
and U33468 (N_33468,N_32833,N_32154);
xnor U33469 (N_33469,N_32170,N_32770);
nor U33470 (N_33470,N_32524,N_32253);
nand U33471 (N_33471,N_32982,N_32763);
and U33472 (N_33472,N_32839,N_32674);
xnor U33473 (N_33473,N_32760,N_32332);
nand U33474 (N_33474,N_32508,N_32233);
or U33475 (N_33475,N_32140,N_32544);
nor U33476 (N_33476,N_32737,N_32145);
xor U33477 (N_33477,N_32421,N_32867);
and U33478 (N_33478,N_32926,N_32515);
xnor U33479 (N_33479,N_32482,N_32664);
or U33480 (N_33480,N_32081,N_32477);
nor U33481 (N_33481,N_32265,N_32176);
xnor U33482 (N_33482,N_32755,N_32961);
nor U33483 (N_33483,N_32299,N_32975);
nor U33484 (N_33484,N_32088,N_32921);
nand U33485 (N_33485,N_32812,N_32263);
nor U33486 (N_33486,N_32498,N_32726);
nand U33487 (N_33487,N_32582,N_32380);
and U33488 (N_33488,N_32974,N_32731);
xnor U33489 (N_33489,N_32718,N_32959);
xor U33490 (N_33490,N_32949,N_32900);
or U33491 (N_33491,N_32618,N_32965);
xnor U33492 (N_33492,N_32888,N_32244);
xnor U33493 (N_33493,N_32587,N_32001);
and U33494 (N_33494,N_32914,N_32540);
or U33495 (N_33495,N_32600,N_32086);
nand U33496 (N_33496,N_32530,N_32871);
nor U33497 (N_33497,N_32717,N_32314);
xnor U33498 (N_33498,N_32510,N_32967);
or U33499 (N_33499,N_32238,N_32922);
nand U33500 (N_33500,N_32005,N_32189);
or U33501 (N_33501,N_32818,N_32874);
nand U33502 (N_33502,N_32655,N_32860);
or U33503 (N_33503,N_32143,N_32826);
xnor U33504 (N_33504,N_32173,N_32402);
nor U33505 (N_33505,N_32914,N_32338);
xnor U33506 (N_33506,N_32234,N_32578);
nand U33507 (N_33507,N_32607,N_32292);
nand U33508 (N_33508,N_32783,N_32808);
nor U33509 (N_33509,N_32590,N_32830);
xnor U33510 (N_33510,N_32889,N_32246);
or U33511 (N_33511,N_32182,N_32236);
xnor U33512 (N_33512,N_32603,N_32048);
nand U33513 (N_33513,N_32738,N_32327);
nor U33514 (N_33514,N_32266,N_32672);
and U33515 (N_33515,N_32621,N_32818);
xnor U33516 (N_33516,N_32614,N_32833);
nand U33517 (N_33517,N_32432,N_32122);
or U33518 (N_33518,N_32589,N_32034);
and U33519 (N_33519,N_32823,N_32915);
nand U33520 (N_33520,N_32843,N_32347);
nand U33521 (N_33521,N_32765,N_32823);
or U33522 (N_33522,N_32995,N_32841);
or U33523 (N_33523,N_32692,N_32058);
or U33524 (N_33524,N_32019,N_32413);
nor U33525 (N_33525,N_32129,N_32187);
xnor U33526 (N_33526,N_32345,N_32980);
or U33527 (N_33527,N_32553,N_32414);
nand U33528 (N_33528,N_32572,N_32482);
or U33529 (N_33529,N_32471,N_32926);
nand U33530 (N_33530,N_32809,N_32968);
xnor U33531 (N_33531,N_32792,N_32691);
or U33532 (N_33532,N_32562,N_32788);
or U33533 (N_33533,N_32907,N_32105);
and U33534 (N_33534,N_32144,N_32595);
and U33535 (N_33535,N_32447,N_32195);
xor U33536 (N_33536,N_32029,N_32071);
and U33537 (N_33537,N_32013,N_32006);
xnor U33538 (N_33538,N_32677,N_32511);
xor U33539 (N_33539,N_32151,N_32660);
nor U33540 (N_33540,N_32020,N_32788);
xnor U33541 (N_33541,N_32429,N_32802);
xor U33542 (N_33542,N_32106,N_32778);
and U33543 (N_33543,N_32644,N_32859);
nor U33544 (N_33544,N_32284,N_32417);
nor U33545 (N_33545,N_32437,N_32638);
nor U33546 (N_33546,N_32707,N_32181);
xor U33547 (N_33547,N_32157,N_32612);
and U33548 (N_33548,N_32635,N_32280);
and U33549 (N_33549,N_32105,N_32264);
nor U33550 (N_33550,N_32809,N_32483);
and U33551 (N_33551,N_32332,N_32301);
nor U33552 (N_33552,N_32419,N_32543);
nor U33553 (N_33553,N_32934,N_32229);
or U33554 (N_33554,N_32324,N_32791);
and U33555 (N_33555,N_32001,N_32496);
and U33556 (N_33556,N_32925,N_32987);
nor U33557 (N_33557,N_32255,N_32038);
nand U33558 (N_33558,N_32601,N_32287);
xnor U33559 (N_33559,N_32744,N_32075);
nor U33560 (N_33560,N_32436,N_32632);
and U33561 (N_33561,N_32938,N_32021);
xor U33562 (N_33562,N_32195,N_32512);
nor U33563 (N_33563,N_32444,N_32373);
nand U33564 (N_33564,N_32903,N_32658);
or U33565 (N_33565,N_32780,N_32044);
or U33566 (N_33566,N_32825,N_32861);
nand U33567 (N_33567,N_32403,N_32439);
and U33568 (N_33568,N_32652,N_32793);
and U33569 (N_33569,N_32094,N_32967);
and U33570 (N_33570,N_32529,N_32507);
nand U33571 (N_33571,N_32169,N_32786);
and U33572 (N_33572,N_32750,N_32015);
or U33573 (N_33573,N_32448,N_32658);
and U33574 (N_33574,N_32395,N_32137);
or U33575 (N_33575,N_32796,N_32760);
and U33576 (N_33576,N_32150,N_32291);
and U33577 (N_33577,N_32818,N_32286);
and U33578 (N_33578,N_32811,N_32058);
xor U33579 (N_33579,N_32739,N_32789);
nand U33580 (N_33580,N_32757,N_32619);
nor U33581 (N_33581,N_32540,N_32963);
and U33582 (N_33582,N_32694,N_32775);
xnor U33583 (N_33583,N_32352,N_32916);
and U33584 (N_33584,N_32396,N_32710);
xnor U33585 (N_33585,N_32937,N_32041);
xor U33586 (N_33586,N_32841,N_32423);
xnor U33587 (N_33587,N_32759,N_32264);
and U33588 (N_33588,N_32081,N_32311);
xnor U33589 (N_33589,N_32409,N_32989);
xor U33590 (N_33590,N_32413,N_32614);
xor U33591 (N_33591,N_32561,N_32727);
or U33592 (N_33592,N_32068,N_32405);
xor U33593 (N_33593,N_32622,N_32406);
and U33594 (N_33594,N_32094,N_32403);
or U33595 (N_33595,N_32030,N_32822);
xor U33596 (N_33596,N_32029,N_32179);
nor U33597 (N_33597,N_32862,N_32459);
nor U33598 (N_33598,N_32921,N_32962);
or U33599 (N_33599,N_32360,N_32883);
or U33600 (N_33600,N_32023,N_32756);
or U33601 (N_33601,N_32836,N_32055);
xor U33602 (N_33602,N_32783,N_32844);
and U33603 (N_33603,N_32660,N_32473);
nand U33604 (N_33604,N_32772,N_32847);
or U33605 (N_33605,N_32218,N_32410);
and U33606 (N_33606,N_32949,N_32007);
and U33607 (N_33607,N_32450,N_32595);
xnor U33608 (N_33608,N_32086,N_32374);
nor U33609 (N_33609,N_32304,N_32995);
nand U33610 (N_33610,N_32341,N_32208);
or U33611 (N_33611,N_32539,N_32681);
or U33612 (N_33612,N_32930,N_32763);
nor U33613 (N_33613,N_32505,N_32709);
and U33614 (N_33614,N_32575,N_32844);
nor U33615 (N_33615,N_32961,N_32202);
nor U33616 (N_33616,N_32762,N_32236);
nor U33617 (N_33617,N_32149,N_32311);
nor U33618 (N_33618,N_32283,N_32868);
nand U33619 (N_33619,N_32068,N_32293);
and U33620 (N_33620,N_32257,N_32721);
nand U33621 (N_33621,N_32155,N_32369);
and U33622 (N_33622,N_32269,N_32969);
nand U33623 (N_33623,N_32784,N_32522);
xor U33624 (N_33624,N_32822,N_32775);
or U33625 (N_33625,N_32197,N_32484);
and U33626 (N_33626,N_32491,N_32972);
nand U33627 (N_33627,N_32087,N_32629);
and U33628 (N_33628,N_32334,N_32055);
or U33629 (N_33629,N_32041,N_32020);
or U33630 (N_33630,N_32617,N_32134);
xor U33631 (N_33631,N_32232,N_32886);
or U33632 (N_33632,N_32534,N_32777);
xor U33633 (N_33633,N_32778,N_32397);
nor U33634 (N_33634,N_32552,N_32938);
nor U33635 (N_33635,N_32778,N_32870);
nand U33636 (N_33636,N_32148,N_32832);
and U33637 (N_33637,N_32951,N_32369);
nand U33638 (N_33638,N_32614,N_32647);
and U33639 (N_33639,N_32069,N_32010);
nand U33640 (N_33640,N_32292,N_32504);
or U33641 (N_33641,N_32887,N_32604);
nor U33642 (N_33642,N_32273,N_32250);
and U33643 (N_33643,N_32077,N_32229);
nor U33644 (N_33644,N_32953,N_32565);
and U33645 (N_33645,N_32444,N_32639);
or U33646 (N_33646,N_32477,N_32953);
nand U33647 (N_33647,N_32209,N_32287);
nor U33648 (N_33648,N_32124,N_32022);
or U33649 (N_33649,N_32887,N_32239);
nand U33650 (N_33650,N_32718,N_32349);
nand U33651 (N_33651,N_32520,N_32834);
and U33652 (N_33652,N_32857,N_32247);
xnor U33653 (N_33653,N_32602,N_32516);
xor U33654 (N_33654,N_32840,N_32367);
nand U33655 (N_33655,N_32286,N_32936);
nor U33656 (N_33656,N_32561,N_32715);
or U33657 (N_33657,N_32189,N_32083);
xor U33658 (N_33658,N_32295,N_32656);
xor U33659 (N_33659,N_32763,N_32257);
nand U33660 (N_33660,N_32867,N_32295);
xor U33661 (N_33661,N_32386,N_32732);
nand U33662 (N_33662,N_32847,N_32871);
xor U33663 (N_33663,N_32569,N_32573);
nand U33664 (N_33664,N_32905,N_32769);
nand U33665 (N_33665,N_32178,N_32296);
and U33666 (N_33666,N_32265,N_32148);
and U33667 (N_33667,N_32283,N_32658);
nor U33668 (N_33668,N_32306,N_32577);
and U33669 (N_33669,N_32098,N_32062);
xor U33670 (N_33670,N_32841,N_32812);
nor U33671 (N_33671,N_32014,N_32526);
nor U33672 (N_33672,N_32878,N_32677);
xnor U33673 (N_33673,N_32893,N_32684);
or U33674 (N_33674,N_32369,N_32473);
xnor U33675 (N_33675,N_32019,N_32865);
xor U33676 (N_33676,N_32318,N_32953);
nand U33677 (N_33677,N_32141,N_32983);
nand U33678 (N_33678,N_32381,N_32123);
xnor U33679 (N_33679,N_32176,N_32248);
nor U33680 (N_33680,N_32712,N_32056);
and U33681 (N_33681,N_32000,N_32857);
nor U33682 (N_33682,N_32108,N_32258);
nor U33683 (N_33683,N_32448,N_32959);
xnor U33684 (N_33684,N_32364,N_32946);
or U33685 (N_33685,N_32785,N_32868);
or U33686 (N_33686,N_32898,N_32736);
and U33687 (N_33687,N_32039,N_32956);
nand U33688 (N_33688,N_32022,N_32950);
and U33689 (N_33689,N_32878,N_32786);
nor U33690 (N_33690,N_32614,N_32900);
xnor U33691 (N_33691,N_32760,N_32914);
nand U33692 (N_33692,N_32932,N_32100);
and U33693 (N_33693,N_32422,N_32888);
and U33694 (N_33694,N_32005,N_32651);
nand U33695 (N_33695,N_32027,N_32803);
or U33696 (N_33696,N_32785,N_32528);
nor U33697 (N_33697,N_32598,N_32191);
or U33698 (N_33698,N_32730,N_32898);
nor U33699 (N_33699,N_32283,N_32528);
and U33700 (N_33700,N_32457,N_32537);
nor U33701 (N_33701,N_32583,N_32735);
nand U33702 (N_33702,N_32664,N_32936);
nand U33703 (N_33703,N_32002,N_32753);
xnor U33704 (N_33704,N_32733,N_32727);
nor U33705 (N_33705,N_32355,N_32331);
xnor U33706 (N_33706,N_32509,N_32847);
nand U33707 (N_33707,N_32054,N_32255);
nor U33708 (N_33708,N_32914,N_32762);
and U33709 (N_33709,N_32310,N_32072);
nor U33710 (N_33710,N_32260,N_32843);
xnor U33711 (N_33711,N_32051,N_32038);
nand U33712 (N_33712,N_32047,N_32894);
xnor U33713 (N_33713,N_32852,N_32114);
or U33714 (N_33714,N_32198,N_32348);
nor U33715 (N_33715,N_32215,N_32645);
xor U33716 (N_33716,N_32521,N_32787);
xor U33717 (N_33717,N_32977,N_32072);
or U33718 (N_33718,N_32054,N_32093);
nor U33719 (N_33719,N_32262,N_32502);
xnor U33720 (N_33720,N_32907,N_32378);
nand U33721 (N_33721,N_32283,N_32909);
and U33722 (N_33722,N_32699,N_32960);
or U33723 (N_33723,N_32974,N_32863);
xnor U33724 (N_33724,N_32934,N_32193);
or U33725 (N_33725,N_32762,N_32727);
xor U33726 (N_33726,N_32119,N_32201);
xor U33727 (N_33727,N_32324,N_32001);
nor U33728 (N_33728,N_32299,N_32907);
or U33729 (N_33729,N_32918,N_32469);
xor U33730 (N_33730,N_32115,N_32087);
or U33731 (N_33731,N_32225,N_32890);
xor U33732 (N_33732,N_32012,N_32667);
nand U33733 (N_33733,N_32606,N_32925);
and U33734 (N_33734,N_32041,N_32921);
xnor U33735 (N_33735,N_32163,N_32254);
xor U33736 (N_33736,N_32597,N_32138);
nor U33737 (N_33737,N_32550,N_32301);
nor U33738 (N_33738,N_32703,N_32828);
and U33739 (N_33739,N_32465,N_32627);
xnor U33740 (N_33740,N_32652,N_32401);
nand U33741 (N_33741,N_32870,N_32754);
or U33742 (N_33742,N_32609,N_32289);
or U33743 (N_33743,N_32640,N_32511);
or U33744 (N_33744,N_32375,N_32818);
nor U33745 (N_33745,N_32277,N_32041);
xnor U33746 (N_33746,N_32063,N_32779);
nand U33747 (N_33747,N_32173,N_32437);
nand U33748 (N_33748,N_32836,N_32126);
xnor U33749 (N_33749,N_32549,N_32403);
nor U33750 (N_33750,N_32579,N_32073);
nor U33751 (N_33751,N_32814,N_32192);
and U33752 (N_33752,N_32639,N_32747);
nand U33753 (N_33753,N_32843,N_32054);
and U33754 (N_33754,N_32734,N_32258);
nor U33755 (N_33755,N_32950,N_32627);
and U33756 (N_33756,N_32912,N_32278);
nand U33757 (N_33757,N_32726,N_32040);
or U33758 (N_33758,N_32992,N_32098);
and U33759 (N_33759,N_32056,N_32543);
or U33760 (N_33760,N_32995,N_32497);
or U33761 (N_33761,N_32636,N_32146);
and U33762 (N_33762,N_32432,N_32657);
nand U33763 (N_33763,N_32191,N_32425);
xnor U33764 (N_33764,N_32302,N_32839);
nor U33765 (N_33765,N_32211,N_32179);
xor U33766 (N_33766,N_32228,N_32052);
xnor U33767 (N_33767,N_32550,N_32383);
xnor U33768 (N_33768,N_32784,N_32349);
or U33769 (N_33769,N_32977,N_32505);
or U33770 (N_33770,N_32326,N_32578);
and U33771 (N_33771,N_32253,N_32289);
and U33772 (N_33772,N_32194,N_32920);
or U33773 (N_33773,N_32290,N_32923);
nor U33774 (N_33774,N_32155,N_32937);
xor U33775 (N_33775,N_32053,N_32030);
xnor U33776 (N_33776,N_32893,N_32054);
nor U33777 (N_33777,N_32602,N_32995);
nor U33778 (N_33778,N_32079,N_32947);
nor U33779 (N_33779,N_32061,N_32025);
or U33780 (N_33780,N_32816,N_32295);
or U33781 (N_33781,N_32267,N_32121);
and U33782 (N_33782,N_32538,N_32770);
nor U33783 (N_33783,N_32882,N_32436);
xnor U33784 (N_33784,N_32423,N_32288);
nor U33785 (N_33785,N_32524,N_32927);
xnor U33786 (N_33786,N_32641,N_32554);
xnor U33787 (N_33787,N_32476,N_32957);
nand U33788 (N_33788,N_32807,N_32341);
or U33789 (N_33789,N_32412,N_32911);
nor U33790 (N_33790,N_32153,N_32530);
or U33791 (N_33791,N_32516,N_32004);
and U33792 (N_33792,N_32646,N_32240);
xnor U33793 (N_33793,N_32387,N_32180);
xor U33794 (N_33794,N_32373,N_32454);
xor U33795 (N_33795,N_32710,N_32462);
or U33796 (N_33796,N_32864,N_32340);
xor U33797 (N_33797,N_32738,N_32667);
nor U33798 (N_33798,N_32632,N_32368);
nand U33799 (N_33799,N_32714,N_32485);
nand U33800 (N_33800,N_32034,N_32639);
or U33801 (N_33801,N_32605,N_32882);
and U33802 (N_33802,N_32165,N_32818);
nand U33803 (N_33803,N_32689,N_32817);
and U33804 (N_33804,N_32799,N_32445);
nor U33805 (N_33805,N_32535,N_32654);
and U33806 (N_33806,N_32341,N_32336);
or U33807 (N_33807,N_32141,N_32558);
and U33808 (N_33808,N_32259,N_32402);
nand U33809 (N_33809,N_32640,N_32830);
nand U33810 (N_33810,N_32655,N_32946);
xor U33811 (N_33811,N_32593,N_32229);
nand U33812 (N_33812,N_32049,N_32560);
or U33813 (N_33813,N_32570,N_32091);
and U33814 (N_33814,N_32446,N_32492);
nand U33815 (N_33815,N_32571,N_32831);
nor U33816 (N_33816,N_32527,N_32759);
and U33817 (N_33817,N_32494,N_32744);
nor U33818 (N_33818,N_32141,N_32603);
xor U33819 (N_33819,N_32134,N_32713);
or U33820 (N_33820,N_32278,N_32011);
and U33821 (N_33821,N_32616,N_32798);
or U33822 (N_33822,N_32073,N_32164);
and U33823 (N_33823,N_32017,N_32526);
nand U33824 (N_33824,N_32872,N_32662);
xnor U33825 (N_33825,N_32082,N_32247);
or U33826 (N_33826,N_32157,N_32545);
or U33827 (N_33827,N_32795,N_32540);
or U33828 (N_33828,N_32297,N_32242);
or U33829 (N_33829,N_32522,N_32745);
xor U33830 (N_33830,N_32597,N_32354);
nand U33831 (N_33831,N_32615,N_32375);
and U33832 (N_33832,N_32151,N_32004);
xor U33833 (N_33833,N_32170,N_32488);
nand U33834 (N_33834,N_32625,N_32084);
nor U33835 (N_33835,N_32303,N_32148);
xnor U33836 (N_33836,N_32329,N_32416);
or U33837 (N_33837,N_32570,N_32550);
nand U33838 (N_33838,N_32618,N_32883);
or U33839 (N_33839,N_32958,N_32368);
xor U33840 (N_33840,N_32575,N_32426);
nor U33841 (N_33841,N_32163,N_32922);
xnor U33842 (N_33842,N_32252,N_32018);
or U33843 (N_33843,N_32625,N_32522);
and U33844 (N_33844,N_32027,N_32272);
nor U33845 (N_33845,N_32558,N_32908);
or U33846 (N_33846,N_32027,N_32332);
and U33847 (N_33847,N_32533,N_32967);
or U33848 (N_33848,N_32909,N_32307);
nand U33849 (N_33849,N_32248,N_32206);
nor U33850 (N_33850,N_32772,N_32373);
and U33851 (N_33851,N_32911,N_32318);
and U33852 (N_33852,N_32328,N_32471);
nand U33853 (N_33853,N_32898,N_32375);
or U33854 (N_33854,N_32548,N_32879);
and U33855 (N_33855,N_32181,N_32119);
nor U33856 (N_33856,N_32164,N_32913);
and U33857 (N_33857,N_32731,N_32424);
or U33858 (N_33858,N_32499,N_32818);
or U33859 (N_33859,N_32693,N_32006);
nand U33860 (N_33860,N_32529,N_32221);
xnor U33861 (N_33861,N_32684,N_32016);
xnor U33862 (N_33862,N_32807,N_32648);
and U33863 (N_33863,N_32821,N_32307);
nor U33864 (N_33864,N_32277,N_32470);
or U33865 (N_33865,N_32692,N_32110);
or U33866 (N_33866,N_32923,N_32991);
or U33867 (N_33867,N_32163,N_32661);
nand U33868 (N_33868,N_32692,N_32756);
nor U33869 (N_33869,N_32744,N_32259);
xnor U33870 (N_33870,N_32895,N_32004);
xor U33871 (N_33871,N_32182,N_32515);
and U33872 (N_33872,N_32771,N_32455);
xnor U33873 (N_33873,N_32947,N_32060);
nand U33874 (N_33874,N_32094,N_32163);
nor U33875 (N_33875,N_32125,N_32295);
nand U33876 (N_33876,N_32083,N_32517);
xor U33877 (N_33877,N_32738,N_32254);
nand U33878 (N_33878,N_32739,N_32308);
nor U33879 (N_33879,N_32363,N_32395);
and U33880 (N_33880,N_32215,N_32882);
xnor U33881 (N_33881,N_32148,N_32105);
nor U33882 (N_33882,N_32657,N_32593);
or U33883 (N_33883,N_32595,N_32948);
nor U33884 (N_33884,N_32659,N_32697);
and U33885 (N_33885,N_32303,N_32863);
nand U33886 (N_33886,N_32619,N_32013);
xor U33887 (N_33887,N_32512,N_32910);
nand U33888 (N_33888,N_32372,N_32344);
nor U33889 (N_33889,N_32036,N_32748);
or U33890 (N_33890,N_32341,N_32621);
nor U33891 (N_33891,N_32521,N_32014);
nor U33892 (N_33892,N_32732,N_32882);
nand U33893 (N_33893,N_32972,N_32687);
nor U33894 (N_33894,N_32324,N_32111);
nor U33895 (N_33895,N_32673,N_32902);
xnor U33896 (N_33896,N_32238,N_32134);
nand U33897 (N_33897,N_32452,N_32552);
xnor U33898 (N_33898,N_32897,N_32444);
xnor U33899 (N_33899,N_32226,N_32082);
xor U33900 (N_33900,N_32061,N_32290);
nor U33901 (N_33901,N_32888,N_32068);
nand U33902 (N_33902,N_32870,N_32081);
or U33903 (N_33903,N_32630,N_32402);
and U33904 (N_33904,N_32195,N_32046);
xnor U33905 (N_33905,N_32007,N_32412);
nand U33906 (N_33906,N_32296,N_32179);
nand U33907 (N_33907,N_32969,N_32827);
nand U33908 (N_33908,N_32901,N_32620);
or U33909 (N_33909,N_32568,N_32736);
xor U33910 (N_33910,N_32832,N_32605);
nand U33911 (N_33911,N_32558,N_32640);
xor U33912 (N_33912,N_32016,N_32187);
xor U33913 (N_33913,N_32504,N_32794);
or U33914 (N_33914,N_32937,N_32785);
xor U33915 (N_33915,N_32309,N_32687);
or U33916 (N_33916,N_32355,N_32745);
nor U33917 (N_33917,N_32993,N_32522);
or U33918 (N_33918,N_32044,N_32809);
xor U33919 (N_33919,N_32188,N_32047);
xnor U33920 (N_33920,N_32096,N_32925);
and U33921 (N_33921,N_32870,N_32619);
or U33922 (N_33922,N_32007,N_32017);
and U33923 (N_33923,N_32824,N_32089);
nor U33924 (N_33924,N_32826,N_32554);
nand U33925 (N_33925,N_32148,N_32005);
nand U33926 (N_33926,N_32069,N_32937);
or U33927 (N_33927,N_32652,N_32703);
nand U33928 (N_33928,N_32274,N_32437);
and U33929 (N_33929,N_32387,N_32891);
xor U33930 (N_33930,N_32356,N_32047);
xnor U33931 (N_33931,N_32198,N_32191);
nand U33932 (N_33932,N_32923,N_32037);
and U33933 (N_33933,N_32073,N_32729);
and U33934 (N_33934,N_32380,N_32800);
xor U33935 (N_33935,N_32580,N_32478);
and U33936 (N_33936,N_32010,N_32120);
and U33937 (N_33937,N_32237,N_32030);
nand U33938 (N_33938,N_32170,N_32061);
nand U33939 (N_33939,N_32871,N_32187);
or U33940 (N_33940,N_32168,N_32829);
nand U33941 (N_33941,N_32710,N_32268);
xnor U33942 (N_33942,N_32183,N_32098);
or U33943 (N_33943,N_32755,N_32173);
nand U33944 (N_33944,N_32706,N_32345);
nor U33945 (N_33945,N_32222,N_32372);
or U33946 (N_33946,N_32327,N_32564);
nand U33947 (N_33947,N_32942,N_32701);
or U33948 (N_33948,N_32979,N_32563);
nand U33949 (N_33949,N_32282,N_32690);
or U33950 (N_33950,N_32058,N_32690);
or U33951 (N_33951,N_32902,N_32186);
xnor U33952 (N_33952,N_32439,N_32188);
xnor U33953 (N_33953,N_32176,N_32228);
and U33954 (N_33954,N_32753,N_32445);
or U33955 (N_33955,N_32983,N_32865);
nand U33956 (N_33956,N_32246,N_32096);
nor U33957 (N_33957,N_32592,N_32579);
xnor U33958 (N_33958,N_32762,N_32055);
or U33959 (N_33959,N_32683,N_32522);
and U33960 (N_33960,N_32508,N_32290);
nor U33961 (N_33961,N_32322,N_32816);
or U33962 (N_33962,N_32608,N_32811);
or U33963 (N_33963,N_32713,N_32437);
and U33964 (N_33964,N_32741,N_32373);
nand U33965 (N_33965,N_32198,N_32742);
nor U33966 (N_33966,N_32213,N_32895);
or U33967 (N_33967,N_32063,N_32266);
or U33968 (N_33968,N_32856,N_32936);
nor U33969 (N_33969,N_32946,N_32218);
and U33970 (N_33970,N_32061,N_32367);
and U33971 (N_33971,N_32277,N_32104);
and U33972 (N_33972,N_32926,N_32767);
nand U33973 (N_33973,N_32286,N_32489);
nor U33974 (N_33974,N_32974,N_32119);
nand U33975 (N_33975,N_32921,N_32621);
nor U33976 (N_33976,N_32373,N_32342);
and U33977 (N_33977,N_32076,N_32986);
or U33978 (N_33978,N_32502,N_32286);
nor U33979 (N_33979,N_32245,N_32692);
and U33980 (N_33980,N_32987,N_32902);
xnor U33981 (N_33981,N_32454,N_32597);
or U33982 (N_33982,N_32700,N_32725);
nand U33983 (N_33983,N_32669,N_32248);
or U33984 (N_33984,N_32052,N_32721);
and U33985 (N_33985,N_32757,N_32898);
or U33986 (N_33986,N_32414,N_32309);
and U33987 (N_33987,N_32853,N_32385);
nor U33988 (N_33988,N_32882,N_32501);
nor U33989 (N_33989,N_32201,N_32572);
xor U33990 (N_33990,N_32220,N_32596);
xor U33991 (N_33991,N_32794,N_32220);
xor U33992 (N_33992,N_32758,N_32641);
xnor U33993 (N_33993,N_32431,N_32957);
or U33994 (N_33994,N_32351,N_32859);
nor U33995 (N_33995,N_32350,N_32920);
or U33996 (N_33996,N_32039,N_32474);
nor U33997 (N_33997,N_32882,N_32221);
and U33998 (N_33998,N_32078,N_32983);
nor U33999 (N_33999,N_32749,N_32811);
nor U34000 (N_34000,N_33918,N_33677);
and U34001 (N_34001,N_33049,N_33633);
nand U34002 (N_34002,N_33964,N_33330);
nor U34003 (N_34003,N_33016,N_33671);
nand U34004 (N_34004,N_33349,N_33515);
xor U34005 (N_34005,N_33422,N_33028);
nand U34006 (N_34006,N_33765,N_33818);
nor U34007 (N_34007,N_33407,N_33745);
xnor U34008 (N_34008,N_33113,N_33066);
or U34009 (N_34009,N_33210,N_33602);
nor U34010 (N_34010,N_33105,N_33891);
xor U34011 (N_34011,N_33548,N_33999);
and U34012 (N_34012,N_33547,N_33424);
or U34013 (N_34013,N_33325,N_33345);
nor U34014 (N_34014,N_33845,N_33592);
nand U34015 (N_34015,N_33796,N_33183);
nand U34016 (N_34016,N_33376,N_33271);
xor U34017 (N_34017,N_33153,N_33604);
nor U34018 (N_34018,N_33539,N_33543);
xor U34019 (N_34019,N_33550,N_33742);
or U34020 (N_34020,N_33162,N_33694);
xor U34021 (N_34021,N_33569,N_33738);
xor U34022 (N_34022,N_33004,N_33428);
and U34023 (N_34023,N_33626,N_33432);
or U34024 (N_34024,N_33879,N_33123);
xnor U34025 (N_34025,N_33563,N_33389);
or U34026 (N_34026,N_33333,N_33744);
or U34027 (N_34027,N_33199,N_33962);
nand U34028 (N_34028,N_33346,N_33926);
and U34029 (N_34029,N_33285,N_33963);
nand U34030 (N_34030,N_33202,N_33776);
and U34031 (N_34031,N_33924,N_33206);
nor U34032 (N_34032,N_33339,N_33618);
nor U34033 (N_34033,N_33807,N_33364);
nor U34034 (N_34034,N_33351,N_33949);
nand U34035 (N_34035,N_33248,N_33201);
or U34036 (N_34036,N_33075,N_33262);
xor U34037 (N_34037,N_33272,N_33519);
nand U34038 (N_34038,N_33590,N_33857);
nor U34039 (N_34039,N_33559,N_33220);
nor U34040 (N_34040,N_33239,N_33021);
and U34041 (N_34041,N_33043,N_33282);
nand U34042 (N_34042,N_33289,N_33082);
or U34043 (N_34043,N_33056,N_33001);
nand U34044 (N_34044,N_33521,N_33758);
xor U34045 (N_34045,N_33904,N_33959);
nor U34046 (N_34046,N_33967,N_33601);
nor U34047 (N_34047,N_33644,N_33275);
or U34048 (N_34048,N_33986,N_33646);
and U34049 (N_34049,N_33363,N_33840);
xnor U34050 (N_34050,N_33484,N_33546);
xor U34051 (N_34051,N_33495,N_33382);
and U34052 (N_34052,N_33794,N_33751);
nand U34053 (N_34053,N_33111,N_33232);
or U34054 (N_34054,N_33994,N_33178);
nor U34055 (N_34055,N_33498,N_33394);
and U34056 (N_34056,N_33425,N_33435);
nor U34057 (N_34057,N_33292,N_33603);
and U34058 (N_34058,N_33854,N_33576);
nor U34059 (N_34059,N_33231,N_33434);
xor U34060 (N_34060,N_33913,N_33561);
nor U34061 (N_34061,N_33530,N_33480);
xnor U34062 (N_34062,N_33409,N_33612);
xnor U34063 (N_34063,N_33290,N_33920);
or U34064 (N_34064,N_33761,N_33577);
and U34065 (N_34065,N_33851,N_33091);
nor U34066 (N_34066,N_33459,N_33584);
xnor U34067 (N_34067,N_33667,N_33130);
xor U34068 (N_34068,N_33946,N_33808);
xor U34069 (N_34069,N_33624,N_33786);
nand U34070 (N_34070,N_33483,N_33855);
and U34071 (N_34071,N_33979,N_33417);
xor U34072 (N_34072,N_33685,N_33412);
nand U34073 (N_34073,N_33340,N_33449);
nand U34074 (N_34074,N_33683,N_33391);
or U34075 (N_34075,N_33229,N_33439);
nand U34076 (N_34076,N_33031,N_33627);
xnor U34077 (N_34077,N_33570,N_33034);
nand U34078 (N_34078,N_33300,N_33128);
xor U34079 (N_34079,N_33771,N_33233);
xor U34080 (N_34080,N_33616,N_33810);
nand U34081 (N_34081,N_33063,N_33298);
or U34082 (N_34082,N_33898,N_33504);
or U34083 (N_34083,N_33752,N_33886);
and U34084 (N_34084,N_33143,N_33064);
and U34085 (N_34085,N_33940,N_33472);
nor U34086 (N_34086,N_33941,N_33301);
nand U34087 (N_34087,N_33370,N_33681);
xor U34088 (N_34088,N_33868,N_33112);
and U34089 (N_34089,N_33533,N_33676);
xor U34090 (N_34090,N_33910,N_33234);
xor U34091 (N_34091,N_33731,N_33485);
xnor U34092 (N_34092,N_33052,N_33534);
or U34093 (N_34093,N_33614,N_33238);
and U34094 (N_34094,N_33544,N_33867);
nand U34095 (N_34095,N_33838,N_33615);
nor U34096 (N_34096,N_33895,N_33585);
or U34097 (N_34097,N_33782,N_33426);
nor U34098 (N_34098,N_33286,N_33606);
and U34099 (N_34099,N_33400,N_33813);
and U34100 (N_34100,N_33702,N_33385);
and U34101 (N_34101,N_33227,N_33102);
nor U34102 (N_34102,N_33656,N_33295);
xor U34103 (N_34103,N_33541,N_33027);
nor U34104 (N_34104,N_33565,N_33674);
xnor U34105 (N_34105,N_33230,N_33655);
nor U34106 (N_34106,N_33287,N_33892);
nor U34107 (N_34107,N_33793,N_33323);
and U34108 (N_34108,N_33664,N_33324);
or U34109 (N_34109,N_33826,N_33416);
or U34110 (N_34110,N_33600,N_33133);
or U34111 (N_34111,N_33925,N_33988);
xor U34112 (N_34112,N_33200,N_33072);
nor U34113 (N_34113,N_33887,N_33155);
or U34114 (N_34114,N_33575,N_33019);
nand U34115 (N_34115,N_33890,N_33916);
nand U34116 (N_34116,N_33101,N_33780);
nor U34117 (N_34117,N_33739,N_33637);
nor U34118 (N_34118,N_33639,N_33799);
or U34119 (N_34119,N_33703,N_33184);
and U34120 (N_34120,N_33591,N_33823);
or U34121 (N_34121,N_33440,N_33724);
and U34122 (N_34122,N_33025,N_33088);
and U34123 (N_34123,N_33746,N_33938);
nor U34124 (N_34124,N_33093,N_33802);
nor U34125 (N_34125,N_33792,N_33454);
xor U34126 (N_34126,N_33023,N_33089);
and U34127 (N_34127,N_33937,N_33686);
nand U34128 (N_34128,N_33789,N_33402);
nor U34129 (N_34129,N_33649,N_33992);
or U34130 (N_34130,N_33573,N_33121);
nand U34131 (N_34131,N_33950,N_33073);
or U34132 (N_34132,N_33359,N_33452);
or U34133 (N_34133,N_33712,N_33215);
and U34134 (N_34134,N_33736,N_33000);
and U34135 (N_34135,N_33873,N_33623);
nor U34136 (N_34136,N_33120,N_33243);
nand U34137 (N_34137,N_33353,N_33368);
xnor U34138 (N_34138,N_33930,N_33993);
and U34139 (N_34139,N_33996,N_33722);
or U34140 (N_34140,N_33837,N_33074);
nor U34141 (N_34141,N_33817,N_33360);
nor U34142 (N_34142,N_33226,N_33866);
nor U34143 (N_34143,N_33247,N_33046);
nand U34144 (N_34144,N_33187,N_33862);
or U34145 (N_34145,N_33728,N_33874);
nor U34146 (N_34146,N_33136,N_33260);
or U34147 (N_34147,N_33321,N_33909);
or U34148 (N_34148,N_33085,N_33297);
and U34149 (N_34149,N_33284,N_33320);
nor U34150 (N_34150,N_33522,N_33582);
xor U34151 (N_34151,N_33291,N_33716);
xnor U34152 (N_34152,N_33939,N_33037);
and U34153 (N_34153,N_33228,N_33216);
and U34154 (N_34154,N_33645,N_33991);
or U34155 (N_34155,N_33399,N_33146);
nor U34156 (N_34156,N_33852,N_33707);
nand U34157 (N_34157,N_33159,N_33441);
xor U34158 (N_34158,N_33915,N_33198);
xnor U34159 (N_34159,N_33772,N_33878);
nor U34160 (N_34160,N_33138,N_33245);
or U34161 (N_34161,N_33068,N_33853);
or U34162 (N_34162,N_33192,N_33989);
xnor U34163 (N_34163,N_33740,N_33557);
and U34164 (N_34164,N_33331,N_33889);
xnor U34165 (N_34165,N_33486,N_33571);
nand U34166 (N_34166,N_33344,N_33847);
and U34167 (N_34167,N_33911,N_33379);
or U34168 (N_34168,N_33551,N_33457);
nor U34169 (N_34169,N_33362,N_33865);
and U34170 (N_34170,N_33475,N_33334);
xnor U34171 (N_34171,N_33191,N_33188);
and U34172 (N_34172,N_33065,N_33253);
and U34173 (N_34173,N_33846,N_33423);
and U34174 (N_34174,N_33901,N_33995);
nand U34175 (N_34175,N_33170,N_33815);
nand U34176 (N_34176,N_33476,N_33084);
nor U34177 (N_34177,N_33437,N_33811);
or U34178 (N_34178,N_33628,N_33270);
or U34179 (N_34179,N_33844,N_33505);
nor U34180 (N_34180,N_33756,N_33933);
nand U34181 (N_34181,N_33494,N_33003);
or U34182 (N_34182,N_33197,N_33668);
or U34183 (N_34183,N_33726,N_33491);
and U34184 (N_34184,N_33354,N_33643);
nand U34185 (N_34185,N_33971,N_33670);
xnor U34186 (N_34186,N_33587,N_33642);
nand U34187 (N_34187,N_33897,N_33833);
nand U34188 (N_34188,N_33473,N_33589);
nor U34189 (N_34189,N_33629,N_33666);
and U34190 (N_34190,N_33134,N_33438);
or U34191 (N_34191,N_33617,N_33358);
nand U34192 (N_34192,N_33267,N_33067);
or U34193 (N_34193,N_33467,N_33958);
and U34194 (N_34194,N_33990,N_33691);
nand U34195 (N_34195,N_33318,N_33393);
or U34196 (N_34196,N_33479,N_33599);
nand U34197 (N_34197,N_33211,N_33922);
and U34198 (N_34198,N_33319,N_33934);
nor U34199 (N_34199,N_33427,N_33302);
xor U34200 (N_34200,N_33875,N_33151);
xnor U34201 (N_34201,N_33970,N_33888);
xor U34202 (N_34202,N_33566,N_33489);
xor U34203 (N_34203,N_33263,N_33766);
nor U34204 (N_34204,N_33662,N_33415);
xor U34205 (N_34205,N_33809,N_33366);
nand U34206 (N_34206,N_33396,N_33255);
nand U34207 (N_34207,N_33715,N_33026);
nor U34208 (N_34208,N_33465,N_33721);
xor U34209 (N_34209,N_33125,N_33581);
nand U34210 (N_34210,N_33157,N_33163);
xnor U34211 (N_34211,N_33743,N_33169);
xor U34212 (N_34212,N_33687,N_33717);
nand U34213 (N_34213,N_33652,N_33160);
or U34214 (N_34214,N_33182,N_33098);
nand U34215 (N_34215,N_33387,N_33936);
and U34216 (N_34216,N_33311,N_33148);
nand U34217 (N_34217,N_33219,N_33347);
and U34218 (N_34218,N_33041,N_33947);
xor U34219 (N_34219,N_33012,N_33516);
nor U34220 (N_34220,N_33675,N_33542);
nor U34221 (N_34221,N_33558,N_33597);
nor U34222 (N_34222,N_33727,N_33132);
nor U34223 (N_34223,N_33078,N_33209);
nor U34224 (N_34224,N_33907,N_33100);
nor U34225 (N_34225,N_33326,N_33212);
or U34226 (N_34226,N_33790,N_33705);
xor U34227 (N_34227,N_33455,N_33981);
nor U34228 (N_34228,N_33880,N_33141);
nor U34229 (N_34229,N_33283,N_33832);
and U34230 (N_34230,N_33024,N_33835);
or U34231 (N_34231,N_33701,N_33147);
nor U34232 (N_34232,N_33378,N_33975);
xor U34233 (N_34233,N_33690,N_33395);
and U34234 (N_34234,N_33179,N_33256);
nand U34235 (N_34235,N_33777,N_33944);
and U34236 (N_34236,N_33729,N_33973);
or U34237 (N_34237,N_33638,N_33536);
xnor U34238 (N_34238,N_33116,N_33266);
xor U34239 (N_34239,N_33118,N_33713);
or U34240 (N_34240,N_33620,N_33696);
nor U34241 (N_34241,N_33942,N_33755);
nor U34242 (N_34242,N_33788,N_33337);
nand U34243 (N_34243,N_33404,N_33564);
nor U34244 (N_34244,N_33115,N_33816);
or U34245 (N_34245,N_33447,N_33493);
xor U34246 (N_34246,N_33278,N_33355);
xnor U34247 (N_34247,N_33175,N_33279);
nand U34248 (N_34248,N_33172,N_33044);
and U34249 (N_34249,N_33408,N_33509);
xnor U34250 (N_34250,N_33069,N_33842);
xnor U34251 (N_34251,N_33672,N_33369);
xnor U34252 (N_34252,N_33237,N_33131);
nand U34253 (N_34253,N_33635,N_33009);
nor U34254 (N_34254,N_33273,N_33831);
nor U34255 (N_34255,N_33503,N_33094);
nand U34256 (N_34256,N_33647,N_33919);
or U34257 (N_34257,N_33773,N_33525);
xnor U34258 (N_34258,N_33092,N_33135);
or U34259 (N_34259,N_33706,N_33126);
nand U34260 (N_34260,N_33429,N_33261);
xor U34261 (N_34261,N_33513,N_33748);
xnor U34262 (N_34262,N_33884,N_33660);
and U34263 (N_34263,N_33650,N_33735);
nand U34264 (N_34264,N_33673,N_33605);
and U34265 (N_34265,N_33552,N_33554);
and U34266 (N_34266,N_33806,N_33371);
nand U34267 (N_34267,N_33622,N_33312);
or U34268 (N_34268,N_33470,N_33572);
and U34269 (N_34269,N_33207,N_33532);
nor U34270 (N_34270,N_33288,N_33529);
nand U34271 (N_34271,N_33152,N_33444);
and U34272 (N_34272,N_33657,N_33974);
nand U34273 (N_34273,N_33787,N_33055);
or U34274 (N_34274,N_33882,N_33413);
nor U34275 (N_34275,N_33520,N_33692);
or U34276 (N_34276,N_33213,N_33960);
or U34277 (N_34277,N_33961,N_33313);
nor U34278 (N_34278,N_33246,N_33625);
or U34279 (N_34279,N_33418,N_33087);
nor U34280 (N_34280,N_33205,N_33167);
nor U34281 (N_34281,N_33537,N_33508);
or U34282 (N_34282,N_33972,N_33456);
nor U34283 (N_34283,N_33779,N_33051);
nand U34284 (N_34284,N_33850,N_33859);
nand U34285 (N_34285,N_33762,N_33086);
xor U34286 (N_34286,N_33952,N_33114);
nand U34287 (N_34287,N_33401,N_33708);
and U34288 (N_34288,N_33770,N_33540);
nor U34289 (N_34289,N_33871,N_33042);
and U34290 (N_34290,N_33471,N_33814);
nor U34291 (N_34291,N_33896,N_33985);
nand U34292 (N_34292,N_33836,N_33124);
nand U34293 (N_34293,N_33365,N_33388);
and U34294 (N_34294,N_33127,N_33678);
nor U34295 (N_34295,N_33805,N_33305);
xor U34296 (N_34296,N_33501,N_33406);
or U34297 (N_34297,N_33224,N_33593);
nor U34298 (N_34298,N_33461,N_33411);
nor U34299 (N_34299,N_33978,N_33140);
xor U34300 (N_34300,N_33142,N_33514);
nand U34301 (N_34301,N_33791,N_33478);
xnor U34302 (N_34302,N_33083,N_33653);
and U34303 (N_34303,N_33870,N_33299);
and U34304 (N_34304,N_33294,N_33214);
nand U34305 (N_34305,N_33883,N_33332);
xor U34306 (N_34306,N_33420,N_33020);
xor U34307 (N_34307,N_33502,N_33030);
or U34308 (N_34308,N_33372,N_33749);
nor U34309 (N_34309,N_33165,N_33906);
and U34310 (N_34310,N_33375,N_33518);
and U34311 (N_34311,N_33511,N_33714);
nand U34312 (N_34312,N_33450,N_33002);
or U34313 (N_34313,N_33442,N_33095);
and U34314 (N_34314,N_33171,N_33497);
nor U34315 (N_34315,N_33469,N_33193);
or U34316 (N_34316,N_33010,N_33586);
nand U34317 (N_34317,N_33381,N_33596);
nand U34318 (N_34318,N_33820,N_33562);
nand U34319 (N_34319,N_33829,N_33733);
and U34320 (N_34320,N_33512,N_33410);
or U34321 (N_34321,N_33693,N_33669);
or U34322 (N_34322,N_33061,N_33535);
nor U34323 (N_34323,N_33309,N_33352);
and U34324 (N_34324,N_33264,N_33968);
xor U34325 (N_34325,N_33338,N_33953);
nand U34326 (N_34326,N_33109,N_33296);
xor U34327 (N_34327,N_33980,N_33356);
nor U34328 (N_34328,N_33062,N_33481);
and U34329 (N_34329,N_33737,N_33161);
or U34330 (N_34330,N_33335,N_33734);
or U34331 (N_34331,N_33899,N_33506);
nor U34332 (N_34332,N_33058,N_33556);
and U34333 (N_34333,N_33553,N_33699);
nand U34334 (N_34334,N_33640,N_33242);
or U34335 (N_34335,N_33856,N_33760);
or U34336 (N_34336,N_33757,N_33704);
and U34337 (N_34337,N_33149,N_33900);
and U34338 (N_34338,N_33763,N_33250);
or U34339 (N_34339,N_33122,N_33386);
or U34340 (N_34340,N_33144,N_33059);
nand U34341 (N_34341,N_33306,N_33801);
xor U34342 (N_34342,N_33150,N_33327);
xnor U34343 (N_34343,N_33310,N_33583);
xnor U34344 (N_34344,N_33221,N_33579);
nand U34345 (N_34345,N_33057,N_33322);
nor U34346 (N_34346,N_33195,N_33164);
and U34347 (N_34347,N_33022,N_33613);
nand U34348 (N_34348,N_33824,N_33621);
nor U34349 (N_34349,N_33281,N_33076);
and U34350 (N_34350,N_33711,N_33464);
nor U34351 (N_34351,N_33307,N_33651);
nand U34352 (N_34352,N_33490,N_33194);
nor U34353 (N_34353,N_33080,N_33500);
nand U34354 (N_34354,N_33775,N_33398);
xor U34355 (N_34355,N_33252,N_33185);
xnor U34356 (N_34356,N_33797,N_33096);
nand U34357 (N_34357,N_33468,N_33610);
and U34358 (N_34358,N_33710,N_33357);
and U34359 (N_34359,N_33917,N_33181);
nor U34360 (N_34360,N_33090,N_33038);
or U34361 (N_34361,N_33106,N_33689);
and U34362 (N_34362,N_33017,N_33932);
nand U34363 (N_34363,N_33035,N_33463);
nor U34364 (N_34364,N_33316,N_33436);
or U34365 (N_34365,N_33720,N_33180);
nand U34366 (N_34366,N_33110,N_33951);
xnor U34367 (N_34367,N_33957,N_33222);
nor U34368 (N_34368,N_33033,N_33390);
xnor U34369 (N_34369,N_33048,N_33108);
xnor U34370 (N_34370,N_33821,N_33013);
nand U34371 (N_34371,N_33217,N_33658);
and U34372 (N_34372,N_33680,N_33166);
or U34373 (N_34373,N_33361,N_33902);
nand U34374 (N_34374,N_33257,N_33218);
nor U34375 (N_34375,N_33139,N_33608);
nand U34376 (N_34376,N_33014,N_33574);
and U34377 (N_34377,N_33036,N_33969);
and U34378 (N_34378,N_33905,N_33783);
and U34379 (N_34379,N_33236,N_33446);
xor U34380 (N_34380,N_33764,N_33631);
or U34381 (N_34381,N_33097,N_33377);
nor U34382 (N_34382,N_33661,N_33923);
or U34383 (N_34383,N_33158,N_33462);
nor U34384 (N_34384,N_33718,N_33825);
and U34385 (N_34385,N_33560,N_33196);
and U34386 (N_34386,N_33419,N_33948);
xor U34387 (N_34387,N_33168,N_33769);
xor U34388 (N_34388,N_33240,N_33040);
nor U34389 (N_34389,N_33881,N_33929);
or U34390 (N_34390,N_33156,N_33258);
xnor U34391 (N_34391,N_33741,N_33293);
xor U34392 (N_34392,N_33443,N_33914);
and U34393 (N_34393,N_33204,N_33137);
xnor U34394 (N_34394,N_33849,N_33528);
xnor U34395 (N_34395,N_33460,N_33695);
nor U34396 (N_34396,N_33119,N_33251);
and U34397 (N_34397,N_33145,N_33632);
and U34398 (N_34398,N_33943,N_33987);
xor U34399 (N_34399,N_33619,N_33594);
and U34400 (N_34400,N_33795,N_33877);
nor U34401 (N_34401,N_33965,N_33531);
nand U34402 (N_34402,N_33630,N_33208);
nand U34403 (N_34403,N_33397,N_33304);
nor U34404 (N_34404,N_33998,N_33774);
nand U34405 (N_34405,N_33079,N_33032);
xor U34406 (N_34406,N_33747,N_33567);
xnor U34407 (N_34407,N_33753,N_33235);
xor U34408 (N_34408,N_33578,N_33314);
nand U34409 (N_34409,N_33723,N_33798);
nand U34410 (N_34410,N_33011,N_33588);
or U34411 (N_34411,N_33822,N_33719);
and U34412 (N_34412,N_33081,N_33510);
nand U34413 (N_34413,N_33496,N_33894);
or U34414 (N_34414,N_33935,N_33474);
nand U34415 (N_34415,N_33329,N_33834);
and U34416 (N_34416,N_33104,N_33380);
xor U34417 (N_34417,N_33893,N_33342);
nor U34418 (N_34418,N_33308,N_33177);
xor U34419 (N_34419,N_33414,N_33580);
and U34420 (N_34420,N_33781,N_33280);
nand U34421 (N_34421,N_33254,N_33174);
or U34422 (N_34422,N_33538,N_33373);
xor U34423 (N_34423,N_33274,N_33863);
nor U34424 (N_34424,N_33977,N_33265);
xor U34425 (N_34425,N_33259,N_33008);
or U34426 (N_34426,N_33709,N_33595);
and U34427 (N_34427,N_33955,N_33315);
nand U34428 (N_34428,N_33350,N_33203);
and U34429 (N_34429,N_33830,N_33700);
xnor U34430 (N_34430,N_33527,N_33641);
xor U34431 (N_34431,N_33269,N_33730);
or U34432 (N_34432,N_33129,N_33956);
or U34433 (N_34433,N_33997,N_33054);
nor U34434 (N_34434,N_33827,N_33006);
and U34435 (N_34435,N_33050,N_33458);
or U34436 (N_34436,N_33249,N_33804);
xnor U34437 (N_34437,N_33445,N_33688);
or U34438 (N_34438,N_33732,N_33492);
or U34439 (N_34439,N_33405,N_33903);
nand U34440 (N_34440,N_33317,N_33908);
nor U34441 (N_34441,N_33384,N_33912);
or U34442 (N_34442,N_33698,N_33984);
nor U34443 (N_34443,N_33966,N_33403);
and U34444 (N_34444,N_33800,N_33117);
nand U34445 (N_34445,N_33099,N_33487);
xor U34446 (N_34446,N_33190,N_33103);
xnor U34447 (N_34447,N_33303,N_33348);
xor U34448 (N_34448,N_33682,N_33785);
nor U34449 (N_34449,N_33778,N_33931);
or U34450 (N_34450,N_33482,N_33018);
nor U34451 (N_34451,N_33665,N_33453);
and U34452 (N_34452,N_33598,N_33392);
nor U34453 (N_34453,N_33725,N_33869);
xnor U34454 (N_34454,N_33477,N_33431);
nand U34455 (N_34455,N_33039,N_33421);
and U34456 (N_34456,N_33611,N_33374);
and U34457 (N_34457,N_33872,N_33225);
xor U34458 (N_34458,N_33241,N_33982);
and U34459 (N_34459,N_33367,N_33858);
xnor U34460 (N_34460,N_33654,N_33154);
xor U34461 (N_34461,N_33983,N_33173);
xnor U34462 (N_34462,N_33861,N_33341);
and U34463 (N_34463,N_33526,N_33276);
nor U34464 (N_34464,N_33451,N_33876);
nor U34465 (N_34465,N_33927,N_33507);
and U34466 (N_34466,N_33843,N_33336);
and U34467 (N_34467,N_33803,N_33077);
and U34468 (N_34468,N_33945,N_33328);
xnor U34469 (N_34469,N_33107,N_33607);
or U34470 (N_34470,N_33555,N_33189);
nor U34471 (N_34471,N_33921,N_33045);
nand U34472 (N_34472,N_33549,N_33383);
and U34473 (N_34473,N_33841,N_33976);
nor U34474 (N_34474,N_33007,N_33684);
xnor U34475 (N_34475,N_33244,N_33679);
or U34476 (N_34476,N_33864,N_33015);
nand U34477 (N_34477,N_33488,N_33659);
or U34478 (N_34478,N_33634,N_33812);
and U34479 (N_34479,N_33545,N_33448);
and U34480 (N_34480,N_33005,N_33433);
xor U34481 (N_34481,N_33186,N_33928);
or U34482 (N_34482,N_33060,N_33343);
nor U34483 (N_34483,N_33277,N_33663);
xnor U34484 (N_34484,N_33568,N_33819);
nor U34485 (N_34485,N_33430,N_33759);
or U34486 (N_34486,N_33648,N_33071);
nand U34487 (N_34487,N_33636,N_33768);
and U34488 (N_34488,N_33954,N_33609);
nand U34489 (N_34489,N_33223,N_33268);
xor U34490 (N_34490,N_33784,N_33848);
xnor U34491 (N_34491,N_33517,N_33053);
or U34492 (N_34492,N_33860,N_33750);
nor U34493 (N_34493,N_33524,N_33466);
nand U34494 (N_34494,N_33499,N_33047);
or U34495 (N_34495,N_33767,N_33828);
and U34496 (N_34496,N_33885,N_33176);
nand U34497 (N_34497,N_33029,N_33697);
and U34498 (N_34498,N_33839,N_33523);
nand U34499 (N_34499,N_33754,N_33070);
or U34500 (N_34500,N_33852,N_33850);
xor U34501 (N_34501,N_33321,N_33460);
nor U34502 (N_34502,N_33126,N_33731);
or U34503 (N_34503,N_33113,N_33998);
or U34504 (N_34504,N_33177,N_33013);
and U34505 (N_34505,N_33370,N_33774);
nor U34506 (N_34506,N_33287,N_33360);
or U34507 (N_34507,N_33814,N_33317);
nor U34508 (N_34508,N_33955,N_33386);
and U34509 (N_34509,N_33882,N_33103);
nand U34510 (N_34510,N_33961,N_33478);
and U34511 (N_34511,N_33018,N_33801);
and U34512 (N_34512,N_33679,N_33830);
nor U34513 (N_34513,N_33100,N_33733);
xor U34514 (N_34514,N_33208,N_33560);
or U34515 (N_34515,N_33298,N_33414);
nor U34516 (N_34516,N_33818,N_33751);
or U34517 (N_34517,N_33328,N_33918);
nand U34518 (N_34518,N_33921,N_33997);
and U34519 (N_34519,N_33519,N_33826);
nor U34520 (N_34520,N_33846,N_33725);
nor U34521 (N_34521,N_33363,N_33472);
xnor U34522 (N_34522,N_33731,N_33177);
or U34523 (N_34523,N_33868,N_33489);
or U34524 (N_34524,N_33667,N_33769);
nand U34525 (N_34525,N_33151,N_33182);
or U34526 (N_34526,N_33697,N_33835);
nand U34527 (N_34527,N_33203,N_33643);
nor U34528 (N_34528,N_33001,N_33014);
nand U34529 (N_34529,N_33927,N_33695);
xor U34530 (N_34530,N_33210,N_33274);
xor U34531 (N_34531,N_33500,N_33050);
or U34532 (N_34532,N_33217,N_33596);
or U34533 (N_34533,N_33728,N_33499);
and U34534 (N_34534,N_33691,N_33737);
nor U34535 (N_34535,N_33334,N_33407);
xnor U34536 (N_34536,N_33339,N_33856);
nand U34537 (N_34537,N_33154,N_33829);
nor U34538 (N_34538,N_33621,N_33964);
and U34539 (N_34539,N_33947,N_33685);
nand U34540 (N_34540,N_33968,N_33325);
and U34541 (N_34541,N_33442,N_33106);
xnor U34542 (N_34542,N_33882,N_33267);
nand U34543 (N_34543,N_33352,N_33040);
or U34544 (N_34544,N_33017,N_33609);
nor U34545 (N_34545,N_33305,N_33877);
or U34546 (N_34546,N_33110,N_33459);
xnor U34547 (N_34547,N_33259,N_33848);
xnor U34548 (N_34548,N_33314,N_33523);
xnor U34549 (N_34549,N_33056,N_33776);
xor U34550 (N_34550,N_33592,N_33435);
nand U34551 (N_34551,N_33465,N_33823);
nor U34552 (N_34552,N_33377,N_33370);
or U34553 (N_34553,N_33421,N_33256);
nand U34554 (N_34554,N_33593,N_33936);
xnor U34555 (N_34555,N_33829,N_33924);
xor U34556 (N_34556,N_33276,N_33590);
nor U34557 (N_34557,N_33114,N_33814);
nand U34558 (N_34558,N_33797,N_33396);
and U34559 (N_34559,N_33801,N_33799);
or U34560 (N_34560,N_33138,N_33338);
and U34561 (N_34561,N_33210,N_33758);
nor U34562 (N_34562,N_33826,N_33389);
nor U34563 (N_34563,N_33542,N_33015);
nand U34564 (N_34564,N_33149,N_33645);
and U34565 (N_34565,N_33561,N_33679);
nand U34566 (N_34566,N_33760,N_33716);
and U34567 (N_34567,N_33910,N_33004);
nor U34568 (N_34568,N_33241,N_33601);
or U34569 (N_34569,N_33270,N_33525);
or U34570 (N_34570,N_33951,N_33190);
nor U34571 (N_34571,N_33655,N_33215);
nand U34572 (N_34572,N_33497,N_33336);
nand U34573 (N_34573,N_33968,N_33887);
xor U34574 (N_34574,N_33818,N_33361);
nand U34575 (N_34575,N_33826,N_33570);
nand U34576 (N_34576,N_33256,N_33348);
or U34577 (N_34577,N_33555,N_33101);
xnor U34578 (N_34578,N_33355,N_33561);
nor U34579 (N_34579,N_33884,N_33118);
or U34580 (N_34580,N_33626,N_33249);
and U34581 (N_34581,N_33727,N_33129);
xor U34582 (N_34582,N_33354,N_33631);
xnor U34583 (N_34583,N_33814,N_33462);
or U34584 (N_34584,N_33321,N_33165);
xnor U34585 (N_34585,N_33429,N_33697);
nand U34586 (N_34586,N_33846,N_33056);
nand U34587 (N_34587,N_33497,N_33116);
xor U34588 (N_34588,N_33229,N_33603);
nand U34589 (N_34589,N_33397,N_33031);
and U34590 (N_34590,N_33049,N_33445);
xnor U34591 (N_34591,N_33102,N_33345);
and U34592 (N_34592,N_33411,N_33056);
nand U34593 (N_34593,N_33487,N_33653);
nor U34594 (N_34594,N_33592,N_33870);
or U34595 (N_34595,N_33480,N_33904);
or U34596 (N_34596,N_33483,N_33936);
nand U34597 (N_34597,N_33753,N_33242);
nand U34598 (N_34598,N_33130,N_33085);
and U34599 (N_34599,N_33034,N_33796);
and U34600 (N_34600,N_33574,N_33779);
or U34601 (N_34601,N_33026,N_33513);
nor U34602 (N_34602,N_33262,N_33113);
nor U34603 (N_34603,N_33775,N_33345);
nand U34604 (N_34604,N_33652,N_33202);
or U34605 (N_34605,N_33137,N_33324);
or U34606 (N_34606,N_33965,N_33334);
or U34607 (N_34607,N_33646,N_33974);
or U34608 (N_34608,N_33211,N_33642);
xor U34609 (N_34609,N_33243,N_33320);
or U34610 (N_34610,N_33601,N_33518);
nand U34611 (N_34611,N_33242,N_33404);
xor U34612 (N_34612,N_33311,N_33473);
or U34613 (N_34613,N_33639,N_33602);
nor U34614 (N_34614,N_33192,N_33058);
nand U34615 (N_34615,N_33877,N_33799);
or U34616 (N_34616,N_33349,N_33136);
xor U34617 (N_34617,N_33446,N_33703);
xor U34618 (N_34618,N_33451,N_33122);
nor U34619 (N_34619,N_33815,N_33785);
xnor U34620 (N_34620,N_33801,N_33260);
nand U34621 (N_34621,N_33958,N_33669);
xor U34622 (N_34622,N_33561,N_33563);
and U34623 (N_34623,N_33921,N_33767);
and U34624 (N_34624,N_33867,N_33225);
nor U34625 (N_34625,N_33336,N_33829);
and U34626 (N_34626,N_33345,N_33105);
nand U34627 (N_34627,N_33114,N_33820);
and U34628 (N_34628,N_33250,N_33009);
or U34629 (N_34629,N_33744,N_33565);
and U34630 (N_34630,N_33466,N_33021);
nor U34631 (N_34631,N_33301,N_33651);
or U34632 (N_34632,N_33130,N_33263);
xor U34633 (N_34633,N_33214,N_33131);
or U34634 (N_34634,N_33947,N_33667);
nor U34635 (N_34635,N_33249,N_33698);
or U34636 (N_34636,N_33354,N_33470);
xor U34637 (N_34637,N_33355,N_33522);
nor U34638 (N_34638,N_33670,N_33715);
nor U34639 (N_34639,N_33658,N_33410);
nor U34640 (N_34640,N_33322,N_33775);
and U34641 (N_34641,N_33368,N_33575);
or U34642 (N_34642,N_33793,N_33492);
nor U34643 (N_34643,N_33433,N_33077);
or U34644 (N_34644,N_33245,N_33207);
or U34645 (N_34645,N_33759,N_33864);
and U34646 (N_34646,N_33877,N_33611);
nor U34647 (N_34647,N_33274,N_33580);
nand U34648 (N_34648,N_33201,N_33206);
nand U34649 (N_34649,N_33703,N_33471);
and U34650 (N_34650,N_33034,N_33486);
or U34651 (N_34651,N_33134,N_33386);
xor U34652 (N_34652,N_33684,N_33168);
and U34653 (N_34653,N_33642,N_33398);
nand U34654 (N_34654,N_33656,N_33921);
xor U34655 (N_34655,N_33639,N_33882);
and U34656 (N_34656,N_33480,N_33522);
or U34657 (N_34657,N_33356,N_33898);
nand U34658 (N_34658,N_33485,N_33069);
or U34659 (N_34659,N_33335,N_33278);
xnor U34660 (N_34660,N_33125,N_33582);
or U34661 (N_34661,N_33494,N_33822);
and U34662 (N_34662,N_33438,N_33985);
or U34663 (N_34663,N_33842,N_33070);
xnor U34664 (N_34664,N_33750,N_33988);
nor U34665 (N_34665,N_33433,N_33401);
xnor U34666 (N_34666,N_33711,N_33584);
nor U34667 (N_34667,N_33010,N_33323);
or U34668 (N_34668,N_33701,N_33165);
nor U34669 (N_34669,N_33701,N_33011);
nor U34670 (N_34670,N_33955,N_33098);
or U34671 (N_34671,N_33745,N_33546);
and U34672 (N_34672,N_33849,N_33598);
or U34673 (N_34673,N_33636,N_33273);
nand U34674 (N_34674,N_33221,N_33195);
xor U34675 (N_34675,N_33421,N_33763);
and U34676 (N_34676,N_33337,N_33274);
or U34677 (N_34677,N_33720,N_33098);
or U34678 (N_34678,N_33226,N_33583);
or U34679 (N_34679,N_33541,N_33926);
or U34680 (N_34680,N_33180,N_33380);
and U34681 (N_34681,N_33078,N_33730);
nor U34682 (N_34682,N_33250,N_33695);
nand U34683 (N_34683,N_33947,N_33520);
nor U34684 (N_34684,N_33527,N_33769);
nor U34685 (N_34685,N_33053,N_33409);
xnor U34686 (N_34686,N_33183,N_33273);
or U34687 (N_34687,N_33329,N_33309);
nand U34688 (N_34688,N_33173,N_33476);
xor U34689 (N_34689,N_33620,N_33764);
nand U34690 (N_34690,N_33316,N_33540);
or U34691 (N_34691,N_33117,N_33796);
xnor U34692 (N_34692,N_33178,N_33576);
nand U34693 (N_34693,N_33442,N_33178);
nor U34694 (N_34694,N_33893,N_33617);
nand U34695 (N_34695,N_33682,N_33489);
or U34696 (N_34696,N_33363,N_33428);
nand U34697 (N_34697,N_33122,N_33025);
and U34698 (N_34698,N_33653,N_33390);
nand U34699 (N_34699,N_33155,N_33702);
xor U34700 (N_34700,N_33920,N_33174);
or U34701 (N_34701,N_33104,N_33699);
nand U34702 (N_34702,N_33043,N_33059);
nand U34703 (N_34703,N_33595,N_33111);
or U34704 (N_34704,N_33439,N_33957);
or U34705 (N_34705,N_33532,N_33945);
nand U34706 (N_34706,N_33791,N_33077);
xor U34707 (N_34707,N_33133,N_33242);
nor U34708 (N_34708,N_33430,N_33334);
and U34709 (N_34709,N_33566,N_33525);
nand U34710 (N_34710,N_33231,N_33451);
xnor U34711 (N_34711,N_33277,N_33012);
nor U34712 (N_34712,N_33729,N_33282);
xnor U34713 (N_34713,N_33065,N_33885);
nand U34714 (N_34714,N_33869,N_33820);
or U34715 (N_34715,N_33809,N_33568);
xnor U34716 (N_34716,N_33094,N_33957);
and U34717 (N_34717,N_33346,N_33178);
xnor U34718 (N_34718,N_33927,N_33156);
or U34719 (N_34719,N_33148,N_33615);
nor U34720 (N_34720,N_33810,N_33040);
nand U34721 (N_34721,N_33507,N_33986);
nor U34722 (N_34722,N_33018,N_33379);
xnor U34723 (N_34723,N_33329,N_33694);
nand U34724 (N_34724,N_33089,N_33063);
and U34725 (N_34725,N_33648,N_33783);
nand U34726 (N_34726,N_33350,N_33800);
nor U34727 (N_34727,N_33722,N_33109);
and U34728 (N_34728,N_33759,N_33051);
and U34729 (N_34729,N_33309,N_33723);
nor U34730 (N_34730,N_33952,N_33201);
or U34731 (N_34731,N_33057,N_33373);
nand U34732 (N_34732,N_33971,N_33986);
or U34733 (N_34733,N_33336,N_33126);
or U34734 (N_34734,N_33066,N_33460);
xor U34735 (N_34735,N_33655,N_33125);
xnor U34736 (N_34736,N_33346,N_33118);
and U34737 (N_34737,N_33844,N_33057);
nand U34738 (N_34738,N_33586,N_33785);
nand U34739 (N_34739,N_33854,N_33232);
nand U34740 (N_34740,N_33609,N_33178);
xnor U34741 (N_34741,N_33635,N_33973);
or U34742 (N_34742,N_33441,N_33823);
and U34743 (N_34743,N_33557,N_33015);
nor U34744 (N_34744,N_33800,N_33909);
nand U34745 (N_34745,N_33012,N_33057);
nor U34746 (N_34746,N_33987,N_33184);
nand U34747 (N_34747,N_33955,N_33867);
nor U34748 (N_34748,N_33905,N_33435);
or U34749 (N_34749,N_33544,N_33951);
nand U34750 (N_34750,N_33621,N_33297);
xnor U34751 (N_34751,N_33177,N_33043);
xnor U34752 (N_34752,N_33251,N_33417);
and U34753 (N_34753,N_33507,N_33052);
nor U34754 (N_34754,N_33345,N_33939);
or U34755 (N_34755,N_33568,N_33695);
nand U34756 (N_34756,N_33442,N_33846);
nand U34757 (N_34757,N_33157,N_33251);
xor U34758 (N_34758,N_33739,N_33047);
nor U34759 (N_34759,N_33072,N_33430);
xnor U34760 (N_34760,N_33786,N_33428);
and U34761 (N_34761,N_33710,N_33418);
xor U34762 (N_34762,N_33813,N_33927);
or U34763 (N_34763,N_33423,N_33562);
nor U34764 (N_34764,N_33325,N_33363);
or U34765 (N_34765,N_33436,N_33276);
nor U34766 (N_34766,N_33151,N_33354);
xnor U34767 (N_34767,N_33256,N_33366);
and U34768 (N_34768,N_33447,N_33677);
and U34769 (N_34769,N_33982,N_33703);
and U34770 (N_34770,N_33126,N_33365);
xnor U34771 (N_34771,N_33864,N_33081);
nand U34772 (N_34772,N_33840,N_33336);
xnor U34773 (N_34773,N_33273,N_33108);
nand U34774 (N_34774,N_33876,N_33250);
nor U34775 (N_34775,N_33388,N_33445);
and U34776 (N_34776,N_33028,N_33782);
nor U34777 (N_34777,N_33034,N_33971);
nand U34778 (N_34778,N_33147,N_33310);
or U34779 (N_34779,N_33332,N_33020);
nand U34780 (N_34780,N_33215,N_33218);
and U34781 (N_34781,N_33003,N_33008);
or U34782 (N_34782,N_33929,N_33462);
nor U34783 (N_34783,N_33988,N_33113);
or U34784 (N_34784,N_33340,N_33773);
or U34785 (N_34785,N_33056,N_33789);
and U34786 (N_34786,N_33899,N_33076);
nand U34787 (N_34787,N_33874,N_33634);
nand U34788 (N_34788,N_33515,N_33759);
xnor U34789 (N_34789,N_33577,N_33243);
and U34790 (N_34790,N_33526,N_33917);
and U34791 (N_34791,N_33988,N_33465);
or U34792 (N_34792,N_33217,N_33377);
xnor U34793 (N_34793,N_33165,N_33125);
nor U34794 (N_34794,N_33949,N_33702);
and U34795 (N_34795,N_33355,N_33265);
and U34796 (N_34796,N_33238,N_33801);
or U34797 (N_34797,N_33797,N_33831);
or U34798 (N_34798,N_33742,N_33663);
nor U34799 (N_34799,N_33697,N_33937);
and U34800 (N_34800,N_33127,N_33860);
and U34801 (N_34801,N_33623,N_33902);
nand U34802 (N_34802,N_33855,N_33563);
nor U34803 (N_34803,N_33732,N_33528);
xor U34804 (N_34804,N_33059,N_33140);
and U34805 (N_34805,N_33969,N_33409);
and U34806 (N_34806,N_33692,N_33706);
nor U34807 (N_34807,N_33882,N_33214);
xnor U34808 (N_34808,N_33687,N_33132);
nand U34809 (N_34809,N_33323,N_33194);
and U34810 (N_34810,N_33098,N_33556);
xnor U34811 (N_34811,N_33336,N_33014);
and U34812 (N_34812,N_33058,N_33447);
nor U34813 (N_34813,N_33326,N_33130);
xor U34814 (N_34814,N_33776,N_33503);
nor U34815 (N_34815,N_33431,N_33882);
and U34816 (N_34816,N_33595,N_33490);
and U34817 (N_34817,N_33306,N_33941);
nand U34818 (N_34818,N_33244,N_33448);
or U34819 (N_34819,N_33581,N_33220);
nand U34820 (N_34820,N_33005,N_33642);
or U34821 (N_34821,N_33995,N_33509);
xnor U34822 (N_34822,N_33589,N_33345);
and U34823 (N_34823,N_33294,N_33753);
or U34824 (N_34824,N_33331,N_33460);
and U34825 (N_34825,N_33192,N_33027);
nor U34826 (N_34826,N_33271,N_33426);
nor U34827 (N_34827,N_33597,N_33247);
nand U34828 (N_34828,N_33157,N_33922);
or U34829 (N_34829,N_33351,N_33913);
and U34830 (N_34830,N_33774,N_33713);
and U34831 (N_34831,N_33880,N_33508);
nand U34832 (N_34832,N_33433,N_33400);
nand U34833 (N_34833,N_33549,N_33318);
nor U34834 (N_34834,N_33139,N_33788);
xor U34835 (N_34835,N_33174,N_33157);
or U34836 (N_34836,N_33422,N_33178);
nand U34837 (N_34837,N_33919,N_33358);
nand U34838 (N_34838,N_33309,N_33243);
and U34839 (N_34839,N_33903,N_33510);
nor U34840 (N_34840,N_33233,N_33266);
and U34841 (N_34841,N_33450,N_33679);
xnor U34842 (N_34842,N_33189,N_33146);
nand U34843 (N_34843,N_33304,N_33437);
and U34844 (N_34844,N_33121,N_33781);
and U34845 (N_34845,N_33912,N_33300);
nor U34846 (N_34846,N_33398,N_33432);
or U34847 (N_34847,N_33182,N_33737);
nor U34848 (N_34848,N_33201,N_33183);
nor U34849 (N_34849,N_33722,N_33929);
or U34850 (N_34850,N_33379,N_33120);
xnor U34851 (N_34851,N_33076,N_33260);
and U34852 (N_34852,N_33082,N_33994);
and U34853 (N_34853,N_33618,N_33310);
xor U34854 (N_34854,N_33777,N_33336);
nor U34855 (N_34855,N_33128,N_33934);
nand U34856 (N_34856,N_33419,N_33130);
xor U34857 (N_34857,N_33144,N_33128);
xor U34858 (N_34858,N_33493,N_33118);
and U34859 (N_34859,N_33886,N_33686);
or U34860 (N_34860,N_33620,N_33205);
nand U34861 (N_34861,N_33708,N_33359);
nand U34862 (N_34862,N_33664,N_33446);
nor U34863 (N_34863,N_33223,N_33521);
and U34864 (N_34864,N_33975,N_33474);
nand U34865 (N_34865,N_33492,N_33972);
nand U34866 (N_34866,N_33852,N_33392);
or U34867 (N_34867,N_33865,N_33923);
nor U34868 (N_34868,N_33072,N_33808);
xnor U34869 (N_34869,N_33923,N_33757);
xor U34870 (N_34870,N_33822,N_33427);
and U34871 (N_34871,N_33089,N_33541);
or U34872 (N_34872,N_33253,N_33468);
nand U34873 (N_34873,N_33394,N_33027);
or U34874 (N_34874,N_33312,N_33780);
and U34875 (N_34875,N_33918,N_33122);
xnor U34876 (N_34876,N_33018,N_33126);
and U34877 (N_34877,N_33485,N_33481);
or U34878 (N_34878,N_33034,N_33969);
or U34879 (N_34879,N_33627,N_33424);
nor U34880 (N_34880,N_33063,N_33276);
or U34881 (N_34881,N_33606,N_33207);
or U34882 (N_34882,N_33296,N_33043);
nand U34883 (N_34883,N_33988,N_33857);
xnor U34884 (N_34884,N_33418,N_33812);
xnor U34885 (N_34885,N_33661,N_33535);
xnor U34886 (N_34886,N_33165,N_33632);
xor U34887 (N_34887,N_33813,N_33977);
and U34888 (N_34888,N_33084,N_33543);
nand U34889 (N_34889,N_33214,N_33549);
nand U34890 (N_34890,N_33936,N_33187);
or U34891 (N_34891,N_33501,N_33859);
and U34892 (N_34892,N_33428,N_33344);
and U34893 (N_34893,N_33322,N_33487);
or U34894 (N_34894,N_33452,N_33951);
nand U34895 (N_34895,N_33227,N_33360);
or U34896 (N_34896,N_33109,N_33897);
or U34897 (N_34897,N_33431,N_33451);
or U34898 (N_34898,N_33303,N_33211);
nor U34899 (N_34899,N_33363,N_33139);
nor U34900 (N_34900,N_33399,N_33144);
nand U34901 (N_34901,N_33339,N_33705);
or U34902 (N_34902,N_33754,N_33654);
nand U34903 (N_34903,N_33572,N_33126);
nor U34904 (N_34904,N_33860,N_33831);
or U34905 (N_34905,N_33902,N_33413);
nor U34906 (N_34906,N_33633,N_33626);
and U34907 (N_34907,N_33400,N_33010);
nand U34908 (N_34908,N_33514,N_33170);
nand U34909 (N_34909,N_33987,N_33146);
or U34910 (N_34910,N_33680,N_33526);
or U34911 (N_34911,N_33785,N_33187);
xnor U34912 (N_34912,N_33627,N_33282);
xnor U34913 (N_34913,N_33339,N_33408);
or U34914 (N_34914,N_33732,N_33677);
nor U34915 (N_34915,N_33449,N_33285);
or U34916 (N_34916,N_33072,N_33710);
xnor U34917 (N_34917,N_33920,N_33221);
and U34918 (N_34918,N_33575,N_33660);
nand U34919 (N_34919,N_33854,N_33010);
nand U34920 (N_34920,N_33841,N_33517);
or U34921 (N_34921,N_33923,N_33502);
nand U34922 (N_34922,N_33510,N_33541);
and U34923 (N_34923,N_33196,N_33543);
xor U34924 (N_34924,N_33597,N_33702);
and U34925 (N_34925,N_33663,N_33789);
nand U34926 (N_34926,N_33867,N_33473);
or U34927 (N_34927,N_33536,N_33027);
nor U34928 (N_34928,N_33254,N_33411);
nor U34929 (N_34929,N_33772,N_33680);
nand U34930 (N_34930,N_33295,N_33307);
and U34931 (N_34931,N_33262,N_33872);
xor U34932 (N_34932,N_33327,N_33643);
and U34933 (N_34933,N_33017,N_33569);
nor U34934 (N_34934,N_33341,N_33260);
and U34935 (N_34935,N_33119,N_33266);
nor U34936 (N_34936,N_33069,N_33496);
and U34937 (N_34937,N_33837,N_33287);
xor U34938 (N_34938,N_33795,N_33710);
xor U34939 (N_34939,N_33248,N_33360);
nand U34940 (N_34940,N_33643,N_33379);
or U34941 (N_34941,N_33765,N_33402);
nor U34942 (N_34942,N_33578,N_33590);
or U34943 (N_34943,N_33597,N_33879);
xnor U34944 (N_34944,N_33435,N_33617);
or U34945 (N_34945,N_33080,N_33324);
or U34946 (N_34946,N_33022,N_33062);
or U34947 (N_34947,N_33162,N_33969);
nor U34948 (N_34948,N_33159,N_33459);
nand U34949 (N_34949,N_33469,N_33090);
xnor U34950 (N_34950,N_33190,N_33559);
nand U34951 (N_34951,N_33242,N_33415);
xor U34952 (N_34952,N_33328,N_33891);
nand U34953 (N_34953,N_33470,N_33980);
xnor U34954 (N_34954,N_33366,N_33615);
or U34955 (N_34955,N_33091,N_33348);
nand U34956 (N_34956,N_33382,N_33132);
or U34957 (N_34957,N_33484,N_33192);
or U34958 (N_34958,N_33228,N_33795);
or U34959 (N_34959,N_33200,N_33607);
xnor U34960 (N_34960,N_33548,N_33684);
nand U34961 (N_34961,N_33567,N_33382);
nor U34962 (N_34962,N_33764,N_33422);
xnor U34963 (N_34963,N_33474,N_33998);
or U34964 (N_34964,N_33240,N_33810);
nand U34965 (N_34965,N_33062,N_33256);
xor U34966 (N_34966,N_33645,N_33209);
nand U34967 (N_34967,N_33282,N_33437);
and U34968 (N_34968,N_33571,N_33949);
xor U34969 (N_34969,N_33232,N_33455);
or U34970 (N_34970,N_33051,N_33512);
or U34971 (N_34971,N_33230,N_33076);
nand U34972 (N_34972,N_33770,N_33626);
nand U34973 (N_34973,N_33931,N_33105);
or U34974 (N_34974,N_33009,N_33631);
nor U34975 (N_34975,N_33255,N_33936);
xor U34976 (N_34976,N_33887,N_33382);
xnor U34977 (N_34977,N_33168,N_33943);
and U34978 (N_34978,N_33779,N_33611);
nor U34979 (N_34979,N_33219,N_33364);
nand U34980 (N_34980,N_33572,N_33267);
or U34981 (N_34981,N_33059,N_33443);
nor U34982 (N_34982,N_33516,N_33220);
nand U34983 (N_34983,N_33264,N_33781);
or U34984 (N_34984,N_33421,N_33847);
nand U34985 (N_34985,N_33906,N_33087);
nand U34986 (N_34986,N_33010,N_33574);
nand U34987 (N_34987,N_33829,N_33750);
nand U34988 (N_34988,N_33714,N_33045);
nand U34989 (N_34989,N_33310,N_33611);
nor U34990 (N_34990,N_33795,N_33315);
or U34991 (N_34991,N_33670,N_33036);
nand U34992 (N_34992,N_33274,N_33040);
xnor U34993 (N_34993,N_33149,N_33543);
or U34994 (N_34994,N_33443,N_33826);
or U34995 (N_34995,N_33362,N_33344);
and U34996 (N_34996,N_33569,N_33933);
or U34997 (N_34997,N_33234,N_33800);
nand U34998 (N_34998,N_33001,N_33238);
nor U34999 (N_34999,N_33681,N_33972);
and U35000 (N_35000,N_34080,N_34193);
xor U35001 (N_35001,N_34467,N_34470);
xor U35002 (N_35002,N_34680,N_34938);
nor U35003 (N_35003,N_34349,N_34290);
xor U35004 (N_35004,N_34119,N_34528);
nand U35005 (N_35005,N_34357,N_34446);
or U35006 (N_35006,N_34718,N_34825);
nor U35007 (N_35007,N_34994,N_34968);
or U35008 (N_35008,N_34147,N_34191);
nor U35009 (N_35009,N_34271,N_34774);
nand U35010 (N_35010,N_34843,N_34242);
nor U35011 (N_35011,N_34034,N_34978);
and U35012 (N_35012,N_34902,N_34494);
nand U35013 (N_35013,N_34218,N_34906);
nor U35014 (N_35014,N_34819,N_34138);
or U35015 (N_35015,N_34237,N_34118);
xnor U35016 (N_35016,N_34610,N_34281);
xor U35017 (N_35017,N_34251,N_34519);
and U35018 (N_35018,N_34256,N_34399);
or U35019 (N_35019,N_34568,N_34581);
or U35020 (N_35020,N_34828,N_34764);
nor U35021 (N_35021,N_34004,N_34327);
xnor U35022 (N_35022,N_34505,N_34612);
nand U35023 (N_35023,N_34223,N_34373);
nand U35024 (N_35024,N_34288,N_34876);
nor U35025 (N_35025,N_34168,N_34779);
xnor U35026 (N_35026,N_34244,N_34411);
nor U35027 (N_35027,N_34189,N_34057);
nand U35028 (N_35028,N_34955,N_34041);
xnor U35029 (N_35029,N_34386,N_34018);
or U35030 (N_35030,N_34420,N_34816);
or U35031 (N_35031,N_34635,N_34884);
nand U35032 (N_35032,N_34712,N_34609);
nor U35033 (N_35033,N_34587,N_34196);
or U35034 (N_35034,N_34973,N_34391);
and U35035 (N_35035,N_34023,N_34835);
and U35036 (N_35036,N_34694,N_34173);
xor U35037 (N_35037,N_34254,N_34472);
nor U35038 (N_35038,N_34940,N_34659);
nand U35039 (N_35039,N_34860,N_34416);
nor U35040 (N_35040,N_34336,N_34997);
or U35041 (N_35041,N_34544,N_34069);
xnor U35042 (N_35042,N_34238,N_34727);
nand U35043 (N_35043,N_34706,N_34880);
xor U35044 (N_35044,N_34353,N_34099);
and U35045 (N_35045,N_34976,N_34947);
xor U35046 (N_35046,N_34967,N_34804);
or U35047 (N_35047,N_34114,N_34499);
or U35048 (N_35048,N_34371,N_34086);
nand U35049 (N_35049,N_34886,N_34527);
or U35050 (N_35050,N_34410,N_34897);
or U35051 (N_35051,N_34056,N_34195);
and U35052 (N_35052,N_34564,N_34423);
nor U35053 (N_35053,N_34582,N_34093);
or U35054 (N_35054,N_34769,N_34401);
xor U35055 (N_35055,N_34275,N_34862);
xor U35056 (N_35056,N_34987,N_34949);
nand U35057 (N_35057,N_34370,N_34224);
and U35058 (N_35058,N_34617,N_34533);
nor U35059 (N_35059,N_34531,N_34982);
and U35060 (N_35060,N_34882,N_34365);
nand U35061 (N_35061,N_34062,N_34044);
nor U35062 (N_35062,N_34012,N_34405);
nor U35063 (N_35063,N_34398,N_34160);
nor U35064 (N_35064,N_34309,N_34717);
or U35065 (N_35065,N_34767,N_34132);
nand U35066 (N_35066,N_34222,N_34143);
xor U35067 (N_35067,N_34338,N_34212);
nand U35068 (N_35068,N_34040,N_34337);
xor U35069 (N_35069,N_34217,N_34347);
xor U35070 (N_35070,N_34765,N_34841);
and U35071 (N_35071,N_34301,N_34546);
or U35072 (N_35072,N_34704,N_34346);
nand U35073 (N_35073,N_34203,N_34507);
and U35074 (N_35074,N_34390,N_34760);
nor U35075 (N_35075,N_34959,N_34632);
xnor U35076 (N_35076,N_34537,N_34891);
nor U35077 (N_35077,N_34125,N_34622);
xor U35078 (N_35078,N_34752,N_34576);
xor U35079 (N_35079,N_34487,N_34356);
nand U35080 (N_35080,N_34434,N_34259);
and U35081 (N_35081,N_34011,N_34594);
or U35082 (N_35082,N_34351,N_34406);
nand U35083 (N_35083,N_34215,N_34321);
xor U35084 (N_35084,N_34059,N_34255);
nor U35085 (N_35085,N_34780,N_34175);
and U35086 (N_35086,N_34444,N_34504);
or U35087 (N_35087,N_34422,N_34042);
and U35088 (N_35088,N_34186,N_34800);
or U35089 (N_35089,N_34087,N_34778);
nand U35090 (N_35090,N_34863,N_34798);
nor U35091 (N_35091,N_34162,N_34851);
xnor U35092 (N_35092,N_34912,N_34895);
or U35093 (N_35093,N_34362,N_34817);
or U35094 (N_35094,N_34993,N_34014);
xor U35095 (N_35095,N_34810,N_34557);
nor U35096 (N_35096,N_34899,N_34685);
or U35097 (N_35097,N_34302,N_34512);
nand U35098 (N_35098,N_34695,N_34079);
xnor U35099 (N_35099,N_34241,N_34358);
or U35100 (N_35100,N_34787,N_34623);
and U35101 (N_35101,N_34793,N_34104);
or U35102 (N_35102,N_34805,N_34318);
nand U35103 (N_35103,N_34269,N_34802);
nand U35104 (N_35104,N_34739,N_34178);
xor U35105 (N_35105,N_34992,N_34952);
nor U35106 (N_35106,N_34131,N_34742);
or U35107 (N_35107,N_34424,N_34204);
xnor U35108 (N_35108,N_34556,N_34293);
xor U35109 (N_35109,N_34231,N_34720);
or U35110 (N_35110,N_34169,N_34698);
and U35111 (N_35111,N_34310,N_34170);
nand U35112 (N_35112,N_34957,N_34484);
or U35113 (N_35113,N_34772,N_34615);
and U35114 (N_35114,N_34672,N_34550);
and U35115 (N_35115,N_34258,N_34154);
nor U35116 (N_35116,N_34171,N_34194);
xnor U35117 (N_35117,N_34654,N_34799);
xor U35118 (N_35118,N_34901,N_34257);
and U35119 (N_35119,N_34482,N_34331);
nand U35120 (N_35120,N_34052,N_34364);
xor U35121 (N_35121,N_34153,N_34511);
and U35122 (N_35122,N_34287,N_34917);
nand U35123 (N_35123,N_34642,N_34524);
xor U35124 (N_35124,N_34105,N_34822);
nor U35125 (N_35125,N_34939,N_34759);
nor U35126 (N_35126,N_34137,N_34664);
and U35127 (N_35127,N_34913,N_34836);
and U35128 (N_35128,N_34380,N_34021);
nand U35129 (N_35129,N_34988,N_34709);
xor U35130 (N_35130,N_34055,N_34181);
xnor U35131 (N_35131,N_34868,N_34784);
nand U35132 (N_35132,N_34015,N_34956);
and U35133 (N_35133,N_34999,N_34001);
nor U35134 (N_35134,N_34812,N_34350);
or U35135 (N_35135,N_34588,N_34716);
nand U35136 (N_35136,N_34239,N_34077);
nor U35137 (N_35137,N_34773,N_34148);
nand U35138 (N_35138,N_34552,N_34155);
nand U35139 (N_35139,N_34864,N_34777);
nand U35140 (N_35140,N_34848,N_34363);
nand U35141 (N_35141,N_34651,N_34120);
nor U35142 (N_35142,N_34000,N_34756);
nor U35143 (N_35143,N_34655,N_34705);
xor U35144 (N_35144,N_34246,N_34885);
or U35145 (N_35145,N_34574,N_34442);
xor U35146 (N_35146,N_34758,N_34316);
or U35147 (N_35147,N_34156,N_34396);
and U35148 (N_35148,N_34413,N_34943);
nor U35149 (N_35149,N_34532,N_34397);
xnor U35150 (N_35150,N_34247,N_34019);
xnor U35151 (N_35151,N_34865,N_34045);
and U35152 (N_35152,N_34834,N_34233);
nor U35153 (N_35153,N_34123,N_34436);
nand U35154 (N_35154,N_34935,N_34094);
nand U35155 (N_35155,N_34749,N_34944);
nand U35156 (N_35156,N_34279,N_34688);
nand U35157 (N_35157,N_34025,N_34916);
nand U35158 (N_35158,N_34963,N_34490);
nor U35159 (N_35159,N_34295,N_34228);
xnor U35160 (N_35160,N_34109,N_34983);
and U35161 (N_35161,N_34996,N_34616);
xnor U35162 (N_35162,N_34549,N_34107);
nor U35163 (N_35163,N_34219,N_34657);
xnor U35164 (N_35164,N_34638,N_34686);
xnor U35165 (N_35165,N_34419,N_34908);
nand U35166 (N_35166,N_34711,N_34343);
or U35167 (N_35167,N_34690,N_34072);
or U35168 (N_35168,N_34268,N_34625);
xnor U35169 (N_35169,N_34469,N_34850);
xnor U35170 (N_35170,N_34185,N_34853);
and U35171 (N_35171,N_34184,N_34207);
nand U35172 (N_35172,N_34547,N_34427);
or U35173 (N_35173,N_34438,N_34746);
xnor U35174 (N_35174,N_34248,N_34394);
xnor U35175 (N_35175,N_34368,N_34971);
nand U35176 (N_35176,N_34307,N_34621);
and U35177 (N_35177,N_34283,N_34262);
xnor U35178 (N_35178,N_34923,N_34395);
xnor U35179 (N_35179,N_34890,N_34869);
and U35180 (N_35180,N_34100,N_34733);
nand U35181 (N_35181,N_34135,N_34921);
xnor U35182 (N_35182,N_34312,N_34946);
or U35183 (N_35183,N_34883,N_34308);
and U35184 (N_35184,N_34545,N_34815);
xnor U35185 (N_35185,N_34639,N_34809);
xor U35186 (N_35186,N_34326,N_34282);
xor U35187 (N_35187,N_34571,N_34763);
nand U35188 (N_35188,N_34907,N_34981);
or U35189 (N_35189,N_34126,N_34329);
nand U35190 (N_35190,N_34333,N_34408);
and U35191 (N_35191,N_34101,N_34381);
and U35192 (N_35192,N_34926,N_34831);
xor U35193 (N_35193,N_34084,N_34180);
or U35194 (N_35194,N_34734,N_34631);
and U35195 (N_35195,N_34474,N_34425);
or U35196 (N_35196,N_34033,N_34274);
nand U35197 (N_35197,N_34061,N_34803);
and U35198 (N_35198,N_34433,N_34342);
and U35199 (N_35199,N_34929,N_34584);
nand U35200 (N_35200,N_34515,N_34529);
nand U35201 (N_35201,N_34790,N_34719);
and U35202 (N_35202,N_34985,N_34775);
xnor U35203 (N_35203,N_34029,N_34782);
nor U35204 (N_35204,N_34620,N_34418);
or U35205 (N_35205,N_34383,N_34048);
xnor U35206 (N_35206,N_34379,N_34280);
and U35207 (N_35207,N_34317,N_34936);
or U35208 (N_35208,N_34745,N_34315);
or U35209 (N_35209,N_34699,N_34506);
or U35210 (N_35210,N_34106,N_34518);
and U35211 (N_35211,N_34950,N_34601);
nand U35212 (N_35212,N_34473,N_34637);
and U35213 (N_35213,N_34412,N_34144);
xor U35214 (N_35214,N_34476,N_34393);
nor U35215 (N_35215,N_34933,N_34047);
nand U35216 (N_35216,N_34960,N_34575);
nor U35217 (N_35217,N_34538,N_34388);
xnor U35218 (N_35218,N_34656,N_34522);
xor U35219 (N_35219,N_34559,N_34867);
nor U35220 (N_35220,N_34503,N_34554);
and U35221 (N_35221,N_34130,N_34569);
nor U35222 (N_35222,N_34201,N_34070);
nor U35223 (N_35223,N_34844,N_34151);
nor U35224 (N_35224,N_34536,N_34035);
xnor U35225 (N_35225,N_34650,N_34791);
xnor U35226 (N_35226,N_34673,N_34796);
and U35227 (N_35227,N_34136,N_34567);
or U35228 (N_35228,N_34296,N_34129);
or U35229 (N_35229,N_34252,N_34965);
and U35230 (N_35230,N_34108,N_34092);
nand U35231 (N_35231,N_34486,N_34592);
xnor U35232 (N_35232,N_34409,N_34932);
nand U35233 (N_35233,N_34771,N_34743);
nand U35234 (N_35234,N_34969,N_34366);
and U35235 (N_35235,N_34236,N_34984);
nor U35236 (N_35236,N_34142,N_34432);
nor U35237 (N_35237,N_34124,N_34437);
or U35238 (N_35238,N_34893,N_34027);
nand U35239 (N_35239,N_34624,N_34022);
nor U35240 (N_35240,N_34896,N_34837);
nand U35241 (N_35241,N_34951,N_34140);
nor U35242 (N_35242,N_34322,N_34874);
nor U35243 (N_35243,N_34873,N_34050);
nand U35244 (N_35244,N_34930,N_34006);
xor U35245 (N_35245,N_34443,N_34483);
and U35246 (N_35246,N_34604,N_34235);
nor U35247 (N_35247,N_34660,N_34485);
nand U35248 (N_35248,N_34513,N_34043);
nand U35249 (N_35249,N_34647,N_34165);
or U35250 (N_35250,N_34666,N_34158);
nand U35251 (N_35251,N_34367,N_34888);
nand U35252 (N_35252,N_34517,N_34009);
nor U35253 (N_35253,N_34465,N_34208);
xnor U35254 (N_35254,N_34008,N_34636);
nor U35255 (N_35255,N_34478,N_34633);
nand U35256 (N_35256,N_34565,N_34210);
xor U35257 (N_35257,N_34498,N_34861);
xnor U35258 (N_35258,N_34243,N_34674);
nor U35259 (N_35259,N_34827,N_34049);
and U35260 (N_35260,N_34500,N_34054);
or U35261 (N_35261,N_34164,N_34691);
and U35262 (N_35262,N_34339,N_34832);
nand U35263 (N_35263,N_34209,N_34313);
nand U35264 (N_35264,N_34440,N_34303);
and U35265 (N_35265,N_34298,N_34064);
or U35266 (N_35266,N_34619,N_34466);
nor U35267 (N_35267,N_34871,N_34927);
and U35268 (N_35268,N_34728,N_34167);
and U35269 (N_35269,N_34786,N_34678);
nor U35270 (N_35270,N_34323,N_34847);
xor U35271 (N_35271,N_34028,N_34492);
and U35272 (N_35272,N_34477,N_34264);
or U35273 (N_35273,N_34788,N_34098);
nand U35274 (N_35274,N_34441,N_34036);
xor U35275 (N_35275,N_34910,N_34017);
xor U35276 (N_35276,N_34455,N_34230);
xnor U35277 (N_35277,N_34128,N_34372);
or U35278 (N_35278,N_34555,N_34352);
and U35279 (N_35279,N_34083,N_34696);
and U35280 (N_35280,N_34270,N_34811);
and U35281 (N_35281,N_34182,N_34875);
xnor U35282 (N_35282,N_34361,N_34038);
or U35283 (N_35283,N_34234,N_34723);
or U35284 (N_35284,N_34345,N_34808);
xnor U35285 (N_35285,N_34894,N_34341);
xnor U35286 (N_35286,N_34192,N_34458);
nor U35287 (N_35287,N_34900,N_34508);
nor U35288 (N_35288,N_34496,N_34989);
xor U35289 (N_35289,N_34954,N_34919);
nor U35290 (N_35290,N_34553,N_34975);
and U35291 (N_35291,N_34082,N_34005);
or U35292 (N_35292,N_34579,N_34495);
xnor U35293 (N_35293,N_34962,N_34431);
nor U35294 (N_35294,N_34648,N_34577);
xor U35295 (N_35295,N_34558,N_34389);
or U35296 (N_35296,N_34998,N_34977);
nor U35297 (N_35297,N_34113,N_34849);
or U35298 (N_35298,N_34789,N_34355);
nor U35299 (N_35299,N_34925,N_34958);
nand U35300 (N_35300,N_34306,N_34475);
and U35301 (N_35301,N_34681,N_34089);
nor U35302 (N_35302,N_34206,N_34598);
nor U35303 (N_35303,N_34272,N_34463);
and U35304 (N_35304,N_34152,N_34260);
xor U35305 (N_35305,N_34330,N_34846);
xor U35306 (N_35306,N_34294,N_34176);
xor U35307 (N_35307,N_34941,N_34721);
nand U35308 (N_35308,N_34768,N_34597);
or U35309 (N_35309,N_34854,N_34889);
or U35310 (N_35310,N_34324,N_34608);
and U35311 (N_35311,N_34284,N_34521);
nand U35312 (N_35312,N_34562,N_34166);
nand U35313 (N_35313,N_34697,N_34117);
nand U35314 (N_35314,N_34725,N_34840);
nor U35315 (N_35315,N_34253,N_34097);
xnor U35316 (N_35316,N_34530,N_34707);
nor U35317 (N_35317,N_34669,N_34676);
xnor U35318 (N_35318,N_34459,N_34814);
xor U35319 (N_35319,N_34149,N_34211);
and U35320 (N_35320,N_34794,N_34514);
nand U35321 (N_35321,N_34911,N_34404);
or U35322 (N_35322,N_34909,N_34179);
xnor U35323 (N_35323,N_34501,N_34599);
nand U35324 (N_35324,N_34964,N_34112);
nor U35325 (N_35325,N_34551,N_34471);
nand U35326 (N_35326,N_34879,N_34920);
nor U35327 (N_35327,N_34359,N_34855);
nor U35328 (N_35328,N_34753,N_34590);
nand U35329 (N_35329,N_34872,N_34539);
nand U35330 (N_35330,N_34007,N_34468);
nand U35331 (N_35331,N_34449,N_34972);
and U35332 (N_35332,N_34400,N_34731);
nor U35333 (N_35333,N_34414,N_34387);
xor U35334 (N_35334,N_34792,N_34710);
nor U35335 (N_35335,N_34813,N_34177);
nand U35336 (N_35336,N_34286,N_34953);
or U35337 (N_35337,N_34526,N_34645);
nand U35338 (N_35338,N_34111,N_34456);
nand U35339 (N_35339,N_34924,N_34190);
xnor U35340 (N_35340,N_34150,N_34051);
and U35341 (N_35341,N_34783,N_34748);
xnor U35342 (N_35342,N_34829,N_34607);
nor U35343 (N_35343,N_34534,N_34945);
nor U35344 (N_35344,N_34377,N_34980);
or U35345 (N_35345,N_34289,N_34003);
xor U35346 (N_35346,N_34634,N_34525);
xnor U35347 (N_35347,N_34741,N_34085);
nand U35348 (N_35348,N_34139,N_34198);
nor U35349 (N_35349,N_34580,N_34606);
nor U35350 (N_35350,N_34214,N_34689);
xnor U35351 (N_35351,N_34523,N_34516);
and U35352 (N_35352,N_34838,N_34626);
or U35353 (N_35353,N_34421,N_34663);
xor U35354 (N_35354,N_34687,N_34375);
nand U35355 (N_35355,N_34677,N_34163);
nor U35356 (N_35356,N_34332,N_34417);
nand U35357 (N_35357,N_34213,N_34770);
or U35358 (N_35358,N_34548,N_34675);
xnor U35359 (N_35359,N_34703,N_34603);
nor U35360 (N_35360,N_34480,N_34754);
or U35361 (N_35361,N_34183,N_34016);
nor U35362 (N_35362,N_34995,N_34278);
or U35363 (N_35363,N_34481,N_34334);
nor U35364 (N_35364,N_34429,N_34785);
and U35365 (N_35365,N_34020,N_34320);
or U35366 (N_35366,N_34451,N_34724);
nor U35367 (N_35367,N_34300,N_34878);
and U35368 (N_35368,N_34172,N_34090);
nor U35369 (N_35369,N_34563,N_34075);
nor U35370 (N_35370,N_34197,N_34134);
and U35371 (N_35371,N_34229,N_34067);
nand U35372 (N_35372,N_34644,N_34668);
and U35373 (N_35373,N_34291,N_34227);
nand U35374 (N_35374,N_34658,N_34751);
and U35375 (N_35375,N_34842,N_34744);
nand U35376 (N_35376,N_34277,N_34216);
nor U35377 (N_35377,N_34961,N_34693);
or U35378 (N_35378,N_34026,N_34948);
nand U35379 (N_35379,N_34187,N_34806);
or U35380 (N_35380,N_34766,N_34966);
and U35381 (N_35381,N_34761,N_34304);
nor U35382 (N_35382,N_34750,N_34073);
or U35383 (N_35383,N_34662,N_34795);
xor U35384 (N_35384,N_34736,N_34646);
nor U35385 (N_35385,N_34205,N_34934);
nor U35386 (N_35386,N_34392,N_34535);
nor U35387 (N_35387,N_34613,N_34068);
nor U35388 (N_35388,N_34266,N_34249);
nor U35389 (N_35389,N_34578,N_34757);
nor U35390 (N_35390,N_34335,N_34922);
nor U35391 (N_35391,N_34314,N_34618);
nand U35392 (N_35392,N_34640,N_34340);
or U35393 (N_35393,N_34781,N_34560);
and U35394 (N_35394,N_34755,N_34701);
nand U35395 (N_35395,N_34708,N_34263);
and U35396 (N_35396,N_34220,N_34833);
or U35397 (N_35397,N_34540,N_34202);
or U35398 (N_35398,N_34328,N_34735);
nand U35399 (N_35399,N_34858,N_34586);
xnor U35400 (N_35400,N_34593,N_34066);
and U35401 (N_35401,N_34489,N_34990);
or U35402 (N_35402,N_34729,N_34488);
xnor U35403 (N_35403,N_34103,N_34060);
nand U35404 (N_35404,N_34058,N_34232);
nor U35405 (N_35405,N_34931,N_34110);
or U35406 (N_35406,N_34820,N_34572);
nor U35407 (N_35407,N_34088,N_34732);
or U35408 (N_35408,N_34145,N_34141);
nand U35409 (N_35409,N_34510,N_34188);
nor U35410 (N_35410,N_34881,N_34845);
xor U35411 (N_35411,N_34877,N_34683);
nand U35412 (N_35412,N_34839,N_34240);
or U35413 (N_35413,N_34614,N_34543);
nor U35414 (N_35414,N_34887,N_34457);
xnor U35415 (N_35415,N_34245,N_34974);
nor U35416 (N_35416,N_34824,N_34852);
or U35417 (N_35417,N_34157,N_34074);
or U35418 (N_35418,N_34561,N_34493);
and U35419 (N_35419,N_34378,N_34602);
nor U35420 (N_35420,N_34122,N_34583);
xnor U35421 (N_35421,N_34311,N_34081);
or U35422 (N_35422,N_34299,N_34573);
xnor U35423 (N_35423,N_34133,N_34589);
and U35424 (N_35424,N_34426,N_34261);
or U35425 (N_35425,N_34903,N_34630);
nor U35426 (N_35426,N_34643,N_34700);
nand U35427 (N_35427,N_34797,N_34305);
xnor U35428 (N_35428,N_34063,N_34830);
nor U35429 (N_35429,N_34199,N_34566);
and U35430 (N_35430,N_34376,N_34096);
xor U35431 (N_35431,N_34200,N_34403);
and U35432 (N_35432,N_34520,N_34801);
nor U35433 (N_35433,N_34402,N_34542);
and U35434 (N_35434,N_34116,N_34276);
or U35435 (N_35435,N_34325,N_34221);
nor U35436 (N_35436,N_34605,N_34611);
and U35437 (N_35437,N_34641,N_34385);
nor U35438 (N_35438,N_34479,N_34986);
nor U35439 (N_35439,N_34870,N_34541);
nand U35440 (N_35440,N_34226,N_34053);
nor U35441 (N_35441,N_34161,N_34918);
nand U35442 (N_35442,N_34502,N_34071);
or U35443 (N_35443,N_34776,N_34024);
and U35444 (N_35444,N_34297,N_34859);
or U35445 (N_35445,N_34714,N_34692);
nor U35446 (N_35446,N_34942,N_34665);
nand U35447 (N_35447,N_34747,N_34095);
xnor U35448 (N_35448,N_34450,N_34453);
xor U35449 (N_35449,N_34031,N_34374);
and U35450 (N_35450,N_34591,N_34740);
and U35451 (N_35451,N_34013,N_34265);
nor U35452 (N_35452,N_34722,N_34857);
and U35453 (N_35453,N_34667,N_34454);
xor U35454 (N_35454,N_34629,N_34670);
xnor U35455 (N_35455,N_34384,N_34596);
and U35456 (N_35456,N_34905,N_34428);
xnor U35457 (N_35457,N_34627,N_34595);
nand U35458 (N_35458,N_34713,N_34121);
and U35459 (N_35459,N_34928,N_34726);
or U35460 (N_35460,N_34032,N_34319);
and U35461 (N_35461,N_34174,N_34826);
nor U35462 (N_35462,N_34682,N_34661);
xnor U35463 (N_35463,N_34344,N_34461);
nor U35464 (N_35464,N_34497,N_34448);
nor U35465 (N_35465,N_34979,N_34679);
nand U35466 (N_35466,N_34991,N_34600);
nor U35467 (N_35467,N_34730,N_34039);
nand U35468 (N_35468,N_34030,N_34937);
xor U35469 (N_35469,N_34348,N_34078);
or U35470 (N_35470,N_34866,N_34354);
and U35471 (N_35471,N_34570,N_34360);
xor U35472 (N_35472,N_34464,N_34127);
or U35473 (N_35473,N_34821,N_34509);
and U35474 (N_35474,N_34273,N_34460);
nor U35475 (N_35475,N_34146,N_34407);
xnor U35476 (N_35476,N_34037,N_34225);
nor U35477 (N_35477,N_34671,N_34369);
nand U35478 (N_35478,N_34898,N_34649);
nand U35479 (N_35479,N_34818,N_34445);
nor U35480 (N_35480,N_34904,N_34065);
nor U35481 (N_35481,N_34684,N_34491);
nand U35482 (N_35482,N_34002,N_34285);
nand U35483 (N_35483,N_34439,N_34585);
or U35484 (N_35484,N_34115,N_34807);
nand U35485 (N_35485,N_34892,N_34452);
nand U35486 (N_35486,N_34250,N_34076);
xnor U35487 (N_35487,N_34738,N_34762);
nor U35488 (N_35488,N_34382,N_34010);
and U35489 (N_35489,N_34435,N_34856);
xnor U35490 (N_35490,N_34652,N_34091);
or U35491 (N_35491,N_34628,N_34046);
and U35492 (N_35492,N_34702,N_34715);
nand U35493 (N_35493,N_34653,N_34970);
and U35494 (N_35494,N_34915,N_34462);
nor U35495 (N_35495,N_34737,N_34823);
or U35496 (N_35496,N_34430,N_34267);
nand U35497 (N_35497,N_34102,N_34447);
and U35498 (N_35498,N_34914,N_34292);
and U35499 (N_35499,N_34415,N_34159);
xnor U35500 (N_35500,N_34392,N_34238);
xor U35501 (N_35501,N_34359,N_34848);
xor U35502 (N_35502,N_34666,N_34865);
and U35503 (N_35503,N_34796,N_34604);
nand U35504 (N_35504,N_34759,N_34526);
and U35505 (N_35505,N_34022,N_34239);
nor U35506 (N_35506,N_34245,N_34199);
nor U35507 (N_35507,N_34070,N_34405);
nor U35508 (N_35508,N_34034,N_34408);
nand U35509 (N_35509,N_34213,N_34268);
nand U35510 (N_35510,N_34365,N_34802);
or U35511 (N_35511,N_34622,N_34926);
or U35512 (N_35512,N_34857,N_34682);
xnor U35513 (N_35513,N_34088,N_34442);
and U35514 (N_35514,N_34115,N_34091);
and U35515 (N_35515,N_34395,N_34595);
nand U35516 (N_35516,N_34795,N_34852);
xnor U35517 (N_35517,N_34699,N_34024);
or U35518 (N_35518,N_34872,N_34485);
and U35519 (N_35519,N_34761,N_34572);
nor U35520 (N_35520,N_34322,N_34521);
xor U35521 (N_35521,N_34130,N_34629);
nor U35522 (N_35522,N_34571,N_34673);
nor U35523 (N_35523,N_34160,N_34032);
or U35524 (N_35524,N_34861,N_34335);
nand U35525 (N_35525,N_34237,N_34440);
nor U35526 (N_35526,N_34584,N_34412);
xor U35527 (N_35527,N_34863,N_34742);
or U35528 (N_35528,N_34342,N_34263);
nor U35529 (N_35529,N_34469,N_34424);
nand U35530 (N_35530,N_34448,N_34814);
xor U35531 (N_35531,N_34220,N_34465);
xnor U35532 (N_35532,N_34550,N_34776);
nand U35533 (N_35533,N_34499,N_34258);
and U35534 (N_35534,N_34761,N_34868);
xor U35535 (N_35535,N_34185,N_34166);
nor U35536 (N_35536,N_34698,N_34440);
xor U35537 (N_35537,N_34672,N_34261);
xor U35538 (N_35538,N_34544,N_34913);
and U35539 (N_35539,N_34132,N_34258);
and U35540 (N_35540,N_34667,N_34309);
xnor U35541 (N_35541,N_34775,N_34120);
nor U35542 (N_35542,N_34826,N_34018);
nand U35543 (N_35543,N_34223,N_34370);
nand U35544 (N_35544,N_34924,N_34221);
nand U35545 (N_35545,N_34747,N_34227);
nand U35546 (N_35546,N_34934,N_34430);
nor U35547 (N_35547,N_34410,N_34319);
nand U35548 (N_35548,N_34690,N_34386);
or U35549 (N_35549,N_34856,N_34152);
and U35550 (N_35550,N_34760,N_34825);
and U35551 (N_35551,N_34258,N_34124);
and U35552 (N_35552,N_34107,N_34575);
xnor U35553 (N_35553,N_34627,N_34986);
nand U35554 (N_35554,N_34294,N_34165);
nor U35555 (N_35555,N_34228,N_34232);
xnor U35556 (N_35556,N_34333,N_34948);
and U35557 (N_35557,N_34005,N_34647);
xnor U35558 (N_35558,N_34548,N_34549);
nor U35559 (N_35559,N_34810,N_34383);
nor U35560 (N_35560,N_34638,N_34438);
or U35561 (N_35561,N_34127,N_34873);
xor U35562 (N_35562,N_34523,N_34243);
or U35563 (N_35563,N_34281,N_34820);
nand U35564 (N_35564,N_34886,N_34245);
or U35565 (N_35565,N_34662,N_34513);
nand U35566 (N_35566,N_34355,N_34720);
nand U35567 (N_35567,N_34000,N_34674);
xnor U35568 (N_35568,N_34120,N_34520);
and U35569 (N_35569,N_34752,N_34561);
xor U35570 (N_35570,N_34175,N_34985);
xor U35571 (N_35571,N_34810,N_34654);
xor U35572 (N_35572,N_34073,N_34342);
or U35573 (N_35573,N_34073,N_34697);
xor U35574 (N_35574,N_34687,N_34888);
nand U35575 (N_35575,N_34086,N_34644);
nand U35576 (N_35576,N_34193,N_34102);
and U35577 (N_35577,N_34115,N_34478);
nand U35578 (N_35578,N_34398,N_34705);
or U35579 (N_35579,N_34503,N_34717);
and U35580 (N_35580,N_34895,N_34449);
nor U35581 (N_35581,N_34424,N_34580);
or U35582 (N_35582,N_34365,N_34618);
nor U35583 (N_35583,N_34766,N_34632);
nor U35584 (N_35584,N_34435,N_34842);
xor U35585 (N_35585,N_34504,N_34901);
nand U35586 (N_35586,N_34792,N_34511);
nand U35587 (N_35587,N_34293,N_34606);
or U35588 (N_35588,N_34124,N_34985);
or U35589 (N_35589,N_34200,N_34542);
nand U35590 (N_35590,N_34701,N_34304);
and U35591 (N_35591,N_34887,N_34389);
or U35592 (N_35592,N_34047,N_34469);
and U35593 (N_35593,N_34360,N_34875);
nand U35594 (N_35594,N_34349,N_34359);
nand U35595 (N_35595,N_34057,N_34312);
xor U35596 (N_35596,N_34857,N_34647);
or U35597 (N_35597,N_34655,N_34822);
nand U35598 (N_35598,N_34270,N_34931);
xor U35599 (N_35599,N_34625,N_34172);
nor U35600 (N_35600,N_34540,N_34974);
and U35601 (N_35601,N_34228,N_34639);
and U35602 (N_35602,N_34625,N_34324);
and U35603 (N_35603,N_34362,N_34027);
or U35604 (N_35604,N_34311,N_34105);
nand U35605 (N_35605,N_34455,N_34065);
nand U35606 (N_35606,N_34707,N_34273);
nor U35607 (N_35607,N_34088,N_34627);
nand U35608 (N_35608,N_34198,N_34050);
nand U35609 (N_35609,N_34144,N_34419);
xnor U35610 (N_35610,N_34461,N_34447);
and U35611 (N_35611,N_34484,N_34056);
nand U35612 (N_35612,N_34831,N_34045);
and U35613 (N_35613,N_34717,N_34223);
nor U35614 (N_35614,N_34387,N_34745);
nand U35615 (N_35615,N_34267,N_34372);
xor U35616 (N_35616,N_34625,N_34033);
nor U35617 (N_35617,N_34650,N_34350);
and U35618 (N_35618,N_34209,N_34108);
nor U35619 (N_35619,N_34840,N_34327);
nor U35620 (N_35620,N_34703,N_34869);
nand U35621 (N_35621,N_34346,N_34255);
and U35622 (N_35622,N_34054,N_34887);
or U35623 (N_35623,N_34978,N_34431);
nor U35624 (N_35624,N_34692,N_34803);
nand U35625 (N_35625,N_34863,N_34795);
or U35626 (N_35626,N_34481,N_34337);
or U35627 (N_35627,N_34416,N_34170);
nand U35628 (N_35628,N_34939,N_34512);
nand U35629 (N_35629,N_34379,N_34900);
nor U35630 (N_35630,N_34751,N_34385);
nor U35631 (N_35631,N_34240,N_34630);
and U35632 (N_35632,N_34004,N_34860);
nand U35633 (N_35633,N_34921,N_34779);
xor U35634 (N_35634,N_34041,N_34500);
or U35635 (N_35635,N_34660,N_34845);
xnor U35636 (N_35636,N_34167,N_34757);
xnor U35637 (N_35637,N_34630,N_34747);
nand U35638 (N_35638,N_34313,N_34525);
or U35639 (N_35639,N_34182,N_34892);
nand U35640 (N_35640,N_34930,N_34212);
nand U35641 (N_35641,N_34492,N_34517);
or U35642 (N_35642,N_34222,N_34428);
nor U35643 (N_35643,N_34716,N_34205);
nand U35644 (N_35644,N_34726,N_34716);
xnor U35645 (N_35645,N_34486,N_34534);
and U35646 (N_35646,N_34632,N_34338);
and U35647 (N_35647,N_34597,N_34428);
nor U35648 (N_35648,N_34687,N_34222);
nand U35649 (N_35649,N_34863,N_34693);
or U35650 (N_35650,N_34722,N_34344);
or U35651 (N_35651,N_34909,N_34904);
nor U35652 (N_35652,N_34395,N_34633);
and U35653 (N_35653,N_34652,N_34566);
nand U35654 (N_35654,N_34050,N_34274);
nand U35655 (N_35655,N_34491,N_34072);
nand U35656 (N_35656,N_34488,N_34564);
nor U35657 (N_35657,N_34950,N_34791);
or U35658 (N_35658,N_34544,N_34136);
or U35659 (N_35659,N_34485,N_34005);
nand U35660 (N_35660,N_34730,N_34347);
xor U35661 (N_35661,N_34675,N_34421);
nor U35662 (N_35662,N_34733,N_34169);
nor U35663 (N_35663,N_34903,N_34174);
or U35664 (N_35664,N_34457,N_34159);
and U35665 (N_35665,N_34351,N_34892);
and U35666 (N_35666,N_34539,N_34769);
or U35667 (N_35667,N_34196,N_34345);
nor U35668 (N_35668,N_34182,N_34358);
nor U35669 (N_35669,N_34117,N_34128);
xor U35670 (N_35670,N_34075,N_34182);
or U35671 (N_35671,N_34726,N_34987);
nor U35672 (N_35672,N_34952,N_34679);
nor U35673 (N_35673,N_34655,N_34441);
and U35674 (N_35674,N_34877,N_34440);
nand U35675 (N_35675,N_34428,N_34533);
nand U35676 (N_35676,N_34522,N_34136);
or U35677 (N_35677,N_34717,N_34569);
nor U35678 (N_35678,N_34869,N_34242);
and U35679 (N_35679,N_34142,N_34765);
and U35680 (N_35680,N_34528,N_34697);
xnor U35681 (N_35681,N_34377,N_34817);
nor U35682 (N_35682,N_34059,N_34254);
nand U35683 (N_35683,N_34910,N_34976);
or U35684 (N_35684,N_34101,N_34670);
and U35685 (N_35685,N_34566,N_34103);
nor U35686 (N_35686,N_34079,N_34638);
or U35687 (N_35687,N_34661,N_34442);
nor U35688 (N_35688,N_34583,N_34831);
xor U35689 (N_35689,N_34820,N_34164);
xor U35690 (N_35690,N_34718,N_34403);
nor U35691 (N_35691,N_34956,N_34189);
or U35692 (N_35692,N_34988,N_34186);
and U35693 (N_35693,N_34333,N_34163);
or U35694 (N_35694,N_34049,N_34231);
nand U35695 (N_35695,N_34629,N_34581);
nand U35696 (N_35696,N_34587,N_34633);
xnor U35697 (N_35697,N_34218,N_34136);
and U35698 (N_35698,N_34510,N_34777);
nand U35699 (N_35699,N_34142,N_34824);
and U35700 (N_35700,N_34759,N_34566);
and U35701 (N_35701,N_34462,N_34058);
nand U35702 (N_35702,N_34135,N_34731);
nand U35703 (N_35703,N_34396,N_34506);
nand U35704 (N_35704,N_34983,N_34494);
or U35705 (N_35705,N_34680,N_34952);
nor U35706 (N_35706,N_34648,N_34724);
and U35707 (N_35707,N_34616,N_34270);
nor U35708 (N_35708,N_34246,N_34421);
nor U35709 (N_35709,N_34386,N_34562);
and U35710 (N_35710,N_34975,N_34008);
or U35711 (N_35711,N_34931,N_34081);
nand U35712 (N_35712,N_34390,N_34278);
nor U35713 (N_35713,N_34892,N_34489);
and U35714 (N_35714,N_34079,N_34002);
and U35715 (N_35715,N_34327,N_34864);
nand U35716 (N_35716,N_34561,N_34326);
xnor U35717 (N_35717,N_34105,N_34451);
nor U35718 (N_35718,N_34949,N_34240);
xnor U35719 (N_35719,N_34042,N_34156);
nand U35720 (N_35720,N_34892,N_34760);
nor U35721 (N_35721,N_34251,N_34384);
nor U35722 (N_35722,N_34941,N_34092);
and U35723 (N_35723,N_34891,N_34584);
or U35724 (N_35724,N_34369,N_34846);
or U35725 (N_35725,N_34303,N_34252);
nand U35726 (N_35726,N_34259,N_34514);
and U35727 (N_35727,N_34135,N_34931);
or U35728 (N_35728,N_34308,N_34587);
nor U35729 (N_35729,N_34996,N_34184);
or U35730 (N_35730,N_34134,N_34226);
nor U35731 (N_35731,N_34675,N_34796);
and U35732 (N_35732,N_34249,N_34294);
or U35733 (N_35733,N_34571,N_34919);
and U35734 (N_35734,N_34262,N_34902);
and U35735 (N_35735,N_34102,N_34807);
nand U35736 (N_35736,N_34142,N_34427);
nand U35737 (N_35737,N_34196,N_34480);
nand U35738 (N_35738,N_34170,N_34972);
nand U35739 (N_35739,N_34669,N_34796);
xor U35740 (N_35740,N_34006,N_34220);
and U35741 (N_35741,N_34171,N_34161);
and U35742 (N_35742,N_34236,N_34240);
xnor U35743 (N_35743,N_34434,N_34719);
or U35744 (N_35744,N_34337,N_34954);
nor U35745 (N_35745,N_34957,N_34918);
nor U35746 (N_35746,N_34769,N_34723);
nor U35747 (N_35747,N_34910,N_34752);
nor U35748 (N_35748,N_34113,N_34753);
xnor U35749 (N_35749,N_34082,N_34055);
nor U35750 (N_35750,N_34333,N_34653);
and U35751 (N_35751,N_34226,N_34992);
nand U35752 (N_35752,N_34962,N_34041);
and U35753 (N_35753,N_34600,N_34998);
and U35754 (N_35754,N_34547,N_34923);
nand U35755 (N_35755,N_34812,N_34318);
and U35756 (N_35756,N_34838,N_34894);
or U35757 (N_35757,N_34874,N_34176);
or U35758 (N_35758,N_34054,N_34569);
or U35759 (N_35759,N_34093,N_34724);
nand U35760 (N_35760,N_34875,N_34089);
nand U35761 (N_35761,N_34554,N_34678);
or U35762 (N_35762,N_34642,N_34603);
and U35763 (N_35763,N_34157,N_34497);
nor U35764 (N_35764,N_34835,N_34879);
and U35765 (N_35765,N_34445,N_34197);
nand U35766 (N_35766,N_34661,N_34395);
or U35767 (N_35767,N_34803,N_34178);
and U35768 (N_35768,N_34224,N_34738);
or U35769 (N_35769,N_34389,N_34573);
xor U35770 (N_35770,N_34265,N_34469);
and U35771 (N_35771,N_34207,N_34093);
xnor U35772 (N_35772,N_34902,N_34817);
nor U35773 (N_35773,N_34571,N_34277);
nand U35774 (N_35774,N_34707,N_34345);
or U35775 (N_35775,N_34192,N_34140);
nand U35776 (N_35776,N_34203,N_34231);
or U35777 (N_35777,N_34727,N_34409);
or U35778 (N_35778,N_34735,N_34441);
and U35779 (N_35779,N_34971,N_34081);
xor U35780 (N_35780,N_34191,N_34831);
nor U35781 (N_35781,N_34196,N_34123);
xor U35782 (N_35782,N_34506,N_34819);
xor U35783 (N_35783,N_34451,N_34234);
nor U35784 (N_35784,N_34809,N_34565);
and U35785 (N_35785,N_34513,N_34719);
xor U35786 (N_35786,N_34346,N_34500);
and U35787 (N_35787,N_34154,N_34586);
xnor U35788 (N_35788,N_34118,N_34934);
and U35789 (N_35789,N_34601,N_34479);
or U35790 (N_35790,N_34843,N_34738);
nand U35791 (N_35791,N_34839,N_34921);
xnor U35792 (N_35792,N_34736,N_34950);
or U35793 (N_35793,N_34598,N_34036);
xnor U35794 (N_35794,N_34558,N_34139);
nor U35795 (N_35795,N_34810,N_34281);
xor U35796 (N_35796,N_34405,N_34889);
or U35797 (N_35797,N_34017,N_34378);
and U35798 (N_35798,N_34374,N_34141);
and U35799 (N_35799,N_34918,N_34871);
xnor U35800 (N_35800,N_34364,N_34457);
or U35801 (N_35801,N_34521,N_34603);
and U35802 (N_35802,N_34238,N_34689);
nor U35803 (N_35803,N_34829,N_34390);
xor U35804 (N_35804,N_34980,N_34694);
nor U35805 (N_35805,N_34115,N_34639);
nor U35806 (N_35806,N_34493,N_34946);
nand U35807 (N_35807,N_34473,N_34525);
nand U35808 (N_35808,N_34028,N_34430);
xnor U35809 (N_35809,N_34478,N_34935);
and U35810 (N_35810,N_34311,N_34188);
or U35811 (N_35811,N_34759,N_34397);
and U35812 (N_35812,N_34037,N_34581);
xnor U35813 (N_35813,N_34061,N_34843);
nor U35814 (N_35814,N_34285,N_34832);
nand U35815 (N_35815,N_34259,N_34333);
or U35816 (N_35816,N_34763,N_34280);
nand U35817 (N_35817,N_34874,N_34733);
and U35818 (N_35818,N_34360,N_34116);
nor U35819 (N_35819,N_34909,N_34860);
or U35820 (N_35820,N_34635,N_34582);
xor U35821 (N_35821,N_34364,N_34892);
xor U35822 (N_35822,N_34785,N_34239);
xor U35823 (N_35823,N_34971,N_34479);
xor U35824 (N_35824,N_34922,N_34539);
nand U35825 (N_35825,N_34040,N_34884);
nand U35826 (N_35826,N_34032,N_34128);
nor U35827 (N_35827,N_34193,N_34198);
nand U35828 (N_35828,N_34877,N_34623);
nor U35829 (N_35829,N_34188,N_34357);
nand U35830 (N_35830,N_34146,N_34336);
nand U35831 (N_35831,N_34179,N_34313);
and U35832 (N_35832,N_34626,N_34033);
and U35833 (N_35833,N_34200,N_34938);
nor U35834 (N_35834,N_34029,N_34862);
nand U35835 (N_35835,N_34838,N_34487);
and U35836 (N_35836,N_34792,N_34282);
nor U35837 (N_35837,N_34150,N_34411);
nor U35838 (N_35838,N_34727,N_34234);
xnor U35839 (N_35839,N_34125,N_34877);
nor U35840 (N_35840,N_34154,N_34657);
xnor U35841 (N_35841,N_34342,N_34656);
and U35842 (N_35842,N_34831,N_34048);
nor U35843 (N_35843,N_34894,N_34778);
xor U35844 (N_35844,N_34266,N_34514);
or U35845 (N_35845,N_34302,N_34538);
and U35846 (N_35846,N_34103,N_34268);
or U35847 (N_35847,N_34652,N_34310);
and U35848 (N_35848,N_34085,N_34607);
or U35849 (N_35849,N_34148,N_34942);
xnor U35850 (N_35850,N_34611,N_34892);
nor U35851 (N_35851,N_34754,N_34777);
xor U35852 (N_35852,N_34419,N_34357);
nor U35853 (N_35853,N_34006,N_34708);
nand U35854 (N_35854,N_34585,N_34321);
or U35855 (N_35855,N_34376,N_34269);
nor U35856 (N_35856,N_34507,N_34413);
xor U35857 (N_35857,N_34591,N_34635);
nor U35858 (N_35858,N_34314,N_34170);
nor U35859 (N_35859,N_34521,N_34967);
and U35860 (N_35860,N_34045,N_34834);
or U35861 (N_35861,N_34580,N_34106);
xor U35862 (N_35862,N_34116,N_34583);
nand U35863 (N_35863,N_34671,N_34735);
and U35864 (N_35864,N_34982,N_34237);
xor U35865 (N_35865,N_34359,N_34215);
nor U35866 (N_35866,N_34048,N_34435);
and U35867 (N_35867,N_34705,N_34687);
xor U35868 (N_35868,N_34063,N_34795);
xnor U35869 (N_35869,N_34467,N_34231);
nor U35870 (N_35870,N_34689,N_34128);
nand U35871 (N_35871,N_34584,N_34770);
nor U35872 (N_35872,N_34986,N_34718);
xor U35873 (N_35873,N_34567,N_34860);
nor U35874 (N_35874,N_34909,N_34814);
xor U35875 (N_35875,N_34741,N_34261);
or U35876 (N_35876,N_34130,N_34926);
nor U35877 (N_35877,N_34908,N_34339);
nand U35878 (N_35878,N_34622,N_34371);
nand U35879 (N_35879,N_34595,N_34799);
or U35880 (N_35880,N_34784,N_34210);
xor U35881 (N_35881,N_34301,N_34067);
xnor U35882 (N_35882,N_34733,N_34677);
xnor U35883 (N_35883,N_34185,N_34467);
nor U35884 (N_35884,N_34055,N_34808);
nor U35885 (N_35885,N_34833,N_34022);
xnor U35886 (N_35886,N_34004,N_34095);
nand U35887 (N_35887,N_34804,N_34459);
nand U35888 (N_35888,N_34221,N_34808);
nor U35889 (N_35889,N_34638,N_34300);
or U35890 (N_35890,N_34219,N_34383);
nand U35891 (N_35891,N_34841,N_34790);
nand U35892 (N_35892,N_34925,N_34156);
and U35893 (N_35893,N_34647,N_34535);
nor U35894 (N_35894,N_34966,N_34531);
or U35895 (N_35895,N_34364,N_34107);
and U35896 (N_35896,N_34555,N_34907);
nor U35897 (N_35897,N_34377,N_34319);
nand U35898 (N_35898,N_34954,N_34496);
or U35899 (N_35899,N_34601,N_34895);
xor U35900 (N_35900,N_34584,N_34896);
or U35901 (N_35901,N_34221,N_34886);
and U35902 (N_35902,N_34382,N_34640);
or U35903 (N_35903,N_34622,N_34013);
xnor U35904 (N_35904,N_34476,N_34720);
nand U35905 (N_35905,N_34239,N_34038);
nor U35906 (N_35906,N_34410,N_34579);
and U35907 (N_35907,N_34229,N_34108);
xor U35908 (N_35908,N_34548,N_34846);
and U35909 (N_35909,N_34956,N_34412);
nand U35910 (N_35910,N_34699,N_34175);
xnor U35911 (N_35911,N_34126,N_34143);
and U35912 (N_35912,N_34847,N_34544);
and U35913 (N_35913,N_34145,N_34548);
or U35914 (N_35914,N_34682,N_34266);
xor U35915 (N_35915,N_34752,N_34019);
xnor U35916 (N_35916,N_34325,N_34297);
xnor U35917 (N_35917,N_34685,N_34184);
xor U35918 (N_35918,N_34781,N_34196);
and U35919 (N_35919,N_34468,N_34922);
and U35920 (N_35920,N_34584,N_34658);
xor U35921 (N_35921,N_34866,N_34704);
and U35922 (N_35922,N_34933,N_34704);
or U35923 (N_35923,N_34394,N_34238);
and U35924 (N_35924,N_34284,N_34516);
or U35925 (N_35925,N_34531,N_34645);
and U35926 (N_35926,N_34458,N_34742);
xnor U35927 (N_35927,N_34884,N_34475);
nor U35928 (N_35928,N_34137,N_34701);
xor U35929 (N_35929,N_34098,N_34768);
xor U35930 (N_35930,N_34786,N_34309);
and U35931 (N_35931,N_34573,N_34353);
and U35932 (N_35932,N_34648,N_34132);
and U35933 (N_35933,N_34029,N_34089);
nor U35934 (N_35934,N_34695,N_34285);
or U35935 (N_35935,N_34571,N_34391);
nand U35936 (N_35936,N_34544,N_34405);
nor U35937 (N_35937,N_34647,N_34006);
nor U35938 (N_35938,N_34287,N_34385);
xnor U35939 (N_35939,N_34838,N_34068);
nand U35940 (N_35940,N_34975,N_34048);
and U35941 (N_35941,N_34419,N_34154);
and U35942 (N_35942,N_34714,N_34530);
nand U35943 (N_35943,N_34434,N_34864);
xnor U35944 (N_35944,N_34598,N_34994);
nand U35945 (N_35945,N_34128,N_34285);
nand U35946 (N_35946,N_34655,N_34604);
and U35947 (N_35947,N_34526,N_34478);
nor U35948 (N_35948,N_34090,N_34811);
or U35949 (N_35949,N_34993,N_34834);
nor U35950 (N_35950,N_34354,N_34588);
and U35951 (N_35951,N_34254,N_34511);
nand U35952 (N_35952,N_34463,N_34500);
nand U35953 (N_35953,N_34902,N_34111);
nand U35954 (N_35954,N_34075,N_34073);
and U35955 (N_35955,N_34345,N_34719);
xor U35956 (N_35956,N_34985,N_34494);
nor U35957 (N_35957,N_34587,N_34017);
and U35958 (N_35958,N_34356,N_34329);
and U35959 (N_35959,N_34240,N_34793);
or U35960 (N_35960,N_34778,N_34981);
nor U35961 (N_35961,N_34542,N_34902);
nand U35962 (N_35962,N_34067,N_34705);
xnor U35963 (N_35963,N_34627,N_34781);
xor U35964 (N_35964,N_34608,N_34165);
nor U35965 (N_35965,N_34276,N_34194);
nor U35966 (N_35966,N_34648,N_34663);
nand U35967 (N_35967,N_34980,N_34865);
xnor U35968 (N_35968,N_34823,N_34742);
or U35969 (N_35969,N_34474,N_34083);
nor U35970 (N_35970,N_34766,N_34073);
or U35971 (N_35971,N_34075,N_34550);
nand U35972 (N_35972,N_34440,N_34604);
or U35973 (N_35973,N_34743,N_34204);
or U35974 (N_35974,N_34004,N_34943);
and U35975 (N_35975,N_34357,N_34890);
xor U35976 (N_35976,N_34044,N_34846);
nand U35977 (N_35977,N_34476,N_34468);
or U35978 (N_35978,N_34488,N_34414);
and U35979 (N_35979,N_34062,N_34881);
nand U35980 (N_35980,N_34114,N_34659);
xor U35981 (N_35981,N_34163,N_34331);
and U35982 (N_35982,N_34163,N_34081);
nor U35983 (N_35983,N_34931,N_34609);
xnor U35984 (N_35984,N_34541,N_34719);
xnor U35985 (N_35985,N_34785,N_34449);
and U35986 (N_35986,N_34560,N_34082);
nor U35987 (N_35987,N_34880,N_34238);
nor U35988 (N_35988,N_34326,N_34598);
and U35989 (N_35989,N_34794,N_34868);
or U35990 (N_35990,N_34848,N_34664);
nand U35991 (N_35991,N_34088,N_34378);
nand U35992 (N_35992,N_34546,N_34181);
nor U35993 (N_35993,N_34121,N_34644);
and U35994 (N_35994,N_34433,N_34653);
and U35995 (N_35995,N_34440,N_34476);
nand U35996 (N_35996,N_34300,N_34876);
nor U35997 (N_35997,N_34798,N_34383);
nand U35998 (N_35998,N_34018,N_34857);
nor U35999 (N_35999,N_34985,N_34726);
nand U36000 (N_36000,N_35954,N_35843);
xor U36001 (N_36001,N_35257,N_35834);
and U36002 (N_36002,N_35025,N_35498);
nand U36003 (N_36003,N_35511,N_35701);
nor U36004 (N_36004,N_35900,N_35094);
xnor U36005 (N_36005,N_35659,N_35279);
xor U36006 (N_36006,N_35083,N_35248);
nand U36007 (N_36007,N_35217,N_35946);
nand U36008 (N_36008,N_35018,N_35532);
nor U36009 (N_36009,N_35499,N_35693);
nor U36010 (N_36010,N_35036,N_35238);
xnor U36011 (N_36011,N_35544,N_35557);
nor U36012 (N_36012,N_35522,N_35576);
nand U36013 (N_36013,N_35844,N_35674);
nand U36014 (N_36014,N_35986,N_35491);
xor U36015 (N_36015,N_35836,N_35420);
xor U36016 (N_36016,N_35088,N_35135);
nor U36017 (N_36017,N_35044,N_35876);
or U36018 (N_36018,N_35479,N_35197);
nand U36019 (N_36019,N_35541,N_35004);
or U36020 (N_36020,N_35097,N_35235);
xor U36021 (N_36021,N_35917,N_35651);
or U36022 (N_36022,N_35289,N_35863);
nand U36023 (N_36023,N_35410,N_35942);
or U36024 (N_36024,N_35333,N_35650);
and U36025 (N_36025,N_35377,N_35294);
or U36026 (N_36026,N_35202,N_35793);
nor U36027 (N_36027,N_35446,N_35787);
xor U36028 (N_36028,N_35928,N_35266);
nand U36029 (N_36029,N_35883,N_35429);
or U36030 (N_36030,N_35280,N_35821);
nor U36031 (N_36031,N_35107,N_35330);
and U36032 (N_36032,N_35108,N_35380);
or U36033 (N_36033,N_35934,N_35551);
or U36034 (N_36034,N_35073,N_35221);
nor U36035 (N_36035,N_35205,N_35345);
xnor U36036 (N_36036,N_35118,N_35148);
and U36037 (N_36037,N_35902,N_35190);
nand U36038 (N_36038,N_35658,N_35966);
and U36039 (N_36039,N_35478,N_35709);
xnor U36040 (N_36040,N_35213,N_35937);
and U36041 (N_36041,N_35791,N_35014);
nand U36042 (N_36042,N_35628,N_35381);
xnor U36043 (N_36043,N_35979,N_35818);
and U36044 (N_36044,N_35944,N_35906);
or U36045 (N_36045,N_35050,N_35058);
xnor U36046 (N_36046,N_35846,N_35936);
nand U36047 (N_36047,N_35458,N_35562);
xor U36048 (N_36048,N_35495,N_35868);
or U36049 (N_36049,N_35961,N_35521);
nor U36050 (N_36050,N_35677,N_35518);
xnor U36051 (N_36051,N_35907,N_35820);
xnor U36052 (N_36052,N_35201,N_35357);
or U36053 (N_36053,N_35375,N_35462);
nor U36054 (N_36054,N_35657,N_35126);
xnor U36055 (N_36055,N_35363,N_35593);
and U36056 (N_36056,N_35922,N_35131);
xor U36057 (N_36057,N_35500,N_35168);
and U36058 (N_36058,N_35655,N_35534);
nand U36059 (N_36059,N_35931,N_35716);
xor U36060 (N_36060,N_35777,N_35840);
and U36061 (N_36061,N_35034,N_35887);
or U36062 (N_36062,N_35372,N_35590);
xnor U36063 (N_36063,N_35851,N_35804);
nand U36064 (N_36064,N_35459,N_35426);
and U36065 (N_36065,N_35340,N_35033);
nor U36066 (N_36066,N_35194,N_35539);
nand U36067 (N_36067,N_35765,N_35595);
or U36068 (N_36068,N_35905,N_35216);
xnor U36069 (N_36069,N_35866,N_35225);
xnor U36070 (N_36070,N_35338,N_35066);
nand U36071 (N_36071,N_35308,N_35435);
nand U36072 (N_36072,N_35618,N_35687);
or U36073 (N_36073,N_35369,N_35412);
and U36074 (N_36074,N_35404,N_35383);
nand U36075 (N_36075,N_35537,N_35466);
nor U36076 (N_36076,N_35461,N_35419);
and U36077 (N_36077,N_35008,N_35886);
xnor U36078 (N_36078,N_35666,N_35797);
or U36079 (N_36079,N_35794,N_35320);
or U36080 (N_36080,N_35231,N_35006);
and U36081 (N_36081,N_35600,N_35542);
and U36082 (N_36082,N_35913,N_35718);
xor U36083 (N_36083,N_35891,N_35304);
and U36084 (N_36084,N_35376,N_35909);
xor U36085 (N_36085,N_35069,N_35012);
xor U36086 (N_36086,N_35915,N_35493);
and U36087 (N_36087,N_35364,N_35224);
and U36088 (N_36088,N_35662,N_35040);
nor U36089 (N_36089,N_35227,N_35188);
or U36090 (N_36090,N_35524,N_35086);
nor U36091 (N_36091,N_35686,N_35047);
nor U36092 (N_36092,N_35776,N_35892);
nand U36093 (N_36093,N_35174,N_35609);
nand U36094 (N_36094,N_35924,N_35995);
nor U36095 (N_36095,N_35564,N_35603);
xnor U36096 (N_36096,N_35469,N_35583);
or U36097 (N_36097,N_35487,N_35315);
xnor U36098 (N_36098,N_35807,N_35943);
nor U36099 (N_36099,N_35212,N_35207);
xnor U36100 (N_36100,N_35795,N_35019);
xor U36101 (N_36101,N_35353,N_35030);
and U36102 (N_36102,N_35855,N_35183);
nand U36103 (N_36103,N_35763,N_35095);
xor U36104 (N_36104,N_35783,N_35623);
and U36105 (N_36105,N_35685,N_35171);
nor U36106 (N_36106,N_35463,N_35325);
nand U36107 (N_36107,N_35262,N_35249);
and U36108 (N_36108,N_35912,N_35156);
and U36109 (N_36109,N_35947,N_35848);
nand U36110 (N_36110,N_35032,N_35789);
nand U36111 (N_36111,N_35114,N_35983);
xnor U36112 (N_36112,N_35167,N_35723);
nor U36113 (N_36113,N_35332,N_35525);
and U36114 (N_36114,N_35373,N_35043);
nand U36115 (N_36115,N_35417,N_35579);
xor U36116 (N_36116,N_35184,N_35334);
xor U36117 (N_36117,N_35626,N_35172);
and U36118 (N_36118,N_35645,N_35170);
nand U36119 (N_36119,N_35281,N_35403);
nor U36120 (N_36120,N_35305,N_35504);
or U36121 (N_36121,N_35189,N_35904);
nand U36122 (N_36122,N_35000,N_35620);
or U36123 (N_36123,N_35864,N_35660);
nand U36124 (N_36124,N_35496,N_35665);
xor U36125 (N_36125,N_35402,N_35240);
and U36126 (N_36126,N_35722,N_35782);
xor U36127 (N_36127,N_35077,N_35215);
xor U36128 (N_36128,N_35884,N_35276);
xor U36129 (N_36129,N_35269,N_35852);
and U36130 (N_36130,N_35144,N_35969);
and U36131 (N_36131,N_35621,N_35523);
or U36132 (N_36132,N_35800,N_35318);
nand U36133 (N_36133,N_35869,N_35298);
nand U36134 (N_36134,N_35672,N_35431);
or U36135 (N_36135,N_35732,N_35393);
nor U36136 (N_36136,N_35336,N_35549);
nor U36137 (N_36137,N_35597,N_35773);
nand U36138 (N_36138,N_35880,N_35878);
nor U36139 (N_36139,N_35053,N_35885);
nand U36140 (N_36140,N_35477,N_35029);
nand U36141 (N_36141,N_35637,N_35124);
nand U36142 (N_36142,N_35175,N_35071);
and U36143 (N_36143,N_35930,N_35903);
or U36144 (N_36144,N_35096,N_35482);
nor U36145 (N_36145,N_35185,N_35853);
xnor U36146 (N_36146,N_35250,N_35313);
or U36147 (N_36147,N_35064,N_35163);
or U36148 (N_36148,N_35195,N_35584);
or U36149 (N_36149,N_35200,N_35631);
xor U36150 (N_36150,N_35920,N_35292);
xnor U36151 (N_36151,N_35165,N_35715);
and U36152 (N_36152,N_35505,N_35953);
and U36153 (N_36153,N_35288,N_35133);
nor U36154 (N_36154,N_35703,N_35490);
nor U36155 (N_36155,N_35519,N_35678);
or U36156 (N_36156,N_35747,N_35870);
and U36157 (N_36157,N_35182,N_35612);
or U36158 (N_36158,N_35245,N_35293);
or U36159 (N_36159,N_35598,N_35873);
and U36160 (N_36160,N_35247,N_35605);
and U36161 (N_36161,N_35100,N_35385);
nand U36162 (N_36162,N_35624,N_35607);
or U36163 (N_36163,N_35384,N_35129);
nand U36164 (N_36164,N_35974,N_35901);
or U36165 (N_36165,N_35606,N_35742);
and U36166 (N_36166,N_35630,N_35625);
nand U36167 (N_36167,N_35186,N_35881);
and U36168 (N_36168,N_35669,N_35919);
xor U36169 (N_36169,N_35398,N_35745);
xor U36170 (N_36170,N_35682,N_35841);
nand U36171 (N_36171,N_35042,N_35571);
nand U36172 (N_36172,N_35652,N_35354);
nand U36173 (N_36173,N_35120,N_35641);
and U36174 (N_36174,N_35287,N_35146);
nand U36175 (N_36175,N_35285,N_35444);
or U36176 (N_36176,N_35158,N_35513);
xor U36177 (N_36177,N_35816,N_35897);
and U36178 (N_36178,N_35286,N_35344);
and U36179 (N_36179,N_35730,N_35358);
xnor U36180 (N_36180,N_35244,N_35152);
xnor U36181 (N_36181,N_35123,N_35312);
nor U36182 (N_36182,N_35255,N_35142);
or U36183 (N_36183,N_35007,N_35492);
nand U36184 (N_36184,N_35858,N_35646);
and U36185 (N_36185,N_35567,N_35990);
or U36186 (N_36186,N_35137,N_35028);
xor U36187 (N_36187,N_35767,N_35076);
nor U36188 (N_36188,N_35604,N_35592);
and U36189 (N_36189,N_35535,N_35411);
and U36190 (N_36190,N_35918,N_35746);
and U36191 (N_36191,N_35991,N_35706);
xnor U36192 (N_36192,N_35988,N_35406);
or U36193 (N_36193,N_35798,N_35688);
and U36194 (N_36194,N_35976,N_35963);
and U36195 (N_36195,N_35486,N_35649);
nor U36196 (N_36196,N_35051,N_35021);
nand U36197 (N_36197,N_35611,N_35485);
nand U36198 (N_36198,N_35517,N_35154);
and U36199 (N_36199,N_35708,N_35675);
and U36200 (N_36200,N_35779,N_35488);
nor U36201 (N_36201,N_35284,N_35448);
or U36202 (N_36202,N_35945,N_35608);
xor U36203 (N_36203,N_35453,N_35483);
or U36204 (N_36204,N_35929,N_35236);
xor U36205 (N_36205,N_35994,N_35845);
nand U36206 (N_36206,N_35617,N_35361);
and U36207 (N_36207,N_35951,N_35140);
nor U36208 (N_36208,N_35379,N_35465);
nand U36209 (N_36209,N_35668,N_35814);
nor U36210 (N_36210,N_35895,N_35982);
and U36211 (N_36211,N_35503,N_35695);
or U36212 (N_36212,N_35531,N_35145);
xnor U36213 (N_36213,N_35468,N_35074);
or U36214 (N_36214,N_35882,N_35515);
or U36215 (N_36215,N_35001,N_35407);
nand U36216 (N_36216,N_35826,N_35998);
and U36217 (N_36217,N_35989,N_35999);
nand U36218 (N_36218,N_35507,N_35049);
xnor U36219 (N_36219,N_35326,N_35356);
and U36220 (N_36220,N_35633,N_35894);
nor U36221 (N_36221,N_35162,N_35967);
nor U36222 (N_36222,N_35940,N_35401);
nor U36223 (N_36223,N_35993,N_35973);
nand U36224 (N_36224,N_35923,N_35965);
and U36225 (N_36225,N_35299,N_35719);
or U36226 (N_36226,N_35740,N_35785);
or U36227 (N_36227,N_35161,N_35057);
nand U36228 (N_36228,N_35437,N_35696);
nand U36229 (N_36229,N_35806,N_35191);
xnor U36230 (N_36230,N_35199,N_35013);
nor U36231 (N_36231,N_35911,N_35387);
and U36232 (N_36232,N_35808,N_35454);
or U36233 (N_36233,N_35449,N_35643);
and U36234 (N_36234,N_35472,N_35689);
or U36235 (N_36235,N_35445,N_35822);
xor U36236 (N_36236,N_35786,N_35022);
nor U36237 (N_36237,N_35075,N_35128);
xnor U36238 (N_36238,N_35093,N_35470);
or U36239 (N_36239,N_35824,N_35041);
and U36240 (N_36240,N_35112,N_35300);
nand U36241 (N_36241,N_35346,N_35935);
xor U36242 (N_36242,N_35311,N_35629);
nor U36243 (N_36243,N_35585,N_35538);
or U36244 (N_36244,N_35169,N_35101);
nor U36245 (N_36245,N_35260,N_35208);
or U36246 (N_36246,N_35817,N_35068);
or U36247 (N_36247,N_35450,N_35342);
nor U36248 (N_36248,N_35751,N_35052);
or U36249 (N_36249,N_35272,N_35038);
nor U36250 (N_36250,N_35638,N_35160);
and U36251 (N_36251,N_35506,N_35065);
xnor U36252 (N_36252,N_35017,N_35424);
xnor U36253 (N_36253,N_35654,N_35770);
and U36254 (N_36254,N_35950,N_35831);
or U36255 (N_36255,N_35414,N_35545);
nor U36256 (N_36256,N_35981,N_35975);
xor U36257 (N_36257,N_35838,N_35516);
xnor U36258 (N_36258,N_35290,N_35087);
nor U36259 (N_36259,N_35543,N_35164);
nor U36260 (N_36260,N_35784,N_35861);
nor U36261 (N_36261,N_35615,N_35602);
nand U36262 (N_36262,N_35319,N_35769);
nand U36263 (N_36263,N_35509,N_35229);
xor U36264 (N_36264,N_35367,N_35771);
or U36265 (N_36265,N_35510,N_35736);
or U36266 (N_36266,N_35705,N_35011);
or U36267 (N_36267,N_35239,N_35737);
nand U36268 (N_36268,N_35889,N_35127);
xor U36269 (N_36269,N_35203,N_35568);
or U36270 (N_36270,N_35875,N_35081);
xnor U36271 (N_36271,N_35177,N_35508);
and U36272 (N_36272,N_35978,N_35520);
and U36273 (N_36273,N_35117,N_35839);
nor U36274 (N_36274,N_35078,N_35653);
nor U36275 (N_36275,N_35992,N_35781);
and U36276 (N_36276,N_35263,N_35540);
and U36277 (N_36277,N_35827,N_35958);
and U36278 (N_36278,N_35024,N_35295);
and U36279 (N_36279,N_35178,N_35233);
or U36280 (N_36280,N_35828,N_35268);
nand U36281 (N_36281,N_35720,N_35147);
or U36282 (N_36282,N_35594,N_35415);
nor U36283 (N_36283,N_35759,N_35382);
nand U36284 (N_36284,N_35408,N_35283);
and U36285 (N_36285,N_35352,N_35790);
nand U36286 (N_36286,N_35634,N_35157);
and U36287 (N_36287,N_35265,N_35390);
xor U36288 (N_36288,N_35209,N_35232);
nand U36289 (N_36289,N_35335,N_35323);
nor U36290 (N_36290,N_35547,N_35099);
nand U36291 (N_36291,N_35091,N_35176);
nand U36292 (N_36292,N_35614,N_35753);
and U36293 (N_36293,N_35589,N_35009);
nor U36294 (N_36294,N_35026,N_35136);
or U36295 (N_36295,N_35721,N_35310);
nand U36296 (N_36296,N_35324,N_35259);
nor U36297 (N_36297,N_35835,N_35351);
nand U36298 (N_36298,N_35690,N_35528);
or U36299 (N_36299,N_35577,N_35728);
and U36300 (N_36300,N_35910,N_35908);
nand U36301 (N_36301,N_35471,N_35704);
and U36302 (N_36302,N_35859,N_35899);
or U36303 (N_36303,N_35581,N_35570);
nand U36304 (N_36304,N_35141,N_35613);
nor U36305 (N_36305,N_35569,N_35251);
xnor U36306 (N_36306,N_35102,N_35258);
or U36307 (N_36307,N_35109,N_35854);
xnor U36308 (N_36308,N_35070,N_35921);
nor U36309 (N_36309,N_35670,N_35374);
nand U36310 (N_36310,N_35683,N_35180);
nand U36311 (N_36311,N_35956,N_35386);
xnor U36312 (N_36312,N_35877,N_35578);
nand U36313 (N_36313,N_35436,N_35580);
and U36314 (N_36314,N_35409,N_35206);
and U36315 (N_36315,N_35927,N_35405);
nand U36316 (N_36316,N_35378,N_35111);
and U36317 (N_36317,N_35481,N_35296);
and U36318 (N_36318,N_35055,N_35278);
nand U36319 (N_36319,N_35309,N_35457);
and U36320 (N_36320,N_35731,N_35327);
and U36321 (N_36321,N_35933,N_35396);
or U36322 (N_36322,N_35512,N_35561);
and U36323 (N_36323,N_35443,N_35226);
xor U36324 (N_36324,N_35241,N_35371);
or U36325 (N_36325,N_35832,N_35741);
or U36326 (N_36326,N_35153,N_35698);
and U36327 (N_36327,N_35764,N_35261);
nand U36328 (N_36328,N_35347,N_35223);
nand U36329 (N_36329,N_35230,N_35467);
or U36330 (N_36330,N_35416,N_35823);
or U36331 (N_36331,N_35627,N_35394);
and U36332 (N_36332,N_35526,N_35341);
and U36333 (N_36333,N_35192,N_35291);
and U36334 (N_36334,N_35711,N_35132);
or U36335 (N_36335,N_35035,N_35389);
or U36336 (N_36336,N_35809,N_35896);
xnor U36337 (N_36337,N_35707,N_35220);
nand U36338 (N_36338,N_35893,N_35159);
nor U36339 (N_36339,N_35328,N_35616);
nor U36340 (N_36340,N_35959,N_35428);
nand U36341 (N_36341,N_35970,N_35438);
xnor U36342 (N_36342,N_35636,N_35761);
xor U36343 (N_36343,N_35270,N_35455);
nor U36344 (N_36344,N_35130,N_35610);
nor U36345 (N_36345,N_35555,N_35805);
and U36346 (N_36346,N_35502,N_35684);
xor U36347 (N_36347,N_35619,N_35103);
nand U36348 (N_36348,N_35368,N_35733);
nand U36349 (N_36349,N_35254,N_35898);
or U36350 (N_36350,N_35775,N_35713);
and U36351 (N_36351,N_35277,N_35768);
xnor U36352 (N_36352,N_35556,N_35559);
nor U36353 (N_36353,N_35214,N_35204);
xor U36354 (N_36354,N_35527,N_35301);
nor U36355 (N_36355,N_35085,N_35273);
nand U36356 (N_36356,N_35766,N_35242);
xnor U36357 (N_36357,N_35890,N_35717);
nand U36358 (N_36358,N_35801,N_35714);
nand U36359 (N_36359,N_35362,N_35536);
and U36360 (N_36360,N_35433,N_35464);
nor U36361 (N_36361,N_35056,N_35925);
or U36362 (N_36362,N_35045,N_35810);
or U36363 (N_36363,N_35957,N_35879);
nand U36364 (N_36364,N_35932,N_35149);
and U36365 (N_36365,N_35181,N_35661);
nor U36366 (N_36366,N_35566,N_35441);
or U36367 (N_36367,N_35725,N_35803);
nand U36368 (N_36368,N_35829,N_35760);
nand U36369 (N_36369,N_35647,N_35811);
nand U36370 (N_36370,N_35048,N_35985);
or U36371 (N_36371,N_35758,N_35274);
nor U36372 (N_36372,N_35681,N_35027);
nor U36373 (N_36373,N_35306,N_35710);
nand U36374 (N_36374,N_35484,N_35002);
xnor U36375 (N_36375,N_35980,N_35090);
xnor U36376 (N_36376,N_35122,N_35622);
xor U36377 (N_36377,N_35252,N_35856);
or U36378 (N_36378,N_35440,N_35774);
and U36379 (N_36379,N_35849,N_35872);
nor U36380 (N_36380,N_35888,N_35360);
or U36381 (N_36381,N_35987,N_35533);
nand U36382 (N_36382,N_35694,N_35587);
and U36383 (N_36383,N_35421,N_35031);
or U36384 (N_36384,N_35514,N_35413);
nand U36385 (N_36385,N_35756,N_35997);
nor U36386 (N_36386,N_35452,N_35348);
or U36387 (N_36387,N_35321,N_35037);
nor U36388 (N_36388,N_35370,N_35480);
nor U36389 (N_36389,N_35780,N_35271);
or U36390 (N_36390,N_35359,N_35546);
or U36391 (N_36391,N_35005,N_35067);
or U36392 (N_36392,N_35939,N_35656);
and U36393 (N_36393,N_35850,N_35871);
xnor U36394 (N_36394,N_35757,N_35228);
and U36395 (N_36395,N_35727,N_35726);
nor U36396 (N_36396,N_35724,N_35530);
nor U36397 (N_36397,N_35139,N_35121);
nor U36398 (N_36398,N_35550,N_35400);
xnor U36399 (N_36399,N_35529,N_35105);
nand U36400 (N_36400,N_35198,N_35084);
xor U36401 (N_36401,N_35489,N_35642);
or U36402 (N_36402,N_35792,N_35560);
xnor U36403 (N_36403,N_35842,N_35392);
xor U36404 (N_36404,N_35586,N_35098);
xor U36405 (N_36405,N_35316,N_35237);
xnor U36406 (N_36406,N_35125,N_35080);
nor U36407 (N_36407,N_35218,N_35427);
xor U36408 (N_36408,N_35574,N_35857);
or U36409 (N_36409,N_35439,N_35635);
and U36410 (N_36410,N_35825,N_35110);
xnor U36411 (N_36411,N_35089,N_35748);
nor U36412 (N_36412,N_35735,N_35072);
or U36413 (N_36413,N_35494,N_35796);
nor U36414 (N_36414,N_35984,N_35676);
nor U36415 (N_36415,N_35442,N_35349);
xnor U36416 (N_36416,N_35106,N_35691);
xnor U36417 (N_36417,N_35926,N_35977);
and U36418 (N_36418,N_35391,N_35632);
or U36419 (N_36419,N_35575,N_35812);
nor U36420 (N_36420,N_35418,N_35234);
xor U36421 (N_36421,N_35476,N_35423);
and U36422 (N_36422,N_35788,N_35833);
nand U36423 (N_36423,N_35151,N_35475);
nand U36424 (N_36424,N_35755,N_35802);
and U36425 (N_36425,N_35734,N_35119);
xor U36426 (N_36426,N_35020,N_35644);
xor U36427 (N_36427,N_35772,N_35501);
and U36428 (N_36428,N_35673,N_35447);
xnor U36429 (N_36429,N_35155,N_35964);
and U36430 (N_36430,N_35874,N_35548);
xor U36431 (N_36431,N_35173,N_35246);
or U36432 (N_36432,N_35743,N_35916);
nand U36433 (N_36433,N_35572,N_35092);
xnor U36434 (N_36434,N_35553,N_35837);
nor U36435 (N_36435,N_35063,N_35565);
or U36436 (N_36436,N_35003,N_35113);
or U36437 (N_36437,N_35815,N_35115);
or U36438 (N_36438,N_35432,N_35303);
xor U36439 (N_36439,N_35253,N_35563);
nand U36440 (N_36440,N_35267,N_35314);
nor U36441 (N_36441,N_35744,N_35640);
and U36442 (N_36442,N_35960,N_35702);
or U36443 (N_36443,N_35813,N_35948);
nand U36444 (N_36444,N_35104,N_35395);
nand U36445 (N_36445,N_35700,N_35497);
nand U36446 (N_36446,N_35712,N_35762);
or U36447 (N_36447,N_35588,N_35972);
xnor U36448 (N_36448,N_35430,N_35996);
or U36449 (N_36449,N_35738,N_35010);
or U36450 (N_36450,N_35599,N_35778);
nand U36451 (N_36451,N_35739,N_35211);
nand U36452 (N_36452,N_35752,N_35282);
nand U36453 (N_36453,N_35264,N_35297);
nand U36454 (N_36454,N_35322,N_35582);
or U36455 (N_36455,N_35434,N_35425);
and U36456 (N_36456,N_35862,N_35680);
xor U36457 (N_36457,N_35116,N_35243);
and U36458 (N_36458,N_35558,N_35952);
and U36459 (N_36459,N_35949,N_35552);
nor U36460 (N_36460,N_35143,N_35302);
or U36461 (N_36461,N_35219,N_35138);
or U36462 (N_36462,N_35365,N_35397);
nor U36463 (N_36463,N_35339,N_35573);
nor U36464 (N_36464,N_35860,N_35971);
nor U36465 (N_36465,N_35061,N_35059);
nor U36466 (N_36466,N_35331,N_35601);
xnor U36467 (N_36467,N_35337,N_35046);
or U36468 (N_36468,N_35938,N_35451);
xnor U36469 (N_36469,N_35193,N_35830);
nor U36470 (N_36470,N_35663,N_35196);
and U36471 (N_36471,N_35015,N_35914);
nor U36472 (N_36472,N_35388,N_35054);
nor U36473 (N_36473,N_35591,N_35474);
or U36474 (N_36474,N_35750,N_35062);
or U36475 (N_36475,N_35968,N_35399);
or U36476 (N_36476,N_35082,N_35679);
and U36477 (N_36477,N_35060,N_35699);
nor U36478 (N_36478,N_35317,N_35664);
or U36479 (N_36479,N_35222,N_35867);
nor U36480 (N_36480,N_35648,N_35639);
or U36481 (N_36481,N_35697,N_35865);
xor U36482 (N_36482,N_35329,N_35671);
and U36483 (N_36483,N_35554,N_35275);
nand U36484 (N_36484,N_35749,N_35366);
and U36485 (N_36485,N_35955,N_35754);
and U36486 (N_36486,N_35079,N_35667);
nand U36487 (N_36487,N_35039,N_35473);
and U36488 (N_36488,N_35422,N_35819);
or U36489 (N_36489,N_35187,N_35941);
and U36490 (N_36490,N_35847,N_35179);
nor U36491 (N_36491,N_35692,N_35343);
and U36492 (N_36492,N_35023,N_35355);
or U36493 (N_36493,N_35729,N_35307);
nand U36494 (N_36494,N_35016,N_35150);
and U36495 (N_36495,N_35134,N_35596);
nor U36496 (N_36496,N_35256,N_35460);
or U36497 (N_36497,N_35350,N_35962);
and U36498 (N_36498,N_35166,N_35799);
or U36499 (N_36499,N_35456,N_35210);
nand U36500 (N_36500,N_35708,N_35504);
nor U36501 (N_36501,N_35346,N_35601);
xor U36502 (N_36502,N_35787,N_35448);
xnor U36503 (N_36503,N_35989,N_35880);
and U36504 (N_36504,N_35312,N_35440);
and U36505 (N_36505,N_35130,N_35431);
and U36506 (N_36506,N_35183,N_35804);
and U36507 (N_36507,N_35502,N_35005);
or U36508 (N_36508,N_35649,N_35915);
or U36509 (N_36509,N_35102,N_35414);
or U36510 (N_36510,N_35504,N_35236);
nor U36511 (N_36511,N_35359,N_35606);
nor U36512 (N_36512,N_35135,N_35823);
nand U36513 (N_36513,N_35021,N_35943);
xnor U36514 (N_36514,N_35796,N_35018);
nand U36515 (N_36515,N_35940,N_35106);
xor U36516 (N_36516,N_35511,N_35962);
and U36517 (N_36517,N_35621,N_35690);
xor U36518 (N_36518,N_35257,N_35554);
nand U36519 (N_36519,N_35267,N_35302);
nand U36520 (N_36520,N_35017,N_35405);
or U36521 (N_36521,N_35241,N_35221);
xor U36522 (N_36522,N_35874,N_35135);
or U36523 (N_36523,N_35270,N_35132);
xnor U36524 (N_36524,N_35185,N_35351);
xor U36525 (N_36525,N_35028,N_35454);
nor U36526 (N_36526,N_35173,N_35528);
and U36527 (N_36527,N_35837,N_35735);
nand U36528 (N_36528,N_35690,N_35424);
xor U36529 (N_36529,N_35167,N_35768);
and U36530 (N_36530,N_35219,N_35865);
nand U36531 (N_36531,N_35616,N_35950);
xnor U36532 (N_36532,N_35504,N_35368);
nand U36533 (N_36533,N_35204,N_35803);
nand U36534 (N_36534,N_35315,N_35939);
nand U36535 (N_36535,N_35677,N_35951);
xnor U36536 (N_36536,N_35912,N_35135);
and U36537 (N_36537,N_35890,N_35251);
and U36538 (N_36538,N_35270,N_35139);
nor U36539 (N_36539,N_35558,N_35028);
xnor U36540 (N_36540,N_35559,N_35141);
and U36541 (N_36541,N_35059,N_35722);
xnor U36542 (N_36542,N_35657,N_35793);
nor U36543 (N_36543,N_35960,N_35802);
and U36544 (N_36544,N_35362,N_35951);
nor U36545 (N_36545,N_35430,N_35920);
and U36546 (N_36546,N_35051,N_35619);
xor U36547 (N_36547,N_35121,N_35420);
or U36548 (N_36548,N_35129,N_35027);
or U36549 (N_36549,N_35204,N_35656);
nor U36550 (N_36550,N_35487,N_35601);
and U36551 (N_36551,N_35686,N_35582);
and U36552 (N_36552,N_35494,N_35704);
nor U36553 (N_36553,N_35251,N_35365);
or U36554 (N_36554,N_35871,N_35114);
or U36555 (N_36555,N_35691,N_35822);
or U36556 (N_36556,N_35847,N_35612);
nand U36557 (N_36557,N_35543,N_35306);
xor U36558 (N_36558,N_35813,N_35186);
xor U36559 (N_36559,N_35899,N_35560);
nand U36560 (N_36560,N_35046,N_35299);
and U36561 (N_36561,N_35028,N_35603);
nor U36562 (N_36562,N_35964,N_35760);
xor U36563 (N_36563,N_35362,N_35384);
xor U36564 (N_36564,N_35745,N_35769);
nand U36565 (N_36565,N_35109,N_35227);
and U36566 (N_36566,N_35392,N_35017);
and U36567 (N_36567,N_35183,N_35321);
nand U36568 (N_36568,N_35675,N_35000);
nor U36569 (N_36569,N_35680,N_35432);
nand U36570 (N_36570,N_35770,N_35543);
xnor U36571 (N_36571,N_35554,N_35083);
and U36572 (N_36572,N_35558,N_35405);
nand U36573 (N_36573,N_35833,N_35118);
xnor U36574 (N_36574,N_35548,N_35258);
nand U36575 (N_36575,N_35972,N_35130);
nand U36576 (N_36576,N_35737,N_35790);
nor U36577 (N_36577,N_35774,N_35409);
xor U36578 (N_36578,N_35115,N_35170);
xnor U36579 (N_36579,N_35288,N_35941);
nor U36580 (N_36580,N_35689,N_35611);
and U36581 (N_36581,N_35359,N_35346);
nand U36582 (N_36582,N_35324,N_35018);
nand U36583 (N_36583,N_35795,N_35249);
and U36584 (N_36584,N_35302,N_35793);
and U36585 (N_36585,N_35528,N_35462);
xnor U36586 (N_36586,N_35356,N_35405);
nand U36587 (N_36587,N_35040,N_35908);
and U36588 (N_36588,N_35112,N_35684);
and U36589 (N_36589,N_35416,N_35991);
nor U36590 (N_36590,N_35457,N_35875);
or U36591 (N_36591,N_35621,N_35965);
and U36592 (N_36592,N_35298,N_35390);
and U36593 (N_36593,N_35200,N_35120);
nand U36594 (N_36594,N_35678,N_35019);
nor U36595 (N_36595,N_35907,N_35888);
nand U36596 (N_36596,N_35240,N_35399);
and U36597 (N_36597,N_35858,N_35640);
nor U36598 (N_36598,N_35586,N_35770);
and U36599 (N_36599,N_35442,N_35949);
and U36600 (N_36600,N_35385,N_35138);
and U36601 (N_36601,N_35682,N_35137);
xnor U36602 (N_36602,N_35301,N_35948);
xor U36603 (N_36603,N_35546,N_35411);
xor U36604 (N_36604,N_35772,N_35466);
nand U36605 (N_36605,N_35813,N_35967);
and U36606 (N_36606,N_35803,N_35087);
nand U36607 (N_36607,N_35895,N_35093);
or U36608 (N_36608,N_35108,N_35430);
nand U36609 (N_36609,N_35291,N_35293);
or U36610 (N_36610,N_35274,N_35946);
nor U36611 (N_36611,N_35829,N_35297);
nand U36612 (N_36612,N_35896,N_35283);
nor U36613 (N_36613,N_35081,N_35609);
or U36614 (N_36614,N_35665,N_35117);
nand U36615 (N_36615,N_35364,N_35089);
nor U36616 (N_36616,N_35889,N_35606);
and U36617 (N_36617,N_35235,N_35201);
and U36618 (N_36618,N_35323,N_35066);
nand U36619 (N_36619,N_35294,N_35037);
nand U36620 (N_36620,N_35863,N_35130);
and U36621 (N_36621,N_35276,N_35745);
xnor U36622 (N_36622,N_35465,N_35229);
nor U36623 (N_36623,N_35317,N_35160);
nand U36624 (N_36624,N_35283,N_35529);
xnor U36625 (N_36625,N_35249,N_35350);
and U36626 (N_36626,N_35737,N_35103);
and U36627 (N_36627,N_35143,N_35486);
xor U36628 (N_36628,N_35024,N_35553);
nor U36629 (N_36629,N_35560,N_35172);
nor U36630 (N_36630,N_35993,N_35897);
or U36631 (N_36631,N_35070,N_35040);
and U36632 (N_36632,N_35946,N_35679);
and U36633 (N_36633,N_35990,N_35384);
nand U36634 (N_36634,N_35760,N_35379);
xor U36635 (N_36635,N_35700,N_35432);
or U36636 (N_36636,N_35272,N_35947);
or U36637 (N_36637,N_35343,N_35151);
or U36638 (N_36638,N_35361,N_35770);
nor U36639 (N_36639,N_35643,N_35028);
or U36640 (N_36640,N_35615,N_35445);
or U36641 (N_36641,N_35079,N_35335);
or U36642 (N_36642,N_35208,N_35705);
and U36643 (N_36643,N_35207,N_35440);
xnor U36644 (N_36644,N_35365,N_35031);
nor U36645 (N_36645,N_35735,N_35071);
or U36646 (N_36646,N_35517,N_35560);
or U36647 (N_36647,N_35966,N_35508);
and U36648 (N_36648,N_35805,N_35542);
or U36649 (N_36649,N_35116,N_35712);
xnor U36650 (N_36650,N_35258,N_35733);
or U36651 (N_36651,N_35285,N_35738);
xor U36652 (N_36652,N_35965,N_35763);
and U36653 (N_36653,N_35508,N_35118);
and U36654 (N_36654,N_35966,N_35366);
and U36655 (N_36655,N_35655,N_35484);
or U36656 (N_36656,N_35421,N_35499);
or U36657 (N_36657,N_35769,N_35885);
nand U36658 (N_36658,N_35631,N_35206);
nand U36659 (N_36659,N_35080,N_35538);
or U36660 (N_36660,N_35918,N_35825);
or U36661 (N_36661,N_35149,N_35832);
nor U36662 (N_36662,N_35682,N_35360);
nand U36663 (N_36663,N_35880,N_35867);
nor U36664 (N_36664,N_35652,N_35294);
nand U36665 (N_36665,N_35573,N_35274);
and U36666 (N_36666,N_35902,N_35538);
nor U36667 (N_36667,N_35232,N_35862);
xor U36668 (N_36668,N_35611,N_35169);
nand U36669 (N_36669,N_35433,N_35543);
xnor U36670 (N_36670,N_35633,N_35477);
nor U36671 (N_36671,N_35691,N_35050);
nand U36672 (N_36672,N_35298,N_35182);
nand U36673 (N_36673,N_35668,N_35683);
nor U36674 (N_36674,N_35815,N_35795);
nor U36675 (N_36675,N_35400,N_35779);
nor U36676 (N_36676,N_35251,N_35685);
nand U36677 (N_36677,N_35958,N_35919);
nand U36678 (N_36678,N_35095,N_35313);
nand U36679 (N_36679,N_35789,N_35004);
nor U36680 (N_36680,N_35453,N_35946);
nand U36681 (N_36681,N_35598,N_35642);
and U36682 (N_36682,N_35179,N_35477);
or U36683 (N_36683,N_35414,N_35877);
nand U36684 (N_36684,N_35420,N_35640);
or U36685 (N_36685,N_35952,N_35738);
or U36686 (N_36686,N_35190,N_35477);
and U36687 (N_36687,N_35393,N_35339);
nor U36688 (N_36688,N_35596,N_35793);
nand U36689 (N_36689,N_35528,N_35505);
or U36690 (N_36690,N_35592,N_35224);
xnor U36691 (N_36691,N_35138,N_35046);
nand U36692 (N_36692,N_35832,N_35432);
and U36693 (N_36693,N_35952,N_35651);
nand U36694 (N_36694,N_35174,N_35784);
xor U36695 (N_36695,N_35656,N_35976);
nand U36696 (N_36696,N_35831,N_35307);
xnor U36697 (N_36697,N_35368,N_35419);
xor U36698 (N_36698,N_35298,N_35302);
or U36699 (N_36699,N_35967,N_35748);
or U36700 (N_36700,N_35815,N_35354);
nand U36701 (N_36701,N_35216,N_35249);
or U36702 (N_36702,N_35988,N_35574);
and U36703 (N_36703,N_35577,N_35799);
or U36704 (N_36704,N_35198,N_35097);
xnor U36705 (N_36705,N_35803,N_35007);
and U36706 (N_36706,N_35965,N_35183);
xor U36707 (N_36707,N_35559,N_35349);
xor U36708 (N_36708,N_35239,N_35570);
nand U36709 (N_36709,N_35132,N_35329);
and U36710 (N_36710,N_35868,N_35911);
and U36711 (N_36711,N_35167,N_35092);
or U36712 (N_36712,N_35320,N_35648);
xor U36713 (N_36713,N_35801,N_35963);
xnor U36714 (N_36714,N_35001,N_35157);
and U36715 (N_36715,N_35805,N_35842);
nor U36716 (N_36716,N_35880,N_35700);
nor U36717 (N_36717,N_35472,N_35688);
or U36718 (N_36718,N_35201,N_35131);
and U36719 (N_36719,N_35395,N_35815);
and U36720 (N_36720,N_35701,N_35918);
nor U36721 (N_36721,N_35026,N_35745);
nand U36722 (N_36722,N_35438,N_35426);
and U36723 (N_36723,N_35840,N_35366);
and U36724 (N_36724,N_35711,N_35627);
and U36725 (N_36725,N_35590,N_35808);
and U36726 (N_36726,N_35924,N_35096);
and U36727 (N_36727,N_35958,N_35677);
and U36728 (N_36728,N_35215,N_35719);
and U36729 (N_36729,N_35595,N_35168);
and U36730 (N_36730,N_35118,N_35253);
nand U36731 (N_36731,N_35757,N_35231);
nand U36732 (N_36732,N_35763,N_35253);
or U36733 (N_36733,N_35279,N_35086);
and U36734 (N_36734,N_35056,N_35618);
and U36735 (N_36735,N_35152,N_35064);
nor U36736 (N_36736,N_35309,N_35323);
and U36737 (N_36737,N_35113,N_35440);
or U36738 (N_36738,N_35239,N_35449);
nor U36739 (N_36739,N_35623,N_35753);
nor U36740 (N_36740,N_35639,N_35844);
nand U36741 (N_36741,N_35988,N_35299);
nor U36742 (N_36742,N_35861,N_35115);
xnor U36743 (N_36743,N_35167,N_35570);
or U36744 (N_36744,N_35861,N_35127);
and U36745 (N_36745,N_35201,N_35327);
and U36746 (N_36746,N_35800,N_35098);
or U36747 (N_36747,N_35388,N_35619);
and U36748 (N_36748,N_35920,N_35170);
nor U36749 (N_36749,N_35083,N_35747);
nand U36750 (N_36750,N_35799,N_35107);
xor U36751 (N_36751,N_35644,N_35846);
or U36752 (N_36752,N_35648,N_35013);
nand U36753 (N_36753,N_35597,N_35685);
or U36754 (N_36754,N_35824,N_35494);
and U36755 (N_36755,N_35262,N_35634);
and U36756 (N_36756,N_35315,N_35959);
xnor U36757 (N_36757,N_35270,N_35385);
or U36758 (N_36758,N_35751,N_35185);
nand U36759 (N_36759,N_35899,N_35499);
and U36760 (N_36760,N_35422,N_35913);
xnor U36761 (N_36761,N_35618,N_35686);
and U36762 (N_36762,N_35241,N_35350);
and U36763 (N_36763,N_35432,N_35397);
and U36764 (N_36764,N_35344,N_35370);
xnor U36765 (N_36765,N_35399,N_35121);
xor U36766 (N_36766,N_35136,N_35357);
xnor U36767 (N_36767,N_35437,N_35231);
nand U36768 (N_36768,N_35667,N_35796);
xor U36769 (N_36769,N_35770,N_35015);
nor U36770 (N_36770,N_35462,N_35786);
nand U36771 (N_36771,N_35762,N_35238);
or U36772 (N_36772,N_35909,N_35065);
nor U36773 (N_36773,N_35081,N_35668);
and U36774 (N_36774,N_35782,N_35506);
or U36775 (N_36775,N_35302,N_35075);
and U36776 (N_36776,N_35872,N_35559);
xnor U36777 (N_36777,N_35873,N_35566);
xor U36778 (N_36778,N_35005,N_35466);
or U36779 (N_36779,N_35894,N_35831);
nor U36780 (N_36780,N_35945,N_35180);
nand U36781 (N_36781,N_35284,N_35250);
xnor U36782 (N_36782,N_35132,N_35033);
or U36783 (N_36783,N_35779,N_35235);
nor U36784 (N_36784,N_35022,N_35113);
nor U36785 (N_36785,N_35502,N_35662);
or U36786 (N_36786,N_35759,N_35166);
nor U36787 (N_36787,N_35546,N_35252);
xnor U36788 (N_36788,N_35840,N_35443);
nor U36789 (N_36789,N_35405,N_35605);
nand U36790 (N_36790,N_35952,N_35927);
nand U36791 (N_36791,N_35408,N_35172);
nand U36792 (N_36792,N_35473,N_35880);
xnor U36793 (N_36793,N_35145,N_35080);
xor U36794 (N_36794,N_35301,N_35620);
nand U36795 (N_36795,N_35704,N_35891);
xor U36796 (N_36796,N_35912,N_35496);
and U36797 (N_36797,N_35526,N_35281);
or U36798 (N_36798,N_35703,N_35311);
xnor U36799 (N_36799,N_35176,N_35390);
and U36800 (N_36800,N_35469,N_35141);
nor U36801 (N_36801,N_35490,N_35693);
or U36802 (N_36802,N_35744,N_35899);
xnor U36803 (N_36803,N_35560,N_35242);
nor U36804 (N_36804,N_35609,N_35565);
nor U36805 (N_36805,N_35312,N_35588);
and U36806 (N_36806,N_35087,N_35337);
or U36807 (N_36807,N_35325,N_35497);
xor U36808 (N_36808,N_35111,N_35935);
or U36809 (N_36809,N_35774,N_35056);
and U36810 (N_36810,N_35239,N_35027);
xnor U36811 (N_36811,N_35717,N_35535);
or U36812 (N_36812,N_35168,N_35334);
or U36813 (N_36813,N_35101,N_35438);
or U36814 (N_36814,N_35179,N_35489);
or U36815 (N_36815,N_35736,N_35219);
nand U36816 (N_36816,N_35078,N_35996);
and U36817 (N_36817,N_35410,N_35639);
and U36818 (N_36818,N_35814,N_35475);
nand U36819 (N_36819,N_35885,N_35289);
or U36820 (N_36820,N_35138,N_35649);
xnor U36821 (N_36821,N_35122,N_35891);
and U36822 (N_36822,N_35469,N_35967);
nor U36823 (N_36823,N_35076,N_35807);
xor U36824 (N_36824,N_35459,N_35539);
nor U36825 (N_36825,N_35666,N_35042);
nor U36826 (N_36826,N_35571,N_35990);
or U36827 (N_36827,N_35149,N_35941);
nor U36828 (N_36828,N_35099,N_35022);
and U36829 (N_36829,N_35117,N_35654);
xor U36830 (N_36830,N_35044,N_35754);
xnor U36831 (N_36831,N_35486,N_35725);
xor U36832 (N_36832,N_35580,N_35287);
or U36833 (N_36833,N_35999,N_35833);
xnor U36834 (N_36834,N_35048,N_35297);
nor U36835 (N_36835,N_35943,N_35892);
and U36836 (N_36836,N_35256,N_35205);
or U36837 (N_36837,N_35373,N_35475);
nor U36838 (N_36838,N_35139,N_35028);
xnor U36839 (N_36839,N_35328,N_35002);
and U36840 (N_36840,N_35398,N_35696);
and U36841 (N_36841,N_35451,N_35771);
or U36842 (N_36842,N_35145,N_35519);
nand U36843 (N_36843,N_35535,N_35241);
xor U36844 (N_36844,N_35481,N_35045);
and U36845 (N_36845,N_35363,N_35182);
or U36846 (N_36846,N_35544,N_35087);
and U36847 (N_36847,N_35551,N_35619);
nor U36848 (N_36848,N_35819,N_35175);
and U36849 (N_36849,N_35281,N_35584);
nor U36850 (N_36850,N_35481,N_35848);
and U36851 (N_36851,N_35542,N_35486);
xor U36852 (N_36852,N_35171,N_35066);
nand U36853 (N_36853,N_35679,N_35865);
xor U36854 (N_36854,N_35122,N_35890);
and U36855 (N_36855,N_35713,N_35631);
and U36856 (N_36856,N_35335,N_35267);
and U36857 (N_36857,N_35540,N_35510);
and U36858 (N_36858,N_35385,N_35989);
or U36859 (N_36859,N_35514,N_35575);
and U36860 (N_36860,N_35075,N_35531);
or U36861 (N_36861,N_35559,N_35956);
or U36862 (N_36862,N_35410,N_35001);
xor U36863 (N_36863,N_35098,N_35827);
nand U36864 (N_36864,N_35409,N_35609);
and U36865 (N_36865,N_35503,N_35965);
nor U36866 (N_36866,N_35822,N_35002);
nand U36867 (N_36867,N_35251,N_35352);
xnor U36868 (N_36868,N_35973,N_35915);
nand U36869 (N_36869,N_35582,N_35981);
xor U36870 (N_36870,N_35999,N_35458);
nand U36871 (N_36871,N_35817,N_35202);
nand U36872 (N_36872,N_35968,N_35233);
xor U36873 (N_36873,N_35248,N_35643);
or U36874 (N_36874,N_35423,N_35990);
nor U36875 (N_36875,N_35188,N_35162);
xnor U36876 (N_36876,N_35234,N_35827);
nand U36877 (N_36877,N_35992,N_35919);
nand U36878 (N_36878,N_35124,N_35497);
xnor U36879 (N_36879,N_35843,N_35522);
nor U36880 (N_36880,N_35443,N_35824);
xnor U36881 (N_36881,N_35337,N_35179);
xnor U36882 (N_36882,N_35002,N_35512);
and U36883 (N_36883,N_35623,N_35403);
or U36884 (N_36884,N_35395,N_35276);
nand U36885 (N_36885,N_35987,N_35313);
nor U36886 (N_36886,N_35823,N_35112);
or U36887 (N_36887,N_35986,N_35192);
or U36888 (N_36888,N_35460,N_35794);
or U36889 (N_36889,N_35175,N_35436);
xor U36890 (N_36890,N_35812,N_35450);
or U36891 (N_36891,N_35116,N_35536);
or U36892 (N_36892,N_35722,N_35081);
and U36893 (N_36893,N_35138,N_35518);
nand U36894 (N_36894,N_35384,N_35998);
xor U36895 (N_36895,N_35619,N_35768);
and U36896 (N_36896,N_35542,N_35791);
xnor U36897 (N_36897,N_35057,N_35409);
or U36898 (N_36898,N_35448,N_35221);
nor U36899 (N_36899,N_35065,N_35157);
nand U36900 (N_36900,N_35051,N_35460);
and U36901 (N_36901,N_35283,N_35074);
xnor U36902 (N_36902,N_35219,N_35747);
nor U36903 (N_36903,N_35718,N_35846);
and U36904 (N_36904,N_35699,N_35343);
or U36905 (N_36905,N_35991,N_35031);
nor U36906 (N_36906,N_35766,N_35784);
nand U36907 (N_36907,N_35471,N_35777);
and U36908 (N_36908,N_35093,N_35012);
or U36909 (N_36909,N_35372,N_35402);
nor U36910 (N_36910,N_35469,N_35233);
nand U36911 (N_36911,N_35976,N_35198);
nand U36912 (N_36912,N_35777,N_35510);
nor U36913 (N_36913,N_35711,N_35415);
nand U36914 (N_36914,N_35858,N_35169);
nor U36915 (N_36915,N_35443,N_35122);
nand U36916 (N_36916,N_35948,N_35448);
nand U36917 (N_36917,N_35466,N_35583);
xor U36918 (N_36918,N_35839,N_35083);
nor U36919 (N_36919,N_35191,N_35837);
xnor U36920 (N_36920,N_35062,N_35887);
and U36921 (N_36921,N_35568,N_35921);
xnor U36922 (N_36922,N_35737,N_35430);
or U36923 (N_36923,N_35636,N_35644);
or U36924 (N_36924,N_35831,N_35502);
nor U36925 (N_36925,N_35752,N_35461);
and U36926 (N_36926,N_35889,N_35227);
and U36927 (N_36927,N_35043,N_35796);
xnor U36928 (N_36928,N_35338,N_35962);
xor U36929 (N_36929,N_35435,N_35914);
nor U36930 (N_36930,N_35265,N_35102);
and U36931 (N_36931,N_35910,N_35968);
and U36932 (N_36932,N_35014,N_35371);
and U36933 (N_36933,N_35485,N_35240);
or U36934 (N_36934,N_35516,N_35726);
xor U36935 (N_36935,N_35238,N_35660);
nor U36936 (N_36936,N_35900,N_35371);
and U36937 (N_36937,N_35724,N_35234);
xor U36938 (N_36938,N_35413,N_35467);
nand U36939 (N_36939,N_35832,N_35109);
xnor U36940 (N_36940,N_35309,N_35358);
and U36941 (N_36941,N_35347,N_35297);
or U36942 (N_36942,N_35897,N_35547);
xor U36943 (N_36943,N_35806,N_35016);
nor U36944 (N_36944,N_35669,N_35829);
or U36945 (N_36945,N_35271,N_35154);
nor U36946 (N_36946,N_35689,N_35127);
and U36947 (N_36947,N_35506,N_35815);
or U36948 (N_36948,N_35135,N_35676);
nand U36949 (N_36949,N_35944,N_35720);
nor U36950 (N_36950,N_35992,N_35505);
nor U36951 (N_36951,N_35095,N_35907);
or U36952 (N_36952,N_35845,N_35271);
or U36953 (N_36953,N_35382,N_35051);
or U36954 (N_36954,N_35772,N_35265);
nand U36955 (N_36955,N_35491,N_35939);
nand U36956 (N_36956,N_35100,N_35921);
nand U36957 (N_36957,N_35696,N_35351);
nor U36958 (N_36958,N_35181,N_35173);
nor U36959 (N_36959,N_35277,N_35349);
nand U36960 (N_36960,N_35919,N_35619);
xor U36961 (N_36961,N_35742,N_35228);
nor U36962 (N_36962,N_35808,N_35896);
and U36963 (N_36963,N_35451,N_35092);
xnor U36964 (N_36964,N_35404,N_35601);
or U36965 (N_36965,N_35589,N_35031);
nor U36966 (N_36966,N_35113,N_35670);
xnor U36967 (N_36967,N_35181,N_35705);
xor U36968 (N_36968,N_35837,N_35821);
xor U36969 (N_36969,N_35541,N_35136);
nor U36970 (N_36970,N_35493,N_35617);
xor U36971 (N_36971,N_35332,N_35183);
xor U36972 (N_36972,N_35104,N_35842);
nor U36973 (N_36973,N_35296,N_35525);
and U36974 (N_36974,N_35676,N_35529);
xor U36975 (N_36975,N_35558,N_35094);
xnor U36976 (N_36976,N_35604,N_35766);
and U36977 (N_36977,N_35189,N_35814);
and U36978 (N_36978,N_35216,N_35993);
nor U36979 (N_36979,N_35239,N_35325);
nand U36980 (N_36980,N_35889,N_35280);
nor U36981 (N_36981,N_35574,N_35016);
or U36982 (N_36982,N_35723,N_35449);
or U36983 (N_36983,N_35093,N_35339);
xor U36984 (N_36984,N_35234,N_35791);
nand U36985 (N_36985,N_35437,N_35655);
and U36986 (N_36986,N_35684,N_35937);
and U36987 (N_36987,N_35167,N_35357);
xnor U36988 (N_36988,N_35353,N_35186);
nor U36989 (N_36989,N_35401,N_35739);
or U36990 (N_36990,N_35940,N_35523);
and U36991 (N_36991,N_35985,N_35449);
and U36992 (N_36992,N_35010,N_35252);
and U36993 (N_36993,N_35507,N_35653);
nor U36994 (N_36994,N_35253,N_35398);
xor U36995 (N_36995,N_35243,N_35226);
or U36996 (N_36996,N_35565,N_35725);
xnor U36997 (N_36997,N_35756,N_35031);
and U36998 (N_36998,N_35433,N_35357);
and U36999 (N_36999,N_35045,N_35280);
nand U37000 (N_37000,N_36326,N_36804);
nor U37001 (N_37001,N_36750,N_36248);
or U37002 (N_37002,N_36337,N_36833);
xnor U37003 (N_37003,N_36288,N_36675);
nor U37004 (N_37004,N_36132,N_36826);
and U37005 (N_37005,N_36117,N_36224);
xnor U37006 (N_37006,N_36740,N_36836);
nand U37007 (N_37007,N_36880,N_36624);
nor U37008 (N_37008,N_36190,N_36981);
nor U37009 (N_37009,N_36491,N_36351);
or U37010 (N_37010,N_36715,N_36828);
nand U37011 (N_37011,N_36523,N_36227);
xor U37012 (N_37012,N_36061,N_36644);
nand U37013 (N_37013,N_36620,N_36287);
nand U37014 (N_37014,N_36781,N_36937);
or U37015 (N_37015,N_36294,N_36371);
nor U37016 (N_37016,N_36674,N_36877);
or U37017 (N_37017,N_36148,N_36438);
xnor U37018 (N_37018,N_36897,N_36367);
and U37019 (N_37019,N_36366,N_36342);
nand U37020 (N_37020,N_36684,N_36830);
or U37021 (N_37021,N_36748,N_36800);
and U37022 (N_37022,N_36409,N_36425);
or U37023 (N_37023,N_36908,N_36894);
and U37024 (N_37024,N_36806,N_36794);
and U37025 (N_37025,N_36980,N_36108);
and U37026 (N_37026,N_36405,N_36305);
and U37027 (N_37027,N_36576,N_36040);
nand U37028 (N_37028,N_36584,N_36668);
nand U37029 (N_37029,N_36430,N_36256);
xor U37030 (N_37030,N_36835,N_36136);
xnor U37031 (N_37031,N_36848,N_36902);
xor U37032 (N_37032,N_36499,N_36608);
nand U37033 (N_37033,N_36501,N_36166);
xnor U37034 (N_37034,N_36859,N_36537);
xor U37035 (N_37035,N_36616,N_36595);
or U37036 (N_37036,N_36555,N_36672);
or U37037 (N_37037,N_36755,N_36269);
nand U37038 (N_37038,N_36001,N_36002);
nand U37039 (N_37039,N_36494,N_36658);
nor U37040 (N_37040,N_36000,N_36015);
nand U37041 (N_37041,N_36741,N_36069);
nor U37042 (N_37042,N_36421,N_36012);
nand U37043 (N_37043,N_36358,N_36770);
or U37044 (N_37044,N_36098,N_36141);
nand U37045 (N_37045,N_36212,N_36474);
xor U37046 (N_37046,N_36298,N_36435);
xnor U37047 (N_37047,N_36129,N_36200);
xor U37048 (N_37048,N_36340,N_36670);
or U37049 (N_37049,N_36912,N_36432);
or U37050 (N_37050,N_36257,N_36119);
xnor U37051 (N_37051,N_36766,N_36946);
nor U37052 (N_37052,N_36872,N_36784);
nand U37053 (N_37053,N_36206,N_36315);
or U37054 (N_37054,N_36303,N_36389);
nand U37055 (N_37055,N_36388,N_36426);
nand U37056 (N_37056,N_36175,N_36921);
nor U37057 (N_37057,N_36732,N_36032);
xnor U37058 (N_37058,N_36538,N_36933);
xnor U37059 (N_37059,N_36522,N_36170);
nand U37060 (N_37060,N_36575,N_36372);
or U37061 (N_37061,N_36037,N_36647);
nor U37062 (N_37062,N_36077,N_36270);
or U37063 (N_37063,N_36102,N_36543);
nand U37064 (N_37064,N_36463,N_36360);
or U37065 (N_37065,N_36111,N_36271);
or U37066 (N_37066,N_36044,N_36733);
xnor U37067 (N_37067,N_36542,N_36791);
xnor U37068 (N_37068,N_36606,N_36498);
and U37069 (N_37069,N_36695,N_36383);
and U37070 (N_37070,N_36824,N_36506);
or U37071 (N_37071,N_36075,N_36602);
xnor U37072 (N_37072,N_36250,N_36539);
nor U37073 (N_37073,N_36837,N_36839);
and U37074 (N_37074,N_36528,N_36599);
nor U37075 (N_37075,N_36530,N_36777);
or U37076 (N_37076,N_36441,N_36384);
xnor U37077 (N_37077,N_36424,N_36920);
nor U37078 (N_37078,N_36890,N_36156);
nor U37079 (N_37079,N_36585,N_36431);
nor U37080 (N_37080,N_36554,N_36645);
or U37081 (N_37081,N_36479,N_36818);
nand U37082 (N_37082,N_36700,N_36725);
nor U37083 (N_37083,N_36423,N_36570);
nor U37084 (N_37084,N_36729,N_36896);
xnor U37085 (N_37085,N_36970,N_36339);
and U37086 (N_37086,N_36134,N_36876);
or U37087 (N_37087,N_36936,N_36944);
and U37088 (N_37088,N_36147,N_36994);
nand U37089 (N_37089,N_36347,N_36184);
or U37090 (N_37090,N_36097,N_36919);
nand U37091 (N_37091,N_36008,N_36116);
xor U37092 (N_37092,N_36513,N_36676);
or U37093 (N_37093,N_36174,N_36359);
nor U37094 (N_37094,N_36406,N_36738);
or U37095 (N_37095,N_36687,N_36247);
or U37096 (N_37096,N_36943,N_36879);
or U37097 (N_37097,N_36254,N_36971);
or U37098 (N_37098,N_36637,N_36734);
or U37099 (N_37099,N_36290,N_36630);
or U37100 (N_37100,N_36039,N_36085);
xnor U37101 (N_37101,N_36251,N_36356);
nor U37102 (N_37102,N_36243,N_36975);
and U37103 (N_37103,N_36051,N_36411);
or U37104 (N_37104,N_36807,N_36100);
nand U37105 (N_37105,N_36625,N_36120);
nor U37106 (N_37106,N_36235,N_36814);
nor U37107 (N_37107,N_36713,N_36547);
nand U37108 (N_37108,N_36666,N_36091);
and U37109 (N_37109,N_36838,N_36278);
or U37110 (N_37110,N_36601,N_36571);
xor U37111 (N_37111,N_36762,N_36022);
nor U37112 (N_37112,N_36133,N_36686);
and U37113 (N_37113,N_36736,N_36756);
nand U37114 (N_37114,N_36495,N_36312);
nor U37115 (N_37115,N_36443,N_36819);
and U37116 (N_37116,N_36983,N_36808);
or U37117 (N_37117,N_36924,N_36241);
nand U37118 (N_37118,N_36245,N_36158);
xnor U37119 (N_37119,N_36285,N_36767);
nand U37120 (N_37120,N_36552,N_36512);
nor U37121 (N_37121,N_36531,N_36314);
or U37122 (N_37122,N_36284,N_36648);
or U37123 (N_37123,N_36357,N_36343);
nor U37124 (N_37124,N_36962,N_36413);
nand U37125 (N_37125,N_36400,N_36950);
and U37126 (N_37126,N_36168,N_36797);
nand U37127 (N_37127,N_36244,N_36151);
nor U37128 (N_37128,N_36948,N_36361);
xor U37129 (N_37129,N_36627,N_36882);
nand U37130 (N_37130,N_36801,N_36619);
nor U37131 (N_37131,N_36353,N_36279);
nor U37132 (N_37132,N_36502,N_36006);
or U37133 (N_37133,N_36153,N_36726);
and U37134 (N_37134,N_36466,N_36930);
nor U37135 (N_37135,N_36336,N_36392);
nand U37136 (N_37136,N_36013,N_36926);
or U37137 (N_37137,N_36350,N_36412);
xor U37138 (N_37138,N_36856,N_36143);
and U37139 (N_37139,N_36829,N_36234);
nor U37140 (N_37140,N_36160,N_36586);
nand U37141 (N_37141,N_36772,N_36354);
nor U37142 (N_37142,N_36817,N_36603);
xnor U37143 (N_37143,N_36963,N_36566);
nor U37144 (N_37144,N_36080,N_36226);
and U37145 (N_37145,N_36987,N_36827);
and U37146 (N_37146,N_36773,N_36311);
nor U37147 (N_37147,N_36678,N_36004);
nor U37148 (N_37148,N_36456,N_36889);
and U37149 (N_37149,N_36060,N_36764);
or U37150 (N_37150,N_36381,N_36949);
nor U37151 (N_37151,N_36723,N_36089);
xnor U37152 (N_37152,N_36988,N_36231);
xor U37153 (N_37153,N_36622,N_36515);
nor U37154 (N_37154,N_36054,N_36149);
xnor U37155 (N_37155,N_36514,N_36855);
xnor U37156 (N_37156,N_36386,N_36870);
nor U37157 (N_37157,N_36107,N_36368);
nor U37158 (N_37158,N_36899,N_36878);
or U37159 (N_37159,N_36544,N_36410);
or U37160 (N_37160,N_36346,N_36395);
nand U37161 (N_37161,N_36179,N_36480);
or U37162 (N_37162,N_36197,N_36783);
nand U37163 (N_37163,N_36209,N_36407);
xor U37164 (N_37164,N_36268,N_36587);
and U37165 (N_37165,N_36364,N_36917);
or U37166 (N_37166,N_36698,N_36786);
xnor U37167 (N_37167,N_36952,N_36562);
nor U37168 (N_37168,N_36671,N_36041);
and U37169 (N_37169,N_36564,N_36313);
and U37170 (N_37170,N_36996,N_36078);
nor U37171 (N_37171,N_36123,N_36984);
and U37172 (N_37172,N_36052,N_36428);
nand U37173 (N_37173,N_36066,N_36594);
xor U37174 (N_37174,N_36913,N_36815);
or U37175 (N_37175,N_36167,N_36344);
xnor U37176 (N_37176,N_36317,N_36187);
nor U37177 (N_37177,N_36639,N_36263);
and U37178 (N_37178,N_36968,N_36296);
nor U37179 (N_37179,N_36292,N_36935);
or U37180 (N_37180,N_36385,N_36655);
xnor U37181 (N_37181,N_36709,N_36592);
nand U37182 (N_37182,N_36802,N_36875);
and U37183 (N_37183,N_36497,N_36568);
xor U37184 (N_37184,N_36799,N_36216);
xnor U37185 (N_37185,N_36795,N_36931);
nand U37186 (N_37186,N_36178,N_36417);
and U37187 (N_37187,N_36613,N_36803);
and U37188 (N_37188,N_36481,N_36934);
nand U37189 (N_37189,N_36633,N_36932);
or U37190 (N_37190,N_36597,N_36653);
nand U37191 (N_37191,N_36205,N_36717);
and U37192 (N_37192,N_36922,N_36898);
nor U37193 (N_37193,N_36977,N_36172);
nor U37194 (N_37194,N_36330,N_36155);
and U37195 (N_37195,N_36549,N_36193);
nand U37196 (N_37196,N_36236,N_36393);
nand U37197 (N_37197,N_36825,N_36103);
nor U37198 (N_37198,N_36654,N_36293);
nor U37199 (N_37199,N_36390,N_36704);
or U37200 (N_37200,N_36272,N_36663);
and U37201 (N_37201,N_36955,N_36883);
xnor U37202 (N_37202,N_36868,N_36403);
nand U37203 (N_37203,N_36535,N_36121);
xnor U37204 (N_37204,N_36452,N_36998);
or U37205 (N_37205,N_36448,N_36192);
nor U37206 (N_37206,N_36517,N_36558);
nor U37207 (N_37207,N_36573,N_36985);
and U37208 (N_37208,N_36334,N_36569);
nor U37209 (N_37209,N_36711,N_36173);
xnor U37210 (N_37210,N_36742,N_36972);
nand U37211 (N_37211,N_36618,N_36034);
nand U37212 (N_37212,N_36861,N_36914);
and U37213 (N_37213,N_36057,N_36691);
or U37214 (N_37214,N_36204,N_36953);
or U37215 (N_37215,N_36679,N_36238);
or U37216 (N_37216,N_36058,N_36685);
xor U37217 (N_37217,N_36778,N_36574);
nand U37218 (N_37218,N_36188,N_36763);
nor U37219 (N_37219,N_36084,N_36532);
nor U37220 (N_37220,N_36050,N_36110);
or U37221 (N_37221,N_36048,N_36140);
or U37222 (N_37222,N_36947,N_36146);
or U37223 (N_37223,N_36112,N_36820);
and U37224 (N_37224,N_36578,N_36163);
or U37225 (N_37225,N_36394,N_36617);
nor U37226 (N_37226,N_36096,N_36901);
and U37227 (N_37227,N_36304,N_36526);
or U37228 (N_37228,N_36477,N_36992);
xor U37229 (N_37229,N_36262,N_36881);
nand U37230 (N_37230,N_36461,N_36527);
xnor U37231 (N_37231,N_36504,N_36708);
nand U37232 (N_37232,N_36813,N_36768);
or U37233 (N_37233,N_36451,N_36928);
nor U37234 (N_37234,N_36959,N_36308);
xor U37235 (N_37235,N_36665,N_36176);
and U37236 (N_37236,N_36707,N_36420);
or U37237 (N_37237,N_36092,N_36553);
or U37238 (N_37238,N_36754,N_36072);
and U37239 (N_37239,N_36490,N_36101);
and U37240 (N_37240,N_36659,N_36476);
or U37241 (N_37241,N_36525,N_36682);
or U37242 (N_37242,N_36455,N_36213);
nor U37243 (N_37243,N_36661,N_36657);
nor U37244 (N_37244,N_36232,N_36775);
nand U37245 (N_37245,N_36169,N_36758);
or U37246 (N_37246,N_36217,N_36960);
and U37247 (N_37247,N_36697,N_36548);
and U37248 (N_37248,N_36472,N_36005);
xor U37249 (N_37249,N_36379,N_36716);
nor U37250 (N_37250,N_36650,N_36858);
and U37251 (N_37251,N_36989,N_36957);
and U37252 (N_37252,N_36995,N_36969);
nor U37253 (N_37253,N_36484,N_36233);
and U37254 (N_37254,N_36246,N_36316);
xnor U37255 (N_37255,N_36918,N_36286);
or U37256 (N_37256,N_36846,N_36677);
nor U37257 (N_37257,N_36218,N_36070);
nor U37258 (N_37258,N_36469,N_36546);
and U37259 (N_37259,N_36701,N_36509);
nand U37260 (N_37260,N_36162,N_36511);
nor U37261 (N_37261,N_36055,N_36871);
nand U37262 (N_37262,N_36332,N_36598);
nor U37263 (N_37263,N_36634,N_36207);
nor U37264 (N_37264,N_36997,N_36788);
nand U37265 (N_37265,N_36266,N_36433);
nand U37266 (N_37266,N_36026,N_36626);
nor U37267 (N_37267,N_36404,N_36321);
or U37268 (N_37268,N_36790,N_36139);
and U37269 (N_37269,N_36399,N_36259);
nor U37270 (N_37270,N_36641,N_36488);
or U37271 (N_37271,N_36699,N_36737);
and U37272 (N_37272,N_36787,N_36915);
or U37273 (N_37273,N_36449,N_36999);
nand U37274 (N_37274,N_36264,N_36122);
nor U37275 (N_37275,N_36581,N_36454);
nand U37276 (N_37276,N_36152,N_36642);
nor U37277 (N_37277,N_36436,N_36727);
nand U37278 (N_37278,N_36299,N_36567);
or U37279 (N_37279,N_36540,N_36593);
nor U37280 (N_37280,N_36370,N_36249);
and U37281 (N_37281,N_36323,N_36604);
nand U37282 (N_37282,N_36047,N_36909);
xnor U37283 (N_37283,N_36018,N_36735);
and U37284 (N_37284,N_36468,N_36805);
or U37285 (N_37285,N_36759,N_36225);
xnor U37286 (N_37286,N_36976,N_36194);
or U37287 (N_37287,N_36482,N_36485);
xor U37288 (N_37288,N_36757,N_36171);
nand U37289 (N_37289,N_36545,N_36028);
nand U37290 (N_37290,N_36518,N_36189);
nand U37291 (N_37291,N_36811,N_36796);
nand U37292 (N_37292,N_36582,N_36688);
and U37293 (N_37293,N_36391,N_36079);
xor U37294 (N_37294,N_36442,N_36789);
and U37295 (N_37295,N_36847,N_36904);
or U37296 (N_37296,N_36589,N_36945);
or U37297 (N_37297,N_36033,N_36062);
xnor U37298 (N_37298,N_36916,N_36074);
nor U37299 (N_37299,N_36021,N_36275);
nand U37300 (N_37300,N_36297,N_36860);
xnor U37301 (N_37301,N_36923,N_36854);
or U37302 (N_37302,N_36752,N_36201);
nor U37303 (N_37303,N_36031,N_36237);
or U37304 (N_37304,N_36503,N_36869);
xor U37305 (N_37305,N_36743,N_36277);
nor U37306 (N_37306,N_36369,N_36591);
or U37307 (N_37307,N_36362,N_36776);
and U37308 (N_37308,N_36487,N_36157);
nand U37309 (N_37309,N_36508,N_36694);
and U37310 (N_37310,N_36265,N_36925);
nor U37311 (N_37311,N_36636,N_36067);
nor U37312 (N_37312,N_36450,N_36907);
xnor U37313 (N_37313,N_36145,N_36942);
nand U37314 (N_37314,N_36185,N_36724);
nor U37315 (N_37315,N_36114,N_36714);
xnor U37316 (N_37316,N_36434,N_36229);
xor U37317 (N_37317,N_36816,N_36534);
xnor U37318 (N_37318,N_36874,N_36705);
nor U37319 (N_37319,N_36220,N_36873);
xor U37320 (N_37320,N_36056,N_36895);
nand U37321 (N_37321,N_36973,N_36387);
xnor U37322 (N_37322,N_36629,N_36842);
nand U37323 (N_37323,N_36186,N_36414);
nand U37324 (N_37324,N_36761,N_36274);
nor U37325 (N_37325,N_36291,N_36774);
or U37326 (N_37326,N_36739,N_36030);
nand U37327 (N_37327,N_36373,N_36090);
nand U37328 (N_37328,N_36845,N_36572);
xor U37329 (N_37329,N_36753,N_36730);
nand U37330 (N_37330,N_36610,N_36956);
nor U37331 (N_37331,N_36492,N_36309);
xor U37332 (N_37332,N_36267,N_36154);
nand U37333 (N_37333,N_36958,N_36809);
xor U37334 (N_37334,N_36095,N_36126);
nand U37335 (N_37335,N_36696,N_36053);
xor U37336 (N_37336,N_36721,N_36380);
and U37337 (N_37337,N_36905,N_36831);
or U37338 (N_37338,N_36024,N_36049);
nor U37339 (N_37339,N_36652,N_36673);
nand U37340 (N_37340,N_36081,N_36559);
and U37341 (N_37341,N_36242,N_36979);
and U37342 (N_37342,N_36144,N_36703);
nor U37343 (N_37343,N_36475,N_36083);
and U37344 (N_37344,N_36834,N_36198);
xor U37345 (N_37345,N_36396,N_36348);
xnor U37346 (N_37346,N_36751,N_36821);
nor U37347 (N_37347,N_36986,N_36020);
or U37348 (N_37348,N_36003,N_36941);
and U37349 (N_37349,N_36780,N_36252);
nor U37350 (N_37350,N_36338,N_36318);
or U37351 (N_37351,N_36483,N_36991);
or U37352 (N_37352,N_36710,N_36556);
nor U37353 (N_37353,N_36223,N_36857);
xnor U37354 (N_37354,N_36664,N_36702);
xor U37355 (N_37355,N_36551,N_36507);
nand U37356 (N_37356,N_36319,N_36722);
or U37357 (N_37357,N_36307,N_36849);
nand U37358 (N_37358,N_36900,N_36043);
and U37359 (N_37359,N_36320,N_36927);
and U37360 (N_37360,N_36439,N_36099);
and U37361 (N_37361,N_36720,N_36844);
xnor U37362 (N_37362,N_36398,N_36341);
or U37363 (N_37363,N_36203,N_36195);
nor U37364 (N_37364,N_36086,N_36408);
and U37365 (N_37365,N_36325,N_36105);
or U37366 (N_37366,N_36891,N_36444);
and U37367 (N_37367,N_36059,N_36533);
nor U37368 (N_37368,N_36521,N_36087);
nand U37369 (N_37369,N_36966,N_36615);
xor U37370 (N_37370,N_36418,N_36010);
nand U37371 (N_37371,N_36215,N_36429);
and U37372 (N_37372,N_36683,N_36331);
nor U37373 (N_37373,N_36982,N_36865);
and U37374 (N_37374,N_36253,N_36689);
nand U37375 (N_37375,N_36939,N_36377);
nand U37376 (N_37376,N_36823,N_36093);
and U37377 (N_37377,N_36255,N_36470);
or U37378 (N_37378,N_36076,N_36524);
or U37379 (N_37379,N_36130,N_36258);
or U37380 (N_37380,N_36306,N_36324);
nor U37381 (N_37381,N_36210,N_36580);
and U37382 (N_37382,N_36221,N_36281);
nor U37383 (N_37383,N_36590,N_36419);
xor U37384 (N_37384,N_36302,N_36561);
xor U37385 (N_37385,N_36866,N_36137);
or U37386 (N_37386,N_36063,N_36329);
nand U37387 (N_37387,N_36138,N_36863);
nand U37388 (N_37388,N_36199,N_36519);
or U37389 (N_37389,N_36437,N_36853);
nor U37390 (N_37390,N_36082,N_36667);
nor U37391 (N_37391,N_36042,N_36965);
and U37392 (N_37392,N_36529,N_36125);
xor U37393 (N_37393,N_36131,N_36577);
nor U37394 (N_37394,N_36669,N_36073);
or U37395 (N_37395,N_36011,N_36027);
and U37396 (N_37396,N_36191,N_36161);
nand U37397 (N_37397,N_36473,N_36583);
and U37398 (N_37398,N_36071,N_36903);
and U37399 (N_37399,N_36609,N_36785);
xor U37400 (N_37400,N_36635,N_36447);
and U37401 (N_37401,N_36632,N_36851);
or U37402 (N_37402,N_36142,N_36036);
nand U37403 (N_37403,N_36023,N_36731);
or U37404 (N_37404,N_36349,N_36745);
nor U37405 (N_37405,N_36841,N_36541);
nand U37406 (N_37406,N_36322,N_36565);
nor U37407 (N_37407,N_36993,N_36280);
and U37408 (N_37408,N_36196,N_36260);
nand U37409 (N_37409,N_36273,N_36579);
and U37410 (N_37410,N_36651,N_36718);
or U37411 (N_37411,N_36211,N_36893);
or U37412 (N_37412,N_36460,N_36640);
and U37413 (N_37413,N_36402,N_36440);
nor U37414 (N_37414,N_36516,N_36464);
nand U37415 (N_37415,N_36025,N_36510);
nand U37416 (N_37416,N_36607,N_36850);
xor U37417 (N_37417,N_36712,N_36911);
nand U37418 (N_37418,N_36822,N_36239);
nor U37419 (N_37419,N_36681,N_36680);
nor U37420 (N_37420,N_36219,N_36746);
xnor U37421 (N_37421,N_36536,N_36401);
or U37422 (N_37422,N_36611,N_36230);
nor U37423 (N_37423,N_36951,N_36938);
or U37424 (N_37424,N_36113,N_36068);
nor U37425 (N_37425,N_36638,N_36940);
xnor U37426 (N_37426,N_36769,N_36124);
nor U37427 (N_37427,N_36415,N_36202);
nor U37428 (N_37428,N_36376,N_36656);
or U37429 (N_37429,N_36065,N_36159);
nand U37430 (N_37430,N_36352,N_36693);
nand U37431 (N_37431,N_36660,N_36690);
or U37432 (N_37432,N_36045,N_36649);
or U37433 (N_37433,N_36843,N_36852);
nand U37434 (N_37434,N_36692,N_36560);
or U37435 (N_37435,N_36888,N_36840);
and U37436 (N_37436,N_36792,N_36588);
xor U37437 (N_37437,N_36150,N_36446);
or U37438 (N_37438,N_36520,N_36550);
nand U37439 (N_37439,N_36064,N_36612);
or U37440 (N_37440,N_36127,N_36600);
or U37441 (N_37441,N_36832,N_36375);
nor U37442 (N_37442,N_36289,N_36261);
xnor U37443 (N_37443,N_36276,N_36623);
nand U37444 (N_37444,N_36458,N_36445);
nand U37445 (N_37445,N_36029,N_36596);
and U37446 (N_37446,N_36115,N_36104);
nor U37447 (N_37447,N_36749,N_36496);
nand U37448 (N_37448,N_36183,N_36135);
nand U37449 (N_37449,N_36214,N_36812);
nor U37450 (N_37450,N_36014,N_36046);
xnor U37451 (N_37451,N_36088,N_36471);
xor U37452 (N_37452,N_36884,N_36867);
nor U37453 (N_37453,N_36614,N_36295);
nand U37454 (N_37454,N_36782,N_36779);
nor U37455 (N_37455,N_36228,N_36810);
or U37456 (N_37456,N_36019,N_36662);
and U37457 (N_37457,N_36240,N_36885);
nor U37458 (N_37458,N_36382,N_36478);
and U37459 (N_37459,N_36557,N_36310);
and U37460 (N_37460,N_36038,N_36886);
and U37461 (N_37461,N_36017,N_36747);
nand U37462 (N_37462,N_36467,N_36282);
or U37463 (N_37463,N_36771,N_36964);
xnor U37464 (N_37464,N_36109,N_36643);
or U37465 (N_37465,N_36961,N_36929);
and U37466 (N_37466,N_36181,N_36128);
xnor U37467 (N_37467,N_36016,N_36793);
and U37468 (N_37468,N_36631,N_36355);
nor U37469 (N_37469,N_36453,N_36283);
nor U37470 (N_37470,N_36628,N_36335);
nor U37471 (N_37471,N_36328,N_36301);
nand U37472 (N_37472,N_36465,N_36505);
or U37473 (N_37473,N_36563,N_36106);
nor U37474 (N_37474,N_36165,N_36798);
and U37475 (N_37475,N_36974,N_36208);
and U37476 (N_37476,N_36978,N_36706);
nand U37477 (N_37477,N_36765,N_36416);
and U37478 (N_37478,N_36094,N_36222);
and U37479 (N_37479,N_36422,N_36954);
xnor U37480 (N_37480,N_36327,N_36365);
and U37481 (N_37481,N_36887,N_36427);
nand U37482 (N_37482,N_36397,N_36910);
nand U37483 (N_37483,N_36906,N_36333);
nor U37484 (N_37484,N_36760,N_36035);
xnor U37485 (N_37485,N_36864,N_36374);
and U37486 (N_37486,N_36378,N_36967);
and U37487 (N_37487,N_36180,N_36345);
and U37488 (N_37488,N_36300,N_36457);
xor U37489 (N_37489,N_36862,N_36182);
or U37490 (N_37490,N_36744,N_36719);
and U37491 (N_37491,N_36493,N_36007);
and U37492 (N_37492,N_36728,N_36009);
nand U37493 (N_37493,N_36489,N_36486);
nand U37494 (N_37494,N_36646,N_36892);
xor U37495 (N_37495,N_36363,N_36462);
and U37496 (N_37496,N_36500,N_36177);
nor U37497 (N_37497,N_36621,N_36459);
or U37498 (N_37498,N_36605,N_36990);
nand U37499 (N_37499,N_36118,N_36164);
or U37500 (N_37500,N_36555,N_36101);
xnor U37501 (N_37501,N_36951,N_36854);
nand U37502 (N_37502,N_36806,N_36552);
xor U37503 (N_37503,N_36174,N_36116);
and U37504 (N_37504,N_36733,N_36908);
nor U37505 (N_37505,N_36185,N_36209);
nand U37506 (N_37506,N_36689,N_36761);
xor U37507 (N_37507,N_36522,N_36548);
nor U37508 (N_37508,N_36345,N_36253);
or U37509 (N_37509,N_36138,N_36991);
and U37510 (N_37510,N_36280,N_36272);
xor U37511 (N_37511,N_36357,N_36517);
nor U37512 (N_37512,N_36015,N_36652);
or U37513 (N_37513,N_36261,N_36285);
and U37514 (N_37514,N_36504,N_36282);
nand U37515 (N_37515,N_36550,N_36043);
nand U37516 (N_37516,N_36712,N_36689);
or U37517 (N_37517,N_36473,N_36288);
or U37518 (N_37518,N_36939,N_36591);
nand U37519 (N_37519,N_36984,N_36574);
nor U37520 (N_37520,N_36172,N_36053);
nand U37521 (N_37521,N_36139,N_36052);
xnor U37522 (N_37522,N_36795,N_36711);
and U37523 (N_37523,N_36162,N_36565);
and U37524 (N_37524,N_36719,N_36105);
and U37525 (N_37525,N_36854,N_36308);
nand U37526 (N_37526,N_36249,N_36733);
xnor U37527 (N_37527,N_36532,N_36757);
or U37528 (N_37528,N_36780,N_36772);
xor U37529 (N_37529,N_36383,N_36026);
nor U37530 (N_37530,N_36855,N_36703);
or U37531 (N_37531,N_36515,N_36065);
nor U37532 (N_37532,N_36946,N_36972);
xor U37533 (N_37533,N_36683,N_36882);
nor U37534 (N_37534,N_36422,N_36749);
nor U37535 (N_37535,N_36709,N_36995);
xnor U37536 (N_37536,N_36087,N_36155);
nor U37537 (N_37537,N_36287,N_36702);
or U37538 (N_37538,N_36815,N_36591);
nand U37539 (N_37539,N_36324,N_36511);
or U37540 (N_37540,N_36291,N_36417);
and U37541 (N_37541,N_36849,N_36440);
nand U37542 (N_37542,N_36487,N_36366);
or U37543 (N_37543,N_36130,N_36870);
or U37544 (N_37544,N_36959,N_36455);
or U37545 (N_37545,N_36695,N_36110);
or U37546 (N_37546,N_36810,N_36849);
xor U37547 (N_37547,N_36278,N_36682);
or U37548 (N_37548,N_36521,N_36306);
nor U37549 (N_37549,N_36183,N_36756);
xor U37550 (N_37550,N_36297,N_36606);
or U37551 (N_37551,N_36716,N_36626);
or U37552 (N_37552,N_36396,N_36944);
and U37553 (N_37553,N_36148,N_36952);
or U37554 (N_37554,N_36345,N_36720);
xnor U37555 (N_37555,N_36110,N_36059);
and U37556 (N_37556,N_36128,N_36702);
or U37557 (N_37557,N_36304,N_36165);
and U37558 (N_37558,N_36458,N_36877);
nand U37559 (N_37559,N_36397,N_36273);
nor U37560 (N_37560,N_36632,N_36951);
or U37561 (N_37561,N_36455,N_36780);
nor U37562 (N_37562,N_36191,N_36498);
xor U37563 (N_37563,N_36298,N_36746);
nand U37564 (N_37564,N_36451,N_36791);
xor U37565 (N_37565,N_36945,N_36973);
and U37566 (N_37566,N_36697,N_36658);
nand U37567 (N_37567,N_36285,N_36536);
nor U37568 (N_37568,N_36076,N_36700);
xor U37569 (N_37569,N_36446,N_36451);
or U37570 (N_37570,N_36361,N_36754);
xor U37571 (N_37571,N_36640,N_36151);
nand U37572 (N_37572,N_36083,N_36209);
nor U37573 (N_37573,N_36159,N_36441);
nor U37574 (N_37574,N_36334,N_36259);
nand U37575 (N_37575,N_36774,N_36916);
nand U37576 (N_37576,N_36304,N_36058);
xnor U37577 (N_37577,N_36365,N_36542);
xnor U37578 (N_37578,N_36019,N_36467);
xor U37579 (N_37579,N_36033,N_36793);
xnor U37580 (N_37580,N_36973,N_36284);
nand U37581 (N_37581,N_36904,N_36307);
xor U37582 (N_37582,N_36914,N_36791);
and U37583 (N_37583,N_36328,N_36436);
xor U37584 (N_37584,N_36264,N_36118);
and U37585 (N_37585,N_36167,N_36061);
nand U37586 (N_37586,N_36905,N_36536);
and U37587 (N_37587,N_36487,N_36243);
and U37588 (N_37588,N_36306,N_36972);
nor U37589 (N_37589,N_36338,N_36670);
and U37590 (N_37590,N_36720,N_36586);
xnor U37591 (N_37591,N_36815,N_36407);
or U37592 (N_37592,N_36186,N_36145);
nand U37593 (N_37593,N_36178,N_36705);
xor U37594 (N_37594,N_36359,N_36261);
or U37595 (N_37595,N_36736,N_36005);
and U37596 (N_37596,N_36808,N_36327);
xnor U37597 (N_37597,N_36906,N_36674);
nand U37598 (N_37598,N_36243,N_36306);
or U37599 (N_37599,N_36033,N_36487);
and U37600 (N_37600,N_36922,N_36578);
nor U37601 (N_37601,N_36942,N_36563);
or U37602 (N_37602,N_36348,N_36824);
xor U37603 (N_37603,N_36244,N_36531);
or U37604 (N_37604,N_36639,N_36500);
and U37605 (N_37605,N_36789,N_36343);
nand U37606 (N_37606,N_36411,N_36191);
nand U37607 (N_37607,N_36930,N_36581);
and U37608 (N_37608,N_36081,N_36611);
nand U37609 (N_37609,N_36571,N_36711);
xor U37610 (N_37610,N_36045,N_36449);
nand U37611 (N_37611,N_36323,N_36065);
nor U37612 (N_37612,N_36770,N_36368);
and U37613 (N_37613,N_36128,N_36792);
nor U37614 (N_37614,N_36836,N_36930);
nand U37615 (N_37615,N_36808,N_36732);
nand U37616 (N_37616,N_36379,N_36082);
nor U37617 (N_37617,N_36566,N_36126);
xnor U37618 (N_37618,N_36767,N_36544);
nor U37619 (N_37619,N_36887,N_36070);
xnor U37620 (N_37620,N_36739,N_36708);
and U37621 (N_37621,N_36735,N_36466);
xnor U37622 (N_37622,N_36736,N_36515);
nor U37623 (N_37623,N_36705,N_36211);
xor U37624 (N_37624,N_36416,N_36244);
and U37625 (N_37625,N_36363,N_36959);
nand U37626 (N_37626,N_36772,N_36905);
and U37627 (N_37627,N_36035,N_36904);
nor U37628 (N_37628,N_36321,N_36920);
or U37629 (N_37629,N_36529,N_36826);
nor U37630 (N_37630,N_36039,N_36537);
nand U37631 (N_37631,N_36397,N_36426);
and U37632 (N_37632,N_36868,N_36406);
nor U37633 (N_37633,N_36189,N_36238);
or U37634 (N_37634,N_36250,N_36938);
nor U37635 (N_37635,N_36278,N_36875);
nand U37636 (N_37636,N_36478,N_36571);
xnor U37637 (N_37637,N_36396,N_36448);
xnor U37638 (N_37638,N_36728,N_36788);
or U37639 (N_37639,N_36122,N_36306);
or U37640 (N_37640,N_36937,N_36848);
xor U37641 (N_37641,N_36378,N_36347);
xnor U37642 (N_37642,N_36103,N_36125);
or U37643 (N_37643,N_36576,N_36459);
and U37644 (N_37644,N_36104,N_36967);
nor U37645 (N_37645,N_36632,N_36943);
or U37646 (N_37646,N_36792,N_36959);
or U37647 (N_37647,N_36726,N_36113);
or U37648 (N_37648,N_36278,N_36429);
nand U37649 (N_37649,N_36465,N_36522);
nor U37650 (N_37650,N_36602,N_36553);
and U37651 (N_37651,N_36029,N_36033);
xnor U37652 (N_37652,N_36419,N_36069);
or U37653 (N_37653,N_36082,N_36435);
nand U37654 (N_37654,N_36804,N_36251);
or U37655 (N_37655,N_36067,N_36899);
xnor U37656 (N_37656,N_36364,N_36990);
nand U37657 (N_37657,N_36157,N_36529);
nor U37658 (N_37658,N_36930,N_36392);
or U37659 (N_37659,N_36124,N_36597);
or U37660 (N_37660,N_36139,N_36319);
nor U37661 (N_37661,N_36902,N_36572);
nor U37662 (N_37662,N_36831,N_36471);
nor U37663 (N_37663,N_36950,N_36845);
nand U37664 (N_37664,N_36664,N_36742);
nand U37665 (N_37665,N_36184,N_36694);
xor U37666 (N_37666,N_36385,N_36092);
nand U37667 (N_37667,N_36550,N_36334);
nand U37668 (N_37668,N_36171,N_36243);
and U37669 (N_37669,N_36116,N_36844);
or U37670 (N_37670,N_36251,N_36159);
xor U37671 (N_37671,N_36120,N_36192);
or U37672 (N_37672,N_36248,N_36215);
and U37673 (N_37673,N_36268,N_36183);
or U37674 (N_37674,N_36882,N_36156);
nand U37675 (N_37675,N_36465,N_36499);
nand U37676 (N_37676,N_36486,N_36215);
xor U37677 (N_37677,N_36214,N_36900);
and U37678 (N_37678,N_36534,N_36006);
or U37679 (N_37679,N_36181,N_36672);
xnor U37680 (N_37680,N_36040,N_36230);
and U37681 (N_37681,N_36360,N_36636);
xor U37682 (N_37682,N_36018,N_36292);
nand U37683 (N_37683,N_36898,N_36153);
and U37684 (N_37684,N_36348,N_36638);
and U37685 (N_37685,N_36906,N_36147);
nand U37686 (N_37686,N_36391,N_36536);
nand U37687 (N_37687,N_36075,N_36972);
or U37688 (N_37688,N_36817,N_36958);
or U37689 (N_37689,N_36738,N_36872);
nand U37690 (N_37690,N_36185,N_36981);
nor U37691 (N_37691,N_36650,N_36504);
and U37692 (N_37692,N_36283,N_36112);
nand U37693 (N_37693,N_36519,N_36652);
and U37694 (N_37694,N_36844,N_36656);
nor U37695 (N_37695,N_36964,N_36605);
nand U37696 (N_37696,N_36745,N_36686);
nand U37697 (N_37697,N_36754,N_36417);
xor U37698 (N_37698,N_36763,N_36670);
nor U37699 (N_37699,N_36821,N_36931);
xor U37700 (N_37700,N_36754,N_36859);
nand U37701 (N_37701,N_36440,N_36769);
nand U37702 (N_37702,N_36660,N_36101);
nand U37703 (N_37703,N_36223,N_36781);
and U37704 (N_37704,N_36029,N_36819);
and U37705 (N_37705,N_36736,N_36690);
nor U37706 (N_37706,N_36123,N_36694);
nor U37707 (N_37707,N_36711,N_36758);
nor U37708 (N_37708,N_36553,N_36792);
nand U37709 (N_37709,N_36361,N_36526);
nand U37710 (N_37710,N_36731,N_36442);
xor U37711 (N_37711,N_36938,N_36597);
nor U37712 (N_37712,N_36601,N_36958);
nor U37713 (N_37713,N_36688,N_36976);
nand U37714 (N_37714,N_36890,N_36508);
xnor U37715 (N_37715,N_36283,N_36588);
xnor U37716 (N_37716,N_36937,N_36036);
nor U37717 (N_37717,N_36715,N_36649);
xor U37718 (N_37718,N_36315,N_36416);
or U37719 (N_37719,N_36662,N_36239);
or U37720 (N_37720,N_36096,N_36178);
xnor U37721 (N_37721,N_36115,N_36752);
nor U37722 (N_37722,N_36750,N_36152);
nor U37723 (N_37723,N_36016,N_36526);
nand U37724 (N_37724,N_36410,N_36756);
or U37725 (N_37725,N_36542,N_36318);
xnor U37726 (N_37726,N_36652,N_36169);
nor U37727 (N_37727,N_36242,N_36667);
nor U37728 (N_37728,N_36052,N_36550);
xor U37729 (N_37729,N_36561,N_36423);
nand U37730 (N_37730,N_36801,N_36222);
and U37731 (N_37731,N_36656,N_36171);
xnor U37732 (N_37732,N_36439,N_36036);
nor U37733 (N_37733,N_36121,N_36769);
xnor U37734 (N_37734,N_36083,N_36970);
nand U37735 (N_37735,N_36314,N_36965);
or U37736 (N_37736,N_36761,N_36491);
xor U37737 (N_37737,N_36981,N_36463);
and U37738 (N_37738,N_36828,N_36212);
nand U37739 (N_37739,N_36458,N_36216);
nor U37740 (N_37740,N_36634,N_36364);
xor U37741 (N_37741,N_36362,N_36556);
or U37742 (N_37742,N_36349,N_36282);
nor U37743 (N_37743,N_36550,N_36629);
or U37744 (N_37744,N_36511,N_36271);
or U37745 (N_37745,N_36929,N_36019);
and U37746 (N_37746,N_36617,N_36614);
nand U37747 (N_37747,N_36962,N_36737);
xnor U37748 (N_37748,N_36260,N_36569);
nor U37749 (N_37749,N_36871,N_36304);
xor U37750 (N_37750,N_36448,N_36318);
xor U37751 (N_37751,N_36858,N_36203);
xnor U37752 (N_37752,N_36859,N_36896);
or U37753 (N_37753,N_36280,N_36290);
nand U37754 (N_37754,N_36524,N_36928);
and U37755 (N_37755,N_36723,N_36798);
nor U37756 (N_37756,N_36329,N_36975);
nand U37757 (N_37757,N_36016,N_36679);
nand U37758 (N_37758,N_36053,N_36820);
xnor U37759 (N_37759,N_36055,N_36299);
nand U37760 (N_37760,N_36121,N_36854);
or U37761 (N_37761,N_36032,N_36425);
nor U37762 (N_37762,N_36054,N_36283);
or U37763 (N_37763,N_36647,N_36192);
nand U37764 (N_37764,N_36133,N_36827);
and U37765 (N_37765,N_36499,N_36668);
or U37766 (N_37766,N_36999,N_36703);
nor U37767 (N_37767,N_36192,N_36749);
and U37768 (N_37768,N_36700,N_36748);
nand U37769 (N_37769,N_36470,N_36730);
xor U37770 (N_37770,N_36390,N_36270);
and U37771 (N_37771,N_36038,N_36789);
and U37772 (N_37772,N_36611,N_36084);
nand U37773 (N_37773,N_36109,N_36821);
nand U37774 (N_37774,N_36852,N_36742);
nand U37775 (N_37775,N_36061,N_36150);
or U37776 (N_37776,N_36336,N_36706);
or U37777 (N_37777,N_36153,N_36972);
or U37778 (N_37778,N_36093,N_36850);
and U37779 (N_37779,N_36018,N_36453);
and U37780 (N_37780,N_36695,N_36584);
nand U37781 (N_37781,N_36343,N_36728);
and U37782 (N_37782,N_36380,N_36525);
nor U37783 (N_37783,N_36683,N_36259);
xor U37784 (N_37784,N_36717,N_36040);
and U37785 (N_37785,N_36861,N_36412);
nand U37786 (N_37786,N_36634,N_36369);
nand U37787 (N_37787,N_36496,N_36455);
nand U37788 (N_37788,N_36448,N_36493);
nand U37789 (N_37789,N_36967,N_36168);
or U37790 (N_37790,N_36307,N_36450);
xnor U37791 (N_37791,N_36342,N_36010);
nand U37792 (N_37792,N_36502,N_36800);
and U37793 (N_37793,N_36771,N_36789);
xnor U37794 (N_37794,N_36746,N_36179);
xor U37795 (N_37795,N_36834,N_36149);
or U37796 (N_37796,N_36795,N_36690);
nand U37797 (N_37797,N_36528,N_36354);
or U37798 (N_37798,N_36201,N_36479);
and U37799 (N_37799,N_36997,N_36028);
xnor U37800 (N_37800,N_36505,N_36427);
nor U37801 (N_37801,N_36105,N_36352);
nor U37802 (N_37802,N_36548,N_36564);
nor U37803 (N_37803,N_36143,N_36534);
and U37804 (N_37804,N_36945,N_36146);
xnor U37805 (N_37805,N_36533,N_36386);
xnor U37806 (N_37806,N_36861,N_36076);
nand U37807 (N_37807,N_36226,N_36681);
and U37808 (N_37808,N_36540,N_36078);
xor U37809 (N_37809,N_36439,N_36682);
and U37810 (N_37810,N_36119,N_36720);
or U37811 (N_37811,N_36832,N_36252);
xor U37812 (N_37812,N_36726,N_36996);
nand U37813 (N_37813,N_36439,N_36746);
or U37814 (N_37814,N_36977,N_36252);
nand U37815 (N_37815,N_36717,N_36082);
nor U37816 (N_37816,N_36468,N_36555);
and U37817 (N_37817,N_36931,N_36149);
nand U37818 (N_37818,N_36842,N_36772);
nand U37819 (N_37819,N_36434,N_36738);
nand U37820 (N_37820,N_36049,N_36935);
nor U37821 (N_37821,N_36066,N_36395);
or U37822 (N_37822,N_36706,N_36207);
nand U37823 (N_37823,N_36233,N_36328);
nand U37824 (N_37824,N_36602,N_36007);
or U37825 (N_37825,N_36715,N_36365);
nor U37826 (N_37826,N_36686,N_36926);
xnor U37827 (N_37827,N_36945,N_36874);
and U37828 (N_37828,N_36142,N_36038);
xnor U37829 (N_37829,N_36211,N_36720);
xnor U37830 (N_37830,N_36334,N_36736);
xor U37831 (N_37831,N_36348,N_36205);
or U37832 (N_37832,N_36699,N_36453);
or U37833 (N_37833,N_36349,N_36472);
and U37834 (N_37834,N_36892,N_36167);
xnor U37835 (N_37835,N_36047,N_36277);
xnor U37836 (N_37836,N_36556,N_36132);
nor U37837 (N_37837,N_36438,N_36702);
and U37838 (N_37838,N_36197,N_36926);
nor U37839 (N_37839,N_36046,N_36542);
nor U37840 (N_37840,N_36004,N_36095);
nor U37841 (N_37841,N_36078,N_36997);
nand U37842 (N_37842,N_36852,N_36428);
and U37843 (N_37843,N_36520,N_36457);
or U37844 (N_37844,N_36748,N_36180);
and U37845 (N_37845,N_36810,N_36687);
xor U37846 (N_37846,N_36604,N_36026);
and U37847 (N_37847,N_36369,N_36339);
nand U37848 (N_37848,N_36986,N_36773);
and U37849 (N_37849,N_36966,N_36147);
and U37850 (N_37850,N_36374,N_36340);
and U37851 (N_37851,N_36810,N_36189);
nand U37852 (N_37852,N_36760,N_36828);
xnor U37853 (N_37853,N_36069,N_36289);
nor U37854 (N_37854,N_36947,N_36822);
xnor U37855 (N_37855,N_36538,N_36814);
nor U37856 (N_37856,N_36600,N_36814);
or U37857 (N_37857,N_36486,N_36859);
xnor U37858 (N_37858,N_36604,N_36123);
or U37859 (N_37859,N_36438,N_36931);
nand U37860 (N_37860,N_36332,N_36077);
xnor U37861 (N_37861,N_36788,N_36276);
nand U37862 (N_37862,N_36496,N_36398);
and U37863 (N_37863,N_36275,N_36265);
and U37864 (N_37864,N_36617,N_36221);
xnor U37865 (N_37865,N_36857,N_36060);
or U37866 (N_37866,N_36243,N_36414);
xor U37867 (N_37867,N_36206,N_36965);
or U37868 (N_37868,N_36532,N_36030);
and U37869 (N_37869,N_36667,N_36803);
and U37870 (N_37870,N_36435,N_36437);
or U37871 (N_37871,N_36866,N_36204);
nand U37872 (N_37872,N_36014,N_36311);
or U37873 (N_37873,N_36406,N_36870);
xnor U37874 (N_37874,N_36001,N_36199);
or U37875 (N_37875,N_36642,N_36939);
or U37876 (N_37876,N_36226,N_36175);
and U37877 (N_37877,N_36060,N_36168);
nor U37878 (N_37878,N_36156,N_36355);
nor U37879 (N_37879,N_36983,N_36035);
nand U37880 (N_37880,N_36845,N_36637);
nor U37881 (N_37881,N_36976,N_36286);
nand U37882 (N_37882,N_36915,N_36895);
xor U37883 (N_37883,N_36071,N_36525);
nor U37884 (N_37884,N_36281,N_36262);
xnor U37885 (N_37885,N_36645,N_36762);
or U37886 (N_37886,N_36502,N_36730);
or U37887 (N_37887,N_36461,N_36613);
or U37888 (N_37888,N_36308,N_36837);
nand U37889 (N_37889,N_36727,N_36662);
nand U37890 (N_37890,N_36294,N_36911);
nor U37891 (N_37891,N_36151,N_36988);
xnor U37892 (N_37892,N_36402,N_36897);
xor U37893 (N_37893,N_36767,N_36140);
xnor U37894 (N_37894,N_36690,N_36048);
nor U37895 (N_37895,N_36369,N_36436);
nand U37896 (N_37896,N_36980,N_36098);
nand U37897 (N_37897,N_36109,N_36701);
nor U37898 (N_37898,N_36584,N_36777);
xnor U37899 (N_37899,N_36690,N_36677);
or U37900 (N_37900,N_36591,N_36410);
and U37901 (N_37901,N_36394,N_36113);
nor U37902 (N_37902,N_36001,N_36108);
nand U37903 (N_37903,N_36196,N_36186);
or U37904 (N_37904,N_36728,N_36230);
and U37905 (N_37905,N_36556,N_36512);
nand U37906 (N_37906,N_36597,N_36749);
nand U37907 (N_37907,N_36997,N_36731);
xor U37908 (N_37908,N_36560,N_36062);
xnor U37909 (N_37909,N_36545,N_36218);
or U37910 (N_37910,N_36082,N_36890);
nor U37911 (N_37911,N_36928,N_36360);
nor U37912 (N_37912,N_36630,N_36380);
nor U37913 (N_37913,N_36773,N_36537);
and U37914 (N_37914,N_36953,N_36939);
nand U37915 (N_37915,N_36376,N_36794);
and U37916 (N_37916,N_36166,N_36372);
nor U37917 (N_37917,N_36760,N_36772);
or U37918 (N_37918,N_36419,N_36107);
nor U37919 (N_37919,N_36889,N_36550);
nor U37920 (N_37920,N_36801,N_36899);
or U37921 (N_37921,N_36454,N_36992);
xor U37922 (N_37922,N_36765,N_36518);
nor U37923 (N_37923,N_36797,N_36531);
and U37924 (N_37924,N_36143,N_36203);
xnor U37925 (N_37925,N_36569,N_36410);
and U37926 (N_37926,N_36210,N_36080);
nand U37927 (N_37927,N_36271,N_36623);
and U37928 (N_37928,N_36017,N_36055);
xnor U37929 (N_37929,N_36506,N_36381);
or U37930 (N_37930,N_36176,N_36703);
and U37931 (N_37931,N_36570,N_36324);
nor U37932 (N_37932,N_36261,N_36911);
or U37933 (N_37933,N_36868,N_36257);
nor U37934 (N_37934,N_36371,N_36670);
or U37935 (N_37935,N_36284,N_36880);
and U37936 (N_37936,N_36600,N_36111);
or U37937 (N_37937,N_36820,N_36114);
nand U37938 (N_37938,N_36385,N_36585);
or U37939 (N_37939,N_36036,N_36920);
nand U37940 (N_37940,N_36148,N_36746);
nand U37941 (N_37941,N_36088,N_36655);
nand U37942 (N_37942,N_36108,N_36493);
nor U37943 (N_37943,N_36442,N_36724);
nand U37944 (N_37944,N_36577,N_36247);
or U37945 (N_37945,N_36602,N_36903);
and U37946 (N_37946,N_36829,N_36434);
xnor U37947 (N_37947,N_36119,N_36175);
or U37948 (N_37948,N_36810,N_36475);
xor U37949 (N_37949,N_36657,N_36358);
or U37950 (N_37950,N_36278,N_36299);
nand U37951 (N_37951,N_36960,N_36789);
xnor U37952 (N_37952,N_36454,N_36837);
nand U37953 (N_37953,N_36614,N_36181);
xnor U37954 (N_37954,N_36233,N_36984);
or U37955 (N_37955,N_36965,N_36986);
nor U37956 (N_37956,N_36444,N_36251);
and U37957 (N_37957,N_36251,N_36591);
nand U37958 (N_37958,N_36833,N_36068);
and U37959 (N_37959,N_36704,N_36846);
or U37960 (N_37960,N_36828,N_36423);
nor U37961 (N_37961,N_36876,N_36617);
and U37962 (N_37962,N_36581,N_36142);
xor U37963 (N_37963,N_36999,N_36629);
nand U37964 (N_37964,N_36582,N_36845);
or U37965 (N_37965,N_36452,N_36811);
and U37966 (N_37966,N_36218,N_36415);
nor U37967 (N_37967,N_36318,N_36172);
nand U37968 (N_37968,N_36186,N_36810);
nand U37969 (N_37969,N_36675,N_36726);
xnor U37970 (N_37970,N_36265,N_36689);
nor U37971 (N_37971,N_36685,N_36546);
and U37972 (N_37972,N_36672,N_36770);
nor U37973 (N_37973,N_36493,N_36383);
nor U37974 (N_37974,N_36213,N_36622);
nor U37975 (N_37975,N_36474,N_36905);
xor U37976 (N_37976,N_36226,N_36334);
xor U37977 (N_37977,N_36532,N_36766);
and U37978 (N_37978,N_36095,N_36331);
nand U37979 (N_37979,N_36186,N_36072);
and U37980 (N_37980,N_36925,N_36147);
or U37981 (N_37981,N_36322,N_36316);
xor U37982 (N_37982,N_36011,N_36265);
nand U37983 (N_37983,N_36417,N_36306);
and U37984 (N_37984,N_36401,N_36621);
xnor U37985 (N_37985,N_36618,N_36396);
and U37986 (N_37986,N_36505,N_36444);
xor U37987 (N_37987,N_36754,N_36577);
and U37988 (N_37988,N_36921,N_36504);
xor U37989 (N_37989,N_36667,N_36733);
or U37990 (N_37990,N_36657,N_36922);
and U37991 (N_37991,N_36586,N_36751);
and U37992 (N_37992,N_36242,N_36976);
and U37993 (N_37993,N_36456,N_36834);
and U37994 (N_37994,N_36803,N_36635);
xor U37995 (N_37995,N_36226,N_36237);
nor U37996 (N_37996,N_36749,N_36731);
or U37997 (N_37997,N_36990,N_36940);
nor U37998 (N_37998,N_36135,N_36615);
nor U37999 (N_37999,N_36683,N_36737);
nand U38000 (N_38000,N_37048,N_37909);
nor U38001 (N_38001,N_37780,N_37747);
nand U38002 (N_38002,N_37585,N_37673);
xor U38003 (N_38003,N_37569,N_37173);
or U38004 (N_38004,N_37665,N_37940);
xor U38005 (N_38005,N_37584,N_37148);
xnor U38006 (N_38006,N_37034,N_37582);
and U38007 (N_38007,N_37746,N_37031);
xnor U38008 (N_38008,N_37768,N_37513);
xnor U38009 (N_38009,N_37955,N_37177);
or U38010 (N_38010,N_37938,N_37823);
nor U38011 (N_38011,N_37033,N_37784);
or U38012 (N_38012,N_37325,N_37101);
nand U38013 (N_38013,N_37680,N_37056);
nand U38014 (N_38014,N_37450,N_37442);
or U38015 (N_38015,N_37428,N_37861);
and U38016 (N_38016,N_37926,N_37968);
or U38017 (N_38017,N_37947,N_37443);
nor U38018 (N_38018,N_37290,N_37781);
nor U38019 (N_38019,N_37255,N_37846);
or U38020 (N_38020,N_37820,N_37767);
and U38021 (N_38021,N_37748,N_37608);
xnor U38022 (N_38022,N_37294,N_37418);
or U38023 (N_38023,N_37809,N_37581);
nand U38024 (N_38024,N_37156,N_37166);
nor U38025 (N_38025,N_37514,N_37457);
xor U38026 (N_38026,N_37007,N_37424);
nor U38027 (N_38027,N_37738,N_37099);
nand U38028 (N_38028,N_37745,N_37228);
xnor U38029 (N_38029,N_37601,N_37465);
xor U38030 (N_38030,N_37836,N_37990);
or U38031 (N_38031,N_37089,N_37610);
nor U38032 (N_38032,N_37519,N_37261);
and U38033 (N_38033,N_37291,N_37460);
nand U38034 (N_38034,N_37941,N_37005);
or U38035 (N_38035,N_37184,N_37198);
and U38036 (N_38036,N_37924,N_37688);
nand U38037 (N_38037,N_37699,N_37501);
nand U38038 (N_38038,N_37730,N_37412);
or U38039 (N_38039,N_37435,N_37835);
nand U38040 (N_38040,N_37329,N_37049);
or U38041 (N_38041,N_37890,N_37201);
xor U38042 (N_38042,N_37011,N_37073);
nand U38043 (N_38043,N_37838,N_37051);
nor U38044 (N_38044,N_37399,N_37742);
nor U38045 (N_38045,N_37119,N_37496);
or U38046 (N_38046,N_37144,N_37625);
nor U38047 (N_38047,N_37817,N_37623);
or U38048 (N_38048,N_37227,N_37546);
and U38049 (N_38049,N_37619,N_37044);
xor U38050 (N_38050,N_37652,N_37620);
nor U38051 (N_38051,N_37196,N_37893);
and U38052 (N_38052,N_37664,N_37984);
and U38053 (N_38053,N_37221,N_37895);
or U38054 (N_38054,N_37482,N_37571);
or U38055 (N_38055,N_37818,N_37212);
nor U38056 (N_38056,N_37320,N_37347);
or U38057 (N_38057,N_37954,N_37485);
and U38058 (N_38058,N_37777,N_37628);
or U38059 (N_38059,N_37392,N_37908);
and U38060 (N_38060,N_37563,N_37591);
nor U38061 (N_38061,N_37481,N_37607);
and U38062 (N_38062,N_37466,N_37650);
xnor U38063 (N_38063,N_37093,N_37606);
or U38064 (N_38064,N_37552,N_37339);
or U38065 (N_38065,N_37079,N_37512);
nand U38066 (N_38066,N_37026,N_37264);
xor U38067 (N_38067,N_37503,N_37659);
or U38068 (N_38068,N_37561,N_37540);
nand U38069 (N_38069,N_37476,N_37276);
nor U38070 (N_38070,N_37704,N_37896);
or U38071 (N_38071,N_37082,N_37762);
or U38072 (N_38072,N_37899,N_37120);
and U38073 (N_38073,N_37888,N_37824);
nand U38074 (N_38074,N_37524,N_37728);
xor U38075 (N_38075,N_37195,N_37914);
nor U38076 (N_38076,N_37475,N_37700);
nand U38077 (N_38077,N_37213,N_37553);
or U38078 (N_38078,N_37887,N_37870);
nor U38079 (N_38079,N_37641,N_37133);
nor U38080 (N_38080,N_37779,N_37168);
and U38081 (N_38081,N_37431,N_37358);
nand U38082 (N_38082,N_37722,N_37630);
nor U38083 (N_38083,N_37706,N_37050);
and U38084 (N_38084,N_37451,N_37361);
nor U38085 (N_38085,N_37074,N_37637);
nand U38086 (N_38086,N_37542,N_37796);
nand U38087 (N_38087,N_37045,N_37807);
nor U38088 (N_38088,N_37520,N_37592);
and U38089 (N_38089,N_37406,N_37530);
nor U38090 (N_38090,N_37225,N_37911);
nand U38091 (N_38091,N_37903,N_37865);
and U38092 (N_38092,N_37981,N_37313);
and U38093 (N_38093,N_37676,N_37245);
or U38094 (N_38094,N_37386,N_37725);
xor U38095 (N_38095,N_37384,N_37960);
or U38096 (N_38096,N_37223,N_37681);
and U38097 (N_38097,N_37980,N_37712);
nand U38098 (N_38098,N_37041,N_37701);
nand U38099 (N_38099,N_37373,N_37178);
nand U38100 (N_38100,N_37027,N_37066);
and U38101 (N_38101,N_37497,N_37928);
xnor U38102 (N_38102,N_37653,N_37535);
and U38103 (N_38103,N_37516,N_37522);
nand U38104 (N_38104,N_37236,N_37898);
or U38105 (N_38105,N_37965,N_37310);
xor U38106 (N_38106,N_37544,N_37023);
and U38107 (N_38107,N_37539,N_37910);
nor U38108 (N_38108,N_37731,N_37797);
or U38109 (N_38109,N_37932,N_37463);
nor U38110 (N_38110,N_37370,N_37286);
or U38111 (N_38111,N_37420,N_37137);
xor U38112 (N_38112,N_37233,N_37977);
nor U38113 (N_38113,N_37032,N_37438);
xnor U38114 (N_38114,N_37307,N_37122);
nor U38115 (N_38115,N_37285,N_37398);
or U38116 (N_38116,N_37827,N_37832);
nor U38117 (N_38117,N_37489,N_37010);
and U38118 (N_38118,N_37423,N_37504);
nand U38119 (N_38119,N_37165,N_37246);
nand U38120 (N_38120,N_37235,N_37605);
xor U38121 (N_38121,N_37739,N_37091);
xor U38122 (N_38122,N_37483,N_37115);
xor U38123 (N_38123,N_37595,N_37309);
nor U38124 (N_38124,N_37287,N_37356);
or U38125 (N_38125,N_37508,N_37249);
and U38126 (N_38126,N_37426,N_37421);
and U38127 (N_38127,N_37929,N_37543);
or U38128 (N_38128,N_37621,N_37464);
nand U38129 (N_38129,N_37643,N_37318);
nand U38130 (N_38130,N_37867,N_37943);
and U38131 (N_38131,N_37743,N_37182);
and U38132 (N_38132,N_37258,N_37646);
nor U38133 (N_38133,N_37132,N_37845);
nand U38134 (N_38134,N_37814,N_37492);
nor U38135 (N_38135,N_37828,N_37289);
nor U38136 (N_38136,N_37169,N_37247);
or U38137 (N_38137,N_37203,N_37798);
nand U38138 (N_38138,N_37877,N_37445);
or U38139 (N_38139,N_37729,N_37419);
nor U38140 (N_38140,N_37302,N_37717);
xnor U38141 (N_38141,N_37087,N_37234);
nand U38142 (N_38142,N_37439,N_37568);
or U38143 (N_38143,N_37557,N_37025);
nand U38144 (N_38144,N_37755,N_37979);
xnor U38145 (N_38145,N_37176,N_37047);
xor U38146 (N_38146,N_37971,N_37869);
and U38147 (N_38147,N_37856,N_37266);
nor U38148 (N_38148,N_37657,N_37952);
or U38149 (N_38149,N_37715,N_37632);
or U38150 (N_38150,N_37912,N_37660);
nor U38151 (N_38151,N_37348,N_37305);
and U38152 (N_38152,N_37702,N_37364);
nand U38153 (N_38153,N_37855,N_37936);
nor U38154 (N_38154,N_37672,N_37456);
or U38155 (N_38155,N_37674,N_37337);
xor U38156 (N_38156,N_37080,N_37905);
nand U38157 (N_38157,N_37160,N_37826);
xor U38158 (N_38158,N_37545,N_37787);
nor U38159 (N_38159,N_37976,N_37024);
xor U38160 (N_38160,N_37612,N_37517);
or U38161 (N_38161,N_37062,N_37139);
nor U38162 (N_38162,N_37242,N_37933);
nand U38163 (N_38163,N_37411,N_37864);
and U38164 (N_38164,N_37920,N_37945);
and U38165 (N_38165,N_37243,N_37316);
nor U38166 (N_38166,N_37494,N_37271);
or U38167 (N_38167,N_37344,N_37939);
and U38168 (N_38168,N_37415,N_37015);
and U38169 (N_38169,N_37351,N_37470);
and U38170 (N_38170,N_37171,N_37417);
nor U38171 (N_38171,N_37360,N_37224);
or U38172 (N_38172,N_37559,N_37104);
xnor U38173 (N_38173,N_37505,N_37741);
nor U38174 (N_38174,N_37782,N_37799);
and U38175 (N_38175,N_37596,N_37837);
nand U38176 (N_38176,N_37829,N_37786);
nand U38177 (N_38177,N_37863,N_37991);
or U38178 (N_38178,N_37640,N_37487);
nor U38179 (N_38179,N_37330,N_37972);
nand U38180 (N_38180,N_37437,N_37108);
xnor U38181 (N_38181,N_37379,N_37397);
and U38182 (N_38182,N_37292,N_37052);
nor U38183 (N_38183,N_37409,N_37434);
nand U38184 (N_38184,N_37352,N_37030);
nand U38185 (N_38185,N_37669,N_37523);
nand U38186 (N_38186,N_37574,N_37978);
and U38187 (N_38187,N_37687,N_37500);
and U38188 (N_38188,N_37155,N_37854);
nand U38189 (N_38189,N_37927,N_37883);
nand U38190 (N_38190,N_37538,N_37121);
xnor U38191 (N_38191,N_37484,N_37260);
xor U38192 (N_38192,N_37711,N_37140);
xnor U38193 (N_38193,N_37708,N_37381);
nor U38194 (N_38194,N_37693,N_37983);
xor U38195 (N_38195,N_37844,N_37562);
nand U38196 (N_38196,N_37805,N_37105);
xor U38197 (N_38197,N_37486,N_37935);
nor U38198 (N_38198,N_37554,N_37853);
nand U38199 (N_38199,N_37186,N_37147);
nand U38200 (N_38200,N_37884,N_37713);
xor U38201 (N_38201,N_37547,N_37267);
and U38202 (N_38202,N_37342,N_37686);
nand U38203 (N_38203,N_37436,N_37962);
nand U38204 (N_38204,N_37858,N_37875);
nor U38205 (N_38205,N_37192,N_37609);
nor U38206 (N_38206,N_37020,N_37006);
nor U38207 (N_38207,N_37263,N_37259);
xnor U38208 (N_38208,N_37391,N_37937);
nor U38209 (N_38209,N_37944,N_37493);
nand U38210 (N_38210,N_37314,N_37262);
xor U38211 (N_38211,N_37449,N_37859);
xnor U38212 (N_38212,N_37705,N_37036);
nor U38213 (N_38213,N_37792,N_37548);
nand U38214 (N_38214,N_37997,N_37885);
and U38215 (N_38215,N_37577,N_37847);
or U38216 (N_38216,N_37275,N_37063);
xnor U38217 (N_38217,N_37014,N_37226);
and U38218 (N_38218,N_37901,N_37580);
nand U38219 (N_38219,N_37998,N_37124);
or U38220 (N_38220,N_37282,N_37793);
xor U38221 (N_38221,N_37841,N_37382);
xnor U38222 (N_38222,N_37112,N_37461);
xnor U38223 (N_38223,N_37679,N_37753);
nor U38224 (N_38224,N_37194,N_37405);
and U38225 (N_38225,N_37018,N_37872);
nor U38226 (N_38226,N_37001,N_37532);
or U38227 (N_38227,N_37422,N_37103);
nand U38228 (N_38228,N_37130,N_37058);
nor U38229 (N_38229,N_37187,N_37413);
and U38230 (N_38230,N_37776,N_37788);
or U38231 (N_38231,N_37537,N_37756);
nand U38232 (N_38232,N_37970,N_37648);
and U38233 (N_38233,N_37240,N_37951);
nand U38234 (N_38234,N_37380,N_37340);
and U38235 (N_38235,N_37749,N_37474);
and U38236 (N_38236,N_37878,N_37447);
or U38237 (N_38237,N_37076,N_37802);
and U38238 (N_38238,N_37279,N_37525);
nand U38239 (N_38239,N_37118,N_37327);
nand U38240 (N_38240,N_37662,N_37175);
nand U38241 (N_38241,N_37953,N_37973);
nor U38242 (N_38242,N_37215,N_37061);
nor U38243 (N_38243,N_37404,N_37647);
or U38244 (N_38244,N_37737,N_37136);
or U38245 (N_38245,N_37987,N_37667);
xor U38246 (N_38246,N_37304,N_37219);
nand U38247 (N_38247,N_37598,N_37432);
nor U38248 (N_38248,N_37860,N_37490);
nand U38249 (N_38249,N_37216,N_37257);
nor U38250 (N_38250,N_37511,N_37763);
and U38251 (N_38251,N_37495,N_37238);
nor U38252 (N_38252,N_37934,N_37232);
xor U38253 (N_38253,N_37624,N_37770);
xor U38254 (N_38254,N_37328,N_37663);
xnor U38255 (N_38255,N_37760,N_37677);
xnor U38256 (N_38256,N_37989,N_37038);
nand U38257 (N_38257,N_37440,N_37109);
xor U38258 (N_38258,N_37564,N_37346);
nor U38259 (N_38259,N_37149,N_37281);
xnor U38260 (N_38260,N_37848,N_37622);
and U38261 (N_38261,N_37761,N_37866);
and U38262 (N_38262,N_37882,N_37879);
and U38263 (N_38263,N_37323,N_37253);
xnor U38264 (N_38264,N_37586,N_37773);
nand U38265 (N_38265,N_37521,N_37654);
xor U38266 (N_38266,N_37956,N_37849);
nor U38267 (N_38267,N_37509,N_37315);
or U38268 (N_38268,N_37806,N_37452);
xnor U38269 (N_38269,N_37433,N_37857);
nor U38270 (N_38270,N_37682,N_37515);
xnor U38271 (N_38271,N_37106,N_37021);
xor U38272 (N_38272,N_37724,N_37576);
nor U38273 (N_38273,N_37597,N_37146);
or U38274 (N_38274,N_37698,N_37174);
or U38275 (N_38275,N_37454,N_37181);
xnor U38276 (N_38276,N_37573,N_37754);
and U38277 (N_38277,N_37029,N_37635);
xor U38278 (N_38278,N_37387,N_37723);
nor U38279 (N_38279,N_37634,N_37239);
nor U38280 (N_38280,N_37090,N_37649);
xor U38281 (N_38281,N_37371,N_37685);
xor U38282 (N_38282,N_37958,N_37378);
or U38283 (N_38283,N_37949,N_37039);
nand U38284 (N_38284,N_37689,N_37163);
and U38285 (N_38285,N_37459,N_37959);
or U38286 (N_38286,N_37800,N_37308);
nand U38287 (N_38287,N_37915,N_37558);
nor U38288 (N_38288,N_37331,N_37046);
nor U38289 (N_38289,N_37498,N_37188);
xnor U38290 (N_38290,N_37094,N_37992);
nand U38291 (N_38291,N_37639,N_37744);
xnor U38292 (N_38292,N_37300,N_37129);
or U38293 (N_38293,N_37009,N_37771);
nand U38294 (N_38294,N_37593,N_37319);
or U38295 (N_38295,N_37790,N_37207);
xnor U38296 (N_38296,N_37288,N_37072);
or U38297 (N_38297,N_37556,N_37566);
xnor U38298 (N_38298,N_37812,N_37703);
or U38299 (N_38299,N_37277,N_37871);
and U38300 (N_38300,N_37611,N_37349);
and U38301 (N_38301,N_37343,N_37335);
or U38302 (N_38302,N_37059,N_37468);
or U38303 (N_38303,N_37633,N_37283);
and U38304 (N_38304,N_37078,N_37057);
nand U38305 (N_38305,N_37734,N_37727);
and U38306 (N_38306,N_37528,N_37720);
and U38307 (N_38307,N_37167,N_37684);
and U38308 (N_38308,N_37158,N_37037);
nand U38309 (N_38309,N_37617,N_37154);
or U38310 (N_38310,N_37383,N_37907);
xor U38311 (N_38311,N_37230,N_37317);
xor U38312 (N_38312,N_37394,N_37638);
and U38313 (N_38313,N_37205,N_37054);
nor U38314 (N_38314,N_37804,N_37472);
xnor U38315 (N_38315,N_37819,N_37811);
xor U38316 (N_38316,N_37709,N_37111);
xor U38317 (N_38317,N_37060,N_37265);
or U38318 (N_38318,N_37092,N_37345);
xor U38319 (N_38319,N_37202,N_37833);
or U38320 (N_38320,N_37488,N_37683);
xnor U38321 (N_38321,N_37085,N_37840);
nand U38322 (N_38322,N_37778,N_37506);
and U38323 (N_38323,N_37003,N_37278);
nand U38324 (N_38324,N_37531,N_37691);
and U38325 (N_38325,N_37068,N_37839);
nor U38326 (N_38326,N_37975,N_37589);
nand U38327 (N_38327,N_37321,N_37813);
nand U38328 (N_38328,N_37107,N_37017);
and U38329 (N_38329,N_37028,N_37529);
and U38330 (N_38330,N_37134,N_37172);
xor U38331 (N_38331,N_37690,N_37471);
xnor U38332 (N_38332,N_37229,N_37189);
or U38333 (N_38333,N_37374,N_37153);
or U38334 (N_38334,N_37390,N_37237);
nand U38335 (N_38335,N_37248,N_37661);
and U38336 (N_38336,N_37135,N_37668);
nor U38337 (N_38337,N_37455,N_37510);
nor U38338 (N_38338,N_37075,N_37388);
nand U38339 (N_38339,N_37268,N_37917);
xnor U38340 (N_38340,N_37332,N_37764);
xor U38341 (N_38341,N_37889,N_37395);
or U38342 (N_38342,N_37179,N_37270);
nor U38343 (N_38343,N_37064,N_37200);
nand U38344 (N_38344,N_37964,N_37241);
nor U38345 (N_38345,N_37923,N_37572);
xor U38346 (N_38346,N_37697,N_37272);
and U38347 (N_38347,N_37750,N_37735);
nor U38348 (N_38348,N_37206,N_37996);
and U38349 (N_38349,N_37694,N_37658);
and U38350 (N_38350,N_37575,N_37966);
and U38351 (N_38351,N_37894,N_37284);
or U38352 (N_38352,N_37312,N_37311);
or U38353 (N_38353,N_37170,N_37204);
and U38354 (N_38354,N_37982,N_37210);
nor U38355 (N_38355,N_37536,N_37324);
and U38356 (N_38356,N_37714,N_37217);
nor U38357 (N_38357,N_37102,N_37602);
and U38358 (N_38358,N_37053,N_37448);
and U38359 (N_38359,N_37393,N_37830);
xnor U38360 (N_38360,N_37906,N_37350);
or U38361 (N_38361,N_37385,N_37721);
xnor U38362 (N_38362,N_37042,N_37071);
nor U38363 (N_38363,N_37583,N_37301);
and U38364 (N_38364,N_37416,N_37043);
nor U38365 (N_38365,N_37815,N_37655);
nand U38366 (N_38366,N_37407,N_37834);
and U38367 (N_38367,N_37696,N_37353);
xnor U38368 (N_38368,N_37916,N_37098);
and U38369 (N_38369,N_37357,N_37218);
xor U38370 (N_38370,N_37222,N_37183);
nand U38371 (N_38371,N_37002,N_37618);
xnor U38372 (N_38372,N_37081,N_37362);
nand U38373 (N_38373,N_37113,N_37671);
nand U38374 (N_38374,N_37366,N_37083);
or U38375 (N_38375,N_37478,N_37019);
xnor U38376 (N_38376,N_37469,N_37891);
xor U38377 (N_38377,N_37719,N_37897);
nor U38378 (N_38378,N_37355,N_37921);
or U38379 (N_38379,N_37070,N_37603);
nand U38380 (N_38380,N_37613,N_37477);
and U38381 (N_38381,N_37040,N_37541);
nand U38382 (N_38382,N_37751,N_37000);
xnor U38383 (N_38383,N_37752,N_37180);
nor U38384 (N_38384,N_37097,N_37013);
or U38385 (N_38385,N_37789,N_37016);
nor U38386 (N_38386,N_37375,N_37651);
nor U38387 (N_38387,N_37502,N_37918);
xnor U38388 (N_38388,N_37892,N_37256);
and U38389 (N_38389,N_37930,N_37850);
nor U38390 (N_38390,N_37785,N_37604);
nand U38391 (N_38391,N_37069,N_37587);
xnor U38392 (N_38392,N_37772,N_37963);
xor U38393 (N_38393,N_37055,N_37533);
nand U38394 (N_38394,N_37142,N_37985);
nand U38395 (N_38395,N_37334,N_37376);
and U38396 (N_38396,N_37957,N_37220);
and U38397 (N_38397,N_37293,N_37244);
or U38398 (N_38398,N_37551,N_37969);
nand U38399 (N_38399,N_37822,N_37141);
nor U38400 (N_38400,N_37534,N_37273);
xnor U38401 (N_38401,N_37707,N_37759);
xor U38402 (N_38402,N_37280,N_37444);
or U38403 (N_38403,N_37151,N_37145);
and U38404 (N_38404,N_37902,N_37880);
nor U38405 (N_38405,N_37616,N_37128);
or U38406 (N_38406,N_37231,N_37303);
and U38407 (N_38407,N_37801,N_37088);
xnor U38408 (N_38408,N_37254,N_37862);
nand U38409 (N_38409,N_37567,N_37925);
nor U38410 (N_38410,N_37695,N_37666);
or U38411 (N_38411,N_37095,N_37816);
or U38412 (N_38412,N_37127,N_37004);
nor U38413 (N_38413,N_37948,N_37579);
or U38414 (N_38414,N_37758,N_37410);
and U38415 (N_38415,N_37157,N_37473);
nor U38416 (N_38416,N_37757,N_37636);
nand U38417 (N_38417,N_37900,N_37365);
or U38418 (N_38418,N_37794,N_37526);
or U38419 (N_38419,N_37499,N_37570);
xnor U38420 (N_38420,N_37994,N_37560);
nor U38421 (N_38421,N_37333,N_37678);
or U38422 (N_38422,N_37590,N_37765);
and U38423 (N_38423,N_37022,N_37555);
or U38424 (N_38424,N_37199,N_37250);
nor U38425 (N_38425,N_37100,N_37326);
or U38426 (N_38426,N_37527,N_37808);
nand U38427 (N_38427,N_37631,N_37831);
xnor U38428 (N_38428,N_37629,N_37297);
nor U38429 (N_38429,N_37642,N_37338);
xnor U38430 (N_38430,N_37726,N_37986);
nor U38431 (N_38431,N_37377,N_37931);
and U38432 (N_38432,N_37123,N_37775);
and U38433 (N_38433,N_37414,N_37550);
xnor U38434 (N_38434,N_37644,N_37269);
xnor U38435 (N_38435,N_37369,N_37067);
or U38436 (N_38436,N_37117,N_37065);
nand U38437 (N_38437,N_37851,N_37159);
xor U38438 (N_38438,N_37252,N_37791);
nor U38439 (N_38439,N_37209,N_37549);
nand U38440 (N_38440,N_37363,N_37408);
and U38441 (N_38441,N_37336,N_37656);
xnor U38442 (N_38442,N_37670,N_37675);
xor U38443 (N_38443,N_37578,N_37185);
or U38444 (N_38444,N_37084,N_37116);
and U38445 (N_38445,N_37402,N_37599);
nand U38446 (N_38446,N_37298,N_37874);
or U38447 (N_38447,N_37821,N_37008);
xor U38448 (N_38448,N_37359,N_37077);
and U38449 (N_38449,N_37732,N_37161);
nand U38450 (N_38450,N_37627,N_37467);
nor U38451 (N_38451,N_37150,N_37716);
nand U38452 (N_38452,N_37458,N_37096);
and U38453 (N_38453,N_37881,N_37740);
xnor U38454 (N_38454,N_37518,N_37427);
nor U38455 (N_38455,N_37479,N_37401);
nor U38456 (N_38456,N_37507,N_37453);
and U38457 (N_38457,N_37995,N_37852);
or U38458 (N_38458,N_37692,N_37446);
and U38459 (N_38459,N_37251,N_37367);
nand U38460 (N_38460,N_37086,N_37600);
xor U38461 (N_38461,N_37614,N_37211);
or U38462 (N_38462,N_37769,N_37718);
nand U38463 (N_38463,N_37368,N_37191);
and U38464 (N_38464,N_37946,N_37626);
nand U38465 (N_38465,N_37999,N_37143);
and U38466 (N_38466,N_37950,N_37162);
nor U38467 (N_38467,N_37299,N_37961);
or U38468 (N_38468,N_37110,N_37138);
or U38469 (N_38469,N_37403,N_37274);
and U38470 (N_38470,N_37429,N_37462);
or U38471 (N_38471,N_37783,N_37354);
xnor U38472 (N_38472,N_37868,N_37131);
xnor U38473 (N_38473,N_37197,N_37594);
and U38474 (N_38474,N_37967,N_37904);
nor U38475 (N_38475,N_37012,N_37441);
or U38476 (N_38476,N_37389,N_37766);
nor U38477 (N_38477,N_37341,N_37615);
nand U38478 (N_38478,N_37190,N_37193);
xor U38479 (N_38479,N_37396,N_37843);
xor U38480 (N_38480,N_37126,N_37825);
and U38481 (N_38481,N_37803,N_37208);
and U38482 (N_38482,N_37922,N_37774);
nor U38483 (N_38483,N_37919,N_37400);
nand U38484 (N_38484,N_37114,N_37565);
or U38485 (N_38485,N_37214,N_37913);
or U38486 (N_38486,N_37322,N_37152);
nand U38487 (N_38487,N_37873,N_37810);
or U38488 (N_38488,N_37988,N_37942);
xnor U38489 (N_38489,N_37736,N_37842);
xor U38490 (N_38490,N_37372,N_37993);
xnor U38491 (N_38491,N_37795,N_37974);
and U38492 (N_38492,N_37480,N_37491);
nand U38493 (N_38493,N_37886,N_37430);
nor U38494 (N_38494,N_37425,N_37295);
nand U38495 (N_38495,N_37125,N_37733);
and U38496 (N_38496,N_37035,N_37645);
and U38497 (N_38497,N_37588,N_37306);
nor U38498 (N_38498,N_37164,N_37710);
or U38499 (N_38499,N_37876,N_37296);
nand U38500 (N_38500,N_37022,N_37364);
nor U38501 (N_38501,N_37846,N_37406);
nor U38502 (N_38502,N_37258,N_37760);
xnor U38503 (N_38503,N_37018,N_37237);
nand U38504 (N_38504,N_37735,N_37616);
or U38505 (N_38505,N_37275,N_37367);
nand U38506 (N_38506,N_37005,N_37462);
nor U38507 (N_38507,N_37779,N_37135);
or U38508 (N_38508,N_37354,N_37156);
nand U38509 (N_38509,N_37387,N_37689);
nor U38510 (N_38510,N_37631,N_37899);
or U38511 (N_38511,N_37334,N_37415);
and U38512 (N_38512,N_37467,N_37036);
nor U38513 (N_38513,N_37195,N_37830);
xnor U38514 (N_38514,N_37180,N_37405);
or U38515 (N_38515,N_37326,N_37916);
or U38516 (N_38516,N_37676,N_37234);
nor U38517 (N_38517,N_37055,N_37081);
nand U38518 (N_38518,N_37848,N_37058);
or U38519 (N_38519,N_37641,N_37637);
nor U38520 (N_38520,N_37821,N_37761);
nor U38521 (N_38521,N_37070,N_37253);
xor U38522 (N_38522,N_37822,N_37025);
xor U38523 (N_38523,N_37180,N_37551);
nor U38524 (N_38524,N_37044,N_37466);
xnor U38525 (N_38525,N_37658,N_37003);
nand U38526 (N_38526,N_37245,N_37590);
nor U38527 (N_38527,N_37940,N_37503);
and U38528 (N_38528,N_37505,N_37742);
or U38529 (N_38529,N_37859,N_37556);
or U38530 (N_38530,N_37040,N_37158);
or U38531 (N_38531,N_37176,N_37208);
xnor U38532 (N_38532,N_37819,N_37726);
or U38533 (N_38533,N_37615,N_37538);
xor U38534 (N_38534,N_37708,N_37945);
xnor U38535 (N_38535,N_37132,N_37997);
nor U38536 (N_38536,N_37110,N_37900);
nor U38537 (N_38537,N_37713,N_37753);
nor U38538 (N_38538,N_37577,N_37694);
or U38539 (N_38539,N_37150,N_37958);
or U38540 (N_38540,N_37651,N_37738);
nor U38541 (N_38541,N_37557,N_37938);
nand U38542 (N_38542,N_37354,N_37866);
xor U38543 (N_38543,N_37897,N_37089);
xor U38544 (N_38544,N_37822,N_37557);
nor U38545 (N_38545,N_37011,N_37198);
nor U38546 (N_38546,N_37650,N_37172);
nor U38547 (N_38547,N_37570,N_37191);
nor U38548 (N_38548,N_37698,N_37936);
nor U38549 (N_38549,N_37506,N_37189);
xnor U38550 (N_38550,N_37445,N_37864);
xor U38551 (N_38551,N_37939,N_37605);
and U38552 (N_38552,N_37918,N_37167);
xnor U38553 (N_38553,N_37403,N_37940);
and U38554 (N_38554,N_37078,N_37652);
nor U38555 (N_38555,N_37636,N_37206);
and U38556 (N_38556,N_37162,N_37396);
and U38557 (N_38557,N_37708,N_37723);
or U38558 (N_38558,N_37087,N_37883);
and U38559 (N_38559,N_37840,N_37688);
or U38560 (N_38560,N_37103,N_37932);
xnor U38561 (N_38561,N_37792,N_37322);
or U38562 (N_38562,N_37675,N_37647);
nor U38563 (N_38563,N_37200,N_37053);
nor U38564 (N_38564,N_37196,N_37294);
xnor U38565 (N_38565,N_37786,N_37254);
nor U38566 (N_38566,N_37956,N_37498);
and U38567 (N_38567,N_37965,N_37162);
nor U38568 (N_38568,N_37740,N_37903);
or U38569 (N_38569,N_37732,N_37914);
or U38570 (N_38570,N_37495,N_37096);
nor U38571 (N_38571,N_37888,N_37518);
nand U38572 (N_38572,N_37182,N_37357);
nor U38573 (N_38573,N_37669,N_37522);
nand U38574 (N_38574,N_37091,N_37423);
nand U38575 (N_38575,N_37476,N_37865);
and U38576 (N_38576,N_37482,N_37612);
or U38577 (N_38577,N_37385,N_37672);
or U38578 (N_38578,N_37610,N_37098);
xor U38579 (N_38579,N_37229,N_37202);
and U38580 (N_38580,N_37990,N_37027);
nand U38581 (N_38581,N_37310,N_37020);
or U38582 (N_38582,N_37142,N_37496);
xor U38583 (N_38583,N_37678,N_37708);
nand U38584 (N_38584,N_37384,N_37262);
nor U38585 (N_38585,N_37906,N_37022);
or U38586 (N_38586,N_37510,N_37119);
and U38587 (N_38587,N_37783,N_37217);
and U38588 (N_38588,N_37077,N_37796);
or U38589 (N_38589,N_37702,N_37128);
nor U38590 (N_38590,N_37507,N_37514);
and U38591 (N_38591,N_37712,N_37895);
nand U38592 (N_38592,N_37178,N_37830);
and U38593 (N_38593,N_37167,N_37185);
xor U38594 (N_38594,N_37043,N_37277);
xor U38595 (N_38595,N_37647,N_37738);
or U38596 (N_38596,N_37447,N_37709);
nand U38597 (N_38597,N_37947,N_37294);
or U38598 (N_38598,N_37431,N_37766);
and U38599 (N_38599,N_37236,N_37464);
or U38600 (N_38600,N_37203,N_37622);
or U38601 (N_38601,N_37460,N_37051);
nand U38602 (N_38602,N_37221,N_37410);
xnor U38603 (N_38603,N_37104,N_37266);
or U38604 (N_38604,N_37864,N_37104);
nand U38605 (N_38605,N_37726,N_37319);
xor U38606 (N_38606,N_37936,N_37841);
and U38607 (N_38607,N_37115,N_37078);
nand U38608 (N_38608,N_37741,N_37041);
or U38609 (N_38609,N_37502,N_37269);
nand U38610 (N_38610,N_37308,N_37090);
or U38611 (N_38611,N_37937,N_37599);
nand U38612 (N_38612,N_37114,N_37193);
nor U38613 (N_38613,N_37809,N_37447);
and U38614 (N_38614,N_37419,N_37034);
and U38615 (N_38615,N_37445,N_37964);
nand U38616 (N_38616,N_37151,N_37793);
nor U38617 (N_38617,N_37869,N_37617);
nor U38618 (N_38618,N_37575,N_37225);
xor U38619 (N_38619,N_37229,N_37713);
and U38620 (N_38620,N_37744,N_37368);
or U38621 (N_38621,N_37649,N_37010);
or U38622 (N_38622,N_37191,N_37654);
or U38623 (N_38623,N_37456,N_37642);
nor U38624 (N_38624,N_37589,N_37959);
nand U38625 (N_38625,N_37388,N_37096);
nand U38626 (N_38626,N_37643,N_37435);
and U38627 (N_38627,N_37859,N_37710);
and U38628 (N_38628,N_37281,N_37796);
or U38629 (N_38629,N_37093,N_37335);
and U38630 (N_38630,N_37130,N_37637);
nor U38631 (N_38631,N_37957,N_37231);
nand U38632 (N_38632,N_37083,N_37730);
or U38633 (N_38633,N_37117,N_37836);
nor U38634 (N_38634,N_37036,N_37309);
xor U38635 (N_38635,N_37342,N_37467);
nand U38636 (N_38636,N_37681,N_37869);
or U38637 (N_38637,N_37407,N_37822);
nand U38638 (N_38638,N_37760,N_37916);
xnor U38639 (N_38639,N_37692,N_37442);
nor U38640 (N_38640,N_37459,N_37287);
nand U38641 (N_38641,N_37448,N_37812);
nand U38642 (N_38642,N_37664,N_37231);
and U38643 (N_38643,N_37090,N_37458);
or U38644 (N_38644,N_37587,N_37055);
xor U38645 (N_38645,N_37527,N_37083);
or U38646 (N_38646,N_37336,N_37597);
nand U38647 (N_38647,N_37376,N_37011);
nor U38648 (N_38648,N_37731,N_37900);
xnor U38649 (N_38649,N_37041,N_37100);
and U38650 (N_38650,N_37881,N_37835);
and U38651 (N_38651,N_37187,N_37730);
and U38652 (N_38652,N_37129,N_37392);
or U38653 (N_38653,N_37753,N_37532);
or U38654 (N_38654,N_37801,N_37993);
xnor U38655 (N_38655,N_37660,N_37262);
nor U38656 (N_38656,N_37673,N_37538);
xor U38657 (N_38657,N_37049,N_37442);
nor U38658 (N_38658,N_37386,N_37073);
nor U38659 (N_38659,N_37722,N_37362);
and U38660 (N_38660,N_37719,N_37798);
nand U38661 (N_38661,N_37137,N_37656);
or U38662 (N_38662,N_37722,N_37191);
nand U38663 (N_38663,N_37312,N_37925);
xor U38664 (N_38664,N_37660,N_37359);
and U38665 (N_38665,N_37302,N_37264);
or U38666 (N_38666,N_37174,N_37664);
and U38667 (N_38667,N_37340,N_37351);
xor U38668 (N_38668,N_37759,N_37528);
xnor U38669 (N_38669,N_37335,N_37188);
nand U38670 (N_38670,N_37093,N_37815);
nor U38671 (N_38671,N_37955,N_37354);
nor U38672 (N_38672,N_37245,N_37824);
nor U38673 (N_38673,N_37109,N_37415);
xnor U38674 (N_38674,N_37573,N_37955);
and U38675 (N_38675,N_37762,N_37990);
or U38676 (N_38676,N_37236,N_37137);
and U38677 (N_38677,N_37061,N_37025);
nand U38678 (N_38678,N_37422,N_37388);
or U38679 (N_38679,N_37082,N_37170);
nor U38680 (N_38680,N_37585,N_37767);
nor U38681 (N_38681,N_37345,N_37656);
nand U38682 (N_38682,N_37696,N_37316);
nand U38683 (N_38683,N_37423,N_37096);
and U38684 (N_38684,N_37381,N_37295);
nand U38685 (N_38685,N_37391,N_37627);
xnor U38686 (N_38686,N_37433,N_37885);
nand U38687 (N_38687,N_37024,N_37141);
nand U38688 (N_38688,N_37503,N_37476);
and U38689 (N_38689,N_37748,N_37960);
nand U38690 (N_38690,N_37906,N_37909);
nor U38691 (N_38691,N_37008,N_37789);
nor U38692 (N_38692,N_37094,N_37734);
nand U38693 (N_38693,N_37875,N_37273);
nor U38694 (N_38694,N_37663,N_37076);
xor U38695 (N_38695,N_37936,N_37800);
xnor U38696 (N_38696,N_37692,N_37638);
and U38697 (N_38697,N_37159,N_37100);
nor U38698 (N_38698,N_37407,N_37153);
xnor U38699 (N_38699,N_37124,N_37373);
nor U38700 (N_38700,N_37058,N_37858);
nor U38701 (N_38701,N_37506,N_37085);
nor U38702 (N_38702,N_37483,N_37290);
nand U38703 (N_38703,N_37072,N_37758);
and U38704 (N_38704,N_37236,N_37421);
or U38705 (N_38705,N_37613,N_37150);
xnor U38706 (N_38706,N_37480,N_37945);
xor U38707 (N_38707,N_37298,N_37569);
xor U38708 (N_38708,N_37125,N_37908);
xor U38709 (N_38709,N_37363,N_37809);
nor U38710 (N_38710,N_37271,N_37809);
and U38711 (N_38711,N_37211,N_37372);
and U38712 (N_38712,N_37549,N_37760);
xor U38713 (N_38713,N_37187,N_37741);
and U38714 (N_38714,N_37131,N_37217);
xnor U38715 (N_38715,N_37613,N_37209);
nand U38716 (N_38716,N_37216,N_37669);
and U38717 (N_38717,N_37917,N_37790);
or U38718 (N_38718,N_37812,N_37697);
nor U38719 (N_38719,N_37911,N_37703);
nand U38720 (N_38720,N_37024,N_37148);
nor U38721 (N_38721,N_37475,N_37449);
and U38722 (N_38722,N_37681,N_37246);
and U38723 (N_38723,N_37945,N_37873);
or U38724 (N_38724,N_37764,N_37195);
nor U38725 (N_38725,N_37360,N_37430);
xor U38726 (N_38726,N_37317,N_37060);
or U38727 (N_38727,N_37147,N_37784);
and U38728 (N_38728,N_37780,N_37050);
or U38729 (N_38729,N_37508,N_37369);
or U38730 (N_38730,N_37742,N_37991);
xnor U38731 (N_38731,N_37964,N_37003);
nand U38732 (N_38732,N_37102,N_37171);
nand U38733 (N_38733,N_37710,N_37626);
nor U38734 (N_38734,N_37107,N_37751);
and U38735 (N_38735,N_37290,N_37285);
and U38736 (N_38736,N_37240,N_37051);
or U38737 (N_38737,N_37004,N_37126);
or U38738 (N_38738,N_37005,N_37514);
or U38739 (N_38739,N_37928,N_37277);
or U38740 (N_38740,N_37323,N_37733);
nand U38741 (N_38741,N_37813,N_37766);
xor U38742 (N_38742,N_37622,N_37553);
and U38743 (N_38743,N_37574,N_37473);
and U38744 (N_38744,N_37493,N_37574);
or U38745 (N_38745,N_37319,N_37831);
xnor U38746 (N_38746,N_37929,N_37159);
or U38747 (N_38747,N_37108,N_37632);
nand U38748 (N_38748,N_37408,N_37594);
nor U38749 (N_38749,N_37034,N_37200);
or U38750 (N_38750,N_37811,N_37387);
or U38751 (N_38751,N_37748,N_37115);
or U38752 (N_38752,N_37827,N_37079);
and U38753 (N_38753,N_37146,N_37868);
or U38754 (N_38754,N_37477,N_37775);
xnor U38755 (N_38755,N_37950,N_37679);
xnor U38756 (N_38756,N_37270,N_37305);
and U38757 (N_38757,N_37117,N_37802);
xnor U38758 (N_38758,N_37154,N_37328);
or U38759 (N_38759,N_37921,N_37123);
or U38760 (N_38760,N_37063,N_37121);
xor U38761 (N_38761,N_37229,N_37805);
or U38762 (N_38762,N_37514,N_37572);
or U38763 (N_38763,N_37377,N_37397);
and U38764 (N_38764,N_37897,N_37422);
xnor U38765 (N_38765,N_37370,N_37112);
nor U38766 (N_38766,N_37087,N_37480);
nand U38767 (N_38767,N_37640,N_37481);
nand U38768 (N_38768,N_37704,N_37985);
or U38769 (N_38769,N_37788,N_37036);
nor U38770 (N_38770,N_37602,N_37756);
nor U38771 (N_38771,N_37415,N_37760);
and U38772 (N_38772,N_37030,N_37766);
and U38773 (N_38773,N_37726,N_37907);
or U38774 (N_38774,N_37660,N_37979);
or U38775 (N_38775,N_37105,N_37916);
nor U38776 (N_38776,N_37823,N_37299);
nand U38777 (N_38777,N_37825,N_37676);
or U38778 (N_38778,N_37024,N_37333);
and U38779 (N_38779,N_37820,N_37682);
nor U38780 (N_38780,N_37558,N_37666);
or U38781 (N_38781,N_37224,N_37364);
xor U38782 (N_38782,N_37167,N_37856);
xnor U38783 (N_38783,N_37530,N_37465);
or U38784 (N_38784,N_37197,N_37455);
or U38785 (N_38785,N_37702,N_37680);
or U38786 (N_38786,N_37865,N_37838);
nor U38787 (N_38787,N_37516,N_37232);
xor U38788 (N_38788,N_37382,N_37729);
xnor U38789 (N_38789,N_37499,N_37841);
xor U38790 (N_38790,N_37916,N_37872);
nand U38791 (N_38791,N_37000,N_37745);
or U38792 (N_38792,N_37400,N_37980);
nand U38793 (N_38793,N_37680,N_37174);
or U38794 (N_38794,N_37263,N_37252);
xnor U38795 (N_38795,N_37748,N_37786);
or U38796 (N_38796,N_37879,N_37139);
nor U38797 (N_38797,N_37149,N_37679);
nand U38798 (N_38798,N_37092,N_37809);
and U38799 (N_38799,N_37121,N_37535);
xor U38800 (N_38800,N_37428,N_37856);
or U38801 (N_38801,N_37051,N_37878);
and U38802 (N_38802,N_37024,N_37311);
nor U38803 (N_38803,N_37315,N_37093);
and U38804 (N_38804,N_37639,N_37915);
xnor U38805 (N_38805,N_37100,N_37787);
nor U38806 (N_38806,N_37257,N_37436);
nand U38807 (N_38807,N_37216,N_37917);
and U38808 (N_38808,N_37438,N_37828);
xnor U38809 (N_38809,N_37808,N_37783);
and U38810 (N_38810,N_37879,N_37553);
nand U38811 (N_38811,N_37694,N_37887);
nor U38812 (N_38812,N_37709,N_37391);
xnor U38813 (N_38813,N_37178,N_37298);
nor U38814 (N_38814,N_37892,N_37420);
xor U38815 (N_38815,N_37313,N_37762);
nand U38816 (N_38816,N_37888,N_37206);
xor U38817 (N_38817,N_37607,N_37834);
nand U38818 (N_38818,N_37272,N_37019);
and U38819 (N_38819,N_37807,N_37662);
and U38820 (N_38820,N_37079,N_37714);
nand U38821 (N_38821,N_37909,N_37481);
nand U38822 (N_38822,N_37914,N_37177);
and U38823 (N_38823,N_37724,N_37307);
nor U38824 (N_38824,N_37474,N_37266);
nand U38825 (N_38825,N_37219,N_37913);
and U38826 (N_38826,N_37636,N_37466);
nand U38827 (N_38827,N_37880,N_37693);
nand U38828 (N_38828,N_37512,N_37550);
xnor U38829 (N_38829,N_37202,N_37375);
xnor U38830 (N_38830,N_37114,N_37628);
and U38831 (N_38831,N_37580,N_37226);
and U38832 (N_38832,N_37306,N_37448);
xnor U38833 (N_38833,N_37769,N_37244);
nor U38834 (N_38834,N_37865,N_37884);
xnor U38835 (N_38835,N_37522,N_37937);
nor U38836 (N_38836,N_37578,N_37210);
nor U38837 (N_38837,N_37498,N_37583);
nand U38838 (N_38838,N_37330,N_37653);
and U38839 (N_38839,N_37316,N_37971);
nand U38840 (N_38840,N_37977,N_37283);
or U38841 (N_38841,N_37836,N_37415);
or U38842 (N_38842,N_37106,N_37950);
xor U38843 (N_38843,N_37439,N_37603);
nand U38844 (N_38844,N_37624,N_37577);
xor U38845 (N_38845,N_37854,N_37024);
nand U38846 (N_38846,N_37080,N_37823);
or U38847 (N_38847,N_37582,N_37377);
nand U38848 (N_38848,N_37583,N_37652);
nor U38849 (N_38849,N_37547,N_37110);
nand U38850 (N_38850,N_37498,N_37285);
nor U38851 (N_38851,N_37263,N_37012);
or U38852 (N_38852,N_37676,N_37308);
nor U38853 (N_38853,N_37255,N_37520);
xor U38854 (N_38854,N_37375,N_37907);
nor U38855 (N_38855,N_37913,N_37096);
or U38856 (N_38856,N_37512,N_37884);
and U38857 (N_38857,N_37365,N_37230);
nor U38858 (N_38858,N_37959,N_37383);
xnor U38859 (N_38859,N_37606,N_37557);
and U38860 (N_38860,N_37143,N_37402);
or U38861 (N_38861,N_37796,N_37220);
nor U38862 (N_38862,N_37357,N_37366);
nor U38863 (N_38863,N_37489,N_37955);
nand U38864 (N_38864,N_37105,N_37716);
nand U38865 (N_38865,N_37866,N_37290);
nor U38866 (N_38866,N_37535,N_37647);
xor U38867 (N_38867,N_37572,N_37883);
xnor U38868 (N_38868,N_37557,N_37596);
nor U38869 (N_38869,N_37741,N_37110);
or U38870 (N_38870,N_37163,N_37216);
and U38871 (N_38871,N_37245,N_37973);
or U38872 (N_38872,N_37636,N_37762);
xnor U38873 (N_38873,N_37873,N_37329);
xor U38874 (N_38874,N_37496,N_37959);
and U38875 (N_38875,N_37766,N_37235);
and U38876 (N_38876,N_37786,N_37712);
nor U38877 (N_38877,N_37220,N_37899);
and U38878 (N_38878,N_37974,N_37278);
and U38879 (N_38879,N_37349,N_37048);
and U38880 (N_38880,N_37125,N_37351);
and U38881 (N_38881,N_37155,N_37093);
nand U38882 (N_38882,N_37619,N_37835);
nor U38883 (N_38883,N_37353,N_37208);
nand U38884 (N_38884,N_37902,N_37034);
or U38885 (N_38885,N_37939,N_37273);
nand U38886 (N_38886,N_37398,N_37080);
nand U38887 (N_38887,N_37082,N_37764);
nor U38888 (N_38888,N_37233,N_37476);
nand U38889 (N_38889,N_37531,N_37346);
nor U38890 (N_38890,N_37066,N_37155);
nand U38891 (N_38891,N_37124,N_37120);
nor U38892 (N_38892,N_37176,N_37241);
xor U38893 (N_38893,N_37691,N_37765);
nor U38894 (N_38894,N_37093,N_37539);
nor U38895 (N_38895,N_37054,N_37588);
nor U38896 (N_38896,N_37021,N_37258);
xor U38897 (N_38897,N_37305,N_37694);
and U38898 (N_38898,N_37464,N_37662);
or U38899 (N_38899,N_37367,N_37880);
xor U38900 (N_38900,N_37774,N_37714);
and U38901 (N_38901,N_37092,N_37916);
nor U38902 (N_38902,N_37714,N_37394);
nor U38903 (N_38903,N_37977,N_37745);
xnor U38904 (N_38904,N_37097,N_37049);
and U38905 (N_38905,N_37461,N_37971);
and U38906 (N_38906,N_37625,N_37237);
or U38907 (N_38907,N_37913,N_37003);
nand U38908 (N_38908,N_37245,N_37758);
or U38909 (N_38909,N_37223,N_37499);
or U38910 (N_38910,N_37152,N_37605);
or U38911 (N_38911,N_37830,N_37158);
and U38912 (N_38912,N_37732,N_37411);
and U38913 (N_38913,N_37885,N_37238);
xnor U38914 (N_38914,N_37930,N_37931);
or U38915 (N_38915,N_37522,N_37749);
and U38916 (N_38916,N_37566,N_37990);
and U38917 (N_38917,N_37921,N_37939);
xnor U38918 (N_38918,N_37527,N_37266);
nand U38919 (N_38919,N_37147,N_37718);
or U38920 (N_38920,N_37681,N_37019);
and U38921 (N_38921,N_37241,N_37846);
or U38922 (N_38922,N_37114,N_37300);
and U38923 (N_38923,N_37689,N_37190);
and U38924 (N_38924,N_37033,N_37416);
xnor U38925 (N_38925,N_37663,N_37313);
and U38926 (N_38926,N_37513,N_37634);
and U38927 (N_38927,N_37102,N_37229);
or U38928 (N_38928,N_37909,N_37386);
and U38929 (N_38929,N_37923,N_37289);
nor U38930 (N_38930,N_37839,N_37518);
and U38931 (N_38931,N_37113,N_37592);
nand U38932 (N_38932,N_37767,N_37346);
nand U38933 (N_38933,N_37794,N_37418);
nand U38934 (N_38934,N_37873,N_37841);
nor U38935 (N_38935,N_37475,N_37705);
or U38936 (N_38936,N_37920,N_37753);
xor U38937 (N_38937,N_37308,N_37466);
xor U38938 (N_38938,N_37643,N_37229);
or U38939 (N_38939,N_37105,N_37651);
nand U38940 (N_38940,N_37123,N_37218);
and U38941 (N_38941,N_37570,N_37112);
or U38942 (N_38942,N_37585,N_37203);
or U38943 (N_38943,N_37858,N_37325);
or U38944 (N_38944,N_37830,N_37249);
xor U38945 (N_38945,N_37523,N_37876);
or U38946 (N_38946,N_37183,N_37928);
and U38947 (N_38947,N_37557,N_37491);
or U38948 (N_38948,N_37636,N_37918);
or U38949 (N_38949,N_37033,N_37052);
nor U38950 (N_38950,N_37871,N_37208);
xnor U38951 (N_38951,N_37303,N_37222);
nor U38952 (N_38952,N_37323,N_37361);
nor U38953 (N_38953,N_37078,N_37482);
nand U38954 (N_38954,N_37928,N_37323);
and U38955 (N_38955,N_37421,N_37252);
nand U38956 (N_38956,N_37595,N_37212);
xnor U38957 (N_38957,N_37321,N_37343);
nor U38958 (N_38958,N_37533,N_37279);
or U38959 (N_38959,N_37258,N_37664);
nor U38960 (N_38960,N_37964,N_37349);
or U38961 (N_38961,N_37845,N_37858);
nor U38962 (N_38962,N_37121,N_37806);
nor U38963 (N_38963,N_37953,N_37483);
nand U38964 (N_38964,N_37136,N_37153);
nand U38965 (N_38965,N_37825,N_37123);
xor U38966 (N_38966,N_37352,N_37687);
and U38967 (N_38967,N_37622,N_37453);
and U38968 (N_38968,N_37459,N_37142);
and U38969 (N_38969,N_37946,N_37871);
nor U38970 (N_38970,N_37931,N_37737);
and U38971 (N_38971,N_37141,N_37547);
nor U38972 (N_38972,N_37638,N_37711);
and U38973 (N_38973,N_37593,N_37607);
or U38974 (N_38974,N_37542,N_37517);
nand U38975 (N_38975,N_37199,N_37159);
nand U38976 (N_38976,N_37040,N_37207);
xor U38977 (N_38977,N_37735,N_37802);
nor U38978 (N_38978,N_37165,N_37680);
nand U38979 (N_38979,N_37207,N_37303);
xor U38980 (N_38980,N_37854,N_37858);
and U38981 (N_38981,N_37259,N_37879);
nand U38982 (N_38982,N_37738,N_37389);
nor U38983 (N_38983,N_37140,N_37647);
or U38984 (N_38984,N_37815,N_37843);
nor U38985 (N_38985,N_37023,N_37011);
nand U38986 (N_38986,N_37206,N_37159);
nand U38987 (N_38987,N_37473,N_37421);
and U38988 (N_38988,N_37954,N_37860);
nand U38989 (N_38989,N_37840,N_37528);
nand U38990 (N_38990,N_37486,N_37926);
xnor U38991 (N_38991,N_37543,N_37578);
xor U38992 (N_38992,N_37366,N_37702);
or U38993 (N_38993,N_37640,N_37983);
or U38994 (N_38994,N_37777,N_37253);
nand U38995 (N_38995,N_37338,N_37274);
or U38996 (N_38996,N_37109,N_37862);
nor U38997 (N_38997,N_37504,N_37466);
and U38998 (N_38998,N_37577,N_37927);
or U38999 (N_38999,N_37880,N_37817);
xor U39000 (N_39000,N_38113,N_38210);
or U39001 (N_39001,N_38613,N_38294);
nand U39002 (N_39002,N_38296,N_38285);
nor U39003 (N_39003,N_38843,N_38736);
nor U39004 (N_39004,N_38855,N_38989);
and U39005 (N_39005,N_38363,N_38487);
nor U39006 (N_39006,N_38637,N_38535);
nor U39007 (N_39007,N_38642,N_38191);
nand U39008 (N_39008,N_38242,N_38035);
xor U39009 (N_39009,N_38782,N_38229);
and U39010 (N_39010,N_38934,N_38721);
nand U39011 (N_39011,N_38972,N_38516);
nor U39012 (N_39012,N_38008,N_38207);
nand U39013 (N_39013,N_38530,N_38791);
and U39014 (N_39014,N_38343,N_38915);
and U39015 (N_39015,N_38331,N_38122);
xnor U39016 (N_39016,N_38981,N_38076);
nor U39017 (N_39017,N_38570,N_38097);
xor U39018 (N_39018,N_38817,N_38978);
or U39019 (N_39019,N_38534,N_38443);
xor U39020 (N_39020,N_38169,N_38785);
or U39021 (N_39021,N_38102,N_38917);
xnor U39022 (N_39022,N_38222,N_38582);
nand U39023 (N_39023,N_38722,N_38953);
or U39024 (N_39024,N_38057,N_38486);
nand U39025 (N_39025,N_38377,N_38248);
nor U39026 (N_39026,N_38970,N_38753);
and U39027 (N_39027,N_38900,N_38876);
nand U39028 (N_39028,N_38490,N_38325);
xor U39029 (N_39029,N_38819,N_38048);
xnor U39030 (N_39030,N_38882,N_38633);
or U39031 (N_39031,N_38653,N_38290);
and U39032 (N_39032,N_38404,N_38686);
xor U39033 (N_39033,N_38946,N_38904);
nand U39034 (N_39034,N_38902,N_38895);
or U39035 (N_39035,N_38383,N_38485);
nand U39036 (N_39036,N_38428,N_38052);
or U39037 (N_39037,N_38245,N_38312);
or U39038 (N_39038,N_38400,N_38279);
or U39039 (N_39039,N_38018,N_38381);
and U39040 (N_39040,N_38963,N_38072);
nor U39041 (N_39041,N_38185,N_38586);
xnor U39042 (N_39042,N_38495,N_38816);
nand U39043 (N_39043,N_38379,N_38778);
nand U39044 (N_39044,N_38051,N_38081);
and U39045 (N_39045,N_38403,N_38803);
xor U39046 (N_39046,N_38837,N_38440);
nand U39047 (N_39047,N_38987,N_38119);
xor U39048 (N_39048,N_38446,N_38992);
nor U39049 (N_39049,N_38725,N_38282);
or U39050 (N_39050,N_38158,N_38905);
xor U39051 (N_39051,N_38339,N_38342);
nor U39052 (N_39052,N_38111,N_38646);
nand U39053 (N_39053,N_38612,N_38459);
xor U39054 (N_39054,N_38644,N_38957);
or U39055 (N_39055,N_38674,N_38859);
xor U39056 (N_39056,N_38761,N_38483);
nor U39057 (N_39057,N_38851,N_38238);
nand U39058 (N_39058,N_38751,N_38489);
nor U39059 (N_39059,N_38519,N_38252);
and U39060 (N_39060,N_38969,N_38541);
or U39061 (N_39061,N_38398,N_38107);
or U39062 (N_39062,N_38512,N_38555);
xor U39063 (N_39063,N_38507,N_38679);
xnor U39064 (N_39064,N_38999,N_38591);
xor U39065 (N_39065,N_38596,N_38986);
nor U39066 (N_39066,N_38743,N_38083);
nor U39067 (N_39067,N_38028,N_38500);
and U39068 (N_39068,N_38773,N_38958);
xor U39069 (N_39069,N_38254,N_38000);
nand U39070 (N_39070,N_38856,N_38406);
or U39071 (N_39071,N_38426,N_38891);
and U39072 (N_39072,N_38645,N_38321);
nand U39073 (N_39073,N_38382,N_38200);
nor U39074 (N_39074,N_38233,N_38177);
or U39075 (N_39075,N_38824,N_38924);
nand U39076 (N_39076,N_38481,N_38409);
xnor U39077 (N_39077,N_38752,N_38874);
nor U39078 (N_39078,N_38421,N_38906);
and U39079 (N_39079,N_38250,N_38606);
or U39080 (N_39080,N_38808,N_38818);
and U39081 (N_39081,N_38871,N_38405);
nor U39082 (N_39082,N_38760,N_38857);
and U39083 (N_39083,N_38730,N_38619);
nor U39084 (N_39084,N_38961,N_38998);
and U39085 (N_39085,N_38356,N_38754);
nand U39086 (N_39086,N_38326,N_38598);
nor U39087 (N_39087,N_38926,N_38190);
nor U39088 (N_39088,N_38355,N_38968);
nand U39089 (N_39089,N_38746,N_38592);
and U39090 (N_39090,N_38231,N_38713);
nand U39091 (N_39091,N_38579,N_38657);
or U39092 (N_39092,N_38162,N_38885);
xor U39093 (N_39093,N_38468,N_38879);
xor U39094 (N_39094,N_38695,N_38246);
or U39095 (N_39095,N_38292,N_38788);
nand U39096 (N_39096,N_38607,N_38304);
nand U39097 (N_39097,N_38228,N_38572);
nor U39098 (N_39098,N_38431,N_38617);
nand U39099 (N_39099,N_38491,N_38236);
and U39100 (N_39100,N_38067,N_38070);
nor U39101 (N_39101,N_38801,N_38576);
and U39102 (N_39102,N_38344,N_38284);
and U39103 (N_39103,N_38216,N_38834);
nor U39104 (N_39104,N_38647,N_38848);
and U39105 (N_39105,N_38389,N_38444);
and U39106 (N_39106,N_38525,N_38849);
nor U39107 (N_39107,N_38029,N_38697);
and U39108 (N_39108,N_38557,N_38365);
or U39109 (N_39109,N_38880,N_38862);
xor U39110 (N_39110,N_38551,N_38194);
nand U39111 (N_39111,N_38449,N_38625);
nand U39112 (N_39112,N_38142,N_38441);
and U39113 (N_39113,N_38967,N_38839);
nor U39114 (N_39114,N_38127,N_38940);
xor U39115 (N_39115,N_38671,N_38451);
nor U39116 (N_39116,N_38407,N_38632);
or U39117 (N_39117,N_38781,N_38120);
xor U39118 (N_39118,N_38765,N_38032);
or U39119 (N_39119,N_38832,N_38826);
or U39120 (N_39120,N_38701,N_38141);
nand U39121 (N_39121,N_38890,N_38241);
and U39122 (N_39122,N_38622,N_38182);
nor U39123 (N_39123,N_38719,N_38694);
nor U39124 (N_39124,N_38706,N_38908);
and U39125 (N_39125,N_38423,N_38681);
and U39126 (N_39126,N_38889,N_38175);
or U39127 (N_39127,N_38584,N_38425);
xnor U39128 (N_39128,N_38023,N_38046);
nand U39129 (N_39129,N_38660,N_38714);
or U39130 (N_39130,N_38501,N_38258);
nand U39131 (N_39131,N_38330,N_38239);
or U39132 (N_39132,N_38410,N_38511);
and U39133 (N_39133,N_38875,N_38827);
and U39134 (N_39134,N_38437,N_38935);
or U39135 (N_39135,N_38505,N_38955);
nor U39136 (N_39136,N_38793,N_38307);
xnor U39137 (N_39137,N_38715,N_38655);
nor U39138 (N_39138,N_38353,N_38422);
and U39139 (N_39139,N_38977,N_38184);
nor U39140 (N_39140,N_38047,N_38792);
nand U39141 (N_39141,N_38213,N_38108);
or U39142 (N_39142,N_38881,N_38395);
nand U39143 (N_39143,N_38916,N_38959);
xor U39144 (N_39144,N_38424,N_38618);
nand U39145 (N_39145,N_38831,N_38698);
and U39146 (N_39146,N_38774,N_38341);
xor U39147 (N_39147,N_38723,N_38869);
nand U39148 (N_39148,N_38347,N_38496);
or U39149 (N_39149,N_38614,N_38259);
and U39150 (N_39150,N_38462,N_38966);
and U39151 (N_39151,N_38615,N_38952);
or U39152 (N_39152,N_38469,N_38894);
nor U39153 (N_39153,N_38965,N_38842);
nand U39154 (N_39154,N_38464,N_38776);
and U39155 (N_39155,N_38772,N_38094);
nor U39156 (N_39156,N_38984,N_38016);
nor U39157 (N_39157,N_38152,N_38962);
and U39158 (N_39158,N_38523,N_38019);
nand U39159 (N_39159,N_38463,N_38669);
or U39160 (N_39160,N_38453,N_38139);
xnor U39161 (N_39161,N_38093,N_38537);
or U39162 (N_39162,N_38274,N_38930);
xnor U39163 (N_39163,N_38771,N_38180);
or U39164 (N_39164,N_38460,N_38100);
nor U39165 (N_39165,N_38375,N_38115);
or U39166 (N_39166,N_38320,N_38610);
nand U39167 (N_39167,N_38936,N_38002);
xor U39168 (N_39168,N_38654,N_38982);
and U39169 (N_39169,N_38477,N_38517);
nor U39170 (N_39170,N_38209,N_38205);
or U39171 (N_39171,N_38049,N_38417);
nand U39172 (N_39172,N_38013,N_38208);
xnor U39173 (N_39173,N_38260,N_38420);
nand U39174 (N_39174,N_38741,N_38638);
or U39175 (N_39175,N_38798,N_38543);
nor U39176 (N_39176,N_38121,N_38080);
nor U39177 (N_39177,N_38004,N_38639);
nor U39178 (N_39178,N_38899,N_38345);
and U39179 (N_39179,N_38063,N_38003);
and U39180 (N_39180,N_38159,N_38281);
nand U39181 (N_39181,N_38418,N_38710);
xnor U39182 (N_39182,N_38357,N_38887);
nor U39183 (N_39183,N_38026,N_38179);
or U39184 (N_39184,N_38867,N_38435);
nand U39185 (N_39185,N_38041,N_38187);
nor U39186 (N_39186,N_38609,N_38058);
or U39187 (N_39187,N_38332,N_38755);
and U39188 (N_39188,N_38696,N_38225);
nand U39189 (N_39189,N_38001,N_38054);
or U39190 (N_39190,N_38560,N_38994);
nor U39191 (N_39191,N_38212,N_38861);
nor U39192 (N_39192,N_38084,N_38457);
or U39193 (N_39193,N_38866,N_38960);
nand U39194 (N_39194,N_38275,N_38183);
or U39195 (N_39195,N_38683,N_38578);
nand U39196 (N_39196,N_38661,N_38739);
nor U39197 (N_39197,N_38524,N_38256);
nand U39198 (N_39198,N_38566,N_38329);
nor U39199 (N_39199,N_38334,N_38430);
and U39200 (N_39200,N_38503,N_38542);
and U39201 (N_39201,N_38744,N_38699);
nor U39202 (N_39202,N_38502,N_38044);
and U39203 (N_39203,N_38295,N_38267);
nor U39204 (N_39204,N_38787,N_38224);
or U39205 (N_39205,N_38547,N_38085);
nor U39206 (N_39206,N_38458,N_38136);
or U39207 (N_39207,N_38948,N_38682);
and U39208 (N_39208,N_38903,N_38473);
or U39209 (N_39209,N_38471,N_38600);
nand U39210 (N_39210,N_38964,N_38797);
nand U39211 (N_39211,N_38309,N_38134);
xor U39212 (N_39212,N_38650,N_38556);
nand U39213 (N_39213,N_38597,N_38214);
xor U39214 (N_39214,N_38945,N_38846);
xor U39215 (N_39215,N_38550,N_38461);
or U39216 (N_39216,N_38075,N_38472);
nand U39217 (N_39217,N_38593,N_38601);
or U39218 (N_39218,N_38763,N_38154);
nor U39219 (N_39219,N_38160,N_38106);
nor U39220 (N_39220,N_38147,N_38769);
nand U39221 (N_39221,N_38039,N_38892);
or U39222 (N_39222,N_38310,N_38865);
or U39223 (N_39223,N_38494,N_38394);
nand U39224 (N_39224,N_38484,N_38221);
nand U39225 (N_39225,N_38372,N_38973);
nor U39226 (N_39226,N_38573,N_38391);
nand U39227 (N_39227,N_38174,N_38621);
or U39228 (N_39228,N_38742,N_38860);
and U39229 (N_39229,N_38884,N_38203);
nand U39230 (N_39230,N_38775,N_38432);
and U39231 (N_39231,N_38604,N_38980);
or U39232 (N_39232,N_38193,N_38515);
nand U39233 (N_39233,N_38131,N_38513);
and U39234 (N_39234,N_38711,N_38411);
nand U39235 (N_39235,N_38186,N_38976);
and U39236 (N_39236,N_38095,N_38812);
xnor U39237 (N_39237,N_38476,N_38204);
nor U39238 (N_39238,N_38358,N_38704);
xnor U39239 (N_39239,N_38171,N_38298);
xnor U39240 (N_39240,N_38918,N_38055);
nor U39241 (N_39241,N_38227,N_38943);
xnor U39242 (N_39242,N_38623,N_38314);
xnor U39243 (N_39243,N_38202,N_38921);
nor U39244 (N_39244,N_38079,N_38361);
or U39245 (N_39245,N_38027,N_38380);
xor U39246 (N_39246,N_38658,N_38036);
nor U39247 (N_39247,N_38868,N_38300);
or U39248 (N_39248,N_38807,N_38678);
nand U39249 (N_39249,N_38488,N_38844);
nand U39250 (N_39250,N_38038,N_38025);
nor U39251 (N_39251,N_38663,N_38168);
and U39252 (N_39252,N_38315,N_38251);
nor U39253 (N_39253,N_38031,N_38732);
or U39254 (N_39254,N_38691,N_38718);
and U39255 (N_39255,N_38814,N_38636);
or U39256 (N_39256,N_38230,N_38338);
or U39257 (N_39257,N_38928,N_38581);
or U39258 (N_39258,N_38983,N_38151);
and U39259 (N_39259,N_38929,N_38143);
xnor U39260 (N_39260,N_38319,N_38043);
xnor U39261 (N_39261,N_38033,N_38863);
and U39262 (N_39262,N_38056,N_38178);
nand U39263 (N_39263,N_38082,N_38217);
xnor U39264 (N_39264,N_38574,N_38901);
and U39265 (N_39265,N_38197,N_38727);
xnor U39266 (N_39266,N_38086,N_38415);
and U39267 (N_39267,N_38764,N_38240);
nor U39268 (N_39268,N_38235,N_38211);
or U39269 (N_39269,N_38497,N_38268);
xnor U39270 (N_39270,N_38132,N_38829);
xnor U39271 (N_39271,N_38408,N_38223);
and U39272 (N_39272,N_38652,N_38700);
and U39273 (N_39273,N_38521,N_38272);
and U39274 (N_39274,N_38749,N_38333);
nand U39275 (N_39275,N_38303,N_38594);
nor U39276 (N_39276,N_38014,N_38323);
nor U39277 (N_39277,N_38092,N_38181);
nand U39278 (N_39278,N_38318,N_38811);
xor U39279 (N_39279,N_38567,N_38112);
and U39280 (N_39280,N_38188,N_38447);
or U39281 (N_39281,N_38071,N_38492);
and U39282 (N_39282,N_38427,N_38724);
and U39283 (N_39283,N_38017,N_38944);
nor U39284 (N_39284,N_38821,N_38634);
xor U39285 (N_39285,N_38931,N_38124);
nor U39286 (N_39286,N_38450,N_38545);
nand U39287 (N_39287,N_38337,N_38909);
nand U39288 (N_39288,N_38089,N_38163);
and U39289 (N_39289,N_38110,N_38133);
or U39290 (N_39290,N_38020,N_38414);
or U39291 (N_39291,N_38933,N_38454);
nor U39292 (N_39292,N_38125,N_38580);
nand U39293 (N_39293,N_38034,N_38273);
nor U39294 (N_39294,N_38011,N_38261);
and U39295 (N_39295,N_38595,N_38288);
or U39296 (N_39296,N_38893,N_38397);
xor U39297 (N_39297,N_38907,N_38583);
and U39298 (N_39298,N_38677,N_38322);
or U39299 (N_39299,N_38243,N_38667);
nand U39300 (N_39300,N_38533,N_38438);
xor U39301 (N_39301,N_38412,N_38206);
nand U39302 (N_39302,N_38116,N_38324);
or U39303 (N_39303,N_38847,N_38413);
nor U39304 (N_39304,N_38308,N_38480);
nand U39305 (N_39305,N_38783,N_38479);
and U39306 (N_39306,N_38841,N_38278);
or U39307 (N_39307,N_38249,N_38030);
or U39308 (N_39308,N_38840,N_38305);
or U39309 (N_39309,N_38226,N_38368);
or U39310 (N_39310,N_38835,N_38616);
or U39311 (N_39311,N_38649,N_38950);
nor U39312 (N_39312,N_38872,N_38804);
or U39313 (N_39313,N_38779,N_38045);
xor U39314 (N_39314,N_38589,N_38280);
nor U39315 (N_39315,N_38378,N_38354);
nand U39316 (N_39316,N_38991,N_38684);
nand U39317 (N_39317,N_38668,N_38351);
xnor U39318 (N_39318,N_38757,N_38734);
nand U39319 (N_39319,N_38923,N_38552);
nor U39320 (N_39320,N_38146,N_38297);
xor U39321 (N_39321,N_38232,N_38135);
nand U39322 (N_39322,N_38703,N_38373);
nor U39323 (N_39323,N_38465,N_38088);
nor U39324 (N_39324,N_38676,N_38369);
and U39325 (N_39325,N_38605,N_38429);
and U39326 (N_39326,N_38506,N_38073);
and U39327 (N_39327,N_38795,N_38470);
or U39328 (N_39328,N_38442,N_38823);
nand U39329 (N_39329,N_38348,N_38687);
xor U39330 (N_39330,N_38629,N_38452);
xor U39331 (N_39331,N_38371,N_38362);
nor U39332 (N_39332,N_38283,N_38590);
and U39333 (N_39333,N_38149,N_38374);
and U39334 (N_39334,N_38201,N_38974);
nand U39335 (N_39335,N_38554,N_38558);
nor U39336 (N_39336,N_38888,N_38006);
xor U39337 (N_39337,N_38467,N_38050);
nand U39338 (N_39338,N_38815,N_38702);
nor U39339 (N_39339,N_38287,N_38705);
xnor U39340 (N_39340,N_38641,N_38833);
or U39341 (N_39341,N_38510,N_38350);
or U39342 (N_39342,N_38302,N_38434);
nand U39343 (N_39343,N_38809,N_38316);
nand U39344 (N_39344,N_38688,N_38564);
and U39345 (N_39345,N_38780,N_38603);
xnor U39346 (N_39346,N_38938,N_38720);
nor U39347 (N_39347,N_38077,N_38099);
xor U39348 (N_39348,N_38820,N_38608);
xnor U39349 (N_39349,N_38810,N_38886);
nor U39350 (N_39350,N_38068,N_38949);
or U39351 (N_39351,N_38393,N_38263);
nor U39352 (N_39352,N_38148,N_38109);
and U39353 (N_39353,N_38789,N_38577);
and U39354 (N_39354,N_38060,N_38009);
nand U39355 (N_39355,N_38173,N_38498);
nand U39356 (N_39356,N_38709,N_38877);
or U39357 (N_39357,N_38954,N_38078);
and U39358 (N_39358,N_38602,N_38898);
nor U39359 (N_39359,N_38640,N_38313);
and U39360 (N_39360,N_38117,N_38651);
nand U39361 (N_39361,N_38482,N_38825);
nor U39362 (N_39362,N_38666,N_38747);
nand U39363 (N_39363,N_38643,N_38198);
or U39364 (N_39364,N_38712,N_38932);
nor U39365 (N_39365,N_38975,N_38777);
or U39366 (N_39366,N_38914,N_38536);
xnor U39367 (N_39367,N_38620,N_38493);
and U39368 (N_39368,N_38024,N_38529);
and U39369 (N_39369,N_38767,N_38140);
or U39370 (N_39370,N_38317,N_38237);
nand U39371 (N_39371,N_38104,N_38768);
xnor U39372 (N_39372,N_38748,N_38144);
xnor U39373 (N_39373,N_38504,N_38830);
nor U39374 (N_39374,N_38707,N_38327);
xnor U39375 (N_39375,N_38247,N_38101);
xnor U39376 (N_39376,N_38897,N_38439);
nor U39377 (N_39377,N_38218,N_38475);
nor U39378 (N_39378,N_38571,N_38074);
or U39379 (N_39379,N_38359,N_38387);
xnor U39380 (N_39380,N_38852,N_38416);
nand U39381 (N_39381,N_38126,N_38951);
nor U39382 (N_39382,N_38277,N_38012);
or U39383 (N_39383,N_38770,N_38137);
or U39384 (N_39384,N_38920,N_38784);
or U39385 (N_39385,N_38386,N_38648);
nor U39386 (N_39386,N_38340,N_38396);
and U39387 (N_39387,N_38262,N_38790);
or U39388 (N_39388,N_38087,N_38360);
xnor U39389 (N_39389,N_38561,N_38123);
nand U39390 (N_39390,N_38005,N_38456);
nor U39391 (N_39391,N_38199,N_38759);
and U39392 (N_39392,N_38522,N_38195);
nor U39393 (N_39393,N_38271,N_38672);
nand U39394 (N_39394,N_38189,N_38390);
xnor U39395 (N_39395,N_38588,N_38433);
nor U39396 (N_39396,N_38499,N_38836);
or U39397 (N_39397,N_38270,N_38685);
nand U39398 (N_39398,N_38170,N_38828);
nor U39399 (N_39399,N_38675,N_38015);
nand U39400 (N_39400,N_38253,N_38166);
nand U39401 (N_39401,N_38883,N_38802);
nand U39402 (N_39402,N_38103,N_38693);
nor U39403 (N_39403,N_38805,N_38010);
or U39404 (N_39404,N_38234,N_38346);
xor U39405 (N_39405,N_38822,N_38587);
nand U39406 (N_39406,N_38167,N_38896);
nand U39407 (N_39407,N_38269,N_38255);
and U39408 (N_39408,N_38064,N_38971);
nor U39409 (N_39409,N_38568,N_38585);
nand U39410 (N_39410,N_38145,N_38153);
nand U39411 (N_39411,N_38455,N_38990);
nand U39412 (N_39412,N_38726,N_38448);
and U39413 (N_39413,N_38392,N_38257);
nor U39414 (N_39414,N_38508,N_38436);
and U39415 (N_39415,N_38664,N_38766);
or U39416 (N_39416,N_38128,N_38911);
or U39417 (N_39417,N_38306,N_38611);
nor U39418 (N_39418,N_38569,N_38873);
or U39419 (N_39419,N_38925,N_38689);
nand U39420 (N_39420,N_38265,N_38670);
xor U39421 (N_39421,N_38528,N_38913);
nand U39422 (N_39422,N_38546,N_38384);
xor U39423 (N_39423,N_38635,N_38367);
nor U39424 (N_39424,N_38090,N_38069);
nand U39425 (N_39425,N_38059,N_38853);
or U39426 (N_39426,N_38690,N_38527);
xor U39427 (N_39427,N_38680,N_38665);
or U39428 (N_39428,N_38445,N_38164);
nand U39429 (N_39429,N_38729,N_38738);
nand U39430 (N_39430,N_38376,N_38165);
nand U39431 (N_39431,N_38737,N_38565);
nand U39432 (N_39432,N_38539,N_38062);
nand U39433 (N_39433,N_38096,N_38399);
or U39434 (N_39434,N_38532,N_38118);
nor U39435 (N_39435,N_38845,N_38289);
nor U39436 (N_39436,N_38708,N_38750);
and U39437 (N_39437,N_38947,N_38286);
nor U39438 (N_39438,N_38518,N_38870);
nor U39439 (N_39439,N_38098,N_38150);
or U39440 (N_39440,N_38910,N_38796);
nor U39441 (N_39441,N_38401,N_38388);
and U39442 (N_39442,N_38786,N_38366);
and U39443 (N_39443,N_38864,N_38402);
or U39444 (N_39444,N_38538,N_38370);
nor U39445 (N_39445,N_38740,N_38756);
and U39446 (N_39446,N_38758,N_38301);
and U39447 (N_39447,N_38673,N_38364);
nand U39448 (N_39448,N_38040,N_38922);
xnor U39449 (N_39449,N_38196,N_38692);
nand U39450 (N_39450,N_38628,N_38176);
or U39451 (N_39451,N_38627,N_38575);
xnor U39452 (N_39452,N_38311,N_38022);
and U39453 (N_39453,N_38352,N_38466);
and U39454 (N_39454,N_38531,N_38540);
nor U39455 (N_39455,N_38912,N_38662);
or U39456 (N_39456,N_38264,N_38996);
or U39457 (N_39457,N_38838,N_38735);
and U39458 (N_39458,N_38878,N_38937);
nor U39459 (N_39459,N_38599,N_38563);
or U39460 (N_39460,N_38385,N_38850);
xor U39461 (N_39461,N_38299,N_38419);
xor U39462 (N_39462,N_38161,N_38220);
nand U39463 (N_39463,N_38942,N_38526);
xnor U39464 (N_39464,N_38559,N_38919);
and U39465 (N_39465,N_38065,N_38474);
and U39466 (N_39466,N_38745,N_38659);
nor U39467 (N_39467,N_38995,N_38105);
nand U39468 (N_39468,N_38129,N_38138);
and U39469 (N_39469,N_38335,N_38172);
nor U39470 (N_39470,N_38155,N_38858);
xnor U39471 (N_39471,N_38349,N_38626);
nor U39472 (N_39472,N_38544,N_38731);
nor U39473 (N_39473,N_38549,N_38061);
xor U39474 (N_39474,N_38114,N_38037);
or U39475 (N_39475,N_38520,N_38656);
nor U39476 (N_39476,N_38762,N_38266);
and U39477 (N_39477,N_38800,N_38007);
xnor U39478 (N_39478,N_38728,N_38328);
nand U39479 (N_39479,N_38794,N_38291);
nor U39480 (N_39480,N_38988,N_38478);
xor U39481 (N_39481,N_38336,N_38717);
xor U39482 (N_39482,N_38806,N_38156);
nor U39483 (N_39483,N_38293,N_38813);
nor U39484 (N_39484,N_38053,N_38553);
and U39485 (N_39485,N_38066,N_38091);
and U39486 (N_39486,N_38799,N_38939);
nand U39487 (N_39487,N_38624,N_38130);
nand U39488 (N_39488,N_38733,N_38562);
xnor U39489 (N_39489,N_38042,N_38021);
and U39490 (N_39490,N_38276,N_38514);
and U39491 (N_39491,N_38854,N_38985);
nand U39492 (N_39492,N_38993,N_38956);
and U39493 (N_39493,N_38548,N_38979);
xor U39494 (N_39494,N_38716,N_38192);
nor U39495 (N_39495,N_38941,N_38997);
nand U39496 (N_39496,N_38927,N_38630);
nand U39497 (N_39497,N_38215,N_38244);
and U39498 (N_39498,N_38219,N_38157);
or U39499 (N_39499,N_38509,N_38631);
or U39500 (N_39500,N_38696,N_38092);
nor U39501 (N_39501,N_38959,N_38873);
or U39502 (N_39502,N_38986,N_38496);
nor U39503 (N_39503,N_38177,N_38035);
xor U39504 (N_39504,N_38461,N_38431);
xnor U39505 (N_39505,N_38933,N_38789);
or U39506 (N_39506,N_38085,N_38102);
xor U39507 (N_39507,N_38230,N_38704);
and U39508 (N_39508,N_38042,N_38442);
nand U39509 (N_39509,N_38211,N_38338);
and U39510 (N_39510,N_38585,N_38873);
nand U39511 (N_39511,N_38540,N_38322);
and U39512 (N_39512,N_38352,N_38626);
and U39513 (N_39513,N_38437,N_38248);
nand U39514 (N_39514,N_38633,N_38987);
xor U39515 (N_39515,N_38315,N_38438);
xor U39516 (N_39516,N_38498,N_38762);
nor U39517 (N_39517,N_38017,N_38931);
nor U39518 (N_39518,N_38621,N_38999);
nor U39519 (N_39519,N_38823,N_38777);
nand U39520 (N_39520,N_38617,N_38926);
nor U39521 (N_39521,N_38990,N_38291);
nand U39522 (N_39522,N_38930,N_38487);
xor U39523 (N_39523,N_38130,N_38431);
and U39524 (N_39524,N_38803,N_38316);
or U39525 (N_39525,N_38458,N_38531);
nor U39526 (N_39526,N_38615,N_38358);
xor U39527 (N_39527,N_38476,N_38505);
nor U39528 (N_39528,N_38474,N_38222);
and U39529 (N_39529,N_38696,N_38402);
and U39530 (N_39530,N_38655,N_38385);
nand U39531 (N_39531,N_38287,N_38877);
xnor U39532 (N_39532,N_38322,N_38372);
nor U39533 (N_39533,N_38690,N_38569);
or U39534 (N_39534,N_38834,N_38014);
nor U39535 (N_39535,N_38970,N_38907);
or U39536 (N_39536,N_38488,N_38551);
and U39537 (N_39537,N_38330,N_38912);
or U39538 (N_39538,N_38852,N_38639);
or U39539 (N_39539,N_38042,N_38653);
xnor U39540 (N_39540,N_38541,N_38806);
and U39541 (N_39541,N_38109,N_38080);
xor U39542 (N_39542,N_38132,N_38750);
xnor U39543 (N_39543,N_38516,N_38112);
or U39544 (N_39544,N_38993,N_38978);
nand U39545 (N_39545,N_38611,N_38510);
and U39546 (N_39546,N_38093,N_38793);
xnor U39547 (N_39547,N_38229,N_38395);
and U39548 (N_39548,N_38239,N_38671);
and U39549 (N_39549,N_38357,N_38587);
and U39550 (N_39550,N_38182,N_38581);
nand U39551 (N_39551,N_38125,N_38898);
and U39552 (N_39552,N_38525,N_38503);
nand U39553 (N_39553,N_38828,N_38444);
or U39554 (N_39554,N_38271,N_38040);
or U39555 (N_39555,N_38915,N_38540);
and U39556 (N_39556,N_38274,N_38725);
and U39557 (N_39557,N_38128,N_38626);
nand U39558 (N_39558,N_38183,N_38766);
and U39559 (N_39559,N_38616,N_38950);
xor U39560 (N_39560,N_38909,N_38647);
nor U39561 (N_39561,N_38171,N_38384);
and U39562 (N_39562,N_38743,N_38918);
or U39563 (N_39563,N_38891,N_38028);
nand U39564 (N_39564,N_38429,N_38819);
or U39565 (N_39565,N_38376,N_38982);
or U39566 (N_39566,N_38582,N_38974);
nand U39567 (N_39567,N_38035,N_38210);
or U39568 (N_39568,N_38091,N_38312);
or U39569 (N_39569,N_38137,N_38199);
nor U39570 (N_39570,N_38735,N_38960);
nor U39571 (N_39571,N_38435,N_38730);
and U39572 (N_39572,N_38117,N_38644);
nor U39573 (N_39573,N_38489,N_38117);
nand U39574 (N_39574,N_38213,N_38904);
and U39575 (N_39575,N_38148,N_38729);
or U39576 (N_39576,N_38463,N_38129);
and U39577 (N_39577,N_38483,N_38425);
nand U39578 (N_39578,N_38408,N_38536);
nor U39579 (N_39579,N_38691,N_38557);
nor U39580 (N_39580,N_38411,N_38713);
nor U39581 (N_39581,N_38846,N_38118);
or U39582 (N_39582,N_38210,N_38050);
or U39583 (N_39583,N_38606,N_38941);
or U39584 (N_39584,N_38863,N_38023);
and U39585 (N_39585,N_38114,N_38554);
and U39586 (N_39586,N_38094,N_38689);
and U39587 (N_39587,N_38755,N_38716);
and U39588 (N_39588,N_38165,N_38180);
nor U39589 (N_39589,N_38309,N_38067);
xor U39590 (N_39590,N_38410,N_38526);
nor U39591 (N_39591,N_38337,N_38082);
nor U39592 (N_39592,N_38213,N_38333);
and U39593 (N_39593,N_38192,N_38199);
and U39594 (N_39594,N_38937,N_38002);
or U39595 (N_39595,N_38094,N_38015);
nand U39596 (N_39596,N_38351,N_38555);
xor U39597 (N_39597,N_38666,N_38203);
nor U39598 (N_39598,N_38759,N_38133);
nor U39599 (N_39599,N_38079,N_38060);
and U39600 (N_39600,N_38183,N_38922);
xnor U39601 (N_39601,N_38780,N_38185);
nand U39602 (N_39602,N_38990,N_38920);
and U39603 (N_39603,N_38399,N_38541);
and U39604 (N_39604,N_38603,N_38417);
and U39605 (N_39605,N_38265,N_38823);
and U39606 (N_39606,N_38566,N_38103);
nand U39607 (N_39607,N_38734,N_38344);
or U39608 (N_39608,N_38383,N_38051);
or U39609 (N_39609,N_38486,N_38474);
and U39610 (N_39610,N_38092,N_38428);
nand U39611 (N_39611,N_38498,N_38658);
nand U39612 (N_39612,N_38707,N_38197);
nand U39613 (N_39613,N_38834,N_38134);
nor U39614 (N_39614,N_38149,N_38782);
xor U39615 (N_39615,N_38041,N_38554);
xnor U39616 (N_39616,N_38445,N_38511);
xor U39617 (N_39617,N_38545,N_38928);
or U39618 (N_39618,N_38700,N_38368);
nand U39619 (N_39619,N_38857,N_38349);
nand U39620 (N_39620,N_38753,N_38816);
or U39621 (N_39621,N_38560,N_38586);
and U39622 (N_39622,N_38482,N_38194);
nor U39623 (N_39623,N_38188,N_38573);
nor U39624 (N_39624,N_38509,N_38900);
nand U39625 (N_39625,N_38221,N_38237);
or U39626 (N_39626,N_38871,N_38220);
xnor U39627 (N_39627,N_38676,N_38189);
or U39628 (N_39628,N_38229,N_38291);
and U39629 (N_39629,N_38542,N_38258);
or U39630 (N_39630,N_38325,N_38746);
and U39631 (N_39631,N_38671,N_38978);
or U39632 (N_39632,N_38870,N_38580);
xor U39633 (N_39633,N_38801,N_38902);
nand U39634 (N_39634,N_38097,N_38217);
nand U39635 (N_39635,N_38889,N_38738);
or U39636 (N_39636,N_38681,N_38881);
xor U39637 (N_39637,N_38442,N_38017);
or U39638 (N_39638,N_38268,N_38773);
xor U39639 (N_39639,N_38168,N_38129);
and U39640 (N_39640,N_38583,N_38121);
xnor U39641 (N_39641,N_38193,N_38492);
or U39642 (N_39642,N_38557,N_38784);
or U39643 (N_39643,N_38079,N_38338);
xnor U39644 (N_39644,N_38097,N_38931);
and U39645 (N_39645,N_38693,N_38955);
nor U39646 (N_39646,N_38961,N_38059);
nor U39647 (N_39647,N_38467,N_38174);
xor U39648 (N_39648,N_38415,N_38929);
or U39649 (N_39649,N_38026,N_38522);
nand U39650 (N_39650,N_38277,N_38285);
and U39651 (N_39651,N_38325,N_38435);
and U39652 (N_39652,N_38465,N_38019);
and U39653 (N_39653,N_38897,N_38527);
nor U39654 (N_39654,N_38818,N_38103);
or U39655 (N_39655,N_38266,N_38452);
nor U39656 (N_39656,N_38687,N_38178);
xor U39657 (N_39657,N_38780,N_38655);
or U39658 (N_39658,N_38088,N_38058);
nand U39659 (N_39659,N_38218,N_38898);
nand U39660 (N_39660,N_38251,N_38365);
and U39661 (N_39661,N_38902,N_38651);
nor U39662 (N_39662,N_38695,N_38310);
or U39663 (N_39663,N_38459,N_38414);
xor U39664 (N_39664,N_38658,N_38969);
xor U39665 (N_39665,N_38564,N_38301);
nand U39666 (N_39666,N_38085,N_38057);
or U39667 (N_39667,N_38827,N_38304);
xor U39668 (N_39668,N_38410,N_38902);
or U39669 (N_39669,N_38169,N_38553);
and U39670 (N_39670,N_38694,N_38745);
nor U39671 (N_39671,N_38569,N_38282);
nor U39672 (N_39672,N_38678,N_38696);
or U39673 (N_39673,N_38085,N_38304);
and U39674 (N_39674,N_38707,N_38387);
xnor U39675 (N_39675,N_38482,N_38812);
and U39676 (N_39676,N_38222,N_38699);
nor U39677 (N_39677,N_38887,N_38915);
xnor U39678 (N_39678,N_38516,N_38735);
nand U39679 (N_39679,N_38304,N_38569);
and U39680 (N_39680,N_38526,N_38045);
nor U39681 (N_39681,N_38325,N_38922);
or U39682 (N_39682,N_38621,N_38833);
xnor U39683 (N_39683,N_38106,N_38141);
xor U39684 (N_39684,N_38720,N_38312);
and U39685 (N_39685,N_38815,N_38765);
xor U39686 (N_39686,N_38676,N_38001);
or U39687 (N_39687,N_38098,N_38818);
nor U39688 (N_39688,N_38893,N_38611);
nand U39689 (N_39689,N_38143,N_38055);
nand U39690 (N_39690,N_38425,N_38406);
or U39691 (N_39691,N_38409,N_38712);
or U39692 (N_39692,N_38870,N_38983);
and U39693 (N_39693,N_38439,N_38342);
xor U39694 (N_39694,N_38569,N_38450);
or U39695 (N_39695,N_38073,N_38960);
nor U39696 (N_39696,N_38586,N_38447);
or U39697 (N_39697,N_38600,N_38964);
nor U39698 (N_39698,N_38390,N_38136);
nand U39699 (N_39699,N_38927,N_38918);
and U39700 (N_39700,N_38122,N_38032);
and U39701 (N_39701,N_38632,N_38775);
and U39702 (N_39702,N_38582,N_38848);
and U39703 (N_39703,N_38128,N_38324);
xnor U39704 (N_39704,N_38413,N_38929);
nand U39705 (N_39705,N_38460,N_38113);
and U39706 (N_39706,N_38343,N_38731);
nor U39707 (N_39707,N_38269,N_38310);
xor U39708 (N_39708,N_38522,N_38419);
and U39709 (N_39709,N_38279,N_38833);
or U39710 (N_39710,N_38882,N_38440);
nand U39711 (N_39711,N_38467,N_38324);
xor U39712 (N_39712,N_38635,N_38405);
xnor U39713 (N_39713,N_38853,N_38630);
nand U39714 (N_39714,N_38729,N_38931);
xor U39715 (N_39715,N_38947,N_38856);
xor U39716 (N_39716,N_38829,N_38514);
xnor U39717 (N_39717,N_38747,N_38827);
or U39718 (N_39718,N_38722,N_38834);
xnor U39719 (N_39719,N_38390,N_38015);
nand U39720 (N_39720,N_38699,N_38370);
or U39721 (N_39721,N_38295,N_38953);
or U39722 (N_39722,N_38294,N_38240);
and U39723 (N_39723,N_38618,N_38223);
or U39724 (N_39724,N_38090,N_38522);
or U39725 (N_39725,N_38121,N_38532);
nand U39726 (N_39726,N_38496,N_38201);
nor U39727 (N_39727,N_38944,N_38335);
or U39728 (N_39728,N_38822,N_38229);
xor U39729 (N_39729,N_38214,N_38608);
and U39730 (N_39730,N_38830,N_38682);
or U39731 (N_39731,N_38341,N_38137);
nor U39732 (N_39732,N_38231,N_38109);
nand U39733 (N_39733,N_38164,N_38373);
nor U39734 (N_39734,N_38580,N_38387);
xor U39735 (N_39735,N_38766,N_38723);
and U39736 (N_39736,N_38860,N_38073);
nand U39737 (N_39737,N_38652,N_38598);
or U39738 (N_39738,N_38742,N_38763);
xor U39739 (N_39739,N_38308,N_38003);
or U39740 (N_39740,N_38478,N_38782);
nand U39741 (N_39741,N_38367,N_38156);
nor U39742 (N_39742,N_38871,N_38457);
nor U39743 (N_39743,N_38464,N_38869);
nand U39744 (N_39744,N_38340,N_38445);
nand U39745 (N_39745,N_38094,N_38288);
or U39746 (N_39746,N_38216,N_38045);
xor U39747 (N_39747,N_38123,N_38577);
or U39748 (N_39748,N_38203,N_38809);
or U39749 (N_39749,N_38504,N_38589);
nor U39750 (N_39750,N_38028,N_38664);
and U39751 (N_39751,N_38807,N_38965);
xnor U39752 (N_39752,N_38977,N_38946);
nor U39753 (N_39753,N_38085,N_38636);
nor U39754 (N_39754,N_38413,N_38126);
or U39755 (N_39755,N_38293,N_38211);
nand U39756 (N_39756,N_38347,N_38750);
and U39757 (N_39757,N_38883,N_38700);
nor U39758 (N_39758,N_38225,N_38591);
nor U39759 (N_39759,N_38785,N_38202);
nor U39760 (N_39760,N_38211,N_38720);
nor U39761 (N_39761,N_38319,N_38580);
xor U39762 (N_39762,N_38692,N_38955);
nor U39763 (N_39763,N_38041,N_38079);
xnor U39764 (N_39764,N_38476,N_38374);
nor U39765 (N_39765,N_38127,N_38736);
xor U39766 (N_39766,N_38186,N_38797);
nand U39767 (N_39767,N_38427,N_38075);
or U39768 (N_39768,N_38144,N_38134);
nor U39769 (N_39769,N_38496,N_38495);
nor U39770 (N_39770,N_38944,N_38080);
nor U39771 (N_39771,N_38160,N_38236);
nand U39772 (N_39772,N_38076,N_38168);
xor U39773 (N_39773,N_38647,N_38216);
and U39774 (N_39774,N_38629,N_38563);
and U39775 (N_39775,N_38409,N_38746);
nor U39776 (N_39776,N_38492,N_38745);
nand U39777 (N_39777,N_38647,N_38538);
and U39778 (N_39778,N_38868,N_38832);
nand U39779 (N_39779,N_38085,N_38392);
and U39780 (N_39780,N_38128,N_38231);
and U39781 (N_39781,N_38732,N_38709);
and U39782 (N_39782,N_38832,N_38472);
and U39783 (N_39783,N_38434,N_38558);
xor U39784 (N_39784,N_38446,N_38852);
xnor U39785 (N_39785,N_38930,N_38212);
or U39786 (N_39786,N_38515,N_38834);
or U39787 (N_39787,N_38764,N_38342);
nor U39788 (N_39788,N_38865,N_38616);
or U39789 (N_39789,N_38494,N_38994);
nor U39790 (N_39790,N_38296,N_38218);
nor U39791 (N_39791,N_38946,N_38183);
nand U39792 (N_39792,N_38386,N_38045);
or U39793 (N_39793,N_38732,N_38385);
or U39794 (N_39794,N_38391,N_38852);
or U39795 (N_39795,N_38755,N_38493);
or U39796 (N_39796,N_38816,N_38472);
or U39797 (N_39797,N_38779,N_38329);
or U39798 (N_39798,N_38369,N_38495);
or U39799 (N_39799,N_38122,N_38863);
nand U39800 (N_39800,N_38602,N_38001);
xor U39801 (N_39801,N_38999,N_38524);
or U39802 (N_39802,N_38824,N_38427);
nor U39803 (N_39803,N_38565,N_38952);
and U39804 (N_39804,N_38647,N_38594);
nand U39805 (N_39805,N_38640,N_38535);
or U39806 (N_39806,N_38796,N_38303);
xor U39807 (N_39807,N_38275,N_38056);
and U39808 (N_39808,N_38014,N_38204);
or U39809 (N_39809,N_38195,N_38656);
or U39810 (N_39810,N_38295,N_38419);
and U39811 (N_39811,N_38740,N_38307);
nor U39812 (N_39812,N_38325,N_38357);
nor U39813 (N_39813,N_38044,N_38298);
or U39814 (N_39814,N_38631,N_38914);
or U39815 (N_39815,N_38162,N_38309);
or U39816 (N_39816,N_38307,N_38977);
xor U39817 (N_39817,N_38545,N_38132);
and U39818 (N_39818,N_38759,N_38952);
nor U39819 (N_39819,N_38141,N_38209);
xnor U39820 (N_39820,N_38861,N_38975);
and U39821 (N_39821,N_38158,N_38955);
nand U39822 (N_39822,N_38460,N_38364);
and U39823 (N_39823,N_38338,N_38851);
and U39824 (N_39824,N_38144,N_38045);
or U39825 (N_39825,N_38128,N_38146);
and U39826 (N_39826,N_38224,N_38858);
nand U39827 (N_39827,N_38782,N_38212);
and U39828 (N_39828,N_38861,N_38607);
or U39829 (N_39829,N_38145,N_38782);
or U39830 (N_39830,N_38207,N_38871);
nand U39831 (N_39831,N_38527,N_38734);
nor U39832 (N_39832,N_38959,N_38874);
xnor U39833 (N_39833,N_38121,N_38562);
and U39834 (N_39834,N_38189,N_38182);
and U39835 (N_39835,N_38926,N_38847);
nor U39836 (N_39836,N_38249,N_38281);
xnor U39837 (N_39837,N_38045,N_38985);
nor U39838 (N_39838,N_38249,N_38613);
or U39839 (N_39839,N_38115,N_38921);
or U39840 (N_39840,N_38211,N_38320);
nand U39841 (N_39841,N_38945,N_38309);
xor U39842 (N_39842,N_38450,N_38122);
or U39843 (N_39843,N_38598,N_38968);
nand U39844 (N_39844,N_38588,N_38251);
xor U39845 (N_39845,N_38605,N_38720);
nand U39846 (N_39846,N_38908,N_38063);
nand U39847 (N_39847,N_38334,N_38012);
xor U39848 (N_39848,N_38534,N_38829);
nand U39849 (N_39849,N_38137,N_38100);
or U39850 (N_39850,N_38434,N_38911);
xnor U39851 (N_39851,N_38627,N_38192);
nor U39852 (N_39852,N_38305,N_38641);
nand U39853 (N_39853,N_38251,N_38533);
nor U39854 (N_39854,N_38590,N_38051);
or U39855 (N_39855,N_38185,N_38886);
and U39856 (N_39856,N_38335,N_38936);
or U39857 (N_39857,N_38540,N_38048);
or U39858 (N_39858,N_38011,N_38233);
and U39859 (N_39859,N_38557,N_38385);
xor U39860 (N_39860,N_38155,N_38099);
or U39861 (N_39861,N_38493,N_38095);
and U39862 (N_39862,N_38101,N_38274);
nor U39863 (N_39863,N_38335,N_38715);
nor U39864 (N_39864,N_38886,N_38589);
or U39865 (N_39865,N_38381,N_38990);
xnor U39866 (N_39866,N_38441,N_38638);
and U39867 (N_39867,N_38227,N_38938);
xor U39868 (N_39868,N_38479,N_38498);
nand U39869 (N_39869,N_38524,N_38853);
and U39870 (N_39870,N_38533,N_38132);
and U39871 (N_39871,N_38295,N_38171);
or U39872 (N_39872,N_38904,N_38570);
xor U39873 (N_39873,N_38888,N_38619);
or U39874 (N_39874,N_38688,N_38760);
nand U39875 (N_39875,N_38117,N_38526);
nand U39876 (N_39876,N_38438,N_38894);
nand U39877 (N_39877,N_38293,N_38003);
xor U39878 (N_39878,N_38181,N_38950);
and U39879 (N_39879,N_38696,N_38029);
or U39880 (N_39880,N_38855,N_38167);
nor U39881 (N_39881,N_38728,N_38621);
xor U39882 (N_39882,N_38000,N_38235);
xnor U39883 (N_39883,N_38104,N_38635);
nor U39884 (N_39884,N_38476,N_38623);
and U39885 (N_39885,N_38124,N_38925);
nor U39886 (N_39886,N_38721,N_38396);
or U39887 (N_39887,N_38604,N_38909);
or U39888 (N_39888,N_38612,N_38818);
or U39889 (N_39889,N_38391,N_38260);
or U39890 (N_39890,N_38882,N_38393);
nor U39891 (N_39891,N_38449,N_38318);
nand U39892 (N_39892,N_38707,N_38678);
and U39893 (N_39893,N_38235,N_38320);
nor U39894 (N_39894,N_38712,N_38153);
xor U39895 (N_39895,N_38437,N_38366);
nand U39896 (N_39896,N_38048,N_38058);
nand U39897 (N_39897,N_38967,N_38763);
or U39898 (N_39898,N_38909,N_38570);
nor U39899 (N_39899,N_38984,N_38559);
nand U39900 (N_39900,N_38946,N_38814);
or U39901 (N_39901,N_38063,N_38087);
nand U39902 (N_39902,N_38103,N_38740);
nor U39903 (N_39903,N_38546,N_38158);
and U39904 (N_39904,N_38947,N_38497);
nor U39905 (N_39905,N_38976,N_38227);
and U39906 (N_39906,N_38583,N_38321);
xor U39907 (N_39907,N_38902,N_38896);
xor U39908 (N_39908,N_38812,N_38699);
nand U39909 (N_39909,N_38455,N_38504);
or U39910 (N_39910,N_38832,N_38308);
and U39911 (N_39911,N_38461,N_38648);
nand U39912 (N_39912,N_38752,N_38531);
and U39913 (N_39913,N_38773,N_38757);
nand U39914 (N_39914,N_38345,N_38359);
and U39915 (N_39915,N_38797,N_38376);
xor U39916 (N_39916,N_38065,N_38075);
or U39917 (N_39917,N_38296,N_38318);
and U39918 (N_39918,N_38873,N_38489);
or U39919 (N_39919,N_38770,N_38302);
nand U39920 (N_39920,N_38582,N_38281);
and U39921 (N_39921,N_38143,N_38646);
nor U39922 (N_39922,N_38524,N_38033);
nor U39923 (N_39923,N_38984,N_38952);
and U39924 (N_39924,N_38874,N_38926);
and U39925 (N_39925,N_38738,N_38961);
or U39926 (N_39926,N_38765,N_38680);
and U39927 (N_39927,N_38657,N_38430);
nor U39928 (N_39928,N_38903,N_38724);
nand U39929 (N_39929,N_38353,N_38052);
nor U39930 (N_39930,N_38662,N_38432);
nor U39931 (N_39931,N_38915,N_38002);
nand U39932 (N_39932,N_38207,N_38588);
xor U39933 (N_39933,N_38347,N_38373);
nor U39934 (N_39934,N_38942,N_38128);
and U39935 (N_39935,N_38209,N_38535);
nor U39936 (N_39936,N_38598,N_38500);
nor U39937 (N_39937,N_38790,N_38581);
nor U39938 (N_39938,N_38644,N_38434);
nand U39939 (N_39939,N_38123,N_38051);
or U39940 (N_39940,N_38527,N_38476);
and U39941 (N_39941,N_38620,N_38887);
or U39942 (N_39942,N_38171,N_38360);
or U39943 (N_39943,N_38034,N_38216);
or U39944 (N_39944,N_38488,N_38252);
xor U39945 (N_39945,N_38946,N_38305);
xor U39946 (N_39946,N_38933,N_38611);
nor U39947 (N_39947,N_38790,N_38355);
and U39948 (N_39948,N_38937,N_38960);
xnor U39949 (N_39949,N_38449,N_38388);
and U39950 (N_39950,N_38429,N_38516);
or U39951 (N_39951,N_38971,N_38079);
or U39952 (N_39952,N_38442,N_38020);
nor U39953 (N_39953,N_38117,N_38846);
nor U39954 (N_39954,N_38444,N_38205);
and U39955 (N_39955,N_38151,N_38937);
nor U39956 (N_39956,N_38248,N_38162);
nand U39957 (N_39957,N_38476,N_38999);
and U39958 (N_39958,N_38781,N_38562);
and U39959 (N_39959,N_38401,N_38931);
nor U39960 (N_39960,N_38431,N_38813);
nand U39961 (N_39961,N_38648,N_38013);
nand U39962 (N_39962,N_38096,N_38517);
or U39963 (N_39963,N_38234,N_38042);
and U39964 (N_39964,N_38879,N_38677);
nand U39965 (N_39965,N_38759,N_38752);
nand U39966 (N_39966,N_38628,N_38490);
and U39967 (N_39967,N_38073,N_38198);
or U39968 (N_39968,N_38661,N_38808);
nor U39969 (N_39969,N_38585,N_38245);
nor U39970 (N_39970,N_38037,N_38992);
nand U39971 (N_39971,N_38750,N_38147);
xnor U39972 (N_39972,N_38743,N_38028);
xor U39973 (N_39973,N_38652,N_38454);
nand U39974 (N_39974,N_38033,N_38228);
and U39975 (N_39975,N_38777,N_38234);
and U39976 (N_39976,N_38606,N_38088);
or U39977 (N_39977,N_38027,N_38015);
or U39978 (N_39978,N_38828,N_38834);
and U39979 (N_39979,N_38116,N_38128);
nor U39980 (N_39980,N_38829,N_38685);
nor U39981 (N_39981,N_38190,N_38804);
or U39982 (N_39982,N_38614,N_38531);
and U39983 (N_39983,N_38752,N_38456);
nor U39984 (N_39984,N_38414,N_38987);
or U39985 (N_39985,N_38510,N_38298);
nand U39986 (N_39986,N_38423,N_38512);
nand U39987 (N_39987,N_38055,N_38674);
nor U39988 (N_39988,N_38539,N_38436);
xor U39989 (N_39989,N_38234,N_38261);
xnor U39990 (N_39990,N_38337,N_38380);
and U39991 (N_39991,N_38475,N_38148);
nand U39992 (N_39992,N_38503,N_38965);
xor U39993 (N_39993,N_38772,N_38623);
xor U39994 (N_39994,N_38350,N_38410);
nand U39995 (N_39995,N_38240,N_38372);
nor U39996 (N_39996,N_38658,N_38707);
and U39997 (N_39997,N_38728,N_38288);
or U39998 (N_39998,N_38572,N_38575);
xnor U39999 (N_39999,N_38909,N_38764);
or U40000 (N_40000,N_39713,N_39437);
and U40001 (N_40001,N_39551,N_39055);
or U40002 (N_40002,N_39368,N_39151);
xnor U40003 (N_40003,N_39159,N_39344);
or U40004 (N_40004,N_39334,N_39410);
or U40005 (N_40005,N_39757,N_39793);
xnor U40006 (N_40006,N_39518,N_39739);
xnor U40007 (N_40007,N_39163,N_39759);
nand U40008 (N_40008,N_39340,N_39767);
and U40009 (N_40009,N_39473,N_39036);
or U40010 (N_40010,N_39084,N_39046);
or U40011 (N_40011,N_39614,N_39965);
and U40012 (N_40012,N_39664,N_39376);
or U40013 (N_40013,N_39206,N_39169);
xnor U40014 (N_40014,N_39471,N_39958);
or U40015 (N_40015,N_39953,N_39364);
and U40016 (N_40016,N_39591,N_39773);
and U40017 (N_40017,N_39039,N_39835);
nor U40018 (N_40018,N_39384,N_39174);
and U40019 (N_40019,N_39913,N_39605);
xor U40020 (N_40020,N_39374,N_39354);
xor U40021 (N_40021,N_39843,N_39270);
xor U40022 (N_40022,N_39540,N_39312);
nor U40023 (N_40023,N_39910,N_39529);
xor U40024 (N_40024,N_39665,N_39610);
or U40025 (N_40025,N_39565,N_39634);
or U40026 (N_40026,N_39676,N_39099);
nand U40027 (N_40027,N_39620,N_39677);
or U40028 (N_40028,N_39592,N_39030);
xor U40029 (N_40029,N_39229,N_39337);
nand U40030 (N_40030,N_39395,N_39137);
or U40031 (N_40031,N_39183,N_39448);
or U40032 (N_40032,N_39116,N_39423);
or U40033 (N_40033,N_39222,N_39477);
nand U40034 (N_40034,N_39747,N_39542);
nor U40035 (N_40035,N_39837,N_39917);
nand U40036 (N_40036,N_39948,N_39988);
xnor U40037 (N_40037,N_39627,N_39916);
xor U40038 (N_40038,N_39439,N_39539);
nor U40039 (N_40039,N_39387,N_39889);
nor U40040 (N_40040,N_39295,N_39588);
and U40041 (N_40041,N_39708,N_39491);
xnor U40042 (N_40042,N_39027,N_39325);
nand U40043 (N_40043,N_39599,N_39303);
and U40044 (N_40044,N_39506,N_39981);
or U40045 (N_40045,N_39125,N_39904);
xor U40046 (N_40046,N_39050,N_39253);
and U40047 (N_40047,N_39435,N_39878);
nand U40048 (N_40048,N_39727,N_39755);
nand U40049 (N_40049,N_39353,N_39262);
nand U40050 (N_40050,N_39153,N_39968);
nand U40051 (N_40051,N_39771,N_39495);
xor U40052 (N_40052,N_39203,N_39415);
nand U40053 (N_40053,N_39121,N_39816);
or U40054 (N_40054,N_39626,N_39937);
xnor U40055 (N_40055,N_39310,N_39349);
nand U40056 (N_40056,N_39586,N_39649);
and U40057 (N_40057,N_39402,N_39556);
xor U40058 (N_40058,N_39386,N_39652);
xnor U40059 (N_40059,N_39298,N_39787);
xor U40060 (N_40060,N_39273,N_39081);
or U40061 (N_40061,N_39894,N_39447);
or U40062 (N_40062,N_39111,N_39500);
and U40063 (N_40063,N_39841,N_39182);
xnor U40064 (N_40064,N_39812,N_39356);
and U40065 (N_40065,N_39636,N_39552);
nor U40066 (N_40066,N_39064,N_39277);
xnor U40067 (N_40067,N_39230,N_39210);
nand U40068 (N_40068,N_39872,N_39839);
and U40069 (N_40069,N_39942,N_39146);
xnor U40070 (N_40070,N_39122,N_39257);
and U40071 (N_40071,N_39849,N_39493);
and U40072 (N_40072,N_39583,N_39675);
and U40073 (N_40073,N_39365,N_39989);
or U40074 (N_40074,N_39920,N_39091);
nor U40075 (N_40075,N_39044,N_39237);
or U40076 (N_40076,N_39720,N_39796);
nand U40077 (N_40077,N_39538,N_39287);
and U40078 (N_40078,N_39895,N_39212);
nor U40079 (N_40079,N_39969,N_39663);
xnor U40080 (N_40080,N_39993,N_39624);
xor U40081 (N_40081,N_39964,N_39528);
or U40082 (N_40082,N_39875,N_39670);
and U40083 (N_40083,N_39346,N_39221);
nand U40084 (N_40084,N_39827,N_39533);
nand U40085 (N_40085,N_39777,N_39840);
xor U40086 (N_40086,N_39233,N_39736);
and U40087 (N_40087,N_39289,N_39416);
or U40088 (N_40088,N_39975,N_39489);
nand U40089 (N_40089,N_39881,N_39095);
nand U40090 (N_40090,N_39004,N_39844);
and U40091 (N_40091,N_39074,N_39502);
and U40092 (N_40092,N_39286,N_39967);
nor U40093 (N_40093,N_39929,N_39276);
nand U40094 (N_40094,N_39445,N_39702);
nor U40095 (N_40095,N_39360,N_39255);
and U40096 (N_40096,N_39772,N_39687);
nand U40097 (N_40097,N_39077,N_39037);
xnor U40098 (N_40098,N_39355,N_39909);
nand U40099 (N_40099,N_39115,N_39748);
nor U40100 (N_40100,N_39570,N_39138);
xnor U40101 (N_40101,N_39654,N_39788);
nor U40102 (N_40102,N_39756,N_39826);
and U40103 (N_40103,N_39519,N_39723);
xor U40104 (N_40104,N_39080,N_39884);
and U40105 (N_40105,N_39347,N_39178);
xnor U40106 (N_40106,N_39822,N_39562);
nor U40107 (N_40107,N_39432,N_39530);
nand U40108 (N_40108,N_39087,N_39561);
xnor U40109 (N_40109,N_39361,N_39585);
nor U40110 (N_40110,N_39828,N_39877);
xor U40111 (N_40111,N_39836,N_39703);
nand U40112 (N_40112,N_39814,N_39128);
xor U40113 (N_40113,N_39243,N_39974);
and U40114 (N_40114,N_39631,N_39573);
and U40115 (N_40115,N_39874,N_39449);
or U40116 (N_40116,N_39526,N_39350);
and U40117 (N_40117,N_39200,N_39582);
nor U40118 (N_40118,N_39375,N_39228);
and U40119 (N_40119,N_39452,N_39770);
xor U40120 (N_40120,N_39763,N_39318);
or U40121 (N_40121,N_39392,N_39005);
and U40122 (N_40122,N_39504,N_39389);
nor U40123 (N_40123,N_39135,N_39003);
xor U40124 (N_40124,N_39915,N_39960);
or U40125 (N_40125,N_39420,N_39048);
or U40126 (N_40126,N_39862,N_39171);
nand U40127 (N_40127,N_39020,N_39443);
and U40128 (N_40128,N_39612,N_39054);
and U40129 (N_40129,N_39886,N_39780);
or U40130 (N_40130,N_39383,N_39083);
nand U40131 (N_40131,N_39370,N_39204);
xnor U40132 (N_40132,N_39069,N_39859);
and U40133 (N_40133,N_39335,N_39532);
nand U40134 (N_40134,N_39743,N_39806);
nor U40135 (N_40135,N_39424,N_39907);
xnor U40136 (N_40136,N_39319,N_39947);
xor U40137 (N_40137,N_39606,N_39934);
nor U40138 (N_40138,N_39466,N_39906);
and U40139 (N_40139,N_39161,N_39774);
and U40140 (N_40140,N_39341,N_39189);
or U40141 (N_40141,N_39698,N_39690);
or U40142 (N_40142,N_39683,N_39805);
xnor U40143 (N_40143,N_39290,N_39701);
and U40144 (N_40144,N_39870,N_39856);
nand U40145 (N_40145,N_39979,N_39052);
and U40146 (N_40146,N_39696,N_39944);
or U40147 (N_40147,N_39602,N_39730);
nand U40148 (N_40148,N_39411,N_39291);
xor U40149 (N_40149,N_39932,N_39373);
or U40150 (N_40150,N_39408,N_39486);
nand U40151 (N_40151,N_39184,N_39018);
nand U40152 (N_40152,N_39170,N_39598);
xnor U40153 (N_40153,N_39674,N_39945);
nor U40154 (N_40154,N_39852,N_39242);
and U40155 (N_40155,N_39363,N_39085);
nor U40156 (N_40156,N_39244,N_39129);
and U40157 (N_40157,N_39110,N_39563);
and U40158 (N_40158,N_39008,N_39750);
or U40159 (N_40159,N_39226,N_39301);
nor U40160 (N_40160,N_39023,N_39499);
nor U40161 (N_40161,N_39554,N_39235);
or U40162 (N_40162,N_39729,N_39791);
and U40163 (N_40163,N_39428,N_39014);
or U40164 (N_40164,N_39058,N_39818);
and U40165 (N_40165,N_39625,N_39234);
and U40166 (N_40166,N_39430,N_39149);
xnor U40167 (N_40167,N_39133,N_39745);
xor U40168 (N_40168,N_39879,N_39207);
nand U40169 (N_40169,N_39692,N_39336);
and U40170 (N_40170,N_39996,N_39117);
nand U40171 (N_40171,N_39684,N_39062);
nor U40172 (N_40172,N_39810,N_39710);
or U40173 (N_40173,N_39901,N_39550);
nand U40174 (N_40174,N_39302,N_39555);
or U40175 (N_40175,N_39782,N_39279);
or U40176 (N_40176,N_39959,N_39446);
and U40177 (N_40177,N_39327,N_39558);
xnor U40178 (N_40178,N_39362,N_39266);
xor U40179 (N_40179,N_39637,N_39492);
and U40180 (N_40180,N_39646,N_39594);
xnor U40181 (N_40181,N_39762,N_39673);
and U40182 (N_40182,N_39078,N_39863);
or U40183 (N_40183,N_39481,N_39127);
and U40184 (N_40184,N_39623,N_39864);
and U40185 (N_40185,N_39735,N_39609);
nor U40186 (N_40186,N_39268,N_39847);
and U40187 (N_40187,N_39248,N_39956);
xor U40188 (N_40188,N_39199,N_39431);
nand U40189 (N_40189,N_39914,N_39966);
or U40190 (N_40190,N_39019,N_39119);
nor U40191 (N_40191,N_39214,N_39453);
and U40192 (N_40192,N_39524,N_39441);
nor U40193 (N_40193,N_39622,N_39252);
nand U40194 (N_40194,N_39267,N_39366);
and U40195 (N_40195,N_39977,N_39067);
or U40196 (N_40196,N_39240,N_39114);
xnor U40197 (N_40197,N_39971,N_39391);
nor U40198 (N_40198,N_39457,N_39783);
nand U40199 (N_40199,N_39196,N_39845);
nand U40200 (N_40200,N_39296,N_39485);
nand U40201 (N_40201,N_39725,N_39854);
xor U40202 (N_40202,N_39232,N_39154);
or U40203 (N_40203,N_39919,N_39251);
nand U40204 (N_40204,N_39238,N_39106);
nor U40205 (N_40205,N_39160,N_39574);
nor U40206 (N_40206,N_39463,N_39292);
nand U40207 (N_40207,N_39145,N_39792);
and U40208 (N_40208,N_39313,N_39032);
nand U40209 (N_40209,N_39508,N_39413);
xor U40210 (N_40210,N_39258,N_39132);
nand U40211 (N_40211,N_39501,N_39165);
nand U40212 (N_40212,N_39850,N_39738);
nor U40213 (N_40213,N_39824,N_39175);
nand U40214 (N_40214,N_39089,N_39997);
xnor U40215 (N_40215,N_39923,N_39579);
nand U40216 (N_40216,N_39007,N_39459);
and U40217 (N_40217,N_39825,N_39815);
xor U40218 (N_40218,N_39247,N_39728);
or U40219 (N_40219,N_39417,N_39926);
xnor U40220 (N_40220,N_39231,N_39903);
nand U40221 (N_40221,N_39571,N_39168);
nand U40222 (N_40222,N_39543,N_39741);
nor U40223 (N_40223,N_39568,N_39525);
nor U40224 (N_40224,N_39744,N_39754);
xnor U40225 (N_40225,N_39405,N_39998);
or U40226 (N_40226,N_39891,N_39288);
nor U40227 (N_40227,N_39666,N_39976);
or U40228 (N_40228,N_39628,N_39250);
and U40229 (N_40229,N_39208,N_39643);
nor U40230 (N_40230,N_39227,N_39015);
nor U40231 (N_40231,N_39479,N_39141);
xor U40232 (N_40232,N_39320,N_39412);
xnor U40233 (N_40233,N_39790,N_39470);
or U40234 (N_40234,N_39496,N_39322);
xnor U40235 (N_40235,N_39461,N_39642);
xnor U40236 (N_40236,N_39660,N_39779);
nor U40237 (N_40237,N_39326,N_39982);
nor U40238 (N_40238,N_39217,N_39472);
nand U40239 (N_40239,N_39398,N_39704);
nor U40240 (N_40240,N_39331,N_39930);
xnor U40241 (N_40241,N_39075,N_39809);
or U40242 (N_40242,N_39686,N_39180);
and U40243 (N_40243,N_39716,N_39404);
nand U40244 (N_40244,N_39369,N_39333);
nand U40245 (N_40245,N_39581,N_39195);
xor U40246 (N_40246,N_39865,N_39259);
and U40247 (N_40247,N_39002,N_39509);
and U40248 (N_40248,N_39962,N_39681);
nor U40249 (N_40249,N_39882,N_39522);
and U40250 (N_40250,N_39892,N_39359);
nand U40251 (N_40251,N_39109,N_39173);
nor U40252 (N_40252,N_39324,N_39980);
nor U40253 (N_40253,N_39742,N_39752);
and U40254 (N_40254,N_39456,N_39450);
and U40255 (N_40255,N_39672,N_39143);
or U40256 (N_40256,N_39158,N_39406);
xnor U40257 (N_40257,N_39534,N_39871);
nor U40258 (N_40258,N_39300,N_39639);
and U40259 (N_40259,N_39352,N_39523);
and U40260 (N_40260,N_39600,N_39434);
nand U40261 (N_40261,N_39897,N_39507);
or U40262 (N_40262,N_39475,N_39024);
nand U40263 (N_40263,N_39147,N_39070);
nor U40264 (N_40264,N_39943,N_39283);
xor U40265 (N_40265,N_39541,N_39516);
or U40266 (N_40266,N_39724,N_39224);
xor U40267 (N_40267,N_39063,N_39113);
nand U40268 (N_40268,N_39700,N_39469);
nand U40269 (N_40269,N_39096,N_39604);
or U40270 (N_40270,N_39817,N_39394);
xor U40271 (N_40271,N_39611,N_39401);
nor U40272 (N_40272,N_39407,N_39607);
nor U40273 (N_40273,N_39821,N_39108);
nand U40274 (N_40274,N_39297,N_39732);
nor U40275 (N_40275,N_39576,N_39963);
nor U40276 (N_40276,N_39832,N_39902);
nand U40277 (N_40277,N_39060,N_39131);
nand U40278 (N_40278,N_39427,N_39645);
nand U40279 (N_40279,N_39876,N_39454);
nand U40280 (N_40280,N_39807,N_39991);
and U40281 (N_40281,N_39465,N_39329);
and U40282 (N_40282,N_39549,N_39572);
or U40283 (N_40283,N_39808,N_39927);
xnor U40284 (N_40284,N_39088,N_39487);
xor U40285 (N_40285,N_39223,N_39012);
xnor U40286 (N_40286,N_39397,N_39630);
and U40287 (N_40287,N_39601,N_39462);
nor U40288 (N_40288,N_39236,N_39198);
xnor U40289 (N_40289,N_39544,N_39651);
or U40290 (N_40290,N_39474,N_39853);
nand U40291 (N_40291,N_39633,N_39488);
and U40292 (N_40292,N_39436,N_39179);
nor U40293 (N_40293,N_39194,N_39061);
and U40294 (N_40294,N_39995,N_39090);
nor U40295 (N_40295,N_39079,N_39668);
or U40296 (N_40296,N_39490,N_39635);
nand U40297 (N_40297,N_39925,N_39804);
or U40298 (N_40298,N_39899,N_39564);
and U40299 (N_40299,N_39107,N_39380);
xnor U40300 (N_40300,N_39714,N_39972);
xnor U40301 (N_40301,N_39045,N_39464);
nor U40302 (N_40302,N_39120,N_39712);
xnor U40303 (N_40303,N_39043,N_39987);
and U40304 (N_40304,N_39990,N_39304);
nand U40305 (N_40305,N_39935,N_39315);
and U40306 (N_40306,N_39803,N_39749);
xor U40307 (N_40307,N_39597,N_39072);
or U40308 (N_40308,N_39284,N_39101);
nand U40309 (N_40309,N_39418,N_39647);
xor U40310 (N_40310,N_39802,N_39890);
and U40311 (N_40311,N_39688,N_39188);
and U40312 (N_40312,N_39309,N_39799);
nand U40313 (N_40313,N_39112,N_39444);
or U40314 (N_40314,N_39691,N_39265);
or U40315 (N_40315,N_39136,N_39467);
nor U40316 (N_40316,N_39706,N_39868);
and U40317 (N_40317,N_39699,N_39225);
xnor U40318 (N_40318,N_39896,N_39928);
or U40319 (N_40319,N_39952,N_39123);
and U40320 (N_40320,N_39026,N_39775);
or U40321 (N_40321,N_39164,N_39984);
nor U40322 (N_40322,N_39105,N_39264);
nand U40323 (N_40323,N_39789,N_39484);
xor U40324 (N_40324,N_39280,N_39396);
xor U40325 (N_40325,N_39314,N_39669);
or U40326 (N_40326,N_39505,N_39186);
nor U40327 (N_40327,N_39241,N_39177);
or U40328 (N_40328,N_39831,N_39946);
nand U40329 (N_40329,N_39883,N_39321);
and U40330 (N_40330,N_39721,N_39753);
xnor U40331 (N_40331,N_39098,N_39857);
xnor U40332 (N_40332,N_39587,N_39185);
nand U40333 (N_40333,N_39269,N_39051);
or U40334 (N_40334,N_39671,N_39261);
or U40335 (N_40335,N_39388,N_39076);
xor U40336 (N_40336,N_39617,N_39094);
nor U40337 (N_40337,N_39000,N_39093);
and U40338 (N_40338,N_39371,N_39794);
nand U40339 (N_40339,N_39978,N_39695);
and U40340 (N_40340,N_39476,N_39851);
xnor U40341 (N_40341,N_39367,N_39148);
xor U40342 (N_40342,N_39842,N_39343);
or U40343 (N_40343,N_39033,N_39042);
nor U40344 (N_40344,N_39577,N_39377);
nor U40345 (N_40345,N_39955,N_39468);
and U40346 (N_40346,N_39211,N_39103);
or U40347 (N_40347,N_39118,N_39025);
nor U40348 (N_40348,N_39679,N_39438);
xnor U40349 (N_40349,N_39379,N_39278);
nor U40350 (N_40350,N_39536,N_39954);
and U40351 (N_40351,N_39905,N_39678);
and U40352 (N_40352,N_39393,N_39339);
and U40353 (N_40353,N_39140,N_39097);
xor U40354 (N_40354,N_39766,N_39992);
nor U40355 (N_40355,N_39722,N_39419);
or U40356 (N_40356,N_39869,N_39442);
and U40357 (N_40357,N_39848,N_39527);
nand U40358 (N_40358,N_39066,N_39638);
xor U40359 (N_40359,N_39192,N_39323);
or U40360 (N_40360,N_39281,N_39205);
nand U40361 (N_40361,N_39545,N_39658);
nor U40362 (N_40362,N_39734,N_39068);
or U40363 (N_40363,N_39034,N_39460);
xnor U40364 (N_40364,N_39422,N_39440);
or U40365 (N_40365,N_39483,N_39838);
nand U40366 (N_40366,N_39006,N_39908);
xor U40367 (N_40367,N_39941,N_39342);
nand U40368 (N_40368,N_39260,N_39715);
xnor U40369 (N_40369,N_39918,N_39559);
nor U40370 (N_40370,N_39245,N_39239);
xor U40371 (N_40371,N_39768,N_39820);
or U40372 (N_40372,N_39167,N_39781);
and U40373 (N_40373,N_39653,N_39059);
nand U40374 (N_40374,N_39390,N_39911);
or U40375 (N_40375,N_39694,N_39589);
and U40376 (N_40376,N_39846,N_39615);
and U40377 (N_40377,N_39640,N_39275);
nor U40378 (N_40378,N_39162,N_39001);
nand U40379 (N_40379,N_39073,N_39049);
nor U40380 (N_40380,N_39433,N_39961);
xor U40381 (N_40381,N_39256,N_39022);
nand U40382 (N_40382,N_39578,N_39512);
nor U40383 (N_40383,N_39482,N_39065);
or U40384 (N_40384,N_39834,N_39426);
nor U40385 (N_40385,N_39662,N_39813);
nand U40386 (N_40386,N_39784,N_39209);
nor U40387 (N_40387,N_39866,N_39801);
nor U40388 (N_40388,N_39880,N_39451);
xor U40389 (N_40389,N_39421,N_39731);
and U40390 (N_40390,N_39938,N_39888);
nor U40391 (N_40391,N_39086,N_39861);
xnor U40392 (N_40392,N_39893,N_39299);
and U40393 (N_40393,N_39317,N_39566);
nor U40394 (N_40394,N_39197,N_39307);
and U40395 (N_40395,N_39282,N_39659);
nand U40396 (N_40396,N_39800,N_39029);
and U40397 (N_40397,N_39621,N_39717);
or U40398 (N_40398,N_39017,N_39590);
and U40399 (N_40399,N_39316,N_39358);
nor U40400 (N_40400,N_39176,N_39092);
or U40401 (N_40401,N_39414,N_39330);
nor U40402 (N_40402,N_39553,N_39013);
nand U40403 (N_40403,N_39521,N_39994);
xnor U40404 (N_40404,N_39758,N_39648);
nor U40405 (N_40405,N_39219,N_39053);
nor U40406 (N_40406,N_39458,N_39513);
nor U40407 (N_40407,N_39047,N_39973);
nand U40408 (N_40408,N_39797,N_39760);
xnor U40409 (N_40409,N_39510,N_39011);
nor U40410 (N_40410,N_39102,N_39274);
nor U40411 (N_40411,N_39385,N_39021);
or U40412 (N_40412,N_39616,N_39305);
nand U40413 (N_40413,N_39531,N_39503);
nand U40414 (N_40414,N_39557,N_39795);
nor U40415 (N_40415,N_39035,N_39372);
nand U40416 (N_40416,N_39139,N_39520);
nor U40417 (N_40417,N_39682,N_39951);
and U40418 (N_40418,N_39400,N_39709);
nand U40419 (N_40419,N_39740,N_39546);
or U40420 (N_40420,N_39608,N_39056);
or U40421 (N_40421,N_39986,N_39381);
and U40422 (N_40422,N_39294,N_39511);
nor U40423 (N_40423,N_39595,N_39833);
nor U40424 (N_40424,N_39898,N_39629);
and U40425 (N_40425,N_39429,N_39764);
nor U40426 (N_40426,N_39497,N_39498);
and U40427 (N_40427,N_39357,N_39547);
xnor U40428 (N_40428,N_39560,N_39746);
or U40429 (N_40429,N_39737,N_39348);
nor U40430 (N_40430,N_39830,N_39921);
and U40431 (N_40431,N_39191,N_39705);
nor U40432 (N_40432,N_39201,N_39769);
nor U40433 (N_40433,N_39776,N_39071);
xnor U40434 (N_40434,N_39970,N_39272);
or U40435 (N_40435,N_39580,N_39811);
nor U40436 (N_40436,N_39718,N_39328);
nor U40437 (N_40437,N_39693,N_39765);
xor U40438 (N_40438,N_39761,N_39306);
and U40439 (N_40439,N_39220,N_39514);
or U40440 (N_40440,N_39213,N_39922);
or U40441 (N_40441,N_39829,N_39040);
xor U40442 (N_40442,N_39172,N_39798);
nor U40443 (N_40443,N_39190,N_39985);
or U40444 (N_40444,N_39537,N_39569);
or U40445 (N_40445,N_39887,N_39719);
nor U40446 (N_40446,N_39936,N_39455);
and U40447 (N_40447,N_39517,N_39819);
xnor U40448 (N_40448,N_39254,N_39409);
and U40449 (N_40449,N_39480,N_39939);
and U40450 (N_40450,N_39478,N_39010);
nand U40451 (N_40451,N_39785,N_39038);
and U40452 (N_40452,N_39641,N_39009);
and U40453 (N_40453,N_39931,N_39940);
and U40454 (N_40454,N_39656,N_39249);
nand U40455 (N_40455,N_39285,N_39613);
nor U40456 (N_40456,N_39382,N_39166);
or U40457 (N_40457,N_39271,N_39603);
xnor U40458 (N_40458,N_39104,N_39150);
nor U40459 (N_40459,N_39751,N_39155);
nand U40460 (N_40460,N_39332,N_39134);
or U40461 (N_40461,N_39144,N_39733);
or U40462 (N_40462,N_39858,N_39100);
nor U40463 (N_40463,N_39425,N_39082);
and U40464 (N_40464,N_39657,N_39293);
nand U40465 (N_40465,N_39697,N_39156);
and U40466 (N_40466,N_39855,N_39584);
or U40467 (N_40467,N_39644,N_39957);
and U40468 (N_40468,N_39823,N_39707);
or U40469 (N_40469,N_39596,N_39667);
nand U40470 (N_40470,N_39057,N_39263);
nand U40471 (N_40471,N_39567,N_39786);
or U40472 (N_40472,N_39193,N_39535);
or U40473 (N_40473,N_39650,N_39950);
nand U40474 (N_40474,N_39548,N_39593);
nand U40475 (N_40475,N_39933,N_39181);
nand U40476 (N_40476,N_39403,N_39126);
and U40477 (N_40477,N_39311,N_39632);
xor U40478 (N_40478,N_39202,N_39999);
nor U40479 (N_40479,N_39778,N_39028);
nor U40480 (N_40480,N_39661,N_39885);
nor U40481 (N_40481,N_39351,N_39860);
and U40482 (N_40482,N_39900,N_39152);
nand U40483 (N_40483,N_39124,N_39726);
nand U40484 (N_40484,N_39399,N_39308);
nor U40485 (N_40485,N_39618,N_39912);
or U40486 (N_40486,N_39575,N_39031);
nor U40487 (N_40487,N_39378,N_39142);
nand U40488 (N_40488,N_39345,N_39187);
nor U40489 (N_40489,N_39949,N_39867);
xnor U40490 (N_40490,N_39873,N_39685);
nor U40491 (N_40491,N_39130,N_39983);
xnor U40492 (N_40492,N_39246,N_39680);
and U40493 (N_40493,N_39157,N_39218);
xor U40494 (N_40494,N_39655,N_39016);
nand U40495 (N_40495,N_39689,N_39041);
or U40496 (N_40496,N_39338,N_39215);
nor U40497 (N_40497,N_39515,N_39711);
and U40498 (N_40498,N_39924,N_39216);
nor U40499 (N_40499,N_39494,N_39619);
or U40500 (N_40500,N_39577,N_39124);
xnor U40501 (N_40501,N_39363,N_39516);
xor U40502 (N_40502,N_39244,N_39587);
xor U40503 (N_40503,N_39772,N_39946);
nand U40504 (N_40504,N_39700,N_39273);
xor U40505 (N_40505,N_39954,N_39290);
nand U40506 (N_40506,N_39741,N_39083);
or U40507 (N_40507,N_39837,N_39501);
or U40508 (N_40508,N_39063,N_39700);
and U40509 (N_40509,N_39282,N_39224);
or U40510 (N_40510,N_39908,N_39359);
and U40511 (N_40511,N_39542,N_39900);
or U40512 (N_40512,N_39964,N_39393);
nand U40513 (N_40513,N_39106,N_39879);
xor U40514 (N_40514,N_39825,N_39691);
nor U40515 (N_40515,N_39337,N_39018);
xnor U40516 (N_40516,N_39263,N_39553);
and U40517 (N_40517,N_39304,N_39596);
or U40518 (N_40518,N_39941,N_39250);
nand U40519 (N_40519,N_39875,N_39859);
xor U40520 (N_40520,N_39148,N_39792);
or U40521 (N_40521,N_39767,N_39385);
xnor U40522 (N_40522,N_39495,N_39324);
and U40523 (N_40523,N_39371,N_39800);
and U40524 (N_40524,N_39857,N_39600);
nor U40525 (N_40525,N_39369,N_39279);
nand U40526 (N_40526,N_39029,N_39310);
xnor U40527 (N_40527,N_39006,N_39819);
nand U40528 (N_40528,N_39802,N_39797);
or U40529 (N_40529,N_39112,N_39365);
nor U40530 (N_40530,N_39089,N_39980);
or U40531 (N_40531,N_39416,N_39332);
or U40532 (N_40532,N_39482,N_39001);
xnor U40533 (N_40533,N_39405,N_39714);
xor U40534 (N_40534,N_39925,N_39068);
nand U40535 (N_40535,N_39945,N_39066);
nand U40536 (N_40536,N_39599,N_39001);
and U40537 (N_40537,N_39533,N_39377);
nor U40538 (N_40538,N_39185,N_39914);
and U40539 (N_40539,N_39447,N_39053);
and U40540 (N_40540,N_39658,N_39966);
xnor U40541 (N_40541,N_39806,N_39273);
xnor U40542 (N_40542,N_39183,N_39064);
or U40543 (N_40543,N_39739,N_39441);
or U40544 (N_40544,N_39623,N_39232);
nor U40545 (N_40545,N_39136,N_39762);
nand U40546 (N_40546,N_39744,N_39405);
nand U40547 (N_40547,N_39630,N_39987);
or U40548 (N_40548,N_39349,N_39812);
nand U40549 (N_40549,N_39529,N_39113);
or U40550 (N_40550,N_39967,N_39190);
nor U40551 (N_40551,N_39564,N_39797);
nor U40552 (N_40552,N_39740,N_39584);
xnor U40553 (N_40553,N_39279,N_39977);
nor U40554 (N_40554,N_39858,N_39467);
nor U40555 (N_40555,N_39710,N_39258);
and U40556 (N_40556,N_39869,N_39921);
nor U40557 (N_40557,N_39532,N_39907);
nand U40558 (N_40558,N_39058,N_39575);
xnor U40559 (N_40559,N_39951,N_39960);
or U40560 (N_40560,N_39163,N_39722);
xnor U40561 (N_40561,N_39359,N_39091);
nor U40562 (N_40562,N_39829,N_39058);
xnor U40563 (N_40563,N_39433,N_39322);
and U40564 (N_40564,N_39038,N_39264);
nor U40565 (N_40565,N_39236,N_39798);
and U40566 (N_40566,N_39476,N_39818);
and U40567 (N_40567,N_39398,N_39128);
nand U40568 (N_40568,N_39757,N_39404);
and U40569 (N_40569,N_39058,N_39352);
nand U40570 (N_40570,N_39537,N_39589);
or U40571 (N_40571,N_39270,N_39148);
nor U40572 (N_40572,N_39732,N_39944);
or U40573 (N_40573,N_39357,N_39088);
or U40574 (N_40574,N_39631,N_39749);
xnor U40575 (N_40575,N_39401,N_39248);
or U40576 (N_40576,N_39847,N_39685);
nor U40577 (N_40577,N_39435,N_39478);
and U40578 (N_40578,N_39700,N_39961);
nor U40579 (N_40579,N_39858,N_39985);
nor U40580 (N_40580,N_39737,N_39722);
nor U40581 (N_40581,N_39955,N_39385);
and U40582 (N_40582,N_39750,N_39838);
or U40583 (N_40583,N_39727,N_39367);
nor U40584 (N_40584,N_39542,N_39175);
nor U40585 (N_40585,N_39403,N_39659);
or U40586 (N_40586,N_39956,N_39597);
and U40587 (N_40587,N_39651,N_39123);
nor U40588 (N_40588,N_39692,N_39541);
nand U40589 (N_40589,N_39227,N_39055);
xnor U40590 (N_40590,N_39706,N_39166);
and U40591 (N_40591,N_39180,N_39988);
xnor U40592 (N_40592,N_39210,N_39992);
and U40593 (N_40593,N_39585,N_39125);
nand U40594 (N_40594,N_39045,N_39895);
and U40595 (N_40595,N_39016,N_39113);
or U40596 (N_40596,N_39385,N_39831);
nor U40597 (N_40597,N_39414,N_39169);
xnor U40598 (N_40598,N_39107,N_39569);
nand U40599 (N_40599,N_39660,N_39009);
nor U40600 (N_40600,N_39815,N_39286);
or U40601 (N_40601,N_39263,N_39227);
nand U40602 (N_40602,N_39528,N_39159);
and U40603 (N_40603,N_39206,N_39811);
or U40604 (N_40604,N_39740,N_39730);
xnor U40605 (N_40605,N_39526,N_39739);
nand U40606 (N_40606,N_39208,N_39702);
xnor U40607 (N_40607,N_39174,N_39683);
or U40608 (N_40608,N_39396,N_39958);
and U40609 (N_40609,N_39791,N_39526);
or U40610 (N_40610,N_39530,N_39743);
nor U40611 (N_40611,N_39606,N_39514);
and U40612 (N_40612,N_39959,N_39852);
nand U40613 (N_40613,N_39941,N_39695);
nand U40614 (N_40614,N_39326,N_39929);
nand U40615 (N_40615,N_39291,N_39267);
and U40616 (N_40616,N_39123,N_39865);
xor U40617 (N_40617,N_39113,N_39766);
xnor U40618 (N_40618,N_39588,N_39280);
nor U40619 (N_40619,N_39369,N_39103);
nand U40620 (N_40620,N_39157,N_39906);
xnor U40621 (N_40621,N_39461,N_39991);
and U40622 (N_40622,N_39714,N_39689);
xnor U40623 (N_40623,N_39930,N_39038);
or U40624 (N_40624,N_39122,N_39937);
and U40625 (N_40625,N_39828,N_39873);
nor U40626 (N_40626,N_39224,N_39455);
nand U40627 (N_40627,N_39332,N_39529);
and U40628 (N_40628,N_39320,N_39610);
xnor U40629 (N_40629,N_39248,N_39203);
or U40630 (N_40630,N_39984,N_39344);
and U40631 (N_40631,N_39976,N_39903);
and U40632 (N_40632,N_39967,N_39928);
nand U40633 (N_40633,N_39930,N_39937);
nand U40634 (N_40634,N_39345,N_39098);
or U40635 (N_40635,N_39452,N_39082);
or U40636 (N_40636,N_39883,N_39427);
xnor U40637 (N_40637,N_39156,N_39195);
nand U40638 (N_40638,N_39297,N_39287);
or U40639 (N_40639,N_39193,N_39846);
and U40640 (N_40640,N_39479,N_39686);
nand U40641 (N_40641,N_39626,N_39950);
xor U40642 (N_40642,N_39468,N_39010);
nor U40643 (N_40643,N_39683,N_39723);
xnor U40644 (N_40644,N_39868,N_39385);
or U40645 (N_40645,N_39986,N_39281);
nor U40646 (N_40646,N_39153,N_39926);
nand U40647 (N_40647,N_39232,N_39772);
nand U40648 (N_40648,N_39601,N_39861);
or U40649 (N_40649,N_39880,N_39823);
nor U40650 (N_40650,N_39145,N_39462);
and U40651 (N_40651,N_39824,N_39271);
nand U40652 (N_40652,N_39066,N_39433);
or U40653 (N_40653,N_39989,N_39579);
or U40654 (N_40654,N_39355,N_39252);
nand U40655 (N_40655,N_39793,N_39584);
nand U40656 (N_40656,N_39809,N_39431);
nor U40657 (N_40657,N_39195,N_39593);
nand U40658 (N_40658,N_39332,N_39090);
or U40659 (N_40659,N_39828,N_39237);
xor U40660 (N_40660,N_39189,N_39919);
or U40661 (N_40661,N_39342,N_39683);
and U40662 (N_40662,N_39128,N_39318);
and U40663 (N_40663,N_39010,N_39743);
or U40664 (N_40664,N_39950,N_39816);
or U40665 (N_40665,N_39322,N_39983);
nand U40666 (N_40666,N_39400,N_39961);
and U40667 (N_40667,N_39037,N_39752);
nor U40668 (N_40668,N_39893,N_39253);
nor U40669 (N_40669,N_39834,N_39300);
nor U40670 (N_40670,N_39546,N_39625);
nand U40671 (N_40671,N_39658,N_39958);
nand U40672 (N_40672,N_39778,N_39223);
or U40673 (N_40673,N_39843,N_39041);
and U40674 (N_40674,N_39607,N_39062);
nor U40675 (N_40675,N_39335,N_39391);
nor U40676 (N_40676,N_39251,N_39380);
nor U40677 (N_40677,N_39032,N_39010);
nand U40678 (N_40678,N_39655,N_39093);
or U40679 (N_40679,N_39734,N_39213);
nand U40680 (N_40680,N_39400,N_39391);
xor U40681 (N_40681,N_39716,N_39028);
nand U40682 (N_40682,N_39405,N_39976);
or U40683 (N_40683,N_39767,N_39957);
xnor U40684 (N_40684,N_39695,N_39267);
and U40685 (N_40685,N_39014,N_39077);
xor U40686 (N_40686,N_39693,N_39507);
nor U40687 (N_40687,N_39859,N_39187);
xor U40688 (N_40688,N_39767,N_39527);
and U40689 (N_40689,N_39762,N_39683);
or U40690 (N_40690,N_39514,N_39394);
or U40691 (N_40691,N_39202,N_39626);
nand U40692 (N_40692,N_39478,N_39511);
nor U40693 (N_40693,N_39347,N_39629);
and U40694 (N_40694,N_39919,N_39826);
xnor U40695 (N_40695,N_39198,N_39947);
nand U40696 (N_40696,N_39427,N_39243);
xor U40697 (N_40697,N_39512,N_39339);
or U40698 (N_40698,N_39406,N_39003);
and U40699 (N_40699,N_39601,N_39238);
and U40700 (N_40700,N_39099,N_39068);
or U40701 (N_40701,N_39002,N_39071);
and U40702 (N_40702,N_39704,N_39737);
nor U40703 (N_40703,N_39686,N_39703);
or U40704 (N_40704,N_39192,N_39419);
nand U40705 (N_40705,N_39743,N_39203);
nand U40706 (N_40706,N_39323,N_39509);
nand U40707 (N_40707,N_39546,N_39690);
and U40708 (N_40708,N_39759,N_39627);
and U40709 (N_40709,N_39932,N_39804);
nor U40710 (N_40710,N_39323,N_39024);
nand U40711 (N_40711,N_39812,N_39624);
nor U40712 (N_40712,N_39231,N_39791);
and U40713 (N_40713,N_39599,N_39549);
nor U40714 (N_40714,N_39297,N_39286);
nor U40715 (N_40715,N_39749,N_39409);
or U40716 (N_40716,N_39082,N_39887);
nor U40717 (N_40717,N_39260,N_39151);
nor U40718 (N_40718,N_39898,N_39884);
nor U40719 (N_40719,N_39789,N_39699);
nor U40720 (N_40720,N_39807,N_39221);
and U40721 (N_40721,N_39629,N_39060);
or U40722 (N_40722,N_39321,N_39305);
and U40723 (N_40723,N_39442,N_39879);
nor U40724 (N_40724,N_39763,N_39739);
xor U40725 (N_40725,N_39510,N_39987);
nor U40726 (N_40726,N_39841,N_39814);
nor U40727 (N_40727,N_39373,N_39039);
nand U40728 (N_40728,N_39982,N_39745);
or U40729 (N_40729,N_39436,N_39690);
and U40730 (N_40730,N_39096,N_39567);
xnor U40731 (N_40731,N_39249,N_39578);
xor U40732 (N_40732,N_39630,N_39215);
and U40733 (N_40733,N_39435,N_39966);
and U40734 (N_40734,N_39416,N_39240);
nand U40735 (N_40735,N_39247,N_39469);
xor U40736 (N_40736,N_39457,N_39361);
xor U40737 (N_40737,N_39146,N_39332);
or U40738 (N_40738,N_39784,N_39271);
or U40739 (N_40739,N_39920,N_39813);
and U40740 (N_40740,N_39128,N_39419);
nor U40741 (N_40741,N_39187,N_39613);
xor U40742 (N_40742,N_39355,N_39284);
xor U40743 (N_40743,N_39389,N_39051);
nand U40744 (N_40744,N_39578,N_39605);
and U40745 (N_40745,N_39418,N_39199);
xnor U40746 (N_40746,N_39294,N_39236);
or U40747 (N_40747,N_39451,N_39219);
xor U40748 (N_40748,N_39465,N_39306);
nor U40749 (N_40749,N_39075,N_39275);
xnor U40750 (N_40750,N_39888,N_39806);
or U40751 (N_40751,N_39716,N_39558);
and U40752 (N_40752,N_39460,N_39780);
nand U40753 (N_40753,N_39093,N_39986);
xnor U40754 (N_40754,N_39383,N_39447);
nor U40755 (N_40755,N_39144,N_39517);
and U40756 (N_40756,N_39831,N_39490);
xor U40757 (N_40757,N_39964,N_39221);
nor U40758 (N_40758,N_39752,N_39541);
or U40759 (N_40759,N_39884,N_39192);
nor U40760 (N_40760,N_39906,N_39813);
and U40761 (N_40761,N_39473,N_39504);
nor U40762 (N_40762,N_39720,N_39073);
nand U40763 (N_40763,N_39380,N_39924);
nor U40764 (N_40764,N_39557,N_39902);
nand U40765 (N_40765,N_39866,N_39216);
nor U40766 (N_40766,N_39297,N_39860);
xor U40767 (N_40767,N_39026,N_39133);
xnor U40768 (N_40768,N_39334,N_39975);
or U40769 (N_40769,N_39583,N_39369);
nand U40770 (N_40770,N_39005,N_39391);
or U40771 (N_40771,N_39038,N_39344);
and U40772 (N_40772,N_39037,N_39183);
and U40773 (N_40773,N_39518,N_39318);
nor U40774 (N_40774,N_39751,N_39821);
xnor U40775 (N_40775,N_39241,N_39769);
xor U40776 (N_40776,N_39816,N_39051);
or U40777 (N_40777,N_39769,N_39811);
nor U40778 (N_40778,N_39176,N_39429);
and U40779 (N_40779,N_39247,N_39113);
nand U40780 (N_40780,N_39655,N_39320);
xor U40781 (N_40781,N_39769,N_39049);
xor U40782 (N_40782,N_39228,N_39942);
or U40783 (N_40783,N_39925,N_39266);
and U40784 (N_40784,N_39929,N_39120);
xor U40785 (N_40785,N_39089,N_39966);
xnor U40786 (N_40786,N_39187,N_39163);
or U40787 (N_40787,N_39468,N_39855);
and U40788 (N_40788,N_39532,N_39443);
and U40789 (N_40789,N_39040,N_39281);
and U40790 (N_40790,N_39660,N_39256);
xor U40791 (N_40791,N_39459,N_39864);
and U40792 (N_40792,N_39729,N_39868);
nor U40793 (N_40793,N_39339,N_39182);
xor U40794 (N_40794,N_39641,N_39939);
and U40795 (N_40795,N_39459,N_39033);
nand U40796 (N_40796,N_39551,N_39433);
nor U40797 (N_40797,N_39355,N_39681);
nor U40798 (N_40798,N_39059,N_39979);
or U40799 (N_40799,N_39111,N_39470);
and U40800 (N_40800,N_39953,N_39797);
nor U40801 (N_40801,N_39071,N_39365);
nand U40802 (N_40802,N_39559,N_39679);
nand U40803 (N_40803,N_39538,N_39637);
nand U40804 (N_40804,N_39338,N_39876);
nand U40805 (N_40805,N_39425,N_39063);
or U40806 (N_40806,N_39127,N_39322);
nand U40807 (N_40807,N_39896,N_39431);
or U40808 (N_40808,N_39533,N_39574);
xor U40809 (N_40809,N_39335,N_39737);
nor U40810 (N_40810,N_39485,N_39591);
xor U40811 (N_40811,N_39140,N_39633);
nor U40812 (N_40812,N_39745,N_39271);
or U40813 (N_40813,N_39596,N_39333);
or U40814 (N_40814,N_39512,N_39336);
xor U40815 (N_40815,N_39938,N_39064);
or U40816 (N_40816,N_39649,N_39143);
and U40817 (N_40817,N_39620,N_39838);
nor U40818 (N_40818,N_39411,N_39991);
nand U40819 (N_40819,N_39478,N_39692);
or U40820 (N_40820,N_39659,N_39139);
nor U40821 (N_40821,N_39686,N_39942);
and U40822 (N_40822,N_39864,N_39611);
or U40823 (N_40823,N_39546,N_39764);
nor U40824 (N_40824,N_39840,N_39916);
and U40825 (N_40825,N_39741,N_39739);
nand U40826 (N_40826,N_39430,N_39058);
or U40827 (N_40827,N_39754,N_39867);
or U40828 (N_40828,N_39374,N_39190);
nand U40829 (N_40829,N_39134,N_39029);
nand U40830 (N_40830,N_39640,N_39215);
or U40831 (N_40831,N_39867,N_39446);
xor U40832 (N_40832,N_39016,N_39963);
and U40833 (N_40833,N_39403,N_39579);
xor U40834 (N_40834,N_39793,N_39016);
xnor U40835 (N_40835,N_39086,N_39796);
nor U40836 (N_40836,N_39645,N_39663);
xor U40837 (N_40837,N_39798,N_39371);
xnor U40838 (N_40838,N_39064,N_39402);
nand U40839 (N_40839,N_39556,N_39808);
xor U40840 (N_40840,N_39699,N_39485);
and U40841 (N_40841,N_39970,N_39630);
xor U40842 (N_40842,N_39663,N_39657);
xor U40843 (N_40843,N_39009,N_39511);
nor U40844 (N_40844,N_39132,N_39232);
nand U40845 (N_40845,N_39511,N_39113);
or U40846 (N_40846,N_39954,N_39120);
and U40847 (N_40847,N_39878,N_39217);
nor U40848 (N_40848,N_39049,N_39742);
nor U40849 (N_40849,N_39418,N_39948);
nand U40850 (N_40850,N_39392,N_39386);
and U40851 (N_40851,N_39859,N_39079);
xor U40852 (N_40852,N_39222,N_39273);
or U40853 (N_40853,N_39080,N_39994);
nand U40854 (N_40854,N_39514,N_39163);
or U40855 (N_40855,N_39778,N_39258);
or U40856 (N_40856,N_39061,N_39163);
nand U40857 (N_40857,N_39053,N_39385);
or U40858 (N_40858,N_39539,N_39707);
nand U40859 (N_40859,N_39701,N_39617);
nor U40860 (N_40860,N_39106,N_39128);
xor U40861 (N_40861,N_39867,N_39476);
nor U40862 (N_40862,N_39895,N_39220);
or U40863 (N_40863,N_39102,N_39911);
and U40864 (N_40864,N_39057,N_39327);
nor U40865 (N_40865,N_39188,N_39927);
nand U40866 (N_40866,N_39842,N_39967);
and U40867 (N_40867,N_39300,N_39152);
or U40868 (N_40868,N_39708,N_39031);
xor U40869 (N_40869,N_39508,N_39447);
nor U40870 (N_40870,N_39520,N_39426);
nor U40871 (N_40871,N_39597,N_39152);
nand U40872 (N_40872,N_39856,N_39064);
nand U40873 (N_40873,N_39553,N_39069);
xor U40874 (N_40874,N_39008,N_39380);
or U40875 (N_40875,N_39357,N_39278);
xnor U40876 (N_40876,N_39217,N_39503);
or U40877 (N_40877,N_39502,N_39315);
xor U40878 (N_40878,N_39467,N_39018);
xor U40879 (N_40879,N_39580,N_39606);
nand U40880 (N_40880,N_39752,N_39456);
and U40881 (N_40881,N_39036,N_39735);
nor U40882 (N_40882,N_39250,N_39064);
and U40883 (N_40883,N_39520,N_39306);
xor U40884 (N_40884,N_39472,N_39721);
or U40885 (N_40885,N_39599,N_39367);
and U40886 (N_40886,N_39729,N_39721);
and U40887 (N_40887,N_39650,N_39696);
xnor U40888 (N_40888,N_39348,N_39835);
nand U40889 (N_40889,N_39338,N_39431);
or U40890 (N_40890,N_39928,N_39603);
nor U40891 (N_40891,N_39019,N_39018);
nor U40892 (N_40892,N_39711,N_39502);
and U40893 (N_40893,N_39247,N_39298);
or U40894 (N_40894,N_39718,N_39513);
nand U40895 (N_40895,N_39999,N_39405);
and U40896 (N_40896,N_39963,N_39442);
xnor U40897 (N_40897,N_39640,N_39297);
and U40898 (N_40898,N_39757,N_39909);
nor U40899 (N_40899,N_39341,N_39320);
nand U40900 (N_40900,N_39952,N_39573);
or U40901 (N_40901,N_39941,N_39706);
and U40902 (N_40902,N_39898,N_39319);
or U40903 (N_40903,N_39279,N_39004);
or U40904 (N_40904,N_39948,N_39623);
and U40905 (N_40905,N_39842,N_39692);
xor U40906 (N_40906,N_39537,N_39130);
or U40907 (N_40907,N_39820,N_39686);
nand U40908 (N_40908,N_39565,N_39328);
nand U40909 (N_40909,N_39725,N_39631);
nand U40910 (N_40910,N_39647,N_39092);
nor U40911 (N_40911,N_39398,N_39154);
and U40912 (N_40912,N_39774,N_39440);
or U40913 (N_40913,N_39358,N_39807);
xnor U40914 (N_40914,N_39697,N_39749);
or U40915 (N_40915,N_39112,N_39273);
nand U40916 (N_40916,N_39815,N_39886);
or U40917 (N_40917,N_39015,N_39269);
or U40918 (N_40918,N_39588,N_39013);
xnor U40919 (N_40919,N_39672,N_39315);
and U40920 (N_40920,N_39476,N_39688);
and U40921 (N_40921,N_39362,N_39806);
nor U40922 (N_40922,N_39134,N_39303);
xor U40923 (N_40923,N_39126,N_39125);
nor U40924 (N_40924,N_39609,N_39301);
xor U40925 (N_40925,N_39380,N_39265);
nor U40926 (N_40926,N_39061,N_39089);
and U40927 (N_40927,N_39586,N_39650);
and U40928 (N_40928,N_39587,N_39472);
nand U40929 (N_40929,N_39733,N_39254);
or U40930 (N_40930,N_39922,N_39215);
nand U40931 (N_40931,N_39350,N_39404);
nand U40932 (N_40932,N_39125,N_39977);
nor U40933 (N_40933,N_39511,N_39335);
nand U40934 (N_40934,N_39499,N_39529);
nor U40935 (N_40935,N_39986,N_39207);
nor U40936 (N_40936,N_39774,N_39280);
xor U40937 (N_40937,N_39260,N_39525);
nand U40938 (N_40938,N_39545,N_39596);
or U40939 (N_40939,N_39616,N_39862);
xor U40940 (N_40940,N_39762,N_39007);
nand U40941 (N_40941,N_39499,N_39314);
xnor U40942 (N_40942,N_39995,N_39633);
and U40943 (N_40943,N_39354,N_39991);
nor U40944 (N_40944,N_39642,N_39498);
nand U40945 (N_40945,N_39541,N_39901);
nor U40946 (N_40946,N_39697,N_39766);
nand U40947 (N_40947,N_39952,N_39048);
or U40948 (N_40948,N_39766,N_39547);
nand U40949 (N_40949,N_39536,N_39656);
xor U40950 (N_40950,N_39690,N_39581);
or U40951 (N_40951,N_39337,N_39658);
nor U40952 (N_40952,N_39570,N_39802);
or U40953 (N_40953,N_39896,N_39420);
or U40954 (N_40954,N_39966,N_39114);
nor U40955 (N_40955,N_39979,N_39925);
xnor U40956 (N_40956,N_39274,N_39630);
xor U40957 (N_40957,N_39573,N_39401);
xor U40958 (N_40958,N_39555,N_39689);
xnor U40959 (N_40959,N_39526,N_39863);
xnor U40960 (N_40960,N_39266,N_39862);
or U40961 (N_40961,N_39031,N_39325);
xor U40962 (N_40962,N_39556,N_39567);
nand U40963 (N_40963,N_39258,N_39378);
nand U40964 (N_40964,N_39974,N_39461);
nand U40965 (N_40965,N_39979,N_39096);
xnor U40966 (N_40966,N_39953,N_39239);
nor U40967 (N_40967,N_39724,N_39690);
xor U40968 (N_40968,N_39091,N_39104);
xor U40969 (N_40969,N_39335,N_39126);
and U40970 (N_40970,N_39521,N_39692);
or U40971 (N_40971,N_39624,N_39982);
or U40972 (N_40972,N_39130,N_39526);
nor U40973 (N_40973,N_39058,N_39119);
nor U40974 (N_40974,N_39750,N_39558);
nor U40975 (N_40975,N_39609,N_39594);
nand U40976 (N_40976,N_39298,N_39165);
nor U40977 (N_40977,N_39386,N_39161);
or U40978 (N_40978,N_39882,N_39777);
nor U40979 (N_40979,N_39160,N_39991);
xnor U40980 (N_40980,N_39793,N_39454);
nor U40981 (N_40981,N_39140,N_39783);
and U40982 (N_40982,N_39994,N_39394);
nand U40983 (N_40983,N_39963,N_39914);
nor U40984 (N_40984,N_39898,N_39002);
or U40985 (N_40985,N_39784,N_39132);
nand U40986 (N_40986,N_39552,N_39312);
and U40987 (N_40987,N_39928,N_39634);
nor U40988 (N_40988,N_39357,N_39782);
nand U40989 (N_40989,N_39270,N_39191);
xnor U40990 (N_40990,N_39688,N_39708);
nor U40991 (N_40991,N_39297,N_39040);
and U40992 (N_40992,N_39299,N_39708);
nand U40993 (N_40993,N_39467,N_39438);
nor U40994 (N_40994,N_39289,N_39438);
nand U40995 (N_40995,N_39928,N_39218);
xor U40996 (N_40996,N_39185,N_39163);
and U40997 (N_40997,N_39564,N_39989);
nand U40998 (N_40998,N_39802,N_39818);
or U40999 (N_40999,N_39623,N_39134);
nand U41000 (N_41000,N_40163,N_40050);
and U41001 (N_41001,N_40158,N_40006);
and U41002 (N_41002,N_40090,N_40615);
nand U41003 (N_41003,N_40371,N_40619);
and U41004 (N_41004,N_40640,N_40466);
or U41005 (N_41005,N_40511,N_40890);
or U41006 (N_41006,N_40148,N_40297);
and U41007 (N_41007,N_40712,N_40273);
or U41008 (N_41008,N_40031,N_40233);
xor U41009 (N_41009,N_40390,N_40026);
and U41010 (N_41010,N_40957,N_40534);
and U41011 (N_41011,N_40405,N_40218);
xnor U41012 (N_41012,N_40682,N_40146);
or U41013 (N_41013,N_40473,N_40345);
nand U41014 (N_41014,N_40452,N_40175);
xnor U41015 (N_41015,N_40036,N_40754);
nor U41016 (N_41016,N_40923,N_40016);
nor U41017 (N_41017,N_40500,N_40424);
xor U41018 (N_41018,N_40654,N_40028);
xor U41019 (N_41019,N_40630,N_40467);
nand U41020 (N_41020,N_40949,N_40816);
xnor U41021 (N_41021,N_40353,N_40337);
and U41022 (N_41022,N_40734,N_40828);
nor U41023 (N_41023,N_40454,N_40625);
and U41024 (N_41024,N_40128,N_40972);
xor U41025 (N_41025,N_40495,N_40237);
or U41026 (N_41026,N_40608,N_40915);
and U41027 (N_41027,N_40303,N_40746);
or U41028 (N_41028,N_40066,N_40341);
or U41029 (N_41029,N_40242,N_40636);
and U41030 (N_41030,N_40496,N_40269);
nand U41031 (N_41031,N_40966,N_40888);
or U41032 (N_41032,N_40839,N_40598);
nand U41033 (N_41033,N_40022,N_40731);
xnor U41034 (N_41034,N_40008,N_40385);
nand U41035 (N_41035,N_40679,N_40898);
nor U41036 (N_41036,N_40662,N_40902);
xnor U41037 (N_41037,N_40781,N_40127);
or U41038 (N_41038,N_40185,N_40650);
xor U41039 (N_41039,N_40751,N_40876);
nor U41040 (N_41040,N_40172,N_40208);
and U41041 (N_41041,N_40577,N_40115);
nand U41042 (N_41042,N_40877,N_40362);
and U41043 (N_41043,N_40271,N_40551);
nand U41044 (N_41044,N_40328,N_40043);
nand U41045 (N_41045,N_40291,N_40100);
xnor U41046 (N_41046,N_40289,N_40699);
xnor U41047 (N_41047,N_40634,N_40716);
xnor U41048 (N_41048,N_40072,N_40344);
or U41049 (N_41049,N_40926,N_40453);
xnor U41050 (N_41050,N_40258,N_40837);
nor U41051 (N_41051,N_40609,N_40510);
nand U41052 (N_41052,N_40098,N_40985);
xor U41053 (N_41053,N_40824,N_40826);
nand U41054 (N_41054,N_40478,N_40783);
and U41055 (N_41055,N_40672,N_40162);
or U41056 (N_41056,N_40874,N_40263);
nand U41057 (N_41057,N_40856,N_40411);
nand U41058 (N_41058,N_40231,N_40339);
xnor U41059 (N_41059,N_40327,N_40363);
nand U41060 (N_41060,N_40181,N_40548);
and U41061 (N_41061,N_40477,N_40338);
and U41062 (N_41062,N_40504,N_40205);
or U41063 (N_41063,N_40546,N_40110);
or U41064 (N_41064,N_40101,N_40914);
or U41065 (N_41065,N_40618,N_40795);
xnor U41066 (N_41066,N_40270,N_40850);
or U41067 (N_41067,N_40536,N_40594);
xor U41068 (N_41068,N_40944,N_40592);
xnor U41069 (N_41069,N_40492,N_40516);
and U41070 (N_41070,N_40917,N_40011);
nor U41071 (N_41071,N_40097,N_40855);
nor U41072 (N_41072,N_40626,N_40800);
xor U41073 (N_41073,N_40203,N_40003);
xor U41074 (N_41074,N_40463,N_40590);
and U41075 (N_41075,N_40843,N_40212);
xnor U41076 (N_41076,N_40535,N_40108);
and U41077 (N_41077,N_40605,N_40964);
or U41078 (N_41078,N_40714,N_40760);
xor U41079 (N_41079,N_40403,N_40829);
xnor U41080 (N_41080,N_40227,N_40204);
and U41081 (N_41081,N_40245,N_40486);
nand U41082 (N_41082,N_40095,N_40659);
nand U41083 (N_41083,N_40152,N_40791);
and U41084 (N_41084,N_40789,N_40429);
or U41085 (N_41085,N_40684,N_40051);
xor U41086 (N_41086,N_40870,N_40431);
nand U41087 (N_41087,N_40210,N_40787);
nor U41088 (N_41088,N_40134,N_40053);
nor U41089 (N_41089,N_40666,N_40275);
and U41090 (N_41090,N_40260,N_40136);
nor U41091 (N_41091,N_40417,N_40696);
nand U41092 (N_41092,N_40343,N_40897);
or U41093 (N_41093,N_40846,N_40907);
nand U41094 (N_41094,N_40241,N_40281);
xor U41095 (N_41095,N_40628,N_40740);
xor U41096 (N_41096,N_40202,N_40295);
nor U41097 (N_41097,N_40419,N_40412);
xnor U41098 (N_41098,N_40566,N_40503);
or U41099 (N_41099,N_40316,N_40280);
xor U41100 (N_41100,N_40934,N_40300);
or U41101 (N_41101,N_40811,N_40767);
nand U41102 (N_41102,N_40235,N_40445);
nor U41103 (N_41103,N_40788,N_40180);
nor U41104 (N_41104,N_40447,N_40644);
or U41105 (N_41105,N_40895,N_40196);
xnor U41106 (N_41106,N_40860,N_40435);
and U41107 (N_41107,N_40436,N_40893);
or U41108 (N_41108,N_40921,N_40188);
and U41109 (N_41109,N_40759,N_40437);
nor U41110 (N_41110,N_40611,N_40414);
nand U41111 (N_41111,N_40284,N_40765);
nand U41112 (N_41112,N_40603,N_40499);
nand U41113 (N_41113,N_40836,N_40970);
nor U41114 (N_41114,N_40963,N_40604);
and U41115 (N_41115,N_40382,N_40621);
or U41116 (N_41116,N_40332,N_40698);
or U41117 (N_41117,N_40918,N_40519);
nand U41118 (N_41118,N_40794,N_40637);
xnor U41119 (N_41119,N_40461,N_40556);
nor U41120 (N_41120,N_40081,N_40039);
and U41121 (N_41121,N_40960,N_40333);
xor U41122 (N_41122,N_40380,N_40935);
or U41123 (N_41123,N_40049,N_40817);
nand U41124 (N_41124,N_40552,N_40543);
or U41125 (N_41125,N_40430,N_40501);
nand U41126 (N_41126,N_40804,N_40361);
or U41127 (N_41127,N_40931,N_40991);
nor U41128 (N_41128,N_40340,N_40497);
xor U41129 (N_41129,N_40773,N_40292);
xnor U41130 (N_41130,N_40267,N_40132);
nor U41131 (N_41131,N_40656,N_40302);
nor U41132 (N_41132,N_40780,N_40190);
or U41133 (N_41133,N_40711,N_40366);
nor U41134 (N_41134,N_40223,N_40715);
nand U41135 (N_41135,N_40434,N_40232);
nor U41136 (N_41136,N_40958,N_40886);
and U41137 (N_41137,N_40784,N_40540);
nor U41138 (N_41138,N_40324,N_40018);
nand U41139 (N_41139,N_40512,N_40624);
nor U41140 (N_41140,N_40950,N_40480);
and U41141 (N_41141,N_40491,N_40655);
or U41142 (N_41142,N_40732,N_40936);
nand U41143 (N_41143,N_40872,N_40847);
xnor U41144 (N_41144,N_40867,N_40080);
or U41145 (N_41145,N_40642,N_40538);
nand U41146 (N_41146,N_40348,N_40755);
and U41147 (N_41147,N_40122,N_40635);
or U41148 (N_41148,N_40472,N_40677);
nor U41149 (N_41149,N_40730,N_40272);
and U41150 (N_41150,N_40588,N_40962);
nor U41151 (N_41151,N_40290,N_40364);
xor U41152 (N_41152,N_40879,N_40299);
xor U41153 (N_41153,N_40941,N_40074);
or U41154 (N_41154,N_40091,N_40213);
and U41155 (N_41155,N_40087,N_40216);
nand U41156 (N_41156,N_40806,N_40660);
xnor U41157 (N_41157,N_40368,N_40733);
and U41158 (N_41158,N_40600,N_40595);
or U41159 (N_41159,N_40415,N_40779);
or U41160 (N_41160,N_40667,N_40307);
or U41161 (N_41161,N_40129,N_40997);
nand U41162 (N_41162,N_40927,N_40040);
and U41163 (N_41163,N_40296,N_40995);
or U41164 (N_41164,N_40124,N_40912);
and U41165 (N_41165,N_40570,N_40597);
and U41166 (N_41166,N_40517,N_40862);
xnor U41167 (N_41167,N_40739,N_40748);
or U41168 (N_41168,N_40520,N_40481);
or U41169 (N_41169,N_40657,N_40671);
xnor U41170 (N_41170,N_40236,N_40614);
or U41171 (N_41171,N_40632,N_40077);
nor U41172 (N_41172,N_40541,N_40703);
nor U41173 (N_41173,N_40537,N_40121);
and U41174 (N_41174,N_40582,N_40880);
nand U41175 (N_41175,N_40211,N_40617);
nor U41176 (N_41176,N_40406,N_40959);
and U41177 (N_41177,N_40903,N_40402);
or U41178 (N_41178,N_40891,N_40919);
nand U41179 (N_41179,N_40736,N_40769);
or U41180 (N_41180,N_40842,N_40017);
nand U41181 (N_41181,N_40401,N_40622);
or U41182 (N_41182,N_40126,N_40356);
nor U41183 (N_41183,N_40854,N_40484);
nor U41184 (N_41184,N_40286,N_40961);
or U41185 (N_41185,N_40764,N_40442);
nor U41186 (N_41186,N_40745,N_40111);
nor U41187 (N_41187,N_40749,N_40974);
nor U41188 (N_41188,N_40351,N_40372);
xnor U41189 (N_41189,N_40825,N_40680);
nand U41190 (N_41190,N_40103,N_40056);
nor U41191 (N_41191,N_40996,N_40981);
xnor U41192 (N_41192,N_40407,N_40584);
and U41193 (N_41193,N_40174,N_40563);
xor U41194 (N_41194,N_40393,N_40485);
or U41195 (N_41195,N_40166,N_40729);
and U41196 (N_41196,N_40845,N_40593);
and U41197 (N_41197,N_40409,N_40325);
or U41198 (N_41198,N_40658,N_40557);
or U41199 (N_41199,N_40612,N_40892);
xor U41200 (N_41200,N_40192,N_40905);
and U41201 (N_41201,N_40085,N_40518);
xnor U41202 (N_41202,N_40306,N_40065);
or U41203 (N_41203,N_40809,N_40195);
and U41204 (N_41204,N_40243,N_40578);
nor U41205 (N_41205,N_40901,N_40579);
and U41206 (N_41206,N_40631,N_40048);
nor U41207 (N_41207,N_40648,N_40864);
and U41208 (N_41208,N_40314,N_40396);
or U41209 (N_41209,N_40147,N_40335);
nand U41210 (N_41210,N_40906,N_40138);
nor U41211 (N_41211,N_40727,N_40940);
and U41212 (N_41212,N_40482,N_40651);
or U41213 (N_41213,N_40186,N_40439);
and U41214 (N_41214,N_40803,N_40287);
nand U41215 (N_41215,N_40792,N_40383);
xnor U41216 (N_41216,N_40665,N_40153);
nand U41217 (N_41217,N_40037,N_40367);
nor U41218 (N_41218,N_40591,N_40820);
nand U41219 (N_41219,N_40268,N_40875);
or U41220 (N_41220,N_40214,N_40399);
and U41221 (N_41221,N_40565,N_40616);
and U41222 (N_41222,N_40882,N_40713);
nand U41223 (N_41223,N_40264,N_40946);
and U41224 (N_41224,N_40564,N_40451);
xnor U41225 (N_41225,N_40157,N_40347);
xnor U41226 (N_41226,N_40060,N_40248);
nor U41227 (N_41227,N_40032,N_40955);
nand U41228 (N_41228,N_40887,N_40379);
and U41229 (N_41229,N_40276,N_40818);
nand U41230 (N_41230,N_40813,N_40130);
nand U41231 (N_41231,N_40596,N_40560);
nor U41232 (N_41232,N_40189,N_40498);
or U41233 (N_41233,N_40278,N_40774);
nand U41234 (N_41234,N_40908,N_40865);
nand U41235 (N_41235,N_40558,N_40425);
nand U41236 (N_41236,N_40222,N_40687);
xnor U41237 (N_41237,N_40848,N_40391);
and U41238 (N_41238,N_40861,N_40513);
xor U41239 (N_41239,N_40525,N_40683);
or U41240 (N_41240,N_40573,N_40691);
nand U41241 (N_41241,N_40164,N_40542);
nand U41242 (N_41242,N_40092,N_40199);
xor U41243 (N_41243,N_40441,N_40140);
xnor U41244 (N_41244,N_40559,N_40045);
nand U41245 (N_41245,N_40827,N_40360);
nand U41246 (N_41246,N_40911,N_40515);
xor U41247 (N_41247,N_40693,N_40724);
nand U41248 (N_41248,N_40853,N_40194);
nand U41249 (N_41249,N_40768,N_40446);
nand U41250 (N_41250,N_40697,N_40661);
nand U41251 (N_41251,N_40885,N_40234);
or U41252 (N_41252,N_40953,N_40823);
nor U41253 (N_41253,N_40775,N_40802);
or U41254 (N_41254,N_40154,N_40322);
nor U41255 (N_41255,N_40722,N_40301);
xor U41256 (N_41256,N_40277,N_40752);
nor U41257 (N_41257,N_40844,N_40082);
xnor U41258 (N_41258,N_40704,N_40990);
xnor U41259 (N_41259,N_40059,N_40020);
nand U41260 (N_41260,N_40514,N_40038);
and U41261 (N_41261,N_40144,N_40455);
and U41262 (N_41262,N_40776,N_40025);
or U41263 (N_41263,N_40553,N_40220);
or U41264 (N_41264,N_40014,N_40173);
or U41265 (N_41265,N_40217,N_40197);
and U41266 (N_41266,N_40329,N_40444);
nor U41267 (N_41267,N_40607,N_40118);
xor U41268 (N_41268,N_40397,N_40968);
nand U41269 (N_41269,N_40283,N_40475);
nor U41270 (N_41270,N_40571,N_40143);
xor U41271 (N_41271,N_40574,N_40330);
xnor U41272 (N_41272,N_40250,N_40613);
nor U41273 (N_41273,N_40975,N_40871);
nand U41274 (N_41274,N_40743,N_40798);
xor U41275 (N_41275,N_40377,N_40058);
xor U41276 (N_41276,N_40531,N_40835);
nor U41277 (N_41277,N_40814,N_40606);
nor U41278 (N_41278,N_40244,N_40061);
xor U41279 (N_41279,N_40352,N_40884);
or U41280 (N_41280,N_40052,N_40471);
nand U41281 (N_41281,N_40954,N_40866);
xnor U41282 (N_41282,N_40527,N_40029);
nor U41283 (N_41283,N_40669,N_40119);
xor U41284 (N_41284,N_40978,N_40801);
or U41285 (N_41285,N_40054,N_40331);
or U41286 (N_41286,N_40965,N_40159);
or U41287 (N_41287,N_40249,N_40423);
nand U41288 (N_41288,N_40742,N_40252);
nor U41289 (N_41289,N_40002,N_40796);
or U41290 (N_41290,N_40388,N_40750);
nor U41291 (N_41291,N_40812,N_40987);
and U41292 (N_41292,N_40178,N_40378);
xnor U41293 (N_41293,N_40834,N_40833);
or U41294 (N_41294,N_40246,N_40469);
nand U41295 (N_41295,N_40488,N_40427);
and U41296 (N_41296,N_40585,N_40323);
or U41297 (N_41297,N_40668,N_40561);
and U41298 (N_41298,N_40418,N_40994);
xor U41299 (N_41299,N_40070,N_40521);
nor U41300 (N_41300,N_40084,N_40530);
or U41301 (N_41301,N_40942,N_40432);
nor U41302 (N_41302,N_40676,N_40062);
nor U41303 (N_41303,N_40096,N_40116);
nor U41304 (N_41304,N_40398,N_40042);
nand U41305 (N_41305,N_40309,N_40448);
and U41306 (N_41306,N_40171,N_40647);
xnor U41307 (N_41307,N_40601,N_40822);
nor U41308 (N_41308,N_40685,N_40544);
and U41309 (N_41309,N_40920,N_40695);
xnor U41310 (N_41310,N_40782,N_40753);
xnor U41311 (N_41311,N_40114,N_40030);
nor U41312 (N_41312,N_40718,N_40365);
or U41313 (N_41313,N_40013,N_40240);
and U41314 (N_41314,N_40373,N_40312);
xor U41315 (N_41315,N_40744,N_40404);
or U41316 (N_41316,N_40161,N_40868);
nand U41317 (N_41317,N_40009,N_40462);
xor U41318 (N_41318,N_40689,N_40044);
nor U41319 (N_41319,N_40456,N_40633);
nand U41320 (N_41320,N_40145,N_40762);
nor U41321 (N_41321,N_40627,N_40089);
xnor U41322 (N_41322,N_40487,N_40641);
or U41323 (N_41323,N_40569,N_40664);
nand U41324 (N_41324,N_40120,N_40165);
or U41325 (N_41325,N_40359,N_40015);
nand U41326 (N_41326,N_40863,N_40977);
nor U41327 (N_41327,N_40988,N_40652);
and U41328 (N_41328,N_40984,N_40725);
nor U41329 (N_41329,N_40394,N_40086);
xor U41330 (N_41330,N_40169,N_40924);
or U41331 (N_41331,N_40758,N_40841);
nand U41332 (N_41332,N_40998,N_40160);
nor U41333 (N_41333,N_40187,N_40012);
and U41334 (N_41334,N_40288,N_40476);
and U41335 (N_41335,N_40034,N_40420);
and U41336 (N_41336,N_40993,N_40150);
nand U41337 (N_41337,N_40468,N_40529);
nor U41338 (N_41338,N_40639,N_40980);
or U41339 (N_41339,N_40149,N_40849);
nand U41340 (N_41340,N_40545,N_40215);
or U41341 (N_41341,N_40810,N_40999);
nor U41342 (N_41342,N_40728,N_40093);
and U41343 (N_41343,N_40900,N_40878);
nand U41344 (N_41344,N_40255,N_40112);
nand U41345 (N_41345,N_40310,N_40673);
nand U41346 (N_41346,N_40719,N_40191);
or U41347 (N_41347,N_40983,N_40073);
and U41348 (N_41348,N_40139,N_40969);
xnor U41349 (N_41349,N_40308,N_40317);
nand U41350 (N_41350,N_40083,N_40643);
nand U41351 (N_41351,N_40021,N_40102);
nand U41352 (N_41352,N_40392,N_40428);
and U41353 (N_41353,N_40135,N_40979);
and U41354 (N_41354,N_40071,N_40830);
xnor U41355 (N_41355,N_40799,N_40620);
xnor U41356 (N_41356,N_40460,N_40088);
nor U41357 (N_41357,N_40443,N_40155);
nand U41358 (N_41358,N_40311,N_40209);
or U41359 (N_41359,N_40479,N_40357);
nand U41360 (N_41360,N_40505,N_40326);
nand U41361 (N_41361,N_40881,N_40770);
nor U41362 (N_41362,N_40395,N_40726);
nor U41363 (N_41363,N_40170,N_40305);
and U41364 (N_41364,N_40939,N_40528);
and U41365 (N_41365,N_40747,N_40449);
nand U41366 (N_41366,N_40678,N_40575);
or U41367 (N_41367,N_40355,N_40674);
and U41368 (N_41368,N_40623,N_40832);
nand U41369 (N_41369,N_40945,N_40221);
nand U41370 (N_41370,N_40230,N_40933);
nor U41371 (N_41371,N_40167,N_40123);
xor U41372 (N_41372,N_40932,N_40433);
xor U41373 (N_41373,N_40757,N_40777);
nor U41374 (N_41374,N_40523,N_40063);
nor U41375 (N_41375,N_40131,N_40156);
or U41376 (N_41376,N_40638,N_40938);
nor U41377 (N_41377,N_40587,N_40710);
nor U41378 (N_41378,N_40438,N_40226);
or U41379 (N_41379,N_40646,N_40986);
nand U41380 (N_41380,N_40251,N_40416);
xor U41381 (N_41381,N_40207,N_40922);
xor U41382 (N_41382,N_40069,N_40735);
nor U41383 (N_41383,N_40738,N_40952);
xor U41384 (N_41384,N_40904,N_40182);
xor U41385 (N_41385,N_40723,N_40334);
nor U41386 (N_41386,N_40894,N_40539);
or U41387 (N_41387,N_40489,N_40198);
nand U41388 (N_41388,N_40000,N_40873);
nor U41389 (N_41389,N_40599,N_40228);
nor U41390 (N_41390,N_40304,N_40247);
and U41391 (N_41391,N_40067,N_40298);
or U41392 (N_41392,N_40522,N_40346);
nor U41393 (N_41393,N_40708,N_40778);
nor U41394 (N_41394,N_40982,N_40282);
or U41395 (N_41395,N_40464,N_40374);
and U41396 (N_41396,N_40688,N_40099);
or U41397 (N_41397,N_40909,N_40450);
nand U41398 (N_41398,N_40265,N_40858);
and U41399 (N_41399,N_40702,N_40075);
or U41400 (N_41400,N_40336,N_40184);
nand U41401 (N_41401,N_40177,N_40686);
and U41402 (N_41402,N_40293,N_40046);
and U41403 (N_41403,N_40319,N_40701);
xor U41404 (N_41404,N_40494,N_40113);
xnor U41405 (N_41405,N_40350,N_40315);
xnor U41406 (N_41406,N_40389,N_40602);
and U41407 (N_41407,N_40193,N_40257);
or U41408 (N_41408,N_40930,N_40001);
or U41409 (N_41409,N_40440,N_40502);
or U41410 (N_41410,N_40109,N_40707);
or U41411 (N_41411,N_40376,N_40400);
and U41412 (N_41412,N_40079,N_40550);
xor U41413 (N_41413,N_40179,N_40151);
and U41414 (N_41414,N_40869,N_40554);
and U41415 (N_41415,N_40470,N_40384);
or U41416 (N_41416,N_40547,N_40386);
or U41417 (N_41417,N_40493,N_40567);
xor U41418 (N_41418,N_40206,N_40422);
and U41419 (N_41419,N_40706,N_40024);
nor U41420 (N_41420,N_40313,N_40610);
nor U41421 (N_41421,N_40943,N_40035);
and U41422 (N_41422,N_40976,N_40705);
nor U41423 (N_41423,N_40709,N_40508);
nor U41424 (N_41424,N_40629,N_40786);
nor U41425 (N_41425,N_40851,N_40266);
and U41426 (N_41426,N_40106,N_40005);
and U41427 (N_41427,N_40805,N_40572);
nand U41428 (N_41428,N_40737,N_40410);
or U41429 (N_41429,N_40007,N_40262);
and U41430 (N_41430,N_40224,N_40318);
xor U41431 (N_41431,N_40229,N_40490);
nor U41432 (N_41432,N_40465,N_40663);
and U41433 (N_41433,N_40375,N_40064);
xor U41434 (N_41434,N_40474,N_40105);
nand U41435 (N_41435,N_40951,N_40690);
and U41436 (N_41436,N_40645,N_40259);
nor U41437 (N_41437,N_40532,N_40720);
and U41438 (N_41438,N_40509,N_40681);
or U41439 (N_41439,N_40771,N_40838);
nor U41440 (N_41440,N_40370,N_40653);
xor U41441 (N_41441,N_40507,N_40785);
nor U41442 (N_41442,N_40041,N_40239);
nand U41443 (N_41443,N_40033,N_40426);
nor U41444 (N_41444,N_40692,N_40852);
xor U41445 (N_41445,N_40225,N_40483);
and U41446 (N_41446,N_40819,N_40256);
and U41447 (N_41447,N_40568,N_40992);
nand U41448 (N_41448,N_40675,N_40142);
and U41449 (N_41449,N_40948,N_40807);
nand U41450 (N_41450,N_40967,N_40790);
xnor U41451 (N_41451,N_40670,N_40506);
and U41452 (N_41452,N_40358,N_40916);
xnor U41453 (N_41453,N_40793,N_40586);
nand U41454 (N_41454,N_40253,N_40925);
and U41455 (N_41455,N_40078,N_40133);
nand U41456 (N_41456,N_40956,N_40889);
nor U41457 (N_41457,N_40381,N_40254);
nor U41458 (N_41458,N_40883,N_40576);
and U41459 (N_41459,N_40354,N_40555);
and U41460 (N_41460,N_40219,N_40928);
nor U41461 (N_41461,N_40458,N_40721);
nand U41462 (N_41462,N_40141,N_40027);
nor U41463 (N_41463,N_40937,N_40700);
xor U41464 (N_41464,N_40408,N_40859);
xnor U41465 (N_41465,N_40176,N_40107);
nand U41466 (N_41466,N_40349,N_40581);
xor U41467 (N_41467,N_40524,N_40387);
or U41468 (N_41468,N_40010,N_40741);
xnor U41469 (N_41469,N_40183,N_40549);
and U41470 (N_41470,N_40533,N_40320);
nor U41471 (N_41471,N_40694,N_40899);
xnor U41472 (N_41472,N_40913,N_40989);
or U41473 (N_41473,N_40459,N_40929);
xor U41474 (N_41474,N_40808,N_40910);
or U41475 (N_41475,N_40831,N_40369);
nor U41476 (N_41476,N_40756,N_40717);
or U41477 (N_41477,N_40285,N_40294);
and U41478 (N_41478,N_40649,N_40526);
xnor U41479 (N_41479,N_40201,N_40973);
nor U41480 (N_41480,N_40583,N_40023);
nand U41481 (N_41481,N_40200,N_40274);
xor U41482 (N_41482,N_40797,N_40094);
and U41483 (N_41483,N_40168,N_40947);
nand U41484 (N_41484,N_40772,N_40971);
or U41485 (N_41485,N_40457,N_40004);
nor U41486 (N_41486,N_40580,N_40076);
or U41487 (N_41487,N_40057,N_40279);
nor U41488 (N_41488,N_40068,N_40821);
xnor U41489 (N_41489,N_40238,N_40562);
nor U41490 (N_41490,N_40766,N_40137);
nand U41491 (N_41491,N_40761,N_40413);
nor U41492 (N_41492,N_40321,N_40421);
and U41493 (N_41493,N_40047,N_40896);
xnor U41494 (N_41494,N_40763,N_40019);
xor U41495 (N_41495,N_40342,N_40055);
and U41496 (N_41496,N_40104,N_40840);
xnor U41497 (N_41497,N_40815,N_40857);
xnor U41498 (N_41498,N_40261,N_40125);
nand U41499 (N_41499,N_40589,N_40117);
nand U41500 (N_41500,N_40785,N_40818);
or U41501 (N_41501,N_40753,N_40250);
nor U41502 (N_41502,N_40693,N_40432);
nand U41503 (N_41503,N_40070,N_40652);
nor U41504 (N_41504,N_40997,N_40226);
nor U41505 (N_41505,N_40480,N_40897);
or U41506 (N_41506,N_40107,N_40926);
xor U41507 (N_41507,N_40036,N_40654);
nand U41508 (N_41508,N_40510,N_40489);
nor U41509 (N_41509,N_40658,N_40799);
or U41510 (N_41510,N_40748,N_40033);
and U41511 (N_41511,N_40877,N_40652);
xor U41512 (N_41512,N_40574,N_40703);
or U41513 (N_41513,N_40249,N_40393);
nor U41514 (N_41514,N_40576,N_40323);
nor U41515 (N_41515,N_40923,N_40293);
xnor U41516 (N_41516,N_40394,N_40410);
and U41517 (N_41517,N_40942,N_40067);
xnor U41518 (N_41518,N_40653,N_40598);
nand U41519 (N_41519,N_40231,N_40670);
nand U41520 (N_41520,N_40042,N_40239);
xor U41521 (N_41521,N_40101,N_40676);
nand U41522 (N_41522,N_40592,N_40488);
nor U41523 (N_41523,N_40282,N_40954);
or U41524 (N_41524,N_40739,N_40230);
xor U41525 (N_41525,N_40867,N_40454);
or U41526 (N_41526,N_40827,N_40434);
and U41527 (N_41527,N_40816,N_40170);
and U41528 (N_41528,N_40409,N_40886);
nor U41529 (N_41529,N_40489,N_40545);
xor U41530 (N_41530,N_40571,N_40147);
xnor U41531 (N_41531,N_40984,N_40844);
and U41532 (N_41532,N_40252,N_40816);
nor U41533 (N_41533,N_40001,N_40830);
and U41534 (N_41534,N_40305,N_40050);
and U41535 (N_41535,N_40093,N_40740);
or U41536 (N_41536,N_40307,N_40841);
or U41537 (N_41537,N_40728,N_40793);
and U41538 (N_41538,N_40625,N_40561);
and U41539 (N_41539,N_40930,N_40505);
and U41540 (N_41540,N_40246,N_40102);
or U41541 (N_41541,N_40538,N_40948);
nand U41542 (N_41542,N_40861,N_40210);
nand U41543 (N_41543,N_40686,N_40294);
and U41544 (N_41544,N_40499,N_40011);
xnor U41545 (N_41545,N_40136,N_40548);
and U41546 (N_41546,N_40784,N_40170);
xnor U41547 (N_41547,N_40669,N_40118);
nor U41548 (N_41548,N_40905,N_40839);
or U41549 (N_41549,N_40671,N_40385);
nor U41550 (N_41550,N_40913,N_40157);
and U41551 (N_41551,N_40131,N_40151);
nand U41552 (N_41552,N_40102,N_40539);
and U41553 (N_41553,N_40719,N_40976);
nor U41554 (N_41554,N_40966,N_40868);
nor U41555 (N_41555,N_40142,N_40266);
or U41556 (N_41556,N_40407,N_40152);
nand U41557 (N_41557,N_40656,N_40843);
xor U41558 (N_41558,N_40077,N_40523);
or U41559 (N_41559,N_40314,N_40269);
nor U41560 (N_41560,N_40878,N_40031);
nor U41561 (N_41561,N_40513,N_40434);
and U41562 (N_41562,N_40260,N_40629);
nor U41563 (N_41563,N_40515,N_40514);
and U41564 (N_41564,N_40860,N_40183);
nand U41565 (N_41565,N_40246,N_40599);
nand U41566 (N_41566,N_40412,N_40981);
or U41567 (N_41567,N_40649,N_40916);
nor U41568 (N_41568,N_40635,N_40593);
or U41569 (N_41569,N_40113,N_40074);
nor U41570 (N_41570,N_40182,N_40154);
nand U41571 (N_41571,N_40292,N_40965);
nand U41572 (N_41572,N_40084,N_40428);
or U41573 (N_41573,N_40013,N_40001);
xor U41574 (N_41574,N_40101,N_40679);
nor U41575 (N_41575,N_40487,N_40698);
nand U41576 (N_41576,N_40201,N_40938);
or U41577 (N_41577,N_40849,N_40421);
nand U41578 (N_41578,N_40996,N_40651);
nor U41579 (N_41579,N_40114,N_40767);
nor U41580 (N_41580,N_40716,N_40455);
nor U41581 (N_41581,N_40627,N_40149);
nor U41582 (N_41582,N_40423,N_40729);
or U41583 (N_41583,N_40682,N_40058);
nor U41584 (N_41584,N_40681,N_40874);
xnor U41585 (N_41585,N_40921,N_40537);
and U41586 (N_41586,N_40646,N_40977);
nor U41587 (N_41587,N_40565,N_40262);
nor U41588 (N_41588,N_40176,N_40747);
nand U41589 (N_41589,N_40526,N_40469);
xnor U41590 (N_41590,N_40059,N_40270);
or U41591 (N_41591,N_40116,N_40583);
and U41592 (N_41592,N_40791,N_40749);
nand U41593 (N_41593,N_40909,N_40393);
xor U41594 (N_41594,N_40474,N_40170);
and U41595 (N_41595,N_40923,N_40719);
nand U41596 (N_41596,N_40828,N_40705);
nor U41597 (N_41597,N_40997,N_40281);
nand U41598 (N_41598,N_40537,N_40755);
and U41599 (N_41599,N_40821,N_40990);
or U41600 (N_41600,N_40799,N_40269);
and U41601 (N_41601,N_40340,N_40279);
or U41602 (N_41602,N_40018,N_40180);
nand U41603 (N_41603,N_40972,N_40896);
and U41604 (N_41604,N_40133,N_40848);
nor U41605 (N_41605,N_40260,N_40137);
nor U41606 (N_41606,N_40332,N_40236);
nor U41607 (N_41607,N_40665,N_40476);
xnor U41608 (N_41608,N_40646,N_40481);
nor U41609 (N_41609,N_40867,N_40982);
nor U41610 (N_41610,N_40785,N_40251);
nand U41611 (N_41611,N_40539,N_40719);
nor U41612 (N_41612,N_40021,N_40535);
nor U41613 (N_41613,N_40839,N_40921);
and U41614 (N_41614,N_40830,N_40895);
and U41615 (N_41615,N_40788,N_40885);
nor U41616 (N_41616,N_40916,N_40758);
and U41617 (N_41617,N_40763,N_40339);
nand U41618 (N_41618,N_40668,N_40160);
nand U41619 (N_41619,N_40977,N_40422);
nand U41620 (N_41620,N_40985,N_40934);
and U41621 (N_41621,N_40441,N_40005);
nand U41622 (N_41622,N_40780,N_40356);
or U41623 (N_41623,N_40441,N_40526);
and U41624 (N_41624,N_40282,N_40868);
nor U41625 (N_41625,N_40885,N_40905);
and U41626 (N_41626,N_40241,N_40509);
and U41627 (N_41627,N_40551,N_40833);
xor U41628 (N_41628,N_40487,N_40006);
and U41629 (N_41629,N_40146,N_40532);
xor U41630 (N_41630,N_40662,N_40377);
nor U41631 (N_41631,N_40274,N_40566);
nor U41632 (N_41632,N_40290,N_40637);
or U41633 (N_41633,N_40186,N_40209);
xor U41634 (N_41634,N_40690,N_40387);
xnor U41635 (N_41635,N_40384,N_40273);
or U41636 (N_41636,N_40826,N_40335);
nor U41637 (N_41637,N_40989,N_40839);
and U41638 (N_41638,N_40607,N_40264);
xnor U41639 (N_41639,N_40850,N_40186);
and U41640 (N_41640,N_40916,N_40501);
or U41641 (N_41641,N_40241,N_40808);
nor U41642 (N_41642,N_40607,N_40460);
nor U41643 (N_41643,N_40557,N_40706);
and U41644 (N_41644,N_40002,N_40397);
nor U41645 (N_41645,N_40562,N_40687);
or U41646 (N_41646,N_40536,N_40709);
and U41647 (N_41647,N_40628,N_40370);
nand U41648 (N_41648,N_40661,N_40763);
xnor U41649 (N_41649,N_40203,N_40804);
nor U41650 (N_41650,N_40395,N_40634);
nand U41651 (N_41651,N_40402,N_40545);
and U41652 (N_41652,N_40669,N_40300);
nor U41653 (N_41653,N_40242,N_40795);
and U41654 (N_41654,N_40891,N_40993);
nand U41655 (N_41655,N_40097,N_40167);
or U41656 (N_41656,N_40103,N_40978);
and U41657 (N_41657,N_40310,N_40239);
xor U41658 (N_41658,N_40041,N_40584);
or U41659 (N_41659,N_40276,N_40573);
and U41660 (N_41660,N_40840,N_40833);
and U41661 (N_41661,N_40026,N_40418);
or U41662 (N_41662,N_40139,N_40706);
and U41663 (N_41663,N_40479,N_40416);
nor U41664 (N_41664,N_40167,N_40076);
and U41665 (N_41665,N_40181,N_40760);
xnor U41666 (N_41666,N_40134,N_40717);
and U41667 (N_41667,N_40808,N_40172);
xor U41668 (N_41668,N_40136,N_40941);
nor U41669 (N_41669,N_40952,N_40168);
nor U41670 (N_41670,N_40170,N_40835);
xor U41671 (N_41671,N_40371,N_40444);
and U41672 (N_41672,N_40919,N_40815);
nand U41673 (N_41673,N_40075,N_40041);
or U41674 (N_41674,N_40707,N_40371);
xnor U41675 (N_41675,N_40762,N_40105);
xor U41676 (N_41676,N_40876,N_40938);
nor U41677 (N_41677,N_40610,N_40420);
and U41678 (N_41678,N_40830,N_40655);
xnor U41679 (N_41679,N_40086,N_40267);
nand U41680 (N_41680,N_40427,N_40200);
nor U41681 (N_41681,N_40809,N_40978);
nor U41682 (N_41682,N_40101,N_40607);
and U41683 (N_41683,N_40336,N_40307);
nor U41684 (N_41684,N_40213,N_40699);
and U41685 (N_41685,N_40468,N_40998);
and U41686 (N_41686,N_40735,N_40943);
xor U41687 (N_41687,N_40836,N_40489);
or U41688 (N_41688,N_40927,N_40037);
xnor U41689 (N_41689,N_40333,N_40994);
and U41690 (N_41690,N_40689,N_40916);
nor U41691 (N_41691,N_40803,N_40115);
or U41692 (N_41692,N_40719,N_40248);
nand U41693 (N_41693,N_40837,N_40602);
nand U41694 (N_41694,N_40543,N_40869);
or U41695 (N_41695,N_40473,N_40559);
and U41696 (N_41696,N_40395,N_40956);
or U41697 (N_41697,N_40065,N_40592);
and U41698 (N_41698,N_40907,N_40125);
and U41699 (N_41699,N_40889,N_40247);
or U41700 (N_41700,N_40846,N_40523);
nor U41701 (N_41701,N_40057,N_40631);
nand U41702 (N_41702,N_40758,N_40229);
or U41703 (N_41703,N_40390,N_40270);
nand U41704 (N_41704,N_40245,N_40190);
nor U41705 (N_41705,N_40413,N_40005);
and U41706 (N_41706,N_40554,N_40953);
and U41707 (N_41707,N_40961,N_40519);
xnor U41708 (N_41708,N_40226,N_40024);
nand U41709 (N_41709,N_40110,N_40377);
or U41710 (N_41710,N_40605,N_40575);
or U41711 (N_41711,N_40812,N_40433);
and U41712 (N_41712,N_40463,N_40884);
and U41713 (N_41713,N_40673,N_40252);
or U41714 (N_41714,N_40330,N_40573);
nand U41715 (N_41715,N_40623,N_40067);
or U41716 (N_41716,N_40763,N_40932);
nor U41717 (N_41717,N_40460,N_40247);
or U41718 (N_41718,N_40241,N_40151);
xnor U41719 (N_41719,N_40006,N_40876);
xor U41720 (N_41720,N_40988,N_40233);
or U41721 (N_41721,N_40360,N_40075);
or U41722 (N_41722,N_40920,N_40300);
nand U41723 (N_41723,N_40930,N_40714);
or U41724 (N_41724,N_40943,N_40196);
nor U41725 (N_41725,N_40326,N_40322);
xor U41726 (N_41726,N_40578,N_40722);
or U41727 (N_41727,N_40669,N_40360);
or U41728 (N_41728,N_40230,N_40349);
and U41729 (N_41729,N_40218,N_40578);
and U41730 (N_41730,N_40405,N_40340);
and U41731 (N_41731,N_40563,N_40461);
nand U41732 (N_41732,N_40274,N_40247);
nor U41733 (N_41733,N_40581,N_40107);
and U41734 (N_41734,N_40344,N_40436);
or U41735 (N_41735,N_40693,N_40973);
nand U41736 (N_41736,N_40982,N_40933);
nand U41737 (N_41737,N_40706,N_40045);
nand U41738 (N_41738,N_40848,N_40351);
and U41739 (N_41739,N_40554,N_40015);
xnor U41740 (N_41740,N_40746,N_40222);
or U41741 (N_41741,N_40207,N_40319);
nand U41742 (N_41742,N_40671,N_40729);
and U41743 (N_41743,N_40612,N_40872);
nor U41744 (N_41744,N_40613,N_40440);
nand U41745 (N_41745,N_40318,N_40744);
and U41746 (N_41746,N_40956,N_40734);
nand U41747 (N_41747,N_40221,N_40235);
and U41748 (N_41748,N_40716,N_40375);
xnor U41749 (N_41749,N_40010,N_40601);
or U41750 (N_41750,N_40331,N_40129);
or U41751 (N_41751,N_40848,N_40678);
xnor U41752 (N_41752,N_40010,N_40927);
or U41753 (N_41753,N_40658,N_40622);
xor U41754 (N_41754,N_40072,N_40940);
nor U41755 (N_41755,N_40916,N_40595);
xor U41756 (N_41756,N_40878,N_40180);
nand U41757 (N_41757,N_40593,N_40648);
nand U41758 (N_41758,N_40376,N_40851);
xor U41759 (N_41759,N_40734,N_40323);
xnor U41760 (N_41760,N_40943,N_40633);
nor U41761 (N_41761,N_40880,N_40968);
nor U41762 (N_41762,N_40043,N_40499);
nor U41763 (N_41763,N_40725,N_40908);
nand U41764 (N_41764,N_40141,N_40177);
nor U41765 (N_41765,N_40895,N_40417);
or U41766 (N_41766,N_40707,N_40860);
xnor U41767 (N_41767,N_40444,N_40036);
nand U41768 (N_41768,N_40008,N_40699);
or U41769 (N_41769,N_40437,N_40761);
nand U41770 (N_41770,N_40180,N_40961);
nand U41771 (N_41771,N_40397,N_40214);
xor U41772 (N_41772,N_40775,N_40719);
nor U41773 (N_41773,N_40702,N_40345);
nor U41774 (N_41774,N_40705,N_40873);
nor U41775 (N_41775,N_40022,N_40140);
xor U41776 (N_41776,N_40167,N_40738);
and U41777 (N_41777,N_40515,N_40987);
xor U41778 (N_41778,N_40974,N_40851);
xor U41779 (N_41779,N_40148,N_40212);
or U41780 (N_41780,N_40351,N_40630);
nand U41781 (N_41781,N_40167,N_40667);
nand U41782 (N_41782,N_40769,N_40745);
or U41783 (N_41783,N_40485,N_40088);
nor U41784 (N_41784,N_40089,N_40280);
xnor U41785 (N_41785,N_40146,N_40448);
and U41786 (N_41786,N_40573,N_40812);
nor U41787 (N_41787,N_40359,N_40074);
and U41788 (N_41788,N_40980,N_40958);
nand U41789 (N_41789,N_40869,N_40263);
nor U41790 (N_41790,N_40927,N_40934);
xor U41791 (N_41791,N_40494,N_40492);
nand U41792 (N_41792,N_40935,N_40161);
nor U41793 (N_41793,N_40044,N_40780);
nand U41794 (N_41794,N_40101,N_40181);
or U41795 (N_41795,N_40090,N_40903);
nor U41796 (N_41796,N_40409,N_40448);
xnor U41797 (N_41797,N_40785,N_40510);
xnor U41798 (N_41798,N_40345,N_40590);
nor U41799 (N_41799,N_40255,N_40854);
and U41800 (N_41800,N_40115,N_40498);
xor U41801 (N_41801,N_40376,N_40690);
xnor U41802 (N_41802,N_40187,N_40947);
nor U41803 (N_41803,N_40904,N_40313);
or U41804 (N_41804,N_40564,N_40915);
xnor U41805 (N_41805,N_40065,N_40399);
or U41806 (N_41806,N_40849,N_40845);
or U41807 (N_41807,N_40079,N_40019);
nor U41808 (N_41808,N_40950,N_40815);
and U41809 (N_41809,N_40047,N_40652);
or U41810 (N_41810,N_40472,N_40709);
nand U41811 (N_41811,N_40834,N_40458);
nand U41812 (N_41812,N_40612,N_40147);
nor U41813 (N_41813,N_40124,N_40011);
nand U41814 (N_41814,N_40924,N_40342);
nand U41815 (N_41815,N_40787,N_40689);
xnor U41816 (N_41816,N_40841,N_40501);
nand U41817 (N_41817,N_40301,N_40677);
and U41818 (N_41818,N_40059,N_40219);
or U41819 (N_41819,N_40064,N_40921);
or U41820 (N_41820,N_40352,N_40355);
nand U41821 (N_41821,N_40388,N_40461);
nand U41822 (N_41822,N_40285,N_40360);
nand U41823 (N_41823,N_40891,N_40282);
and U41824 (N_41824,N_40837,N_40711);
and U41825 (N_41825,N_40594,N_40283);
nor U41826 (N_41826,N_40949,N_40190);
xnor U41827 (N_41827,N_40077,N_40860);
and U41828 (N_41828,N_40813,N_40611);
or U41829 (N_41829,N_40197,N_40278);
and U41830 (N_41830,N_40029,N_40367);
xor U41831 (N_41831,N_40970,N_40413);
nor U41832 (N_41832,N_40508,N_40324);
nand U41833 (N_41833,N_40670,N_40383);
nor U41834 (N_41834,N_40947,N_40961);
nor U41835 (N_41835,N_40984,N_40909);
nand U41836 (N_41836,N_40498,N_40702);
nand U41837 (N_41837,N_40959,N_40556);
nand U41838 (N_41838,N_40600,N_40359);
nor U41839 (N_41839,N_40486,N_40853);
nand U41840 (N_41840,N_40782,N_40310);
xnor U41841 (N_41841,N_40029,N_40689);
xor U41842 (N_41842,N_40072,N_40036);
and U41843 (N_41843,N_40815,N_40651);
nor U41844 (N_41844,N_40250,N_40558);
xor U41845 (N_41845,N_40541,N_40503);
xnor U41846 (N_41846,N_40255,N_40889);
nor U41847 (N_41847,N_40046,N_40036);
or U41848 (N_41848,N_40290,N_40527);
nor U41849 (N_41849,N_40609,N_40551);
or U41850 (N_41850,N_40789,N_40649);
or U41851 (N_41851,N_40551,N_40008);
and U41852 (N_41852,N_40118,N_40771);
nand U41853 (N_41853,N_40755,N_40450);
and U41854 (N_41854,N_40373,N_40413);
or U41855 (N_41855,N_40696,N_40595);
nand U41856 (N_41856,N_40233,N_40362);
xor U41857 (N_41857,N_40926,N_40892);
nand U41858 (N_41858,N_40334,N_40508);
xnor U41859 (N_41859,N_40826,N_40089);
nand U41860 (N_41860,N_40952,N_40108);
or U41861 (N_41861,N_40138,N_40809);
nand U41862 (N_41862,N_40170,N_40018);
nand U41863 (N_41863,N_40786,N_40500);
nand U41864 (N_41864,N_40604,N_40901);
and U41865 (N_41865,N_40612,N_40869);
and U41866 (N_41866,N_40380,N_40491);
nor U41867 (N_41867,N_40699,N_40408);
nand U41868 (N_41868,N_40631,N_40754);
nor U41869 (N_41869,N_40612,N_40635);
and U41870 (N_41870,N_40668,N_40563);
or U41871 (N_41871,N_40639,N_40985);
and U41872 (N_41872,N_40431,N_40539);
nand U41873 (N_41873,N_40058,N_40152);
nand U41874 (N_41874,N_40751,N_40665);
nor U41875 (N_41875,N_40568,N_40978);
or U41876 (N_41876,N_40999,N_40243);
nor U41877 (N_41877,N_40876,N_40796);
xnor U41878 (N_41878,N_40512,N_40189);
and U41879 (N_41879,N_40298,N_40434);
nor U41880 (N_41880,N_40447,N_40670);
xor U41881 (N_41881,N_40965,N_40910);
or U41882 (N_41882,N_40959,N_40616);
xor U41883 (N_41883,N_40761,N_40687);
and U41884 (N_41884,N_40407,N_40224);
and U41885 (N_41885,N_40768,N_40805);
and U41886 (N_41886,N_40177,N_40274);
and U41887 (N_41887,N_40598,N_40237);
xor U41888 (N_41888,N_40276,N_40135);
or U41889 (N_41889,N_40604,N_40815);
nor U41890 (N_41890,N_40265,N_40868);
xor U41891 (N_41891,N_40591,N_40885);
and U41892 (N_41892,N_40088,N_40796);
xor U41893 (N_41893,N_40848,N_40716);
xnor U41894 (N_41894,N_40462,N_40224);
and U41895 (N_41895,N_40963,N_40790);
xnor U41896 (N_41896,N_40257,N_40666);
nand U41897 (N_41897,N_40578,N_40047);
nand U41898 (N_41898,N_40394,N_40209);
nor U41899 (N_41899,N_40157,N_40301);
nor U41900 (N_41900,N_40228,N_40015);
and U41901 (N_41901,N_40385,N_40107);
xor U41902 (N_41902,N_40177,N_40316);
nor U41903 (N_41903,N_40280,N_40974);
nand U41904 (N_41904,N_40637,N_40454);
xor U41905 (N_41905,N_40964,N_40990);
nor U41906 (N_41906,N_40220,N_40256);
and U41907 (N_41907,N_40807,N_40360);
xor U41908 (N_41908,N_40240,N_40211);
xnor U41909 (N_41909,N_40231,N_40479);
nor U41910 (N_41910,N_40176,N_40971);
nor U41911 (N_41911,N_40774,N_40900);
or U41912 (N_41912,N_40273,N_40266);
xnor U41913 (N_41913,N_40382,N_40377);
and U41914 (N_41914,N_40775,N_40477);
nand U41915 (N_41915,N_40108,N_40129);
xor U41916 (N_41916,N_40081,N_40929);
nand U41917 (N_41917,N_40471,N_40620);
nand U41918 (N_41918,N_40893,N_40145);
and U41919 (N_41919,N_40698,N_40245);
xor U41920 (N_41920,N_40144,N_40889);
nand U41921 (N_41921,N_40138,N_40079);
or U41922 (N_41922,N_40858,N_40905);
and U41923 (N_41923,N_40704,N_40319);
and U41924 (N_41924,N_40339,N_40184);
nand U41925 (N_41925,N_40381,N_40419);
nor U41926 (N_41926,N_40065,N_40846);
nand U41927 (N_41927,N_40817,N_40667);
and U41928 (N_41928,N_40444,N_40445);
nand U41929 (N_41929,N_40170,N_40646);
nand U41930 (N_41930,N_40414,N_40927);
nand U41931 (N_41931,N_40318,N_40393);
and U41932 (N_41932,N_40616,N_40480);
and U41933 (N_41933,N_40830,N_40801);
or U41934 (N_41934,N_40098,N_40506);
xnor U41935 (N_41935,N_40597,N_40471);
or U41936 (N_41936,N_40399,N_40031);
or U41937 (N_41937,N_40801,N_40440);
xor U41938 (N_41938,N_40602,N_40591);
nor U41939 (N_41939,N_40117,N_40934);
xnor U41940 (N_41940,N_40576,N_40819);
and U41941 (N_41941,N_40040,N_40374);
xnor U41942 (N_41942,N_40996,N_40021);
or U41943 (N_41943,N_40195,N_40080);
nor U41944 (N_41944,N_40559,N_40668);
nand U41945 (N_41945,N_40862,N_40451);
xnor U41946 (N_41946,N_40591,N_40113);
xnor U41947 (N_41947,N_40593,N_40399);
nor U41948 (N_41948,N_40497,N_40543);
nor U41949 (N_41949,N_40765,N_40191);
xor U41950 (N_41950,N_40578,N_40857);
or U41951 (N_41951,N_40520,N_40632);
xnor U41952 (N_41952,N_40674,N_40358);
and U41953 (N_41953,N_40280,N_40474);
nor U41954 (N_41954,N_40833,N_40217);
xnor U41955 (N_41955,N_40006,N_40024);
or U41956 (N_41956,N_40637,N_40664);
xnor U41957 (N_41957,N_40476,N_40855);
nor U41958 (N_41958,N_40500,N_40358);
and U41959 (N_41959,N_40312,N_40660);
or U41960 (N_41960,N_40452,N_40061);
nor U41961 (N_41961,N_40412,N_40853);
and U41962 (N_41962,N_40744,N_40101);
nor U41963 (N_41963,N_40741,N_40443);
or U41964 (N_41964,N_40311,N_40872);
xor U41965 (N_41965,N_40813,N_40883);
and U41966 (N_41966,N_40150,N_40317);
or U41967 (N_41967,N_40155,N_40069);
and U41968 (N_41968,N_40802,N_40859);
or U41969 (N_41969,N_40087,N_40319);
xnor U41970 (N_41970,N_40921,N_40866);
nand U41971 (N_41971,N_40922,N_40151);
or U41972 (N_41972,N_40486,N_40033);
or U41973 (N_41973,N_40265,N_40514);
or U41974 (N_41974,N_40978,N_40336);
and U41975 (N_41975,N_40905,N_40520);
xor U41976 (N_41976,N_40479,N_40761);
or U41977 (N_41977,N_40762,N_40827);
nor U41978 (N_41978,N_40211,N_40823);
nor U41979 (N_41979,N_40461,N_40255);
nor U41980 (N_41980,N_40772,N_40847);
or U41981 (N_41981,N_40472,N_40364);
or U41982 (N_41982,N_40896,N_40307);
xor U41983 (N_41983,N_40421,N_40642);
and U41984 (N_41984,N_40923,N_40274);
or U41985 (N_41985,N_40627,N_40844);
nor U41986 (N_41986,N_40411,N_40314);
or U41987 (N_41987,N_40123,N_40998);
and U41988 (N_41988,N_40924,N_40580);
nor U41989 (N_41989,N_40524,N_40212);
xor U41990 (N_41990,N_40487,N_40528);
or U41991 (N_41991,N_40838,N_40124);
nand U41992 (N_41992,N_40631,N_40795);
nor U41993 (N_41993,N_40984,N_40125);
nor U41994 (N_41994,N_40341,N_40642);
xnor U41995 (N_41995,N_40254,N_40552);
xnor U41996 (N_41996,N_40994,N_40291);
or U41997 (N_41997,N_40804,N_40175);
or U41998 (N_41998,N_40066,N_40668);
nand U41999 (N_41999,N_40323,N_40251);
xnor U42000 (N_42000,N_41598,N_41370);
xor U42001 (N_42001,N_41941,N_41653);
and U42002 (N_42002,N_41338,N_41620);
or U42003 (N_42003,N_41515,N_41557);
and U42004 (N_42004,N_41851,N_41174);
xor U42005 (N_42005,N_41177,N_41938);
nor U42006 (N_42006,N_41816,N_41696);
and U42007 (N_42007,N_41982,N_41301);
nor U42008 (N_42008,N_41670,N_41424);
and U42009 (N_42009,N_41224,N_41155);
nor U42010 (N_42010,N_41541,N_41498);
or U42011 (N_42011,N_41256,N_41580);
nor U42012 (N_42012,N_41343,N_41025);
or U42013 (N_42013,N_41348,N_41698);
nand U42014 (N_42014,N_41173,N_41278);
and U42015 (N_42015,N_41780,N_41464);
nor U42016 (N_42016,N_41112,N_41877);
and U42017 (N_42017,N_41794,N_41054);
nand U42018 (N_42018,N_41164,N_41907);
and U42019 (N_42019,N_41835,N_41600);
nand U42020 (N_42020,N_41086,N_41789);
and U42021 (N_42021,N_41657,N_41380);
and U42022 (N_42022,N_41355,N_41171);
xnor U42023 (N_42023,N_41477,N_41300);
and U42024 (N_42024,N_41944,N_41373);
or U42025 (N_42025,N_41248,N_41975);
or U42026 (N_42026,N_41873,N_41189);
or U42027 (N_42027,N_41628,N_41429);
and U42028 (N_42028,N_41209,N_41716);
xor U42029 (N_42029,N_41753,N_41317);
and U42030 (N_42030,N_41798,N_41947);
nand U42031 (N_42031,N_41743,N_41267);
or U42032 (N_42032,N_41096,N_41900);
or U42033 (N_42033,N_41455,N_41147);
and U42034 (N_42034,N_41148,N_41239);
xor U42035 (N_42035,N_41472,N_41140);
xor U42036 (N_42036,N_41074,N_41020);
nand U42037 (N_42037,N_41918,N_41956);
xor U42038 (N_42038,N_41690,N_41245);
or U42039 (N_42039,N_41230,N_41058);
and U42040 (N_42040,N_41970,N_41269);
and U42041 (N_42041,N_41930,N_41675);
and U42042 (N_42042,N_41638,N_41759);
nor U42043 (N_42043,N_41181,N_41803);
or U42044 (N_42044,N_41559,N_41687);
or U42045 (N_42045,N_41917,N_41099);
xor U42046 (N_42046,N_41492,N_41972);
nand U42047 (N_42047,N_41506,N_41996);
nor U42048 (N_42048,N_41097,N_41481);
nor U42049 (N_42049,N_41289,N_41280);
and U42050 (N_42050,N_41213,N_41735);
nand U42051 (N_42051,N_41952,N_41118);
xnor U42052 (N_42052,N_41190,N_41881);
xor U42053 (N_42053,N_41644,N_41511);
or U42054 (N_42054,N_41457,N_41346);
xor U42055 (N_42055,N_41402,N_41252);
nor U42056 (N_42056,N_41535,N_41195);
and U42057 (N_42057,N_41840,N_41616);
xor U42058 (N_42058,N_41255,N_41612);
nor U42059 (N_42059,N_41888,N_41211);
or U42060 (N_42060,N_41218,N_41825);
xor U42061 (N_42061,N_41351,N_41114);
xor U42062 (N_42062,N_41078,N_41981);
and U42063 (N_42063,N_41850,N_41805);
and U42064 (N_42064,N_41589,N_41066);
nand U42065 (N_42065,N_41408,N_41971);
and U42066 (N_42066,N_41852,N_41369);
nor U42067 (N_42067,N_41647,N_41602);
and U42068 (N_42068,N_41809,N_41146);
and U42069 (N_42069,N_41861,N_41622);
xor U42070 (N_42070,N_41503,N_41661);
and U42071 (N_42071,N_41166,N_41621);
nand U42072 (N_42072,N_41636,N_41340);
and U42073 (N_42073,N_41185,N_41491);
nor U42074 (N_42074,N_41531,N_41694);
or U42075 (N_42075,N_41282,N_41225);
nor U42076 (N_42076,N_41149,N_41766);
or U42077 (N_42077,N_41257,N_41920);
or U42078 (N_42078,N_41067,N_41308);
nor U42079 (N_42079,N_41395,N_41710);
or U42080 (N_42080,N_41847,N_41795);
and U42081 (N_42081,N_41111,N_41427);
and U42082 (N_42082,N_41757,N_41456);
or U42083 (N_42083,N_41201,N_41529);
nor U42084 (N_42084,N_41057,N_41889);
and U42085 (N_42085,N_41823,N_41948);
nor U42086 (N_42086,N_41957,N_41186);
xnor U42087 (N_42087,N_41534,N_41578);
nor U42088 (N_42088,N_41352,N_41490);
and U42089 (N_42089,N_41782,N_41232);
and U42090 (N_42090,N_41431,N_41196);
xnor U42091 (N_42091,N_41231,N_41188);
nand U42092 (N_42092,N_41311,N_41389);
and U42093 (N_42093,N_41765,N_41295);
nand U42094 (N_42094,N_41413,N_41671);
and U42095 (N_42095,N_41502,N_41379);
or U42096 (N_42096,N_41932,N_41206);
xnor U42097 (N_42097,N_41946,N_41375);
and U42098 (N_42098,N_41162,N_41762);
xor U42099 (N_42099,N_41899,N_41144);
xnor U42100 (N_42100,N_41568,N_41163);
nor U42101 (N_42101,N_41995,N_41629);
xor U42102 (N_42102,N_41951,N_41715);
nand U42103 (N_42103,N_41411,N_41243);
or U42104 (N_42104,N_41180,N_41482);
nand U42105 (N_42105,N_41279,N_41247);
or U42106 (N_42106,N_41294,N_41228);
xor U42107 (N_42107,N_41770,N_41922);
and U42108 (N_42108,N_41980,N_41883);
and U42109 (N_42109,N_41198,N_41599);
and U42110 (N_42110,N_41539,N_41626);
nand U42111 (N_42111,N_41959,N_41746);
xnor U42112 (N_42112,N_41550,N_41409);
nor U42113 (N_42113,N_41242,N_41912);
xnor U42114 (N_42114,N_41864,N_41854);
nor U42115 (N_42115,N_41674,N_41719);
or U42116 (N_42116,N_41420,N_41625);
and U42117 (N_42117,N_41652,N_41070);
nor U42118 (N_42118,N_41082,N_41736);
nor U42119 (N_42119,N_41264,N_41662);
and U42120 (N_42120,N_41226,N_41128);
or U42121 (N_42121,N_41812,N_41993);
or U42122 (N_42122,N_41131,N_41569);
nand U42123 (N_42123,N_41042,N_41838);
xor U42124 (N_42124,N_41421,N_41500);
and U42125 (N_42125,N_41358,N_41940);
xnor U42126 (N_42126,N_41634,N_41479);
xnor U42127 (N_42127,N_41771,N_41718);
xnor U42128 (N_42128,N_41648,N_41315);
and U42129 (N_42129,N_41514,N_41032);
and U42130 (N_42130,N_41513,N_41640);
and U42131 (N_42131,N_41496,N_41035);
xnor U42132 (N_42132,N_41867,N_41229);
xnor U42133 (N_42133,N_41385,N_41688);
or U42134 (N_42134,N_41274,N_41281);
and U42135 (N_42135,N_41565,N_41160);
and U42136 (N_42136,N_41808,N_41319);
nand U42137 (N_42137,N_41566,N_41637);
and U42138 (N_42138,N_41132,N_41283);
nor U42139 (N_42139,N_41724,N_41656);
xor U42140 (N_42140,N_41183,N_41799);
xnor U42141 (N_42141,N_41756,N_41235);
xor U42142 (N_42142,N_41702,N_41588);
or U42143 (N_42143,N_41334,N_41775);
and U42144 (N_42144,N_41668,N_41894);
xnor U42145 (N_42145,N_41669,N_41158);
and U42146 (N_42146,N_41543,N_41448);
nor U42147 (N_42147,N_41037,N_41459);
nor U42148 (N_42148,N_41890,N_41141);
xnor U42149 (N_42149,N_41341,N_41992);
xor U42150 (N_42150,N_41570,N_41839);
nor U42151 (N_42151,N_41489,N_41695);
and U42152 (N_42152,N_41773,N_41071);
and U42153 (N_42153,N_41501,N_41246);
or U42154 (N_42154,N_41707,N_41837);
or U42155 (N_42155,N_41592,N_41654);
nand U42156 (N_42156,N_41574,N_41085);
or U42157 (N_42157,N_41567,N_41007);
or U42158 (N_42158,N_41785,N_41857);
or U42159 (N_42159,N_41721,N_41265);
or U42160 (N_42160,N_41874,N_41296);
and U42161 (N_42161,N_41404,N_41223);
nand U42162 (N_42162,N_41764,N_41792);
nand U42163 (N_42163,N_41901,N_41813);
and U42164 (N_42164,N_41554,N_41556);
and U42165 (N_42165,N_41540,N_41415);
or U42166 (N_42166,N_41327,N_41023);
xor U42167 (N_42167,N_41328,N_41614);
nor U42168 (N_42168,N_41056,N_41843);
nor U42169 (N_42169,N_41649,N_41494);
nor U42170 (N_42170,N_41088,N_41509);
nor U42171 (N_42171,N_41987,N_41488);
and U42172 (N_42172,N_41525,N_41005);
nor U42173 (N_42173,N_41989,N_41030);
and U42174 (N_42174,N_41277,N_41898);
nand U42175 (N_42175,N_41329,N_41318);
and U42176 (N_42176,N_41471,N_41965);
nand U42177 (N_42177,N_41312,N_41586);
xnor U42178 (N_42178,N_41806,N_41768);
nor U42179 (N_42179,N_41682,N_41214);
and U42180 (N_42180,N_41862,N_41168);
xnor U42181 (N_42181,N_41110,N_41821);
nor U42182 (N_42182,N_41444,N_41828);
and U42183 (N_42183,N_41394,N_41137);
nor U42184 (N_42184,N_41655,N_41686);
xor U42185 (N_42185,N_41609,N_41572);
xor U42186 (N_42186,N_41933,N_41726);
nor U42187 (N_42187,N_41276,N_41422);
nand U42188 (N_42188,N_41522,N_41776);
and U42189 (N_42189,N_41432,N_41596);
and U42190 (N_42190,N_41203,N_41884);
nand U42191 (N_42191,N_41019,N_41967);
xnor U42192 (N_42192,N_41306,N_41018);
or U42193 (N_42193,N_41635,N_41752);
or U42194 (N_42194,N_41446,N_41016);
and U42195 (N_42195,N_41709,N_41673);
xnor U42196 (N_42196,N_41055,N_41363);
xnor U42197 (N_42197,N_41704,N_41299);
xor U42198 (N_42198,N_41610,N_41049);
and U42199 (N_42199,N_41259,N_41191);
nand U42200 (N_42200,N_41512,N_41858);
and U42201 (N_42201,N_41953,N_41676);
nand U42202 (N_42202,N_41094,N_41630);
nor U42203 (N_42203,N_41357,N_41065);
xnor U42204 (N_42204,N_41095,N_41476);
or U42205 (N_42205,N_41571,N_41663);
and U42206 (N_42206,N_41107,N_41439);
nor U42207 (N_42207,N_41249,N_41273);
nand U42208 (N_42208,N_41542,N_41154);
or U42209 (N_42209,N_41712,N_41216);
nor U42210 (N_42210,N_41205,N_41855);
nand U42211 (N_42211,N_41084,N_41935);
nand U42212 (N_42212,N_41466,N_41961);
nor U42213 (N_42213,N_41820,N_41014);
or U42214 (N_42214,N_41558,N_41165);
and U42215 (N_42215,N_41923,N_41270);
nor U42216 (N_42216,N_41790,N_41703);
or U42217 (N_42217,N_41193,N_41116);
xor U42218 (N_42218,N_41560,N_41927);
nor U42219 (N_42219,N_41928,N_41774);
nand U42220 (N_42220,N_41555,N_41182);
nor U42221 (N_42221,N_41842,N_41293);
xor U42222 (N_42222,N_41802,N_41659);
nand U42223 (N_42223,N_41606,N_41916);
xnor U42224 (N_42224,N_41848,N_41263);
and U42225 (N_42225,N_41639,N_41123);
or U42226 (N_42226,N_41344,N_41129);
nor U42227 (N_42227,N_41119,N_41079);
nand U42228 (N_42228,N_41650,N_41692);
xnor U42229 (N_42229,N_41860,N_41262);
xnor U42230 (N_42230,N_41321,N_41038);
xnor U42231 (N_42231,N_41031,N_41573);
or U42232 (N_42232,N_41331,N_41194);
xnor U42233 (N_42233,N_41651,N_41966);
xor U42234 (N_42234,N_41210,N_41913);
and U42235 (N_42235,N_41043,N_41000);
and U42236 (N_42236,N_41760,N_41997);
nor U42237 (N_42237,N_41608,N_41978);
or U42238 (N_42238,N_41749,N_41495);
and U42239 (N_42239,N_41977,N_41865);
nor U42240 (N_42240,N_41863,N_41903);
or U42241 (N_42241,N_41791,N_41271);
nor U42242 (N_42242,N_41219,N_41544);
xor U42243 (N_42243,N_41098,N_41130);
or U42244 (N_42244,N_41125,N_41699);
nand U42245 (N_42245,N_41104,N_41062);
nor U42246 (N_42246,N_41335,N_41426);
nor U42247 (N_42247,N_41581,N_41151);
and U42248 (N_42248,N_41388,N_41212);
and U42249 (N_42249,N_41562,N_41442);
and U42250 (N_42250,N_41258,N_41347);
or U42251 (N_42251,N_41391,N_41002);
xor U42252 (N_42252,N_41367,N_41516);
or U42253 (N_42253,N_41725,N_41006);
xnor U42254 (N_42254,N_41458,N_41868);
xnor U42255 (N_42255,N_41800,N_41684);
nor U42256 (N_42256,N_41126,N_41763);
xor U42257 (N_42257,N_41430,N_41728);
and U42258 (N_42258,N_41607,N_41172);
nand U42259 (N_42259,N_41241,N_41632);
xor U42260 (N_42260,N_41666,N_41605);
nor U42261 (N_42261,N_41383,N_41199);
and U42262 (N_42262,N_41701,N_41063);
and U42263 (N_42263,N_41991,N_41026);
nor U42264 (N_42264,N_41286,N_41364);
xnor U42265 (N_42265,N_41325,N_41505);
nand U42266 (N_42266,N_41937,N_41410);
nand U42267 (N_42267,N_41885,N_41819);
and U42268 (N_42268,N_41804,N_41870);
xor U42269 (N_42269,N_41548,N_41115);
nand U42270 (N_42270,N_41679,N_41053);
nand U42271 (N_42271,N_41717,N_41484);
or U42272 (N_42272,N_41487,N_41538);
nor U42273 (N_42273,N_41117,N_41939);
xnor U42274 (N_42274,N_41577,N_41926);
and U42275 (N_42275,N_41135,N_41984);
nand U42276 (N_42276,N_41127,N_41817);
xor U42277 (N_42277,N_41244,N_41170);
and U42278 (N_42278,N_41733,N_41504);
and U42279 (N_42279,N_41841,N_41075);
nand U42280 (N_42280,N_41934,N_41452);
nor U42281 (N_42281,N_41462,N_41093);
or U42282 (N_42282,N_41896,N_41371);
nand U42283 (N_42283,N_41121,N_41011);
and U42284 (N_42284,N_41138,N_41553);
or U42285 (N_42285,N_41474,N_41398);
and U42286 (N_42286,N_41473,N_41897);
or U42287 (N_42287,N_41323,N_41382);
nand U42288 (N_42288,N_41302,N_41526);
nand U42289 (N_42289,N_41366,N_41400);
xor U42290 (N_42290,N_41576,N_41027);
nand U42291 (N_42291,N_41354,N_41460);
or U42292 (N_42292,N_41983,N_41931);
and U42293 (N_42293,N_41092,N_41478);
xor U42294 (N_42294,N_41708,N_41386);
xnor U42295 (N_42295,N_41461,N_41184);
xnor U42296 (N_42296,N_41664,N_41958);
nand U42297 (N_42297,N_41960,N_41309);
nand U42298 (N_42298,N_41849,N_41012);
and U42299 (N_42299,N_41611,N_41204);
or U42300 (N_42300,N_41872,N_41061);
and U42301 (N_42301,N_41254,N_41374);
and U42302 (N_42302,N_41748,N_41875);
and U42303 (N_42303,N_41985,N_41046);
nand U42304 (N_42304,N_41642,N_41833);
nand U42305 (N_42305,N_41905,N_41152);
or U42306 (N_42306,N_41705,N_41167);
nand U42307 (N_42307,N_41683,N_41585);
and U42308 (N_42308,N_41040,N_41830);
xnor U42309 (N_42309,N_41113,N_41266);
or U42310 (N_42310,N_41832,N_41986);
xnor U42311 (N_42311,N_41039,N_41545);
xor U42312 (N_42312,N_41250,N_41467);
or U42313 (N_42313,N_41624,N_41449);
or U42314 (N_42314,N_41313,N_41051);
nand U42315 (N_42315,N_41807,N_41024);
nor U42316 (N_42316,N_41551,N_41142);
nor U42317 (N_42317,N_41416,N_41356);
or U42318 (N_42318,N_41595,N_41594);
or U42319 (N_42319,N_41010,N_41015);
and U42320 (N_42320,N_41779,N_41451);
xnor U42321 (N_42321,N_41200,N_41290);
nand U42322 (N_42322,N_41059,N_41909);
nor U42323 (N_42323,N_41758,N_41326);
or U42324 (N_42324,N_41742,N_41237);
xor U42325 (N_42325,N_41999,N_41134);
xor U42326 (N_42326,N_41829,N_41822);
and U42327 (N_42327,N_41387,N_41564);
nor U42328 (N_42328,N_41929,N_41122);
and U42329 (N_42329,N_41871,N_41485);
nand U42330 (N_42330,N_41349,N_41103);
or U42331 (N_42331,N_41310,N_41150);
xor U42332 (N_42332,N_41305,N_41597);
xor U42333 (N_42333,N_41994,N_41463);
or U42334 (N_42334,N_41145,N_41251);
and U42335 (N_42335,N_41272,N_41445);
or U42336 (N_42336,N_41962,N_41836);
xor U42337 (N_42337,N_41723,N_41510);
nand U42338 (N_42338,N_41493,N_41261);
or U42339 (N_42339,N_41083,N_41175);
and U42340 (N_42340,N_41453,N_41672);
nor U42341 (N_42341,N_41869,N_41641);
nor U42342 (N_42342,N_41304,N_41009);
nand U42343 (N_42343,N_41781,N_41797);
nand U42344 (N_42344,N_41633,N_41827);
and U42345 (N_42345,N_41973,N_41613);
and U42346 (N_42346,N_41552,N_41745);
xor U42347 (N_42347,N_41465,N_41217);
xnor U42348 (N_42348,N_41811,N_41017);
and U42349 (N_42349,N_41751,N_41974);
and U42350 (N_42350,N_41615,N_41969);
xor U42351 (N_42351,N_41072,N_41878);
or U42352 (N_42352,N_41480,N_41603);
and U42353 (N_42353,N_41895,N_41810);
or U42354 (N_42354,N_41631,N_41524);
nor U42355 (N_42355,N_41440,N_41866);
xnor U42356 (N_42356,N_41178,N_41443);
nor U42357 (N_42357,N_41845,N_41976);
xnor U42358 (N_42358,N_41236,N_41406);
and U42359 (N_42359,N_41815,N_41988);
nor U42360 (N_42360,N_41441,N_41508);
and U42361 (N_42361,N_41073,N_41234);
nand U42362 (N_42362,N_41579,N_41793);
or U42363 (N_42363,N_41192,N_41530);
nor U42364 (N_42364,N_41108,N_41880);
or U42365 (N_42365,N_41914,N_41739);
and U42366 (N_42366,N_41680,N_41052);
nand U42367 (N_42367,N_41253,N_41519);
nor U42368 (N_42368,N_41392,N_41527);
nand U42369 (N_42369,N_41220,N_41968);
nand U42370 (N_42370,N_41617,N_41143);
xor U42371 (N_42371,N_41001,N_41233);
and U42372 (N_42372,N_41499,N_41412);
nand U42373 (N_42373,N_41711,N_41433);
xnor U42374 (N_42374,N_41518,N_41755);
or U42375 (N_42375,N_41998,N_41068);
or U42376 (N_42376,N_41081,N_41906);
nand U42377 (N_42377,N_41322,N_41731);
nand U42378 (N_42378,N_41292,N_41425);
or U42379 (N_42379,N_41238,N_41284);
and U42380 (N_42380,N_41853,N_41824);
nor U42381 (N_42381,N_41050,N_41008);
nand U42382 (N_42382,N_41330,N_41393);
nor U42383 (N_42383,N_41590,N_41750);
nand U42384 (N_42384,N_41777,N_41438);
and U42385 (N_42385,N_41423,N_41507);
or U42386 (N_42386,N_41036,N_41563);
and U42387 (N_42387,N_41646,N_41450);
xor U42388 (N_42388,N_41483,N_41908);
xnor U42389 (N_42389,N_41044,N_41660);
and U42390 (N_42390,N_41950,N_41399);
nor U42391 (N_42391,N_41287,N_41623);
nand U42392 (N_42392,N_41727,N_41744);
xor U42393 (N_42393,N_41834,N_41910);
xor U42394 (N_42394,N_41076,N_41090);
xor U42395 (N_42395,N_41936,N_41796);
and U42396 (N_42396,N_41697,N_41197);
or U42397 (N_42397,N_41333,N_41619);
and U42398 (N_42398,N_41497,N_41990);
or U42399 (N_42399,N_41921,N_41732);
nor U42400 (N_42400,N_41060,N_41911);
nand U42401 (N_42401,N_41080,N_41643);
nand U42402 (N_42402,N_41470,N_41893);
or U42403 (N_42403,N_41136,N_41691);
xnor U42404 (N_42404,N_41202,N_41887);
and U42405 (N_42405,N_41100,N_41353);
xnor U42406 (N_42406,N_41437,N_41943);
or U42407 (N_42407,N_41316,N_41260);
and U42408 (N_42408,N_41077,N_41741);
and U42409 (N_42409,N_41778,N_41285);
and U42410 (N_42410,N_41298,N_41275);
nand U42411 (N_42411,N_41783,N_41362);
nand U42412 (N_42412,N_41720,N_41291);
nand U42413 (N_42413,N_41013,N_41713);
or U42414 (N_42414,N_41734,N_41029);
or U42415 (N_42415,N_41879,N_41361);
or U42416 (N_42416,N_41109,N_41368);
nand U42417 (N_42417,N_41157,N_41475);
and U42418 (N_42418,N_41949,N_41786);
nor U42419 (N_42419,N_41468,N_41658);
nor U42420 (N_42420,N_41737,N_41583);
or U42421 (N_42421,N_41892,N_41376);
xnor U42422 (N_42422,N_41963,N_41390);
nor U42423 (N_42423,N_41179,N_41447);
and U42424 (N_42424,N_41268,N_41722);
xor U42425 (N_42425,N_41520,N_41549);
xnor U42426 (N_42426,N_41045,N_41955);
xor U42427 (N_42427,N_41297,N_41919);
or U42428 (N_42428,N_41378,N_41034);
nor U42429 (N_42429,N_41332,N_41339);
nor U42430 (N_42430,N_41324,N_41593);
xnor U42431 (N_42431,N_41693,N_41730);
or U42432 (N_42432,N_41105,N_41207);
xnor U42433 (N_42433,N_41587,N_41767);
and U42434 (N_42434,N_41945,N_41665);
nor U42435 (N_42435,N_41729,N_41288);
or U42436 (N_42436,N_41436,N_41964);
or U42437 (N_42437,N_41831,N_41384);
nand U42438 (N_42438,N_41915,N_41153);
and U42439 (N_42439,N_41396,N_41754);
nand U42440 (N_42440,N_41582,N_41761);
xor U42441 (N_42441,N_41882,N_41547);
nand U42442 (N_42442,N_41747,N_41350);
xnor U42443 (N_42443,N_41517,N_41575);
nand U42444 (N_42444,N_41047,N_41004);
or U42445 (N_42445,N_41414,N_41365);
nand U42446 (N_42446,N_41801,N_41561);
nand U42447 (N_42447,N_41069,N_41700);
and U42448 (N_42448,N_41091,N_41064);
nor U42449 (N_42449,N_41022,N_41418);
nor U42450 (N_42450,N_41601,N_41401);
xnor U42451 (N_42451,N_41089,N_41859);
or U42452 (N_42452,N_41738,N_41902);
or U42453 (N_42453,N_41156,N_41667);
and U42454 (N_42454,N_41904,N_41689);
nor U42455 (N_42455,N_41087,N_41533);
nand U42456 (N_42456,N_41604,N_41714);
and U42457 (N_42457,N_41407,N_41124);
nand U42458 (N_42458,N_41048,N_41788);
or U42459 (N_42459,N_41546,N_41215);
or U42460 (N_42460,N_41954,N_41314);
nand U42461 (N_42461,N_41924,N_41307);
nor U42462 (N_42462,N_41886,N_41337);
and U42463 (N_42463,N_41176,N_41856);
nor U42464 (N_42464,N_41120,N_41161);
nor U42465 (N_42465,N_41360,N_41033);
xor U42466 (N_42466,N_41101,N_41784);
and U42467 (N_42467,N_41685,N_41320);
nand U42468 (N_42468,N_41627,N_41706);
nor U42469 (N_42469,N_41221,N_41405);
nor U42470 (N_42470,N_41826,N_41486);
nand U42471 (N_42471,N_41469,N_41041);
nand U42472 (N_42472,N_41342,N_41532);
nor U42473 (N_42473,N_41979,N_41187);
or U42474 (N_42474,N_41677,N_41345);
xnor U42475 (N_42475,N_41133,N_41102);
nor U42476 (N_42476,N_41521,N_41419);
and U42477 (N_42477,N_41106,N_41222);
xor U42478 (N_42478,N_41435,N_41227);
or U42479 (N_42479,N_41159,N_41536);
nand U42480 (N_42480,N_41303,N_41240);
and U42481 (N_42481,N_41769,N_41403);
and U42482 (N_42482,N_41814,N_41925);
and U42483 (N_42483,N_41876,N_41678);
and U42484 (N_42484,N_41381,N_41740);
nand U42485 (N_42485,N_41428,N_41681);
nand U42486 (N_42486,N_41772,N_41359);
or U42487 (N_42487,N_41787,N_41021);
and U42488 (N_42488,N_41537,N_41891);
nor U42489 (N_42489,N_41434,N_41454);
nor U42490 (N_42490,N_41645,N_41028);
or U42491 (N_42491,N_41372,N_41377);
nor U42492 (N_42492,N_41844,N_41584);
xor U42493 (N_42493,N_41591,N_41528);
xor U42494 (N_42494,N_41208,N_41942);
xnor U42495 (N_42495,N_41846,N_41336);
or U42496 (N_42496,N_41397,N_41139);
xor U42497 (N_42497,N_41818,N_41523);
or U42498 (N_42498,N_41003,N_41169);
xor U42499 (N_42499,N_41417,N_41618);
nand U42500 (N_42500,N_41097,N_41887);
and U42501 (N_42501,N_41693,N_41716);
and U42502 (N_42502,N_41904,N_41385);
xnor U42503 (N_42503,N_41238,N_41171);
and U42504 (N_42504,N_41524,N_41411);
xor U42505 (N_42505,N_41754,N_41320);
or U42506 (N_42506,N_41787,N_41096);
xor U42507 (N_42507,N_41927,N_41829);
xor U42508 (N_42508,N_41677,N_41725);
xnor U42509 (N_42509,N_41704,N_41317);
nand U42510 (N_42510,N_41530,N_41089);
xnor U42511 (N_42511,N_41178,N_41785);
or U42512 (N_42512,N_41811,N_41238);
or U42513 (N_42513,N_41023,N_41200);
nand U42514 (N_42514,N_41980,N_41578);
nor U42515 (N_42515,N_41813,N_41899);
nand U42516 (N_42516,N_41194,N_41802);
nand U42517 (N_42517,N_41670,N_41076);
or U42518 (N_42518,N_41377,N_41091);
nand U42519 (N_42519,N_41446,N_41987);
and U42520 (N_42520,N_41908,N_41175);
xnor U42521 (N_42521,N_41344,N_41474);
xor U42522 (N_42522,N_41177,N_41011);
or U42523 (N_42523,N_41460,N_41953);
nand U42524 (N_42524,N_41494,N_41879);
or U42525 (N_42525,N_41232,N_41795);
xnor U42526 (N_42526,N_41173,N_41258);
xnor U42527 (N_42527,N_41430,N_41493);
or U42528 (N_42528,N_41599,N_41449);
and U42529 (N_42529,N_41626,N_41054);
nand U42530 (N_42530,N_41109,N_41331);
nor U42531 (N_42531,N_41326,N_41776);
xor U42532 (N_42532,N_41545,N_41553);
or U42533 (N_42533,N_41213,N_41591);
nand U42534 (N_42534,N_41581,N_41373);
nor U42535 (N_42535,N_41588,N_41649);
xor U42536 (N_42536,N_41926,N_41489);
and U42537 (N_42537,N_41375,N_41556);
xor U42538 (N_42538,N_41813,N_41054);
and U42539 (N_42539,N_41629,N_41010);
or U42540 (N_42540,N_41620,N_41881);
or U42541 (N_42541,N_41976,N_41414);
nor U42542 (N_42542,N_41534,N_41880);
xor U42543 (N_42543,N_41064,N_41341);
xnor U42544 (N_42544,N_41458,N_41584);
xnor U42545 (N_42545,N_41316,N_41330);
or U42546 (N_42546,N_41014,N_41252);
nand U42547 (N_42547,N_41254,N_41757);
and U42548 (N_42548,N_41785,N_41356);
xor U42549 (N_42549,N_41300,N_41623);
and U42550 (N_42550,N_41040,N_41206);
nand U42551 (N_42551,N_41645,N_41372);
xnor U42552 (N_42552,N_41679,N_41097);
and U42553 (N_42553,N_41809,N_41924);
nor U42554 (N_42554,N_41380,N_41032);
and U42555 (N_42555,N_41592,N_41174);
or U42556 (N_42556,N_41073,N_41208);
nor U42557 (N_42557,N_41507,N_41301);
and U42558 (N_42558,N_41265,N_41052);
or U42559 (N_42559,N_41155,N_41274);
and U42560 (N_42560,N_41658,N_41592);
nand U42561 (N_42561,N_41595,N_41649);
xor U42562 (N_42562,N_41807,N_41628);
and U42563 (N_42563,N_41457,N_41354);
and U42564 (N_42564,N_41076,N_41001);
nand U42565 (N_42565,N_41378,N_41366);
nand U42566 (N_42566,N_41063,N_41381);
nor U42567 (N_42567,N_41745,N_41191);
xnor U42568 (N_42568,N_41856,N_41077);
and U42569 (N_42569,N_41464,N_41441);
and U42570 (N_42570,N_41647,N_41561);
and U42571 (N_42571,N_41795,N_41639);
xnor U42572 (N_42572,N_41160,N_41911);
or U42573 (N_42573,N_41691,N_41960);
and U42574 (N_42574,N_41679,N_41964);
or U42575 (N_42575,N_41716,N_41856);
nand U42576 (N_42576,N_41480,N_41484);
nand U42577 (N_42577,N_41536,N_41002);
xnor U42578 (N_42578,N_41972,N_41955);
and U42579 (N_42579,N_41481,N_41366);
nand U42580 (N_42580,N_41779,N_41106);
nand U42581 (N_42581,N_41752,N_41190);
and U42582 (N_42582,N_41027,N_41351);
xor U42583 (N_42583,N_41769,N_41131);
nor U42584 (N_42584,N_41801,N_41325);
nand U42585 (N_42585,N_41795,N_41129);
nor U42586 (N_42586,N_41247,N_41602);
and U42587 (N_42587,N_41755,N_41568);
or U42588 (N_42588,N_41004,N_41293);
xor U42589 (N_42589,N_41058,N_41354);
xor U42590 (N_42590,N_41732,N_41714);
and U42591 (N_42591,N_41805,N_41257);
nand U42592 (N_42592,N_41142,N_41719);
nor U42593 (N_42593,N_41499,N_41826);
nand U42594 (N_42594,N_41670,N_41191);
nor U42595 (N_42595,N_41695,N_41843);
or U42596 (N_42596,N_41305,N_41881);
nand U42597 (N_42597,N_41141,N_41590);
nor U42598 (N_42598,N_41970,N_41464);
xnor U42599 (N_42599,N_41902,N_41380);
xor U42600 (N_42600,N_41666,N_41791);
and U42601 (N_42601,N_41538,N_41352);
xor U42602 (N_42602,N_41957,N_41137);
nor U42603 (N_42603,N_41569,N_41198);
nand U42604 (N_42604,N_41903,N_41037);
or U42605 (N_42605,N_41853,N_41604);
nor U42606 (N_42606,N_41385,N_41102);
or U42607 (N_42607,N_41047,N_41530);
or U42608 (N_42608,N_41193,N_41453);
nand U42609 (N_42609,N_41297,N_41461);
or U42610 (N_42610,N_41434,N_41421);
nor U42611 (N_42611,N_41918,N_41799);
and U42612 (N_42612,N_41000,N_41090);
xnor U42613 (N_42613,N_41347,N_41868);
xnor U42614 (N_42614,N_41906,N_41953);
xnor U42615 (N_42615,N_41143,N_41908);
xnor U42616 (N_42616,N_41059,N_41803);
or U42617 (N_42617,N_41735,N_41039);
or U42618 (N_42618,N_41416,N_41230);
or U42619 (N_42619,N_41793,N_41697);
and U42620 (N_42620,N_41544,N_41561);
nand U42621 (N_42621,N_41569,N_41379);
nor U42622 (N_42622,N_41404,N_41104);
nor U42623 (N_42623,N_41903,N_41559);
xnor U42624 (N_42624,N_41947,N_41926);
nor U42625 (N_42625,N_41720,N_41370);
or U42626 (N_42626,N_41744,N_41726);
and U42627 (N_42627,N_41800,N_41649);
nand U42628 (N_42628,N_41882,N_41185);
nor U42629 (N_42629,N_41127,N_41962);
and U42630 (N_42630,N_41745,N_41856);
and U42631 (N_42631,N_41055,N_41427);
and U42632 (N_42632,N_41360,N_41916);
or U42633 (N_42633,N_41946,N_41271);
or U42634 (N_42634,N_41541,N_41666);
xnor U42635 (N_42635,N_41434,N_41993);
xor U42636 (N_42636,N_41306,N_41427);
or U42637 (N_42637,N_41167,N_41372);
or U42638 (N_42638,N_41514,N_41285);
or U42639 (N_42639,N_41951,N_41803);
and U42640 (N_42640,N_41446,N_41796);
nor U42641 (N_42641,N_41135,N_41968);
xor U42642 (N_42642,N_41084,N_41462);
nor U42643 (N_42643,N_41664,N_41796);
xor U42644 (N_42644,N_41761,N_41802);
nor U42645 (N_42645,N_41223,N_41370);
xor U42646 (N_42646,N_41808,N_41711);
xnor U42647 (N_42647,N_41114,N_41558);
nor U42648 (N_42648,N_41479,N_41085);
nand U42649 (N_42649,N_41889,N_41754);
xor U42650 (N_42650,N_41911,N_41834);
and U42651 (N_42651,N_41326,N_41673);
xor U42652 (N_42652,N_41754,N_41191);
and U42653 (N_42653,N_41680,N_41565);
or U42654 (N_42654,N_41600,N_41524);
nor U42655 (N_42655,N_41238,N_41973);
xnor U42656 (N_42656,N_41273,N_41355);
and U42657 (N_42657,N_41633,N_41357);
and U42658 (N_42658,N_41412,N_41907);
xnor U42659 (N_42659,N_41557,N_41463);
nand U42660 (N_42660,N_41249,N_41286);
or U42661 (N_42661,N_41289,N_41599);
nand U42662 (N_42662,N_41714,N_41756);
nand U42663 (N_42663,N_41487,N_41720);
or U42664 (N_42664,N_41842,N_41752);
nand U42665 (N_42665,N_41733,N_41514);
and U42666 (N_42666,N_41617,N_41811);
or U42667 (N_42667,N_41256,N_41050);
nor U42668 (N_42668,N_41284,N_41370);
nand U42669 (N_42669,N_41021,N_41552);
or U42670 (N_42670,N_41511,N_41840);
nor U42671 (N_42671,N_41363,N_41313);
xor U42672 (N_42672,N_41095,N_41523);
xor U42673 (N_42673,N_41720,N_41161);
xnor U42674 (N_42674,N_41847,N_41727);
nand U42675 (N_42675,N_41277,N_41729);
nand U42676 (N_42676,N_41605,N_41894);
and U42677 (N_42677,N_41787,N_41439);
xnor U42678 (N_42678,N_41789,N_41202);
and U42679 (N_42679,N_41649,N_41613);
nor U42680 (N_42680,N_41415,N_41172);
nand U42681 (N_42681,N_41717,N_41592);
and U42682 (N_42682,N_41582,N_41061);
nor U42683 (N_42683,N_41839,N_41196);
or U42684 (N_42684,N_41112,N_41497);
and U42685 (N_42685,N_41392,N_41794);
and U42686 (N_42686,N_41901,N_41969);
nand U42687 (N_42687,N_41639,N_41218);
or U42688 (N_42688,N_41656,N_41722);
nand U42689 (N_42689,N_41728,N_41543);
and U42690 (N_42690,N_41502,N_41859);
xnor U42691 (N_42691,N_41657,N_41543);
nand U42692 (N_42692,N_41924,N_41458);
xnor U42693 (N_42693,N_41094,N_41868);
or U42694 (N_42694,N_41983,N_41518);
nand U42695 (N_42695,N_41281,N_41771);
xnor U42696 (N_42696,N_41294,N_41366);
xor U42697 (N_42697,N_41073,N_41147);
nor U42698 (N_42698,N_41156,N_41132);
xnor U42699 (N_42699,N_41659,N_41481);
or U42700 (N_42700,N_41858,N_41761);
xor U42701 (N_42701,N_41499,N_41815);
or U42702 (N_42702,N_41423,N_41984);
and U42703 (N_42703,N_41329,N_41861);
nor U42704 (N_42704,N_41238,N_41353);
and U42705 (N_42705,N_41953,N_41066);
xor U42706 (N_42706,N_41559,N_41312);
nand U42707 (N_42707,N_41324,N_41680);
xor U42708 (N_42708,N_41754,N_41842);
nand U42709 (N_42709,N_41453,N_41612);
and U42710 (N_42710,N_41057,N_41645);
nand U42711 (N_42711,N_41402,N_41289);
xnor U42712 (N_42712,N_41105,N_41366);
nor U42713 (N_42713,N_41990,N_41045);
xnor U42714 (N_42714,N_41342,N_41566);
and U42715 (N_42715,N_41139,N_41307);
xor U42716 (N_42716,N_41266,N_41561);
nand U42717 (N_42717,N_41545,N_41945);
xor U42718 (N_42718,N_41667,N_41713);
or U42719 (N_42719,N_41226,N_41216);
nor U42720 (N_42720,N_41823,N_41081);
xnor U42721 (N_42721,N_41563,N_41822);
and U42722 (N_42722,N_41269,N_41660);
nor U42723 (N_42723,N_41602,N_41226);
nand U42724 (N_42724,N_41556,N_41098);
nand U42725 (N_42725,N_41176,N_41338);
nor U42726 (N_42726,N_41632,N_41379);
or U42727 (N_42727,N_41847,N_41635);
nor U42728 (N_42728,N_41357,N_41939);
and U42729 (N_42729,N_41975,N_41341);
nand U42730 (N_42730,N_41562,N_41455);
and U42731 (N_42731,N_41109,N_41672);
nor U42732 (N_42732,N_41222,N_41121);
xor U42733 (N_42733,N_41949,N_41980);
or U42734 (N_42734,N_41969,N_41807);
nand U42735 (N_42735,N_41359,N_41428);
nor U42736 (N_42736,N_41461,N_41668);
or U42737 (N_42737,N_41077,N_41525);
and U42738 (N_42738,N_41720,N_41753);
or U42739 (N_42739,N_41586,N_41183);
xnor U42740 (N_42740,N_41127,N_41206);
nand U42741 (N_42741,N_41793,N_41537);
nand U42742 (N_42742,N_41122,N_41057);
xor U42743 (N_42743,N_41812,N_41765);
nor U42744 (N_42744,N_41663,N_41022);
xor U42745 (N_42745,N_41287,N_41305);
and U42746 (N_42746,N_41906,N_41484);
nand U42747 (N_42747,N_41894,N_41776);
and U42748 (N_42748,N_41830,N_41536);
and U42749 (N_42749,N_41332,N_41722);
and U42750 (N_42750,N_41434,N_41409);
nand U42751 (N_42751,N_41841,N_41274);
nand U42752 (N_42752,N_41221,N_41844);
nand U42753 (N_42753,N_41945,N_41095);
and U42754 (N_42754,N_41070,N_41150);
nor U42755 (N_42755,N_41835,N_41247);
nand U42756 (N_42756,N_41493,N_41878);
and U42757 (N_42757,N_41370,N_41629);
or U42758 (N_42758,N_41544,N_41188);
xor U42759 (N_42759,N_41589,N_41791);
nand U42760 (N_42760,N_41104,N_41328);
or U42761 (N_42761,N_41901,N_41783);
xnor U42762 (N_42762,N_41426,N_41515);
nand U42763 (N_42763,N_41809,N_41539);
nand U42764 (N_42764,N_41972,N_41317);
and U42765 (N_42765,N_41780,N_41892);
nand U42766 (N_42766,N_41511,N_41288);
and U42767 (N_42767,N_41889,N_41679);
xor U42768 (N_42768,N_41411,N_41780);
nand U42769 (N_42769,N_41239,N_41433);
and U42770 (N_42770,N_41866,N_41370);
and U42771 (N_42771,N_41840,N_41559);
xor U42772 (N_42772,N_41738,N_41065);
nand U42773 (N_42773,N_41236,N_41282);
xor U42774 (N_42774,N_41501,N_41121);
nor U42775 (N_42775,N_41837,N_41549);
nor U42776 (N_42776,N_41883,N_41167);
or U42777 (N_42777,N_41566,N_41200);
nand U42778 (N_42778,N_41923,N_41536);
or U42779 (N_42779,N_41859,N_41919);
nand U42780 (N_42780,N_41261,N_41138);
nand U42781 (N_42781,N_41662,N_41790);
xor U42782 (N_42782,N_41966,N_41691);
nand U42783 (N_42783,N_41198,N_41536);
and U42784 (N_42784,N_41351,N_41093);
or U42785 (N_42785,N_41561,N_41413);
xnor U42786 (N_42786,N_41245,N_41360);
or U42787 (N_42787,N_41720,N_41582);
or U42788 (N_42788,N_41985,N_41899);
nor U42789 (N_42789,N_41466,N_41401);
nor U42790 (N_42790,N_41390,N_41956);
or U42791 (N_42791,N_41729,N_41532);
xnor U42792 (N_42792,N_41675,N_41101);
xnor U42793 (N_42793,N_41427,N_41778);
xnor U42794 (N_42794,N_41299,N_41705);
xnor U42795 (N_42795,N_41046,N_41357);
xnor U42796 (N_42796,N_41776,N_41929);
nand U42797 (N_42797,N_41057,N_41663);
nor U42798 (N_42798,N_41542,N_41726);
and U42799 (N_42799,N_41669,N_41288);
nor U42800 (N_42800,N_41287,N_41740);
nor U42801 (N_42801,N_41663,N_41544);
xnor U42802 (N_42802,N_41568,N_41224);
and U42803 (N_42803,N_41906,N_41615);
nand U42804 (N_42804,N_41730,N_41980);
xor U42805 (N_42805,N_41109,N_41055);
and U42806 (N_42806,N_41866,N_41525);
or U42807 (N_42807,N_41707,N_41725);
or U42808 (N_42808,N_41943,N_41249);
xnor U42809 (N_42809,N_41537,N_41508);
nor U42810 (N_42810,N_41287,N_41683);
or U42811 (N_42811,N_41148,N_41033);
nand U42812 (N_42812,N_41750,N_41347);
and U42813 (N_42813,N_41774,N_41294);
or U42814 (N_42814,N_41305,N_41818);
and U42815 (N_42815,N_41026,N_41080);
or U42816 (N_42816,N_41453,N_41694);
xnor U42817 (N_42817,N_41934,N_41177);
nor U42818 (N_42818,N_41329,N_41420);
xor U42819 (N_42819,N_41610,N_41257);
nor U42820 (N_42820,N_41065,N_41591);
xnor U42821 (N_42821,N_41778,N_41857);
and U42822 (N_42822,N_41644,N_41871);
nand U42823 (N_42823,N_41054,N_41436);
and U42824 (N_42824,N_41254,N_41209);
nor U42825 (N_42825,N_41766,N_41312);
and U42826 (N_42826,N_41721,N_41922);
or U42827 (N_42827,N_41608,N_41697);
nand U42828 (N_42828,N_41900,N_41842);
nor U42829 (N_42829,N_41237,N_41784);
xnor U42830 (N_42830,N_41537,N_41122);
xor U42831 (N_42831,N_41428,N_41176);
and U42832 (N_42832,N_41561,N_41642);
xor U42833 (N_42833,N_41043,N_41973);
nand U42834 (N_42834,N_41159,N_41204);
or U42835 (N_42835,N_41188,N_41260);
or U42836 (N_42836,N_41341,N_41059);
xor U42837 (N_42837,N_41097,N_41580);
nor U42838 (N_42838,N_41595,N_41674);
nor U42839 (N_42839,N_41711,N_41696);
or U42840 (N_42840,N_41962,N_41010);
xor U42841 (N_42841,N_41852,N_41787);
or U42842 (N_42842,N_41828,N_41276);
nand U42843 (N_42843,N_41871,N_41334);
or U42844 (N_42844,N_41296,N_41511);
nor U42845 (N_42845,N_41068,N_41002);
nand U42846 (N_42846,N_41432,N_41329);
nand U42847 (N_42847,N_41264,N_41789);
and U42848 (N_42848,N_41274,N_41067);
xor U42849 (N_42849,N_41129,N_41734);
xnor U42850 (N_42850,N_41141,N_41689);
and U42851 (N_42851,N_41862,N_41979);
and U42852 (N_42852,N_41223,N_41496);
nor U42853 (N_42853,N_41597,N_41232);
xor U42854 (N_42854,N_41951,N_41376);
or U42855 (N_42855,N_41677,N_41722);
nor U42856 (N_42856,N_41477,N_41736);
and U42857 (N_42857,N_41796,N_41626);
xnor U42858 (N_42858,N_41438,N_41173);
nand U42859 (N_42859,N_41643,N_41648);
or U42860 (N_42860,N_41048,N_41698);
and U42861 (N_42861,N_41421,N_41834);
nand U42862 (N_42862,N_41943,N_41905);
nor U42863 (N_42863,N_41834,N_41278);
nand U42864 (N_42864,N_41849,N_41776);
nand U42865 (N_42865,N_41946,N_41640);
and U42866 (N_42866,N_41649,N_41619);
nand U42867 (N_42867,N_41494,N_41307);
nor U42868 (N_42868,N_41296,N_41411);
nand U42869 (N_42869,N_41900,N_41474);
and U42870 (N_42870,N_41036,N_41551);
nand U42871 (N_42871,N_41423,N_41417);
and U42872 (N_42872,N_41885,N_41937);
xor U42873 (N_42873,N_41168,N_41522);
and U42874 (N_42874,N_41375,N_41276);
and U42875 (N_42875,N_41381,N_41341);
xor U42876 (N_42876,N_41219,N_41903);
nand U42877 (N_42877,N_41097,N_41348);
and U42878 (N_42878,N_41606,N_41523);
xnor U42879 (N_42879,N_41734,N_41985);
or U42880 (N_42880,N_41803,N_41642);
and U42881 (N_42881,N_41647,N_41936);
xor U42882 (N_42882,N_41209,N_41173);
and U42883 (N_42883,N_41597,N_41661);
or U42884 (N_42884,N_41591,N_41533);
nand U42885 (N_42885,N_41686,N_41072);
nand U42886 (N_42886,N_41896,N_41190);
nor U42887 (N_42887,N_41813,N_41815);
and U42888 (N_42888,N_41172,N_41249);
nor U42889 (N_42889,N_41560,N_41470);
nor U42890 (N_42890,N_41887,N_41129);
xor U42891 (N_42891,N_41389,N_41369);
nand U42892 (N_42892,N_41638,N_41970);
nor U42893 (N_42893,N_41508,N_41190);
nand U42894 (N_42894,N_41545,N_41122);
xor U42895 (N_42895,N_41341,N_41447);
or U42896 (N_42896,N_41033,N_41337);
nand U42897 (N_42897,N_41239,N_41548);
nor U42898 (N_42898,N_41070,N_41889);
or U42899 (N_42899,N_41365,N_41374);
nand U42900 (N_42900,N_41528,N_41223);
nor U42901 (N_42901,N_41045,N_41489);
nor U42902 (N_42902,N_41386,N_41159);
nand U42903 (N_42903,N_41996,N_41877);
and U42904 (N_42904,N_41205,N_41551);
xor U42905 (N_42905,N_41682,N_41506);
or U42906 (N_42906,N_41118,N_41583);
xnor U42907 (N_42907,N_41722,N_41592);
nand U42908 (N_42908,N_41204,N_41510);
and U42909 (N_42909,N_41118,N_41098);
and U42910 (N_42910,N_41621,N_41903);
nand U42911 (N_42911,N_41246,N_41961);
nand U42912 (N_42912,N_41441,N_41789);
xnor U42913 (N_42913,N_41401,N_41226);
nor U42914 (N_42914,N_41865,N_41033);
nor U42915 (N_42915,N_41043,N_41241);
and U42916 (N_42916,N_41704,N_41553);
nor U42917 (N_42917,N_41094,N_41363);
nor U42918 (N_42918,N_41906,N_41201);
nand U42919 (N_42919,N_41180,N_41490);
or U42920 (N_42920,N_41192,N_41865);
or U42921 (N_42921,N_41766,N_41132);
nand U42922 (N_42922,N_41051,N_41031);
or U42923 (N_42923,N_41308,N_41902);
and U42924 (N_42924,N_41486,N_41644);
xnor U42925 (N_42925,N_41824,N_41264);
nor U42926 (N_42926,N_41002,N_41763);
xnor U42927 (N_42927,N_41016,N_41642);
xor U42928 (N_42928,N_41062,N_41759);
nor U42929 (N_42929,N_41742,N_41206);
nand U42930 (N_42930,N_41129,N_41946);
or U42931 (N_42931,N_41373,N_41016);
xor U42932 (N_42932,N_41441,N_41337);
nor U42933 (N_42933,N_41281,N_41606);
nand U42934 (N_42934,N_41483,N_41492);
xnor U42935 (N_42935,N_41239,N_41739);
and U42936 (N_42936,N_41760,N_41914);
or U42937 (N_42937,N_41401,N_41214);
xnor U42938 (N_42938,N_41613,N_41063);
xor U42939 (N_42939,N_41844,N_41383);
or U42940 (N_42940,N_41407,N_41919);
nor U42941 (N_42941,N_41057,N_41799);
nand U42942 (N_42942,N_41749,N_41648);
or U42943 (N_42943,N_41860,N_41455);
nor U42944 (N_42944,N_41168,N_41396);
and U42945 (N_42945,N_41781,N_41251);
or U42946 (N_42946,N_41068,N_41033);
and U42947 (N_42947,N_41125,N_41593);
or U42948 (N_42948,N_41513,N_41128);
xnor U42949 (N_42949,N_41354,N_41259);
and U42950 (N_42950,N_41170,N_41083);
or U42951 (N_42951,N_41193,N_41777);
xnor U42952 (N_42952,N_41219,N_41951);
xor U42953 (N_42953,N_41153,N_41363);
and U42954 (N_42954,N_41857,N_41402);
nor U42955 (N_42955,N_41789,N_41101);
xnor U42956 (N_42956,N_41568,N_41190);
or U42957 (N_42957,N_41471,N_41300);
and U42958 (N_42958,N_41234,N_41585);
xor U42959 (N_42959,N_41401,N_41074);
and U42960 (N_42960,N_41071,N_41715);
and U42961 (N_42961,N_41511,N_41044);
or U42962 (N_42962,N_41615,N_41840);
nand U42963 (N_42963,N_41773,N_41591);
nand U42964 (N_42964,N_41683,N_41185);
xnor U42965 (N_42965,N_41079,N_41107);
nand U42966 (N_42966,N_41193,N_41527);
nand U42967 (N_42967,N_41742,N_41380);
or U42968 (N_42968,N_41969,N_41026);
or U42969 (N_42969,N_41632,N_41982);
and U42970 (N_42970,N_41131,N_41119);
nand U42971 (N_42971,N_41951,N_41717);
and U42972 (N_42972,N_41609,N_41921);
nor U42973 (N_42973,N_41696,N_41615);
and U42974 (N_42974,N_41146,N_41605);
and U42975 (N_42975,N_41227,N_41884);
or U42976 (N_42976,N_41854,N_41100);
nand U42977 (N_42977,N_41028,N_41541);
xnor U42978 (N_42978,N_41001,N_41435);
or U42979 (N_42979,N_41615,N_41441);
or U42980 (N_42980,N_41608,N_41337);
nor U42981 (N_42981,N_41796,N_41525);
and U42982 (N_42982,N_41167,N_41085);
nand U42983 (N_42983,N_41530,N_41305);
xor U42984 (N_42984,N_41525,N_41031);
or U42985 (N_42985,N_41586,N_41498);
and U42986 (N_42986,N_41662,N_41512);
or U42987 (N_42987,N_41888,N_41147);
xor U42988 (N_42988,N_41611,N_41568);
nand U42989 (N_42989,N_41153,N_41373);
xor U42990 (N_42990,N_41766,N_41749);
nand U42991 (N_42991,N_41527,N_41046);
xnor U42992 (N_42992,N_41560,N_41480);
nor U42993 (N_42993,N_41942,N_41638);
and U42994 (N_42994,N_41724,N_41576);
xor U42995 (N_42995,N_41929,N_41895);
nand U42996 (N_42996,N_41899,N_41219);
nand U42997 (N_42997,N_41760,N_41011);
nor U42998 (N_42998,N_41160,N_41163);
or U42999 (N_42999,N_41642,N_41865);
xnor U43000 (N_43000,N_42412,N_42347);
xor U43001 (N_43001,N_42780,N_42728);
and U43002 (N_43002,N_42127,N_42556);
and U43003 (N_43003,N_42094,N_42875);
or U43004 (N_43004,N_42241,N_42585);
xnor U43005 (N_43005,N_42679,N_42055);
nor U43006 (N_43006,N_42735,N_42515);
or U43007 (N_43007,N_42617,N_42719);
nor U43008 (N_43008,N_42032,N_42958);
nand U43009 (N_43009,N_42286,N_42653);
nand U43010 (N_43010,N_42114,N_42611);
and U43011 (N_43011,N_42501,N_42165);
and U43012 (N_43012,N_42090,N_42764);
nand U43013 (N_43013,N_42152,N_42861);
nand U43014 (N_43014,N_42065,N_42253);
xnor U43015 (N_43015,N_42524,N_42684);
or U43016 (N_43016,N_42011,N_42818);
nor U43017 (N_43017,N_42627,N_42411);
nor U43018 (N_43018,N_42647,N_42095);
nand U43019 (N_43019,N_42405,N_42690);
or U43020 (N_43020,N_42419,N_42354);
and U43021 (N_43021,N_42193,N_42900);
or U43022 (N_43022,N_42837,N_42722);
xor U43023 (N_43023,N_42358,N_42705);
and U43024 (N_43024,N_42079,N_42991);
and U43025 (N_43025,N_42004,N_42480);
nand U43026 (N_43026,N_42484,N_42163);
nand U43027 (N_43027,N_42208,N_42450);
or U43028 (N_43028,N_42022,N_42709);
nand U43029 (N_43029,N_42268,N_42896);
or U43030 (N_43030,N_42188,N_42021);
nor U43031 (N_43031,N_42260,N_42276);
nand U43032 (N_43032,N_42579,N_42797);
nor U43033 (N_43033,N_42031,N_42905);
xor U43034 (N_43034,N_42969,N_42911);
nor U43035 (N_43035,N_42944,N_42568);
or U43036 (N_43036,N_42409,N_42945);
and U43037 (N_43037,N_42870,N_42441);
xnor U43038 (N_43038,N_42695,N_42227);
or U43039 (N_43039,N_42202,N_42319);
nand U43040 (N_43040,N_42345,N_42996);
xor U43041 (N_43041,N_42424,N_42586);
nand U43042 (N_43042,N_42015,N_42646);
xnor U43043 (N_43043,N_42348,N_42103);
and U43044 (N_43044,N_42306,N_42746);
and U43045 (N_43045,N_42481,N_42661);
nor U43046 (N_43046,N_42597,N_42561);
nor U43047 (N_43047,N_42659,N_42619);
nand U43048 (N_43048,N_42217,N_42964);
xor U43049 (N_43049,N_42939,N_42576);
and U43050 (N_43050,N_42249,N_42003);
or U43051 (N_43051,N_42883,N_42080);
nor U43052 (N_43052,N_42739,N_42804);
xor U43053 (N_43053,N_42102,N_42057);
and U43054 (N_43054,N_42670,N_42063);
or U43055 (N_43055,N_42731,N_42935);
nand U43056 (N_43056,N_42398,N_42142);
nand U43057 (N_43057,N_42242,N_42457);
nor U43058 (N_43058,N_42064,N_42546);
xor U43059 (N_43059,N_42821,N_42040);
nand U43060 (N_43060,N_42018,N_42651);
nor U43061 (N_43061,N_42461,N_42074);
xnor U43062 (N_43062,N_42421,N_42187);
and U43063 (N_43063,N_42541,N_42186);
and U43064 (N_43064,N_42706,N_42362);
and U43065 (N_43065,N_42360,N_42342);
or U43066 (N_43066,N_42938,N_42898);
and U43067 (N_43067,N_42971,N_42236);
and U43068 (N_43068,N_42060,N_42869);
or U43069 (N_43069,N_42698,N_42234);
and U43070 (N_43070,N_42558,N_42762);
and U43071 (N_43071,N_42331,N_42582);
or U43072 (N_43072,N_42263,N_42274);
xnor U43073 (N_43073,N_42367,N_42917);
and U43074 (N_43074,N_42547,N_42321);
and U43075 (N_43075,N_42085,N_42049);
nor U43076 (N_43076,N_42271,N_42552);
nor U43077 (N_43077,N_42554,N_42959);
nor U43078 (N_43078,N_42589,N_42785);
nand U43079 (N_43079,N_42769,N_42406);
and U43080 (N_43080,N_42766,N_42191);
or U43081 (N_43081,N_42140,N_42575);
nand U43082 (N_43082,N_42963,N_42178);
and U43083 (N_43083,N_42696,N_42282);
xor U43084 (N_43084,N_42951,N_42291);
xor U43085 (N_43085,N_42867,N_42046);
nand U43086 (N_43086,N_42506,N_42244);
or U43087 (N_43087,N_42609,N_42929);
nor U43088 (N_43088,N_42516,N_42431);
or U43089 (N_43089,N_42363,N_42304);
or U43090 (N_43090,N_42510,N_42239);
xor U43091 (N_43091,N_42596,N_42614);
xor U43092 (N_43092,N_42717,N_42564);
nor U43093 (N_43093,N_42344,N_42529);
nand U43094 (N_43094,N_42000,N_42933);
nor U43095 (N_43095,N_42810,N_42452);
or U43096 (N_43096,N_42654,N_42125);
nor U43097 (N_43097,N_42136,N_42738);
nand U43098 (N_43098,N_42451,N_42711);
nor U43099 (N_43099,N_42396,N_42350);
or U43100 (N_43100,N_42429,N_42872);
and U43101 (N_43101,N_42976,N_42774);
and U43102 (N_43102,N_42625,N_42508);
xnor U43103 (N_43103,N_42068,N_42028);
nor U43104 (N_43104,N_42594,N_42427);
nand U43105 (N_43105,N_42889,N_42744);
nor U43106 (N_43106,N_42885,N_42414);
or U43107 (N_43107,N_42311,N_42496);
and U43108 (N_43108,N_42098,N_42300);
xor U43109 (N_43109,N_42866,N_42838);
and U43110 (N_43110,N_42394,N_42841);
and U43111 (N_43111,N_42397,N_42981);
xnor U43112 (N_43112,N_42482,N_42091);
nor U43113 (N_43113,N_42144,N_42305);
or U43114 (N_43114,N_42848,N_42814);
nand U43115 (N_43115,N_42148,N_42726);
nor U43116 (N_43116,N_42381,N_42952);
or U43117 (N_43117,N_42308,N_42834);
and U43118 (N_43118,N_42824,N_42608);
xnor U43119 (N_43119,N_42833,N_42827);
and U43120 (N_43120,N_42954,N_42198);
nor U43121 (N_43121,N_42519,N_42968);
xor U43122 (N_43122,N_42873,N_42538);
xnor U43123 (N_43123,N_42544,N_42469);
and U43124 (N_43124,N_42732,N_42030);
nor U43125 (N_43125,N_42047,N_42357);
and U43126 (N_43126,N_42113,N_42270);
nor U43127 (N_43127,N_42649,N_42545);
or U43128 (N_43128,N_42323,N_42328);
nor U43129 (N_43129,N_42395,N_42806);
and U43130 (N_43130,N_42920,N_42168);
nor U43131 (N_43131,N_42007,N_42631);
and U43132 (N_43132,N_42967,N_42225);
or U43133 (N_43133,N_42216,N_42026);
xnor U43134 (N_43134,N_42602,N_42509);
nor U43135 (N_43135,N_42598,N_42855);
and U43136 (N_43136,N_42630,N_42283);
nand U43137 (N_43137,N_42449,N_42555);
and U43138 (N_43138,N_42111,N_42039);
nor U43139 (N_43139,N_42259,N_42445);
xor U43140 (N_43140,N_42928,N_42024);
or U43141 (N_43141,N_42658,N_42009);
and U43142 (N_43142,N_42822,N_42708);
nor U43143 (N_43143,N_42408,N_42389);
nor U43144 (N_43144,N_42418,N_42563);
nand U43145 (N_43145,N_42237,N_42688);
xnor U43146 (N_43146,N_42641,N_42560);
nand U43147 (N_43147,N_42874,N_42448);
or U43148 (N_43148,N_42084,N_42226);
xor U43149 (N_43149,N_42666,N_42209);
or U43150 (N_43150,N_42580,N_42668);
nand U43151 (N_43151,N_42423,N_42703);
or U43152 (N_43152,N_42845,N_42511);
or U43153 (N_43153,N_42212,N_42017);
and U43154 (N_43154,N_42200,N_42776);
nor U43155 (N_43155,N_42789,N_42203);
xnor U43156 (N_43156,N_42061,N_42836);
nor U43157 (N_43157,N_42486,N_42010);
xor U43158 (N_43158,N_42373,N_42131);
xor U43159 (N_43159,N_42779,N_42685);
or U43160 (N_43160,N_42376,N_42336);
xor U43161 (N_43161,N_42196,N_42638);
nor U43162 (N_43162,N_42391,N_42995);
nand U43163 (N_43163,N_42553,N_42264);
or U43164 (N_43164,N_42218,N_42067);
xor U43165 (N_43165,N_42077,N_42669);
and U43166 (N_43166,N_42223,N_42603);
xnor U43167 (N_43167,N_42158,N_42904);
nand U43168 (N_43168,N_42923,N_42134);
xor U43169 (N_43169,N_42941,N_42574);
nand U43170 (N_43170,N_42890,N_42346);
and U43171 (N_43171,N_42133,N_42924);
nor U43172 (N_43172,N_42862,N_42371);
and U43173 (N_43173,N_42364,N_42536);
xnor U43174 (N_43174,N_42686,N_42674);
and U43175 (N_43175,N_42856,N_42813);
and U43176 (N_43176,N_42124,N_42587);
nor U43177 (N_43177,N_42689,N_42310);
and U43178 (N_43178,N_42466,N_42499);
or U43179 (N_43179,N_42707,N_42416);
and U43180 (N_43180,N_42853,N_42730);
or U43181 (N_43181,N_42915,N_42712);
nor U43182 (N_43182,N_42453,N_42372);
xnor U43183 (N_43183,N_42167,N_42878);
or U43184 (N_43184,N_42784,N_42830);
nor U43185 (N_43185,N_42792,N_42369);
nor U43186 (N_43186,N_42219,N_42143);
xnor U43187 (N_43187,N_42807,N_42037);
and U43188 (N_43188,N_42301,N_42072);
and U43189 (N_43189,N_42128,N_42577);
xor U43190 (N_43190,N_42736,N_42288);
nand U43191 (N_43191,N_42337,N_42643);
or U43192 (N_43192,N_42020,N_42543);
nor U43193 (N_43193,N_42044,N_42432);
nand U43194 (N_43194,N_42153,N_42392);
xnor U43195 (N_43195,N_42338,N_42622);
and U43196 (N_43196,N_42897,N_42341);
nand U43197 (N_43197,N_42989,N_42982);
nor U43198 (N_43198,N_42206,N_42156);
xnor U43199 (N_43199,N_42335,N_42333);
xor U43200 (N_43200,N_42663,N_42793);
xnor U43201 (N_43201,N_42737,N_42317);
or U43202 (N_43202,N_42812,N_42468);
xor U43203 (N_43203,N_42652,N_42704);
nor U43204 (N_43204,N_42994,N_42116);
xor U43205 (N_43205,N_42718,N_42520);
xor U43206 (N_43206,N_42887,N_42471);
nand U43207 (N_43207,N_42492,N_42682);
or U43208 (N_43208,N_42475,N_42681);
nand U43209 (N_43209,N_42906,N_42016);
and U43210 (N_43210,N_42045,N_42680);
xor U43211 (N_43211,N_42247,N_42697);
xor U43212 (N_43212,N_42566,N_42087);
nand U43213 (N_43213,N_42415,N_42041);
nand U43214 (N_43214,N_42595,N_42801);
and U43215 (N_43215,N_42059,N_42303);
nor U43216 (N_43216,N_42176,N_42562);
and U43217 (N_43217,N_42727,N_42368);
xor U43218 (N_43218,N_42527,N_42166);
nor U43219 (N_43219,N_42925,N_42962);
nor U43220 (N_43220,N_42284,N_42811);
nor U43221 (N_43221,N_42246,N_42447);
nor U43222 (N_43222,N_42851,N_42375);
and U43223 (N_43223,N_42184,N_42699);
nand U43224 (N_43224,N_42950,N_42639);
xnor U43225 (N_43225,N_42593,N_42361);
and U43226 (N_43226,N_42002,N_42177);
nand U43227 (N_43227,N_42235,N_42076);
xnor U43228 (N_43228,N_42477,N_42840);
and U43229 (N_43229,N_42642,N_42458);
nor U43230 (N_43230,N_42472,N_42075);
xor U43231 (N_43231,N_42295,N_42353);
nor U43232 (N_43232,N_42694,N_42782);
and U43233 (N_43233,N_42488,N_42565);
nor U43234 (N_43234,N_42921,N_42023);
nor U43235 (N_43235,N_42693,N_42384);
and U43236 (N_43236,N_42997,N_42135);
or U43237 (N_43237,N_42370,N_42755);
or U43238 (N_43238,N_42279,N_42465);
nand U43239 (N_43239,N_42388,N_42828);
nand U43240 (N_43240,N_42894,N_42729);
or U43241 (N_43241,N_42112,N_42473);
or U43242 (N_43242,N_42985,N_42220);
or U43243 (N_43243,N_42498,N_42322);
nand U43244 (N_43244,N_42352,N_42528);
nor U43245 (N_43245,N_42359,N_42761);
and U43246 (N_43246,N_42132,N_42294);
nand U43247 (N_43247,N_42355,N_42474);
nor U43248 (N_43248,N_42001,N_42459);
and U43249 (N_43249,N_42145,N_42365);
or U43250 (N_43250,N_42932,N_42919);
and U43251 (N_43251,N_42960,N_42926);
or U43252 (N_43252,N_42988,N_42417);
or U43253 (N_43253,N_42146,N_42559);
and U43254 (N_43254,N_42808,N_42185);
xnor U43255 (N_43255,N_42990,N_42050);
nand U43256 (N_43256,N_42129,N_42460);
nor U43257 (N_43257,N_42918,N_42390);
nor U43258 (N_43258,N_42831,N_42507);
and U43259 (N_43259,N_42787,N_42588);
xor U43260 (N_43260,N_42826,N_42318);
xor U43261 (N_43261,N_42036,N_42772);
nand U43262 (N_43262,N_42986,N_42750);
nor U43263 (N_43263,N_42182,N_42604);
nand U43264 (N_43264,N_42307,N_42850);
nor U43265 (N_43265,N_42343,N_42623);
nand U43266 (N_43266,N_42118,N_42179);
nor U43267 (N_43267,N_42993,N_42590);
xnor U43268 (N_43268,N_42854,N_42832);
nor U43269 (N_43269,N_42446,N_42891);
nor U43270 (N_43270,N_42635,N_42181);
or U43271 (N_43271,N_42513,N_42281);
xnor U43272 (N_43272,N_42108,N_42914);
and U43273 (N_43273,N_42999,N_42083);
nand U43274 (N_43274,N_42800,N_42266);
nor U43275 (N_43275,N_42846,N_42073);
xnor U43276 (N_43276,N_42115,N_42734);
xnor U43277 (N_43277,N_42403,N_42671);
nor U43278 (N_43278,N_42913,N_42640);
nor U43279 (N_43279,N_42410,N_42799);
nor U43280 (N_43280,N_42664,N_42314);
xor U43281 (N_43281,N_42716,N_42940);
nand U43282 (N_43282,N_42204,N_42215);
nand U43283 (N_43283,N_42296,N_42387);
nand U43284 (N_43284,N_42299,N_42700);
nor U43285 (N_43285,N_42329,N_42916);
and U43286 (N_43286,N_42230,N_42183);
nand U43287 (N_43287,N_42297,N_42042);
and U43288 (N_43288,N_42942,N_42549);
nand U43289 (N_43289,N_42667,N_42790);
or U43290 (N_43290,N_42277,N_42164);
xor U43291 (N_43291,N_42616,N_42105);
or U43292 (N_43292,N_42422,N_42823);
nand U43293 (N_43293,N_42927,N_42530);
or U43294 (N_43294,N_42953,N_42006);
and U43295 (N_43295,N_42526,N_42197);
and U43296 (N_43296,N_42213,N_42287);
nand U43297 (N_43297,N_42765,N_42535);
nor U43298 (N_43298,N_42442,N_42691);
nor U43299 (N_43299,N_42678,N_42816);
nand U43300 (N_43300,N_42443,N_42171);
nand U43301 (N_43301,N_42402,N_42798);
xor U43302 (N_43302,N_42882,N_42683);
or U43303 (N_43303,N_42992,N_42910);
and U43304 (N_43304,N_42612,N_42272);
and U43305 (N_43305,N_42089,N_42071);
nor U43306 (N_43306,N_42819,N_42238);
and U43307 (N_43307,N_42521,N_42313);
nand U43308 (N_43308,N_42636,N_42749);
or U43309 (N_43309,N_42435,N_42839);
and U43310 (N_43310,N_42551,N_42759);
xnor U43311 (N_43311,N_42008,N_42880);
or U43312 (N_43312,N_42934,N_42650);
or U43313 (N_43313,N_42503,N_42302);
xnor U43314 (N_43314,N_42487,N_42634);
or U43315 (N_43315,N_42504,N_42339);
nor U43316 (N_43316,N_42676,N_42835);
nand U43317 (N_43317,N_42907,N_42485);
or U43318 (N_43318,N_42280,N_42753);
and U43319 (N_43319,N_42325,N_42326);
nor U43320 (N_43320,N_42518,N_42232);
xor U43321 (N_43321,N_42251,N_42380);
or U43322 (N_43322,N_42123,N_42657);
xor U43323 (N_43323,N_42805,N_42413);
nor U43324 (N_43324,N_42931,N_42748);
nand U43325 (N_43325,N_42970,N_42399);
nor U43326 (N_43326,N_42285,N_42626);
nor U43327 (N_43327,N_42881,N_42600);
xor U43328 (N_43328,N_42456,N_42298);
nand U43329 (N_43329,N_42138,N_42721);
nand U43330 (N_43330,N_42628,N_42888);
xor U43331 (N_43331,N_42201,N_42386);
nor U43332 (N_43332,N_42438,N_42439);
xor U43333 (N_43333,N_42385,N_42902);
xnor U43334 (N_43334,N_42444,N_42591);
nor U43335 (N_43335,N_42351,N_42137);
or U43336 (N_43336,N_42523,N_42803);
xor U43337 (N_43337,N_42497,N_42194);
or U43338 (N_43338,N_42309,N_42884);
nand U43339 (N_43339,N_42871,N_42278);
xor U43340 (N_43340,N_42713,N_42930);
and U43341 (N_43341,N_42231,N_42005);
nand U43342 (N_43342,N_42978,N_42240);
or U43343 (N_43343,N_42532,N_42093);
or U43344 (N_43344,N_42760,N_42618);
nand U43345 (N_43345,N_42768,N_42578);
nor U43346 (N_43346,N_42425,N_42956);
and U43347 (N_43347,N_42829,N_42788);
nor U43348 (N_43348,N_42715,N_42817);
or U43349 (N_43349,N_42211,N_42615);
or U43350 (N_43350,N_42100,N_42710);
xnor U43351 (N_43351,N_42292,N_42975);
and U43352 (N_43352,N_42864,N_42190);
xnor U43353 (N_43353,N_42781,N_42228);
nand U43354 (N_43354,N_42273,N_42092);
nand U43355 (N_43355,N_42675,N_42013);
nor U43356 (N_43356,N_42665,N_42983);
and U43357 (N_43357,N_42379,N_42437);
nor U43358 (N_43358,N_42229,N_42633);
nand U43359 (N_43359,N_42464,N_42078);
nor U43360 (N_43360,N_42195,N_42033);
nor U43361 (N_43361,N_42054,N_42791);
or U43362 (N_43362,N_42058,N_42052);
or U43363 (N_43363,N_42248,N_42533);
xnor U43364 (N_43364,N_42027,N_42895);
and U43365 (N_43365,N_42644,N_42802);
xnor U43366 (N_43366,N_42154,N_42783);
or U43367 (N_43367,N_42767,N_42624);
nand U43368 (N_43368,N_42210,N_42147);
and U43369 (N_43369,N_42025,N_42070);
nand U43370 (N_43370,N_42757,N_42893);
nor U43371 (N_43371,N_42778,N_42069);
nor U43372 (N_43372,N_42860,N_42955);
or U43373 (N_43373,N_42610,N_42479);
or U43374 (N_43374,N_42815,N_42943);
nor U43375 (N_43375,N_42972,N_42601);
or U43376 (N_43376,N_42572,N_42170);
and U43377 (N_43377,N_42099,N_42692);
xor U43378 (N_43378,N_42843,N_42275);
nand U43379 (N_43379,N_42998,N_42502);
xor U43380 (N_43380,N_42428,N_42569);
or U43381 (N_43381,N_42677,N_42672);
and U43382 (N_43382,N_42901,N_42687);
xor U43383 (N_43383,N_42775,N_42632);
nor U43384 (N_43384,N_42965,N_42258);
nand U43385 (N_43385,N_42120,N_42723);
xor U43386 (N_43386,N_42557,N_42796);
nand U43387 (N_43387,N_42426,N_42908);
nand U43388 (N_43388,N_42517,N_42648);
xnor U43389 (N_43389,N_42374,N_42849);
or U43390 (N_43390,N_42320,N_42974);
xor U43391 (N_43391,N_42117,N_42293);
or U43392 (N_43392,N_42493,N_42570);
and U43393 (N_43393,N_42289,N_42122);
and U43394 (N_43394,N_42483,N_42786);
nor U43395 (N_43395,N_42756,N_42868);
xnor U43396 (N_43396,N_42262,N_42899);
or U43397 (N_43397,N_42062,N_42673);
nand U43398 (N_43398,N_42495,N_42106);
xor U43399 (N_43399,N_42420,N_42257);
and U43400 (N_43400,N_42514,N_42252);
or U43401 (N_43401,N_42101,N_42973);
and U43402 (N_43402,N_42629,N_42316);
xnor U43403 (N_43403,N_42876,N_42733);
or U43404 (N_43404,N_42107,N_42470);
nand U43405 (N_43405,N_42491,N_42548);
and U43406 (N_43406,N_42404,N_42909);
nand U43407 (N_43407,N_42221,N_42531);
or U43408 (N_43408,N_42947,N_42014);
and U43409 (N_43409,N_42795,N_42606);
or U43410 (N_43410,N_42637,N_42349);
or U43411 (N_43411,N_42327,N_42957);
or U43412 (N_43412,N_42332,N_42583);
nand U43413 (N_43413,N_42747,N_42500);
xor U43414 (N_43414,N_42189,N_42987);
or U43415 (N_43415,N_42751,N_42243);
or U43416 (N_43416,N_42607,N_42490);
nand U43417 (N_43417,N_42400,N_42537);
or U43418 (N_43418,N_42740,N_42984);
nor U43419 (N_43419,N_42567,N_42852);
or U43420 (N_43420,N_42222,N_42139);
xor U43421 (N_43421,N_42773,N_42038);
and U43422 (N_43422,N_42255,N_42467);
nor U43423 (N_43423,N_42174,N_42662);
nor U43424 (N_43424,N_42724,N_42150);
and U43425 (N_43425,N_42126,N_42771);
nor U43426 (N_43426,N_42043,N_42645);
or U43427 (N_43427,N_42540,N_42130);
nor U43428 (N_43428,N_42454,N_42613);
xnor U43429 (N_43429,N_42088,N_42478);
nand U43430 (N_43430,N_42082,N_42119);
xnor U43431 (N_43431,N_42254,N_42573);
or U43432 (N_43432,N_42401,N_42159);
nor U43433 (N_43433,N_42892,N_42290);
nor U43434 (N_43434,N_42173,N_42382);
or U43435 (N_43435,N_42324,N_42256);
and U43436 (N_43436,N_42584,N_42366);
xnor U43437 (N_43437,N_42315,N_42720);
xor U43438 (N_43438,N_42051,N_42175);
or U43439 (N_43439,N_42199,N_42539);
nor U43440 (N_43440,N_42110,N_42525);
and U43441 (N_43441,N_42157,N_42269);
or U43442 (N_43442,N_42702,N_42462);
xor U43443 (N_43443,N_42592,N_42656);
or U43444 (N_43444,N_42961,N_42312);
or U43445 (N_43445,N_42621,N_42489);
and U43446 (N_43446,N_42056,N_42109);
or U43447 (N_43447,N_42233,N_42741);
xor U43448 (N_43448,N_42250,N_42035);
nand U43449 (N_43449,N_42777,N_42754);
nand U43450 (N_43450,N_42267,N_42378);
and U43451 (N_43451,N_42393,N_42012);
xor U43452 (N_43452,N_42214,N_42752);
xor U43453 (N_43453,N_42066,N_42192);
or U43454 (N_43454,N_42407,N_42980);
nor U43455 (N_43455,N_42340,N_42053);
or U43456 (N_43456,N_42794,N_42161);
nor U43457 (N_43457,N_42104,N_42966);
and U43458 (N_43458,N_42436,N_42261);
xnor U43459 (N_43459,N_42440,N_42505);
nand U43460 (N_43460,N_42151,N_42714);
nand U43461 (N_43461,N_42863,N_42857);
and U43462 (N_43462,N_42745,N_42912);
or U43463 (N_43463,N_42330,N_42937);
or U43464 (N_43464,N_42701,N_42356);
nor U43465 (N_43465,N_42180,N_42476);
xor U43466 (N_43466,N_42770,N_42434);
xor U43467 (N_43467,N_42809,N_42494);
and U43468 (N_43468,N_42847,N_42149);
xnor U43469 (N_43469,N_42743,N_42463);
or U43470 (N_43470,N_42865,N_42946);
xor U43471 (N_43471,N_42245,N_42820);
and U43472 (N_43472,N_42169,N_42948);
and U43473 (N_43473,N_42534,N_42844);
and U43474 (N_43474,N_42581,N_42034);
or U43475 (N_43475,N_42842,N_42858);
or U43476 (N_43476,N_42725,N_42086);
nor U43477 (N_43477,N_42430,N_42605);
nor U43478 (N_43478,N_42879,N_42433);
nor U43479 (N_43479,N_42825,N_42141);
and U43480 (N_43480,N_42949,N_42859);
nor U43481 (N_43481,N_42903,N_42265);
nand U43482 (N_43482,N_42224,N_42571);
xnor U43483 (N_43483,N_42096,N_42979);
and U43484 (N_43484,N_42742,N_42936);
and U43485 (N_43485,N_42048,N_42019);
nor U43486 (N_43486,N_42886,N_42121);
and U43487 (N_43487,N_42550,N_42160);
xnor U43488 (N_43488,N_42877,N_42207);
nor U43489 (N_43489,N_42512,N_42763);
nor U43490 (N_43490,N_42620,N_42655);
or U43491 (N_43491,N_42081,N_42455);
or U43492 (N_43492,N_42097,N_42377);
xor U43493 (N_43493,N_42383,N_42977);
xnor U43494 (N_43494,N_42155,N_42162);
xnor U43495 (N_43495,N_42599,N_42922);
nor U43496 (N_43496,N_42029,N_42172);
nor U43497 (N_43497,N_42334,N_42660);
or U43498 (N_43498,N_42542,N_42758);
or U43499 (N_43499,N_42522,N_42205);
xnor U43500 (N_43500,N_42833,N_42337);
or U43501 (N_43501,N_42410,N_42797);
or U43502 (N_43502,N_42530,N_42994);
nand U43503 (N_43503,N_42822,N_42578);
xnor U43504 (N_43504,N_42910,N_42661);
and U43505 (N_43505,N_42971,N_42736);
or U43506 (N_43506,N_42504,N_42311);
nand U43507 (N_43507,N_42346,N_42817);
nor U43508 (N_43508,N_42185,N_42129);
and U43509 (N_43509,N_42610,N_42766);
and U43510 (N_43510,N_42050,N_42152);
and U43511 (N_43511,N_42544,N_42004);
and U43512 (N_43512,N_42085,N_42589);
or U43513 (N_43513,N_42446,N_42921);
nor U43514 (N_43514,N_42504,N_42158);
nand U43515 (N_43515,N_42730,N_42841);
nand U43516 (N_43516,N_42234,N_42335);
nand U43517 (N_43517,N_42291,N_42379);
and U43518 (N_43518,N_42070,N_42671);
xor U43519 (N_43519,N_42598,N_42488);
or U43520 (N_43520,N_42107,N_42166);
or U43521 (N_43521,N_42196,N_42081);
nand U43522 (N_43522,N_42832,N_42615);
nand U43523 (N_43523,N_42840,N_42364);
nand U43524 (N_43524,N_42873,N_42879);
xor U43525 (N_43525,N_42903,N_42668);
xnor U43526 (N_43526,N_42219,N_42318);
xnor U43527 (N_43527,N_42532,N_42086);
or U43528 (N_43528,N_42664,N_42401);
or U43529 (N_43529,N_42081,N_42143);
nor U43530 (N_43530,N_42579,N_42445);
nand U43531 (N_43531,N_42079,N_42546);
and U43532 (N_43532,N_42167,N_42115);
xnor U43533 (N_43533,N_42327,N_42014);
xor U43534 (N_43534,N_42745,N_42169);
nand U43535 (N_43535,N_42775,N_42148);
or U43536 (N_43536,N_42828,N_42953);
xor U43537 (N_43537,N_42278,N_42792);
xor U43538 (N_43538,N_42597,N_42773);
and U43539 (N_43539,N_42021,N_42757);
xnor U43540 (N_43540,N_42522,N_42800);
nor U43541 (N_43541,N_42328,N_42008);
nand U43542 (N_43542,N_42848,N_42279);
or U43543 (N_43543,N_42083,N_42733);
and U43544 (N_43544,N_42473,N_42239);
xor U43545 (N_43545,N_42227,N_42263);
and U43546 (N_43546,N_42475,N_42693);
or U43547 (N_43547,N_42572,N_42946);
and U43548 (N_43548,N_42189,N_42683);
or U43549 (N_43549,N_42824,N_42152);
nor U43550 (N_43550,N_42757,N_42124);
nor U43551 (N_43551,N_42942,N_42459);
nor U43552 (N_43552,N_42204,N_42338);
or U43553 (N_43553,N_42189,N_42156);
nor U43554 (N_43554,N_42591,N_42820);
or U43555 (N_43555,N_42689,N_42203);
nand U43556 (N_43556,N_42004,N_42333);
xnor U43557 (N_43557,N_42894,N_42025);
and U43558 (N_43558,N_42031,N_42882);
or U43559 (N_43559,N_42525,N_42935);
xor U43560 (N_43560,N_42988,N_42460);
and U43561 (N_43561,N_42951,N_42906);
and U43562 (N_43562,N_42165,N_42950);
xnor U43563 (N_43563,N_42977,N_42870);
nor U43564 (N_43564,N_42804,N_42351);
xnor U43565 (N_43565,N_42817,N_42585);
or U43566 (N_43566,N_42404,N_42668);
nor U43567 (N_43567,N_42596,N_42096);
nor U43568 (N_43568,N_42051,N_42661);
nor U43569 (N_43569,N_42700,N_42050);
xnor U43570 (N_43570,N_42059,N_42080);
or U43571 (N_43571,N_42548,N_42946);
nor U43572 (N_43572,N_42853,N_42963);
nand U43573 (N_43573,N_42968,N_42125);
nand U43574 (N_43574,N_42878,N_42335);
and U43575 (N_43575,N_42957,N_42291);
xnor U43576 (N_43576,N_42858,N_42885);
nor U43577 (N_43577,N_42194,N_42238);
and U43578 (N_43578,N_42671,N_42392);
nand U43579 (N_43579,N_42215,N_42075);
nand U43580 (N_43580,N_42038,N_42586);
or U43581 (N_43581,N_42297,N_42951);
nor U43582 (N_43582,N_42625,N_42991);
or U43583 (N_43583,N_42735,N_42873);
nor U43584 (N_43584,N_42318,N_42882);
nor U43585 (N_43585,N_42896,N_42412);
and U43586 (N_43586,N_42615,N_42755);
nand U43587 (N_43587,N_42073,N_42286);
and U43588 (N_43588,N_42026,N_42608);
nand U43589 (N_43589,N_42866,N_42467);
xor U43590 (N_43590,N_42584,N_42281);
and U43591 (N_43591,N_42073,N_42769);
nand U43592 (N_43592,N_42926,N_42794);
xor U43593 (N_43593,N_42145,N_42783);
nor U43594 (N_43594,N_42589,N_42172);
or U43595 (N_43595,N_42588,N_42408);
and U43596 (N_43596,N_42440,N_42642);
or U43597 (N_43597,N_42481,N_42124);
nor U43598 (N_43598,N_42465,N_42542);
xor U43599 (N_43599,N_42743,N_42897);
or U43600 (N_43600,N_42441,N_42580);
and U43601 (N_43601,N_42577,N_42828);
nor U43602 (N_43602,N_42099,N_42416);
or U43603 (N_43603,N_42272,N_42583);
nand U43604 (N_43604,N_42192,N_42146);
and U43605 (N_43605,N_42911,N_42625);
and U43606 (N_43606,N_42090,N_42036);
nor U43607 (N_43607,N_42682,N_42463);
and U43608 (N_43608,N_42298,N_42123);
and U43609 (N_43609,N_42087,N_42260);
xor U43610 (N_43610,N_42915,N_42475);
or U43611 (N_43611,N_42953,N_42726);
or U43612 (N_43612,N_42801,N_42941);
or U43613 (N_43613,N_42978,N_42892);
nand U43614 (N_43614,N_42115,N_42768);
and U43615 (N_43615,N_42991,N_42758);
nor U43616 (N_43616,N_42280,N_42251);
xnor U43617 (N_43617,N_42375,N_42283);
xor U43618 (N_43618,N_42234,N_42896);
or U43619 (N_43619,N_42576,N_42589);
and U43620 (N_43620,N_42092,N_42636);
or U43621 (N_43621,N_42616,N_42347);
and U43622 (N_43622,N_42147,N_42485);
nand U43623 (N_43623,N_42006,N_42303);
nor U43624 (N_43624,N_42256,N_42133);
xor U43625 (N_43625,N_42113,N_42248);
or U43626 (N_43626,N_42671,N_42348);
and U43627 (N_43627,N_42066,N_42402);
or U43628 (N_43628,N_42284,N_42456);
nand U43629 (N_43629,N_42865,N_42025);
nor U43630 (N_43630,N_42828,N_42076);
nor U43631 (N_43631,N_42444,N_42391);
and U43632 (N_43632,N_42601,N_42514);
or U43633 (N_43633,N_42487,N_42850);
nor U43634 (N_43634,N_42427,N_42588);
nor U43635 (N_43635,N_42904,N_42850);
and U43636 (N_43636,N_42801,N_42686);
nor U43637 (N_43637,N_42963,N_42347);
nand U43638 (N_43638,N_42657,N_42576);
or U43639 (N_43639,N_42054,N_42988);
xnor U43640 (N_43640,N_42006,N_42976);
nor U43641 (N_43641,N_42761,N_42030);
nor U43642 (N_43642,N_42328,N_42211);
nor U43643 (N_43643,N_42500,N_42577);
xor U43644 (N_43644,N_42691,N_42236);
nand U43645 (N_43645,N_42797,N_42289);
nor U43646 (N_43646,N_42605,N_42646);
nor U43647 (N_43647,N_42049,N_42031);
and U43648 (N_43648,N_42434,N_42253);
or U43649 (N_43649,N_42152,N_42297);
nor U43650 (N_43650,N_42866,N_42294);
or U43651 (N_43651,N_42916,N_42908);
nand U43652 (N_43652,N_42855,N_42965);
and U43653 (N_43653,N_42474,N_42965);
or U43654 (N_43654,N_42310,N_42874);
xor U43655 (N_43655,N_42644,N_42937);
nor U43656 (N_43656,N_42004,N_42486);
xor U43657 (N_43657,N_42527,N_42807);
nor U43658 (N_43658,N_42761,N_42733);
nor U43659 (N_43659,N_42406,N_42057);
or U43660 (N_43660,N_42583,N_42973);
or U43661 (N_43661,N_42121,N_42774);
or U43662 (N_43662,N_42555,N_42584);
nor U43663 (N_43663,N_42862,N_42688);
or U43664 (N_43664,N_42527,N_42105);
nor U43665 (N_43665,N_42419,N_42489);
nand U43666 (N_43666,N_42828,N_42608);
nand U43667 (N_43667,N_42300,N_42385);
nand U43668 (N_43668,N_42201,N_42671);
nand U43669 (N_43669,N_42651,N_42379);
and U43670 (N_43670,N_42366,N_42309);
nor U43671 (N_43671,N_42617,N_42954);
and U43672 (N_43672,N_42193,N_42981);
or U43673 (N_43673,N_42874,N_42010);
nand U43674 (N_43674,N_42518,N_42808);
and U43675 (N_43675,N_42800,N_42071);
xor U43676 (N_43676,N_42721,N_42588);
or U43677 (N_43677,N_42860,N_42585);
and U43678 (N_43678,N_42142,N_42772);
nand U43679 (N_43679,N_42055,N_42421);
nor U43680 (N_43680,N_42373,N_42146);
xnor U43681 (N_43681,N_42169,N_42484);
or U43682 (N_43682,N_42546,N_42909);
xnor U43683 (N_43683,N_42662,N_42276);
nand U43684 (N_43684,N_42522,N_42100);
nor U43685 (N_43685,N_42650,N_42198);
and U43686 (N_43686,N_42047,N_42108);
xnor U43687 (N_43687,N_42496,N_42131);
or U43688 (N_43688,N_42081,N_42253);
nand U43689 (N_43689,N_42156,N_42864);
and U43690 (N_43690,N_42510,N_42273);
nand U43691 (N_43691,N_42270,N_42853);
or U43692 (N_43692,N_42634,N_42505);
or U43693 (N_43693,N_42804,N_42299);
nand U43694 (N_43694,N_42436,N_42478);
nor U43695 (N_43695,N_42600,N_42610);
nor U43696 (N_43696,N_42611,N_42007);
nor U43697 (N_43697,N_42258,N_42465);
or U43698 (N_43698,N_42329,N_42296);
or U43699 (N_43699,N_42345,N_42562);
xor U43700 (N_43700,N_42937,N_42003);
nand U43701 (N_43701,N_42962,N_42616);
xor U43702 (N_43702,N_42379,N_42325);
and U43703 (N_43703,N_42831,N_42223);
nor U43704 (N_43704,N_42618,N_42774);
nand U43705 (N_43705,N_42009,N_42948);
nor U43706 (N_43706,N_42335,N_42640);
and U43707 (N_43707,N_42001,N_42552);
or U43708 (N_43708,N_42000,N_42001);
or U43709 (N_43709,N_42448,N_42135);
nor U43710 (N_43710,N_42242,N_42789);
and U43711 (N_43711,N_42785,N_42555);
or U43712 (N_43712,N_42986,N_42893);
nand U43713 (N_43713,N_42881,N_42928);
nand U43714 (N_43714,N_42862,N_42227);
xnor U43715 (N_43715,N_42993,N_42620);
nor U43716 (N_43716,N_42003,N_42789);
or U43717 (N_43717,N_42643,N_42180);
xor U43718 (N_43718,N_42098,N_42293);
or U43719 (N_43719,N_42471,N_42531);
nand U43720 (N_43720,N_42966,N_42432);
nor U43721 (N_43721,N_42232,N_42265);
nand U43722 (N_43722,N_42589,N_42602);
and U43723 (N_43723,N_42348,N_42693);
and U43724 (N_43724,N_42436,N_42308);
xor U43725 (N_43725,N_42515,N_42617);
and U43726 (N_43726,N_42664,N_42537);
nand U43727 (N_43727,N_42925,N_42908);
xor U43728 (N_43728,N_42694,N_42784);
nand U43729 (N_43729,N_42649,N_42514);
and U43730 (N_43730,N_42765,N_42750);
nor U43731 (N_43731,N_42630,N_42430);
nand U43732 (N_43732,N_42273,N_42708);
or U43733 (N_43733,N_42129,N_42652);
or U43734 (N_43734,N_42590,N_42291);
nand U43735 (N_43735,N_42679,N_42097);
and U43736 (N_43736,N_42409,N_42524);
xor U43737 (N_43737,N_42395,N_42134);
nand U43738 (N_43738,N_42936,N_42373);
xnor U43739 (N_43739,N_42026,N_42173);
or U43740 (N_43740,N_42949,N_42022);
nor U43741 (N_43741,N_42109,N_42780);
and U43742 (N_43742,N_42651,N_42314);
and U43743 (N_43743,N_42905,N_42669);
or U43744 (N_43744,N_42942,N_42070);
or U43745 (N_43745,N_42653,N_42865);
nand U43746 (N_43746,N_42676,N_42169);
xnor U43747 (N_43747,N_42466,N_42799);
xor U43748 (N_43748,N_42205,N_42477);
and U43749 (N_43749,N_42859,N_42805);
or U43750 (N_43750,N_42779,N_42321);
and U43751 (N_43751,N_42462,N_42339);
nand U43752 (N_43752,N_42348,N_42316);
or U43753 (N_43753,N_42431,N_42664);
or U43754 (N_43754,N_42797,N_42111);
nor U43755 (N_43755,N_42942,N_42389);
and U43756 (N_43756,N_42111,N_42986);
and U43757 (N_43757,N_42536,N_42401);
nor U43758 (N_43758,N_42705,N_42676);
or U43759 (N_43759,N_42379,N_42702);
nor U43760 (N_43760,N_42012,N_42820);
and U43761 (N_43761,N_42703,N_42849);
and U43762 (N_43762,N_42886,N_42505);
or U43763 (N_43763,N_42426,N_42454);
nor U43764 (N_43764,N_42678,N_42805);
nor U43765 (N_43765,N_42329,N_42419);
and U43766 (N_43766,N_42255,N_42632);
nand U43767 (N_43767,N_42274,N_42007);
xor U43768 (N_43768,N_42412,N_42184);
nand U43769 (N_43769,N_42520,N_42149);
and U43770 (N_43770,N_42646,N_42056);
and U43771 (N_43771,N_42910,N_42450);
nor U43772 (N_43772,N_42449,N_42487);
and U43773 (N_43773,N_42985,N_42280);
nand U43774 (N_43774,N_42980,N_42262);
nor U43775 (N_43775,N_42860,N_42008);
nand U43776 (N_43776,N_42564,N_42809);
and U43777 (N_43777,N_42360,N_42030);
and U43778 (N_43778,N_42458,N_42577);
or U43779 (N_43779,N_42896,N_42170);
nor U43780 (N_43780,N_42468,N_42056);
and U43781 (N_43781,N_42298,N_42933);
and U43782 (N_43782,N_42532,N_42629);
nand U43783 (N_43783,N_42697,N_42131);
nor U43784 (N_43784,N_42106,N_42901);
and U43785 (N_43785,N_42297,N_42399);
nand U43786 (N_43786,N_42449,N_42645);
nor U43787 (N_43787,N_42980,N_42369);
or U43788 (N_43788,N_42620,N_42712);
or U43789 (N_43789,N_42513,N_42611);
or U43790 (N_43790,N_42107,N_42560);
or U43791 (N_43791,N_42606,N_42391);
and U43792 (N_43792,N_42379,N_42611);
xnor U43793 (N_43793,N_42515,N_42878);
and U43794 (N_43794,N_42802,N_42827);
and U43795 (N_43795,N_42977,N_42105);
nand U43796 (N_43796,N_42716,N_42115);
or U43797 (N_43797,N_42435,N_42933);
xnor U43798 (N_43798,N_42943,N_42934);
and U43799 (N_43799,N_42850,N_42482);
xor U43800 (N_43800,N_42494,N_42637);
or U43801 (N_43801,N_42380,N_42825);
and U43802 (N_43802,N_42301,N_42387);
and U43803 (N_43803,N_42283,N_42810);
nand U43804 (N_43804,N_42897,N_42771);
or U43805 (N_43805,N_42039,N_42982);
or U43806 (N_43806,N_42781,N_42074);
nor U43807 (N_43807,N_42483,N_42845);
nand U43808 (N_43808,N_42312,N_42722);
nor U43809 (N_43809,N_42549,N_42634);
or U43810 (N_43810,N_42200,N_42965);
xor U43811 (N_43811,N_42830,N_42038);
and U43812 (N_43812,N_42782,N_42523);
nor U43813 (N_43813,N_42153,N_42423);
nor U43814 (N_43814,N_42884,N_42861);
or U43815 (N_43815,N_42185,N_42178);
xor U43816 (N_43816,N_42491,N_42798);
and U43817 (N_43817,N_42584,N_42305);
nor U43818 (N_43818,N_42606,N_42389);
or U43819 (N_43819,N_42074,N_42865);
xnor U43820 (N_43820,N_42699,N_42808);
xnor U43821 (N_43821,N_42727,N_42058);
or U43822 (N_43822,N_42853,N_42387);
nand U43823 (N_43823,N_42054,N_42875);
nor U43824 (N_43824,N_42829,N_42865);
or U43825 (N_43825,N_42077,N_42196);
and U43826 (N_43826,N_42445,N_42869);
nand U43827 (N_43827,N_42951,N_42342);
nor U43828 (N_43828,N_42858,N_42775);
and U43829 (N_43829,N_42451,N_42195);
nand U43830 (N_43830,N_42163,N_42822);
nor U43831 (N_43831,N_42780,N_42186);
and U43832 (N_43832,N_42794,N_42439);
nor U43833 (N_43833,N_42907,N_42433);
and U43834 (N_43834,N_42144,N_42762);
xnor U43835 (N_43835,N_42911,N_42853);
xnor U43836 (N_43836,N_42583,N_42901);
nand U43837 (N_43837,N_42362,N_42703);
nand U43838 (N_43838,N_42718,N_42963);
xnor U43839 (N_43839,N_42053,N_42279);
nor U43840 (N_43840,N_42626,N_42764);
xor U43841 (N_43841,N_42056,N_42039);
xnor U43842 (N_43842,N_42597,N_42724);
or U43843 (N_43843,N_42558,N_42367);
xnor U43844 (N_43844,N_42497,N_42394);
or U43845 (N_43845,N_42299,N_42785);
and U43846 (N_43846,N_42045,N_42411);
nor U43847 (N_43847,N_42420,N_42894);
and U43848 (N_43848,N_42787,N_42747);
nor U43849 (N_43849,N_42993,N_42613);
xor U43850 (N_43850,N_42199,N_42066);
or U43851 (N_43851,N_42269,N_42170);
and U43852 (N_43852,N_42986,N_42873);
or U43853 (N_43853,N_42717,N_42009);
nor U43854 (N_43854,N_42854,N_42815);
nor U43855 (N_43855,N_42371,N_42973);
nand U43856 (N_43856,N_42094,N_42160);
xor U43857 (N_43857,N_42542,N_42089);
nor U43858 (N_43858,N_42340,N_42548);
nor U43859 (N_43859,N_42050,N_42956);
and U43860 (N_43860,N_42555,N_42310);
xor U43861 (N_43861,N_42163,N_42323);
or U43862 (N_43862,N_42568,N_42392);
nand U43863 (N_43863,N_42431,N_42110);
nand U43864 (N_43864,N_42198,N_42015);
and U43865 (N_43865,N_42345,N_42754);
and U43866 (N_43866,N_42064,N_42880);
nand U43867 (N_43867,N_42826,N_42248);
or U43868 (N_43868,N_42272,N_42396);
xnor U43869 (N_43869,N_42437,N_42030);
or U43870 (N_43870,N_42701,N_42543);
and U43871 (N_43871,N_42547,N_42085);
xor U43872 (N_43872,N_42022,N_42672);
xor U43873 (N_43873,N_42720,N_42980);
and U43874 (N_43874,N_42619,N_42931);
nand U43875 (N_43875,N_42521,N_42285);
or U43876 (N_43876,N_42839,N_42205);
or U43877 (N_43877,N_42850,N_42911);
nor U43878 (N_43878,N_42857,N_42909);
nor U43879 (N_43879,N_42488,N_42413);
or U43880 (N_43880,N_42909,N_42758);
nor U43881 (N_43881,N_42247,N_42188);
nor U43882 (N_43882,N_42158,N_42316);
or U43883 (N_43883,N_42681,N_42034);
nor U43884 (N_43884,N_42991,N_42196);
and U43885 (N_43885,N_42295,N_42006);
nand U43886 (N_43886,N_42915,N_42572);
or U43887 (N_43887,N_42055,N_42404);
xor U43888 (N_43888,N_42274,N_42559);
and U43889 (N_43889,N_42559,N_42142);
or U43890 (N_43890,N_42981,N_42159);
and U43891 (N_43891,N_42839,N_42790);
xor U43892 (N_43892,N_42039,N_42557);
and U43893 (N_43893,N_42242,N_42671);
nand U43894 (N_43894,N_42190,N_42169);
and U43895 (N_43895,N_42294,N_42665);
xnor U43896 (N_43896,N_42667,N_42960);
nand U43897 (N_43897,N_42362,N_42068);
nand U43898 (N_43898,N_42087,N_42036);
and U43899 (N_43899,N_42577,N_42109);
nor U43900 (N_43900,N_42678,N_42819);
and U43901 (N_43901,N_42064,N_42721);
nor U43902 (N_43902,N_42597,N_42219);
nand U43903 (N_43903,N_42476,N_42533);
nand U43904 (N_43904,N_42732,N_42618);
or U43905 (N_43905,N_42163,N_42057);
xnor U43906 (N_43906,N_42735,N_42135);
and U43907 (N_43907,N_42987,N_42040);
nand U43908 (N_43908,N_42095,N_42782);
and U43909 (N_43909,N_42033,N_42548);
nor U43910 (N_43910,N_42210,N_42655);
or U43911 (N_43911,N_42809,N_42276);
nor U43912 (N_43912,N_42416,N_42178);
and U43913 (N_43913,N_42312,N_42887);
or U43914 (N_43914,N_42486,N_42948);
and U43915 (N_43915,N_42592,N_42674);
or U43916 (N_43916,N_42982,N_42001);
xor U43917 (N_43917,N_42792,N_42757);
nor U43918 (N_43918,N_42771,N_42237);
or U43919 (N_43919,N_42593,N_42339);
and U43920 (N_43920,N_42309,N_42843);
nor U43921 (N_43921,N_42417,N_42821);
xnor U43922 (N_43922,N_42838,N_42575);
nor U43923 (N_43923,N_42115,N_42086);
xor U43924 (N_43924,N_42176,N_42500);
or U43925 (N_43925,N_42612,N_42308);
and U43926 (N_43926,N_42411,N_42639);
and U43927 (N_43927,N_42487,N_42448);
nand U43928 (N_43928,N_42085,N_42314);
and U43929 (N_43929,N_42630,N_42458);
nand U43930 (N_43930,N_42391,N_42965);
nor U43931 (N_43931,N_42397,N_42177);
or U43932 (N_43932,N_42187,N_42681);
nor U43933 (N_43933,N_42186,N_42501);
or U43934 (N_43934,N_42140,N_42870);
nor U43935 (N_43935,N_42159,N_42735);
or U43936 (N_43936,N_42228,N_42065);
or U43937 (N_43937,N_42360,N_42521);
xnor U43938 (N_43938,N_42269,N_42320);
xor U43939 (N_43939,N_42052,N_42569);
xnor U43940 (N_43940,N_42693,N_42779);
nor U43941 (N_43941,N_42152,N_42216);
nand U43942 (N_43942,N_42234,N_42041);
xnor U43943 (N_43943,N_42753,N_42726);
and U43944 (N_43944,N_42672,N_42080);
nor U43945 (N_43945,N_42910,N_42272);
and U43946 (N_43946,N_42760,N_42031);
or U43947 (N_43947,N_42353,N_42244);
nor U43948 (N_43948,N_42709,N_42673);
or U43949 (N_43949,N_42450,N_42885);
nand U43950 (N_43950,N_42883,N_42224);
nand U43951 (N_43951,N_42535,N_42400);
and U43952 (N_43952,N_42586,N_42208);
xor U43953 (N_43953,N_42401,N_42065);
and U43954 (N_43954,N_42809,N_42349);
nand U43955 (N_43955,N_42665,N_42750);
xnor U43956 (N_43956,N_42212,N_42426);
or U43957 (N_43957,N_42397,N_42068);
or U43958 (N_43958,N_42306,N_42781);
nor U43959 (N_43959,N_42597,N_42619);
nor U43960 (N_43960,N_42131,N_42511);
nand U43961 (N_43961,N_42789,N_42743);
and U43962 (N_43962,N_42293,N_42237);
and U43963 (N_43963,N_42548,N_42287);
nor U43964 (N_43964,N_42637,N_42599);
nor U43965 (N_43965,N_42110,N_42418);
xnor U43966 (N_43966,N_42668,N_42507);
or U43967 (N_43967,N_42171,N_42278);
or U43968 (N_43968,N_42236,N_42067);
xor U43969 (N_43969,N_42006,N_42028);
xor U43970 (N_43970,N_42644,N_42679);
and U43971 (N_43971,N_42188,N_42881);
xor U43972 (N_43972,N_42825,N_42592);
xnor U43973 (N_43973,N_42486,N_42173);
xnor U43974 (N_43974,N_42674,N_42481);
and U43975 (N_43975,N_42734,N_42652);
xnor U43976 (N_43976,N_42082,N_42081);
nand U43977 (N_43977,N_42527,N_42051);
xor U43978 (N_43978,N_42223,N_42269);
and U43979 (N_43979,N_42672,N_42901);
xor U43980 (N_43980,N_42670,N_42784);
nor U43981 (N_43981,N_42667,N_42320);
and U43982 (N_43982,N_42160,N_42168);
nand U43983 (N_43983,N_42243,N_42231);
and U43984 (N_43984,N_42761,N_42664);
xnor U43985 (N_43985,N_42513,N_42209);
nor U43986 (N_43986,N_42248,N_42032);
and U43987 (N_43987,N_42353,N_42184);
xor U43988 (N_43988,N_42580,N_42905);
nor U43989 (N_43989,N_42019,N_42269);
xor U43990 (N_43990,N_42824,N_42733);
or U43991 (N_43991,N_42457,N_42771);
or U43992 (N_43992,N_42756,N_42131);
nor U43993 (N_43993,N_42129,N_42321);
nand U43994 (N_43994,N_42209,N_42891);
and U43995 (N_43995,N_42610,N_42940);
and U43996 (N_43996,N_42353,N_42417);
or U43997 (N_43997,N_42491,N_42151);
nand U43998 (N_43998,N_42964,N_42080);
nor U43999 (N_43999,N_42557,N_42124);
and U44000 (N_44000,N_43161,N_43266);
and U44001 (N_44001,N_43476,N_43379);
or U44002 (N_44002,N_43876,N_43365);
nand U44003 (N_44003,N_43736,N_43226);
xor U44004 (N_44004,N_43628,N_43335);
and U44005 (N_44005,N_43905,N_43245);
nor U44006 (N_44006,N_43268,N_43375);
xor U44007 (N_44007,N_43507,N_43349);
nor U44008 (N_44008,N_43851,N_43612);
nand U44009 (N_44009,N_43009,N_43844);
nand U44010 (N_44010,N_43216,N_43119);
nand U44011 (N_44011,N_43105,N_43630);
or U44012 (N_44012,N_43897,N_43000);
or U44013 (N_44013,N_43451,N_43635);
xor U44014 (N_44014,N_43791,N_43038);
xnor U44015 (N_44015,N_43445,N_43819);
and U44016 (N_44016,N_43544,N_43713);
or U44017 (N_44017,N_43735,N_43985);
or U44018 (N_44018,N_43106,N_43881);
or U44019 (N_44019,N_43475,N_43043);
or U44020 (N_44020,N_43502,N_43575);
nand U44021 (N_44021,N_43351,N_43213);
and U44022 (N_44022,N_43925,N_43298);
or U44023 (N_44023,N_43163,N_43899);
nand U44024 (N_44024,N_43829,N_43966);
nor U44025 (N_44025,N_43199,N_43793);
or U44026 (N_44026,N_43164,N_43509);
and U44027 (N_44027,N_43439,N_43825);
nand U44028 (N_44028,N_43267,N_43595);
xor U44029 (N_44029,N_43091,N_43691);
or U44030 (N_44030,N_43323,N_43577);
nand U44031 (N_44031,N_43535,N_43926);
nand U44032 (N_44032,N_43399,N_43328);
nand U44033 (N_44033,N_43653,N_43688);
nor U44034 (N_44034,N_43907,N_43121);
xnor U44035 (N_44035,N_43376,N_43358);
or U44036 (N_44036,N_43209,N_43046);
xor U44037 (N_44037,N_43415,N_43466);
or U44038 (N_44038,N_43553,N_43811);
or U44039 (N_44039,N_43533,N_43703);
and U44040 (N_44040,N_43371,N_43025);
nand U44041 (N_44041,N_43668,N_43240);
and U44042 (N_44042,N_43940,N_43711);
nand U44043 (N_44043,N_43853,N_43814);
nand U44044 (N_44044,N_43879,N_43370);
and U44045 (N_44045,N_43434,N_43319);
or U44046 (N_44046,N_43112,N_43249);
nand U44047 (N_44047,N_43798,N_43422);
xor U44048 (N_44048,N_43387,N_43759);
xor U44049 (N_44049,N_43331,N_43783);
xor U44050 (N_44050,N_43457,N_43887);
or U44051 (N_44051,N_43638,N_43733);
nor U44052 (N_44052,N_43598,N_43524);
and U44053 (N_44053,N_43490,N_43229);
or U44054 (N_44054,N_43311,N_43952);
and U44055 (N_44055,N_43421,N_43377);
nand U44056 (N_44056,N_43781,N_43418);
nor U44057 (N_44057,N_43359,N_43130);
and U44058 (N_44058,N_43679,N_43823);
nor U44059 (N_44059,N_43145,N_43054);
nor U44060 (N_44060,N_43655,N_43676);
and U44061 (N_44061,N_43090,N_43010);
nand U44062 (N_44062,N_43045,N_43522);
and U44063 (N_44063,N_43016,N_43546);
and U44064 (N_44064,N_43231,N_43717);
or U44065 (N_44065,N_43693,N_43132);
or U44066 (N_44066,N_43860,N_43114);
nand U44067 (N_44067,N_43945,N_43198);
and U44068 (N_44068,N_43013,N_43435);
nor U44069 (N_44069,N_43604,N_43083);
nand U44070 (N_44070,N_43067,N_43280);
or U44071 (N_44071,N_43382,N_43797);
or U44072 (N_44072,N_43874,N_43287);
nor U44073 (N_44073,N_43545,N_43726);
nor U44074 (N_44074,N_43138,N_43963);
xnor U44075 (N_44075,N_43867,N_43386);
nor U44076 (N_44076,N_43183,N_43714);
xor U44077 (N_44077,N_43766,N_43915);
or U44078 (N_44078,N_43018,N_43888);
or U44079 (N_44079,N_43957,N_43603);
nor U44080 (N_44080,N_43217,N_43548);
and U44081 (N_44081,N_43710,N_43931);
nand U44082 (N_44082,N_43086,N_43592);
and U44083 (N_44083,N_43750,N_43519);
or U44084 (N_44084,N_43402,N_43568);
nor U44085 (N_44085,N_43123,N_43656);
xnor U44086 (N_44086,N_43060,N_43803);
and U44087 (N_44087,N_43618,N_43185);
or U44088 (N_44088,N_43234,N_43134);
nor U44089 (N_44089,N_43196,N_43020);
or U44090 (N_44090,N_43409,N_43005);
nor U44091 (N_44091,N_43725,N_43934);
nand U44092 (N_44092,N_43184,N_43982);
nand U44093 (N_44093,N_43412,N_43109);
or U44094 (N_44094,N_43983,N_43933);
nor U44095 (N_44095,N_43133,N_43317);
nand U44096 (N_44096,N_43702,N_43274);
xor U44097 (N_44097,N_43030,N_43650);
nand U44098 (N_44098,N_43305,N_43450);
nand U44099 (N_44099,N_43805,N_43143);
nand U44100 (N_44100,N_43877,N_43828);
nand U44101 (N_44101,N_43673,N_43687);
or U44102 (N_44102,N_43340,N_43935);
nand U44103 (N_44103,N_43378,N_43438);
xnor U44104 (N_44104,N_43153,N_43115);
nor U44105 (N_44105,N_43707,N_43589);
nor U44106 (N_44106,N_43219,N_43740);
xnor U44107 (N_44107,N_43525,N_43116);
xor U44108 (N_44108,N_43355,N_43330);
nor U44109 (N_44109,N_43472,N_43316);
and U44110 (N_44110,N_43663,N_43389);
and U44111 (N_44111,N_43547,N_43858);
nor U44112 (N_44112,N_43523,N_43738);
nand U44113 (N_44113,N_43039,N_43639);
nor U44114 (N_44114,N_43100,N_43346);
nor U44115 (N_44115,N_43055,N_43194);
nand U44116 (N_44116,N_43747,N_43168);
or U44117 (N_44117,N_43843,N_43824);
nand U44118 (N_44118,N_43799,N_43079);
xnor U44119 (N_44119,N_43660,N_43596);
nand U44120 (N_44120,N_43066,N_43255);
and U44121 (N_44121,N_43857,N_43357);
and U44122 (N_44122,N_43873,N_43667);
or U44123 (N_44123,N_43428,N_43372);
nor U44124 (N_44124,N_43689,N_43871);
xnor U44125 (N_44125,N_43260,N_43125);
nand U44126 (N_44126,N_43035,N_43403);
and U44127 (N_44127,N_43930,N_43141);
or U44128 (N_44128,N_43098,N_43580);
or U44129 (N_44129,N_43302,N_43579);
xor U44130 (N_44130,N_43962,N_43795);
xor U44131 (N_44131,N_43006,N_43356);
nand U44132 (N_44132,N_43373,N_43481);
or U44133 (N_44133,N_43773,N_43835);
nor U44134 (N_44134,N_43051,N_43752);
and U44135 (N_44135,N_43980,N_43654);
and U44136 (N_44136,N_43836,N_43352);
and U44137 (N_44137,N_43761,N_43210);
nand U44138 (N_44138,N_43608,N_43891);
xor U44139 (N_44139,N_43426,N_43406);
nand U44140 (N_44140,N_43777,N_43631);
or U44141 (N_44141,N_43584,N_43642);
and U44142 (N_44142,N_43669,N_43646);
or U44143 (N_44143,N_43447,N_43276);
and U44144 (N_44144,N_43151,N_43961);
xor U44145 (N_44145,N_43901,N_43776);
and U44146 (N_44146,N_43671,N_43674);
and U44147 (N_44147,N_43498,N_43609);
nand U44148 (N_44148,N_43221,N_43363);
or U44149 (N_44149,N_43032,N_43895);
and U44150 (N_44150,N_43692,N_43413);
or U44151 (N_44151,N_43062,N_43444);
and U44152 (N_44152,N_43503,N_43237);
or U44153 (N_44153,N_43162,N_43566);
or U44154 (N_44154,N_43479,N_43286);
xor U44155 (N_44155,N_43753,N_43859);
xnor U44156 (N_44156,N_43520,N_43576);
and U44157 (N_44157,N_43064,N_43206);
xor U44158 (N_44158,N_43443,N_43456);
nand U44159 (N_44159,N_43970,N_43094);
and U44160 (N_44160,N_43549,N_43588);
or U44161 (N_44161,N_43212,N_43353);
or U44162 (N_44162,N_43607,N_43890);
or U44163 (N_44163,N_43366,N_43977);
or U44164 (N_44164,N_43556,N_43265);
nor U44165 (N_44165,N_43801,N_43361);
and U44166 (N_44166,N_43527,N_43807);
nor U44167 (N_44167,N_43581,N_43227);
and U44168 (N_44168,N_43611,N_43495);
xor U44169 (N_44169,N_43658,N_43170);
nor U44170 (N_44170,N_43284,N_43385);
xnor U44171 (N_44171,N_43492,N_43336);
or U44172 (N_44172,N_43437,N_43820);
nor U44173 (N_44173,N_43939,N_43263);
or U44174 (N_44174,N_43880,N_43754);
nor U44175 (N_44175,N_43312,N_43041);
nand U44176 (N_44176,N_43292,N_43780);
or U44177 (N_44177,N_43313,N_43069);
and U44178 (N_44178,N_43176,N_43900);
nor U44179 (N_44179,N_43026,N_43560);
and U44180 (N_44180,N_43295,N_43892);
nor U44181 (N_44181,N_43281,N_43306);
nand U44182 (N_44182,N_43433,N_43345);
nand U44183 (N_44183,N_43414,N_43918);
nand U44184 (N_44184,N_43526,N_43827);
or U44185 (N_44185,N_43465,N_43728);
nand U44186 (N_44186,N_43474,N_43214);
and U44187 (N_44187,N_43137,N_43790);
or U44188 (N_44188,N_43037,N_43657);
nor U44189 (N_44189,N_43264,N_43486);
or U44190 (N_44190,N_43193,N_43028);
and U44191 (N_44191,N_43104,N_43648);
and U44192 (N_44192,N_43369,N_43582);
nor U44193 (N_44193,N_43448,N_43171);
nor U44194 (N_44194,N_43076,N_43324);
xor U44195 (N_44195,N_43429,N_43716);
xor U44196 (N_44196,N_43022,N_43297);
nor U44197 (N_44197,N_43454,N_43757);
xor U44198 (N_44198,N_43056,N_43001);
xnor U44199 (N_44199,N_43570,N_43246);
xnor U44200 (N_44200,N_43937,N_43273);
xor U44201 (N_44201,N_43911,N_43529);
xnor U44202 (N_44202,N_43861,N_43508);
and U44203 (N_44203,N_43473,N_43742);
nor U44204 (N_44204,N_43616,N_43468);
and U44205 (N_44205,N_43626,N_43124);
or U44206 (N_44206,N_43845,N_43909);
nor U44207 (N_44207,N_43511,N_43749);
nand U44208 (N_44208,N_43211,N_43620);
nor U44209 (N_44209,N_43694,N_43951);
and U44210 (N_44210,N_43586,N_43459);
xor U44211 (N_44211,N_43131,N_43659);
or U44212 (N_44212,N_43597,N_43169);
or U44213 (N_44213,N_43095,N_43093);
nand U44214 (N_44214,N_43097,N_43649);
and U44215 (N_44215,N_43397,N_43826);
nor U44216 (N_44216,N_43117,N_43774);
xnor U44217 (N_44217,N_43622,N_43243);
nand U44218 (N_44218,N_43103,N_43269);
or U44219 (N_44219,N_43082,N_43247);
and U44220 (N_44220,N_43436,N_43070);
xor U44221 (N_44221,N_43325,N_43561);
xnor U44222 (N_44222,N_43721,N_43441);
and U44223 (N_44223,N_43470,N_43758);
nor U44224 (N_44224,N_43973,N_43496);
xnor U44225 (N_44225,N_43763,N_43239);
or U44226 (N_44226,N_43233,N_43883);
xor U44227 (N_44227,N_43021,N_43619);
or U44228 (N_44228,N_43555,N_43380);
or U44229 (N_44229,N_43917,N_43333);
xor U44230 (N_44230,N_43965,N_43849);
or U44231 (N_44231,N_43381,N_43613);
and U44232 (N_44232,N_43984,N_43338);
nor U44233 (N_44233,N_43585,N_43832);
and U44234 (N_44234,N_43680,N_43583);
and U44235 (N_44235,N_43995,N_43411);
or U44236 (N_44236,N_43257,N_43099);
nand U44237 (N_44237,N_43539,N_43870);
nand U44238 (N_44238,N_43610,N_43019);
nand U44239 (N_44239,N_43187,N_43310);
or U44240 (N_44240,N_43731,N_43727);
xor U44241 (N_44241,N_43485,N_43572);
xor U44242 (N_44242,N_43948,N_43174);
nor U44243 (N_44243,N_43856,N_43218);
xor U44244 (N_44244,N_43499,N_43894);
xor U44245 (N_44245,N_43606,N_43244);
xor U44246 (N_44246,N_43514,N_43990);
nand U44247 (N_44247,N_43532,N_43782);
nor U44248 (N_44248,N_43347,N_43512);
nand U44249 (N_44249,N_43953,N_43500);
nand U44250 (N_44250,N_43329,N_43388);
xor U44251 (N_44251,N_43912,N_43815);
or U44252 (N_44252,N_43812,N_43741);
nor U44253 (N_44253,N_43664,N_43339);
xor U44254 (N_44254,N_43775,N_43755);
and U44255 (N_44255,N_43943,N_43154);
or U44256 (N_44256,N_43368,N_43075);
nor U44257 (N_44257,N_43061,N_43991);
or U44258 (N_44258,N_43182,N_43932);
or U44259 (N_44259,N_43872,N_43573);
xor U44260 (N_44260,N_43241,N_43981);
or U44261 (N_44261,N_43559,N_43924);
nor U44262 (N_44262,N_43308,N_43960);
or U44263 (N_44263,N_43954,N_43487);
nand U44264 (N_44264,N_43294,N_43250);
nor U44265 (N_44265,N_43040,N_43967);
and U44266 (N_44266,N_43108,N_43847);
nand U44267 (N_44267,N_43551,N_43684);
or U44268 (N_44268,N_43031,N_43304);
and U44269 (N_44269,N_43959,N_43629);
nor U44270 (N_44270,N_43863,N_43748);
and U44271 (N_44271,N_43751,N_43955);
and U44272 (N_44272,N_43947,N_43665);
nor U44273 (N_44273,N_43530,N_43065);
and U44274 (N_44274,N_43334,N_43878);
and U44275 (N_44275,N_43173,N_43446);
or U44276 (N_44276,N_43299,N_43223);
nor U44277 (N_44277,N_43600,N_43969);
and U44278 (N_44278,N_43786,N_43148);
or U44279 (N_44279,N_43567,N_43279);
nor U44280 (N_44280,N_43166,N_43192);
and U44281 (N_44281,N_43842,N_43057);
nand U44282 (N_44282,N_43675,N_43698);
nor U44283 (N_44283,N_43362,N_43706);
nor U44284 (N_44284,N_43332,N_43073);
xor U44285 (N_44285,N_43813,N_43405);
or U44286 (N_44286,N_43278,N_43391);
nor U44287 (N_44287,N_43058,N_43146);
or U44288 (N_44288,N_43404,N_43913);
and U44289 (N_44289,N_43623,N_43569);
and U44290 (N_44290,N_43225,N_43126);
nor U44291 (N_44291,N_43200,N_43467);
nand U44292 (N_44292,N_43550,N_43804);
xnor U44293 (N_44293,N_43762,N_43140);
or U44294 (N_44294,N_43477,N_43175);
and U44295 (N_44295,N_43601,N_43301);
or U44296 (N_44296,N_43928,N_43017);
or U44297 (N_44297,N_43998,N_43833);
nor U44298 (N_44298,N_43430,N_43427);
nor U44299 (N_44299,N_43886,N_43158);
nor U44300 (N_44300,N_43997,N_43846);
and U44301 (N_44301,N_43270,N_43723);
or U44302 (N_44302,N_43670,N_43760);
nand U44303 (N_44303,N_43864,N_43855);
nor U44304 (N_44304,N_43767,N_43700);
nand U44305 (N_44305,N_43516,N_43699);
nor U44306 (N_44306,N_43591,N_43189);
nor U44307 (N_44307,N_43191,N_43293);
or U44308 (N_44308,N_43341,N_43033);
and U44309 (N_44309,N_43096,N_43578);
or U44310 (N_44310,N_43205,N_43645);
nor U44311 (N_44311,N_43921,N_43142);
nor U44312 (N_44312,N_43077,N_43734);
nand U44313 (N_44313,N_43722,N_43528);
nand U44314 (N_44314,N_43431,N_43197);
or U44315 (N_44315,N_43252,N_43074);
or U44316 (N_44316,N_43557,N_43398);
and U44317 (N_44317,N_43806,N_43204);
and U44318 (N_44318,N_43882,N_43838);
xnor U44319 (N_44319,N_43417,N_43682);
and U44320 (N_44320,N_43558,N_43034);
or U44321 (N_44321,N_43541,N_43690);
or U44322 (N_44322,N_43986,N_43203);
nand U44323 (N_44323,N_43617,N_43309);
or U44324 (N_44324,N_43283,N_43666);
xor U44325 (N_44325,N_43364,N_43460);
or U44326 (N_44326,N_43464,N_43513);
and U44327 (N_44327,N_43300,N_43071);
or U44328 (N_44328,N_43012,N_43809);
and U44329 (N_44329,N_43420,N_43615);
nand U44330 (N_44330,N_43230,N_43469);
nor U44331 (N_44331,N_43136,N_43342);
and U44332 (N_44332,N_43976,N_43718);
and U44333 (N_44333,N_43261,N_43303);
xnor U44334 (N_44334,N_43181,N_43936);
nor U44335 (N_44335,N_43228,N_43172);
nand U44336 (N_44336,N_43150,N_43662);
nand U44337 (N_44337,N_43400,N_43408);
nor U44338 (N_44338,N_43686,N_43078);
nor U44339 (N_44339,N_43709,N_43044);
and U44340 (N_44340,N_43903,N_43517);
nor U44341 (N_44341,N_43251,N_43188);
xor U44342 (N_44342,N_43552,N_43452);
xnor U44343 (N_44343,N_43092,N_43139);
xor U44344 (N_44344,N_43157,N_43587);
xor U44345 (N_44345,N_43875,N_43272);
nor U44346 (N_44346,N_43705,N_43993);
nand U44347 (N_44347,N_43994,N_43730);
nand U44348 (N_44348,N_43484,N_43506);
nand U44349 (N_44349,N_43180,N_43023);
nor U44350 (N_44350,N_43633,N_43048);
or U44351 (N_44351,N_43854,N_43215);
nand U44352 (N_44352,N_43177,N_43771);
and U44353 (N_44353,N_43968,N_43958);
xnor U44354 (N_44354,N_43063,N_43564);
nor U44355 (N_44355,N_43049,N_43536);
nand U44356 (N_44356,N_43015,N_43908);
xnor U44357 (N_44357,N_43808,N_43964);
and U44358 (N_44358,N_43478,N_43831);
nor U44359 (N_44359,N_43505,N_43321);
or U44360 (N_44360,N_43636,N_43111);
nand U44361 (N_44361,N_43322,N_43393);
nand U44362 (N_44362,N_43396,N_43354);
and U44363 (N_44363,N_43384,N_43974);
or U44364 (N_44364,N_43110,N_43080);
nand U44365 (N_44365,N_43565,N_43971);
xnor U44366 (N_44366,N_43765,N_43314);
nor U44367 (N_44367,N_43036,N_43785);
and U44368 (N_44368,N_43120,N_43160);
nand U44369 (N_44369,N_43254,N_43344);
xnor U44370 (N_44370,N_43769,N_43236);
nor U44371 (N_44371,N_43916,N_43839);
or U44372 (N_44372,N_43594,N_43850);
nor U44373 (N_44373,N_43944,N_43195);
or U44374 (N_44374,N_43089,N_43996);
or U44375 (N_44375,N_43271,N_43003);
xnor U44376 (N_44376,N_43896,N_43992);
or U44377 (N_44377,N_43778,N_43374);
or U44378 (N_44378,N_43852,N_43571);
xor U44379 (N_44379,N_43802,N_43866);
nand U44380 (N_44380,N_43988,N_43817);
xor U44381 (N_44381,N_43059,N_43461);
nand U44382 (N_44382,N_43898,N_43834);
nor U44383 (N_44383,N_43122,N_43701);
and U44384 (N_44384,N_43326,N_43220);
xor U44385 (N_44385,N_43602,N_43149);
and U44386 (N_44386,N_43350,N_43772);
nand U44387 (N_44387,N_43462,N_43488);
or U44388 (N_44388,N_43737,N_43262);
xor U44389 (N_44389,N_43590,N_43614);
or U44390 (N_44390,N_43296,N_43764);
nor U44391 (N_44391,N_43989,N_43489);
nand U44392 (N_44392,N_43914,N_43455);
and U44393 (N_44393,N_43315,N_43885);
nor U44394 (N_44394,N_43789,N_43410);
and U44395 (N_44395,N_43238,N_43837);
nand U44396 (N_44396,N_43922,N_43841);
or U44397 (N_44397,N_43088,N_43232);
and U44398 (N_44398,N_43956,N_43715);
nor U44399 (N_44399,N_43190,N_43416);
or U44400 (N_44400,N_43792,N_43949);
and U44401 (N_44401,N_43796,N_43178);
nor U44402 (N_44402,N_43179,N_43155);
xor U44403 (N_44403,N_43307,N_43128);
and U44404 (N_44404,N_43840,N_43643);
xnor U44405 (N_44405,N_43756,N_43637);
nand U44406 (N_44406,N_43927,N_43599);
or U44407 (N_44407,N_43862,N_43563);
or U44408 (N_44408,N_43222,N_43493);
xnor U44409 (N_44409,N_43147,N_43027);
xor U44410 (N_44410,N_43050,N_43343);
nand U44411 (N_44411,N_43007,N_43652);
nor U44412 (N_44412,N_43542,N_43129);
or U44413 (N_44413,N_43562,N_43113);
or U44414 (N_44414,N_43784,N_43440);
and U44415 (N_44415,N_43975,N_43681);
or U44416 (N_44416,N_43685,N_43004);
and U44417 (N_44417,N_43515,N_43830);
or U44418 (N_44418,N_43739,N_43906);
xor U44419 (N_44419,N_43661,N_43282);
nand U44420 (N_44420,N_43938,N_43729);
or U44421 (N_44421,N_43395,N_43256);
xnor U44422 (N_44422,N_43627,N_43518);
xor U44423 (N_44423,N_43208,N_43770);
and U44424 (N_44424,N_43538,N_43081);
xor U44425 (N_44425,N_43288,N_43248);
nor U44426 (N_44426,N_43869,N_43253);
and U44427 (N_44427,N_43102,N_43677);
and U44428 (N_44428,N_43678,N_43695);
nand U44429 (N_44429,N_43107,N_43242);
nor U44430 (N_44430,N_43442,N_43320);
nor U44431 (N_44431,N_43543,N_43712);
xor U44432 (N_44432,N_43640,N_43053);
or U44433 (N_44433,N_43011,N_43024);
and U44434 (N_44434,N_43165,N_43497);
nor U44435 (N_44435,N_43978,N_43277);
nand U44436 (N_44436,N_43072,N_43534);
xnor U44437 (N_44437,N_43085,N_43144);
nand U44438 (N_44438,N_43821,N_43779);
or U44439 (N_44439,N_43014,N_43697);
nand U44440 (N_44440,N_43720,N_43127);
and U44441 (N_44441,N_43482,N_43624);
xnor U44442 (N_44442,N_43979,N_43008);
nand U44443 (N_44443,N_43800,N_43290);
xnor U44444 (N_44444,N_43383,N_43367);
and U44445 (N_44445,N_43491,N_43647);
xnor U44446 (N_44446,N_43152,N_43285);
nor U44447 (N_44447,N_43719,N_43794);
nor U44448 (N_44448,N_43818,N_43101);
nor U44449 (N_44449,N_43327,N_43787);
or U44450 (N_44450,N_43425,N_43291);
and U44451 (N_44451,N_43724,N_43972);
and U44452 (N_44452,N_43593,N_43202);
nand U44453 (N_44453,N_43480,N_43118);
nor U44454 (N_44454,N_43704,N_43651);
nor U44455 (N_44455,N_43946,N_43531);
nand U44456 (N_44456,N_43167,N_43625);
and U44457 (N_44457,N_43999,N_43942);
nand U44458 (N_44458,N_43463,N_43390);
nand U44459 (N_44459,N_43458,N_43510);
or U44460 (N_44460,N_43159,N_43904);
or U44461 (N_44461,N_43521,N_43068);
xnor U44462 (N_44462,N_43893,N_43941);
nand U44463 (N_44463,N_43258,N_43052);
nand U44464 (N_44464,N_43047,N_43042);
xnor U44465 (N_44465,N_43186,N_43224);
nand U44466 (N_44466,N_43453,N_43848);
or U44467 (N_44467,N_43424,N_43449);
nand U44468 (N_44468,N_43884,N_43407);
xnor U44469 (N_44469,N_43201,N_43360);
nand U44470 (N_44470,N_43494,N_43275);
nand U44471 (N_44471,N_43683,N_43923);
xor U44472 (N_44472,N_43289,N_43135);
nor U44473 (N_44473,N_43337,N_43394);
nand U44474 (N_44474,N_43696,N_43259);
nand U44475 (N_44475,N_43348,N_43029);
or U44476 (N_44476,N_43574,N_43621);
xnor U44477 (N_44477,N_43540,N_43641);
nand U44478 (N_44478,N_43605,N_43919);
and U44479 (N_44479,N_43889,N_43920);
xor U44480 (N_44480,N_43235,N_43392);
xnor U44481 (N_44481,N_43554,N_43419);
and U44482 (N_44482,N_43744,N_43087);
or U44483 (N_44483,N_43207,N_43432);
and U44484 (N_44484,N_43632,N_43788);
and U44485 (N_44485,N_43483,N_43987);
and U44486 (N_44486,N_43501,N_43156);
xor U44487 (N_44487,N_43810,N_43708);
nand U44488 (N_44488,N_43537,N_43084);
nor U44489 (N_44489,N_43822,N_43318);
and U44490 (N_44490,N_43002,N_43865);
xnor U44491 (N_44491,N_43746,N_43743);
nor U44492 (N_44492,N_43950,N_43816);
and U44493 (N_44493,N_43634,N_43868);
nor U44494 (N_44494,N_43732,N_43644);
nand U44495 (N_44495,N_43929,N_43401);
xnor U44496 (N_44496,N_43423,N_43745);
and U44497 (N_44497,N_43768,N_43504);
and U44498 (N_44498,N_43902,N_43471);
or U44499 (N_44499,N_43672,N_43910);
nand U44500 (N_44500,N_43889,N_43150);
xnor U44501 (N_44501,N_43260,N_43043);
or U44502 (N_44502,N_43249,N_43752);
or U44503 (N_44503,N_43198,N_43894);
nor U44504 (N_44504,N_43959,N_43892);
nor U44505 (N_44505,N_43360,N_43925);
and U44506 (N_44506,N_43953,N_43085);
nand U44507 (N_44507,N_43634,N_43150);
and U44508 (N_44508,N_43178,N_43709);
or U44509 (N_44509,N_43021,N_43865);
nor U44510 (N_44510,N_43700,N_43529);
and U44511 (N_44511,N_43471,N_43402);
xor U44512 (N_44512,N_43213,N_43994);
or U44513 (N_44513,N_43916,N_43659);
or U44514 (N_44514,N_43424,N_43648);
xor U44515 (N_44515,N_43740,N_43368);
or U44516 (N_44516,N_43239,N_43621);
and U44517 (N_44517,N_43245,N_43166);
or U44518 (N_44518,N_43171,N_43424);
and U44519 (N_44519,N_43791,N_43079);
xnor U44520 (N_44520,N_43431,N_43166);
and U44521 (N_44521,N_43375,N_43317);
xor U44522 (N_44522,N_43393,N_43034);
xnor U44523 (N_44523,N_43298,N_43946);
nand U44524 (N_44524,N_43106,N_43724);
or U44525 (N_44525,N_43769,N_43594);
xor U44526 (N_44526,N_43279,N_43682);
or U44527 (N_44527,N_43246,N_43521);
xnor U44528 (N_44528,N_43541,N_43669);
and U44529 (N_44529,N_43288,N_43173);
xnor U44530 (N_44530,N_43640,N_43437);
nor U44531 (N_44531,N_43932,N_43881);
nor U44532 (N_44532,N_43110,N_43069);
or U44533 (N_44533,N_43267,N_43867);
xor U44534 (N_44534,N_43261,N_43662);
nor U44535 (N_44535,N_43756,N_43702);
or U44536 (N_44536,N_43357,N_43387);
xor U44537 (N_44537,N_43734,N_43841);
xor U44538 (N_44538,N_43227,N_43405);
nor U44539 (N_44539,N_43767,N_43518);
nand U44540 (N_44540,N_43748,N_43035);
nor U44541 (N_44541,N_43637,N_43113);
or U44542 (N_44542,N_43022,N_43750);
nor U44543 (N_44543,N_43164,N_43871);
or U44544 (N_44544,N_43817,N_43854);
or U44545 (N_44545,N_43407,N_43215);
and U44546 (N_44546,N_43655,N_43553);
and U44547 (N_44547,N_43648,N_43804);
nor U44548 (N_44548,N_43065,N_43642);
nor U44549 (N_44549,N_43944,N_43425);
nand U44550 (N_44550,N_43680,N_43828);
or U44551 (N_44551,N_43485,N_43881);
nor U44552 (N_44552,N_43440,N_43967);
xnor U44553 (N_44553,N_43319,N_43828);
xor U44554 (N_44554,N_43101,N_43325);
xor U44555 (N_44555,N_43141,N_43476);
nor U44556 (N_44556,N_43866,N_43848);
nor U44557 (N_44557,N_43252,N_43928);
xnor U44558 (N_44558,N_43769,N_43945);
xor U44559 (N_44559,N_43607,N_43500);
xnor U44560 (N_44560,N_43120,N_43781);
or U44561 (N_44561,N_43732,N_43388);
and U44562 (N_44562,N_43345,N_43277);
or U44563 (N_44563,N_43891,N_43298);
or U44564 (N_44564,N_43999,N_43687);
nand U44565 (N_44565,N_43330,N_43252);
or U44566 (N_44566,N_43136,N_43641);
nand U44567 (N_44567,N_43032,N_43827);
xnor U44568 (N_44568,N_43017,N_43060);
nand U44569 (N_44569,N_43997,N_43671);
xnor U44570 (N_44570,N_43820,N_43384);
xor U44571 (N_44571,N_43828,N_43250);
xor U44572 (N_44572,N_43756,N_43834);
nor U44573 (N_44573,N_43353,N_43889);
and U44574 (N_44574,N_43372,N_43016);
or U44575 (N_44575,N_43960,N_43275);
nand U44576 (N_44576,N_43654,N_43882);
or U44577 (N_44577,N_43201,N_43037);
and U44578 (N_44578,N_43870,N_43268);
nand U44579 (N_44579,N_43181,N_43420);
or U44580 (N_44580,N_43644,N_43999);
xnor U44581 (N_44581,N_43599,N_43078);
or U44582 (N_44582,N_43780,N_43489);
xnor U44583 (N_44583,N_43340,N_43094);
xor U44584 (N_44584,N_43202,N_43922);
and U44585 (N_44585,N_43212,N_43972);
and U44586 (N_44586,N_43723,N_43740);
and U44587 (N_44587,N_43188,N_43191);
and U44588 (N_44588,N_43608,N_43469);
and U44589 (N_44589,N_43463,N_43158);
nor U44590 (N_44590,N_43840,N_43243);
and U44591 (N_44591,N_43705,N_43597);
nand U44592 (N_44592,N_43627,N_43488);
and U44593 (N_44593,N_43807,N_43233);
nand U44594 (N_44594,N_43513,N_43081);
xnor U44595 (N_44595,N_43932,N_43548);
and U44596 (N_44596,N_43661,N_43708);
nor U44597 (N_44597,N_43160,N_43118);
and U44598 (N_44598,N_43833,N_43168);
or U44599 (N_44599,N_43287,N_43817);
or U44600 (N_44600,N_43786,N_43168);
nor U44601 (N_44601,N_43380,N_43841);
nor U44602 (N_44602,N_43592,N_43966);
xor U44603 (N_44603,N_43639,N_43121);
and U44604 (N_44604,N_43642,N_43594);
xnor U44605 (N_44605,N_43363,N_43339);
nand U44606 (N_44606,N_43758,N_43621);
xor U44607 (N_44607,N_43484,N_43109);
and U44608 (N_44608,N_43176,N_43867);
or U44609 (N_44609,N_43230,N_43982);
nand U44610 (N_44610,N_43540,N_43901);
and U44611 (N_44611,N_43151,N_43285);
xor U44612 (N_44612,N_43437,N_43165);
nand U44613 (N_44613,N_43601,N_43419);
or U44614 (N_44614,N_43907,N_43145);
nand U44615 (N_44615,N_43941,N_43085);
xor U44616 (N_44616,N_43865,N_43738);
nor U44617 (N_44617,N_43766,N_43075);
nor U44618 (N_44618,N_43011,N_43056);
nand U44619 (N_44619,N_43641,N_43188);
or U44620 (N_44620,N_43509,N_43161);
and U44621 (N_44621,N_43739,N_43813);
and U44622 (N_44622,N_43575,N_43556);
and U44623 (N_44623,N_43300,N_43891);
and U44624 (N_44624,N_43425,N_43410);
and U44625 (N_44625,N_43522,N_43114);
nor U44626 (N_44626,N_43136,N_43396);
and U44627 (N_44627,N_43835,N_43963);
and U44628 (N_44628,N_43362,N_43669);
or U44629 (N_44629,N_43194,N_43756);
or U44630 (N_44630,N_43484,N_43111);
xnor U44631 (N_44631,N_43561,N_43507);
or U44632 (N_44632,N_43691,N_43040);
nor U44633 (N_44633,N_43685,N_43562);
nor U44634 (N_44634,N_43662,N_43891);
nand U44635 (N_44635,N_43454,N_43776);
nor U44636 (N_44636,N_43321,N_43893);
or U44637 (N_44637,N_43059,N_43755);
or U44638 (N_44638,N_43319,N_43537);
nor U44639 (N_44639,N_43580,N_43035);
nand U44640 (N_44640,N_43381,N_43228);
xor U44641 (N_44641,N_43841,N_43846);
nor U44642 (N_44642,N_43907,N_43150);
nor U44643 (N_44643,N_43470,N_43916);
or U44644 (N_44644,N_43572,N_43685);
xor U44645 (N_44645,N_43889,N_43255);
xor U44646 (N_44646,N_43597,N_43898);
nand U44647 (N_44647,N_43714,N_43992);
xnor U44648 (N_44648,N_43359,N_43727);
and U44649 (N_44649,N_43112,N_43070);
and U44650 (N_44650,N_43279,N_43975);
xnor U44651 (N_44651,N_43214,N_43073);
or U44652 (N_44652,N_43792,N_43454);
xor U44653 (N_44653,N_43247,N_43348);
and U44654 (N_44654,N_43687,N_43503);
or U44655 (N_44655,N_43744,N_43509);
and U44656 (N_44656,N_43434,N_43645);
nand U44657 (N_44657,N_43181,N_43522);
or U44658 (N_44658,N_43704,N_43298);
and U44659 (N_44659,N_43427,N_43564);
nand U44660 (N_44660,N_43541,N_43995);
xnor U44661 (N_44661,N_43804,N_43966);
or U44662 (N_44662,N_43437,N_43579);
xor U44663 (N_44663,N_43172,N_43842);
nor U44664 (N_44664,N_43760,N_43711);
xor U44665 (N_44665,N_43998,N_43075);
nor U44666 (N_44666,N_43694,N_43481);
nor U44667 (N_44667,N_43575,N_43838);
xnor U44668 (N_44668,N_43857,N_43907);
nor U44669 (N_44669,N_43512,N_43516);
nor U44670 (N_44670,N_43803,N_43686);
and U44671 (N_44671,N_43175,N_43533);
and U44672 (N_44672,N_43006,N_43934);
nor U44673 (N_44673,N_43789,N_43703);
or U44674 (N_44674,N_43421,N_43438);
nor U44675 (N_44675,N_43907,N_43140);
nor U44676 (N_44676,N_43410,N_43436);
and U44677 (N_44677,N_43332,N_43887);
or U44678 (N_44678,N_43545,N_43246);
nand U44679 (N_44679,N_43534,N_43516);
and U44680 (N_44680,N_43849,N_43440);
and U44681 (N_44681,N_43053,N_43421);
and U44682 (N_44682,N_43466,N_43149);
and U44683 (N_44683,N_43865,N_43753);
nor U44684 (N_44684,N_43073,N_43506);
or U44685 (N_44685,N_43375,N_43281);
nor U44686 (N_44686,N_43512,N_43207);
or U44687 (N_44687,N_43659,N_43023);
or U44688 (N_44688,N_43063,N_43668);
and U44689 (N_44689,N_43350,N_43288);
xor U44690 (N_44690,N_43934,N_43580);
or U44691 (N_44691,N_43610,N_43724);
nand U44692 (N_44692,N_43421,N_43593);
xnor U44693 (N_44693,N_43897,N_43053);
nor U44694 (N_44694,N_43353,N_43643);
nor U44695 (N_44695,N_43731,N_43138);
and U44696 (N_44696,N_43419,N_43174);
xnor U44697 (N_44697,N_43758,N_43354);
xnor U44698 (N_44698,N_43024,N_43575);
nand U44699 (N_44699,N_43328,N_43684);
xor U44700 (N_44700,N_43684,N_43289);
xor U44701 (N_44701,N_43535,N_43005);
nor U44702 (N_44702,N_43912,N_43115);
and U44703 (N_44703,N_43447,N_43465);
and U44704 (N_44704,N_43739,N_43231);
and U44705 (N_44705,N_43819,N_43017);
nand U44706 (N_44706,N_43653,N_43996);
or U44707 (N_44707,N_43620,N_43593);
nor U44708 (N_44708,N_43168,N_43665);
xnor U44709 (N_44709,N_43887,N_43765);
or U44710 (N_44710,N_43140,N_43849);
or U44711 (N_44711,N_43454,N_43952);
nor U44712 (N_44712,N_43867,N_43754);
nor U44713 (N_44713,N_43938,N_43575);
or U44714 (N_44714,N_43264,N_43911);
xnor U44715 (N_44715,N_43613,N_43992);
nand U44716 (N_44716,N_43045,N_43872);
xor U44717 (N_44717,N_43270,N_43721);
nor U44718 (N_44718,N_43677,N_43348);
nor U44719 (N_44719,N_43581,N_43150);
xnor U44720 (N_44720,N_43317,N_43077);
nor U44721 (N_44721,N_43750,N_43676);
xor U44722 (N_44722,N_43255,N_43170);
nor U44723 (N_44723,N_43334,N_43572);
and U44724 (N_44724,N_43888,N_43452);
nand U44725 (N_44725,N_43970,N_43043);
or U44726 (N_44726,N_43639,N_43958);
or U44727 (N_44727,N_43906,N_43493);
or U44728 (N_44728,N_43465,N_43105);
xnor U44729 (N_44729,N_43421,N_43321);
nor U44730 (N_44730,N_43914,N_43681);
or U44731 (N_44731,N_43757,N_43730);
or U44732 (N_44732,N_43734,N_43158);
and U44733 (N_44733,N_43415,N_43266);
or U44734 (N_44734,N_43257,N_43591);
or U44735 (N_44735,N_43275,N_43286);
xor U44736 (N_44736,N_43790,N_43358);
and U44737 (N_44737,N_43008,N_43107);
nor U44738 (N_44738,N_43748,N_43003);
xor U44739 (N_44739,N_43307,N_43599);
nand U44740 (N_44740,N_43102,N_43048);
and U44741 (N_44741,N_43046,N_43793);
and U44742 (N_44742,N_43037,N_43197);
or U44743 (N_44743,N_43768,N_43917);
or U44744 (N_44744,N_43198,N_43313);
nand U44745 (N_44745,N_43686,N_43613);
xor U44746 (N_44746,N_43163,N_43917);
nor U44747 (N_44747,N_43283,N_43961);
and U44748 (N_44748,N_43186,N_43476);
nand U44749 (N_44749,N_43339,N_43083);
and U44750 (N_44750,N_43255,N_43999);
xnor U44751 (N_44751,N_43742,N_43824);
nand U44752 (N_44752,N_43634,N_43824);
nand U44753 (N_44753,N_43423,N_43453);
nand U44754 (N_44754,N_43607,N_43446);
nor U44755 (N_44755,N_43076,N_43894);
xor U44756 (N_44756,N_43297,N_43058);
nor U44757 (N_44757,N_43531,N_43813);
xor U44758 (N_44758,N_43979,N_43624);
nand U44759 (N_44759,N_43775,N_43686);
xor U44760 (N_44760,N_43462,N_43221);
nand U44761 (N_44761,N_43212,N_43768);
xor U44762 (N_44762,N_43502,N_43451);
or U44763 (N_44763,N_43981,N_43917);
and U44764 (N_44764,N_43149,N_43716);
or U44765 (N_44765,N_43123,N_43557);
or U44766 (N_44766,N_43539,N_43590);
nor U44767 (N_44767,N_43332,N_43936);
and U44768 (N_44768,N_43572,N_43493);
or U44769 (N_44769,N_43368,N_43892);
nand U44770 (N_44770,N_43750,N_43179);
nor U44771 (N_44771,N_43522,N_43425);
and U44772 (N_44772,N_43032,N_43789);
or U44773 (N_44773,N_43627,N_43912);
or U44774 (N_44774,N_43709,N_43668);
xnor U44775 (N_44775,N_43303,N_43131);
or U44776 (N_44776,N_43366,N_43325);
and U44777 (N_44777,N_43258,N_43677);
nor U44778 (N_44778,N_43981,N_43777);
and U44779 (N_44779,N_43183,N_43049);
xor U44780 (N_44780,N_43838,N_43531);
nand U44781 (N_44781,N_43101,N_43380);
nand U44782 (N_44782,N_43079,N_43453);
nand U44783 (N_44783,N_43917,N_43640);
nor U44784 (N_44784,N_43743,N_43470);
or U44785 (N_44785,N_43561,N_43458);
nor U44786 (N_44786,N_43246,N_43384);
or U44787 (N_44787,N_43938,N_43890);
and U44788 (N_44788,N_43209,N_43680);
and U44789 (N_44789,N_43650,N_43316);
nand U44790 (N_44790,N_43271,N_43623);
and U44791 (N_44791,N_43708,N_43057);
or U44792 (N_44792,N_43587,N_43009);
and U44793 (N_44793,N_43247,N_43383);
and U44794 (N_44794,N_43532,N_43006);
xnor U44795 (N_44795,N_43732,N_43359);
nand U44796 (N_44796,N_43442,N_43037);
nor U44797 (N_44797,N_43273,N_43862);
or U44798 (N_44798,N_43073,N_43580);
and U44799 (N_44799,N_43252,N_43964);
xnor U44800 (N_44800,N_43163,N_43249);
nand U44801 (N_44801,N_43332,N_43629);
xor U44802 (N_44802,N_43701,N_43080);
nand U44803 (N_44803,N_43640,N_43044);
nand U44804 (N_44804,N_43922,N_43275);
nor U44805 (N_44805,N_43437,N_43347);
or U44806 (N_44806,N_43087,N_43966);
nand U44807 (N_44807,N_43783,N_43407);
and U44808 (N_44808,N_43429,N_43564);
xnor U44809 (N_44809,N_43806,N_43025);
nand U44810 (N_44810,N_43042,N_43358);
nor U44811 (N_44811,N_43825,N_43053);
and U44812 (N_44812,N_43166,N_43889);
or U44813 (N_44813,N_43671,N_43693);
nand U44814 (N_44814,N_43798,N_43706);
xor U44815 (N_44815,N_43789,N_43463);
xor U44816 (N_44816,N_43072,N_43796);
or U44817 (N_44817,N_43348,N_43430);
xnor U44818 (N_44818,N_43008,N_43576);
and U44819 (N_44819,N_43282,N_43213);
or U44820 (N_44820,N_43768,N_43276);
or U44821 (N_44821,N_43914,N_43236);
nand U44822 (N_44822,N_43189,N_43703);
xor U44823 (N_44823,N_43317,N_43248);
nor U44824 (N_44824,N_43961,N_43139);
and U44825 (N_44825,N_43077,N_43028);
nor U44826 (N_44826,N_43883,N_43982);
nor U44827 (N_44827,N_43418,N_43495);
nand U44828 (N_44828,N_43345,N_43907);
xnor U44829 (N_44829,N_43774,N_43656);
nor U44830 (N_44830,N_43186,N_43767);
xor U44831 (N_44831,N_43885,N_43738);
nand U44832 (N_44832,N_43563,N_43091);
xor U44833 (N_44833,N_43035,N_43769);
xor U44834 (N_44834,N_43305,N_43416);
nor U44835 (N_44835,N_43812,N_43864);
nor U44836 (N_44836,N_43485,N_43606);
and U44837 (N_44837,N_43027,N_43870);
nor U44838 (N_44838,N_43657,N_43926);
nor U44839 (N_44839,N_43311,N_43576);
nor U44840 (N_44840,N_43883,N_43656);
or U44841 (N_44841,N_43122,N_43775);
xor U44842 (N_44842,N_43823,N_43610);
xor U44843 (N_44843,N_43176,N_43484);
nor U44844 (N_44844,N_43864,N_43476);
nor U44845 (N_44845,N_43445,N_43455);
or U44846 (N_44846,N_43015,N_43823);
nand U44847 (N_44847,N_43737,N_43676);
xnor U44848 (N_44848,N_43072,N_43572);
nor U44849 (N_44849,N_43388,N_43495);
xor U44850 (N_44850,N_43247,N_43733);
or U44851 (N_44851,N_43530,N_43347);
nor U44852 (N_44852,N_43013,N_43155);
and U44853 (N_44853,N_43419,N_43395);
nand U44854 (N_44854,N_43482,N_43144);
and U44855 (N_44855,N_43802,N_43541);
xnor U44856 (N_44856,N_43353,N_43328);
and U44857 (N_44857,N_43914,N_43219);
nand U44858 (N_44858,N_43368,N_43009);
xor U44859 (N_44859,N_43575,N_43794);
nor U44860 (N_44860,N_43292,N_43978);
nor U44861 (N_44861,N_43599,N_43948);
or U44862 (N_44862,N_43243,N_43672);
or U44863 (N_44863,N_43939,N_43593);
xor U44864 (N_44864,N_43085,N_43729);
and U44865 (N_44865,N_43715,N_43375);
nor U44866 (N_44866,N_43240,N_43075);
or U44867 (N_44867,N_43247,N_43081);
nand U44868 (N_44868,N_43050,N_43838);
xor U44869 (N_44869,N_43774,N_43252);
nand U44870 (N_44870,N_43693,N_43512);
or U44871 (N_44871,N_43287,N_43721);
and U44872 (N_44872,N_43293,N_43899);
and U44873 (N_44873,N_43884,N_43822);
nand U44874 (N_44874,N_43697,N_43225);
nor U44875 (N_44875,N_43648,N_43588);
nand U44876 (N_44876,N_43678,N_43823);
or U44877 (N_44877,N_43358,N_43078);
or U44878 (N_44878,N_43159,N_43551);
or U44879 (N_44879,N_43354,N_43737);
nor U44880 (N_44880,N_43520,N_43228);
xnor U44881 (N_44881,N_43494,N_43608);
nand U44882 (N_44882,N_43834,N_43706);
xnor U44883 (N_44883,N_43980,N_43419);
nor U44884 (N_44884,N_43505,N_43348);
nand U44885 (N_44885,N_43955,N_43125);
and U44886 (N_44886,N_43473,N_43226);
xor U44887 (N_44887,N_43195,N_43855);
nand U44888 (N_44888,N_43272,N_43772);
and U44889 (N_44889,N_43457,N_43272);
nor U44890 (N_44890,N_43068,N_43702);
or U44891 (N_44891,N_43477,N_43032);
xor U44892 (N_44892,N_43859,N_43833);
nor U44893 (N_44893,N_43226,N_43327);
nor U44894 (N_44894,N_43131,N_43670);
and U44895 (N_44895,N_43668,N_43356);
or U44896 (N_44896,N_43361,N_43082);
xnor U44897 (N_44897,N_43087,N_43523);
and U44898 (N_44898,N_43781,N_43462);
or U44899 (N_44899,N_43730,N_43921);
and U44900 (N_44900,N_43508,N_43295);
and U44901 (N_44901,N_43086,N_43031);
and U44902 (N_44902,N_43552,N_43859);
xnor U44903 (N_44903,N_43716,N_43399);
nor U44904 (N_44904,N_43444,N_43437);
and U44905 (N_44905,N_43696,N_43608);
and U44906 (N_44906,N_43402,N_43211);
and U44907 (N_44907,N_43228,N_43215);
nor U44908 (N_44908,N_43754,N_43896);
xor U44909 (N_44909,N_43978,N_43618);
nor U44910 (N_44910,N_43482,N_43892);
or U44911 (N_44911,N_43012,N_43019);
and U44912 (N_44912,N_43339,N_43004);
or U44913 (N_44913,N_43990,N_43662);
and U44914 (N_44914,N_43143,N_43564);
nand U44915 (N_44915,N_43997,N_43876);
and U44916 (N_44916,N_43447,N_43203);
or U44917 (N_44917,N_43909,N_43436);
nand U44918 (N_44918,N_43499,N_43422);
and U44919 (N_44919,N_43699,N_43315);
nand U44920 (N_44920,N_43487,N_43241);
nor U44921 (N_44921,N_43510,N_43927);
and U44922 (N_44922,N_43348,N_43453);
xor U44923 (N_44923,N_43500,N_43825);
nand U44924 (N_44924,N_43477,N_43022);
nand U44925 (N_44925,N_43696,N_43906);
or U44926 (N_44926,N_43437,N_43083);
nor U44927 (N_44927,N_43971,N_43567);
or U44928 (N_44928,N_43581,N_43623);
nand U44929 (N_44929,N_43380,N_43060);
and U44930 (N_44930,N_43473,N_43117);
nand U44931 (N_44931,N_43318,N_43548);
xnor U44932 (N_44932,N_43860,N_43068);
and U44933 (N_44933,N_43604,N_43208);
xor U44934 (N_44934,N_43457,N_43899);
xnor U44935 (N_44935,N_43746,N_43349);
xnor U44936 (N_44936,N_43263,N_43817);
nor U44937 (N_44937,N_43023,N_43956);
and U44938 (N_44938,N_43784,N_43638);
nand U44939 (N_44939,N_43209,N_43190);
nor U44940 (N_44940,N_43678,N_43918);
nand U44941 (N_44941,N_43512,N_43986);
and U44942 (N_44942,N_43508,N_43043);
or U44943 (N_44943,N_43810,N_43314);
and U44944 (N_44944,N_43891,N_43155);
and U44945 (N_44945,N_43065,N_43058);
xnor U44946 (N_44946,N_43905,N_43731);
and U44947 (N_44947,N_43921,N_43607);
and U44948 (N_44948,N_43283,N_43050);
and U44949 (N_44949,N_43305,N_43481);
and U44950 (N_44950,N_43376,N_43516);
xnor U44951 (N_44951,N_43525,N_43819);
or U44952 (N_44952,N_43478,N_43966);
xnor U44953 (N_44953,N_43886,N_43414);
nand U44954 (N_44954,N_43757,N_43756);
xnor U44955 (N_44955,N_43196,N_43510);
nand U44956 (N_44956,N_43898,N_43700);
and U44957 (N_44957,N_43479,N_43371);
or U44958 (N_44958,N_43390,N_43282);
xor U44959 (N_44959,N_43308,N_43400);
xnor U44960 (N_44960,N_43753,N_43470);
xor U44961 (N_44961,N_43240,N_43531);
and U44962 (N_44962,N_43282,N_43830);
xnor U44963 (N_44963,N_43570,N_43497);
and U44964 (N_44964,N_43901,N_43682);
nand U44965 (N_44965,N_43642,N_43355);
nand U44966 (N_44966,N_43279,N_43179);
or U44967 (N_44967,N_43090,N_43930);
and U44968 (N_44968,N_43232,N_43961);
xnor U44969 (N_44969,N_43127,N_43659);
and U44970 (N_44970,N_43151,N_43195);
xnor U44971 (N_44971,N_43225,N_43065);
and U44972 (N_44972,N_43069,N_43199);
or U44973 (N_44973,N_43859,N_43043);
nor U44974 (N_44974,N_43527,N_43180);
or U44975 (N_44975,N_43920,N_43842);
nand U44976 (N_44976,N_43952,N_43638);
xnor U44977 (N_44977,N_43790,N_43935);
nand U44978 (N_44978,N_43518,N_43929);
nand U44979 (N_44979,N_43691,N_43124);
xnor U44980 (N_44980,N_43376,N_43897);
nand U44981 (N_44981,N_43588,N_43405);
or U44982 (N_44982,N_43028,N_43661);
nor U44983 (N_44983,N_43485,N_43438);
nor U44984 (N_44984,N_43780,N_43961);
nand U44985 (N_44985,N_43080,N_43280);
xnor U44986 (N_44986,N_43299,N_43363);
nor U44987 (N_44987,N_43438,N_43974);
and U44988 (N_44988,N_43947,N_43644);
xnor U44989 (N_44989,N_43472,N_43064);
nand U44990 (N_44990,N_43528,N_43856);
and U44991 (N_44991,N_43644,N_43938);
and U44992 (N_44992,N_43313,N_43972);
and U44993 (N_44993,N_43077,N_43989);
and U44994 (N_44994,N_43452,N_43388);
and U44995 (N_44995,N_43973,N_43283);
xor U44996 (N_44996,N_43952,N_43850);
and U44997 (N_44997,N_43505,N_43447);
nand U44998 (N_44998,N_43353,N_43396);
xor U44999 (N_44999,N_43141,N_43164);
and U45000 (N_45000,N_44997,N_44460);
nand U45001 (N_45001,N_44746,N_44233);
xnor U45002 (N_45002,N_44383,N_44718);
or U45003 (N_45003,N_44815,N_44712);
and U45004 (N_45004,N_44584,N_44222);
and U45005 (N_45005,N_44881,N_44902);
or U45006 (N_45006,N_44887,N_44281);
and U45007 (N_45007,N_44094,N_44347);
and U45008 (N_45008,N_44249,N_44948);
xor U45009 (N_45009,N_44111,N_44609);
and U45010 (N_45010,N_44365,N_44106);
nand U45011 (N_45011,N_44015,N_44100);
and U45012 (N_45012,N_44357,N_44433);
nand U45013 (N_45013,N_44048,N_44481);
or U45014 (N_45014,N_44361,N_44827);
and U45015 (N_45015,N_44499,N_44127);
or U45016 (N_45016,N_44781,N_44714);
or U45017 (N_45017,N_44445,N_44080);
nor U45018 (N_45018,N_44913,N_44770);
nor U45019 (N_45019,N_44364,N_44400);
xnor U45020 (N_45020,N_44920,N_44469);
xnor U45021 (N_45021,N_44856,N_44638);
nand U45022 (N_45022,N_44200,N_44651);
and U45023 (N_45023,N_44268,N_44497);
or U45024 (N_45024,N_44672,N_44244);
or U45025 (N_45025,N_44680,N_44483);
nor U45026 (N_45026,N_44424,N_44501);
xnor U45027 (N_45027,N_44141,N_44387);
or U45028 (N_45028,N_44086,N_44337);
or U45029 (N_45029,N_44318,N_44510);
or U45030 (N_45030,N_44555,N_44980);
and U45031 (N_45031,N_44486,N_44264);
xor U45032 (N_45032,N_44967,N_44076);
xor U45033 (N_45033,N_44284,N_44208);
nand U45034 (N_45034,N_44403,N_44182);
nand U45035 (N_45035,N_44704,N_44578);
nor U45036 (N_45036,N_44265,N_44198);
nand U45037 (N_45037,N_44346,N_44761);
and U45038 (N_45038,N_44049,N_44278);
and U45039 (N_45039,N_44331,N_44126);
or U45040 (N_45040,N_44861,N_44294);
xnor U45041 (N_45041,N_44426,N_44889);
and U45042 (N_45042,N_44814,N_44969);
and U45043 (N_45043,N_44267,N_44779);
nor U45044 (N_45044,N_44479,N_44930);
xor U45045 (N_45045,N_44175,N_44859);
xor U45046 (N_45046,N_44062,N_44464);
xor U45047 (N_45047,N_44514,N_44994);
and U45048 (N_45048,N_44134,N_44971);
nand U45049 (N_45049,N_44248,N_44467);
nand U45050 (N_45050,N_44791,N_44897);
or U45051 (N_45051,N_44275,N_44984);
nor U45052 (N_45052,N_44298,N_44652);
or U45053 (N_45053,N_44676,N_44325);
nand U45054 (N_45054,N_44288,N_44345);
nor U45055 (N_45055,N_44798,N_44098);
nand U45056 (N_45056,N_44922,N_44561);
and U45057 (N_45057,N_44556,N_44334);
nor U45058 (N_45058,N_44031,N_44371);
or U45059 (N_45059,N_44420,N_44181);
xnor U45060 (N_45060,N_44719,N_44549);
and U45061 (N_45061,N_44137,N_44941);
and U45062 (N_45062,N_44225,N_44104);
nor U45063 (N_45063,N_44805,N_44545);
or U45064 (N_45064,N_44604,N_44522);
and U45065 (N_45065,N_44505,N_44133);
and U45066 (N_45066,N_44614,N_44115);
or U45067 (N_45067,N_44550,N_44147);
nor U45068 (N_45068,N_44576,N_44860);
or U45069 (N_45069,N_44670,N_44329);
nor U45070 (N_45070,N_44165,N_44730);
and U45071 (N_45071,N_44257,N_44053);
nor U45072 (N_45072,N_44579,N_44091);
or U45073 (N_45073,N_44903,N_44082);
and U45074 (N_45074,N_44146,N_44663);
or U45075 (N_45075,N_44794,N_44707);
and U45076 (N_45076,N_44241,N_44051);
xor U45077 (N_45077,N_44946,N_44336);
and U45078 (N_45078,N_44456,N_44187);
nand U45079 (N_45079,N_44837,N_44066);
nand U45080 (N_45080,N_44709,N_44037);
or U45081 (N_45081,N_44532,N_44145);
nor U45082 (N_45082,N_44885,N_44523);
or U45083 (N_45083,N_44963,N_44940);
nor U45084 (N_45084,N_44724,N_44934);
nor U45085 (N_45085,N_44942,N_44711);
nand U45086 (N_45086,N_44769,N_44011);
xor U45087 (N_45087,N_44759,N_44074);
nor U45088 (N_45088,N_44723,N_44368);
nor U45089 (N_45089,N_44277,N_44119);
nor U45090 (N_45090,N_44192,N_44435);
and U45091 (N_45091,N_44698,N_44312);
or U45092 (N_45092,N_44907,N_44362);
or U45093 (N_45093,N_44485,N_44418);
xor U45094 (N_45094,N_44664,N_44880);
or U45095 (N_45095,N_44321,N_44517);
and U45096 (N_45096,N_44454,N_44474);
or U45097 (N_45097,N_44307,N_44964);
and U45098 (N_45098,N_44995,N_44434);
and U45099 (N_45099,N_44219,N_44909);
nand U45100 (N_45100,N_44637,N_44436);
nand U45101 (N_45101,N_44201,N_44702);
nor U45102 (N_45102,N_44188,N_44810);
or U45103 (N_45103,N_44197,N_44996);
or U45104 (N_45104,N_44527,N_44973);
nand U45105 (N_45105,N_44087,N_44605);
or U45106 (N_45106,N_44045,N_44531);
xor U45107 (N_45107,N_44694,N_44229);
or U45108 (N_45108,N_44461,N_44720);
nand U45109 (N_45109,N_44613,N_44804);
nor U45110 (N_45110,N_44957,N_44109);
and U45111 (N_45111,N_44803,N_44121);
and U45112 (N_45112,N_44540,N_44910);
xor U45113 (N_45113,N_44819,N_44220);
xnor U45114 (N_45114,N_44758,N_44577);
xnor U45115 (N_45115,N_44895,N_44826);
xnor U45116 (N_45116,N_44841,N_44239);
nor U45117 (N_45117,N_44754,N_44245);
nor U45118 (N_45118,N_44449,N_44713);
and U45119 (N_45119,N_44982,N_44524);
xor U45120 (N_45120,N_44085,N_44904);
or U45121 (N_45121,N_44872,N_44726);
xnor U45122 (N_45122,N_44040,N_44833);
and U45123 (N_45123,N_44925,N_44283);
xnor U45124 (N_45124,N_44390,N_44618);
and U45125 (N_45125,N_44731,N_44752);
or U45126 (N_45126,N_44046,N_44343);
or U45127 (N_45127,N_44915,N_44866);
and U45128 (N_45128,N_44828,N_44102);
or U45129 (N_45129,N_44839,N_44843);
nor U45130 (N_45130,N_44742,N_44305);
nand U45131 (N_45131,N_44060,N_44039);
nand U45132 (N_45132,N_44128,N_44835);
and U45133 (N_45133,N_44666,N_44322);
nor U45134 (N_45134,N_44554,N_44447);
xnor U45135 (N_45135,N_44263,N_44246);
and U45136 (N_45136,N_44630,N_44675);
nand U45137 (N_45137,N_44627,N_44097);
nor U45138 (N_45138,N_44050,N_44956);
or U45139 (N_45139,N_44430,N_44189);
nor U45140 (N_45140,N_44944,N_44689);
nor U45141 (N_45141,N_44162,N_44071);
nand U45142 (N_45142,N_44582,N_44224);
and U45143 (N_45143,N_44854,N_44206);
and U45144 (N_45144,N_44533,N_44421);
xor U45145 (N_45145,N_44251,N_44685);
nand U45146 (N_45146,N_44414,N_44802);
nand U45147 (N_45147,N_44632,N_44480);
nand U45148 (N_45148,N_44848,N_44811);
or U45149 (N_45149,N_44767,N_44033);
nor U45150 (N_45150,N_44475,N_44542);
and U45151 (N_45151,N_44906,N_44335);
nor U45152 (N_45152,N_44161,N_44772);
or U45153 (N_45153,N_44844,N_44491);
and U45154 (N_45154,N_44358,N_44306);
nor U45155 (N_45155,N_44732,N_44124);
and U45156 (N_45156,N_44110,N_44615);
and U45157 (N_45157,N_44693,N_44196);
and U45158 (N_45158,N_44393,N_44027);
or U45159 (N_45159,N_44455,N_44255);
xor U45160 (N_45160,N_44961,N_44093);
nand U45161 (N_45161,N_44324,N_44417);
nor U45162 (N_45162,N_44226,N_44747);
and U45163 (N_45163,N_44933,N_44007);
nor U45164 (N_45164,N_44657,N_44478);
and U45165 (N_45165,N_44945,N_44620);
xnor U45166 (N_45166,N_44800,N_44653);
and U45167 (N_45167,N_44047,N_44825);
or U45168 (N_45168,N_44507,N_44728);
xnor U45169 (N_45169,N_44431,N_44024);
and U45170 (N_45170,N_44450,N_44308);
nand U45171 (N_45171,N_44349,N_44061);
nand U45172 (N_45172,N_44309,N_44156);
or U45173 (N_45173,N_44799,N_44112);
nand U45174 (N_45174,N_44649,N_44778);
xor U45175 (N_45175,N_44587,N_44935);
nand U45176 (N_45176,N_44882,N_44429);
nor U45177 (N_45177,N_44869,N_44338);
or U45178 (N_45178,N_44564,N_44697);
nand U45179 (N_45179,N_44428,N_44612);
and U45180 (N_45180,N_44590,N_44459);
or U45181 (N_45181,N_44375,N_44842);
and U45182 (N_45182,N_44737,N_44269);
xnor U45183 (N_45183,N_44557,N_44059);
nor U45184 (N_45184,N_44817,N_44397);
nand U45185 (N_45185,N_44955,N_44008);
and U45186 (N_45186,N_44003,N_44727);
xnor U45187 (N_45187,N_44378,N_44760);
nor U45188 (N_45188,N_44144,N_44756);
and U45189 (N_45189,N_44568,N_44927);
nand U45190 (N_45190,N_44316,N_44359);
or U45191 (N_45191,N_44688,N_44487);
nand U45192 (N_45192,N_44256,N_44422);
and U45193 (N_45193,N_44589,N_44153);
and U45194 (N_45194,N_44541,N_44068);
nand U45195 (N_45195,N_44072,N_44502);
or U45196 (N_45196,N_44928,N_44315);
xor U45197 (N_45197,N_44721,N_44809);
or U45198 (N_45198,N_44979,N_44660);
nor U45199 (N_45199,N_44865,N_44089);
nand U45200 (N_45200,N_44512,N_44936);
or U45201 (N_45201,N_44290,N_44640);
nand U45202 (N_45202,N_44585,N_44395);
nor U45203 (N_45203,N_44125,N_44656);
or U45204 (N_45204,N_44981,N_44559);
nand U45205 (N_45205,N_44706,N_44212);
nor U45206 (N_45206,N_44855,N_44914);
nand U45207 (N_45207,N_44782,N_44753);
xor U45208 (N_45208,N_44939,N_44287);
and U45209 (N_45209,N_44509,N_44539);
nor U45210 (N_45210,N_44734,N_44634);
nand U45211 (N_45211,N_44621,N_44836);
nor U45212 (N_45212,N_44818,N_44427);
xor U45213 (N_45213,N_44966,N_44506);
xor U45214 (N_45214,N_44820,N_44525);
xor U45215 (N_45215,N_44178,N_44518);
xor U45216 (N_45216,N_44641,N_44551);
and U45217 (N_45217,N_44235,N_44304);
nand U45218 (N_45218,N_44372,N_44873);
or U45219 (N_45219,N_44311,N_44138);
or U45220 (N_45220,N_44477,N_44254);
and U45221 (N_45221,N_44195,N_44566);
xnor U45222 (N_45222,N_44784,N_44291);
and U45223 (N_45223,N_44991,N_44847);
nand U45224 (N_45224,N_44838,N_44056);
and U45225 (N_45225,N_44622,N_44592);
or U45226 (N_45226,N_44215,N_44270);
and U45227 (N_45227,N_44296,N_44139);
nor U45228 (N_45228,N_44645,N_44004);
and U45229 (N_45229,N_44292,N_44367);
or U45230 (N_45230,N_44647,N_44705);
nor U45231 (N_45231,N_44684,N_44157);
and U45232 (N_45232,N_44896,N_44776);
or U45233 (N_45233,N_44073,N_44191);
and U45234 (N_45234,N_44992,N_44888);
xnor U45235 (N_45235,N_44667,N_44691);
and U45236 (N_45236,N_44136,N_44924);
and U45237 (N_45237,N_44238,N_44832);
nor U45238 (N_45238,N_44735,N_44105);
xnor U45239 (N_45239,N_44028,N_44293);
or U45240 (N_45240,N_44503,N_44333);
nor U45241 (N_45241,N_44999,N_44870);
nand U45242 (N_45242,N_44905,N_44923);
nand U45243 (N_45243,N_44926,N_44314);
nor U45244 (N_45244,N_44415,N_44526);
xor U45245 (N_45245,N_44849,N_44912);
and U45246 (N_45246,N_44030,N_44356);
xnor U45247 (N_45247,N_44065,N_44001);
xor U45248 (N_45248,N_44552,N_44588);
nand U45249 (N_45249,N_44179,N_44699);
or U45250 (N_45250,N_44247,N_44376);
nor U45251 (N_45251,N_44987,N_44968);
nor U45252 (N_45252,N_44567,N_44813);
or U45253 (N_45253,N_44757,N_44272);
or U45254 (N_45254,N_44583,N_44214);
xnor U45255 (N_45255,N_44710,N_44722);
or U45256 (N_45256,N_44608,N_44029);
and U45257 (N_45257,N_44044,N_44185);
nor U45258 (N_45258,N_44052,N_44026);
or U45259 (N_45259,N_44690,N_44107);
and U45260 (N_45260,N_44686,N_44570);
nand U45261 (N_45261,N_44890,N_44186);
or U45262 (N_45262,N_44317,N_44299);
nor U45263 (N_45263,N_44831,N_44862);
nand U45264 (N_45264,N_44412,N_44016);
and U45265 (N_45265,N_44611,N_44899);
and U45266 (N_45266,N_44673,N_44452);
nor U45267 (N_45267,N_44681,N_44183);
nor U45268 (N_45268,N_44389,N_44227);
nor U45269 (N_45269,N_44339,N_44626);
and U45270 (N_45270,N_44406,N_44687);
and U45271 (N_45271,N_44374,N_44801);
or U45272 (N_45272,N_44210,N_44211);
or U45273 (N_45273,N_44565,N_44385);
xor U45274 (N_45274,N_44332,N_44571);
nand U45275 (N_45275,N_44425,N_44009);
and U45276 (N_45276,N_44300,N_44750);
and U45277 (N_45277,N_44413,N_44432);
xor U45278 (N_45278,N_44642,N_44289);
and U45279 (N_45279,N_44000,N_44853);
or U45280 (N_45280,N_44745,N_44633);
and U45281 (N_45281,N_44977,N_44950);
and U45282 (N_45282,N_44092,N_44019);
or U45283 (N_45283,N_44636,N_44204);
xor U45284 (N_45284,N_44038,N_44352);
and U45285 (N_45285,N_44232,N_44768);
or U45286 (N_45286,N_44142,N_44373);
nand U45287 (N_45287,N_44863,N_44949);
nand U45288 (N_45288,N_44310,N_44118);
nand U45289 (N_45289,N_44993,N_44603);
nor U45290 (N_45290,N_44736,N_44190);
nand U45291 (N_45291,N_44473,N_44279);
nor U45292 (N_45292,N_44598,N_44840);
and U45293 (N_45293,N_44205,N_44678);
and U45294 (N_45294,N_44569,N_44851);
xnor U45295 (N_45295,N_44738,N_44492);
nor U45296 (N_45296,N_44682,N_44323);
nand U45297 (N_45297,N_44610,N_44807);
or U45298 (N_45298,N_44398,N_44563);
nor U45299 (N_45299,N_44005,N_44261);
or U45300 (N_45300,N_44574,N_44231);
nand U45301 (N_45301,N_44797,N_44273);
nand U45302 (N_45302,N_44488,N_44380);
xnor U45303 (N_45303,N_44871,N_44320);
xor U45304 (N_45304,N_44386,N_44536);
nand U45305 (N_45305,N_44116,N_44143);
nor U45306 (N_45306,N_44845,N_44160);
nor U45307 (N_45307,N_44063,N_44500);
xnor U45308 (N_45308,N_44017,N_44864);
xor U45309 (N_45309,N_44780,N_44703);
nand U45310 (N_45310,N_44444,N_44643);
and U45311 (N_45311,N_44654,N_44276);
or U45312 (N_45312,N_44282,N_44965);
xor U45313 (N_45313,N_44164,N_44103);
nand U45314 (N_45314,N_44765,N_44985);
nand U45315 (N_45315,N_44974,N_44867);
nor U45316 (N_45316,N_44058,N_44593);
or U45317 (N_45317,N_44792,N_44023);
nand U45318 (N_45318,N_44891,N_44465);
xor U45319 (N_45319,N_44295,N_44408);
nand U45320 (N_45320,N_44919,N_44528);
and U45321 (N_45321,N_44983,N_44504);
nand U45322 (N_45322,N_44490,N_44602);
and U45323 (N_45323,N_44020,N_44534);
and U45324 (N_45324,N_44596,N_44113);
xnor U45325 (N_45325,N_44580,N_44874);
and U45326 (N_45326,N_44237,N_44679);
or U45327 (N_45327,N_44476,N_44823);
or U45328 (N_45328,N_44619,N_44057);
nand U45329 (N_45329,N_44716,N_44537);
nand U45330 (N_45330,N_44242,N_44631);
nor U45331 (N_45331,N_44771,N_44516);
xor U45332 (N_45332,N_44440,N_44929);
nor U45333 (N_45333,N_44377,N_44055);
nor U45334 (N_45334,N_44744,N_44482);
nor U45335 (N_45335,N_44101,N_44508);
nor U45336 (N_45336,N_44898,N_44159);
or U45337 (N_45337,N_44472,N_44793);
nand U45338 (N_45338,N_44351,N_44850);
xor U45339 (N_45339,N_44259,N_44193);
or U45340 (N_45340,N_44457,N_44370);
nor U45341 (N_45341,N_44174,N_44096);
nand U45342 (N_45342,N_44354,N_44083);
nand U45343 (N_45343,N_44658,N_44171);
nor U45344 (N_45344,N_44821,N_44606);
xnor U45345 (N_45345,N_44886,N_44013);
nand U45346 (N_45346,N_44830,N_44280);
or U45347 (N_45347,N_44313,N_44253);
or U45348 (N_45348,N_44700,N_44150);
or U45349 (N_45349,N_44773,N_44366);
nand U45350 (N_45350,N_44749,N_44668);
xor U45351 (N_45351,N_44513,N_44169);
nor U45352 (N_45352,N_44441,N_44496);
or U45353 (N_45353,N_44018,N_44976);
xor U45354 (N_45354,N_44022,N_44725);
nand U45355 (N_45355,N_44054,N_44947);
nand U45356 (N_45356,N_44117,N_44879);
or U45357 (N_45357,N_44132,N_44209);
xor U45358 (N_45358,N_44410,N_44808);
nor U45359 (N_45359,N_44327,N_44893);
xor U45360 (N_45360,N_44152,N_44547);
xor U45361 (N_45361,N_44114,N_44035);
and U45362 (N_45362,N_44741,N_44494);
xor U45363 (N_45363,N_44399,N_44766);
xnor U45364 (N_45364,N_44795,N_44868);
nor U45365 (N_45365,N_44597,N_44230);
and U45366 (N_45366,N_44070,N_44755);
nand U45367 (N_45367,N_44529,N_44095);
xnor U45368 (N_45368,N_44172,N_44203);
xnor U45369 (N_45369,N_44774,N_44916);
and U45370 (N_45370,N_44671,N_44543);
xnor U45371 (N_45371,N_44123,N_44489);
xnor U45372 (N_45372,N_44646,N_44151);
and U45373 (N_45373,N_44519,N_44648);
and U45374 (N_45374,N_44025,N_44404);
and U45375 (N_45375,N_44363,N_44546);
or U45376 (N_45376,N_44443,N_44986);
nand U45377 (N_45377,N_44355,N_44786);
xnor U45378 (N_45378,N_44184,N_44701);
nor U45379 (N_45379,N_44900,N_44350);
and U45380 (N_45380,N_44901,N_44846);
and U45381 (N_45381,N_44069,N_44975);
or U45382 (N_45382,N_44170,N_44453);
nand U45383 (N_45383,N_44562,N_44884);
nor U45384 (N_45384,N_44908,N_44129);
nor U45385 (N_45385,N_44341,N_44135);
xnor U45386 (N_45386,N_44498,N_44423);
and U45387 (N_45387,N_44154,N_44953);
xor U45388 (N_45388,N_44829,N_44034);
and U45389 (N_45389,N_44243,N_44140);
nand U45390 (N_45390,N_44990,N_44852);
nor U45391 (N_45391,N_44194,N_44493);
or U45392 (N_45392,N_44696,N_44108);
xor U45393 (N_45393,N_44409,N_44623);
or U45394 (N_45394,N_44442,N_44931);
or U45395 (N_45395,N_44388,N_44739);
xnor U45396 (N_45396,N_44495,N_44834);
nand U45397 (N_45397,N_44816,N_44067);
and U45398 (N_45398,N_44674,N_44553);
or U45399 (N_45399,N_44439,N_44624);
xnor U45400 (N_45400,N_44591,N_44382);
or U45401 (N_45401,N_44575,N_44548);
or U45402 (N_45402,N_44883,N_44616);
and U45403 (N_45403,N_44748,N_44733);
nand U45404 (N_45404,N_44344,N_44163);
or U45405 (N_45405,N_44328,N_44790);
nor U45406 (N_45406,N_44348,N_44951);
nand U45407 (N_45407,N_44607,N_44360);
or U45408 (N_45408,N_44777,N_44216);
nor U45409 (N_45409,N_44451,N_44075);
xor U45410 (N_45410,N_44462,N_44695);
nor U45411 (N_45411,N_44659,N_44260);
nand U45412 (N_45412,N_44878,N_44471);
or U45413 (N_45413,N_44391,N_44099);
nand U45414 (N_45414,N_44952,N_44958);
nor U45415 (N_45415,N_44402,N_44405);
nor U45416 (N_45416,N_44635,N_44202);
nand U45417 (N_45417,N_44988,N_44297);
xor U45418 (N_45418,N_44876,N_44970);
xor U45419 (N_45419,N_44010,N_44463);
xor U45420 (N_45420,N_44708,N_44286);
and U45421 (N_45421,N_44396,N_44644);
xor U45422 (N_45422,N_44665,N_44894);
or U45423 (N_45423,N_44599,N_44892);
xor U45424 (N_45424,N_44081,N_44628);
nor U45425 (N_45425,N_44743,N_44381);
or U45426 (N_45426,N_44629,N_44763);
nand U45427 (N_45427,N_44573,N_44043);
nor U45428 (N_45428,N_44875,N_44252);
xnor U45429 (N_45429,N_44729,N_44662);
and U45430 (N_45430,N_44954,N_44560);
xnor U45431 (N_45431,N_44006,N_44303);
or U45432 (N_45432,N_44937,N_44617);
nand U45433 (N_45433,N_44148,N_44521);
and U45434 (N_45434,N_44921,N_44787);
nor U45435 (N_45435,N_44978,N_44715);
xor U45436 (N_45436,N_44600,N_44032);
and U45437 (N_45437,N_44824,N_44207);
nand U45438 (N_45438,N_44812,N_44079);
and U45439 (N_45439,N_44088,N_44581);
xnor U45440 (N_45440,N_44213,N_44236);
and U45441 (N_45441,N_44319,N_44661);
nor U45442 (N_45442,N_44595,N_44470);
nor U45443 (N_45443,N_44692,N_44601);
or U45444 (N_45444,N_44960,N_44911);
nor U45445 (N_45445,N_44064,N_44535);
nand U45446 (N_45446,N_44989,N_44938);
nor U45447 (N_45447,N_44130,N_44530);
and U45448 (N_45448,N_44639,N_44458);
and U45449 (N_45449,N_44544,N_44234);
nand U45450 (N_45450,N_44218,N_44511);
xor U45451 (N_45451,N_44419,N_44416);
or U45452 (N_45452,N_44258,N_44586);
or U45453 (N_45453,N_44158,N_44041);
nand U45454 (N_45454,N_44669,N_44788);
and U45455 (N_45455,N_44330,N_44149);
xnor U45456 (N_45456,N_44301,N_44340);
and U45457 (N_45457,N_44655,N_44437);
nand U45458 (N_45458,N_44250,N_44783);
xor U45459 (N_45459,N_44271,N_44806);
and U45460 (N_45460,N_44036,N_44077);
nor U45461 (N_45461,N_44520,N_44572);
and U45462 (N_45462,N_44877,N_44012);
nor U45463 (N_45463,N_44084,N_44796);
nor U45464 (N_45464,N_44384,N_44468);
xor U45465 (N_45465,N_44221,N_44677);
nor U45466 (N_45466,N_44021,N_44392);
or U45467 (N_45467,N_44717,N_44262);
nor U45468 (N_45468,N_44302,N_44762);
or U45469 (N_45469,N_44764,N_44918);
nand U45470 (N_45470,N_44131,N_44625);
and U45471 (N_45471,N_44090,N_44326);
nor U45472 (N_45472,N_44167,N_44446);
or U45473 (N_45473,N_44353,N_44407);
nand U45474 (N_45474,N_44177,N_44122);
nor U45475 (N_45475,N_44173,N_44002);
and U45476 (N_45476,N_44785,N_44857);
xor U45477 (N_45477,N_44448,N_44217);
nand U45478 (N_45478,N_44155,N_44789);
nor U45479 (N_45479,N_44740,N_44285);
nand U45480 (N_45480,N_44538,N_44775);
xnor U45481 (N_45481,N_44223,N_44411);
xor U45482 (N_45482,N_44515,N_44466);
nand U45483 (N_45483,N_44166,N_44484);
nand U45484 (N_45484,N_44932,N_44228);
nand U45485 (N_45485,N_44274,N_44120);
or U45486 (N_45486,N_44401,N_44342);
and U45487 (N_45487,N_44558,N_44180);
xnor U45488 (N_45488,N_44394,N_44369);
nor U45489 (N_45489,N_44168,N_44594);
nand U45490 (N_45490,N_44379,N_44199);
or U45491 (N_45491,N_44078,N_44962);
and U45492 (N_45492,N_44650,N_44176);
nand U45493 (N_45493,N_44683,N_44943);
and U45494 (N_45494,N_44438,N_44751);
or U45495 (N_45495,N_44240,N_44858);
and U45496 (N_45496,N_44972,N_44042);
or U45497 (N_45497,N_44959,N_44014);
xnor U45498 (N_45498,N_44917,N_44998);
nand U45499 (N_45499,N_44822,N_44266);
and U45500 (N_45500,N_44470,N_44852);
nand U45501 (N_45501,N_44599,N_44948);
or U45502 (N_45502,N_44349,N_44292);
nor U45503 (N_45503,N_44386,N_44821);
xor U45504 (N_45504,N_44519,N_44558);
or U45505 (N_45505,N_44771,N_44884);
and U45506 (N_45506,N_44121,N_44194);
or U45507 (N_45507,N_44733,N_44732);
nor U45508 (N_45508,N_44503,N_44804);
xnor U45509 (N_45509,N_44934,N_44866);
xor U45510 (N_45510,N_44219,N_44338);
xnor U45511 (N_45511,N_44875,N_44787);
or U45512 (N_45512,N_44803,N_44819);
xor U45513 (N_45513,N_44776,N_44780);
xnor U45514 (N_45514,N_44807,N_44783);
nand U45515 (N_45515,N_44030,N_44929);
xor U45516 (N_45516,N_44393,N_44097);
or U45517 (N_45517,N_44972,N_44579);
and U45518 (N_45518,N_44435,N_44688);
nand U45519 (N_45519,N_44517,N_44706);
nand U45520 (N_45520,N_44406,N_44241);
nand U45521 (N_45521,N_44152,N_44802);
nor U45522 (N_45522,N_44432,N_44592);
or U45523 (N_45523,N_44311,N_44982);
nand U45524 (N_45524,N_44942,N_44594);
or U45525 (N_45525,N_44110,N_44016);
nand U45526 (N_45526,N_44999,N_44302);
xor U45527 (N_45527,N_44530,N_44531);
nor U45528 (N_45528,N_44460,N_44749);
nor U45529 (N_45529,N_44619,N_44775);
nor U45530 (N_45530,N_44533,N_44275);
or U45531 (N_45531,N_44498,N_44715);
xnor U45532 (N_45532,N_44242,N_44961);
or U45533 (N_45533,N_44462,N_44122);
xnor U45534 (N_45534,N_44979,N_44191);
xnor U45535 (N_45535,N_44270,N_44194);
or U45536 (N_45536,N_44910,N_44886);
and U45537 (N_45537,N_44109,N_44380);
nor U45538 (N_45538,N_44010,N_44415);
and U45539 (N_45539,N_44086,N_44601);
xnor U45540 (N_45540,N_44116,N_44726);
and U45541 (N_45541,N_44573,N_44030);
or U45542 (N_45542,N_44843,N_44507);
nand U45543 (N_45543,N_44114,N_44036);
nor U45544 (N_45544,N_44379,N_44471);
xor U45545 (N_45545,N_44638,N_44850);
nand U45546 (N_45546,N_44775,N_44402);
or U45547 (N_45547,N_44775,N_44501);
or U45548 (N_45548,N_44494,N_44470);
and U45549 (N_45549,N_44768,N_44270);
nand U45550 (N_45550,N_44557,N_44110);
nand U45551 (N_45551,N_44125,N_44042);
and U45552 (N_45552,N_44538,N_44477);
xnor U45553 (N_45553,N_44716,N_44070);
and U45554 (N_45554,N_44595,N_44308);
and U45555 (N_45555,N_44874,N_44248);
and U45556 (N_45556,N_44051,N_44675);
or U45557 (N_45557,N_44992,N_44083);
nand U45558 (N_45558,N_44821,N_44086);
nand U45559 (N_45559,N_44083,N_44845);
nor U45560 (N_45560,N_44008,N_44560);
nor U45561 (N_45561,N_44209,N_44903);
or U45562 (N_45562,N_44149,N_44054);
and U45563 (N_45563,N_44507,N_44462);
nand U45564 (N_45564,N_44422,N_44980);
nor U45565 (N_45565,N_44446,N_44030);
and U45566 (N_45566,N_44276,N_44278);
nor U45567 (N_45567,N_44635,N_44732);
nor U45568 (N_45568,N_44700,N_44082);
nand U45569 (N_45569,N_44066,N_44651);
and U45570 (N_45570,N_44494,N_44090);
nor U45571 (N_45571,N_44131,N_44837);
xor U45572 (N_45572,N_44667,N_44317);
nor U45573 (N_45573,N_44428,N_44371);
and U45574 (N_45574,N_44992,N_44182);
xor U45575 (N_45575,N_44745,N_44266);
nand U45576 (N_45576,N_44898,N_44150);
nor U45577 (N_45577,N_44893,N_44036);
xor U45578 (N_45578,N_44612,N_44647);
xnor U45579 (N_45579,N_44518,N_44706);
nor U45580 (N_45580,N_44204,N_44010);
or U45581 (N_45581,N_44038,N_44758);
xnor U45582 (N_45582,N_44754,N_44360);
nor U45583 (N_45583,N_44023,N_44041);
nand U45584 (N_45584,N_44359,N_44071);
xnor U45585 (N_45585,N_44519,N_44729);
nand U45586 (N_45586,N_44589,N_44512);
xnor U45587 (N_45587,N_44937,N_44982);
nand U45588 (N_45588,N_44521,N_44331);
nor U45589 (N_45589,N_44558,N_44676);
nand U45590 (N_45590,N_44052,N_44733);
nor U45591 (N_45591,N_44378,N_44640);
and U45592 (N_45592,N_44243,N_44778);
and U45593 (N_45593,N_44354,N_44129);
xor U45594 (N_45594,N_44153,N_44174);
xor U45595 (N_45595,N_44590,N_44232);
xnor U45596 (N_45596,N_44384,N_44327);
and U45597 (N_45597,N_44051,N_44343);
nand U45598 (N_45598,N_44462,N_44278);
xor U45599 (N_45599,N_44023,N_44475);
and U45600 (N_45600,N_44789,N_44572);
nor U45601 (N_45601,N_44755,N_44244);
nor U45602 (N_45602,N_44301,N_44776);
or U45603 (N_45603,N_44306,N_44614);
or U45604 (N_45604,N_44717,N_44491);
or U45605 (N_45605,N_44463,N_44980);
and U45606 (N_45606,N_44903,N_44078);
xnor U45607 (N_45607,N_44034,N_44612);
and U45608 (N_45608,N_44167,N_44556);
nor U45609 (N_45609,N_44129,N_44659);
or U45610 (N_45610,N_44622,N_44472);
xnor U45611 (N_45611,N_44464,N_44860);
xnor U45612 (N_45612,N_44039,N_44734);
and U45613 (N_45613,N_44465,N_44381);
nor U45614 (N_45614,N_44006,N_44696);
nor U45615 (N_45615,N_44085,N_44088);
nand U45616 (N_45616,N_44777,N_44711);
nor U45617 (N_45617,N_44162,N_44032);
and U45618 (N_45618,N_44844,N_44706);
and U45619 (N_45619,N_44696,N_44411);
nor U45620 (N_45620,N_44901,N_44426);
nand U45621 (N_45621,N_44723,N_44650);
or U45622 (N_45622,N_44306,N_44754);
nor U45623 (N_45623,N_44126,N_44248);
or U45624 (N_45624,N_44784,N_44622);
and U45625 (N_45625,N_44790,N_44149);
nor U45626 (N_45626,N_44496,N_44400);
and U45627 (N_45627,N_44642,N_44708);
and U45628 (N_45628,N_44098,N_44212);
nor U45629 (N_45629,N_44783,N_44233);
nand U45630 (N_45630,N_44652,N_44010);
or U45631 (N_45631,N_44940,N_44373);
nor U45632 (N_45632,N_44170,N_44439);
and U45633 (N_45633,N_44916,N_44070);
and U45634 (N_45634,N_44342,N_44795);
or U45635 (N_45635,N_44163,N_44025);
or U45636 (N_45636,N_44442,N_44375);
or U45637 (N_45637,N_44553,N_44073);
xnor U45638 (N_45638,N_44633,N_44365);
and U45639 (N_45639,N_44769,N_44538);
xor U45640 (N_45640,N_44495,N_44269);
nand U45641 (N_45641,N_44391,N_44887);
or U45642 (N_45642,N_44412,N_44894);
and U45643 (N_45643,N_44131,N_44390);
and U45644 (N_45644,N_44987,N_44426);
nand U45645 (N_45645,N_44467,N_44968);
or U45646 (N_45646,N_44858,N_44751);
nor U45647 (N_45647,N_44805,N_44853);
or U45648 (N_45648,N_44446,N_44534);
or U45649 (N_45649,N_44238,N_44776);
and U45650 (N_45650,N_44036,N_44851);
nand U45651 (N_45651,N_44925,N_44346);
nor U45652 (N_45652,N_44139,N_44105);
or U45653 (N_45653,N_44569,N_44672);
nor U45654 (N_45654,N_44786,N_44904);
nor U45655 (N_45655,N_44281,N_44052);
and U45656 (N_45656,N_44748,N_44437);
nor U45657 (N_45657,N_44423,N_44207);
and U45658 (N_45658,N_44371,N_44890);
and U45659 (N_45659,N_44140,N_44320);
nor U45660 (N_45660,N_44830,N_44017);
xnor U45661 (N_45661,N_44528,N_44167);
nand U45662 (N_45662,N_44396,N_44289);
nor U45663 (N_45663,N_44187,N_44670);
xor U45664 (N_45664,N_44979,N_44942);
and U45665 (N_45665,N_44982,N_44215);
or U45666 (N_45666,N_44352,N_44923);
nand U45667 (N_45667,N_44611,N_44225);
xor U45668 (N_45668,N_44941,N_44928);
nand U45669 (N_45669,N_44785,N_44406);
nand U45670 (N_45670,N_44108,N_44047);
xor U45671 (N_45671,N_44872,N_44109);
nand U45672 (N_45672,N_44449,N_44059);
or U45673 (N_45673,N_44904,N_44816);
and U45674 (N_45674,N_44257,N_44363);
nor U45675 (N_45675,N_44701,N_44458);
nand U45676 (N_45676,N_44153,N_44463);
nand U45677 (N_45677,N_44658,N_44495);
xor U45678 (N_45678,N_44225,N_44466);
and U45679 (N_45679,N_44457,N_44996);
xnor U45680 (N_45680,N_44925,N_44415);
and U45681 (N_45681,N_44071,N_44329);
or U45682 (N_45682,N_44763,N_44640);
nor U45683 (N_45683,N_44189,N_44629);
nand U45684 (N_45684,N_44634,N_44865);
xnor U45685 (N_45685,N_44811,N_44592);
and U45686 (N_45686,N_44827,N_44904);
xor U45687 (N_45687,N_44747,N_44688);
nand U45688 (N_45688,N_44894,N_44799);
and U45689 (N_45689,N_44348,N_44455);
nor U45690 (N_45690,N_44283,N_44540);
or U45691 (N_45691,N_44507,N_44051);
nand U45692 (N_45692,N_44367,N_44670);
nor U45693 (N_45693,N_44810,N_44471);
nand U45694 (N_45694,N_44304,N_44089);
xnor U45695 (N_45695,N_44791,N_44143);
nand U45696 (N_45696,N_44518,N_44323);
xnor U45697 (N_45697,N_44300,N_44909);
nor U45698 (N_45698,N_44902,N_44307);
nor U45699 (N_45699,N_44752,N_44464);
nand U45700 (N_45700,N_44790,N_44165);
nor U45701 (N_45701,N_44664,N_44630);
or U45702 (N_45702,N_44954,N_44120);
or U45703 (N_45703,N_44034,N_44538);
nand U45704 (N_45704,N_44129,N_44272);
and U45705 (N_45705,N_44795,N_44729);
xor U45706 (N_45706,N_44017,N_44909);
or U45707 (N_45707,N_44395,N_44539);
or U45708 (N_45708,N_44419,N_44040);
nor U45709 (N_45709,N_44571,N_44139);
and U45710 (N_45710,N_44986,N_44702);
or U45711 (N_45711,N_44141,N_44940);
nand U45712 (N_45712,N_44524,N_44515);
nand U45713 (N_45713,N_44026,N_44035);
nand U45714 (N_45714,N_44774,N_44153);
or U45715 (N_45715,N_44738,N_44886);
nand U45716 (N_45716,N_44804,N_44193);
xor U45717 (N_45717,N_44815,N_44111);
or U45718 (N_45718,N_44503,N_44610);
xnor U45719 (N_45719,N_44543,N_44569);
and U45720 (N_45720,N_44473,N_44609);
and U45721 (N_45721,N_44699,N_44807);
and U45722 (N_45722,N_44124,N_44747);
or U45723 (N_45723,N_44956,N_44994);
or U45724 (N_45724,N_44856,N_44677);
or U45725 (N_45725,N_44308,N_44210);
nand U45726 (N_45726,N_44518,N_44498);
nor U45727 (N_45727,N_44257,N_44986);
or U45728 (N_45728,N_44038,N_44791);
nor U45729 (N_45729,N_44079,N_44152);
or U45730 (N_45730,N_44095,N_44171);
xor U45731 (N_45731,N_44715,N_44872);
or U45732 (N_45732,N_44823,N_44721);
nand U45733 (N_45733,N_44885,N_44197);
or U45734 (N_45734,N_44556,N_44330);
and U45735 (N_45735,N_44031,N_44574);
nand U45736 (N_45736,N_44585,N_44720);
or U45737 (N_45737,N_44509,N_44714);
and U45738 (N_45738,N_44968,N_44762);
nand U45739 (N_45739,N_44053,N_44360);
nand U45740 (N_45740,N_44087,N_44561);
or U45741 (N_45741,N_44791,N_44458);
nand U45742 (N_45742,N_44127,N_44109);
nand U45743 (N_45743,N_44152,N_44196);
or U45744 (N_45744,N_44252,N_44137);
xor U45745 (N_45745,N_44523,N_44589);
xnor U45746 (N_45746,N_44297,N_44832);
or U45747 (N_45747,N_44711,N_44213);
or U45748 (N_45748,N_44948,N_44151);
nand U45749 (N_45749,N_44078,N_44853);
or U45750 (N_45750,N_44166,N_44598);
and U45751 (N_45751,N_44689,N_44295);
nor U45752 (N_45752,N_44426,N_44983);
and U45753 (N_45753,N_44843,N_44225);
xnor U45754 (N_45754,N_44172,N_44571);
and U45755 (N_45755,N_44215,N_44623);
nand U45756 (N_45756,N_44609,N_44413);
and U45757 (N_45757,N_44641,N_44337);
xor U45758 (N_45758,N_44414,N_44272);
xor U45759 (N_45759,N_44313,N_44152);
nor U45760 (N_45760,N_44109,N_44966);
xnor U45761 (N_45761,N_44721,N_44817);
and U45762 (N_45762,N_44058,N_44179);
nor U45763 (N_45763,N_44797,N_44698);
or U45764 (N_45764,N_44029,N_44962);
xnor U45765 (N_45765,N_44701,N_44716);
or U45766 (N_45766,N_44239,N_44774);
xnor U45767 (N_45767,N_44995,N_44228);
or U45768 (N_45768,N_44928,N_44072);
xnor U45769 (N_45769,N_44144,N_44338);
nor U45770 (N_45770,N_44062,N_44946);
xnor U45771 (N_45771,N_44619,N_44784);
nand U45772 (N_45772,N_44361,N_44600);
or U45773 (N_45773,N_44099,N_44253);
nand U45774 (N_45774,N_44339,N_44523);
or U45775 (N_45775,N_44772,N_44073);
or U45776 (N_45776,N_44928,N_44028);
and U45777 (N_45777,N_44203,N_44339);
and U45778 (N_45778,N_44575,N_44937);
or U45779 (N_45779,N_44100,N_44312);
or U45780 (N_45780,N_44076,N_44851);
and U45781 (N_45781,N_44543,N_44771);
nand U45782 (N_45782,N_44191,N_44890);
or U45783 (N_45783,N_44555,N_44084);
nor U45784 (N_45784,N_44176,N_44212);
nor U45785 (N_45785,N_44931,N_44286);
nand U45786 (N_45786,N_44316,N_44678);
nor U45787 (N_45787,N_44516,N_44319);
and U45788 (N_45788,N_44890,N_44507);
nor U45789 (N_45789,N_44447,N_44597);
xor U45790 (N_45790,N_44440,N_44157);
or U45791 (N_45791,N_44211,N_44082);
xor U45792 (N_45792,N_44356,N_44517);
xnor U45793 (N_45793,N_44399,N_44763);
xor U45794 (N_45794,N_44137,N_44656);
nand U45795 (N_45795,N_44846,N_44420);
xor U45796 (N_45796,N_44080,N_44205);
and U45797 (N_45797,N_44690,N_44614);
xor U45798 (N_45798,N_44635,N_44755);
and U45799 (N_45799,N_44154,N_44122);
xor U45800 (N_45800,N_44373,N_44569);
nor U45801 (N_45801,N_44762,N_44563);
nand U45802 (N_45802,N_44348,N_44118);
xnor U45803 (N_45803,N_44637,N_44744);
xor U45804 (N_45804,N_44702,N_44129);
or U45805 (N_45805,N_44685,N_44607);
xnor U45806 (N_45806,N_44848,N_44215);
nor U45807 (N_45807,N_44853,N_44876);
xnor U45808 (N_45808,N_44662,N_44183);
or U45809 (N_45809,N_44824,N_44050);
nand U45810 (N_45810,N_44053,N_44738);
nand U45811 (N_45811,N_44143,N_44931);
nor U45812 (N_45812,N_44968,N_44815);
nand U45813 (N_45813,N_44620,N_44942);
or U45814 (N_45814,N_44115,N_44220);
and U45815 (N_45815,N_44796,N_44498);
and U45816 (N_45816,N_44811,N_44999);
nor U45817 (N_45817,N_44923,N_44685);
or U45818 (N_45818,N_44476,N_44985);
or U45819 (N_45819,N_44164,N_44930);
nor U45820 (N_45820,N_44670,N_44603);
nor U45821 (N_45821,N_44602,N_44239);
nor U45822 (N_45822,N_44269,N_44058);
nand U45823 (N_45823,N_44483,N_44271);
xor U45824 (N_45824,N_44813,N_44129);
and U45825 (N_45825,N_44119,N_44921);
or U45826 (N_45826,N_44467,N_44209);
or U45827 (N_45827,N_44487,N_44669);
xor U45828 (N_45828,N_44458,N_44015);
xnor U45829 (N_45829,N_44433,N_44553);
and U45830 (N_45830,N_44405,N_44021);
nand U45831 (N_45831,N_44781,N_44744);
nand U45832 (N_45832,N_44780,N_44044);
nand U45833 (N_45833,N_44933,N_44046);
and U45834 (N_45834,N_44028,N_44329);
xnor U45835 (N_45835,N_44879,N_44303);
and U45836 (N_45836,N_44380,N_44683);
nand U45837 (N_45837,N_44188,N_44824);
and U45838 (N_45838,N_44887,N_44899);
and U45839 (N_45839,N_44468,N_44305);
nor U45840 (N_45840,N_44735,N_44291);
xnor U45841 (N_45841,N_44152,N_44403);
and U45842 (N_45842,N_44846,N_44927);
nand U45843 (N_45843,N_44003,N_44925);
and U45844 (N_45844,N_44379,N_44753);
nor U45845 (N_45845,N_44302,N_44289);
nor U45846 (N_45846,N_44557,N_44276);
or U45847 (N_45847,N_44992,N_44594);
and U45848 (N_45848,N_44795,N_44686);
xnor U45849 (N_45849,N_44937,N_44577);
and U45850 (N_45850,N_44424,N_44910);
and U45851 (N_45851,N_44888,N_44178);
nand U45852 (N_45852,N_44624,N_44325);
nand U45853 (N_45853,N_44351,N_44037);
nand U45854 (N_45854,N_44716,N_44149);
nand U45855 (N_45855,N_44264,N_44533);
nor U45856 (N_45856,N_44223,N_44318);
or U45857 (N_45857,N_44908,N_44659);
nor U45858 (N_45858,N_44553,N_44976);
nor U45859 (N_45859,N_44849,N_44475);
xor U45860 (N_45860,N_44300,N_44110);
nor U45861 (N_45861,N_44085,N_44283);
nand U45862 (N_45862,N_44809,N_44105);
or U45863 (N_45863,N_44579,N_44490);
nand U45864 (N_45864,N_44429,N_44228);
and U45865 (N_45865,N_44772,N_44586);
nand U45866 (N_45866,N_44919,N_44827);
xnor U45867 (N_45867,N_44154,N_44667);
and U45868 (N_45868,N_44872,N_44012);
nand U45869 (N_45869,N_44922,N_44189);
xnor U45870 (N_45870,N_44279,N_44081);
nand U45871 (N_45871,N_44971,N_44445);
nor U45872 (N_45872,N_44828,N_44972);
or U45873 (N_45873,N_44763,N_44491);
nand U45874 (N_45874,N_44783,N_44855);
xnor U45875 (N_45875,N_44505,N_44392);
or U45876 (N_45876,N_44813,N_44569);
and U45877 (N_45877,N_44394,N_44311);
and U45878 (N_45878,N_44689,N_44542);
or U45879 (N_45879,N_44572,N_44418);
xnor U45880 (N_45880,N_44932,N_44143);
or U45881 (N_45881,N_44482,N_44281);
xnor U45882 (N_45882,N_44892,N_44724);
or U45883 (N_45883,N_44901,N_44801);
and U45884 (N_45884,N_44864,N_44918);
nor U45885 (N_45885,N_44806,N_44466);
nand U45886 (N_45886,N_44162,N_44990);
and U45887 (N_45887,N_44614,N_44692);
and U45888 (N_45888,N_44304,N_44414);
or U45889 (N_45889,N_44803,N_44584);
xnor U45890 (N_45890,N_44226,N_44378);
and U45891 (N_45891,N_44522,N_44495);
nand U45892 (N_45892,N_44417,N_44503);
or U45893 (N_45893,N_44375,N_44230);
nand U45894 (N_45894,N_44968,N_44419);
nand U45895 (N_45895,N_44171,N_44871);
and U45896 (N_45896,N_44304,N_44696);
or U45897 (N_45897,N_44546,N_44157);
nand U45898 (N_45898,N_44744,N_44305);
and U45899 (N_45899,N_44957,N_44287);
or U45900 (N_45900,N_44065,N_44920);
or U45901 (N_45901,N_44418,N_44334);
or U45902 (N_45902,N_44335,N_44758);
nor U45903 (N_45903,N_44148,N_44389);
and U45904 (N_45904,N_44990,N_44031);
or U45905 (N_45905,N_44942,N_44065);
or U45906 (N_45906,N_44660,N_44398);
nand U45907 (N_45907,N_44168,N_44689);
nand U45908 (N_45908,N_44552,N_44593);
and U45909 (N_45909,N_44532,N_44751);
nand U45910 (N_45910,N_44858,N_44655);
nor U45911 (N_45911,N_44236,N_44769);
xor U45912 (N_45912,N_44168,N_44578);
or U45913 (N_45913,N_44000,N_44671);
xor U45914 (N_45914,N_44925,N_44015);
nor U45915 (N_45915,N_44995,N_44620);
and U45916 (N_45916,N_44036,N_44002);
nand U45917 (N_45917,N_44319,N_44722);
nor U45918 (N_45918,N_44007,N_44081);
xor U45919 (N_45919,N_44702,N_44182);
nand U45920 (N_45920,N_44936,N_44943);
nor U45921 (N_45921,N_44783,N_44484);
and U45922 (N_45922,N_44487,N_44444);
xor U45923 (N_45923,N_44822,N_44651);
nor U45924 (N_45924,N_44878,N_44541);
nand U45925 (N_45925,N_44174,N_44794);
or U45926 (N_45926,N_44625,N_44847);
and U45927 (N_45927,N_44959,N_44574);
nand U45928 (N_45928,N_44979,N_44169);
xnor U45929 (N_45929,N_44218,N_44333);
nand U45930 (N_45930,N_44858,N_44563);
and U45931 (N_45931,N_44044,N_44498);
and U45932 (N_45932,N_44230,N_44073);
nor U45933 (N_45933,N_44780,N_44254);
or U45934 (N_45934,N_44736,N_44445);
xnor U45935 (N_45935,N_44476,N_44098);
and U45936 (N_45936,N_44504,N_44584);
nand U45937 (N_45937,N_44837,N_44702);
nand U45938 (N_45938,N_44181,N_44380);
or U45939 (N_45939,N_44902,N_44059);
xnor U45940 (N_45940,N_44621,N_44363);
nor U45941 (N_45941,N_44092,N_44889);
and U45942 (N_45942,N_44122,N_44143);
and U45943 (N_45943,N_44746,N_44316);
nand U45944 (N_45944,N_44975,N_44038);
nand U45945 (N_45945,N_44972,N_44939);
or U45946 (N_45946,N_44240,N_44162);
or U45947 (N_45947,N_44887,N_44072);
nor U45948 (N_45948,N_44971,N_44085);
or U45949 (N_45949,N_44602,N_44227);
nor U45950 (N_45950,N_44127,N_44196);
xnor U45951 (N_45951,N_44178,N_44275);
nand U45952 (N_45952,N_44119,N_44166);
nand U45953 (N_45953,N_44434,N_44404);
or U45954 (N_45954,N_44218,N_44320);
xor U45955 (N_45955,N_44562,N_44185);
and U45956 (N_45956,N_44110,N_44364);
nor U45957 (N_45957,N_44459,N_44326);
nor U45958 (N_45958,N_44558,N_44576);
or U45959 (N_45959,N_44846,N_44556);
nand U45960 (N_45960,N_44201,N_44943);
nor U45961 (N_45961,N_44021,N_44848);
nand U45962 (N_45962,N_44822,N_44084);
and U45963 (N_45963,N_44167,N_44686);
xor U45964 (N_45964,N_44293,N_44342);
or U45965 (N_45965,N_44169,N_44624);
nand U45966 (N_45966,N_44806,N_44293);
xnor U45967 (N_45967,N_44123,N_44294);
and U45968 (N_45968,N_44674,N_44193);
or U45969 (N_45969,N_44231,N_44368);
nor U45970 (N_45970,N_44644,N_44187);
nor U45971 (N_45971,N_44564,N_44769);
nor U45972 (N_45972,N_44457,N_44696);
and U45973 (N_45973,N_44554,N_44097);
nor U45974 (N_45974,N_44582,N_44721);
or U45975 (N_45975,N_44185,N_44784);
nand U45976 (N_45976,N_44970,N_44375);
and U45977 (N_45977,N_44599,N_44402);
xor U45978 (N_45978,N_44528,N_44071);
or U45979 (N_45979,N_44621,N_44782);
and U45980 (N_45980,N_44356,N_44773);
or U45981 (N_45981,N_44872,N_44759);
nand U45982 (N_45982,N_44987,N_44880);
or U45983 (N_45983,N_44380,N_44944);
xor U45984 (N_45984,N_44240,N_44001);
and U45985 (N_45985,N_44902,N_44548);
nor U45986 (N_45986,N_44427,N_44325);
and U45987 (N_45987,N_44271,N_44734);
and U45988 (N_45988,N_44421,N_44500);
nor U45989 (N_45989,N_44331,N_44242);
and U45990 (N_45990,N_44101,N_44042);
nor U45991 (N_45991,N_44057,N_44575);
nor U45992 (N_45992,N_44843,N_44900);
xor U45993 (N_45993,N_44595,N_44740);
xnor U45994 (N_45994,N_44942,N_44314);
nor U45995 (N_45995,N_44145,N_44313);
and U45996 (N_45996,N_44076,N_44714);
and U45997 (N_45997,N_44801,N_44001);
or U45998 (N_45998,N_44438,N_44402);
or U45999 (N_45999,N_44046,N_44857);
nand U46000 (N_46000,N_45310,N_45687);
xnor U46001 (N_46001,N_45425,N_45524);
or U46002 (N_46002,N_45428,N_45673);
xnor U46003 (N_46003,N_45419,N_45364);
xnor U46004 (N_46004,N_45485,N_45194);
and U46005 (N_46005,N_45289,N_45674);
and U46006 (N_46006,N_45470,N_45216);
xor U46007 (N_46007,N_45671,N_45219);
and U46008 (N_46008,N_45004,N_45058);
and U46009 (N_46009,N_45884,N_45938);
and U46010 (N_46010,N_45923,N_45521);
nand U46011 (N_46011,N_45082,N_45015);
or U46012 (N_46012,N_45784,N_45456);
nor U46013 (N_46013,N_45440,N_45800);
nand U46014 (N_46014,N_45110,N_45823);
or U46015 (N_46015,N_45556,N_45877);
or U46016 (N_46016,N_45706,N_45436);
nand U46017 (N_46017,N_45595,N_45757);
and U46018 (N_46018,N_45492,N_45870);
nand U46019 (N_46019,N_45410,N_45933);
xnor U46020 (N_46020,N_45718,N_45430);
and U46021 (N_46021,N_45891,N_45481);
and U46022 (N_46022,N_45463,N_45628);
nor U46023 (N_46023,N_45368,N_45005);
nand U46024 (N_46024,N_45383,N_45078);
xnor U46025 (N_46025,N_45531,N_45063);
and U46026 (N_46026,N_45947,N_45061);
xnor U46027 (N_46027,N_45291,N_45306);
and U46028 (N_46028,N_45772,N_45262);
nor U46029 (N_46029,N_45159,N_45208);
nand U46030 (N_46030,N_45661,N_45105);
nand U46031 (N_46031,N_45014,N_45789);
xnor U46032 (N_46032,N_45722,N_45518);
xnor U46033 (N_46033,N_45894,N_45442);
nor U46034 (N_46034,N_45948,N_45809);
and U46035 (N_46035,N_45545,N_45685);
or U46036 (N_46036,N_45587,N_45163);
nand U46037 (N_46037,N_45259,N_45824);
nor U46038 (N_46038,N_45752,N_45804);
or U46039 (N_46039,N_45856,N_45966);
xor U46040 (N_46040,N_45953,N_45267);
or U46041 (N_46041,N_45094,N_45618);
nor U46042 (N_46042,N_45901,N_45801);
or U46043 (N_46043,N_45986,N_45557);
and U46044 (N_46044,N_45125,N_45406);
xor U46045 (N_46045,N_45820,N_45853);
nand U46046 (N_46046,N_45493,N_45985);
xnor U46047 (N_46047,N_45220,N_45715);
and U46048 (N_46048,N_45304,N_45756);
nor U46049 (N_46049,N_45630,N_45994);
xor U46050 (N_46050,N_45731,N_45039);
xnor U46051 (N_46051,N_45995,N_45051);
or U46052 (N_46052,N_45583,N_45249);
xnor U46053 (N_46053,N_45904,N_45581);
or U46054 (N_46054,N_45975,N_45598);
and U46055 (N_46055,N_45634,N_45132);
xor U46056 (N_46056,N_45644,N_45530);
and U46057 (N_46057,N_45964,N_45234);
nor U46058 (N_46058,N_45192,N_45026);
nand U46059 (N_46059,N_45504,N_45010);
and U46060 (N_46060,N_45501,N_45137);
nand U46061 (N_46061,N_45865,N_45505);
nor U46062 (N_46062,N_45596,N_45754);
nor U46063 (N_46063,N_45251,N_45957);
nor U46064 (N_46064,N_45069,N_45832);
and U46065 (N_46065,N_45777,N_45164);
nor U46066 (N_46066,N_45215,N_45882);
or U46067 (N_46067,N_45334,N_45041);
xnor U46068 (N_46068,N_45317,N_45427);
nand U46069 (N_46069,N_45211,N_45792);
xnor U46070 (N_46070,N_45560,N_45639);
nand U46071 (N_46071,N_45315,N_45897);
nor U46072 (N_46072,N_45303,N_45418);
xnor U46073 (N_46073,N_45642,N_45741);
nor U46074 (N_46074,N_45799,N_45072);
xor U46075 (N_46075,N_45200,N_45511);
nand U46076 (N_46076,N_45042,N_45247);
xor U46077 (N_46077,N_45539,N_45830);
and U46078 (N_46078,N_45305,N_45815);
nand U46079 (N_46079,N_45478,N_45765);
nand U46080 (N_46080,N_45950,N_45468);
nand U46081 (N_46081,N_45389,N_45561);
nor U46082 (N_46082,N_45030,N_45028);
xor U46083 (N_46083,N_45136,N_45935);
nand U46084 (N_46084,N_45198,N_45623);
or U46085 (N_46085,N_45180,N_45373);
and U46086 (N_46086,N_45625,N_45532);
or U46087 (N_46087,N_45977,N_45467);
and U46088 (N_46088,N_45140,N_45697);
and U46089 (N_46089,N_45817,N_45483);
nand U46090 (N_46090,N_45878,N_45096);
nor U46091 (N_46091,N_45274,N_45664);
nand U46092 (N_46092,N_45747,N_45038);
nand U46093 (N_46093,N_45086,N_45496);
and U46094 (N_46094,N_45860,N_45896);
and U46095 (N_46095,N_45759,N_45678);
or U46096 (N_46096,N_45265,N_45112);
nor U46097 (N_46097,N_45502,N_45775);
nor U46098 (N_46098,N_45057,N_45528);
nor U46099 (N_46099,N_45764,N_45139);
xnor U46100 (N_46100,N_45808,N_45812);
xor U46101 (N_46101,N_45450,N_45121);
or U46102 (N_46102,N_45490,N_45133);
or U46103 (N_46103,N_45308,N_45827);
nand U46104 (N_46104,N_45189,N_45095);
nand U46105 (N_46105,N_45349,N_45423);
xor U46106 (N_46106,N_45847,N_45783);
nor U46107 (N_46107,N_45537,N_45340);
nor U46108 (N_46108,N_45512,N_45184);
nand U46109 (N_46109,N_45321,N_45118);
nand U46110 (N_46110,N_45700,N_45647);
nor U46111 (N_46111,N_45908,N_45543);
and U46112 (N_46112,N_45148,N_45793);
or U46113 (N_46113,N_45965,N_45941);
nor U46114 (N_46114,N_45873,N_45367);
nor U46115 (N_46115,N_45365,N_45407);
or U46116 (N_46116,N_45395,N_45107);
and U46117 (N_46117,N_45721,N_45233);
nor U46118 (N_46118,N_45602,N_45971);
nor U46119 (N_46119,N_45314,N_45239);
nor U46120 (N_46120,N_45930,N_45093);
nor U46121 (N_46121,N_45613,N_45982);
and U46122 (N_46122,N_45144,N_45952);
nand U46123 (N_46123,N_45869,N_45175);
nand U46124 (N_46124,N_45185,N_45236);
xor U46125 (N_46125,N_45085,N_45655);
xnor U46126 (N_46126,N_45191,N_45196);
xor U46127 (N_46127,N_45210,N_45794);
xor U46128 (N_46128,N_45569,N_45115);
nor U46129 (N_46129,N_45988,N_45577);
nand U46130 (N_46130,N_45600,N_45143);
and U46131 (N_46131,N_45465,N_45646);
or U46132 (N_46132,N_45282,N_45513);
xor U46133 (N_46133,N_45405,N_45199);
and U46134 (N_46134,N_45393,N_45857);
or U46135 (N_46135,N_45762,N_45432);
and U46136 (N_46136,N_45842,N_45221);
nand U46137 (N_46137,N_45408,N_45173);
and U46138 (N_46138,N_45566,N_45920);
xnor U46139 (N_46139,N_45302,N_45424);
or U46140 (N_46140,N_45202,N_45052);
xor U46141 (N_46141,N_45134,N_45795);
nor U46142 (N_46142,N_45962,N_45377);
nand U46143 (N_46143,N_45796,N_45912);
nand U46144 (N_46144,N_45821,N_45846);
nor U46145 (N_46145,N_45029,N_45593);
xor U46146 (N_46146,N_45227,N_45811);
and U46147 (N_46147,N_45611,N_45346);
and U46148 (N_46148,N_45361,N_45854);
xnor U46149 (N_46149,N_45711,N_45044);
xnor U46150 (N_46150,N_45100,N_45620);
nor U46151 (N_46151,N_45914,N_45120);
nor U46152 (N_46152,N_45619,N_45769);
xnor U46153 (N_46153,N_45260,N_45209);
nand U46154 (N_46154,N_45043,N_45339);
and U46155 (N_46155,N_45983,N_45165);
or U46156 (N_46156,N_45401,N_45714);
nand U46157 (N_46157,N_45375,N_45328);
xnor U46158 (N_46158,N_45129,N_45855);
or U46159 (N_46159,N_45515,N_45932);
and U46160 (N_46160,N_45222,N_45807);
xnor U46161 (N_46161,N_45244,N_45659);
xor U46162 (N_46162,N_45391,N_45025);
or U46163 (N_46163,N_45437,N_45936);
nor U46164 (N_46164,N_45763,N_45183);
xnor U46165 (N_46165,N_45997,N_45974);
xnor U46166 (N_46166,N_45875,N_45381);
nand U46167 (N_46167,N_45411,N_45895);
xnor U46168 (N_46168,N_45555,N_45152);
nand U46169 (N_46169,N_45802,N_45122);
and U46170 (N_46170,N_45048,N_45636);
nor U46171 (N_46171,N_45273,N_45226);
xor U46172 (N_46172,N_45774,N_45670);
nand U46173 (N_46173,N_45441,N_45024);
xnor U46174 (N_46174,N_45961,N_45476);
xnor U46175 (N_46175,N_45336,N_45937);
nor U46176 (N_46176,N_45154,N_45240);
nor U46177 (N_46177,N_45751,N_45522);
nor U46178 (N_46178,N_45635,N_45667);
nand U46179 (N_46179,N_45307,N_45461);
nand U46180 (N_46180,N_45197,N_45352);
xor U46181 (N_46181,N_45167,N_45263);
nor U46182 (N_46182,N_45068,N_45387);
xor U46183 (N_46183,N_45797,N_45235);
nand U46184 (N_46184,N_45392,N_45416);
and U46185 (N_46185,N_45867,N_45370);
and U46186 (N_46186,N_45420,N_45733);
nand U46187 (N_46187,N_45980,N_45178);
nand U46188 (N_46188,N_45627,N_45926);
nor U46189 (N_46189,N_45444,N_45839);
xor U46190 (N_46190,N_45519,N_45651);
or U46191 (N_46191,N_45770,N_45089);
and U46192 (N_46192,N_45360,N_45160);
nand U46193 (N_46193,N_45541,N_45217);
and U46194 (N_46194,N_45604,N_45905);
and U46195 (N_46195,N_45347,N_45939);
nand U46196 (N_46196,N_45059,N_45656);
and U46197 (N_46197,N_45993,N_45978);
or U46198 (N_46198,N_45924,N_45325);
or U46199 (N_46199,N_45149,N_45617);
and U46200 (N_46200,N_45699,N_45323);
nand U46201 (N_46201,N_45172,N_45117);
or U46202 (N_46202,N_45469,N_45091);
and U46203 (N_46203,N_45327,N_45248);
xnor U46204 (N_46204,N_45145,N_45443);
or U46205 (N_46205,N_45818,N_45934);
nand U46206 (N_46206,N_45535,N_45421);
or U46207 (N_46207,N_45214,N_45701);
and U46208 (N_46208,N_45500,N_45998);
or U46209 (N_46209,N_45987,N_45626);
xor U46210 (N_46210,N_45119,N_45009);
nor U46211 (N_46211,N_45527,N_45076);
nor U46212 (N_46212,N_45679,N_45445);
and U46213 (N_46213,N_45071,N_45633);
and U46214 (N_46214,N_45771,N_45487);
nand U46215 (N_46215,N_45237,N_45554);
and U46216 (N_46216,N_45562,N_45653);
nand U46217 (N_46217,N_45768,N_45023);
nand U46218 (N_46218,N_45850,N_45288);
nand U46219 (N_46219,N_45459,N_45745);
nand U46220 (N_46220,N_45454,N_45438);
nand U46221 (N_46221,N_45312,N_45886);
and U46222 (N_46222,N_45065,N_45313);
and U46223 (N_46223,N_45296,N_45081);
or U46224 (N_46224,N_45447,N_45640);
xnor U46225 (N_46225,N_45195,N_45969);
nor U46226 (N_46226,N_45147,N_45879);
or U46227 (N_46227,N_45669,N_45637);
xnor U46228 (N_46228,N_45477,N_45422);
nand U46229 (N_46229,N_45999,N_45691);
xnor U46230 (N_46230,N_45471,N_45694);
nor U46231 (N_46231,N_45666,N_45177);
or U46232 (N_46232,N_45020,N_45601);
nand U46233 (N_46233,N_45413,N_45169);
xor U46234 (N_46234,N_45786,N_45371);
nand U46235 (N_46235,N_45123,N_45036);
or U46236 (N_46236,N_45675,N_45648);
or U46237 (N_46237,N_45482,N_45355);
or U46238 (N_46238,N_45663,N_45458);
and U46239 (N_46239,N_45337,N_45275);
xnor U46240 (N_46240,N_45689,N_45736);
or U46241 (N_46241,N_45698,N_45344);
xor U46242 (N_46242,N_45429,N_45403);
and U46243 (N_46243,N_45060,N_45106);
and U46244 (N_46244,N_45677,N_45351);
nand U46245 (N_46245,N_45358,N_45206);
xor U46246 (N_46246,N_45097,N_45281);
and U46247 (N_46247,N_45079,N_45001);
xnor U46248 (N_46248,N_45271,N_45942);
nor U46249 (N_46249,N_45074,N_45342);
nor U46250 (N_46250,N_45622,N_45798);
or U46251 (N_46251,N_45514,N_45890);
nor U46252 (N_46252,N_45725,N_45976);
or U46253 (N_46253,N_45826,N_45376);
or U46254 (N_46254,N_45567,N_45055);
or U46255 (N_46255,N_45297,N_45256);
nor U46256 (N_46256,N_45399,N_45766);
nor U46257 (N_46257,N_45668,N_45844);
nor U46258 (N_46258,N_45868,N_45650);
and U46259 (N_46259,N_45050,N_45610);
and U46260 (N_46260,N_45494,N_45520);
nor U46261 (N_46261,N_45728,N_45146);
or U46262 (N_46262,N_45084,N_45362);
nor U46263 (N_46263,N_45991,N_45290);
nand U46264 (N_46264,N_45047,N_45828);
nor U46265 (N_46265,N_45755,N_45021);
nand U46266 (N_46266,N_45729,N_45128);
nor U46267 (N_46267,N_45300,N_45474);
nor U46268 (N_46268,N_45298,N_45054);
nor U46269 (N_46269,N_45921,N_45584);
or U46270 (N_46270,N_45466,N_45283);
nor U46271 (N_46271,N_45131,N_45831);
nor U46272 (N_46272,N_45603,N_45124);
nand U46273 (N_46273,N_45922,N_45384);
and U46274 (N_46274,N_45907,N_45187);
nor U46275 (N_46275,N_45268,N_45951);
nand U46276 (N_46276,N_45205,N_45077);
nand U46277 (N_46277,N_45223,N_45254);
nand U46278 (N_46278,N_45067,N_45092);
xnor U46279 (N_46279,N_45909,N_45301);
nor U46280 (N_46280,N_45724,N_45785);
nand U46281 (N_46281,N_45981,N_45404);
nor U46282 (N_46282,N_45819,N_45088);
xor U46283 (N_46283,N_45871,N_45130);
nand U46284 (N_46284,N_45643,N_45286);
nand U46285 (N_46285,N_45435,N_45155);
nor U46286 (N_46286,N_45887,N_45484);
xnor U46287 (N_46287,N_45350,N_45734);
or U46288 (N_46288,N_45585,N_45898);
and U46289 (N_46289,N_45900,N_45324);
nor U46290 (N_46290,N_45838,N_45954);
or U46291 (N_46291,N_45616,N_45990);
and U46292 (N_46292,N_45564,N_45848);
or U46293 (N_46293,N_45386,N_45712);
nor U46294 (N_46294,N_45503,N_45586);
or U46295 (N_46295,N_45565,N_45621);
xnor U46296 (N_46296,N_45695,N_45388);
and U46297 (N_46297,N_45885,N_45707);
xor U46298 (N_46298,N_45012,N_45902);
xor U46299 (N_46299,N_45116,N_45207);
nand U46300 (N_46300,N_45927,N_45665);
nand U46301 (N_46301,N_45176,N_45692);
nand U46302 (N_46302,N_45166,N_45426);
nand U46303 (N_46303,N_45672,N_45135);
or U46304 (N_46304,N_45333,N_45737);
and U46305 (N_46305,N_45582,N_45016);
or U46306 (N_46306,N_45753,N_45533);
nor U46307 (N_46307,N_45141,N_45363);
nor U46308 (N_46308,N_45473,N_45758);
or U46309 (N_46309,N_45780,N_45446);
nand U46310 (N_46310,N_45790,N_45491);
xor U46311 (N_46311,N_45967,N_45017);
and U46312 (N_46312,N_45833,N_45781);
xnor U46313 (N_46313,N_45385,N_45917);
xor U46314 (N_46314,N_45657,N_45835);
or U46315 (N_46315,N_45632,N_45114);
nor U46316 (N_46316,N_45309,N_45874);
or U46317 (N_46317,N_45919,N_45099);
or U46318 (N_46318,N_45190,N_45179);
xor U46319 (N_46319,N_45609,N_45536);
or U46320 (N_46320,N_45615,N_45931);
nor U46321 (N_46321,N_45412,N_45834);
or U46322 (N_46322,N_45479,N_45318);
xor U46323 (N_46323,N_45335,N_45040);
nand U46324 (N_46324,N_45726,N_45959);
nor U46325 (N_46325,N_45480,N_45322);
xnor U46326 (N_46326,N_45570,N_45013);
and U46327 (N_46327,N_45242,N_45683);
nand U46328 (N_46328,N_45744,N_45488);
and U46329 (N_46329,N_45153,N_45398);
xnor U46330 (N_46330,N_45910,N_45238);
nor U46331 (N_46331,N_45498,N_45066);
nand U46332 (N_46332,N_45574,N_45778);
and U46333 (N_46333,N_45973,N_45658);
or U46334 (N_46334,N_45472,N_45285);
nor U46335 (N_46335,N_45022,N_45127);
xnor U46336 (N_46336,N_45279,N_45080);
or U46337 (N_46337,N_45918,N_45944);
or U46338 (N_46338,N_45649,N_45203);
and U46339 (N_46339,N_45433,N_45645);
and U46340 (N_46340,N_45805,N_45849);
xor U46341 (N_46341,N_45767,N_45270);
or U46342 (N_46342,N_45027,N_45588);
and U46343 (N_46343,N_45292,N_45031);
nor U46344 (N_46344,N_45348,N_45045);
nor U46345 (N_46345,N_45552,N_45578);
xnor U46346 (N_46346,N_45686,N_45837);
nand U46347 (N_46347,N_45864,N_45558);
nor U46348 (N_46348,N_45453,N_45002);
nor U46349 (N_46349,N_45193,N_45546);
nand U46350 (N_46350,N_45224,N_45580);
nor U46351 (N_46351,N_45703,N_45157);
nand U46352 (N_46352,N_45813,N_45330);
or U46353 (N_46353,N_45353,N_45508);
nand U46354 (N_46354,N_45963,N_45597);
nand U46355 (N_46355,N_45989,N_45892);
or U46356 (N_46356,N_45538,N_45840);
nand U46357 (N_46357,N_45161,N_45229);
nand U46358 (N_46358,N_45046,N_45573);
xnor U46359 (N_46359,N_45250,N_45571);
and U46360 (N_46360,N_45378,N_45186);
and U46361 (N_46361,N_45006,N_45380);
nand U46362 (N_46362,N_45594,N_45563);
and U46363 (N_46363,N_45329,N_45037);
xor U46364 (N_46364,N_45320,N_45409);
xnor U46365 (N_46365,N_45782,N_45497);
nor U46366 (N_46366,N_45277,N_45319);
and U46367 (N_46367,N_45690,N_45641);
or U46368 (N_46368,N_45851,N_45280);
nor U46369 (N_46369,N_45579,N_45572);
nand U46370 (N_46370,N_45943,N_45624);
and U46371 (N_46371,N_45181,N_45899);
nand U46372 (N_46372,N_45742,N_45032);
xnor U46373 (N_46373,N_45372,N_45204);
nand U46374 (N_46374,N_45019,N_45761);
xnor U46375 (N_46375,N_45232,N_45760);
or U46376 (N_46376,N_45863,N_45970);
and U46377 (N_46377,N_45499,N_45684);
nand U46378 (N_46378,N_45822,N_45652);
xor U46379 (N_46379,N_45956,N_45568);
xor U46380 (N_46380,N_45269,N_45101);
nor U46381 (N_46381,N_45979,N_45748);
nand U46382 (N_46382,N_45676,N_45607);
nand U46383 (N_46383,N_45743,N_45911);
and U46384 (N_46384,N_45083,N_45170);
or U46385 (N_46385,N_45266,N_45916);
nand U46386 (N_46386,N_45218,N_45287);
nand U46387 (N_46387,N_45495,N_45738);
and U46388 (N_46388,N_45608,N_45551);
and U46389 (N_46389,N_45893,N_45462);
nand U46390 (N_46390,N_45968,N_45258);
or U46391 (N_46391,N_45787,N_45548);
and U46392 (N_46392,N_45230,N_45201);
nor U46393 (N_46393,N_45311,N_45704);
xnor U46394 (N_46394,N_45862,N_45841);
nand U46395 (N_46395,N_45246,N_45845);
and U46396 (N_46396,N_45168,N_45984);
xnor U46397 (N_46397,N_45188,N_45278);
or U46398 (N_46398,N_45245,N_45241);
or U46399 (N_46399,N_45379,N_45606);
nor U46400 (N_46400,N_45612,N_45925);
nand U46401 (N_46401,N_45660,N_45688);
and U46402 (N_46402,N_45814,N_45903);
nor U46403 (N_46403,N_45090,N_45880);
nor U46404 (N_46404,N_45946,N_45872);
nor U46405 (N_46405,N_45151,N_45705);
nand U46406 (N_46406,N_45889,N_45575);
and U46407 (N_46407,N_45171,N_45945);
nand U46408 (N_46408,N_45605,N_45272);
xor U46409 (N_46409,N_45033,N_45331);
xnor U46410 (N_46410,N_45174,N_45517);
nor U46411 (N_46411,N_45382,N_45225);
nand U46412 (N_46412,N_45400,N_45727);
nor U46413 (N_46413,N_45464,N_45915);
nor U46414 (N_46414,N_45709,N_45662);
nand U46415 (N_46415,N_45070,N_45680);
nor U46416 (N_46416,N_45111,N_45011);
nand U46417 (N_46417,N_45414,N_45779);
and U46418 (N_46418,N_45859,N_45452);
nand U46419 (N_46419,N_45955,N_45791);
or U46420 (N_46420,N_45631,N_45261);
nand U46421 (N_46421,N_45750,N_45150);
or U46422 (N_46422,N_45591,N_45843);
or U46423 (N_46423,N_45906,N_45213);
xor U46424 (N_46424,N_45509,N_45374);
xor U46425 (N_46425,N_45341,N_45776);
xnor U46426 (N_46426,N_45888,N_45345);
or U46427 (N_46427,N_45053,N_45018);
nand U46428 (N_46428,N_45866,N_45996);
or U46429 (N_46429,N_45876,N_45294);
xor U46430 (N_46430,N_45434,N_45702);
or U46431 (N_46431,N_45449,N_45293);
xor U46432 (N_46432,N_45460,N_45534);
and U46433 (N_46433,N_45252,N_45559);
xor U46434 (N_46434,N_45682,N_45062);
nor U46435 (N_46435,N_45087,N_45696);
xnor U46436 (N_46436,N_45913,N_45212);
nand U46437 (N_46437,N_45264,N_45356);
nand U46438 (N_46438,N_45506,N_45730);
xnor U46439 (N_46439,N_45681,N_45858);
and U46440 (N_46440,N_45836,N_45654);
nor U46441 (N_46441,N_45881,N_45158);
nand U46442 (N_46442,N_45576,N_45369);
nor U46443 (N_46443,N_45929,N_45056);
or U46444 (N_46444,N_45861,N_45883);
nor U46445 (N_46445,N_45773,N_45717);
nor U46446 (N_46446,N_45710,N_45544);
xor U46447 (N_46447,N_45525,N_45732);
nand U46448 (N_46448,N_45486,N_45960);
nand U46449 (N_46449,N_45540,N_45803);
nand U46450 (N_46450,N_45708,N_45402);
and U46451 (N_46451,N_45231,N_45394);
nand U46452 (N_46452,N_45138,N_45550);
nand U46453 (N_46453,N_45940,N_45735);
nor U46454 (N_46454,N_45113,N_45589);
nand U46455 (N_46455,N_45825,N_45357);
xnor U46456 (N_46456,N_45299,N_45713);
or U46457 (N_46457,N_45949,N_45316);
and U46458 (N_46458,N_45338,N_45523);
xnor U46459 (N_46459,N_45390,N_45507);
nand U46460 (N_46460,N_45720,N_45098);
and U46461 (N_46461,N_45284,N_45049);
nor U46462 (N_46462,N_45716,N_45034);
nand U46463 (N_46463,N_45788,N_45516);
nand U46464 (N_46464,N_45739,N_45629);
nand U46465 (N_46465,N_45276,N_45104);
nor U46466 (N_46466,N_45542,N_45156);
nand U46467 (N_46467,N_45003,N_45992);
nand U46468 (N_46468,N_45599,N_45638);
nor U46469 (N_46469,N_45852,N_45719);
nand U46470 (N_46470,N_45035,N_45972);
nor U46471 (N_46471,N_45332,N_45489);
xnor U46472 (N_46472,N_45526,N_45243);
or U46473 (N_46473,N_45397,N_45354);
or U46474 (N_46474,N_45928,N_45142);
xor U46475 (N_46475,N_45475,N_45228);
and U46476 (N_46476,N_45326,N_45108);
and U46477 (N_46477,N_45126,N_45359);
xor U46478 (N_46478,N_45257,N_45806);
nand U46479 (N_46479,N_45162,N_45547);
nor U46480 (N_46480,N_45109,N_45749);
and U46481 (N_46481,N_45439,N_45451);
nor U46482 (N_46482,N_45592,N_45295);
and U46483 (N_46483,N_45343,N_45958);
xnor U46484 (N_46484,N_45529,N_45075);
nand U46485 (N_46485,N_45740,N_45553);
nor U46486 (N_46486,N_45510,N_45103);
xnor U46487 (N_46487,N_45417,N_45816);
nand U46488 (N_46488,N_45008,N_45448);
and U46489 (N_46489,N_45746,N_45829);
nand U46490 (N_46490,N_45366,N_45693);
nand U46491 (N_46491,N_45000,N_45723);
and U46492 (N_46492,N_45007,N_45590);
or U46493 (N_46493,N_45810,N_45614);
or U46494 (N_46494,N_45073,N_45415);
xnor U46495 (N_46495,N_45182,N_45253);
and U46496 (N_46496,N_45396,N_45255);
and U46497 (N_46497,N_45457,N_45549);
and U46498 (N_46498,N_45431,N_45102);
nand U46499 (N_46499,N_45064,N_45455);
nand U46500 (N_46500,N_45259,N_45995);
xor U46501 (N_46501,N_45286,N_45413);
xnor U46502 (N_46502,N_45845,N_45377);
nand U46503 (N_46503,N_45205,N_45484);
or U46504 (N_46504,N_45750,N_45752);
nand U46505 (N_46505,N_45395,N_45513);
xor U46506 (N_46506,N_45764,N_45860);
and U46507 (N_46507,N_45759,N_45517);
nand U46508 (N_46508,N_45395,N_45234);
xnor U46509 (N_46509,N_45603,N_45801);
nand U46510 (N_46510,N_45563,N_45308);
xor U46511 (N_46511,N_45784,N_45619);
and U46512 (N_46512,N_45343,N_45102);
or U46513 (N_46513,N_45887,N_45836);
nand U46514 (N_46514,N_45753,N_45505);
nor U46515 (N_46515,N_45905,N_45488);
nand U46516 (N_46516,N_45992,N_45598);
xor U46517 (N_46517,N_45411,N_45882);
nand U46518 (N_46518,N_45403,N_45813);
nor U46519 (N_46519,N_45976,N_45701);
nor U46520 (N_46520,N_45888,N_45462);
or U46521 (N_46521,N_45370,N_45521);
and U46522 (N_46522,N_45146,N_45254);
or U46523 (N_46523,N_45423,N_45659);
nor U46524 (N_46524,N_45954,N_45569);
nor U46525 (N_46525,N_45671,N_45928);
xnor U46526 (N_46526,N_45888,N_45610);
and U46527 (N_46527,N_45856,N_45992);
nor U46528 (N_46528,N_45008,N_45015);
and U46529 (N_46529,N_45185,N_45458);
xnor U46530 (N_46530,N_45975,N_45128);
xor U46531 (N_46531,N_45830,N_45398);
or U46532 (N_46532,N_45021,N_45680);
and U46533 (N_46533,N_45458,N_45487);
xor U46534 (N_46534,N_45736,N_45767);
nor U46535 (N_46535,N_45704,N_45050);
and U46536 (N_46536,N_45170,N_45008);
and U46537 (N_46537,N_45480,N_45691);
xnor U46538 (N_46538,N_45344,N_45061);
xor U46539 (N_46539,N_45679,N_45514);
or U46540 (N_46540,N_45206,N_45263);
nor U46541 (N_46541,N_45246,N_45406);
nor U46542 (N_46542,N_45132,N_45032);
and U46543 (N_46543,N_45074,N_45119);
or U46544 (N_46544,N_45593,N_45767);
xor U46545 (N_46545,N_45126,N_45732);
nand U46546 (N_46546,N_45219,N_45737);
and U46547 (N_46547,N_45493,N_45626);
xnor U46548 (N_46548,N_45586,N_45371);
nor U46549 (N_46549,N_45223,N_45766);
nand U46550 (N_46550,N_45142,N_45793);
nand U46551 (N_46551,N_45164,N_45139);
or U46552 (N_46552,N_45139,N_45050);
nand U46553 (N_46553,N_45167,N_45129);
or U46554 (N_46554,N_45042,N_45005);
or U46555 (N_46555,N_45212,N_45957);
xor U46556 (N_46556,N_45581,N_45726);
nand U46557 (N_46557,N_45366,N_45455);
nor U46558 (N_46558,N_45413,N_45933);
nor U46559 (N_46559,N_45159,N_45123);
xnor U46560 (N_46560,N_45327,N_45752);
and U46561 (N_46561,N_45714,N_45225);
xor U46562 (N_46562,N_45034,N_45462);
or U46563 (N_46563,N_45042,N_45826);
or U46564 (N_46564,N_45336,N_45984);
nor U46565 (N_46565,N_45313,N_45737);
nand U46566 (N_46566,N_45337,N_45670);
nor U46567 (N_46567,N_45150,N_45104);
and U46568 (N_46568,N_45326,N_45797);
nand U46569 (N_46569,N_45894,N_45575);
or U46570 (N_46570,N_45738,N_45422);
and U46571 (N_46571,N_45489,N_45844);
or U46572 (N_46572,N_45487,N_45502);
and U46573 (N_46573,N_45881,N_45416);
nor U46574 (N_46574,N_45143,N_45705);
nand U46575 (N_46575,N_45801,N_45248);
nand U46576 (N_46576,N_45551,N_45196);
nand U46577 (N_46577,N_45714,N_45725);
and U46578 (N_46578,N_45588,N_45241);
and U46579 (N_46579,N_45257,N_45638);
nor U46580 (N_46580,N_45547,N_45751);
nand U46581 (N_46581,N_45800,N_45998);
xor U46582 (N_46582,N_45222,N_45763);
nor U46583 (N_46583,N_45438,N_45362);
or U46584 (N_46584,N_45438,N_45472);
nor U46585 (N_46585,N_45748,N_45722);
and U46586 (N_46586,N_45783,N_45795);
and U46587 (N_46587,N_45080,N_45321);
nand U46588 (N_46588,N_45533,N_45714);
xnor U46589 (N_46589,N_45981,N_45089);
and U46590 (N_46590,N_45578,N_45475);
nand U46591 (N_46591,N_45961,N_45698);
xnor U46592 (N_46592,N_45592,N_45109);
xor U46593 (N_46593,N_45646,N_45325);
nand U46594 (N_46594,N_45286,N_45545);
nand U46595 (N_46595,N_45112,N_45183);
nor U46596 (N_46596,N_45284,N_45344);
and U46597 (N_46597,N_45154,N_45747);
xor U46598 (N_46598,N_45872,N_45730);
nand U46599 (N_46599,N_45927,N_45494);
or U46600 (N_46600,N_45285,N_45363);
nor U46601 (N_46601,N_45359,N_45184);
and U46602 (N_46602,N_45427,N_45899);
or U46603 (N_46603,N_45454,N_45694);
or U46604 (N_46604,N_45867,N_45722);
xor U46605 (N_46605,N_45321,N_45923);
xor U46606 (N_46606,N_45088,N_45778);
or U46607 (N_46607,N_45087,N_45342);
nor U46608 (N_46608,N_45808,N_45490);
nor U46609 (N_46609,N_45580,N_45091);
nor U46610 (N_46610,N_45312,N_45997);
or U46611 (N_46611,N_45987,N_45461);
xnor U46612 (N_46612,N_45883,N_45985);
and U46613 (N_46613,N_45124,N_45294);
nand U46614 (N_46614,N_45264,N_45842);
xnor U46615 (N_46615,N_45022,N_45081);
nand U46616 (N_46616,N_45708,N_45248);
and U46617 (N_46617,N_45537,N_45027);
nand U46618 (N_46618,N_45971,N_45584);
nor U46619 (N_46619,N_45361,N_45771);
xnor U46620 (N_46620,N_45022,N_45166);
xnor U46621 (N_46621,N_45846,N_45302);
nand U46622 (N_46622,N_45634,N_45267);
nand U46623 (N_46623,N_45303,N_45936);
nor U46624 (N_46624,N_45162,N_45899);
xnor U46625 (N_46625,N_45902,N_45977);
xor U46626 (N_46626,N_45603,N_45048);
xnor U46627 (N_46627,N_45090,N_45934);
xnor U46628 (N_46628,N_45042,N_45557);
xor U46629 (N_46629,N_45345,N_45413);
or U46630 (N_46630,N_45641,N_45531);
and U46631 (N_46631,N_45663,N_45604);
nand U46632 (N_46632,N_45933,N_45393);
and U46633 (N_46633,N_45838,N_45994);
nand U46634 (N_46634,N_45105,N_45148);
and U46635 (N_46635,N_45048,N_45173);
and U46636 (N_46636,N_45430,N_45907);
nand U46637 (N_46637,N_45753,N_45608);
nand U46638 (N_46638,N_45264,N_45055);
nor U46639 (N_46639,N_45114,N_45753);
xor U46640 (N_46640,N_45719,N_45150);
nor U46641 (N_46641,N_45346,N_45407);
xor U46642 (N_46642,N_45211,N_45271);
and U46643 (N_46643,N_45976,N_45866);
and U46644 (N_46644,N_45403,N_45001);
nand U46645 (N_46645,N_45853,N_45790);
nand U46646 (N_46646,N_45693,N_45880);
nor U46647 (N_46647,N_45612,N_45335);
xnor U46648 (N_46648,N_45098,N_45572);
xnor U46649 (N_46649,N_45504,N_45109);
nand U46650 (N_46650,N_45247,N_45923);
nor U46651 (N_46651,N_45756,N_45604);
nor U46652 (N_46652,N_45247,N_45831);
xnor U46653 (N_46653,N_45711,N_45512);
and U46654 (N_46654,N_45451,N_45106);
xor U46655 (N_46655,N_45760,N_45112);
xnor U46656 (N_46656,N_45410,N_45372);
nand U46657 (N_46657,N_45211,N_45137);
or U46658 (N_46658,N_45322,N_45154);
nand U46659 (N_46659,N_45411,N_45649);
nor U46660 (N_46660,N_45797,N_45545);
and U46661 (N_46661,N_45058,N_45588);
or U46662 (N_46662,N_45185,N_45629);
or U46663 (N_46663,N_45424,N_45027);
nor U46664 (N_46664,N_45934,N_45733);
nor U46665 (N_46665,N_45100,N_45807);
nor U46666 (N_46666,N_45397,N_45715);
nand U46667 (N_46667,N_45570,N_45926);
or U46668 (N_46668,N_45759,N_45487);
xor U46669 (N_46669,N_45394,N_45993);
xor U46670 (N_46670,N_45949,N_45827);
nor U46671 (N_46671,N_45112,N_45270);
and U46672 (N_46672,N_45602,N_45976);
xor U46673 (N_46673,N_45165,N_45592);
xor U46674 (N_46674,N_45774,N_45489);
and U46675 (N_46675,N_45366,N_45534);
nand U46676 (N_46676,N_45741,N_45539);
xnor U46677 (N_46677,N_45723,N_45222);
and U46678 (N_46678,N_45158,N_45826);
or U46679 (N_46679,N_45355,N_45975);
or U46680 (N_46680,N_45930,N_45303);
xnor U46681 (N_46681,N_45082,N_45694);
or U46682 (N_46682,N_45992,N_45527);
or U46683 (N_46683,N_45350,N_45555);
or U46684 (N_46684,N_45979,N_45729);
or U46685 (N_46685,N_45163,N_45618);
nand U46686 (N_46686,N_45964,N_45077);
or U46687 (N_46687,N_45124,N_45246);
nand U46688 (N_46688,N_45881,N_45883);
nand U46689 (N_46689,N_45583,N_45510);
or U46690 (N_46690,N_45413,N_45806);
xor U46691 (N_46691,N_45372,N_45480);
and U46692 (N_46692,N_45547,N_45137);
xnor U46693 (N_46693,N_45105,N_45700);
nand U46694 (N_46694,N_45895,N_45505);
nor U46695 (N_46695,N_45421,N_45818);
nor U46696 (N_46696,N_45002,N_45226);
nor U46697 (N_46697,N_45931,N_45138);
nor U46698 (N_46698,N_45829,N_45343);
nand U46699 (N_46699,N_45292,N_45331);
nor U46700 (N_46700,N_45097,N_45637);
nor U46701 (N_46701,N_45536,N_45972);
nor U46702 (N_46702,N_45360,N_45762);
nor U46703 (N_46703,N_45278,N_45021);
nor U46704 (N_46704,N_45539,N_45700);
or U46705 (N_46705,N_45250,N_45146);
xor U46706 (N_46706,N_45031,N_45212);
and U46707 (N_46707,N_45699,N_45759);
nor U46708 (N_46708,N_45597,N_45576);
or U46709 (N_46709,N_45228,N_45115);
nor U46710 (N_46710,N_45237,N_45637);
xnor U46711 (N_46711,N_45855,N_45360);
xnor U46712 (N_46712,N_45633,N_45750);
xor U46713 (N_46713,N_45426,N_45440);
or U46714 (N_46714,N_45843,N_45599);
xnor U46715 (N_46715,N_45258,N_45359);
nor U46716 (N_46716,N_45314,N_45660);
xor U46717 (N_46717,N_45728,N_45366);
and U46718 (N_46718,N_45388,N_45624);
nand U46719 (N_46719,N_45847,N_45267);
nor U46720 (N_46720,N_45388,N_45539);
and U46721 (N_46721,N_45278,N_45996);
nor U46722 (N_46722,N_45267,N_45450);
nor U46723 (N_46723,N_45863,N_45501);
or U46724 (N_46724,N_45679,N_45316);
nand U46725 (N_46725,N_45397,N_45999);
and U46726 (N_46726,N_45528,N_45167);
or U46727 (N_46727,N_45650,N_45183);
xor U46728 (N_46728,N_45891,N_45746);
xnor U46729 (N_46729,N_45801,N_45592);
nor U46730 (N_46730,N_45171,N_45217);
or U46731 (N_46731,N_45440,N_45693);
or U46732 (N_46732,N_45744,N_45948);
nand U46733 (N_46733,N_45404,N_45617);
nor U46734 (N_46734,N_45237,N_45816);
nor U46735 (N_46735,N_45873,N_45376);
and U46736 (N_46736,N_45745,N_45992);
nand U46737 (N_46737,N_45478,N_45268);
xnor U46738 (N_46738,N_45061,N_45870);
xor U46739 (N_46739,N_45472,N_45562);
xor U46740 (N_46740,N_45644,N_45272);
or U46741 (N_46741,N_45536,N_45993);
xor U46742 (N_46742,N_45138,N_45323);
and U46743 (N_46743,N_45799,N_45267);
xor U46744 (N_46744,N_45383,N_45411);
or U46745 (N_46745,N_45859,N_45801);
and U46746 (N_46746,N_45269,N_45196);
or U46747 (N_46747,N_45255,N_45493);
or U46748 (N_46748,N_45388,N_45685);
and U46749 (N_46749,N_45575,N_45929);
xor U46750 (N_46750,N_45761,N_45071);
and U46751 (N_46751,N_45385,N_45062);
or U46752 (N_46752,N_45465,N_45828);
or U46753 (N_46753,N_45827,N_45526);
nand U46754 (N_46754,N_45930,N_45184);
nor U46755 (N_46755,N_45288,N_45169);
nor U46756 (N_46756,N_45947,N_45662);
xnor U46757 (N_46757,N_45614,N_45971);
nor U46758 (N_46758,N_45309,N_45306);
and U46759 (N_46759,N_45557,N_45761);
nor U46760 (N_46760,N_45898,N_45516);
nand U46761 (N_46761,N_45716,N_45234);
and U46762 (N_46762,N_45968,N_45636);
or U46763 (N_46763,N_45726,N_45979);
xor U46764 (N_46764,N_45165,N_45340);
or U46765 (N_46765,N_45877,N_45710);
nand U46766 (N_46766,N_45984,N_45475);
xnor U46767 (N_46767,N_45383,N_45963);
or U46768 (N_46768,N_45075,N_45610);
nor U46769 (N_46769,N_45595,N_45486);
xnor U46770 (N_46770,N_45401,N_45957);
or U46771 (N_46771,N_45656,N_45996);
xnor U46772 (N_46772,N_45561,N_45042);
or U46773 (N_46773,N_45208,N_45294);
nor U46774 (N_46774,N_45070,N_45529);
nor U46775 (N_46775,N_45365,N_45292);
xnor U46776 (N_46776,N_45884,N_45992);
nor U46777 (N_46777,N_45636,N_45049);
and U46778 (N_46778,N_45397,N_45898);
nand U46779 (N_46779,N_45633,N_45731);
nand U46780 (N_46780,N_45317,N_45882);
nand U46781 (N_46781,N_45866,N_45758);
nand U46782 (N_46782,N_45179,N_45290);
or U46783 (N_46783,N_45895,N_45002);
nand U46784 (N_46784,N_45343,N_45514);
xor U46785 (N_46785,N_45042,N_45614);
and U46786 (N_46786,N_45528,N_45768);
nor U46787 (N_46787,N_45194,N_45077);
nand U46788 (N_46788,N_45950,N_45593);
xor U46789 (N_46789,N_45089,N_45392);
and U46790 (N_46790,N_45051,N_45223);
and U46791 (N_46791,N_45201,N_45137);
nand U46792 (N_46792,N_45362,N_45654);
or U46793 (N_46793,N_45785,N_45159);
nand U46794 (N_46794,N_45495,N_45477);
or U46795 (N_46795,N_45897,N_45616);
xnor U46796 (N_46796,N_45972,N_45158);
nand U46797 (N_46797,N_45561,N_45680);
or U46798 (N_46798,N_45938,N_45641);
nand U46799 (N_46799,N_45071,N_45676);
or U46800 (N_46800,N_45179,N_45191);
nor U46801 (N_46801,N_45172,N_45970);
or U46802 (N_46802,N_45198,N_45734);
nand U46803 (N_46803,N_45341,N_45928);
xor U46804 (N_46804,N_45850,N_45802);
and U46805 (N_46805,N_45780,N_45293);
and U46806 (N_46806,N_45567,N_45100);
nand U46807 (N_46807,N_45491,N_45932);
nand U46808 (N_46808,N_45411,N_45601);
or U46809 (N_46809,N_45354,N_45133);
and U46810 (N_46810,N_45451,N_45506);
xor U46811 (N_46811,N_45835,N_45745);
nand U46812 (N_46812,N_45979,N_45980);
and U46813 (N_46813,N_45153,N_45097);
xnor U46814 (N_46814,N_45466,N_45397);
nand U46815 (N_46815,N_45494,N_45007);
and U46816 (N_46816,N_45988,N_45644);
nand U46817 (N_46817,N_45389,N_45050);
nand U46818 (N_46818,N_45590,N_45211);
xnor U46819 (N_46819,N_45707,N_45645);
and U46820 (N_46820,N_45221,N_45428);
and U46821 (N_46821,N_45338,N_45678);
or U46822 (N_46822,N_45480,N_45428);
nand U46823 (N_46823,N_45680,N_45117);
and U46824 (N_46824,N_45438,N_45122);
nand U46825 (N_46825,N_45872,N_45505);
nand U46826 (N_46826,N_45228,N_45306);
or U46827 (N_46827,N_45460,N_45014);
nor U46828 (N_46828,N_45266,N_45426);
nor U46829 (N_46829,N_45015,N_45925);
or U46830 (N_46830,N_45193,N_45181);
nand U46831 (N_46831,N_45294,N_45347);
xor U46832 (N_46832,N_45720,N_45701);
and U46833 (N_46833,N_45900,N_45408);
nor U46834 (N_46834,N_45730,N_45010);
xor U46835 (N_46835,N_45726,N_45829);
nor U46836 (N_46836,N_45411,N_45043);
and U46837 (N_46837,N_45894,N_45840);
nor U46838 (N_46838,N_45876,N_45814);
and U46839 (N_46839,N_45850,N_45729);
xor U46840 (N_46840,N_45346,N_45039);
and U46841 (N_46841,N_45296,N_45336);
or U46842 (N_46842,N_45485,N_45051);
and U46843 (N_46843,N_45051,N_45896);
nor U46844 (N_46844,N_45356,N_45778);
and U46845 (N_46845,N_45279,N_45335);
nor U46846 (N_46846,N_45920,N_45036);
or U46847 (N_46847,N_45807,N_45067);
xor U46848 (N_46848,N_45919,N_45861);
xor U46849 (N_46849,N_45564,N_45820);
xnor U46850 (N_46850,N_45815,N_45557);
and U46851 (N_46851,N_45251,N_45402);
nor U46852 (N_46852,N_45932,N_45165);
or U46853 (N_46853,N_45199,N_45980);
xor U46854 (N_46854,N_45487,N_45278);
or U46855 (N_46855,N_45573,N_45625);
nor U46856 (N_46856,N_45090,N_45960);
nor U46857 (N_46857,N_45331,N_45540);
nor U46858 (N_46858,N_45297,N_45099);
nand U46859 (N_46859,N_45976,N_45047);
nand U46860 (N_46860,N_45048,N_45590);
or U46861 (N_46861,N_45302,N_45640);
nor U46862 (N_46862,N_45744,N_45648);
xor U46863 (N_46863,N_45928,N_45208);
xnor U46864 (N_46864,N_45943,N_45311);
and U46865 (N_46865,N_45716,N_45057);
nand U46866 (N_46866,N_45422,N_45637);
or U46867 (N_46867,N_45359,N_45464);
nand U46868 (N_46868,N_45872,N_45014);
nor U46869 (N_46869,N_45664,N_45736);
xnor U46870 (N_46870,N_45927,N_45384);
xor U46871 (N_46871,N_45495,N_45504);
or U46872 (N_46872,N_45399,N_45388);
nor U46873 (N_46873,N_45137,N_45172);
nor U46874 (N_46874,N_45271,N_45360);
xor U46875 (N_46875,N_45061,N_45010);
nand U46876 (N_46876,N_45261,N_45865);
nor U46877 (N_46877,N_45010,N_45278);
and U46878 (N_46878,N_45916,N_45043);
nand U46879 (N_46879,N_45559,N_45938);
nand U46880 (N_46880,N_45065,N_45328);
nor U46881 (N_46881,N_45206,N_45108);
or U46882 (N_46882,N_45314,N_45853);
xor U46883 (N_46883,N_45681,N_45223);
xnor U46884 (N_46884,N_45500,N_45380);
nand U46885 (N_46885,N_45636,N_45323);
xnor U46886 (N_46886,N_45627,N_45612);
nand U46887 (N_46887,N_45458,N_45093);
nand U46888 (N_46888,N_45183,N_45379);
xor U46889 (N_46889,N_45848,N_45113);
xor U46890 (N_46890,N_45006,N_45503);
and U46891 (N_46891,N_45879,N_45811);
xnor U46892 (N_46892,N_45454,N_45710);
xor U46893 (N_46893,N_45839,N_45422);
and U46894 (N_46894,N_45575,N_45397);
or U46895 (N_46895,N_45013,N_45407);
or U46896 (N_46896,N_45775,N_45587);
nor U46897 (N_46897,N_45349,N_45876);
or U46898 (N_46898,N_45522,N_45369);
xnor U46899 (N_46899,N_45735,N_45971);
and U46900 (N_46900,N_45861,N_45608);
and U46901 (N_46901,N_45012,N_45871);
xnor U46902 (N_46902,N_45627,N_45365);
or U46903 (N_46903,N_45098,N_45717);
nand U46904 (N_46904,N_45015,N_45530);
xnor U46905 (N_46905,N_45486,N_45287);
nand U46906 (N_46906,N_45506,N_45860);
xnor U46907 (N_46907,N_45095,N_45283);
and U46908 (N_46908,N_45376,N_45592);
and U46909 (N_46909,N_45323,N_45480);
or U46910 (N_46910,N_45599,N_45378);
and U46911 (N_46911,N_45297,N_45339);
or U46912 (N_46912,N_45645,N_45157);
nand U46913 (N_46913,N_45973,N_45286);
or U46914 (N_46914,N_45993,N_45122);
nor U46915 (N_46915,N_45993,N_45798);
nor U46916 (N_46916,N_45066,N_45268);
nor U46917 (N_46917,N_45479,N_45601);
nand U46918 (N_46918,N_45990,N_45417);
or U46919 (N_46919,N_45102,N_45114);
nor U46920 (N_46920,N_45380,N_45381);
or U46921 (N_46921,N_45555,N_45633);
nor U46922 (N_46922,N_45533,N_45860);
and U46923 (N_46923,N_45922,N_45547);
xnor U46924 (N_46924,N_45013,N_45148);
xor U46925 (N_46925,N_45340,N_45128);
or U46926 (N_46926,N_45704,N_45832);
and U46927 (N_46927,N_45064,N_45980);
xor U46928 (N_46928,N_45527,N_45893);
xnor U46929 (N_46929,N_45824,N_45541);
xnor U46930 (N_46930,N_45869,N_45835);
and U46931 (N_46931,N_45992,N_45680);
xor U46932 (N_46932,N_45289,N_45544);
or U46933 (N_46933,N_45628,N_45473);
xnor U46934 (N_46934,N_45393,N_45403);
xor U46935 (N_46935,N_45570,N_45650);
nor U46936 (N_46936,N_45085,N_45706);
and U46937 (N_46937,N_45239,N_45685);
or U46938 (N_46938,N_45045,N_45600);
nor U46939 (N_46939,N_45831,N_45193);
or U46940 (N_46940,N_45688,N_45689);
xnor U46941 (N_46941,N_45857,N_45346);
and U46942 (N_46942,N_45453,N_45409);
nand U46943 (N_46943,N_45983,N_45254);
nand U46944 (N_46944,N_45043,N_45167);
and U46945 (N_46945,N_45234,N_45731);
nand U46946 (N_46946,N_45075,N_45567);
or U46947 (N_46947,N_45366,N_45874);
nor U46948 (N_46948,N_45677,N_45772);
and U46949 (N_46949,N_45611,N_45005);
xor U46950 (N_46950,N_45180,N_45490);
or U46951 (N_46951,N_45240,N_45441);
xnor U46952 (N_46952,N_45010,N_45463);
xnor U46953 (N_46953,N_45513,N_45743);
or U46954 (N_46954,N_45005,N_45968);
xnor U46955 (N_46955,N_45571,N_45080);
and U46956 (N_46956,N_45756,N_45760);
or U46957 (N_46957,N_45161,N_45789);
nand U46958 (N_46958,N_45243,N_45932);
nor U46959 (N_46959,N_45070,N_45788);
nor U46960 (N_46960,N_45923,N_45443);
xor U46961 (N_46961,N_45206,N_45065);
nand U46962 (N_46962,N_45837,N_45047);
or U46963 (N_46963,N_45342,N_45218);
nand U46964 (N_46964,N_45979,N_45756);
nor U46965 (N_46965,N_45707,N_45038);
nor U46966 (N_46966,N_45983,N_45084);
nand U46967 (N_46967,N_45850,N_45764);
nor U46968 (N_46968,N_45125,N_45680);
or U46969 (N_46969,N_45943,N_45467);
nor U46970 (N_46970,N_45391,N_45427);
nand U46971 (N_46971,N_45157,N_45743);
and U46972 (N_46972,N_45624,N_45905);
nor U46973 (N_46973,N_45273,N_45179);
or U46974 (N_46974,N_45472,N_45196);
and U46975 (N_46975,N_45151,N_45544);
nand U46976 (N_46976,N_45214,N_45115);
nor U46977 (N_46977,N_45777,N_45224);
xor U46978 (N_46978,N_45455,N_45039);
or U46979 (N_46979,N_45906,N_45465);
or U46980 (N_46980,N_45840,N_45364);
nand U46981 (N_46981,N_45716,N_45276);
or U46982 (N_46982,N_45014,N_45283);
nand U46983 (N_46983,N_45887,N_45406);
xor U46984 (N_46984,N_45604,N_45343);
or U46985 (N_46985,N_45218,N_45263);
or U46986 (N_46986,N_45434,N_45496);
or U46987 (N_46987,N_45008,N_45920);
and U46988 (N_46988,N_45242,N_45626);
or U46989 (N_46989,N_45502,N_45141);
xor U46990 (N_46990,N_45446,N_45294);
nor U46991 (N_46991,N_45489,N_45373);
and U46992 (N_46992,N_45991,N_45246);
nand U46993 (N_46993,N_45945,N_45132);
xnor U46994 (N_46994,N_45713,N_45135);
or U46995 (N_46995,N_45521,N_45032);
and U46996 (N_46996,N_45528,N_45784);
and U46997 (N_46997,N_45866,N_45792);
nand U46998 (N_46998,N_45863,N_45813);
nand U46999 (N_46999,N_45629,N_45946);
nand U47000 (N_47000,N_46785,N_46445);
nand U47001 (N_47001,N_46519,N_46352);
nand U47002 (N_47002,N_46506,N_46198);
or U47003 (N_47003,N_46042,N_46769);
nand U47004 (N_47004,N_46789,N_46203);
or U47005 (N_47005,N_46383,N_46708);
nor U47006 (N_47006,N_46979,N_46053);
xnor U47007 (N_47007,N_46263,N_46653);
or U47008 (N_47008,N_46533,N_46786);
and U47009 (N_47009,N_46814,N_46110);
or U47010 (N_47010,N_46711,N_46036);
or U47011 (N_47011,N_46123,N_46562);
xnor U47012 (N_47012,N_46087,N_46799);
nor U47013 (N_47013,N_46540,N_46964);
and U47014 (N_47014,N_46116,N_46144);
and U47015 (N_47015,N_46176,N_46894);
or U47016 (N_47016,N_46621,N_46248);
nor U47017 (N_47017,N_46508,N_46566);
xor U47018 (N_47018,N_46570,N_46579);
nor U47019 (N_47019,N_46007,N_46730);
nand U47020 (N_47020,N_46732,N_46090);
xnor U47021 (N_47021,N_46738,N_46705);
and U47022 (N_47022,N_46867,N_46006);
nor U47023 (N_47023,N_46221,N_46495);
xor U47024 (N_47024,N_46490,N_46431);
xnor U47025 (N_47025,N_46780,N_46525);
nand U47026 (N_47026,N_46100,N_46948);
or U47027 (N_47027,N_46505,N_46312);
nor U47028 (N_47028,N_46073,N_46417);
xnor U47029 (N_47029,N_46832,N_46085);
nor U47030 (N_47030,N_46402,N_46603);
or U47031 (N_47031,N_46145,N_46464);
nand U47032 (N_47032,N_46324,N_46120);
nor U47033 (N_47033,N_46912,N_46457);
xnor U47034 (N_47034,N_46611,N_46432);
and U47035 (N_47035,N_46493,N_46152);
xnor U47036 (N_47036,N_46401,N_46368);
xnor U47037 (N_47037,N_46781,N_46960);
or U47038 (N_47038,N_46453,N_46716);
xnor U47039 (N_47039,N_46082,N_46807);
nand U47040 (N_47040,N_46925,N_46550);
nor U47041 (N_47041,N_46949,N_46450);
and U47042 (N_47042,N_46625,N_46749);
or U47043 (N_47043,N_46886,N_46530);
nand U47044 (N_47044,N_46397,N_46596);
and U47045 (N_47045,N_46788,N_46645);
or U47046 (N_47046,N_46808,N_46595);
and U47047 (N_47047,N_46454,N_46673);
or U47048 (N_47048,N_46816,N_46651);
nand U47049 (N_47049,N_46213,N_46900);
xnor U47050 (N_47050,N_46469,N_46794);
xor U47051 (N_47051,N_46336,N_46634);
or U47052 (N_47052,N_46823,N_46726);
or U47053 (N_47053,N_46989,N_46011);
nand U47054 (N_47054,N_46180,N_46486);
xor U47055 (N_47055,N_46833,N_46237);
nand U47056 (N_47056,N_46171,N_46154);
or U47057 (N_47057,N_46952,N_46970);
or U47058 (N_47058,N_46020,N_46284);
xnor U47059 (N_47059,N_46062,N_46172);
nor U47060 (N_47060,N_46386,N_46641);
and U47061 (N_47061,N_46555,N_46329);
or U47062 (N_47062,N_46366,N_46325);
or U47063 (N_47063,N_46390,N_46906);
nand U47064 (N_47064,N_46547,N_46019);
nor U47065 (N_47065,N_46442,N_46622);
and U47066 (N_47066,N_46648,N_46939);
xor U47067 (N_47067,N_46168,N_46323);
nor U47068 (N_47068,N_46755,N_46733);
xor U47069 (N_47069,N_46911,N_46838);
nor U47070 (N_47070,N_46182,N_46690);
nand U47071 (N_47071,N_46276,N_46600);
nand U47072 (N_47072,N_46111,N_46881);
or U47073 (N_47073,N_46029,N_46360);
and U47074 (N_47074,N_46935,N_46063);
or U47075 (N_47075,N_46338,N_46872);
nand U47076 (N_47076,N_46700,N_46423);
nand U47077 (N_47077,N_46689,N_46660);
or U47078 (N_47078,N_46984,N_46656);
xnor U47079 (N_47079,N_46850,N_46267);
and U47080 (N_47080,N_46847,N_46305);
nand U47081 (N_47081,N_46842,N_46617);
and U47082 (N_47082,N_46688,N_46418);
xnor U47083 (N_47083,N_46956,N_46633);
nand U47084 (N_47084,N_46797,N_46941);
nor U47085 (N_47085,N_46008,N_46005);
or U47086 (N_47086,N_46119,N_46370);
nor U47087 (N_47087,N_46723,N_46015);
or U47088 (N_47088,N_46387,N_46942);
or U47089 (N_47089,N_46576,N_46040);
or U47090 (N_47090,N_46848,N_46016);
or U47091 (N_47091,N_46902,N_46452);
and U47092 (N_47092,N_46420,N_46861);
nor U47093 (N_47093,N_46114,N_46663);
xnor U47094 (N_47094,N_46434,N_46404);
or U47095 (N_47095,N_46410,N_46300);
and U47096 (N_47096,N_46281,N_46422);
xnor U47097 (N_47097,N_46269,N_46717);
nand U47098 (N_47098,N_46943,N_46279);
nor U47099 (N_47099,N_46936,N_46855);
xor U47100 (N_47100,N_46270,N_46715);
and U47101 (N_47101,N_46129,N_46577);
and U47102 (N_47102,N_46985,N_46548);
and U47103 (N_47103,N_46558,N_46262);
nor U47104 (N_47104,N_46871,N_46542);
and U47105 (N_47105,N_46544,N_46583);
nor U47106 (N_47106,N_46585,N_46578);
xor U47107 (N_47107,N_46181,N_46398);
nand U47108 (N_47108,N_46987,N_46869);
or U47109 (N_47109,N_46817,N_46408);
nand U47110 (N_47110,N_46208,N_46158);
or U47111 (N_47111,N_46148,N_46271);
xor U47112 (N_47112,N_46125,N_46889);
nor U47113 (N_47113,N_46677,N_46374);
and U47114 (N_47114,N_46497,N_46591);
nand U47115 (N_47115,N_46975,N_46244);
and U47116 (N_47116,N_46257,N_46779);
xnor U47117 (N_47117,N_46230,N_46680);
and U47118 (N_47118,N_46350,N_46915);
and U47119 (N_47119,N_46013,N_46655);
nor U47120 (N_47120,N_46793,N_46295);
or U47121 (N_47121,N_46862,N_46783);
nor U47122 (N_47122,N_46274,N_46472);
or U47123 (N_47123,N_46031,N_46130);
nand U47124 (N_47124,N_46938,N_46156);
or U47125 (N_47125,N_46344,N_46170);
and U47126 (N_47126,N_46478,N_46974);
and U47127 (N_47127,N_46612,N_46299);
or U47128 (N_47128,N_46384,N_46986);
nor U47129 (N_47129,N_46804,N_46509);
xor U47130 (N_47130,N_46455,N_46223);
or U47131 (N_47131,N_46630,N_46863);
nor U47132 (N_47132,N_46242,N_46033);
xnor U47133 (N_47133,N_46065,N_46475);
and U47134 (N_47134,N_46801,N_46777);
and U47135 (N_47135,N_46534,N_46724);
nor U47136 (N_47136,N_46843,N_46860);
xnor U47137 (N_47137,N_46400,N_46205);
or U47138 (N_47138,N_46683,N_46999);
or U47139 (N_47139,N_46880,N_46907);
nand U47140 (N_47140,N_46997,N_46414);
nor U47141 (N_47141,N_46055,N_46030);
and U47142 (N_47142,N_46758,N_46131);
and U47143 (N_47143,N_46520,N_46235);
nor U47144 (N_47144,N_46895,N_46415);
nor U47145 (N_47145,N_46760,N_46892);
or U47146 (N_47146,N_46538,N_46927);
nand U47147 (N_47147,N_46481,N_46682);
or U47148 (N_47148,N_46694,N_46084);
and U47149 (N_47149,N_46845,N_46865);
xor U47150 (N_47150,N_46669,N_46365);
nand U47151 (N_47151,N_46037,N_46759);
and U47152 (N_47152,N_46396,N_46896);
nor U47153 (N_47153,N_46304,N_46095);
xor U47154 (N_47154,N_46851,N_46291);
nand U47155 (N_47155,N_46479,N_46664);
nand U47156 (N_47156,N_46640,N_46297);
xnor U47157 (N_47157,N_46381,N_46772);
nor U47158 (N_47158,N_46092,N_46556);
nand U47159 (N_47159,N_46606,N_46972);
nand U47160 (N_47160,N_46592,N_46990);
or U47161 (N_47161,N_46736,N_46018);
nand U47162 (N_47162,N_46275,N_46311);
nor U47163 (N_47163,N_46194,N_46501);
and U47164 (N_47164,N_46255,N_46891);
and U47165 (N_47165,N_46768,N_46955);
nand U47166 (N_47166,N_46245,N_46572);
and U47167 (N_47167,N_46601,N_46340);
nor U47168 (N_47168,N_46916,N_46128);
nor U47169 (N_47169,N_46070,N_46476);
xnor U47170 (N_47170,N_46764,N_46272);
nand U47171 (N_47171,N_46060,N_46320);
or U47172 (N_47172,N_46670,N_46686);
nand U47173 (N_47173,N_46593,N_46588);
xor U47174 (N_47174,N_46347,N_46977);
or U47175 (N_47175,N_46098,N_46959);
xnor U47176 (N_47176,N_46504,N_46000);
xor U47177 (N_47177,N_46898,N_46824);
and U47178 (N_47178,N_46088,N_46623);
and U47179 (N_47179,N_46214,N_46189);
xor U47180 (N_47180,N_46602,N_46810);
xnor U47181 (N_47181,N_46049,N_46526);
and U47182 (N_47182,N_46587,N_46458);
and U47183 (N_47183,N_46157,N_46613);
or U47184 (N_47184,N_46259,N_46568);
nand U47185 (N_47185,N_46903,N_46210);
nand U47186 (N_47186,N_46913,N_46932);
and U47187 (N_47187,N_46962,N_46953);
or U47188 (N_47188,N_46028,N_46460);
nand U47189 (N_47189,N_46358,N_46691);
and U47190 (N_47190,N_46561,N_46200);
nor U47191 (N_47191,N_46830,N_46122);
or U47192 (N_47192,N_46322,N_46333);
or U47193 (N_47193,N_46888,N_46190);
and U47194 (N_47194,N_46193,N_46106);
nor U47195 (N_47195,N_46254,N_46175);
or U47196 (N_47196,N_46108,N_46598);
or U47197 (N_47197,N_46039,N_46767);
xor U47198 (N_47198,N_46136,N_46341);
or U47199 (N_47199,N_46061,N_46674);
xor U47200 (N_47200,N_46419,N_46004);
and U47201 (N_47201,N_46032,N_46580);
nand U47202 (N_47202,N_46864,N_46474);
nor U47203 (N_47203,N_46770,N_46775);
nor U47204 (N_47204,N_46695,N_46626);
or U47205 (N_47205,N_46192,N_46380);
nand U47206 (N_47206,N_46378,N_46307);
or U47207 (N_47207,N_46806,N_46346);
and U47208 (N_47208,N_46224,N_46468);
nand U47209 (N_47209,N_46294,N_46620);
xor U47210 (N_47210,N_46355,N_46910);
xor U47211 (N_47211,N_46107,N_46051);
xnor U47212 (N_47212,N_46251,N_46776);
xor U47213 (N_47213,N_46043,N_46480);
nand U47214 (N_47214,N_46405,N_46206);
and U47215 (N_47215,N_46687,N_46348);
and U47216 (N_47216,N_46052,N_46980);
nor U47217 (N_47217,N_46316,N_46236);
nand U47218 (N_47218,N_46289,N_46115);
nor U47219 (N_47219,N_46126,N_46513);
nand U47220 (N_47220,N_46188,N_46089);
and U47221 (N_47221,N_46047,N_46283);
and U47222 (N_47222,N_46345,N_46109);
and U47223 (N_47223,N_46652,N_46662);
and U47224 (N_47224,N_46151,N_46826);
and U47225 (N_47225,N_46339,N_46083);
and U47226 (N_47226,N_46335,N_46080);
and U47227 (N_47227,N_46564,N_46721);
and U47228 (N_47228,N_46812,N_46491);
or U47229 (N_47229,N_46178,N_46787);
and U47230 (N_47230,N_46743,N_46071);
nor U47231 (N_47231,N_46658,N_46800);
xnor U47232 (N_47232,N_46437,N_46642);
xnor U47233 (N_47233,N_46565,N_46228);
or U47234 (N_47234,N_46522,N_46908);
and U47235 (N_47235,N_46958,N_46961);
or U47236 (N_47236,N_46427,N_46334);
or U47237 (N_47237,N_46449,N_46649);
nand U47238 (N_47238,N_46499,N_46866);
nor U47239 (N_47239,N_46978,N_46552);
nand U47240 (N_47240,N_46597,N_46536);
nor U47241 (N_47241,N_46516,N_46003);
nor U47242 (N_47242,N_46357,N_46142);
nor U47243 (N_47243,N_46412,N_46354);
xnor U47244 (N_47244,N_46132,N_46153);
nor U47245 (N_47245,N_46310,N_46735);
or U47246 (N_47246,N_46435,N_46429);
xor U47247 (N_47247,N_46027,N_46009);
xnor U47248 (N_47248,N_46976,N_46921);
nand U47249 (N_47249,N_46059,N_46696);
nand U47250 (N_47250,N_46337,N_46933);
and U47251 (N_47251,N_46146,N_46757);
and U47252 (N_47252,N_46951,N_46438);
and U47253 (N_47253,N_46638,N_46155);
xor U47254 (N_47254,N_46928,N_46240);
and U47255 (N_47255,N_46376,N_46492);
nor U47256 (N_47256,N_46829,N_46367);
nand U47257 (N_47257,N_46433,N_46639);
and U47258 (N_47258,N_46046,N_46258);
xnor U47259 (N_47259,N_46950,N_46278);
xnor U47260 (N_47260,N_46720,N_46466);
nor U47261 (N_47261,N_46428,N_46922);
and U47262 (N_47262,N_46543,N_46097);
and U47263 (N_47263,N_46118,N_46774);
xor U47264 (N_47264,N_46728,N_46233);
xor U47265 (N_47265,N_46795,N_46559);
nand U47266 (N_47266,N_46002,N_46313);
or U47267 (N_47267,N_46571,N_46841);
and U47268 (N_47268,N_46684,N_46856);
nand U47269 (N_47269,N_46239,N_46447);
nand U47270 (N_47270,N_46919,N_46615);
nor U47271 (N_47271,N_46605,N_46105);
nor U47272 (N_47272,N_46388,N_46840);
nor U47273 (N_47273,N_46463,N_46671);
nand U47274 (N_47274,N_46072,N_46676);
xor U47275 (N_47275,N_46058,N_46470);
xnor U47276 (N_47276,N_46748,N_46822);
or U47277 (N_47277,N_46803,N_46854);
or U47278 (N_47278,N_46483,N_46563);
nand U47279 (N_47279,N_46746,N_46424);
nand U47280 (N_47280,N_46740,N_46878);
nand U47281 (N_47281,N_46298,N_46331);
nor U47282 (N_47282,N_46440,N_46473);
and U47283 (N_47283,N_46992,N_46859);
nand U47284 (N_47284,N_46394,N_46837);
and U47285 (N_47285,N_46609,N_46675);
nand U47286 (N_47286,N_46379,N_46988);
and U47287 (N_47287,N_46503,N_46698);
or U47288 (N_47288,N_46582,N_46624);
nor U47289 (N_47289,N_46280,N_46288);
nor U47290 (N_47290,N_46947,N_46968);
or U47291 (N_47291,N_46104,N_46586);
nor U47292 (N_47292,N_46186,N_46818);
or U47293 (N_47293,N_46426,N_46870);
and U47294 (N_47294,N_46025,N_46931);
and U47295 (N_47295,N_46103,N_46995);
xor U47296 (N_47296,N_46372,N_46375);
and U47297 (N_47297,N_46904,N_46231);
nor U47298 (N_47298,N_46608,N_46135);
xnor U47299 (N_47299,N_46584,N_46884);
xor U47300 (N_47300,N_46629,N_46195);
nor U47301 (N_47301,N_46734,N_46858);
nand U47302 (N_47302,N_46782,N_46117);
xor U47303 (N_47303,N_46754,N_46981);
and U47304 (N_47304,N_46389,N_46517);
nor U47305 (N_47305,N_46706,N_46177);
nand U47306 (N_47306,N_46569,N_46050);
nor U47307 (N_47307,N_46849,N_46184);
and U47308 (N_47308,N_46187,N_46202);
or U47309 (N_47309,N_46277,N_46699);
and U47310 (N_47310,N_46727,N_46885);
nand U47311 (N_47311,N_46197,N_46646);
xnor U47312 (N_47312,N_46714,N_46436);
nand U47313 (N_47313,N_46531,N_46139);
and U47314 (N_47314,N_46439,N_46361);
nand U47315 (N_47315,N_46247,N_46141);
or U47316 (N_47316,N_46731,N_46409);
or U47317 (N_47317,N_46659,N_46668);
or U47318 (N_47318,N_46074,N_46369);
and U47319 (N_47319,N_46930,N_46166);
xnor U47320 (N_47320,N_46905,N_46994);
or U47321 (N_47321,N_46012,N_46332);
and U47322 (N_47322,N_46619,N_46737);
nor U47323 (N_47323,N_46512,N_46326);
nor U47324 (N_47324,N_46678,N_46140);
or U47325 (N_47325,N_46725,N_46893);
or U47326 (N_47326,N_46399,N_46599);
or U47327 (N_47327,N_46147,N_46234);
nor U47328 (N_47328,N_46742,N_46616);
or U47329 (N_47329,N_46448,N_46351);
or U47330 (N_47330,N_46553,N_46207);
nand U47331 (N_47331,N_46484,N_46243);
and U47332 (N_47332,N_46001,N_46253);
nand U47333 (N_47333,N_46343,N_46229);
nor U47334 (N_47334,N_46353,N_46461);
nand U47335 (N_47335,N_46196,N_46441);
nor U47336 (N_47336,N_46496,N_46672);
nand U47337 (N_47337,N_46926,N_46024);
xnor U47338 (N_47338,N_46741,N_46167);
xnor U47339 (N_47339,N_46308,N_46637);
nand U47340 (N_47340,N_46707,N_46765);
and U47341 (N_47341,N_46518,N_46963);
nand U47342 (N_47342,N_46996,N_46756);
nor U47343 (N_47343,N_46303,N_46430);
xnor U47344 (N_47344,N_46101,N_46138);
nand U47345 (N_47345,N_46831,N_46590);
nor U47346 (N_47346,N_46681,N_46967);
or U47347 (N_47347,N_46853,N_46068);
nand U47348 (N_47348,N_46957,N_46163);
xor U47349 (N_47349,N_46798,N_46382);
xor U47350 (N_47350,N_46567,N_46077);
or U47351 (N_47351,N_46834,N_46546);
nand U47352 (N_47352,N_46502,N_46041);
or U47353 (N_47353,N_46747,N_46667);
nand U47354 (N_47354,N_46614,N_46796);
or U47355 (N_47355,N_46969,N_46581);
and U47356 (N_47356,N_46456,N_46521);
or U47357 (N_47357,N_46709,N_46554);
or U47358 (N_47358,N_46159,N_46589);
nand U47359 (N_47359,N_46879,N_46252);
and U47360 (N_47360,N_46852,N_46778);
and U47361 (N_47361,N_46647,N_46017);
nand U47362 (N_47362,N_46679,N_46643);
nand U47363 (N_47363,N_46945,N_46446);
or U47364 (N_47364,N_46791,N_46594);
xor U47365 (N_47365,N_46661,N_46314);
and U47366 (N_47366,N_46890,N_46371);
or U47367 (N_47367,N_46693,N_46809);
or U47368 (N_47368,N_46330,N_46815);
nor U47369 (N_47369,N_46532,N_46462);
nand U47370 (N_47370,N_46421,N_46607);
nor U47371 (N_47371,N_46983,N_46813);
nand U47372 (N_47372,N_46160,N_46821);
nand U47373 (N_47373,N_46836,N_46739);
xor U47374 (N_47374,N_46477,N_46164);
nand U47375 (N_47375,N_46215,N_46318);
and U47376 (N_47376,N_46287,N_46574);
or U47377 (N_47377,N_46752,N_46296);
or U47378 (N_47378,N_46882,N_46811);
and U47379 (N_47379,N_46056,N_46745);
and U47380 (N_47380,N_46704,N_46183);
xnor U47381 (N_47381,N_46363,N_46857);
xnor U47382 (N_47382,N_46161,N_46222);
xnor U47383 (N_47383,N_46362,N_46549);
nor U47384 (N_47384,N_46321,N_46887);
nor U47385 (N_47385,N_46185,N_46685);
xor U47386 (N_47386,N_46666,N_46744);
nand U47387 (N_47387,N_46137,N_46573);
and U47388 (N_47388,N_46249,N_46524);
nand U47389 (N_47389,N_46225,N_46628);
and U47390 (N_47390,N_46523,N_46064);
nor U47391 (N_47391,N_46527,N_46306);
nor U47392 (N_47392,N_46026,N_46819);
or U47393 (N_47393,N_46873,N_46124);
or U47394 (N_47394,N_46844,N_46407);
and U47395 (N_47395,N_46529,N_46766);
xnor U47396 (N_47396,N_46048,N_46557);
and U47397 (N_47397,N_46246,N_46971);
or U47398 (N_47398,N_46165,N_46924);
or U47399 (N_47399,N_46471,N_46729);
nand U47400 (N_47400,N_46069,N_46023);
xnor U47401 (N_47401,N_46217,N_46067);
nor U47402 (N_47402,N_46846,N_46162);
or U47403 (N_47403,N_46909,N_46150);
nor U47404 (N_47404,N_46507,N_46373);
and U47405 (N_47405,N_46697,N_46459);
and U47406 (N_47406,N_46514,N_46763);
nand U47407 (N_47407,N_46790,N_46965);
and U47408 (N_47408,N_46075,N_46883);
or U47409 (N_47409,N_46038,N_46081);
xor U47410 (N_47410,N_46511,N_46954);
xor U47411 (N_47411,N_46631,N_46057);
and U47412 (N_47412,N_46485,N_46899);
and U47413 (N_47413,N_46293,N_46875);
and U47414 (N_47414,N_46839,N_46391);
and U47415 (N_47415,N_46292,N_46143);
xnor U47416 (N_47416,N_46635,N_46266);
and U47417 (N_47417,N_46528,N_46500);
nand U47418 (N_47418,N_46537,N_46218);
nand U47419 (N_47419,N_46966,N_46487);
and U47420 (N_47420,N_46359,N_46627);
and U47421 (N_47421,N_46998,N_46022);
nand U47422 (N_47422,N_46920,N_46703);
xnor U47423 (N_47423,N_46174,N_46250);
nand U47424 (N_47424,N_46632,N_46494);
and U47425 (N_47425,N_46692,N_46403);
nor U47426 (N_47426,N_46636,N_46086);
and U47427 (N_47427,N_46535,N_46282);
xnor U47428 (N_47428,N_46268,N_46179);
nand U47429 (N_47429,N_46877,N_46465);
nor U47430 (N_47430,N_46771,N_46078);
nand U47431 (N_47431,N_46260,N_46551);
or U47432 (N_47432,N_46993,N_46079);
or U47433 (N_47433,N_46918,N_46356);
or U47434 (N_47434,N_46315,N_46169);
xnor U47435 (N_47435,N_46488,N_46991);
or U47436 (N_47436,N_46385,N_46076);
and U47437 (N_47437,N_46393,N_46946);
and U47438 (N_47438,N_46377,N_46874);
xor U47439 (N_47439,N_46761,N_46868);
nand U47440 (N_47440,N_46451,N_46710);
or U47441 (N_47441,N_46876,N_46014);
and U47442 (N_47442,N_46498,N_46545);
nor U47443 (N_47443,N_46201,N_46515);
xnor U47444 (N_47444,N_46784,N_46121);
or U47445 (N_47445,N_46364,N_46094);
or U47446 (N_47446,N_46897,N_46191);
xor U47447 (N_47447,N_46173,N_46657);
or U47448 (N_47448,N_46718,N_46113);
or U47449 (N_47449,N_46406,N_46828);
nor U47450 (N_47450,N_46035,N_46982);
or U47451 (N_47451,N_46560,N_46940);
nand U47452 (N_47452,N_46091,N_46820);
nand U47453 (N_47453,N_46219,N_46149);
xor U47454 (N_47454,N_46238,N_46216);
nor U47455 (N_47455,N_46973,N_46204);
and U47456 (N_47456,N_46917,N_46273);
nand U47457 (N_47457,N_46342,N_46328);
nand U47458 (N_47458,N_46066,N_46241);
nand U47459 (N_47459,N_46618,N_46701);
nor U47460 (N_47460,N_46209,N_46127);
nor U47461 (N_47461,N_46712,N_46264);
or U47462 (N_47462,N_46226,N_46301);
nor U47463 (N_47463,N_46914,N_46411);
nor U47464 (N_47464,N_46654,N_46575);
nor U47465 (N_47465,N_46290,N_46792);
and U47466 (N_47466,N_46302,N_46650);
nand U47467 (N_47467,N_46034,N_46349);
xnor U47468 (N_47468,N_46610,N_46199);
nor U47469 (N_47469,N_46112,N_46702);
xor U47470 (N_47470,N_46416,N_46443);
xor U47471 (N_47471,N_46539,N_46762);
nor U47472 (N_47472,N_46934,N_46265);
nand U47473 (N_47473,N_46750,N_46327);
nand U47474 (N_47474,N_46054,N_46232);
nand U47475 (N_47475,N_46467,N_46444);
or U47476 (N_47476,N_46261,N_46482);
nand U47477 (N_47477,N_46644,N_46773);
xnor U47478 (N_47478,N_46319,N_46044);
nor U47479 (N_47479,N_46827,N_46665);
and U47480 (N_47480,N_46802,N_46929);
or U47481 (N_47481,N_46021,N_46093);
nor U47482 (N_47482,N_46413,N_46102);
xnor U47483 (N_47483,N_46753,N_46309);
nor U47484 (N_47484,N_46133,N_46256);
xor U47485 (N_47485,N_46395,N_46489);
or U47486 (N_47486,N_46212,N_46286);
and U47487 (N_47487,N_46010,N_46134);
or U47488 (N_47488,N_46713,N_46285);
xnor U47489 (N_47489,N_46045,N_46805);
or U47490 (N_47490,N_46719,N_46751);
or U47491 (N_47491,N_46835,N_46901);
nand U47492 (N_47492,N_46510,N_46425);
or U47493 (N_47493,N_46944,N_46227);
xnor U47494 (N_47494,N_46937,N_46099);
nand U47495 (N_47495,N_46722,N_46392);
xor U47496 (N_47496,N_46317,N_46211);
nand U47497 (N_47497,N_46923,N_46541);
nand U47498 (N_47498,N_46825,N_46220);
or U47499 (N_47499,N_46604,N_46096);
and U47500 (N_47500,N_46553,N_46865);
xor U47501 (N_47501,N_46609,N_46672);
xor U47502 (N_47502,N_46700,N_46660);
nand U47503 (N_47503,N_46038,N_46696);
or U47504 (N_47504,N_46292,N_46796);
xnor U47505 (N_47505,N_46017,N_46245);
nor U47506 (N_47506,N_46586,N_46256);
or U47507 (N_47507,N_46213,N_46352);
nor U47508 (N_47508,N_46455,N_46895);
nand U47509 (N_47509,N_46038,N_46586);
nand U47510 (N_47510,N_46568,N_46340);
or U47511 (N_47511,N_46673,N_46427);
nor U47512 (N_47512,N_46186,N_46297);
and U47513 (N_47513,N_46134,N_46018);
and U47514 (N_47514,N_46214,N_46534);
and U47515 (N_47515,N_46899,N_46725);
or U47516 (N_47516,N_46336,N_46257);
and U47517 (N_47517,N_46462,N_46604);
and U47518 (N_47518,N_46744,N_46402);
xnor U47519 (N_47519,N_46662,N_46415);
and U47520 (N_47520,N_46002,N_46680);
nand U47521 (N_47521,N_46228,N_46116);
xnor U47522 (N_47522,N_46561,N_46448);
and U47523 (N_47523,N_46571,N_46560);
xnor U47524 (N_47524,N_46854,N_46758);
xnor U47525 (N_47525,N_46174,N_46746);
xor U47526 (N_47526,N_46001,N_46421);
xnor U47527 (N_47527,N_46254,N_46677);
and U47528 (N_47528,N_46794,N_46789);
nor U47529 (N_47529,N_46956,N_46096);
nor U47530 (N_47530,N_46982,N_46828);
nor U47531 (N_47531,N_46635,N_46576);
nor U47532 (N_47532,N_46605,N_46998);
xnor U47533 (N_47533,N_46039,N_46656);
xnor U47534 (N_47534,N_46670,N_46327);
and U47535 (N_47535,N_46388,N_46935);
nand U47536 (N_47536,N_46253,N_46727);
nor U47537 (N_47537,N_46232,N_46000);
xnor U47538 (N_47538,N_46144,N_46785);
nor U47539 (N_47539,N_46181,N_46035);
or U47540 (N_47540,N_46613,N_46040);
xnor U47541 (N_47541,N_46903,N_46816);
nand U47542 (N_47542,N_46678,N_46172);
and U47543 (N_47543,N_46337,N_46074);
and U47544 (N_47544,N_46978,N_46504);
xnor U47545 (N_47545,N_46380,N_46333);
and U47546 (N_47546,N_46904,N_46417);
nand U47547 (N_47547,N_46724,N_46529);
nor U47548 (N_47548,N_46369,N_46613);
or U47549 (N_47549,N_46496,N_46107);
nor U47550 (N_47550,N_46406,N_46019);
xnor U47551 (N_47551,N_46129,N_46362);
nor U47552 (N_47552,N_46740,N_46260);
or U47553 (N_47553,N_46193,N_46469);
and U47554 (N_47554,N_46219,N_46173);
and U47555 (N_47555,N_46821,N_46437);
nor U47556 (N_47556,N_46824,N_46755);
nand U47557 (N_47557,N_46053,N_46086);
xor U47558 (N_47558,N_46799,N_46195);
or U47559 (N_47559,N_46167,N_46385);
and U47560 (N_47560,N_46252,N_46506);
nor U47561 (N_47561,N_46925,N_46180);
or U47562 (N_47562,N_46806,N_46815);
nor U47563 (N_47563,N_46230,N_46257);
xor U47564 (N_47564,N_46839,N_46143);
xnor U47565 (N_47565,N_46267,N_46105);
nand U47566 (N_47566,N_46875,N_46630);
and U47567 (N_47567,N_46468,N_46564);
xor U47568 (N_47568,N_46779,N_46088);
and U47569 (N_47569,N_46158,N_46795);
and U47570 (N_47570,N_46025,N_46405);
nand U47571 (N_47571,N_46570,N_46315);
and U47572 (N_47572,N_46821,N_46287);
or U47573 (N_47573,N_46792,N_46031);
or U47574 (N_47574,N_46732,N_46367);
xor U47575 (N_47575,N_46950,N_46623);
nor U47576 (N_47576,N_46487,N_46179);
or U47577 (N_47577,N_46991,N_46466);
nand U47578 (N_47578,N_46244,N_46497);
or U47579 (N_47579,N_46439,N_46882);
nand U47580 (N_47580,N_46697,N_46017);
nand U47581 (N_47581,N_46275,N_46550);
and U47582 (N_47582,N_46305,N_46474);
and U47583 (N_47583,N_46964,N_46485);
nor U47584 (N_47584,N_46214,N_46549);
nor U47585 (N_47585,N_46291,N_46378);
and U47586 (N_47586,N_46595,N_46883);
or U47587 (N_47587,N_46238,N_46180);
or U47588 (N_47588,N_46075,N_46377);
and U47589 (N_47589,N_46735,N_46329);
or U47590 (N_47590,N_46938,N_46015);
xor U47591 (N_47591,N_46527,N_46349);
nand U47592 (N_47592,N_46320,N_46945);
nor U47593 (N_47593,N_46966,N_46387);
nor U47594 (N_47594,N_46914,N_46305);
nand U47595 (N_47595,N_46287,N_46820);
xnor U47596 (N_47596,N_46173,N_46843);
and U47597 (N_47597,N_46032,N_46381);
xor U47598 (N_47598,N_46091,N_46664);
or U47599 (N_47599,N_46051,N_46918);
nor U47600 (N_47600,N_46703,N_46190);
nand U47601 (N_47601,N_46905,N_46555);
or U47602 (N_47602,N_46253,N_46719);
or U47603 (N_47603,N_46856,N_46928);
nor U47604 (N_47604,N_46329,N_46410);
and U47605 (N_47605,N_46291,N_46061);
xnor U47606 (N_47606,N_46456,N_46339);
and U47607 (N_47607,N_46366,N_46296);
xor U47608 (N_47608,N_46308,N_46876);
xor U47609 (N_47609,N_46250,N_46952);
xor U47610 (N_47610,N_46710,N_46121);
or U47611 (N_47611,N_46022,N_46997);
nand U47612 (N_47612,N_46035,N_46264);
or U47613 (N_47613,N_46064,N_46699);
nor U47614 (N_47614,N_46521,N_46770);
nor U47615 (N_47615,N_46883,N_46290);
nand U47616 (N_47616,N_46591,N_46411);
xor U47617 (N_47617,N_46339,N_46302);
or U47618 (N_47618,N_46312,N_46805);
or U47619 (N_47619,N_46181,N_46566);
and U47620 (N_47620,N_46290,N_46878);
nor U47621 (N_47621,N_46805,N_46201);
and U47622 (N_47622,N_46024,N_46734);
nand U47623 (N_47623,N_46271,N_46664);
or U47624 (N_47624,N_46900,N_46449);
xnor U47625 (N_47625,N_46219,N_46201);
nor U47626 (N_47626,N_46665,N_46747);
nand U47627 (N_47627,N_46289,N_46924);
and U47628 (N_47628,N_46633,N_46654);
nor U47629 (N_47629,N_46528,N_46181);
or U47630 (N_47630,N_46505,N_46450);
nor U47631 (N_47631,N_46624,N_46283);
or U47632 (N_47632,N_46559,N_46742);
xnor U47633 (N_47633,N_46230,N_46866);
nand U47634 (N_47634,N_46513,N_46091);
xnor U47635 (N_47635,N_46281,N_46291);
and U47636 (N_47636,N_46599,N_46327);
nor U47637 (N_47637,N_46553,N_46222);
and U47638 (N_47638,N_46278,N_46023);
nand U47639 (N_47639,N_46050,N_46448);
nor U47640 (N_47640,N_46089,N_46076);
nand U47641 (N_47641,N_46516,N_46521);
nand U47642 (N_47642,N_46458,N_46507);
xor U47643 (N_47643,N_46191,N_46330);
nand U47644 (N_47644,N_46946,N_46816);
or U47645 (N_47645,N_46175,N_46138);
nor U47646 (N_47646,N_46377,N_46296);
and U47647 (N_47647,N_46898,N_46517);
and U47648 (N_47648,N_46968,N_46854);
nor U47649 (N_47649,N_46101,N_46239);
nor U47650 (N_47650,N_46626,N_46072);
xnor U47651 (N_47651,N_46326,N_46641);
nor U47652 (N_47652,N_46801,N_46152);
and U47653 (N_47653,N_46759,N_46131);
nand U47654 (N_47654,N_46673,N_46809);
xor U47655 (N_47655,N_46911,N_46586);
nand U47656 (N_47656,N_46832,N_46365);
or U47657 (N_47657,N_46820,N_46256);
nand U47658 (N_47658,N_46130,N_46696);
xor U47659 (N_47659,N_46130,N_46297);
and U47660 (N_47660,N_46674,N_46559);
xor U47661 (N_47661,N_46747,N_46298);
nand U47662 (N_47662,N_46438,N_46048);
nand U47663 (N_47663,N_46476,N_46648);
xor U47664 (N_47664,N_46142,N_46392);
and U47665 (N_47665,N_46312,N_46190);
xnor U47666 (N_47666,N_46770,N_46357);
nor U47667 (N_47667,N_46092,N_46656);
xnor U47668 (N_47668,N_46628,N_46804);
nand U47669 (N_47669,N_46405,N_46949);
and U47670 (N_47670,N_46879,N_46449);
xor U47671 (N_47671,N_46378,N_46449);
nor U47672 (N_47672,N_46629,N_46855);
nand U47673 (N_47673,N_46479,N_46928);
nand U47674 (N_47674,N_46356,N_46464);
xnor U47675 (N_47675,N_46840,N_46673);
or U47676 (N_47676,N_46705,N_46116);
or U47677 (N_47677,N_46812,N_46011);
xnor U47678 (N_47678,N_46096,N_46655);
nand U47679 (N_47679,N_46441,N_46134);
xor U47680 (N_47680,N_46898,N_46187);
nor U47681 (N_47681,N_46592,N_46814);
nand U47682 (N_47682,N_46728,N_46178);
nor U47683 (N_47683,N_46523,N_46444);
or U47684 (N_47684,N_46879,N_46797);
nand U47685 (N_47685,N_46195,N_46684);
and U47686 (N_47686,N_46015,N_46764);
and U47687 (N_47687,N_46962,N_46031);
nor U47688 (N_47688,N_46881,N_46812);
xnor U47689 (N_47689,N_46456,N_46276);
or U47690 (N_47690,N_46545,N_46623);
nor U47691 (N_47691,N_46764,N_46643);
nor U47692 (N_47692,N_46144,N_46071);
nand U47693 (N_47693,N_46379,N_46807);
nor U47694 (N_47694,N_46726,N_46932);
nand U47695 (N_47695,N_46976,N_46743);
and U47696 (N_47696,N_46588,N_46857);
xor U47697 (N_47697,N_46733,N_46473);
nand U47698 (N_47698,N_46552,N_46888);
nand U47699 (N_47699,N_46446,N_46401);
xor U47700 (N_47700,N_46385,N_46721);
or U47701 (N_47701,N_46838,N_46639);
xnor U47702 (N_47702,N_46433,N_46808);
and U47703 (N_47703,N_46904,N_46882);
and U47704 (N_47704,N_46053,N_46378);
xor U47705 (N_47705,N_46819,N_46646);
nand U47706 (N_47706,N_46106,N_46091);
nor U47707 (N_47707,N_46534,N_46895);
and U47708 (N_47708,N_46564,N_46692);
nor U47709 (N_47709,N_46035,N_46342);
nand U47710 (N_47710,N_46432,N_46608);
nor U47711 (N_47711,N_46875,N_46136);
nand U47712 (N_47712,N_46141,N_46931);
nor U47713 (N_47713,N_46138,N_46963);
nand U47714 (N_47714,N_46431,N_46827);
nor U47715 (N_47715,N_46879,N_46637);
xnor U47716 (N_47716,N_46898,N_46331);
or U47717 (N_47717,N_46059,N_46781);
xor U47718 (N_47718,N_46382,N_46583);
nor U47719 (N_47719,N_46039,N_46281);
or U47720 (N_47720,N_46209,N_46276);
nand U47721 (N_47721,N_46576,N_46035);
xor U47722 (N_47722,N_46644,N_46040);
and U47723 (N_47723,N_46295,N_46468);
and U47724 (N_47724,N_46111,N_46135);
nor U47725 (N_47725,N_46181,N_46885);
and U47726 (N_47726,N_46646,N_46309);
and U47727 (N_47727,N_46502,N_46864);
or U47728 (N_47728,N_46883,N_46630);
or U47729 (N_47729,N_46396,N_46014);
and U47730 (N_47730,N_46610,N_46775);
or U47731 (N_47731,N_46573,N_46233);
nand U47732 (N_47732,N_46150,N_46120);
and U47733 (N_47733,N_46633,N_46849);
and U47734 (N_47734,N_46240,N_46301);
nor U47735 (N_47735,N_46383,N_46123);
xnor U47736 (N_47736,N_46099,N_46262);
nor U47737 (N_47737,N_46825,N_46614);
xnor U47738 (N_47738,N_46866,N_46301);
and U47739 (N_47739,N_46125,N_46885);
nor U47740 (N_47740,N_46356,N_46658);
nor U47741 (N_47741,N_46423,N_46247);
nor U47742 (N_47742,N_46620,N_46159);
nor U47743 (N_47743,N_46795,N_46811);
xnor U47744 (N_47744,N_46637,N_46917);
nor U47745 (N_47745,N_46695,N_46544);
or U47746 (N_47746,N_46772,N_46261);
xnor U47747 (N_47747,N_46969,N_46580);
xor U47748 (N_47748,N_46258,N_46145);
nand U47749 (N_47749,N_46255,N_46091);
or U47750 (N_47750,N_46618,N_46839);
xor U47751 (N_47751,N_46474,N_46348);
nor U47752 (N_47752,N_46380,N_46840);
nor U47753 (N_47753,N_46747,N_46495);
or U47754 (N_47754,N_46321,N_46529);
or U47755 (N_47755,N_46144,N_46668);
and U47756 (N_47756,N_46479,N_46468);
and U47757 (N_47757,N_46447,N_46162);
nor U47758 (N_47758,N_46512,N_46952);
nand U47759 (N_47759,N_46301,N_46937);
and U47760 (N_47760,N_46397,N_46449);
or U47761 (N_47761,N_46765,N_46513);
or U47762 (N_47762,N_46433,N_46414);
xnor U47763 (N_47763,N_46456,N_46471);
and U47764 (N_47764,N_46693,N_46050);
nand U47765 (N_47765,N_46617,N_46537);
and U47766 (N_47766,N_46756,N_46400);
xnor U47767 (N_47767,N_46680,N_46876);
nor U47768 (N_47768,N_46610,N_46511);
and U47769 (N_47769,N_46974,N_46399);
xnor U47770 (N_47770,N_46889,N_46619);
xnor U47771 (N_47771,N_46179,N_46411);
and U47772 (N_47772,N_46853,N_46617);
nand U47773 (N_47773,N_46765,N_46759);
or U47774 (N_47774,N_46615,N_46352);
nand U47775 (N_47775,N_46779,N_46690);
or U47776 (N_47776,N_46778,N_46941);
nor U47777 (N_47777,N_46664,N_46364);
nor U47778 (N_47778,N_46809,N_46062);
and U47779 (N_47779,N_46672,N_46279);
xnor U47780 (N_47780,N_46575,N_46184);
nor U47781 (N_47781,N_46974,N_46312);
xor U47782 (N_47782,N_46048,N_46890);
xor U47783 (N_47783,N_46162,N_46319);
nand U47784 (N_47784,N_46695,N_46777);
xor U47785 (N_47785,N_46110,N_46134);
xnor U47786 (N_47786,N_46986,N_46429);
xor U47787 (N_47787,N_46014,N_46912);
or U47788 (N_47788,N_46416,N_46121);
xnor U47789 (N_47789,N_46473,N_46137);
and U47790 (N_47790,N_46875,N_46472);
nor U47791 (N_47791,N_46466,N_46697);
or U47792 (N_47792,N_46050,N_46700);
or U47793 (N_47793,N_46737,N_46656);
xor U47794 (N_47794,N_46576,N_46750);
and U47795 (N_47795,N_46351,N_46298);
nor U47796 (N_47796,N_46188,N_46866);
nor U47797 (N_47797,N_46158,N_46513);
nand U47798 (N_47798,N_46904,N_46968);
nor U47799 (N_47799,N_46599,N_46534);
nand U47800 (N_47800,N_46182,N_46785);
nand U47801 (N_47801,N_46492,N_46226);
nor U47802 (N_47802,N_46097,N_46989);
and U47803 (N_47803,N_46015,N_46781);
xnor U47804 (N_47804,N_46029,N_46243);
and U47805 (N_47805,N_46701,N_46463);
or U47806 (N_47806,N_46341,N_46454);
nor U47807 (N_47807,N_46489,N_46121);
and U47808 (N_47808,N_46084,N_46706);
nor U47809 (N_47809,N_46471,N_46392);
nand U47810 (N_47810,N_46032,N_46838);
and U47811 (N_47811,N_46621,N_46105);
xnor U47812 (N_47812,N_46645,N_46647);
or U47813 (N_47813,N_46502,N_46323);
nand U47814 (N_47814,N_46957,N_46818);
nor U47815 (N_47815,N_46897,N_46108);
nand U47816 (N_47816,N_46487,N_46744);
nand U47817 (N_47817,N_46967,N_46345);
xor U47818 (N_47818,N_46456,N_46353);
and U47819 (N_47819,N_46712,N_46284);
and U47820 (N_47820,N_46449,N_46211);
and U47821 (N_47821,N_46580,N_46668);
or U47822 (N_47822,N_46650,N_46137);
and U47823 (N_47823,N_46014,N_46546);
and U47824 (N_47824,N_46784,N_46976);
xor U47825 (N_47825,N_46250,N_46416);
nor U47826 (N_47826,N_46935,N_46942);
or U47827 (N_47827,N_46661,N_46126);
nand U47828 (N_47828,N_46976,N_46838);
or U47829 (N_47829,N_46429,N_46557);
or U47830 (N_47830,N_46646,N_46552);
xnor U47831 (N_47831,N_46664,N_46058);
or U47832 (N_47832,N_46704,N_46448);
xnor U47833 (N_47833,N_46305,N_46855);
or U47834 (N_47834,N_46423,N_46664);
and U47835 (N_47835,N_46690,N_46871);
or U47836 (N_47836,N_46846,N_46643);
or U47837 (N_47837,N_46854,N_46416);
nand U47838 (N_47838,N_46844,N_46153);
xnor U47839 (N_47839,N_46528,N_46860);
nand U47840 (N_47840,N_46450,N_46526);
or U47841 (N_47841,N_46006,N_46281);
nor U47842 (N_47842,N_46710,N_46611);
nand U47843 (N_47843,N_46862,N_46944);
or U47844 (N_47844,N_46870,N_46536);
and U47845 (N_47845,N_46061,N_46003);
nor U47846 (N_47846,N_46052,N_46309);
nor U47847 (N_47847,N_46439,N_46259);
and U47848 (N_47848,N_46726,N_46501);
xor U47849 (N_47849,N_46563,N_46400);
nand U47850 (N_47850,N_46795,N_46456);
nor U47851 (N_47851,N_46953,N_46663);
nor U47852 (N_47852,N_46866,N_46733);
and U47853 (N_47853,N_46192,N_46484);
xor U47854 (N_47854,N_46151,N_46058);
or U47855 (N_47855,N_46421,N_46436);
and U47856 (N_47856,N_46200,N_46422);
nor U47857 (N_47857,N_46054,N_46991);
nand U47858 (N_47858,N_46499,N_46948);
or U47859 (N_47859,N_46650,N_46058);
nor U47860 (N_47860,N_46689,N_46265);
and U47861 (N_47861,N_46671,N_46030);
and U47862 (N_47862,N_46949,N_46688);
nor U47863 (N_47863,N_46922,N_46552);
nand U47864 (N_47864,N_46507,N_46834);
nand U47865 (N_47865,N_46453,N_46725);
nor U47866 (N_47866,N_46980,N_46895);
or U47867 (N_47867,N_46305,N_46603);
nand U47868 (N_47868,N_46372,N_46165);
and U47869 (N_47869,N_46021,N_46520);
nor U47870 (N_47870,N_46005,N_46416);
xnor U47871 (N_47871,N_46014,N_46986);
nor U47872 (N_47872,N_46548,N_46338);
and U47873 (N_47873,N_46787,N_46587);
xnor U47874 (N_47874,N_46744,N_46330);
xnor U47875 (N_47875,N_46969,N_46866);
and U47876 (N_47876,N_46630,N_46224);
xor U47877 (N_47877,N_46787,N_46841);
and U47878 (N_47878,N_46225,N_46910);
xnor U47879 (N_47879,N_46596,N_46352);
and U47880 (N_47880,N_46699,N_46193);
or U47881 (N_47881,N_46461,N_46360);
nand U47882 (N_47882,N_46315,N_46767);
nor U47883 (N_47883,N_46281,N_46667);
nor U47884 (N_47884,N_46618,N_46367);
nor U47885 (N_47885,N_46931,N_46282);
and U47886 (N_47886,N_46149,N_46617);
nor U47887 (N_47887,N_46932,N_46220);
nor U47888 (N_47888,N_46716,N_46821);
xor U47889 (N_47889,N_46586,N_46452);
xnor U47890 (N_47890,N_46140,N_46012);
and U47891 (N_47891,N_46369,N_46407);
nand U47892 (N_47892,N_46776,N_46279);
nor U47893 (N_47893,N_46976,N_46176);
or U47894 (N_47894,N_46716,N_46518);
xor U47895 (N_47895,N_46536,N_46652);
nand U47896 (N_47896,N_46035,N_46034);
and U47897 (N_47897,N_46477,N_46022);
and U47898 (N_47898,N_46469,N_46833);
nor U47899 (N_47899,N_46572,N_46479);
and U47900 (N_47900,N_46858,N_46638);
nand U47901 (N_47901,N_46499,N_46367);
or U47902 (N_47902,N_46668,N_46419);
nor U47903 (N_47903,N_46268,N_46662);
and U47904 (N_47904,N_46971,N_46152);
or U47905 (N_47905,N_46691,N_46850);
and U47906 (N_47906,N_46955,N_46604);
nand U47907 (N_47907,N_46620,N_46857);
nor U47908 (N_47908,N_46449,N_46141);
and U47909 (N_47909,N_46769,N_46814);
and U47910 (N_47910,N_46634,N_46369);
nand U47911 (N_47911,N_46261,N_46644);
and U47912 (N_47912,N_46375,N_46592);
nor U47913 (N_47913,N_46732,N_46839);
nand U47914 (N_47914,N_46663,N_46908);
xor U47915 (N_47915,N_46900,N_46078);
nor U47916 (N_47916,N_46369,N_46665);
nor U47917 (N_47917,N_46082,N_46971);
and U47918 (N_47918,N_46323,N_46429);
or U47919 (N_47919,N_46815,N_46754);
or U47920 (N_47920,N_46921,N_46833);
nor U47921 (N_47921,N_46531,N_46535);
nand U47922 (N_47922,N_46207,N_46839);
and U47923 (N_47923,N_46232,N_46897);
nor U47924 (N_47924,N_46351,N_46566);
nand U47925 (N_47925,N_46746,N_46843);
nor U47926 (N_47926,N_46300,N_46485);
nand U47927 (N_47927,N_46732,N_46348);
xnor U47928 (N_47928,N_46209,N_46753);
xor U47929 (N_47929,N_46038,N_46326);
nor U47930 (N_47930,N_46861,N_46905);
xor U47931 (N_47931,N_46349,N_46685);
or U47932 (N_47932,N_46577,N_46628);
nand U47933 (N_47933,N_46456,N_46180);
or U47934 (N_47934,N_46631,N_46615);
nor U47935 (N_47935,N_46539,N_46710);
or U47936 (N_47936,N_46247,N_46979);
and U47937 (N_47937,N_46233,N_46801);
or U47938 (N_47938,N_46029,N_46620);
and U47939 (N_47939,N_46306,N_46604);
or U47940 (N_47940,N_46968,N_46773);
xor U47941 (N_47941,N_46635,N_46500);
nor U47942 (N_47942,N_46249,N_46498);
or U47943 (N_47943,N_46864,N_46763);
and U47944 (N_47944,N_46899,N_46688);
or U47945 (N_47945,N_46752,N_46722);
nor U47946 (N_47946,N_46620,N_46348);
nand U47947 (N_47947,N_46045,N_46741);
and U47948 (N_47948,N_46515,N_46444);
or U47949 (N_47949,N_46552,N_46716);
or U47950 (N_47950,N_46373,N_46303);
nor U47951 (N_47951,N_46506,N_46105);
xnor U47952 (N_47952,N_46511,N_46366);
nand U47953 (N_47953,N_46455,N_46782);
nor U47954 (N_47954,N_46330,N_46650);
and U47955 (N_47955,N_46677,N_46651);
and U47956 (N_47956,N_46109,N_46439);
or U47957 (N_47957,N_46398,N_46244);
and U47958 (N_47958,N_46906,N_46457);
nand U47959 (N_47959,N_46013,N_46744);
or U47960 (N_47960,N_46500,N_46643);
nand U47961 (N_47961,N_46467,N_46801);
nor U47962 (N_47962,N_46528,N_46448);
nor U47963 (N_47963,N_46495,N_46525);
and U47964 (N_47964,N_46854,N_46721);
xor U47965 (N_47965,N_46430,N_46358);
nand U47966 (N_47966,N_46961,N_46787);
and U47967 (N_47967,N_46171,N_46368);
xor U47968 (N_47968,N_46159,N_46907);
nand U47969 (N_47969,N_46899,N_46616);
nor U47970 (N_47970,N_46207,N_46765);
nand U47971 (N_47971,N_46049,N_46879);
nand U47972 (N_47972,N_46678,N_46245);
xor U47973 (N_47973,N_46137,N_46726);
or U47974 (N_47974,N_46599,N_46009);
nand U47975 (N_47975,N_46646,N_46841);
and U47976 (N_47976,N_46955,N_46614);
nand U47977 (N_47977,N_46847,N_46406);
nand U47978 (N_47978,N_46211,N_46246);
and U47979 (N_47979,N_46019,N_46095);
xor U47980 (N_47980,N_46691,N_46101);
nand U47981 (N_47981,N_46744,N_46789);
xor U47982 (N_47982,N_46575,N_46113);
or U47983 (N_47983,N_46237,N_46920);
nor U47984 (N_47984,N_46132,N_46171);
or U47985 (N_47985,N_46840,N_46523);
xor U47986 (N_47986,N_46370,N_46890);
nand U47987 (N_47987,N_46465,N_46894);
xnor U47988 (N_47988,N_46963,N_46913);
nor U47989 (N_47989,N_46885,N_46829);
xnor U47990 (N_47990,N_46719,N_46957);
or U47991 (N_47991,N_46240,N_46453);
and U47992 (N_47992,N_46224,N_46672);
nand U47993 (N_47993,N_46303,N_46840);
xnor U47994 (N_47994,N_46239,N_46803);
or U47995 (N_47995,N_46673,N_46890);
xnor U47996 (N_47996,N_46987,N_46908);
or U47997 (N_47997,N_46914,N_46272);
and U47998 (N_47998,N_46965,N_46651);
or U47999 (N_47999,N_46587,N_46000);
or U48000 (N_48000,N_47842,N_47705);
or U48001 (N_48001,N_47216,N_47794);
and U48002 (N_48002,N_47424,N_47582);
xnor U48003 (N_48003,N_47097,N_47007);
or U48004 (N_48004,N_47947,N_47348);
nand U48005 (N_48005,N_47665,N_47089);
or U48006 (N_48006,N_47963,N_47503);
and U48007 (N_48007,N_47179,N_47881);
or U48008 (N_48008,N_47144,N_47683);
or U48009 (N_48009,N_47676,N_47324);
xnor U48010 (N_48010,N_47129,N_47235);
nor U48011 (N_48011,N_47560,N_47205);
nand U48012 (N_48012,N_47112,N_47780);
and U48013 (N_48013,N_47158,N_47702);
nand U48014 (N_48014,N_47069,N_47633);
or U48015 (N_48015,N_47987,N_47398);
or U48016 (N_48016,N_47020,N_47209);
xor U48017 (N_48017,N_47653,N_47903);
and U48018 (N_48018,N_47717,N_47625);
nand U48019 (N_48019,N_47631,N_47293);
xnor U48020 (N_48020,N_47461,N_47298);
nand U48021 (N_48021,N_47978,N_47237);
and U48022 (N_48022,N_47678,N_47056);
xnor U48023 (N_48023,N_47621,N_47051);
and U48024 (N_48024,N_47491,N_47327);
xor U48025 (N_48025,N_47090,N_47677);
nor U48026 (N_48026,N_47851,N_47386);
or U48027 (N_48027,N_47896,N_47308);
or U48028 (N_48028,N_47151,N_47382);
and U48029 (N_48029,N_47040,N_47006);
nand U48030 (N_48030,N_47068,N_47243);
or U48031 (N_48031,N_47379,N_47866);
xor U48032 (N_48032,N_47303,N_47604);
nand U48033 (N_48033,N_47688,N_47085);
or U48034 (N_48034,N_47497,N_47536);
xnor U48035 (N_48035,N_47302,N_47787);
nand U48036 (N_48036,N_47409,N_47356);
nand U48037 (N_48037,N_47605,N_47574);
nor U48038 (N_48038,N_47728,N_47516);
and U48039 (N_48039,N_47519,N_47742);
nand U48040 (N_48040,N_47091,N_47354);
xnor U48041 (N_48041,N_47583,N_47325);
nor U48042 (N_48042,N_47626,N_47443);
or U48043 (N_48043,N_47732,N_47811);
and U48044 (N_48044,N_47912,N_47101);
and U48045 (N_48045,N_47171,N_47393);
or U48046 (N_48046,N_47817,N_47161);
xor U48047 (N_48047,N_47652,N_47092);
or U48048 (N_48048,N_47707,N_47288);
or U48049 (N_48049,N_47149,N_47062);
nor U48050 (N_48050,N_47370,N_47390);
or U48051 (N_48051,N_47154,N_47425);
xor U48052 (N_48052,N_47444,N_47814);
and U48053 (N_48053,N_47744,N_47966);
nor U48054 (N_48054,N_47697,N_47788);
or U48055 (N_48055,N_47537,N_47615);
or U48056 (N_48056,N_47271,N_47834);
nor U48057 (N_48057,N_47180,N_47982);
or U48058 (N_48058,N_47862,N_47534);
nand U48059 (N_48059,N_47291,N_47859);
or U48060 (N_48060,N_47614,N_47523);
or U48061 (N_48061,N_47945,N_47545);
xor U48062 (N_48062,N_47646,N_47266);
xnor U48063 (N_48063,N_47353,N_47185);
or U48064 (N_48064,N_47385,N_47973);
xnor U48065 (N_48065,N_47400,N_47964);
xnor U48066 (N_48066,N_47925,N_47558);
and U48067 (N_48067,N_47512,N_47808);
and U48068 (N_48068,N_47643,N_47577);
and U48069 (N_48069,N_47720,N_47207);
xor U48070 (N_48070,N_47992,N_47478);
and U48071 (N_48071,N_47823,N_47182);
nand U48072 (N_48072,N_47969,N_47220);
nand U48073 (N_48073,N_47907,N_47367);
nor U48074 (N_48074,N_47566,N_47835);
xor U48075 (N_48075,N_47190,N_47289);
nor U48076 (N_48076,N_47886,N_47706);
or U48077 (N_48077,N_47977,N_47957);
nor U48078 (N_48078,N_47195,N_47900);
nor U48079 (N_48079,N_47052,N_47251);
nor U48080 (N_48080,N_47622,N_47448);
or U48081 (N_48081,N_47918,N_47338);
xnor U48082 (N_48082,N_47781,N_47562);
nor U48083 (N_48083,N_47402,N_47230);
nand U48084 (N_48084,N_47596,N_47273);
nand U48085 (N_48085,N_47058,N_47684);
and U48086 (N_48086,N_47698,N_47740);
nand U48087 (N_48087,N_47313,N_47831);
nand U48088 (N_48088,N_47261,N_47021);
nand U48089 (N_48089,N_47247,N_47726);
and U48090 (N_48090,N_47135,N_47752);
and U48091 (N_48091,N_47113,N_47471);
nand U48092 (N_48092,N_47428,N_47989);
or U48093 (N_48093,N_47829,N_47024);
nand U48094 (N_48094,N_47259,N_47334);
or U48095 (N_48095,N_47733,N_47368);
or U48096 (N_48096,N_47713,N_47380);
nor U48097 (N_48097,N_47347,N_47768);
nand U48098 (N_48098,N_47679,N_47087);
nor U48099 (N_48099,N_47399,N_47609);
nor U48100 (N_48100,N_47258,N_47522);
nand U48101 (N_48101,N_47505,N_47724);
xor U48102 (N_48102,N_47839,N_47295);
or U48103 (N_48103,N_47847,N_47240);
xnor U48104 (N_48104,N_47983,N_47563);
nor U48105 (N_48105,N_47818,N_47875);
nand U48106 (N_48106,N_47958,N_47580);
and U48107 (N_48107,N_47594,N_47476);
nand U48108 (N_48108,N_47120,N_47730);
nand U48109 (N_48109,N_47454,N_47821);
xor U48110 (N_48110,N_47198,N_47208);
xnor U48111 (N_48111,N_47692,N_47392);
nand U48112 (N_48112,N_47283,N_47714);
or U48113 (N_48113,N_47268,N_47634);
xnor U48114 (N_48114,N_47433,N_47890);
or U48115 (N_48115,N_47070,N_47877);
or U48116 (N_48116,N_47736,N_47670);
xnor U48117 (N_48117,N_47304,N_47828);
nand U48118 (N_48118,N_47943,N_47009);
or U48119 (N_48119,N_47806,N_47319);
and U48120 (N_48120,N_47483,N_47311);
xor U48121 (N_48121,N_47538,N_47836);
nand U48122 (N_48122,N_47718,N_47294);
nand U48123 (N_48123,N_47529,N_47355);
nor U48124 (N_48124,N_47329,N_47406);
or U48125 (N_48125,N_47146,N_47553);
xor U48126 (N_48126,N_47559,N_47739);
nand U48127 (N_48127,N_47822,N_47830);
nand U48128 (N_48128,N_47194,N_47929);
xnor U48129 (N_48129,N_47300,N_47447);
nand U48130 (N_48130,N_47126,N_47920);
nor U48131 (N_48131,N_47429,N_47515);
nor U48132 (N_48132,N_47915,N_47793);
nor U48133 (N_48133,N_47939,N_47466);
and U48134 (N_48134,N_47513,N_47954);
nand U48135 (N_48135,N_47778,N_47979);
nor U48136 (N_48136,N_47949,N_47723);
or U48137 (N_48137,N_47280,N_47910);
xor U48138 (N_48138,N_47388,N_47123);
or U48139 (N_48139,N_47776,N_47879);
and U48140 (N_48140,N_47629,N_47164);
nor U48141 (N_48141,N_47500,N_47548);
nand U48142 (N_48142,N_47172,N_47043);
xnor U48143 (N_48143,N_47581,N_47326);
nor U48144 (N_48144,N_47250,N_47639);
or U48145 (N_48145,N_47944,N_47997);
or U48146 (N_48146,N_47961,N_47800);
xnor U48147 (N_48147,N_47239,N_47016);
or U48148 (N_48148,N_47140,N_47215);
nor U48149 (N_48149,N_47673,N_47391);
nor U48150 (N_48150,N_47991,N_47077);
xor U48151 (N_48151,N_47033,N_47850);
xnor U48152 (N_48152,N_47034,N_47318);
or U48153 (N_48153,N_47103,N_47663);
and U48154 (N_48154,N_47246,N_47312);
or U48155 (N_48155,N_47932,N_47597);
xor U48156 (N_48156,N_47467,N_47064);
nand U48157 (N_48157,N_47893,N_47975);
or U48158 (N_48158,N_47131,N_47843);
nand U48159 (N_48159,N_47018,N_47061);
xnor U48160 (N_48160,N_47395,N_47366);
or U48161 (N_48161,N_47286,N_47008);
or U48162 (N_48162,N_47420,N_47544);
and U48163 (N_48163,N_47186,N_47122);
nor U48164 (N_48164,N_47813,N_47328);
nand U48165 (N_48165,N_47438,N_47946);
nor U48166 (N_48166,N_47712,N_47244);
nand U48167 (N_48167,N_47446,N_47242);
nor U48168 (N_48168,N_47786,N_47801);
nand U48169 (N_48169,N_47825,N_47098);
or U48170 (N_48170,N_47317,N_47521);
nor U48171 (N_48171,N_47542,N_47254);
xor U48172 (N_48172,N_47919,N_47602);
nand U48173 (N_48173,N_47297,N_47490);
nand U48174 (N_48174,N_47134,N_47369);
nand U48175 (N_48175,N_47022,N_47114);
nor U48176 (N_48176,N_47985,N_47265);
nor U48177 (N_48177,N_47407,N_47066);
nor U48178 (N_48178,N_47193,N_47440);
nor U48179 (N_48179,N_47591,N_47050);
and U48180 (N_48180,N_47690,N_47869);
and U48181 (N_48181,N_47059,N_47054);
or U48182 (N_48182,N_47887,N_47322);
xnor U48183 (N_48183,N_47725,N_47014);
nor U48184 (N_48184,N_47231,N_47485);
xor U48185 (N_48185,N_47867,N_47856);
xor U48186 (N_48186,N_47660,N_47037);
nand U48187 (N_48187,N_47346,N_47555);
xor U48188 (N_48188,N_47854,N_47272);
nand U48189 (N_48189,N_47727,N_47403);
nand U48190 (N_48190,N_47990,N_47635);
and U48191 (N_48191,N_47188,N_47894);
or U48192 (N_48192,N_47870,N_47387);
and U48193 (N_48193,N_47816,N_47671);
xnor U48194 (N_48194,N_47422,N_47249);
or U48195 (N_48195,N_47238,N_47518);
and U48196 (N_48196,N_47674,N_47948);
nor U48197 (N_48197,N_47189,N_47248);
nand U48198 (N_48198,N_47108,N_47832);
xnor U48199 (N_48199,N_47695,N_47371);
xnor U48200 (N_48200,N_47155,N_47873);
xor U48201 (N_48201,N_47549,N_47613);
xor U48202 (N_48202,N_47750,N_47359);
nand U48203 (N_48203,N_47032,N_47861);
and U48204 (N_48204,N_47133,N_47649);
xor U48205 (N_48205,N_47612,N_47796);
xnor U48206 (N_48206,N_47000,N_47415);
nor U48207 (N_48207,N_47252,N_47459);
nand U48208 (N_48208,N_47405,N_47372);
nand U48209 (N_48209,N_47775,N_47524);
xnor U48210 (N_48210,N_47262,N_47655);
xnor U48211 (N_48211,N_47735,N_47445);
nand U48212 (N_48212,N_47658,N_47936);
nor U48213 (N_48213,N_47082,N_47715);
or U48214 (N_48214,N_47804,N_47528);
nand U48215 (N_48215,N_47756,N_47603);
or U48216 (N_48216,N_47901,N_47965);
nor U48217 (N_48217,N_47586,N_47229);
and U48218 (N_48218,N_47908,N_47116);
xor U48219 (N_48219,N_47437,N_47026);
and U48220 (N_48220,N_47336,N_47691);
xnor U48221 (N_48221,N_47351,N_47373);
and U48222 (N_48222,N_47426,N_47860);
xnor U48223 (N_48223,N_47567,N_47340);
or U48224 (N_48224,N_47645,N_47748);
or U48225 (N_48225,N_47427,N_47410);
xor U48226 (N_48226,N_47759,N_47441);
and U48227 (N_48227,N_47417,N_47951);
nand U48228 (N_48228,N_47130,N_47075);
nand U48229 (N_48229,N_47094,N_47938);
or U48230 (N_48230,N_47928,N_47457);
or U48231 (N_48231,N_47472,N_47275);
nor U48232 (N_48232,N_47914,N_47320);
and U48233 (N_48233,N_47330,N_47974);
or U48234 (N_48234,N_47510,N_47587);
xor U48235 (N_48235,N_47227,N_47079);
nand U48236 (N_48236,N_47960,N_47197);
or U48237 (N_48237,N_47853,N_47119);
xor U48238 (N_48238,N_47620,N_47905);
xnor U48239 (N_48239,N_47526,N_47934);
nor U48240 (N_48240,N_47669,N_47554);
nand U48241 (N_48241,N_47274,N_47520);
nand U48242 (N_48242,N_47078,N_47153);
or U48243 (N_48243,N_47001,N_47412);
or U48244 (N_48244,N_47159,N_47530);
or U48245 (N_48245,N_47093,N_47588);
or U48246 (N_48246,N_47540,N_47342);
nand U48247 (N_48247,N_47502,N_47199);
and U48248 (N_48248,N_47086,N_47865);
xor U48249 (N_48249,N_47637,N_47999);
nor U48250 (N_48250,N_47228,N_47281);
nand U48251 (N_48251,N_47686,N_47290);
or U48252 (N_48252,N_47572,N_47600);
or U48253 (N_48253,N_47644,N_47143);
and U48254 (N_48254,N_47111,N_47494);
xnor U48255 (N_48255,N_47798,N_47270);
nand U48256 (N_48256,N_47616,N_47088);
nand U48257 (N_48257,N_47942,N_47439);
xor U48258 (N_48258,N_47771,N_47004);
and U48259 (N_48259,N_47165,N_47333);
nor U48260 (N_48260,N_47384,N_47307);
or U48261 (N_48261,N_47305,N_47871);
or U48262 (N_48262,N_47511,N_47508);
nor U48263 (N_48263,N_47408,N_47592);
nand U48264 (N_48264,N_47028,N_47880);
nand U48265 (N_48265,N_47765,N_47442);
nor U48266 (N_48266,N_47475,N_47221);
xor U48267 (N_48267,N_47651,N_47118);
and U48268 (N_48268,N_47301,N_47699);
nor U48269 (N_48269,N_47223,N_47046);
or U48270 (N_48270,N_47096,N_47783);
nor U48271 (N_48271,N_47824,N_47498);
or U48272 (N_48272,N_47891,N_47343);
nor U48273 (N_48273,N_47256,N_47257);
and U48274 (N_48274,N_47121,N_47998);
and U48275 (N_48275,N_47469,N_47414);
nor U48276 (N_48276,N_47202,N_47166);
nor U48277 (N_48277,N_47263,N_47858);
xnor U48278 (N_48278,N_47138,N_47152);
nand U48279 (N_48279,N_47374,N_47909);
xor U48280 (N_48280,N_47922,N_47535);
nor U48281 (N_48281,N_47729,N_47045);
nor U48282 (N_48282,N_47504,N_47496);
nand U48283 (N_48283,N_47168,N_47940);
nand U48284 (N_48284,N_47364,N_47589);
nor U48285 (N_48285,N_47036,N_47852);
nand U48286 (N_48286,N_47255,N_47971);
or U48287 (N_48287,N_47309,N_47685);
and U48288 (N_48288,N_47815,N_47777);
and U48289 (N_48289,N_47795,N_47279);
nand U48290 (N_48290,N_47003,N_47187);
nand U48291 (N_48291,N_47352,N_47627);
or U48292 (N_48292,N_47984,N_47421);
nor U48293 (N_48293,N_47394,N_47277);
nand U48294 (N_48294,N_47264,N_47745);
nor U48295 (N_48295,N_47953,N_47917);
or U48296 (N_48296,N_47218,N_47565);
and U48297 (N_48297,N_47100,N_47864);
and U48298 (N_48298,N_47701,N_47737);
xnor U48299 (N_48299,N_47299,N_47682);
nor U48300 (N_48300,N_47623,N_47487);
nand U48301 (N_48301,N_47023,N_47749);
nor U48302 (N_48302,N_47225,N_47477);
nand U48303 (N_48303,N_47716,N_47206);
or U48304 (N_48304,N_47995,N_47930);
nor U48305 (N_48305,N_47610,N_47640);
or U48306 (N_48306,N_47315,N_47527);
xnor U48307 (N_48307,N_47601,N_47770);
or U48308 (N_48308,N_47878,N_47234);
nand U48309 (N_48309,N_47630,N_47576);
and U48310 (N_48310,N_47618,N_47063);
xnor U48311 (N_48311,N_47377,N_47766);
xnor U48312 (N_48312,N_47889,N_47196);
nor U48313 (N_48313,N_47042,N_47672);
xor U48314 (N_48314,N_47556,N_47647);
nor U48315 (N_48315,N_47784,N_47902);
and U48316 (N_48316,N_47950,N_47285);
xor U48317 (N_48317,N_47191,N_47650);
nand U48318 (N_48318,N_47782,N_47048);
nor U48319 (N_48319,N_47065,N_47452);
and U48320 (N_48320,N_47245,N_47762);
or U48321 (N_48321,N_47696,N_47287);
nor U48322 (N_48322,N_47167,N_47711);
nand U48323 (N_48323,N_47057,N_47430);
nor U48324 (N_48324,N_47492,N_47840);
xor U48325 (N_48325,N_47080,N_47809);
nand U48326 (N_48326,N_47774,N_47599);
nor U48327 (N_48327,N_47418,N_47731);
and U48328 (N_48328,N_47358,N_47769);
nor U48329 (N_48329,N_47470,N_47213);
nand U48330 (N_48330,N_47175,N_47976);
and U48331 (N_48331,N_47656,N_47224);
xor U48332 (N_48332,N_47413,N_47332);
and U48333 (N_48333,N_47968,N_47150);
nor U48334 (N_48334,N_47177,N_47173);
nor U48335 (N_48335,N_47148,N_47017);
xor U48336 (N_48336,N_47642,N_47719);
and U48337 (N_48337,N_47758,N_47137);
or U48338 (N_48338,N_47125,N_47361);
or U48339 (N_48339,N_47106,N_47986);
and U48340 (N_48340,N_47827,N_47031);
or U48341 (N_48341,N_47904,N_47884);
and U48342 (N_48342,N_47060,N_47451);
or U48343 (N_48343,N_47109,N_47010);
and U48344 (N_48344,N_47204,N_47906);
nor U48345 (N_48345,N_47797,N_47139);
and U48346 (N_48346,N_47431,N_47509);
nor U48347 (N_48347,N_47575,N_47792);
nor U48348 (N_48348,N_47105,N_47005);
or U48349 (N_48349,N_47753,N_47269);
or U48350 (N_48350,N_47345,N_47619);
or U48351 (N_48351,N_47462,N_47331);
xnor U48352 (N_48352,N_47668,N_47363);
and U48353 (N_48353,N_47002,N_47099);
and U48354 (N_48354,N_47826,N_47585);
and U48355 (N_48355,N_47981,N_47927);
or U48356 (N_48356,N_47226,N_47767);
nor U48357 (N_48357,N_47694,N_47241);
and U48358 (N_48358,N_47550,N_47617);
or U48359 (N_48359,N_47030,N_47807);
and U48360 (N_48360,N_47799,N_47874);
or U48361 (N_48361,N_47067,N_47110);
nor U48362 (N_48362,N_47757,N_47200);
nor U48363 (N_48363,N_47675,N_47474);
and U48364 (N_48364,N_47136,N_47785);
nand U48365 (N_48365,N_47899,N_47924);
xnor U48366 (N_48366,N_47460,N_47708);
or U48367 (N_48367,N_47011,N_47480);
or U48368 (N_48368,N_47606,N_47608);
and U48369 (N_48369,N_47595,N_47872);
or U48370 (N_48370,N_47038,N_47156);
xor U48371 (N_48371,N_47803,N_47641);
nor U48372 (N_48372,N_47763,N_47959);
nor U48373 (N_48373,N_47183,N_47624);
nand U48374 (N_48374,N_47681,N_47547);
xnor U48375 (N_48375,N_47479,N_47423);
or U48376 (N_48376,N_47169,N_47081);
or U48377 (N_48377,N_47552,N_47754);
or U48378 (N_48378,N_47115,N_47276);
nand U48379 (N_48379,N_47214,N_47913);
xor U48380 (N_48380,N_47898,N_47638);
nand U48381 (N_48381,N_47482,N_47689);
xor U48382 (N_48382,N_47855,N_47436);
nor U48383 (N_48383,N_47306,N_47632);
and U48384 (N_48384,N_47260,N_47564);
or U48385 (N_48385,N_47012,N_47734);
nand U48386 (N_48386,N_47570,N_47489);
nand U48387 (N_48387,N_47779,N_47233);
nand U48388 (N_48388,N_47885,N_47453);
nor U48389 (N_48389,N_47411,N_47344);
xor U48390 (N_48390,N_47703,N_47027);
nor U48391 (N_48391,N_47802,N_47868);
nand U48392 (N_48392,N_47212,N_47141);
nor U48393 (N_48393,N_47972,N_47365);
nand U48394 (N_48394,N_47755,N_47278);
xor U48395 (N_48395,N_47071,N_47076);
or U48396 (N_48396,N_47941,N_47435);
nor U48397 (N_48397,N_47389,N_47967);
and U48398 (N_48398,N_47506,N_47841);
and U48399 (N_48399,N_47284,N_47956);
nand U48400 (N_48400,N_47693,N_47219);
nand U48401 (N_48401,N_47211,N_47911);
nand U48402 (N_48402,N_47019,N_47882);
nor U48403 (N_48403,N_47107,N_47751);
nor U48404 (N_48404,N_47292,N_47937);
nor U48405 (N_48405,N_47531,N_47310);
and U48406 (N_48406,N_47486,N_47499);
xnor U48407 (N_48407,N_47222,N_47493);
xor U48408 (N_48408,N_47047,N_47095);
and U48409 (N_48409,N_47721,N_47514);
or U48410 (N_48410,N_47145,N_47162);
and U48411 (N_48411,N_47988,N_47517);
or U48412 (N_48412,N_47473,N_47142);
nand U48413 (N_48413,N_47041,N_47848);
nor U48414 (N_48414,N_47654,N_47184);
or U48415 (N_48415,N_47383,N_47636);
and U48416 (N_48416,N_47738,N_47084);
nor U48417 (N_48417,N_47741,N_47743);
nand U48418 (N_48418,N_47760,N_47434);
and U48419 (N_48419,N_47666,N_47539);
nand U48420 (N_48420,N_47895,N_47584);
nor U48421 (N_48421,N_47128,N_47579);
nand U48422 (N_48422,N_47104,N_47931);
nor U48423 (N_48423,N_47844,N_47747);
or U48424 (N_48424,N_47661,N_47812);
or U48425 (N_48425,N_47532,N_47049);
nor U48426 (N_48426,N_47072,N_47568);
nor U48427 (N_48427,N_47419,N_47837);
xor U48428 (N_48428,N_47456,N_47362);
and U48429 (N_48429,N_47933,N_47700);
nand U48430 (N_48430,N_47236,N_47449);
nor U48431 (N_48431,N_47996,N_47029);
nor U48432 (N_48432,N_47955,N_47192);
or U48433 (N_48433,N_47764,N_47892);
and U48434 (N_48434,N_47464,N_47450);
or U48435 (N_48435,N_47217,N_47883);
and U48436 (N_48436,N_47124,N_47117);
or U48437 (N_48437,N_47375,N_47296);
nor U48438 (N_48438,N_47176,N_47484);
xor U48439 (N_48439,N_47102,N_47127);
nor U48440 (N_48440,N_47455,N_47888);
nand U48441 (N_48441,N_47339,N_47035);
or U48442 (N_48442,N_47833,N_47013);
and U48443 (N_48443,N_47335,N_47857);
and U48444 (N_48444,N_47160,N_47863);
nand U48445 (N_48445,N_47657,N_47337);
or U48446 (N_48446,N_47845,N_47667);
nand U48447 (N_48447,N_47357,N_47463);
and U48448 (N_48448,N_47132,N_47598);
xor U48449 (N_48449,N_47432,N_47397);
xor U48450 (N_48450,N_47316,N_47571);
nor U48451 (N_48451,N_47789,N_47210);
or U48452 (N_48452,N_47525,N_47541);
nor U48453 (N_48453,N_47607,N_47282);
nand U48454 (N_48454,N_47015,N_47593);
xnor U48455 (N_48455,N_47926,N_47628);
or U48456 (N_48456,N_47849,N_47350);
xor U48457 (N_48457,N_47025,N_47897);
xor U48458 (N_48458,N_47994,N_47314);
or U48459 (N_48459,N_47819,N_47321);
nand U48460 (N_48460,N_47232,N_47488);
nor U48461 (N_48461,N_47147,N_47381);
or U48462 (N_48462,N_47501,N_47341);
or U48463 (N_48463,N_47952,N_47044);
nand U48464 (N_48464,N_47662,N_47935);
and U48465 (N_48465,N_47546,N_47970);
and U48466 (N_48466,N_47323,N_47923);
or U48467 (N_48467,N_47772,N_47962);
nand U48468 (N_48468,N_47773,N_47201);
nor U48469 (N_48469,N_47495,N_47846);
or U48470 (N_48470,N_47074,N_47710);
and U48471 (N_48471,N_47790,N_47349);
xor U48472 (N_48472,N_47396,N_47178);
nand U48473 (N_48473,N_47543,N_47791);
xor U48474 (N_48474,N_47611,N_47468);
nor U48475 (N_48475,N_47704,N_47163);
or U48476 (N_48476,N_47253,N_47203);
xnor U48477 (N_48477,N_47980,N_47507);
xnor U48478 (N_48478,N_47838,N_47073);
nor U48479 (N_48479,N_47481,N_47170);
nor U48480 (N_48480,N_47820,N_47181);
or U48481 (N_48481,N_47267,N_47404);
xnor U48482 (N_48482,N_47039,N_47687);
nor U48483 (N_48483,N_47916,N_47416);
or U48484 (N_48484,N_47680,N_47557);
or U48485 (N_48485,N_47805,N_47578);
nand U48486 (N_48486,N_47569,N_47083);
xor U48487 (N_48487,N_47810,N_47590);
and U48488 (N_48488,N_47533,N_47053);
nand U48489 (N_48489,N_47465,N_47458);
xor U48490 (N_48490,N_47876,N_47551);
and U48491 (N_48491,N_47561,N_47746);
nand U48492 (N_48492,N_47648,N_47055);
nand U48493 (N_48493,N_47664,N_47722);
or U48494 (N_48494,N_47157,N_47993);
and U48495 (N_48495,N_47709,N_47659);
xor U48496 (N_48496,N_47360,N_47378);
or U48497 (N_48497,N_47573,N_47761);
nand U48498 (N_48498,N_47921,N_47174);
and U48499 (N_48499,N_47376,N_47401);
and U48500 (N_48500,N_47760,N_47269);
nand U48501 (N_48501,N_47160,N_47001);
and U48502 (N_48502,N_47078,N_47436);
nand U48503 (N_48503,N_47925,N_47196);
nand U48504 (N_48504,N_47593,N_47544);
and U48505 (N_48505,N_47631,N_47489);
nand U48506 (N_48506,N_47684,N_47442);
or U48507 (N_48507,N_47413,N_47036);
nor U48508 (N_48508,N_47149,N_47386);
nor U48509 (N_48509,N_47750,N_47368);
or U48510 (N_48510,N_47563,N_47747);
xor U48511 (N_48511,N_47683,N_47955);
xor U48512 (N_48512,N_47213,N_47913);
and U48513 (N_48513,N_47175,N_47034);
and U48514 (N_48514,N_47727,N_47320);
or U48515 (N_48515,N_47169,N_47025);
nand U48516 (N_48516,N_47031,N_47484);
or U48517 (N_48517,N_47094,N_47761);
and U48518 (N_48518,N_47929,N_47387);
xnor U48519 (N_48519,N_47572,N_47901);
or U48520 (N_48520,N_47222,N_47238);
and U48521 (N_48521,N_47626,N_47460);
or U48522 (N_48522,N_47689,N_47352);
xnor U48523 (N_48523,N_47573,N_47450);
nand U48524 (N_48524,N_47902,N_47899);
nand U48525 (N_48525,N_47632,N_47040);
and U48526 (N_48526,N_47125,N_47516);
nor U48527 (N_48527,N_47030,N_47133);
nand U48528 (N_48528,N_47501,N_47705);
xnor U48529 (N_48529,N_47648,N_47782);
and U48530 (N_48530,N_47488,N_47409);
and U48531 (N_48531,N_47521,N_47519);
xnor U48532 (N_48532,N_47536,N_47271);
nand U48533 (N_48533,N_47805,N_47312);
and U48534 (N_48534,N_47744,N_47030);
or U48535 (N_48535,N_47246,N_47123);
or U48536 (N_48536,N_47650,N_47051);
or U48537 (N_48537,N_47955,N_47229);
or U48538 (N_48538,N_47003,N_47803);
or U48539 (N_48539,N_47214,N_47508);
or U48540 (N_48540,N_47558,N_47515);
or U48541 (N_48541,N_47459,N_47631);
or U48542 (N_48542,N_47489,N_47196);
and U48543 (N_48543,N_47587,N_47842);
xor U48544 (N_48544,N_47474,N_47143);
and U48545 (N_48545,N_47693,N_47809);
or U48546 (N_48546,N_47155,N_47498);
nor U48547 (N_48547,N_47114,N_47479);
nand U48548 (N_48548,N_47083,N_47961);
nor U48549 (N_48549,N_47244,N_47574);
or U48550 (N_48550,N_47860,N_47340);
and U48551 (N_48551,N_47748,N_47931);
nand U48552 (N_48552,N_47379,N_47234);
or U48553 (N_48553,N_47089,N_47904);
nor U48554 (N_48554,N_47961,N_47586);
nand U48555 (N_48555,N_47316,N_47416);
and U48556 (N_48556,N_47511,N_47954);
xnor U48557 (N_48557,N_47436,N_47527);
nor U48558 (N_48558,N_47603,N_47936);
xor U48559 (N_48559,N_47557,N_47207);
or U48560 (N_48560,N_47853,N_47794);
nor U48561 (N_48561,N_47419,N_47530);
and U48562 (N_48562,N_47442,N_47316);
xor U48563 (N_48563,N_47971,N_47705);
xor U48564 (N_48564,N_47686,N_47915);
xor U48565 (N_48565,N_47155,N_47759);
nand U48566 (N_48566,N_47836,N_47888);
nor U48567 (N_48567,N_47676,N_47972);
xor U48568 (N_48568,N_47262,N_47470);
nor U48569 (N_48569,N_47005,N_47659);
nor U48570 (N_48570,N_47656,N_47752);
nor U48571 (N_48571,N_47329,N_47019);
or U48572 (N_48572,N_47845,N_47823);
xor U48573 (N_48573,N_47650,N_47953);
and U48574 (N_48574,N_47315,N_47144);
nand U48575 (N_48575,N_47545,N_47135);
or U48576 (N_48576,N_47952,N_47219);
nor U48577 (N_48577,N_47507,N_47679);
and U48578 (N_48578,N_47994,N_47172);
xnor U48579 (N_48579,N_47832,N_47340);
and U48580 (N_48580,N_47398,N_47885);
and U48581 (N_48581,N_47499,N_47359);
xor U48582 (N_48582,N_47860,N_47867);
and U48583 (N_48583,N_47424,N_47181);
or U48584 (N_48584,N_47722,N_47571);
or U48585 (N_48585,N_47086,N_47184);
nand U48586 (N_48586,N_47666,N_47161);
nor U48587 (N_48587,N_47290,N_47354);
and U48588 (N_48588,N_47262,N_47198);
xor U48589 (N_48589,N_47397,N_47198);
and U48590 (N_48590,N_47633,N_47653);
and U48591 (N_48591,N_47632,N_47789);
nor U48592 (N_48592,N_47692,N_47675);
nand U48593 (N_48593,N_47733,N_47152);
or U48594 (N_48594,N_47872,N_47541);
and U48595 (N_48595,N_47098,N_47338);
or U48596 (N_48596,N_47234,N_47442);
xor U48597 (N_48597,N_47344,N_47038);
or U48598 (N_48598,N_47959,N_47955);
or U48599 (N_48599,N_47208,N_47076);
or U48600 (N_48600,N_47461,N_47825);
nor U48601 (N_48601,N_47011,N_47797);
or U48602 (N_48602,N_47314,N_47861);
and U48603 (N_48603,N_47037,N_47477);
or U48604 (N_48604,N_47313,N_47877);
nand U48605 (N_48605,N_47881,N_47819);
nor U48606 (N_48606,N_47584,N_47581);
nor U48607 (N_48607,N_47669,N_47130);
xnor U48608 (N_48608,N_47664,N_47833);
xor U48609 (N_48609,N_47440,N_47890);
xor U48610 (N_48610,N_47162,N_47251);
nand U48611 (N_48611,N_47563,N_47285);
nand U48612 (N_48612,N_47063,N_47861);
and U48613 (N_48613,N_47643,N_47776);
xnor U48614 (N_48614,N_47363,N_47512);
and U48615 (N_48615,N_47492,N_47580);
xor U48616 (N_48616,N_47503,N_47190);
or U48617 (N_48617,N_47656,N_47136);
nand U48618 (N_48618,N_47206,N_47065);
xor U48619 (N_48619,N_47076,N_47750);
nor U48620 (N_48620,N_47158,N_47731);
or U48621 (N_48621,N_47481,N_47047);
and U48622 (N_48622,N_47252,N_47384);
xor U48623 (N_48623,N_47196,N_47251);
nor U48624 (N_48624,N_47423,N_47077);
or U48625 (N_48625,N_47820,N_47445);
and U48626 (N_48626,N_47599,N_47791);
nand U48627 (N_48627,N_47319,N_47830);
and U48628 (N_48628,N_47087,N_47202);
nand U48629 (N_48629,N_47623,N_47709);
nor U48630 (N_48630,N_47522,N_47824);
xor U48631 (N_48631,N_47665,N_47601);
nand U48632 (N_48632,N_47502,N_47421);
nand U48633 (N_48633,N_47596,N_47875);
xor U48634 (N_48634,N_47915,N_47554);
xnor U48635 (N_48635,N_47153,N_47480);
nor U48636 (N_48636,N_47069,N_47817);
xnor U48637 (N_48637,N_47494,N_47184);
nand U48638 (N_48638,N_47600,N_47382);
xnor U48639 (N_48639,N_47756,N_47780);
xnor U48640 (N_48640,N_47957,N_47803);
nor U48641 (N_48641,N_47012,N_47003);
nand U48642 (N_48642,N_47242,N_47159);
and U48643 (N_48643,N_47380,N_47637);
or U48644 (N_48644,N_47227,N_47818);
nor U48645 (N_48645,N_47931,N_47740);
xnor U48646 (N_48646,N_47210,N_47256);
or U48647 (N_48647,N_47517,N_47584);
nand U48648 (N_48648,N_47994,N_47084);
nor U48649 (N_48649,N_47953,N_47286);
nor U48650 (N_48650,N_47444,N_47470);
or U48651 (N_48651,N_47732,N_47685);
xnor U48652 (N_48652,N_47400,N_47921);
nor U48653 (N_48653,N_47095,N_47996);
or U48654 (N_48654,N_47038,N_47253);
or U48655 (N_48655,N_47301,N_47425);
nand U48656 (N_48656,N_47403,N_47847);
and U48657 (N_48657,N_47630,N_47164);
or U48658 (N_48658,N_47408,N_47419);
xor U48659 (N_48659,N_47220,N_47818);
and U48660 (N_48660,N_47327,N_47670);
or U48661 (N_48661,N_47374,N_47593);
and U48662 (N_48662,N_47428,N_47026);
xnor U48663 (N_48663,N_47157,N_47115);
or U48664 (N_48664,N_47240,N_47935);
and U48665 (N_48665,N_47830,N_47389);
and U48666 (N_48666,N_47108,N_47956);
nor U48667 (N_48667,N_47072,N_47659);
or U48668 (N_48668,N_47099,N_47770);
xor U48669 (N_48669,N_47144,N_47019);
xor U48670 (N_48670,N_47719,N_47927);
and U48671 (N_48671,N_47706,N_47957);
nor U48672 (N_48672,N_47534,N_47743);
xnor U48673 (N_48673,N_47981,N_47728);
nor U48674 (N_48674,N_47160,N_47746);
or U48675 (N_48675,N_47333,N_47494);
or U48676 (N_48676,N_47208,N_47943);
nand U48677 (N_48677,N_47551,N_47477);
and U48678 (N_48678,N_47681,N_47559);
nand U48679 (N_48679,N_47710,N_47125);
and U48680 (N_48680,N_47490,N_47031);
nand U48681 (N_48681,N_47145,N_47531);
nand U48682 (N_48682,N_47272,N_47894);
nand U48683 (N_48683,N_47856,N_47933);
nor U48684 (N_48684,N_47526,N_47145);
xor U48685 (N_48685,N_47154,N_47156);
and U48686 (N_48686,N_47837,N_47592);
nor U48687 (N_48687,N_47887,N_47072);
nor U48688 (N_48688,N_47493,N_47600);
nand U48689 (N_48689,N_47742,N_47606);
xnor U48690 (N_48690,N_47690,N_47831);
or U48691 (N_48691,N_47429,N_47621);
or U48692 (N_48692,N_47380,N_47264);
xnor U48693 (N_48693,N_47030,N_47639);
nand U48694 (N_48694,N_47269,N_47202);
and U48695 (N_48695,N_47031,N_47888);
and U48696 (N_48696,N_47564,N_47417);
nor U48697 (N_48697,N_47653,N_47135);
xor U48698 (N_48698,N_47479,N_47727);
or U48699 (N_48699,N_47879,N_47249);
xnor U48700 (N_48700,N_47439,N_47123);
xor U48701 (N_48701,N_47262,N_47995);
xnor U48702 (N_48702,N_47288,N_47133);
nor U48703 (N_48703,N_47408,N_47341);
nand U48704 (N_48704,N_47356,N_47991);
or U48705 (N_48705,N_47601,N_47062);
nand U48706 (N_48706,N_47141,N_47214);
or U48707 (N_48707,N_47716,N_47044);
xnor U48708 (N_48708,N_47293,N_47250);
nor U48709 (N_48709,N_47229,N_47197);
or U48710 (N_48710,N_47683,N_47257);
and U48711 (N_48711,N_47209,N_47796);
nor U48712 (N_48712,N_47898,N_47058);
xor U48713 (N_48713,N_47034,N_47824);
xor U48714 (N_48714,N_47500,N_47440);
nor U48715 (N_48715,N_47010,N_47654);
xor U48716 (N_48716,N_47767,N_47156);
nor U48717 (N_48717,N_47620,N_47110);
and U48718 (N_48718,N_47736,N_47713);
or U48719 (N_48719,N_47105,N_47072);
nor U48720 (N_48720,N_47240,N_47679);
xor U48721 (N_48721,N_47424,N_47472);
nand U48722 (N_48722,N_47926,N_47879);
and U48723 (N_48723,N_47657,N_47423);
xnor U48724 (N_48724,N_47708,N_47156);
or U48725 (N_48725,N_47897,N_47122);
or U48726 (N_48726,N_47937,N_47950);
and U48727 (N_48727,N_47376,N_47448);
nor U48728 (N_48728,N_47122,N_47747);
nand U48729 (N_48729,N_47909,N_47671);
nor U48730 (N_48730,N_47824,N_47208);
and U48731 (N_48731,N_47578,N_47752);
nor U48732 (N_48732,N_47293,N_47269);
or U48733 (N_48733,N_47922,N_47081);
nor U48734 (N_48734,N_47149,N_47425);
and U48735 (N_48735,N_47095,N_47307);
nand U48736 (N_48736,N_47222,N_47492);
or U48737 (N_48737,N_47077,N_47091);
xnor U48738 (N_48738,N_47062,N_47129);
xor U48739 (N_48739,N_47837,N_47805);
or U48740 (N_48740,N_47001,N_47491);
xnor U48741 (N_48741,N_47140,N_47383);
xor U48742 (N_48742,N_47593,N_47396);
nor U48743 (N_48743,N_47333,N_47334);
nand U48744 (N_48744,N_47655,N_47228);
nor U48745 (N_48745,N_47772,N_47577);
or U48746 (N_48746,N_47141,N_47170);
nand U48747 (N_48747,N_47107,N_47396);
and U48748 (N_48748,N_47165,N_47310);
xor U48749 (N_48749,N_47725,N_47609);
and U48750 (N_48750,N_47593,N_47185);
or U48751 (N_48751,N_47408,N_47334);
and U48752 (N_48752,N_47637,N_47301);
or U48753 (N_48753,N_47293,N_47373);
or U48754 (N_48754,N_47282,N_47439);
nor U48755 (N_48755,N_47487,N_47285);
or U48756 (N_48756,N_47224,N_47835);
nor U48757 (N_48757,N_47334,N_47350);
or U48758 (N_48758,N_47316,N_47928);
xor U48759 (N_48759,N_47255,N_47682);
or U48760 (N_48760,N_47261,N_47186);
nand U48761 (N_48761,N_47750,N_47081);
nand U48762 (N_48762,N_47342,N_47417);
or U48763 (N_48763,N_47657,N_47833);
and U48764 (N_48764,N_47374,N_47210);
nor U48765 (N_48765,N_47657,N_47011);
xnor U48766 (N_48766,N_47069,N_47758);
and U48767 (N_48767,N_47566,N_47767);
nand U48768 (N_48768,N_47523,N_47252);
or U48769 (N_48769,N_47000,N_47337);
or U48770 (N_48770,N_47123,N_47083);
xor U48771 (N_48771,N_47141,N_47583);
or U48772 (N_48772,N_47554,N_47992);
nand U48773 (N_48773,N_47133,N_47986);
or U48774 (N_48774,N_47059,N_47850);
and U48775 (N_48775,N_47605,N_47460);
or U48776 (N_48776,N_47289,N_47991);
nor U48777 (N_48777,N_47453,N_47511);
and U48778 (N_48778,N_47083,N_47038);
nor U48779 (N_48779,N_47368,N_47167);
nor U48780 (N_48780,N_47620,N_47146);
or U48781 (N_48781,N_47441,N_47831);
xnor U48782 (N_48782,N_47383,N_47679);
and U48783 (N_48783,N_47305,N_47689);
xor U48784 (N_48784,N_47994,N_47037);
and U48785 (N_48785,N_47521,N_47375);
nor U48786 (N_48786,N_47590,N_47865);
or U48787 (N_48787,N_47817,N_47028);
xor U48788 (N_48788,N_47843,N_47559);
or U48789 (N_48789,N_47062,N_47856);
nor U48790 (N_48790,N_47081,N_47442);
or U48791 (N_48791,N_47624,N_47684);
and U48792 (N_48792,N_47990,N_47026);
nand U48793 (N_48793,N_47387,N_47969);
nor U48794 (N_48794,N_47706,N_47346);
and U48795 (N_48795,N_47387,N_47071);
or U48796 (N_48796,N_47448,N_47393);
xnor U48797 (N_48797,N_47765,N_47741);
xor U48798 (N_48798,N_47966,N_47156);
nor U48799 (N_48799,N_47309,N_47294);
or U48800 (N_48800,N_47502,N_47754);
nor U48801 (N_48801,N_47846,N_47027);
nor U48802 (N_48802,N_47062,N_47862);
nor U48803 (N_48803,N_47682,N_47898);
or U48804 (N_48804,N_47665,N_47585);
nor U48805 (N_48805,N_47326,N_47792);
xnor U48806 (N_48806,N_47292,N_47413);
nand U48807 (N_48807,N_47602,N_47281);
nand U48808 (N_48808,N_47502,N_47726);
or U48809 (N_48809,N_47355,N_47934);
nor U48810 (N_48810,N_47879,N_47157);
nand U48811 (N_48811,N_47262,N_47163);
nor U48812 (N_48812,N_47536,N_47014);
or U48813 (N_48813,N_47656,N_47476);
nand U48814 (N_48814,N_47586,N_47010);
or U48815 (N_48815,N_47752,N_47698);
nand U48816 (N_48816,N_47979,N_47089);
or U48817 (N_48817,N_47180,N_47862);
or U48818 (N_48818,N_47643,N_47308);
xor U48819 (N_48819,N_47455,N_47117);
nor U48820 (N_48820,N_47227,N_47059);
or U48821 (N_48821,N_47621,N_47661);
xor U48822 (N_48822,N_47317,N_47201);
and U48823 (N_48823,N_47368,N_47206);
nor U48824 (N_48824,N_47955,N_47115);
and U48825 (N_48825,N_47582,N_47255);
or U48826 (N_48826,N_47322,N_47045);
or U48827 (N_48827,N_47757,N_47042);
or U48828 (N_48828,N_47718,N_47185);
xnor U48829 (N_48829,N_47173,N_47128);
xnor U48830 (N_48830,N_47117,N_47556);
or U48831 (N_48831,N_47555,N_47018);
nand U48832 (N_48832,N_47215,N_47167);
or U48833 (N_48833,N_47119,N_47444);
and U48834 (N_48834,N_47784,N_47097);
xor U48835 (N_48835,N_47361,N_47414);
or U48836 (N_48836,N_47354,N_47039);
or U48837 (N_48837,N_47714,N_47129);
or U48838 (N_48838,N_47274,N_47252);
nor U48839 (N_48839,N_47500,N_47486);
nand U48840 (N_48840,N_47577,N_47370);
xor U48841 (N_48841,N_47866,N_47214);
nand U48842 (N_48842,N_47180,N_47920);
and U48843 (N_48843,N_47642,N_47412);
or U48844 (N_48844,N_47456,N_47384);
xnor U48845 (N_48845,N_47919,N_47931);
xnor U48846 (N_48846,N_47813,N_47681);
or U48847 (N_48847,N_47354,N_47674);
nor U48848 (N_48848,N_47491,N_47638);
xor U48849 (N_48849,N_47917,N_47208);
and U48850 (N_48850,N_47527,N_47905);
nor U48851 (N_48851,N_47097,N_47810);
nor U48852 (N_48852,N_47761,N_47498);
nand U48853 (N_48853,N_47435,N_47539);
and U48854 (N_48854,N_47705,N_47538);
or U48855 (N_48855,N_47173,N_47524);
or U48856 (N_48856,N_47916,N_47886);
and U48857 (N_48857,N_47367,N_47193);
and U48858 (N_48858,N_47745,N_47665);
and U48859 (N_48859,N_47040,N_47387);
xnor U48860 (N_48860,N_47780,N_47590);
nor U48861 (N_48861,N_47553,N_47691);
xnor U48862 (N_48862,N_47621,N_47533);
xnor U48863 (N_48863,N_47869,N_47993);
or U48864 (N_48864,N_47465,N_47101);
and U48865 (N_48865,N_47098,N_47418);
nor U48866 (N_48866,N_47427,N_47090);
nand U48867 (N_48867,N_47887,N_47432);
and U48868 (N_48868,N_47438,N_47696);
nand U48869 (N_48869,N_47343,N_47208);
and U48870 (N_48870,N_47321,N_47287);
and U48871 (N_48871,N_47538,N_47968);
and U48872 (N_48872,N_47275,N_47116);
nor U48873 (N_48873,N_47813,N_47453);
or U48874 (N_48874,N_47327,N_47580);
and U48875 (N_48875,N_47310,N_47872);
xor U48876 (N_48876,N_47466,N_47648);
nand U48877 (N_48877,N_47372,N_47504);
nor U48878 (N_48878,N_47077,N_47779);
or U48879 (N_48879,N_47279,N_47202);
nand U48880 (N_48880,N_47396,N_47062);
xor U48881 (N_48881,N_47605,N_47220);
nand U48882 (N_48882,N_47705,N_47222);
nand U48883 (N_48883,N_47796,N_47654);
xnor U48884 (N_48884,N_47703,N_47816);
and U48885 (N_48885,N_47671,N_47593);
or U48886 (N_48886,N_47334,N_47716);
nand U48887 (N_48887,N_47432,N_47643);
xnor U48888 (N_48888,N_47231,N_47968);
nor U48889 (N_48889,N_47778,N_47476);
and U48890 (N_48890,N_47525,N_47054);
xnor U48891 (N_48891,N_47893,N_47502);
or U48892 (N_48892,N_47942,N_47578);
xor U48893 (N_48893,N_47956,N_47597);
nand U48894 (N_48894,N_47877,N_47801);
nand U48895 (N_48895,N_47355,N_47605);
and U48896 (N_48896,N_47720,N_47242);
nor U48897 (N_48897,N_47423,N_47785);
and U48898 (N_48898,N_47817,N_47697);
or U48899 (N_48899,N_47868,N_47804);
xnor U48900 (N_48900,N_47953,N_47466);
xnor U48901 (N_48901,N_47925,N_47735);
and U48902 (N_48902,N_47789,N_47529);
and U48903 (N_48903,N_47000,N_47836);
nand U48904 (N_48904,N_47924,N_47317);
nand U48905 (N_48905,N_47315,N_47691);
and U48906 (N_48906,N_47964,N_47799);
nand U48907 (N_48907,N_47257,N_47215);
xor U48908 (N_48908,N_47208,N_47931);
nand U48909 (N_48909,N_47699,N_47706);
or U48910 (N_48910,N_47047,N_47530);
or U48911 (N_48911,N_47691,N_47985);
xnor U48912 (N_48912,N_47440,N_47499);
and U48913 (N_48913,N_47097,N_47015);
or U48914 (N_48914,N_47227,N_47060);
nand U48915 (N_48915,N_47500,N_47475);
xnor U48916 (N_48916,N_47224,N_47467);
nand U48917 (N_48917,N_47128,N_47221);
or U48918 (N_48918,N_47932,N_47816);
xnor U48919 (N_48919,N_47682,N_47819);
nand U48920 (N_48920,N_47227,N_47363);
xor U48921 (N_48921,N_47129,N_47305);
nand U48922 (N_48922,N_47160,N_47869);
and U48923 (N_48923,N_47605,N_47240);
nand U48924 (N_48924,N_47564,N_47164);
nor U48925 (N_48925,N_47125,N_47651);
and U48926 (N_48926,N_47279,N_47332);
nor U48927 (N_48927,N_47881,N_47377);
nand U48928 (N_48928,N_47895,N_47338);
nor U48929 (N_48929,N_47547,N_47154);
nor U48930 (N_48930,N_47212,N_47511);
nor U48931 (N_48931,N_47248,N_47446);
and U48932 (N_48932,N_47447,N_47499);
or U48933 (N_48933,N_47551,N_47626);
nor U48934 (N_48934,N_47542,N_47552);
and U48935 (N_48935,N_47654,N_47308);
nor U48936 (N_48936,N_47911,N_47707);
or U48937 (N_48937,N_47662,N_47395);
nor U48938 (N_48938,N_47833,N_47598);
and U48939 (N_48939,N_47693,N_47796);
and U48940 (N_48940,N_47319,N_47211);
and U48941 (N_48941,N_47157,N_47097);
or U48942 (N_48942,N_47651,N_47678);
nor U48943 (N_48943,N_47155,N_47204);
or U48944 (N_48944,N_47355,N_47047);
or U48945 (N_48945,N_47236,N_47121);
and U48946 (N_48946,N_47249,N_47678);
and U48947 (N_48947,N_47903,N_47395);
xnor U48948 (N_48948,N_47083,N_47760);
xor U48949 (N_48949,N_47340,N_47682);
and U48950 (N_48950,N_47731,N_47905);
nand U48951 (N_48951,N_47415,N_47261);
or U48952 (N_48952,N_47222,N_47014);
xnor U48953 (N_48953,N_47260,N_47936);
nor U48954 (N_48954,N_47896,N_47131);
and U48955 (N_48955,N_47670,N_47639);
and U48956 (N_48956,N_47045,N_47151);
and U48957 (N_48957,N_47859,N_47745);
or U48958 (N_48958,N_47529,N_47727);
or U48959 (N_48959,N_47138,N_47611);
or U48960 (N_48960,N_47188,N_47946);
nand U48961 (N_48961,N_47152,N_47188);
nor U48962 (N_48962,N_47429,N_47770);
nand U48963 (N_48963,N_47893,N_47238);
or U48964 (N_48964,N_47904,N_47567);
nand U48965 (N_48965,N_47992,N_47531);
or U48966 (N_48966,N_47198,N_47189);
and U48967 (N_48967,N_47145,N_47267);
nand U48968 (N_48968,N_47313,N_47893);
and U48969 (N_48969,N_47082,N_47983);
or U48970 (N_48970,N_47337,N_47346);
xor U48971 (N_48971,N_47179,N_47262);
nor U48972 (N_48972,N_47957,N_47008);
and U48973 (N_48973,N_47228,N_47132);
nand U48974 (N_48974,N_47966,N_47227);
xnor U48975 (N_48975,N_47045,N_47996);
nand U48976 (N_48976,N_47723,N_47342);
and U48977 (N_48977,N_47379,N_47844);
xnor U48978 (N_48978,N_47193,N_47570);
nor U48979 (N_48979,N_47083,N_47523);
and U48980 (N_48980,N_47383,N_47753);
nand U48981 (N_48981,N_47961,N_47473);
and U48982 (N_48982,N_47217,N_47655);
nor U48983 (N_48983,N_47869,N_47755);
xor U48984 (N_48984,N_47093,N_47752);
and U48985 (N_48985,N_47149,N_47640);
and U48986 (N_48986,N_47761,N_47913);
nand U48987 (N_48987,N_47425,N_47957);
and U48988 (N_48988,N_47423,N_47257);
and U48989 (N_48989,N_47628,N_47101);
nor U48990 (N_48990,N_47462,N_47668);
xnor U48991 (N_48991,N_47105,N_47006);
or U48992 (N_48992,N_47751,N_47746);
nor U48993 (N_48993,N_47508,N_47180);
nand U48994 (N_48994,N_47310,N_47968);
nor U48995 (N_48995,N_47521,N_47727);
and U48996 (N_48996,N_47677,N_47298);
nor U48997 (N_48997,N_47143,N_47632);
xor U48998 (N_48998,N_47409,N_47743);
nor U48999 (N_48999,N_47647,N_47472);
and U49000 (N_49000,N_48666,N_48514);
nor U49001 (N_49001,N_48534,N_48753);
or U49002 (N_49002,N_48496,N_48809);
and U49003 (N_49003,N_48600,N_48213);
or U49004 (N_49004,N_48913,N_48491);
xnor U49005 (N_49005,N_48970,N_48106);
nor U49006 (N_49006,N_48903,N_48900);
and U49007 (N_49007,N_48373,N_48902);
xor U49008 (N_49008,N_48751,N_48549);
or U49009 (N_49009,N_48065,N_48450);
nand U49010 (N_49010,N_48570,N_48252);
xor U49011 (N_49011,N_48795,N_48104);
or U49012 (N_49012,N_48352,N_48303);
xor U49013 (N_49013,N_48461,N_48687);
xnor U49014 (N_49014,N_48827,N_48038);
nand U49015 (N_49015,N_48342,N_48931);
nor U49016 (N_49016,N_48710,N_48173);
nor U49017 (N_49017,N_48770,N_48925);
nand U49018 (N_49018,N_48228,N_48441);
and U49019 (N_49019,N_48421,N_48611);
and U49020 (N_49020,N_48608,N_48553);
and U49021 (N_49021,N_48136,N_48046);
nand U49022 (N_49022,N_48143,N_48281);
xnor U49023 (N_49023,N_48322,N_48802);
nand U49024 (N_49024,N_48062,N_48616);
or U49025 (N_49025,N_48420,N_48327);
nor U49026 (N_49026,N_48187,N_48276);
and U49027 (N_49027,N_48750,N_48885);
nor U49028 (N_49028,N_48166,N_48181);
nand U49029 (N_49029,N_48008,N_48694);
and U49030 (N_49030,N_48575,N_48851);
xor U49031 (N_49031,N_48305,N_48004);
and U49032 (N_49032,N_48935,N_48587);
xor U49033 (N_49033,N_48701,N_48888);
or U49034 (N_49034,N_48444,N_48474);
and U49035 (N_49035,N_48357,N_48929);
nor U49036 (N_49036,N_48560,N_48153);
nor U49037 (N_49037,N_48845,N_48740);
nand U49038 (N_49038,N_48861,N_48384);
and U49039 (N_49039,N_48140,N_48977);
xor U49040 (N_49040,N_48240,N_48400);
and U49041 (N_49041,N_48531,N_48957);
nand U49042 (N_49042,N_48500,N_48951);
xor U49043 (N_49043,N_48264,N_48224);
or U49044 (N_49044,N_48538,N_48773);
nand U49045 (N_49045,N_48998,N_48026);
nand U49046 (N_49046,N_48088,N_48048);
or U49047 (N_49047,N_48547,N_48675);
and U49048 (N_49048,N_48348,N_48454);
nor U49049 (N_49049,N_48346,N_48719);
nand U49050 (N_49050,N_48519,N_48179);
xor U49051 (N_49051,N_48162,N_48163);
nand U49052 (N_49052,N_48098,N_48016);
and U49053 (N_49053,N_48457,N_48979);
xor U49054 (N_49054,N_48854,N_48294);
nor U49055 (N_49055,N_48639,N_48101);
nand U49056 (N_49056,N_48437,N_48172);
nor U49057 (N_49057,N_48954,N_48190);
nor U49058 (N_49058,N_48697,N_48473);
nand U49059 (N_49059,N_48508,N_48337);
xor U49060 (N_49060,N_48061,N_48222);
nor U49061 (N_49061,N_48469,N_48145);
or U49062 (N_49062,N_48664,N_48070);
and U49063 (N_49063,N_48386,N_48476);
and U49064 (N_49064,N_48663,N_48270);
and U49065 (N_49065,N_48040,N_48049);
or U49066 (N_49066,N_48653,N_48927);
or U49067 (N_49067,N_48440,N_48909);
or U49068 (N_49068,N_48882,N_48391);
or U49069 (N_49069,N_48335,N_48219);
nor U49070 (N_49070,N_48746,N_48878);
nand U49071 (N_49071,N_48269,N_48843);
or U49072 (N_49072,N_48949,N_48898);
nand U49073 (N_49073,N_48170,N_48388);
xnor U49074 (N_49074,N_48124,N_48520);
nor U49075 (N_49075,N_48555,N_48074);
or U49076 (N_49076,N_48550,N_48881);
xnor U49077 (N_49077,N_48063,N_48915);
or U49078 (N_49078,N_48150,N_48435);
nor U49079 (N_49079,N_48051,N_48695);
nand U49080 (N_49080,N_48486,N_48083);
or U49081 (N_49081,N_48054,N_48811);
xnor U49082 (N_49082,N_48632,N_48956);
nor U49083 (N_49083,N_48546,N_48076);
or U49084 (N_49084,N_48947,N_48395);
nand U49085 (N_49085,N_48418,N_48928);
or U49086 (N_49086,N_48527,N_48196);
xor U49087 (N_49087,N_48626,N_48498);
nand U49088 (N_49088,N_48064,N_48630);
nand U49089 (N_49089,N_48573,N_48238);
and U49090 (N_49090,N_48297,N_48960);
or U49091 (N_49091,N_48250,N_48197);
nor U49092 (N_49092,N_48880,N_48168);
nand U49093 (N_49093,N_48073,N_48955);
nor U49094 (N_49094,N_48620,N_48409);
nand U49095 (N_49095,N_48594,N_48146);
nand U49096 (N_49096,N_48100,N_48952);
nor U49097 (N_49097,N_48522,N_48152);
xor U49098 (N_49098,N_48511,N_48011);
nand U49099 (N_49099,N_48981,N_48612);
xor U49100 (N_49100,N_48483,N_48938);
or U49101 (N_49101,N_48313,N_48732);
xor U49102 (N_49102,N_48381,N_48462);
xor U49103 (N_49103,N_48636,N_48923);
xor U49104 (N_49104,N_48245,N_48424);
xnor U49105 (N_49105,N_48368,N_48926);
and U49106 (N_49106,N_48225,N_48661);
nor U49107 (N_49107,N_48304,N_48438);
and U49108 (N_49108,N_48963,N_48962);
and U49109 (N_49109,N_48579,N_48082);
nor U49110 (N_49110,N_48985,N_48964);
or U49111 (N_49111,N_48353,N_48613);
xor U49112 (N_49112,N_48984,N_48633);
nand U49113 (N_49113,N_48236,N_48904);
or U49114 (N_49114,N_48832,N_48265);
nand U49115 (N_49115,N_48220,N_48988);
and U49116 (N_49116,N_48227,N_48488);
and U49117 (N_49117,N_48212,N_48109);
xor U49118 (N_49118,N_48967,N_48422);
or U49119 (N_49119,N_48261,N_48071);
nand U49120 (N_49120,N_48433,N_48393);
nor U49121 (N_49121,N_48300,N_48248);
and U49122 (N_49122,N_48918,N_48119);
nor U49123 (N_49123,N_48157,N_48115);
nand U49124 (N_49124,N_48234,N_48356);
nor U49125 (N_49125,N_48079,N_48336);
or U49126 (N_49126,N_48419,N_48058);
nand U49127 (N_49127,N_48816,N_48922);
or U49128 (N_49128,N_48521,N_48426);
nand U49129 (N_49129,N_48287,N_48141);
nor U49130 (N_49130,N_48286,N_48897);
nand U49131 (N_49131,N_48586,N_48721);
xnor U49132 (N_49132,N_48764,N_48097);
and U49133 (N_49133,N_48425,N_48863);
nor U49134 (N_49134,N_48599,N_48595);
nor U49135 (N_49135,N_48370,N_48862);
and U49136 (N_49136,N_48059,N_48315);
and U49137 (N_49137,N_48278,N_48708);
nor U49138 (N_49138,N_48293,N_48249);
and U49139 (N_49139,N_48602,N_48841);
xor U49140 (N_49140,N_48013,N_48257);
or U49141 (N_49141,N_48510,N_48509);
xnor U49142 (N_49142,N_48349,N_48323);
nor U49143 (N_49143,N_48601,N_48911);
nand U49144 (N_49144,N_48057,N_48413);
or U49145 (N_49145,N_48518,N_48397);
xnor U49146 (N_49146,N_48254,N_48377);
or U49147 (N_49147,N_48333,N_48012);
and U49148 (N_49148,N_48939,N_48908);
nor U49149 (N_49149,N_48582,N_48699);
nand U49150 (N_49150,N_48554,N_48712);
nor U49151 (N_49151,N_48975,N_48670);
and U49152 (N_49152,N_48319,N_48330);
and U49153 (N_49153,N_48855,N_48536);
nor U49154 (N_49154,N_48644,N_48472);
nor U49155 (N_49155,N_48756,N_48379);
xnor U49156 (N_49156,N_48316,N_48726);
xnor U49157 (N_49157,N_48369,N_48321);
or U49158 (N_49158,N_48598,N_48134);
nor U49159 (N_49159,N_48090,N_48635);
and U49160 (N_49160,N_48320,N_48730);
xor U49161 (N_49161,N_48609,N_48188);
and U49162 (N_49162,N_48762,N_48255);
xnor U49163 (N_49163,N_48271,N_48408);
nor U49164 (N_49164,N_48788,N_48385);
nand U49165 (N_49165,N_48752,N_48724);
nand U49166 (N_49166,N_48544,N_48530);
and U49167 (N_49167,N_48195,N_48912);
nand U49168 (N_49168,N_48649,N_48765);
xnor U49169 (N_49169,N_48785,N_48551);
xnor U49170 (N_49170,N_48763,N_48492);
or U49171 (N_49171,N_48541,N_48571);
nor U49172 (N_49172,N_48731,N_48358);
and U49173 (N_49173,N_48452,N_48506);
or U49174 (N_49174,N_48858,N_48623);
xor U49175 (N_49175,N_48799,N_48468);
xnor U49176 (N_49176,N_48482,N_48275);
nor U49177 (N_49177,N_48883,N_48189);
nor U49178 (N_49178,N_48332,N_48113);
or U49179 (N_49179,N_48365,N_48993);
nand U49180 (N_49180,N_48637,N_48375);
and U49181 (N_49181,N_48801,N_48047);
nor U49182 (N_49182,N_48971,N_48149);
xnor U49183 (N_49183,N_48629,N_48820);
xnor U49184 (N_49184,N_48127,N_48010);
nor U49185 (N_49185,N_48007,N_48091);
or U49186 (N_49186,N_48487,N_48338);
or U49187 (N_49187,N_48658,N_48060);
nor U49188 (N_49188,N_48873,N_48376);
and U49189 (N_49189,N_48345,N_48133);
xor U49190 (N_49190,N_48449,N_48754);
nor U49191 (N_49191,N_48737,N_48154);
and U49192 (N_49192,N_48705,N_48259);
xnor U49193 (N_49193,N_48410,N_48000);
and U49194 (N_49194,N_48481,N_48680);
nor U49195 (N_49195,N_48273,N_48703);
nand U49196 (N_49196,N_48849,N_48148);
and U49197 (N_49197,N_48879,N_48577);
and U49198 (N_49198,N_48470,N_48648);
nor U49199 (N_49199,N_48806,N_48009);
and U49200 (N_49200,N_48621,N_48308);
xnor U49201 (N_49201,N_48976,N_48362);
nand U49202 (N_49202,N_48990,N_48326);
xnor U49203 (N_49203,N_48242,N_48822);
nor U49204 (N_49204,N_48736,N_48757);
nor U49205 (N_49205,N_48184,N_48738);
and U49206 (N_49206,N_48796,N_48036);
or U49207 (N_49207,N_48745,N_48607);
xor U49208 (N_49208,N_48574,N_48974);
and U49209 (N_49209,N_48445,N_48485);
or U49210 (N_49210,N_48256,N_48285);
or U49211 (N_49211,N_48859,N_48218);
and U49212 (N_49212,N_48006,N_48033);
or U49213 (N_49213,N_48117,N_48589);
nor U49214 (N_49214,N_48089,N_48371);
nand U49215 (N_49215,N_48673,N_48451);
xor U49216 (N_49216,N_48053,N_48235);
nor U49217 (N_49217,N_48361,N_48367);
and U49218 (N_49218,N_48593,N_48355);
nor U49219 (N_49219,N_48994,N_48032);
and U49220 (N_49220,N_48704,N_48122);
xor U49221 (N_49221,N_48453,N_48944);
or U49222 (N_49222,N_48556,N_48041);
nand U49223 (N_49223,N_48792,N_48894);
nand U49224 (N_49224,N_48233,N_48210);
nand U49225 (N_49225,N_48480,N_48776);
nand U49226 (N_49226,N_48340,N_48202);
nor U49227 (N_49227,N_48789,N_48512);
or U49228 (N_49228,N_48605,N_48842);
nand U49229 (N_49229,N_48847,N_48005);
or U49230 (N_49230,N_48290,N_48713);
xnor U49231 (N_49231,N_48359,N_48907);
or U49232 (N_49232,N_48545,N_48786);
xor U49233 (N_49233,N_48456,N_48344);
nand U49234 (N_49234,N_48982,N_48874);
nand U49235 (N_49235,N_48299,N_48941);
and U49236 (N_49236,N_48229,N_48158);
nand U49237 (N_49237,N_48934,N_48436);
xor U49238 (N_49238,N_48965,N_48211);
and U49239 (N_49239,N_48432,N_48996);
nand U49240 (N_49240,N_48997,N_48564);
or U49241 (N_49241,N_48728,N_48537);
or U49242 (N_49242,N_48516,N_48031);
and U49243 (N_49243,N_48077,N_48258);
nand U49244 (N_49244,N_48884,N_48568);
nand U49245 (N_49245,N_48475,N_48110);
or U49246 (N_49246,N_48347,N_48830);
nor U49247 (N_49247,N_48204,N_48698);
nand U49248 (N_49248,N_48775,N_48583);
or U49249 (N_49249,N_48787,N_48479);
xor U49250 (N_49250,N_48107,N_48209);
nor U49251 (N_49251,N_48099,N_48654);
nand U49252 (N_49252,N_48584,N_48590);
and U49253 (N_49253,N_48552,N_48852);
nor U49254 (N_49254,N_48237,N_48804);
nor U49255 (N_49255,N_48194,N_48423);
nand U49256 (N_49256,N_48018,N_48042);
nor U49257 (N_49257,N_48251,N_48991);
xor U49258 (N_49258,N_48191,N_48727);
nand U49259 (N_49259,N_48180,N_48241);
nor U49260 (N_49260,N_48945,N_48857);
nand U49261 (N_49261,N_48085,N_48489);
nand U49262 (N_49262,N_48864,N_48690);
xor U49263 (N_49263,N_48364,N_48813);
or U49264 (N_49264,N_48328,N_48095);
nand U49265 (N_49265,N_48614,N_48147);
or U49266 (N_49266,N_48182,N_48646);
nor U49267 (N_49267,N_48442,N_48374);
and U49268 (N_49268,N_48592,N_48382);
nor U49269 (N_49269,N_48354,N_48282);
and U49270 (N_49270,N_48120,N_48341);
nand U49271 (N_49271,N_48428,N_48615);
nor U49272 (N_49272,N_48019,N_48958);
nor U49273 (N_49273,N_48490,N_48893);
nand U49274 (N_49274,N_48688,N_48114);
nand U49275 (N_49275,N_48777,N_48023);
and U49276 (N_49276,N_48950,N_48803);
and U49277 (N_49277,N_48890,N_48284);
nand U49278 (N_49278,N_48129,N_48742);
xor U49279 (N_49279,N_48138,N_48467);
and U49280 (N_49280,N_48749,N_48378);
and U49281 (N_49281,N_48403,N_48797);
xnor U49282 (N_49282,N_48072,N_48302);
and U49283 (N_49283,N_48798,N_48723);
and U49284 (N_49284,N_48891,N_48659);
nand U49285 (N_49285,N_48668,N_48910);
or U49286 (N_49286,N_48411,N_48856);
nor U49287 (N_49287,N_48360,N_48768);
or U49288 (N_49288,N_48681,N_48696);
or U49289 (N_49289,N_48144,N_48266);
or U49290 (N_49290,N_48747,N_48755);
nor U49291 (N_49291,N_48683,N_48831);
nand U49292 (N_49292,N_48105,N_48669);
xor U49293 (N_49293,N_48678,N_48706);
xor U49294 (N_49294,N_48933,N_48406);
nor U49295 (N_49295,N_48513,N_48532);
nand U49296 (N_49296,N_48231,N_48260);
nor U49297 (N_49297,N_48989,N_48735);
and U49298 (N_49298,N_48709,N_48263);
xnor U49299 (N_49299,N_48494,N_48244);
xor U49300 (N_49300,N_48020,N_48691);
xor U49301 (N_49301,N_48142,N_48387);
and U49302 (N_49302,N_48790,N_48643);
nor U49303 (N_49303,N_48094,N_48183);
and U49304 (N_49304,N_48528,N_48292);
nand U49305 (N_49305,N_48200,N_48096);
and U49306 (N_49306,N_48325,N_48940);
xor U49307 (N_49307,N_48992,N_48921);
and U49308 (N_49308,N_48298,N_48800);
nand U49309 (N_49309,N_48662,N_48622);
xor U49310 (N_49310,N_48959,N_48930);
and U49311 (N_49311,N_48999,N_48734);
nand U49312 (N_49312,N_48216,N_48034);
nand U49313 (N_49313,N_48176,N_48657);
nor U49314 (N_49314,N_48567,N_48446);
xnor U49315 (N_49315,N_48390,N_48682);
xnor U49316 (N_49316,N_48507,N_48092);
xor U49317 (N_49317,N_48447,N_48867);
nor U49318 (N_49318,N_48484,N_48192);
xor U49319 (N_49319,N_48833,N_48201);
nand U49320 (N_49320,N_48131,N_48674);
or U49321 (N_49321,N_48980,N_48924);
nand U49322 (N_49322,N_48716,N_48539);
and U49323 (N_49323,N_48718,N_48618);
xnor U49324 (N_49324,N_48686,N_48001);
nor U49325 (N_49325,N_48987,N_48280);
nor U49326 (N_49326,N_48875,N_48558);
nor U49327 (N_49327,N_48937,N_48837);
nand U49328 (N_49328,N_48164,N_48246);
and U49329 (N_49329,N_48892,N_48853);
nor U49330 (N_49330,N_48078,N_48022);
and U49331 (N_49331,N_48239,N_48986);
nor U49332 (N_49332,N_48744,N_48283);
nor U49333 (N_49333,N_48784,N_48093);
or U49334 (N_49334,N_48399,N_48203);
and U49335 (N_49335,N_48651,N_48103);
and U49336 (N_49336,N_48156,N_48068);
nand U49337 (N_49337,N_48983,N_48819);
xnor U49338 (N_49338,N_48081,N_48112);
and U49339 (N_49339,N_48052,N_48580);
or U49340 (N_49340,N_48917,N_48279);
xnor U49341 (N_49341,N_48814,N_48230);
nor U49342 (N_49342,N_48717,N_48021);
xnor U49343 (N_49343,N_48459,N_48331);
nor U49344 (N_49344,N_48501,N_48310);
and U49345 (N_49345,N_48017,N_48471);
xor U49346 (N_49346,N_48850,N_48464);
xnor U49347 (N_49347,N_48404,N_48693);
nor U49348 (N_49348,N_48848,N_48306);
xor U49349 (N_49349,N_48953,N_48961);
and U49350 (N_49350,N_48645,N_48808);
nor U49351 (N_49351,N_48366,N_48414);
nand U49352 (N_49352,N_48267,N_48434);
xor U49353 (N_49353,N_48014,N_48178);
xnor U49354 (N_49354,N_48679,N_48037);
nor U49355 (N_49355,N_48030,N_48761);
nor U49356 (N_49356,N_48024,N_48667);
nor U49357 (N_49357,N_48161,N_48606);
or U49358 (N_49358,N_48493,N_48155);
nor U49359 (N_49359,N_48585,N_48692);
nand U49360 (N_49360,N_48039,N_48886);
nand U49361 (N_49361,N_48860,N_48714);
nor U49362 (N_49362,N_48137,N_48372);
nor U49363 (N_49363,N_48624,N_48272);
nand U49364 (N_49364,N_48660,N_48067);
nand U49365 (N_49365,N_48477,N_48504);
nor U49366 (N_49366,N_48221,N_48121);
xor U49367 (N_49367,N_48767,N_48151);
or U49368 (N_49368,N_48919,N_48309);
xor U49369 (N_49369,N_48817,N_48417);
nand U49370 (N_49370,N_48748,N_48655);
and U49371 (N_49371,N_48412,N_48715);
xnor U49372 (N_49372,N_48596,N_48783);
or U49373 (N_49373,N_48995,N_48650);
xor U49374 (N_49374,N_48588,N_48318);
nor U49375 (N_49375,N_48086,N_48215);
xor U49376 (N_49376,N_48407,N_48430);
or U49377 (N_49377,N_48029,N_48311);
nand U49378 (N_49378,N_48836,N_48887);
nor U49379 (N_49379,N_48050,N_48810);
nor U49380 (N_49380,N_48771,N_48415);
nand U49381 (N_49381,N_48314,N_48942);
nor U49382 (N_49382,N_48631,N_48916);
nor U49383 (N_49383,N_48523,N_48563);
xnor U49384 (N_49384,N_48821,N_48572);
nor U49385 (N_49385,N_48834,N_48812);
xor U49386 (N_49386,N_48043,N_48416);
nand U49387 (N_49387,N_48495,N_48642);
xnor U49388 (N_49388,N_48948,N_48169);
xnor U49389 (N_49389,N_48656,N_48055);
xor U49390 (N_49390,N_48296,N_48460);
or U49391 (N_49391,N_48394,N_48126);
or U49392 (N_49392,N_48232,N_48247);
xor U49393 (N_49393,N_48478,N_48289);
and U49394 (N_49394,N_48102,N_48465);
or U49395 (N_49395,N_48872,N_48778);
and U49396 (N_49396,N_48805,N_48253);
or U49397 (N_49397,N_48617,N_48725);
xor U49398 (N_49398,N_48002,N_48439);
nor U49399 (N_49399,N_48758,N_48463);
nand U49400 (N_49400,N_48610,N_48760);
and U49401 (N_49401,N_48274,N_48497);
nor U49402 (N_49402,N_48186,N_48720);
nor U49403 (N_49403,N_48966,N_48317);
xnor U49404 (N_49404,N_48533,N_48581);
or U49405 (N_49405,N_48003,N_48823);
nand U49406 (N_49406,N_48206,N_48401);
and U49407 (N_49407,N_48540,N_48217);
or U49408 (N_49408,N_48877,N_48226);
xnor U49409 (N_49409,N_48329,N_48689);
nor U49410 (N_49410,N_48791,N_48932);
xnor U49411 (N_49411,N_48807,N_48978);
and U49412 (N_49412,N_48535,N_48548);
nor U49413 (N_49413,N_48700,N_48035);
nand U49414 (N_49414,N_48069,N_48135);
and U49415 (N_49415,N_48604,N_48402);
and U49416 (N_49416,N_48628,N_48641);
nor U49417 (N_49417,N_48167,N_48844);
and U49418 (N_49418,N_48524,N_48174);
or U49419 (N_49419,N_48543,N_48936);
and U49420 (N_49420,N_48324,N_48427);
xnor U49421 (N_49421,N_48561,N_48351);
and U49422 (N_49422,N_48307,N_48045);
xor U49423 (N_49423,N_48665,N_48634);
and U49424 (N_49424,N_48044,N_48268);
nor U49425 (N_49425,N_48780,N_48243);
or U49426 (N_49426,N_48108,N_48901);
or U49427 (N_49427,N_48116,N_48739);
or U49428 (N_49428,N_48502,N_48208);
nand U49429 (N_49429,N_48815,N_48128);
or U49430 (N_49430,N_48199,N_48565);
or U49431 (N_49431,N_48779,N_48343);
nand U49432 (N_49432,N_48363,N_48334);
and U49433 (N_49433,N_48896,N_48676);
and U49434 (N_49434,N_48130,N_48625);
nor U49435 (N_49435,N_48825,N_48895);
xor U49436 (N_49436,N_48647,N_48542);
nand U49437 (N_49437,N_48295,N_48899);
nand U49438 (N_49438,N_48868,N_48627);
nand U49439 (N_49439,N_48870,N_48448);
or U49440 (N_49440,N_48392,N_48591);
and U49441 (N_49441,N_48025,N_48671);
nor U49442 (N_49442,N_48027,N_48466);
nor U49443 (N_49443,N_48207,N_48288);
or U49444 (N_49444,N_48741,N_48685);
xor U49445 (N_49445,N_48906,N_48165);
xnor U49446 (N_49446,N_48132,N_48389);
or U49447 (N_49447,N_48566,N_48223);
nand U49448 (N_49448,N_48759,N_48702);
nor U49449 (N_49449,N_48301,N_48015);
or U49450 (N_49450,N_48865,N_48794);
and U49451 (N_49451,N_48111,N_48383);
and U49452 (N_49452,N_48603,N_48943);
and U49453 (N_49453,N_48969,N_48835);
or U49454 (N_49454,N_48866,N_48443);
nand U49455 (N_49455,N_48905,N_48291);
nor U49456 (N_49456,N_48559,N_48968);
and U49457 (N_49457,N_48529,N_48139);
and U49458 (N_49458,N_48840,N_48920);
nand U49459 (N_49459,N_48505,N_48499);
or U49460 (N_49460,N_48125,N_48350);
nor U49461 (N_49461,N_48638,N_48177);
or U49462 (N_49462,N_48946,N_48515);
nand U49463 (N_49463,N_48159,N_48517);
xnor U49464 (N_49464,N_48793,N_48672);
or U49465 (N_49465,N_48455,N_48198);
xor U49466 (N_49466,N_48569,N_48677);
and U49467 (N_49467,N_48576,N_48828);
or U49468 (N_49468,N_48889,N_48729);
nand U49469 (N_49469,N_48525,N_48557);
nand U49470 (N_49470,N_48684,N_48743);
nor U49471 (N_49471,N_48869,N_48619);
nor U49472 (N_49472,N_48056,N_48972);
and U49473 (N_49473,N_48312,N_48818);
and U49474 (N_49474,N_48722,N_48838);
or U49475 (N_49475,N_48080,N_48846);
or U49476 (N_49476,N_48175,N_48277);
and U49477 (N_49477,N_48205,N_48262);
and U49478 (N_49478,N_48084,N_48597);
nand U49479 (N_49479,N_48578,N_48185);
nand U49480 (N_49480,N_48118,N_48829);
nand U49481 (N_49481,N_48640,N_48398);
nand U49482 (N_49482,N_48826,N_48526);
nand U49483 (N_49483,N_48652,N_48839);
nor U49484 (N_49484,N_48711,N_48396);
xor U49485 (N_49485,N_48772,N_48781);
and U49486 (N_49486,N_48707,N_48123);
or U49487 (N_49487,N_48876,N_48871);
nand U49488 (N_49488,N_48782,N_48733);
xor U49489 (N_49489,N_48087,N_48380);
and U49490 (N_49490,N_48973,N_48429);
nand U49491 (N_49491,N_48075,N_48431);
nand U49492 (N_49492,N_48028,N_48824);
and U49493 (N_49493,N_48193,N_48339);
nor U49494 (N_49494,N_48160,N_48066);
nor U49495 (N_49495,N_48914,N_48171);
and U49496 (N_49496,N_48769,N_48774);
nand U49497 (N_49497,N_48503,N_48458);
nor U49498 (N_49498,N_48405,N_48766);
nand U49499 (N_49499,N_48562,N_48214);
xor U49500 (N_49500,N_48883,N_48047);
nor U49501 (N_49501,N_48340,N_48540);
nor U49502 (N_49502,N_48002,N_48359);
nand U49503 (N_49503,N_48556,N_48017);
and U49504 (N_49504,N_48241,N_48750);
or U49505 (N_49505,N_48224,N_48043);
xor U49506 (N_49506,N_48764,N_48343);
nand U49507 (N_49507,N_48567,N_48998);
and U49508 (N_49508,N_48554,N_48358);
nand U49509 (N_49509,N_48027,N_48386);
and U49510 (N_49510,N_48677,N_48367);
and U49511 (N_49511,N_48267,N_48185);
xnor U49512 (N_49512,N_48245,N_48804);
nor U49513 (N_49513,N_48794,N_48595);
or U49514 (N_49514,N_48554,N_48504);
xor U49515 (N_49515,N_48017,N_48189);
nand U49516 (N_49516,N_48696,N_48973);
xnor U49517 (N_49517,N_48815,N_48997);
and U49518 (N_49518,N_48662,N_48112);
nor U49519 (N_49519,N_48799,N_48030);
nand U49520 (N_49520,N_48378,N_48253);
xnor U49521 (N_49521,N_48419,N_48663);
nand U49522 (N_49522,N_48419,N_48357);
xnor U49523 (N_49523,N_48596,N_48713);
and U49524 (N_49524,N_48689,N_48664);
and U49525 (N_49525,N_48772,N_48377);
nor U49526 (N_49526,N_48390,N_48086);
nand U49527 (N_49527,N_48539,N_48714);
xor U49528 (N_49528,N_48303,N_48444);
or U49529 (N_49529,N_48873,N_48913);
or U49530 (N_49530,N_48559,N_48388);
or U49531 (N_49531,N_48373,N_48169);
xnor U49532 (N_49532,N_48048,N_48751);
nor U49533 (N_49533,N_48808,N_48896);
nand U49534 (N_49534,N_48044,N_48442);
xor U49535 (N_49535,N_48514,N_48581);
xor U49536 (N_49536,N_48592,N_48599);
xor U49537 (N_49537,N_48045,N_48548);
nor U49538 (N_49538,N_48498,N_48137);
nand U49539 (N_49539,N_48958,N_48615);
nor U49540 (N_49540,N_48066,N_48573);
xor U49541 (N_49541,N_48039,N_48384);
xnor U49542 (N_49542,N_48127,N_48842);
nand U49543 (N_49543,N_48627,N_48603);
xnor U49544 (N_49544,N_48979,N_48208);
nand U49545 (N_49545,N_48536,N_48352);
or U49546 (N_49546,N_48471,N_48356);
nor U49547 (N_49547,N_48102,N_48696);
or U49548 (N_49548,N_48004,N_48077);
or U49549 (N_49549,N_48073,N_48803);
xnor U49550 (N_49550,N_48519,N_48036);
nand U49551 (N_49551,N_48747,N_48247);
xnor U49552 (N_49552,N_48845,N_48660);
nor U49553 (N_49553,N_48797,N_48118);
and U49554 (N_49554,N_48857,N_48333);
and U49555 (N_49555,N_48103,N_48159);
nand U49556 (N_49556,N_48317,N_48105);
xnor U49557 (N_49557,N_48542,N_48079);
nor U49558 (N_49558,N_48718,N_48952);
xor U49559 (N_49559,N_48112,N_48207);
nor U49560 (N_49560,N_48385,N_48015);
nand U49561 (N_49561,N_48986,N_48755);
xor U49562 (N_49562,N_48375,N_48110);
nor U49563 (N_49563,N_48519,N_48816);
nor U49564 (N_49564,N_48820,N_48974);
or U49565 (N_49565,N_48254,N_48450);
or U49566 (N_49566,N_48678,N_48160);
nand U49567 (N_49567,N_48188,N_48107);
xnor U49568 (N_49568,N_48402,N_48087);
or U49569 (N_49569,N_48347,N_48857);
nand U49570 (N_49570,N_48569,N_48938);
or U49571 (N_49571,N_48298,N_48018);
nor U49572 (N_49572,N_48236,N_48612);
nor U49573 (N_49573,N_48084,N_48817);
nand U49574 (N_49574,N_48937,N_48770);
xnor U49575 (N_49575,N_48655,N_48657);
or U49576 (N_49576,N_48426,N_48934);
xor U49577 (N_49577,N_48266,N_48184);
xor U49578 (N_49578,N_48166,N_48723);
xnor U49579 (N_49579,N_48078,N_48868);
nand U49580 (N_49580,N_48075,N_48934);
nand U49581 (N_49581,N_48265,N_48589);
nor U49582 (N_49582,N_48745,N_48376);
nand U49583 (N_49583,N_48046,N_48629);
nor U49584 (N_49584,N_48838,N_48393);
nor U49585 (N_49585,N_48962,N_48711);
xnor U49586 (N_49586,N_48186,N_48951);
xnor U49587 (N_49587,N_48453,N_48796);
nand U49588 (N_49588,N_48216,N_48771);
and U49589 (N_49589,N_48171,N_48689);
nand U49590 (N_49590,N_48869,N_48492);
or U49591 (N_49591,N_48809,N_48350);
nand U49592 (N_49592,N_48392,N_48421);
nor U49593 (N_49593,N_48412,N_48205);
and U49594 (N_49594,N_48568,N_48917);
xor U49595 (N_49595,N_48502,N_48655);
nor U49596 (N_49596,N_48805,N_48403);
or U49597 (N_49597,N_48943,N_48244);
xnor U49598 (N_49598,N_48167,N_48227);
and U49599 (N_49599,N_48470,N_48485);
nor U49600 (N_49600,N_48073,N_48723);
nand U49601 (N_49601,N_48758,N_48018);
nand U49602 (N_49602,N_48655,N_48005);
nor U49603 (N_49603,N_48001,N_48070);
nor U49604 (N_49604,N_48443,N_48935);
xor U49605 (N_49605,N_48879,N_48878);
and U49606 (N_49606,N_48713,N_48089);
nand U49607 (N_49607,N_48846,N_48735);
or U49608 (N_49608,N_48148,N_48592);
nor U49609 (N_49609,N_48084,N_48857);
nor U49610 (N_49610,N_48951,N_48607);
nand U49611 (N_49611,N_48351,N_48954);
or U49612 (N_49612,N_48886,N_48226);
nor U49613 (N_49613,N_48237,N_48927);
and U49614 (N_49614,N_48987,N_48739);
nor U49615 (N_49615,N_48293,N_48697);
nand U49616 (N_49616,N_48929,N_48455);
and U49617 (N_49617,N_48453,N_48230);
xnor U49618 (N_49618,N_48092,N_48539);
or U49619 (N_49619,N_48047,N_48613);
and U49620 (N_49620,N_48707,N_48509);
nor U49621 (N_49621,N_48541,N_48129);
nor U49622 (N_49622,N_48405,N_48394);
xnor U49623 (N_49623,N_48837,N_48409);
nor U49624 (N_49624,N_48455,N_48088);
nand U49625 (N_49625,N_48812,N_48481);
or U49626 (N_49626,N_48329,N_48027);
nand U49627 (N_49627,N_48462,N_48264);
nand U49628 (N_49628,N_48125,N_48363);
xor U49629 (N_49629,N_48748,N_48983);
nand U49630 (N_49630,N_48748,N_48407);
xor U49631 (N_49631,N_48923,N_48893);
nor U49632 (N_49632,N_48763,N_48137);
nand U49633 (N_49633,N_48333,N_48984);
nor U49634 (N_49634,N_48668,N_48980);
xor U49635 (N_49635,N_48991,N_48614);
nand U49636 (N_49636,N_48174,N_48375);
nor U49637 (N_49637,N_48976,N_48320);
or U49638 (N_49638,N_48933,N_48403);
xnor U49639 (N_49639,N_48102,N_48596);
nand U49640 (N_49640,N_48935,N_48782);
and U49641 (N_49641,N_48093,N_48670);
xor U49642 (N_49642,N_48115,N_48625);
or U49643 (N_49643,N_48549,N_48903);
nand U49644 (N_49644,N_48419,N_48287);
xnor U49645 (N_49645,N_48580,N_48484);
nand U49646 (N_49646,N_48657,N_48920);
nand U49647 (N_49647,N_48410,N_48657);
or U49648 (N_49648,N_48256,N_48615);
and U49649 (N_49649,N_48874,N_48622);
and U49650 (N_49650,N_48304,N_48195);
xor U49651 (N_49651,N_48551,N_48995);
or U49652 (N_49652,N_48153,N_48886);
or U49653 (N_49653,N_48426,N_48443);
or U49654 (N_49654,N_48355,N_48377);
nand U49655 (N_49655,N_48942,N_48802);
nor U49656 (N_49656,N_48669,N_48381);
or U49657 (N_49657,N_48557,N_48449);
xor U49658 (N_49658,N_48110,N_48699);
and U49659 (N_49659,N_48029,N_48066);
xnor U49660 (N_49660,N_48384,N_48863);
and U49661 (N_49661,N_48463,N_48145);
nand U49662 (N_49662,N_48623,N_48969);
or U49663 (N_49663,N_48717,N_48296);
xnor U49664 (N_49664,N_48685,N_48795);
nor U49665 (N_49665,N_48131,N_48877);
and U49666 (N_49666,N_48419,N_48116);
nand U49667 (N_49667,N_48047,N_48630);
xnor U49668 (N_49668,N_48378,N_48523);
nor U49669 (N_49669,N_48933,N_48694);
or U49670 (N_49670,N_48093,N_48246);
nand U49671 (N_49671,N_48265,N_48466);
nand U49672 (N_49672,N_48053,N_48869);
nor U49673 (N_49673,N_48178,N_48657);
nand U49674 (N_49674,N_48657,N_48945);
nand U49675 (N_49675,N_48108,N_48339);
xor U49676 (N_49676,N_48640,N_48860);
nor U49677 (N_49677,N_48903,N_48667);
nor U49678 (N_49678,N_48312,N_48324);
nor U49679 (N_49679,N_48330,N_48858);
or U49680 (N_49680,N_48725,N_48986);
and U49681 (N_49681,N_48202,N_48549);
and U49682 (N_49682,N_48794,N_48644);
xnor U49683 (N_49683,N_48894,N_48577);
xnor U49684 (N_49684,N_48016,N_48183);
and U49685 (N_49685,N_48975,N_48107);
nor U49686 (N_49686,N_48447,N_48045);
nand U49687 (N_49687,N_48236,N_48443);
or U49688 (N_49688,N_48265,N_48040);
nor U49689 (N_49689,N_48332,N_48195);
or U49690 (N_49690,N_48967,N_48740);
and U49691 (N_49691,N_48100,N_48968);
nor U49692 (N_49692,N_48694,N_48857);
or U49693 (N_49693,N_48439,N_48601);
and U49694 (N_49694,N_48179,N_48713);
and U49695 (N_49695,N_48070,N_48723);
nor U49696 (N_49696,N_48443,N_48471);
or U49697 (N_49697,N_48824,N_48605);
and U49698 (N_49698,N_48849,N_48259);
or U49699 (N_49699,N_48989,N_48011);
nand U49700 (N_49700,N_48185,N_48281);
and U49701 (N_49701,N_48544,N_48146);
nor U49702 (N_49702,N_48959,N_48909);
nor U49703 (N_49703,N_48581,N_48038);
or U49704 (N_49704,N_48881,N_48353);
nand U49705 (N_49705,N_48626,N_48439);
nand U49706 (N_49706,N_48292,N_48407);
nand U49707 (N_49707,N_48604,N_48834);
or U49708 (N_49708,N_48072,N_48206);
nor U49709 (N_49709,N_48097,N_48072);
nand U49710 (N_49710,N_48401,N_48124);
nand U49711 (N_49711,N_48888,N_48307);
nand U49712 (N_49712,N_48889,N_48182);
xor U49713 (N_49713,N_48077,N_48222);
nor U49714 (N_49714,N_48209,N_48848);
or U49715 (N_49715,N_48703,N_48129);
xor U49716 (N_49716,N_48177,N_48182);
and U49717 (N_49717,N_48518,N_48604);
nor U49718 (N_49718,N_48574,N_48610);
nor U49719 (N_49719,N_48522,N_48258);
and U49720 (N_49720,N_48646,N_48754);
and U49721 (N_49721,N_48321,N_48178);
xor U49722 (N_49722,N_48475,N_48307);
nand U49723 (N_49723,N_48259,N_48415);
nor U49724 (N_49724,N_48056,N_48125);
nand U49725 (N_49725,N_48667,N_48732);
nor U49726 (N_49726,N_48341,N_48213);
nand U49727 (N_49727,N_48068,N_48050);
or U49728 (N_49728,N_48118,N_48788);
nor U49729 (N_49729,N_48845,N_48083);
or U49730 (N_49730,N_48960,N_48440);
or U49731 (N_49731,N_48149,N_48898);
nand U49732 (N_49732,N_48349,N_48640);
or U49733 (N_49733,N_48764,N_48480);
or U49734 (N_49734,N_48374,N_48269);
or U49735 (N_49735,N_48840,N_48887);
nand U49736 (N_49736,N_48851,N_48141);
nand U49737 (N_49737,N_48096,N_48177);
xor U49738 (N_49738,N_48733,N_48021);
xnor U49739 (N_49739,N_48989,N_48963);
and U49740 (N_49740,N_48325,N_48648);
or U49741 (N_49741,N_48504,N_48886);
or U49742 (N_49742,N_48021,N_48901);
nor U49743 (N_49743,N_48603,N_48463);
nor U49744 (N_49744,N_48115,N_48804);
or U49745 (N_49745,N_48335,N_48550);
nand U49746 (N_49746,N_48810,N_48040);
and U49747 (N_49747,N_48670,N_48746);
xnor U49748 (N_49748,N_48438,N_48073);
or U49749 (N_49749,N_48540,N_48192);
or U49750 (N_49750,N_48021,N_48410);
nor U49751 (N_49751,N_48919,N_48580);
or U49752 (N_49752,N_48819,N_48436);
and U49753 (N_49753,N_48733,N_48589);
xnor U49754 (N_49754,N_48068,N_48759);
nor U49755 (N_49755,N_48825,N_48706);
and U49756 (N_49756,N_48833,N_48752);
nand U49757 (N_49757,N_48049,N_48964);
nor U49758 (N_49758,N_48083,N_48115);
nand U49759 (N_49759,N_48783,N_48567);
or U49760 (N_49760,N_48564,N_48198);
and U49761 (N_49761,N_48610,N_48436);
nand U49762 (N_49762,N_48890,N_48560);
xor U49763 (N_49763,N_48016,N_48013);
nand U49764 (N_49764,N_48728,N_48451);
nor U49765 (N_49765,N_48319,N_48131);
and U49766 (N_49766,N_48082,N_48674);
and U49767 (N_49767,N_48425,N_48768);
nand U49768 (N_49768,N_48589,N_48887);
and U49769 (N_49769,N_48319,N_48394);
nor U49770 (N_49770,N_48674,N_48837);
xnor U49771 (N_49771,N_48122,N_48879);
nor U49772 (N_49772,N_48140,N_48251);
nand U49773 (N_49773,N_48996,N_48906);
xor U49774 (N_49774,N_48468,N_48430);
xnor U49775 (N_49775,N_48814,N_48173);
nor U49776 (N_49776,N_48785,N_48796);
nor U49777 (N_49777,N_48096,N_48578);
nor U49778 (N_49778,N_48127,N_48823);
xor U49779 (N_49779,N_48325,N_48785);
or U49780 (N_49780,N_48137,N_48813);
nor U49781 (N_49781,N_48308,N_48543);
and U49782 (N_49782,N_48010,N_48112);
xor U49783 (N_49783,N_48097,N_48653);
xnor U49784 (N_49784,N_48910,N_48160);
and U49785 (N_49785,N_48034,N_48453);
or U49786 (N_49786,N_48012,N_48217);
xnor U49787 (N_49787,N_48134,N_48263);
or U49788 (N_49788,N_48390,N_48982);
or U49789 (N_49789,N_48677,N_48929);
or U49790 (N_49790,N_48114,N_48067);
and U49791 (N_49791,N_48947,N_48943);
xor U49792 (N_49792,N_48650,N_48601);
and U49793 (N_49793,N_48698,N_48330);
and U49794 (N_49794,N_48587,N_48714);
nand U49795 (N_49795,N_48559,N_48451);
or U49796 (N_49796,N_48700,N_48042);
and U49797 (N_49797,N_48706,N_48221);
or U49798 (N_49798,N_48352,N_48016);
xor U49799 (N_49799,N_48407,N_48345);
xor U49800 (N_49800,N_48112,N_48847);
nor U49801 (N_49801,N_48178,N_48606);
nand U49802 (N_49802,N_48215,N_48021);
nor U49803 (N_49803,N_48173,N_48282);
nor U49804 (N_49804,N_48306,N_48133);
xor U49805 (N_49805,N_48705,N_48468);
xor U49806 (N_49806,N_48528,N_48043);
nor U49807 (N_49807,N_48328,N_48162);
nor U49808 (N_49808,N_48727,N_48821);
or U49809 (N_49809,N_48503,N_48051);
nor U49810 (N_49810,N_48858,N_48470);
xnor U49811 (N_49811,N_48688,N_48861);
nor U49812 (N_49812,N_48701,N_48034);
nor U49813 (N_49813,N_48207,N_48130);
or U49814 (N_49814,N_48703,N_48550);
and U49815 (N_49815,N_48331,N_48991);
xnor U49816 (N_49816,N_48152,N_48193);
xnor U49817 (N_49817,N_48259,N_48670);
nand U49818 (N_49818,N_48774,N_48819);
xnor U49819 (N_49819,N_48304,N_48135);
xor U49820 (N_49820,N_48598,N_48246);
and U49821 (N_49821,N_48150,N_48882);
and U49822 (N_49822,N_48925,N_48776);
nor U49823 (N_49823,N_48948,N_48033);
nand U49824 (N_49824,N_48493,N_48258);
xnor U49825 (N_49825,N_48449,N_48053);
or U49826 (N_49826,N_48012,N_48660);
or U49827 (N_49827,N_48333,N_48618);
nand U49828 (N_49828,N_48171,N_48947);
xor U49829 (N_49829,N_48732,N_48118);
nand U49830 (N_49830,N_48807,N_48166);
or U49831 (N_49831,N_48655,N_48286);
and U49832 (N_49832,N_48781,N_48171);
and U49833 (N_49833,N_48462,N_48922);
or U49834 (N_49834,N_48969,N_48607);
and U49835 (N_49835,N_48101,N_48058);
xor U49836 (N_49836,N_48789,N_48532);
and U49837 (N_49837,N_48940,N_48127);
or U49838 (N_49838,N_48345,N_48421);
and U49839 (N_49839,N_48719,N_48119);
and U49840 (N_49840,N_48266,N_48596);
xor U49841 (N_49841,N_48215,N_48292);
or U49842 (N_49842,N_48126,N_48434);
or U49843 (N_49843,N_48863,N_48652);
nand U49844 (N_49844,N_48055,N_48975);
nand U49845 (N_49845,N_48604,N_48709);
nand U49846 (N_49846,N_48655,N_48630);
nand U49847 (N_49847,N_48115,N_48162);
nor U49848 (N_49848,N_48932,N_48881);
and U49849 (N_49849,N_48459,N_48615);
nor U49850 (N_49850,N_48178,N_48819);
and U49851 (N_49851,N_48507,N_48272);
xnor U49852 (N_49852,N_48920,N_48352);
xor U49853 (N_49853,N_48068,N_48341);
nand U49854 (N_49854,N_48235,N_48335);
and U49855 (N_49855,N_48636,N_48822);
nand U49856 (N_49856,N_48271,N_48405);
nor U49857 (N_49857,N_48124,N_48289);
nor U49858 (N_49858,N_48679,N_48224);
and U49859 (N_49859,N_48523,N_48764);
and U49860 (N_49860,N_48084,N_48870);
and U49861 (N_49861,N_48235,N_48168);
nand U49862 (N_49862,N_48597,N_48439);
or U49863 (N_49863,N_48216,N_48272);
nor U49864 (N_49864,N_48513,N_48079);
nor U49865 (N_49865,N_48091,N_48051);
nand U49866 (N_49866,N_48752,N_48572);
and U49867 (N_49867,N_48089,N_48956);
and U49868 (N_49868,N_48899,N_48184);
and U49869 (N_49869,N_48337,N_48496);
nand U49870 (N_49870,N_48925,N_48439);
or U49871 (N_49871,N_48032,N_48381);
xnor U49872 (N_49872,N_48066,N_48695);
nand U49873 (N_49873,N_48856,N_48316);
nor U49874 (N_49874,N_48835,N_48025);
nor U49875 (N_49875,N_48910,N_48550);
nor U49876 (N_49876,N_48989,N_48161);
and U49877 (N_49877,N_48242,N_48950);
and U49878 (N_49878,N_48277,N_48512);
nor U49879 (N_49879,N_48562,N_48670);
and U49880 (N_49880,N_48164,N_48207);
nand U49881 (N_49881,N_48311,N_48157);
or U49882 (N_49882,N_48156,N_48140);
and U49883 (N_49883,N_48072,N_48671);
and U49884 (N_49884,N_48528,N_48529);
nand U49885 (N_49885,N_48950,N_48866);
nor U49886 (N_49886,N_48014,N_48537);
or U49887 (N_49887,N_48108,N_48892);
or U49888 (N_49888,N_48574,N_48704);
nor U49889 (N_49889,N_48981,N_48947);
xor U49890 (N_49890,N_48377,N_48066);
nand U49891 (N_49891,N_48213,N_48804);
xnor U49892 (N_49892,N_48723,N_48233);
xnor U49893 (N_49893,N_48612,N_48454);
xor U49894 (N_49894,N_48195,N_48153);
xor U49895 (N_49895,N_48332,N_48811);
nor U49896 (N_49896,N_48331,N_48659);
nor U49897 (N_49897,N_48231,N_48386);
nor U49898 (N_49898,N_48268,N_48295);
or U49899 (N_49899,N_48822,N_48361);
and U49900 (N_49900,N_48376,N_48002);
and U49901 (N_49901,N_48475,N_48352);
or U49902 (N_49902,N_48193,N_48930);
xor U49903 (N_49903,N_48096,N_48055);
nand U49904 (N_49904,N_48201,N_48368);
nand U49905 (N_49905,N_48505,N_48496);
nor U49906 (N_49906,N_48750,N_48757);
xnor U49907 (N_49907,N_48628,N_48586);
nand U49908 (N_49908,N_48491,N_48767);
nor U49909 (N_49909,N_48759,N_48522);
xor U49910 (N_49910,N_48028,N_48690);
nand U49911 (N_49911,N_48923,N_48303);
xor U49912 (N_49912,N_48158,N_48532);
xor U49913 (N_49913,N_48856,N_48787);
and U49914 (N_49914,N_48924,N_48672);
nand U49915 (N_49915,N_48385,N_48709);
and U49916 (N_49916,N_48163,N_48765);
and U49917 (N_49917,N_48357,N_48387);
xor U49918 (N_49918,N_48937,N_48020);
nor U49919 (N_49919,N_48186,N_48654);
nor U49920 (N_49920,N_48339,N_48567);
xor U49921 (N_49921,N_48447,N_48480);
or U49922 (N_49922,N_48606,N_48786);
nor U49923 (N_49923,N_48886,N_48191);
or U49924 (N_49924,N_48538,N_48777);
or U49925 (N_49925,N_48032,N_48585);
and U49926 (N_49926,N_48789,N_48414);
xnor U49927 (N_49927,N_48760,N_48445);
nor U49928 (N_49928,N_48511,N_48256);
xor U49929 (N_49929,N_48034,N_48766);
or U49930 (N_49930,N_48746,N_48216);
and U49931 (N_49931,N_48961,N_48744);
and U49932 (N_49932,N_48786,N_48356);
nand U49933 (N_49933,N_48065,N_48297);
and U49934 (N_49934,N_48165,N_48388);
or U49935 (N_49935,N_48193,N_48765);
nor U49936 (N_49936,N_48773,N_48948);
nand U49937 (N_49937,N_48147,N_48258);
and U49938 (N_49938,N_48710,N_48217);
xnor U49939 (N_49939,N_48067,N_48143);
nor U49940 (N_49940,N_48449,N_48989);
nor U49941 (N_49941,N_48729,N_48915);
nor U49942 (N_49942,N_48087,N_48620);
or U49943 (N_49943,N_48364,N_48228);
nand U49944 (N_49944,N_48045,N_48702);
nand U49945 (N_49945,N_48425,N_48993);
xnor U49946 (N_49946,N_48951,N_48873);
nand U49947 (N_49947,N_48940,N_48297);
nor U49948 (N_49948,N_48399,N_48131);
nand U49949 (N_49949,N_48559,N_48747);
or U49950 (N_49950,N_48529,N_48171);
xnor U49951 (N_49951,N_48612,N_48122);
and U49952 (N_49952,N_48998,N_48941);
and U49953 (N_49953,N_48918,N_48002);
or U49954 (N_49954,N_48558,N_48948);
nor U49955 (N_49955,N_48398,N_48095);
xnor U49956 (N_49956,N_48322,N_48846);
xnor U49957 (N_49957,N_48611,N_48506);
and U49958 (N_49958,N_48386,N_48506);
nor U49959 (N_49959,N_48580,N_48118);
nand U49960 (N_49960,N_48587,N_48487);
nor U49961 (N_49961,N_48071,N_48826);
or U49962 (N_49962,N_48634,N_48189);
nand U49963 (N_49963,N_48951,N_48071);
nand U49964 (N_49964,N_48769,N_48589);
or U49965 (N_49965,N_48540,N_48891);
nand U49966 (N_49966,N_48178,N_48660);
or U49967 (N_49967,N_48217,N_48007);
and U49968 (N_49968,N_48549,N_48200);
or U49969 (N_49969,N_48154,N_48129);
nor U49970 (N_49970,N_48526,N_48719);
and U49971 (N_49971,N_48229,N_48312);
nand U49972 (N_49972,N_48924,N_48153);
xnor U49973 (N_49973,N_48186,N_48632);
xnor U49974 (N_49974,N_48346,N_48864);
nor U49975 (N_49975,N_48354,N_48028);
nand U49976 (N_49976,N_48283,N_48061);
or U49977 (N_49977,N_48528,N_48037);
or U49978 (N_49978,N_48343,N_48887);
or U49979 (N_49979,N_48536,N_48905);
and U49980 (N_49980,N_48464,N_48276);
and U49981 (N_49981,N_48698,N_48802);
xnor U49982 (N_49982,N_48411,N_48390);
xor U49983 (N_49983,N_48893,N_48683);
nand U49984 (N_49984,N_48736,N_48455);
and U49985 (N_49985,N_48486,N_48562);
and U49986 (N_49986,N_48569,N_48681);
xor U49987 (N_49987,N_48140,N_48410);
xor U49988 (N_49988,N_48416,N_48237);
nand U49989 (N_49989,N_48024,N_48197);
nor U49990 (N_49990,N_48695,N_48957);
nor U49991 (N_49991,N_48244,N_48507);
nor U49992 (N_49992,N_48592,N_48869);
or U49993 (N_49993,N_48877,N_48857);
and U49994 (N_49994,N_48595,N_48356);
nand U49995 (N_49995,N_48823,N_48856);
nor U49996 (N_49996,N_48275,N_48846);
xor U49997 (N_49997,N_48108,N_48578);
or U49998 (N_49998,N_48844,N_48499);
nor U49999 (N_49999,N_48877,N_48719);
nand UO_0 (O_0,N_49295,N_49221);
or UO_1 (O_1,N_49785,N_49126);
and UO_2 (O_2,N_49561,N_49335);
and UO_3 (O_3,N_49465,N_49754);
or UO_4 (O_4,N_49676,N_49764);
or UO_5 (O_5,N_49951,N_49058);
nor UO_6 (O_6,N_49244,N_49652);
nand UO_7 (O_7,N_49877,N_49899);
nand UO_8 (O_8,N_49635,N_49059);
nor UO_9 (O_9,N_49849,N_49495);
or UO_10 (O_10,N_49287,N_49095);
nand UO_11 (O_11,N_49001,N_49460);
or UO_12 (O_12,N_49422,N_49817);
nor UO_13 (O_13,N_49227,N_49511);
nand UO_14 (O_14,N_49284,N_49205);
xor UO_15 (O_15,N_49309,N_49722);
nand UO_16 (O_16,N_49346,N_49163);
or UO_17 (O_17,N_49254,N_49992);
nor UO_18 (O_18,N_49612,N_49779);
nor UO_19 (O_19,N_49609,N_49149);
or UO_20 (O_20,N_49861,N_49680);
nor UO_21 (O_21,N_49709,N_49049);
or UO_22 (O_22,N_49539,N_49397);
and UO_23 (O_23,N_49203,N_49316);
and UO_24 (O_24,N_49223,N_49050);
and UO_25 (O_25,N_49351,N_49989);
nor UO_26 (O_26,N_49554,N_49690);
nor UO_27 (O_27,N_49837,N_49536);
nor UO_28 (O_28,N_49915,N_49831);
xor UO_29 (O_29,N_49751,N_49454);
xnor UO_30 (O_30,N_49990,N_49256);
or UO_31 (O_31,N_49273,N_49655);
nor UO_32 (O_32,N_49175,N_49540);
nor UO_33 (O_33,N_49400,N_49304);
nor UO_34 (O_34,N_49482,N_49937);
and UO_35 (O_35,N_49427,N_49296);
and UO_36 (O_36,N_49542,N_49041);
and UO_37 (O_37,N_49546,N_49399);
nand UO_38 (O_38,N_49171,N_49130);
nor UO_39 (O_39,N_49199,N_49865);
nor UO_40 (O_40,N_49177,N_49017);
nand UO_41 (O_41,N_49696,N_49693);
or UO_42 (O_42,N_49802,N_49288);
xor UO_43 (O_43,N_49337,N_49329);
and UO_44 (O_44,N_49068,N_49241);
or UO_45 (O_45,N_49900,N_49201);
or UO_46 (O_46,N_49863,N_49154);
nor UO_47 (O_47,N_49891,N_49769);
nor UO_48 (O_48,N_49759,N_49851);
nand UO_49 (O_49,N_49219,N_49667);
xor UO_50 (O_50,N_49305,N_49846);
nor UO_51 (O_51,N_49767,N_49641);
xnor UO_52 (O_52,N_49470,N_49942);
or UO_53 (O_53,N_49557,N_49020);
nor UO_54 (O_54,N_49710,N_49172);
nand UO_55 (O_55,N_49982,N_49210);
xor UO_56 (O_56,N_49164,N_49114);
and UO_57 (O_57,N_49517,N_49286);
nand UO_58 (O_58,N_49645,N_49189);
xnor UO_59 (O_59,N_49396,N_49193);
xor UO_60 (O_60,N_49531,N_49463);
nor UO_61 (O_61,N_49515,N_49842);
and UO_62 (O_62,N_49883,N_49448);
nor UO_63 (O_63,N_49650,N_49372);
nand UO_64 (O_64,N_49505,N_49739);
or UO_65 (O_65,N_49753,N_49004);
nor UO_66 (O_66,N_49333,N_49191);
nor UO_67 (O_67,N_49721,N_49852);
nand UO_68 (O_68,N_49800,N_49875);
and UO_69 (O_69,N_49012,N_49995);
and UO_70 (O_70,N_49322,N_49508);
and UO_71 (O_71,N_49468,N_49647);
nor UO_72 (O_72,N_49027,N_49317);
nor UO_73 (O_73,N_49057,N_49594);
xnor UO_74 (O_74,N_49220,N_49222);
xnor UO_75 (O_75,N_49692,N_49549);
xor UO_76 (O_76,N_49474,N_49858);
or UO_77 (O_77,N_49748,N_49357);
and UO_78 (O_78,N_49161,N_49360);
xor UO_79 (O_79,N_49098,N_49872);
nand UO_80 (O_80,N_49662,N_49786);
nor UO_81 (O_81,N_49055,N_49890);
xor UO_82 (O_82,N_49046,N_49019);
xor UO_83 (O_83,N_49311,N_49781);
xnor UO_84 (O_84,N_49906,N_49209);
xor UO_85 (O_85,N_49487,N_49620);
or UO_86 (O_86,N_49701,N_49242);
and UO_87 (O_87,N_49051,N_49010);
xnor UO_88 (O_88,N_49815,N_49668);
or UO_89 (O_89,N_49099,N_49332);
and UO_90 (O_90,N_49484,N_49720);
and UO_91 (O_91,N_49887,N_49853);
and UO_92 (O_92,N_49375,N_49587);
or UO_93 (O_93,N_49509,N_49471);
xor UO_94 (O_94,N_49477,N_49718);
or UO_95 (O_95,N_49884,N_49566);
xor UO_96 (O_96,N_49898,N_49829);
xnor UO_97 (O_97,N_49871,N_49541);
and UO_98 (O_98,N_49121,N_49791);
nor UO_99 (O_99,N_49847,N_49708);
nor UO_100 (O_100,N_49874,N_49778);
nand UO_101 (O_101,N_49530,N_49499);
xor UO_102 (O_102,N_49606,N_49231);
nand UO_103 (O_103,N_49081,N_49741);
and UO_104 (O_104,N_49535,N_49386);
and UO_105 (O_105,N_49763,N_49651);
nor UO_106 (O_106,N_49383,N_49233);
or UO_107 (O_107,N_49799,N_49673);
xor UO_108 (O_108,N_49324,N_49715);
xnor UO_109 (O_109,N_49052,N_49678);
and UO_110 (O_110,N_49133,N_49925);
nand UO_111 (O_111,N_49331,N_49596);
nor UO_112 (O_112,N_49994,N_49101);
nor UO_113 (O_113,N_49270,N_49263);
nor UO_114 (O_114,N_49129,N_49731);
and UO_115 (O_115,N_49611,N_49644);
xor UO_116 (O_116,N_49502,N_49965);
xor UO_117 (O_117,N_49476,N_49525);
or UO_118 (O_118,N_49090,N_49239);
or UO_119 (O_119,N_49868,N_49117);
and UO_120 (O_120,N_49380,N_49355);
nor UO_121 (O_121,N_49870,N_49336);
nand UO_122 (O_122,N_49366,N_49921);
and UO_123 (O_123,N_49637,N_49134);
nor UO_124 (O_124,N_49638,N_49077);
nor UO_125 (O_125,N_49569,N_49005);
nand UO_126 (O_126,N_49736,N_49473);
xnor UO_127 (O_127,N_49600,N_49737);
nand UO_128 (O_128,N_49192,N_49354);
nand UO_129 (O_129,N_49727,N_49719);
and UO_130 (O_130,N_49479,N_49573);
and UO_131 (O_131,N_49553,N_49766);
and UO_132 (O_132,N_49728,N_49840);
xor UO_133 (O_133,N_49971,N_49584);
or UO_134 (O_134,N_49744,N_49094);
xor UO_135 (O_135,N_49803,N_49136);
nand UO_136 (O_136,N_49089,N_49809);
and UO_137 (O_137,N_49603,N_49774);
nor UO_138 (O_138,N_49480,N_49216);
nor UO_139 (O_139,N_49342,N_49810);
xnor UO_140 (O_140,N_49901,N_49570);
nand UO_141 (O_141,N_49626,N_49087);
nor UO_142 (O_142,N_49128,N_49376);
nand UO_143 (O_143,N_49949,N_49957);
nor UO_144 (O_144,N_49956,N_49602);
nor UO_145 (O_145,N_49862,N_49249);
or UO_146 (O_146,N_49691,N_49008);
or UO_147 (O_147,N_49827,N_49729);
nand UO_148 (O_148,N_49776,N_49389);
nand UO_149 (O_149,N_49880,N_49705);
or UO_150 (O_150,N_49026,N_49439);
or UO_151 (O_151,N_49518,N_49973);
and UO_152 (O_152,N_49500,N_49440);
nor UO_153 (O_153,N_49271,N_49923);
nand UO_154 (O_154,N_49688,N_49371);
nand UO_155 (O_155,N_49856,N_49895);
nand UO_156 (O_156,N_49469,N_49462);
or UO_157 (O_157,N_49202,N_49092);
nand UO_158 (O_158,N_49974,N_49628);
xnor UO_159 (O_159,N_49677,N_49653);
xnor UO_160 (O_160,N_49850,N_49631);
nor UO_161 (O_161,N_49293,N_49946);
nand UO_162 (O_162,N_49167,N_49031);
nand UO_163 (O_163,N_49416,N_49493);
nor UO_164 (O_164,N_49586,N_49006);
and UO_165 (O_165,N_49443,N_49037);
and UO_166 (O_166,N_49893,N_49624);
and UO_167 (O_167,N_49580,N_49327);
nand UO_168 (O_168,N_49124,N_49713);
nor UO_169 (O_169,N_49639,N_49401);
nand UO_170 (O_170,N_49621,N_49155);
xnor UO_171 (O_171,N_49208,N_49243);
and UO_172 (O_172,N_49168,N_49732);
nor UO_173 (O_173,N_49083,N_49836);
nand UO_174 (O_174,N_49913,N_49053);
or UO_175 (O_175,N_49986,N_49016);
nand UO_176 (O_176,N_49929,N_49707);
and UO_177 (O_177,N_49504,N_49262);
nand UO_178 (O_178,N_49523,N_49844);
nor UO_179 (O_179,N_49784,N_49738);
or UO_180 (O_180,N_49072,N_49105);
or UO_181 (O_181,N_49733,N_49402);
nand UO_182 (O_182,N_49137,N_49093);
nand UO_183 (O_183,N_49218,N_49537);
nand UO_184 (O_184,N_49816,N_49259);
and UO_185 (O_185,N_49240,N_49200);
xnor UO_186 (O_186,N_49833,N_49265);
and UO_187 (O_187,N_49977,N_49987);
or UO_188 (O_188,N_49217,N_49301);
or UO_189 (O_189,N_49984,N_49808);
or UO_190 (O_190,N_49697,N_49555);
nor UO_191 (O_191,N_49467,N_49552);
or UO_192 (O_192,N_49415,N_49466);
or UO_193 (O_193,N_49165,N_49023);
xor UO_194 (O_194,N_49792,N_49151);
or UO_195 (O_195,N_49176,N_49740);
xnor UO_196 (O_196,N_49771,N_49365);
nand UO_197 (O_197,N_49746,N_49654);
and UO_198 (O_198,N_49250,N_49486);
xor UO_199 (O_199,N_49993,N_49437);
nor UO_200 (O_200,N_49689,N_49078);
or UO_201 (O_201,N_49079,N_49014);
and UO_202 (O_202,N_49257,N_49576);
or UO_203 (O_203,N_49015,N_49830);
nor UO_204 (O_204,N_49166,N_49675);
and UO_205 (O_205,N_49773,N_49181);
and UO_206 (O_206,N_49060,N_49275);
nand UO_207 (O_207,N_49714,N_49512);
and UO_208 (O_208,N_49266,N_49581);
and UO_209 (O_209,N_49312,N_49418);
nand UO_210 (O_210,N_49866,N_49116);
xnor UO_211 (O_211,N_49700,N_49524);
nand UO_212 (O_212,N_49459,N_49935);
xnor UO_213 (O_213,N_49451,N_49048);
or UO_214 (O_214,N_49762,N_49356);
xnor UO_215 (O_215,N_49393,N_49567);
nand UO_216 (O_216,N_49247,N_49490);
xor UO_217 (O_217,N_49319,N_49104);
nor UO_218 (O_218,N_49648,N_49142);
nor UO_219 (O_219,N_49757,N_49796);
xor UO_220 (O_220,N_49981,N_49343);
xnor UO_221 (O_221,N_49395,N_49604);
nor UO_222 (O_222,N_49267,N_49869);
or UO_223 (O_223,N_49933,N_49909);
nand UO_224 (O_224,N_49002,N_49622);
and UO_225 (O_225,N_49966,N_49007);
xnor UO_226 (O_226,N_49283,N_49873);
or UO_227 (O_227,N_49962,N_49723);
xnor UO_228 (O_228,N_49601,N_49528);
or UO_229 (O_229,N_49444,N_49119);
and UO_230 (O_230,N_49634,N_49406);
or UO_231 (O_231,N_49889,N_49533);
xnor UO_232 (O_232,N_49350,N_49967);
nor UO_233 (O_233,N_49353,N_49794);
and UO_234 (O_234,N_49712,N_49497);
nand UO_235 (O_235,N_49627,N_49029);
xor UO_236 (O_236,N_49907,N_49507);
nor UO_237 (O_237,N_49063,N_49003);
and UO_238 (O_238,N_49384,N_49173);
xor UO_239 (O_239,N_49591,N_49922);
and UO_240 (O_240,N_49423,N_49941);
or UO_241 (O_241,N_49562,N_49228);
and UO_242 (O_242,N_49629,N_49464);
xnor UO_243 (O_243,N_49761,N_49588);
nand UO_244 (O_244,N_49436,N_49153);
and UO_245 (O_245,N_49103,N_49657);
nor UO_246 (O_246,N_49320,N_49408);
nor UO_247 (O_247,N_49742,N_49716);
nor UO_248 (O_248,N_49407,N_49954);
xor UO_249 (O_249,N_49107,N_49914);
or UO_250 (O_250,N_49377,N_49503);
xor UO_251 (O_251,N_49091,N_49752);
nor UO_252 (O_252,N_49750,N_49843);
nor UO_253 (O_253,N_49281,N_49881);
nand UO_254 (O_254,N_49717,N_49636);
xor UO_255 (O_255,N_49032,N_49532);
xor UO_256 (O_256,N_49340,N_49447);
or UO_257 (O_257,N_49894,N_49062);
or UO_258 (O_258,N_49760,N_49080);
or UO_259 (O_259,N_49857,N_49456);
nand UO_260 (O_260,N_49328,N_49972);
and UO_261 (O_261,N_49968,N_49413);
xor UO_262 (O_262,N_49663,N_49429);
nand UO_263 (O_263,N_49488,N_49226);
nand UO_264 (O_264,N_49940,N_49110);
nor UO_265 (O_265,N_49790,N_49959);
and UO_266 (O_266,N_49428,N_49806);
xnor UO_267 (O_267,N_49326,N_49123);
or UO_268 (O_268,N_49777,N_49449);
or UO_269 (O_269,N_49607,N_49264);
and UO_270 (O_270,N_49315,N_49882);
nand UO_271 (O_271,N_49349,N_49640);
or UO_272 (O_272,N_49585,N_49127);
or UO_273 (O_273,N_49088,N_49577);
nand UO_274 (O_274,N_49338,N_49358);
and UO_275 (O_275,N_49630,N_49255);
xnor UO_276 (O_276,N_49261,N_49302);
and UO_277 (O_277,N_49671,N_49282);
xor UO_278 (O_278,N_49845,N_49445);
xnor UO_279 (O_279,N_49985,N_49252);
xor UO_280 (O_280,N_49197,N_49952);
and UO_281 (O_281,N_49521,N_49102);
or UO_282 (O_282,N_49361,N_49684);
and UO_283 (O_283,N_49135,N_49698);
xnor UO_284 (O_284,N_49162,N_49224);
nor UO_285 (O_285,N_49410,N_49411);
or UO_286 (O_286,N_49185,N_49550);
nor UO_287 (O_287,N_49724,N_49735);
nand UO_288 (O_288,N_49426,N_49100);
and UO_289 (O_289,N_49156,N_49278);
xor UO_290 (O_290,N_49695,N_49614);
nor UO_291 (O_291,N_49623,N_49314);
nand UO_292 (O_292,N_49325,N_49294);
nand UO_293 (O_293,N_49298,N_49021);
nor UO_294 (O_294,N_49483,N_49927);
nand UO_295 (O_295,N_49417,N_49146);
and UO_296 (O_296,N_49211,N_49685);
xnor UO_297 (O_297,N_49076,N_49373);
xor UO_298 (O_298,N_49948,N_49681);
nand UO_299 (O_299,N_49308,N_49944);
nand UO_300 (O_300,N_49303,N_49825);
nand UO_301 (O_301,N_49330,N_49132);
xnor UO_302 (O_302,N_49187,N_49307);
and UO_303 (O_303,N_49054,N_49387);
or UO_304 (O_304,N_49248,N_49919);
and UO_305 (O_305,N_49788,N_49073);
and UO_306 (O_306,N_49818,N_49547);
or UO_307 (O_307,N_49280,N_49633);
or UO_308 (O_308,N_49323,N_49498);
xor UO_309 (O_309,N_49043,N_49649);
or UO_310 (O_310,N_49666,N_49074);
nand UO_311 (O_311,N_49207,N_49139);
or UO_312 (O_312,N_49924,N_49501);
nor UO_313 (O_313,N_49572,N_49616);
or UO_314 (O_314,N_49159,N_49359);
nor UO_315 (O_315,N_49034,N_49822);
nand UO_316 (O_316,N_49215,N_49598);
xor UO_317 (O_317,N_49183,N_49213);
nor UO_318 (O_318,N_49075,N_49352);
and UO_319 (O_319,N_49425,N_49421);
or UO_320 (O_320,N_49605,N_49938);
xor UO_321 (O_321,N_49999,N_49196);
or UO_322 (O_322,N_49782,N_49318);
or UO_323 (O_323,N_49832,N_49939);
or UO_324 (O_324,N_49613,N_49022);
or UO_325 (O_325,N_49238,N_49589);
nor UO_326 (O_326,N_49038,N_49169);
or UO_327 (O_327,N_49235,N_49147);
or UO_328 (O_328,N_49268,N_49279);
nor UO_329 (O_329,N_49122,N_49450);
and UO_330 (O_330,N_49225,N_49787);
nor UO_331 (O_331,N_49912,N_49615);
nor UO_332 (O_332,N_49699,N_49886);
xnor UO_333 (O_333,N_49475,N_49979);
xnor UO_334 (O_334,N_49180,N_49814);
xor UO_335 (O_335,N_49028,N_49198);
nand UO_336 (O_336,N_49378,N_49398);
or UO_337 (O_337,N_49859,N_49930);
nand UO_338 (O_338,N_49885,N_49527);
and UO_339 (O_339,N_49823,N_49775);
or UO_340 (O_340,N_49253,N_49683);
xnor UO_341 (O_341,N_49042,N_49140);
or UO_342 (O_342,N_49011,N_49903);
nor UO_343 (O_343,N_49260,N_49364);
and UO_344 (O_344,N_49839,N_49195);
nand UO_345 (O_345,N_49348,N_49807);
or UO_346 (O_346,N_49047,N_49583);
nand UO_347 (O_347,N_49506,N_49457);
and UO_348 (O_348,N_49452,N_49489);
and UO_349 (O_349,N_49370,N_49064);
nand UO_350 (O_350,N_49141,N_49947);
nor UO_351 (O_351,N_49686,N_49381);
nor UO_352 (O_352,N_49433,N_49341);
xor UO_353 (O_353,N_49496,N_49108);
and UO_354 (O_354,N_49412,N_49682);
or UO_355 (O_355,N_49747,N_49113);
xnor UO_356 (O_356,N_49519,N_49069);
nor UO_357 (O_357,N_49625,N_49902);
and UO_358 (O_358,N_49970,N_49820);
nor UO_359 (O_359,N_49190,N_49526);
xor UO_360 (O_360,N_49290,N_49595);
and UO_361 (O_361,N_49904,N_49963);
nor UO_362 (O_362,N_49755,N_49559);
or UO_363 (O_363,N_49409,N_49204);
and UO_364 (O_364,N_49855,N_49665);
or UO_365 (O_365,N_49556,N_49659);
xnor UO_366 (O_366,N_49976,N_49246);
and UO_367 (O_367,N_49975,N_49579);
or UO_368 (O_368,N_49367,N_49955);
xor UO_369 (O_369,N_49274,N_49749);
or UO_370 (O_370,N_49000,N_49656);
xor UO_371 (O_371,N_49194,N_49170);
nand UO_372 (O_372,N_49251,N_49131);
xor UO_373 (O_373,N_49908,N_49404);
xnor UO_374 (O_374,N_49642,N_49916);
nand UO_375 (O_375,N_49988,N_49953);
xnor UO_376 (O_376,N_49632,N_49578);
and UO_377 (O_377,N_49996,N_49661);
or UO_378 (O_378,N_49812,N_49430);
nand UO_379 (O_379,N_49258,N_49044);
nand UO_380 (O_380,N_49212,N_49795);
xnor UO_381 (O_381,N_49392,N_49910);
nor UO_382 (O_382,N_49148,N_49565);
nand UO_383 (O_383,N_49980,N_49545);
xor UO_384 (O_384,N_49670,N_49819);
xnor UO_385 (O_385,N_49961,N_49236);
nor UO_386 (O_386,N_49179,N_49096);
and UO_387 (O_387,N_49453,N_49382);
and UO_388 (O_388,N_49813,N_49431);
nand UO_389 (O_389,N_49998,N_49514);
nor UO_390 (O_390,N_49013,N_49983);
or UO_391 (O_391,N_49801,N_49403);
nand UO_392 (O_392,N_49560,N_49593);
nor UO_393 (O_393,N_49936,N_49568);
or UO_394 (O_394,N_49276,N_49854);
xnor UO_395 (O_395,N_49897,N_49481);
and UO_396 (O_396,N_49888,N_49610);
nand UO_397 (O_397,N_49285,N_49574);
nor UO_398 (O_398,N_49793,N_49056);
and UO_399 (O_399,N_49405,N_49188);
xnor UO_400 (O_400,N_49563,N_49478);
nor UO_401 (O_401,N_49943,N_49841);
xnor UO_402 (O_402,N_49300,N_49391);
or UO_403 (O_403,N_49687,N_49472);
and UO_404 (O_404,N_49878,N_49726);
nor UO_405 (O_405,N_49932,N_49066);
nand UO_406 (O_406,N_49144,N_49379);
or UO_407 (O_407,N_49118,N_49798);
or UO_408 (O_408,N_49510,N_49571);
xnor UO_409 (O_409,N_49125,N_49374);
and UO_410 (O_410,N_49071,N_49269);
nand UO_411 (O_411,N_49905,N_49544);
nor UO_412 (O_412,N_49033,N_49917);
xor UO_413 (O_413,N_49797,N_49234);
and UO_414 (O_414,N_49230,N_49237);
or UO_415 (O_415,N_49551,N_49679);
nor UO_416 (O_416,N_49964,N_49706);
xnor UO_417 (O_417,N_49592,N_49458);
nor UO_418 (O_418,N_49834,N_49978);
nand UO_419 (O_419,N_49920,N_49082);
and UO_420 (O_420,N_49674,N_49485);
or UO_421 (O_421,N_49804,N_49896);
xor UO_422 (O_422,N_49520,N_49385);
or UO_423 (O_423,N_49711,N_49321);
nor UO_424 (O_424,N_49120,N_49435);
xnor UO_425 (O_425,N_49522,N_49867);
nor UO_426 (O_426,N_49768,N_49918);
or UO_427 (O_427,N_49772,N_49424);
xor UO_428 (O_428,N_49950,N_49035);
nand UO_429 (O_429,N_49145,N_49826);
xor UO_430 (O_430,N_49743,N_49297);
xnor UO_431 (O_431,N_49643,N_49025);
xor UO_432 (O_432,N_49660,N_49931);
and UO_433 (O_433,N_49420,N_49835);
and UO_434 (O_434,N_49926,N_49494);
or UO_435 (O_435,N_49065,N_49097);
or UO_436 (O_436,N_49824,N_49368);
and UO_437 (O_437,N_49548,N_49725);
nor UO_438 (O_438,N_49617,N_49045);
or UO_439 (O_439,N_49811,N_49529);
and UO_440 (O_440,N_49214,N_49441);
nand UO_441 (O_441,N_49455,N_49960);
or UO_442 (O_442,N_49702,N_49369);
or UO_443 (O_443,N_49182,N_49582);
or UO_444 (O_444,N_49160,N_49911);
xnor UO_445 (O_445,N_49783,N_49313);
xnor UO_446 (O_446,N_49860,N_49277);
and UO_447 (O_447,N_49438,N_49143);
nand UO_448 (O_448,N_49184,N_49291);
nor UO_449 (O_449,N_49491,N_49229);
nand UO_450 (O_450,N_49086,N_49150);
and UO_451 (O_451,N_49516,N_49765);
xor UO_452 (O_452,N_49513,N_49009);
or UO_453 (O_453,N_49534,N_49590);
xor UO_454 (O_454,N_49958,N_49805);
or UO_455 (O_455,N_49672,N_49111);
nand UO_456 (O_456,N_49599,N_49344);
and UO_457 (O_457,N_49363,N_49543);
xor UO_458 (O_458,N_49669,N_49292);
and UO_459 (O_459,N_49564,N_49703);
or UO_460 (O_460,N_49558,N_49024);
or UO_461 (O_461,N_49339,N_49152);
or UO_462 (O_462,N_49997,N_49934);
or UO_463 (O_463,N_49848,N_49394);
nor UO_464 (O_464,N_49206,N_49362);
xor UO_465 (O_465,N_49084,N_49538);
nor UO_466 (O_466,N_49174,N_49969);
and UO_467 (O_467,N_49419,N_49345);
xnor UO_468 (O_468,N_49414,N_49040);
nor UO_469 (O_469,N_49070,N_49347);
xor UO_470 (O_470,N_49299,N_49704);
xnor UO_471 (O_471,N_49758,N_49945);
xnor UO_472 (O_472,N_49730,N_49838);
nand UO_473 (O_473,N_49608,N_49664);
nor UO_474 (O_474,N_49694,N_49789);
nand UO_475 (O_475,N_49864,N_49432);
or UO_476 (O_476,N_49442,N_49390);
nor UO_477 (O_477,N_49178,N_49388);
nand UO_478 (O_478,N_49106,N_49756);
or UO_479 (O_479,N_49067,N_49245);
and UO_480 (O_480,N_49446,N_49289);
and UO_481 (O_481,N_49828,N_49306);
and UO_482 (O_482,N_49158,N_49039);
or UO_483 (O_483,N_49821,N_49138);
nand UO_484 (O_484,N_49310,N_49109);
and UO_485 (O_485,N_49492,N_49115);
nor UO_486 (O_486,N_49434,N_49061);
and UO_487 (O_487,N_49112,N_49157);
xor UO_488 (O_488,N_49619,N_49232);
or UO_489 (O_489,N_49892,N_49770);
and UO_490 (O_490,N_49618,N_49272);
xnor UO_491 (O_491,N_49186,N_49018);
xnor UO_492 (O_492,N_49334,N_49575);
nand UO_493 (O_493,N_49734,N_49461);
nand UO_494 (O_494,N_49780,N_49745);
or UO_495 (O_495,N_49085,N_49030);
nor UO_496 (O_496,N_49036,N_49597);
xor UO_497 (O_497,N_49646,N_49928);
xor UO_498 (O_498,N_49658,N_49991);
xnor UO_499 (O_499,N_49876,N_49879);
xor UO_500 (O_500,N_49535,N_49572);
nor UO_501 (O_501,N_49514,N_49903);
nor UO_502 (O_502,N_49594,N_49490);
nor UO_503 (O_503,N_49652,N_49804);
or UO_504 (O_504,N_49653,N_49934);
xor UO_505 (O_505,N_49853,N_49572);
and UO_506 (O_506,N_49269,N_49754);
or UO_507 (O_507,N_49075,N_49128);
nand UO_508 (O_508,N_49885,N_49595);
or UO_509 (O_509,N_49614,N_49952);
nor UO_510 (O_510,N_49108,N_49615);
and UO_511 (O_511,N_49272,N_49975);
nand UO_512 (O_512,N_49592,N_49208);
nand UO_513 (O_513,N_49076,N_49217);
nand UO_514 (O_514,N_49531,N_49422);
xor UO_515 (O_515,N_49002,N_49385);
nor UO_516 (O_516,N_49269,N_49640);
nor UO_517 (O_517,N_49163,N_49600);
nand UO_518 (O_518,N_49129,N_49988);
or UO_519 (O_519,N_49418,N_49172);
nor UO_520 (O_520,N_49424,N_49762);
xnor UO_521 (O_521,N_49036,N_49374);
xnor UO_522 (O_522,N_49913,N_49879);
and UO_523 (O_523,N_49241,N_49339);
xor UO_524 (O_524,N_49419,N_49992);
xnor UO_525 (O_525,N_49241,N_49569);
and UO_526 (O_526,N_49463,N_49523);
or UO_527 (O_527,N_49598,N_49517);
or UO_528 (O_528,N_49312,N_49592);
and UO_529 (O_529,N_49934,N_49005);
nand UO_530 (O_530,N_49178,N_49092);
xor UO_531 (O_531,N_49900,N_49606);
xor UO_532 (O_532,N_49456,N_49600);
xnor UO_533 (O_533,N_49434,N_49264);
nand UO_534 (O_534,N_49219,N_49619);
and UO_535 (O_535,N_49478,N_49718);
and UO_536 (O_536,N_49067,N_49529);
nor UO_537 (O_537,N_49817,N_49921);
xor UO_538 (O_538,N_49719,N_49193);
or UO_539 (O_539,N_49015,N_49560);
or UO_540 (O_540,N_49615,N_49126);
nand UO_541 (O_541,N_49693,N_49048);
nand UO_542 (O_542,N_49824,N_49095);
and UO_543 (O_543,N_49419,N_49725);
and UO_544 (O_544,N_49881,N_49417);
xnor UO_545 (O_545,N_49458,N_49148);
and UO_546 (O_546,N_49381,N_49560);
nor UO_547 (O_547,N_49503,N_49337);
nor UO_548 (O_548,N_49538,N_49729);
or UO_549 (O_549,N_49614,N_49262);
nand UO_550 (O_550,N_49356,N_49559);
nand UO_551 (O_551,N_49040,N_49839);
nor UO_552 (O_552,N_49170,N_49927);
and UO_553 (O_553,N_49251,N_49581);
and UO_554 (O_554,N_49463,N_49125);
nand UO_555 (O_555,N_49856,N_49353);
xor UO_556 (O_556,N_49199,N_49787);
or UO_557 (O_557,N_49000,N_49651);
or UO_558 (O_558,N_49420,N_49313);
nor UO_559 (O_559,N_49420,N_49999);
xnor UO_560 (O_560,N_49973,N_49477);
nor UO_561 (O_561,N_49577,N_49424);
xnor UO_562 (O_562,N_49739,N_49007);
nand UO_563 (O_563,N_49218,N_49005);
and UO_564 (O_564,N_49210,N_49944);
nand UO_565 (O_565,N_49526,N_49445);
and UO_566 (O_566,N_49435,N_49740);
or UO_567 (O_567,N_49252,N_49535);
nand UO_568 (O_568,N_49624,N_49139);
or UO_569 (O_569,N_49095,N_49745);
nand UO_570 (O_570,N_49667,N_49723);
nor UO_571 (O_571,N_49304,N_49138);
and UO_572 (O_572,N_49842,N_49044);
nand UO_573 (O_573,N_49859,N_49717);
nor UO_574 (O_574,N_49412,N_49386);
or UO_575 (O_575,N_49076,N_49990);
nor UO_576 (O_576,N_49418,N_49897);
xnor UO_577 (O_577,N_49376,N_49309);
or UO_578 (O_578,N_49161,N_49392);
or UO_579 (O_579,N_49299,N_49982);
and UO_580 (O_580,N_49989,N_49682);
and UO_581 (O_581,N_49610,N_49185);
or UO_582 (O_582,N_49306,N_49870);
and UO_583 (O_583,N_49598,N_49390);
or UO_584 (O_584,N_49285,N_49294);
nand UO_585 (O_585,N_49650,N_49529);
or UO_586 (O_586,N_49959,N_49958);
nand UO_587 (O_587,N_49901,N_49274);
or UO_588 (O_588,N_49306,N_49737);
xnor UO_589 (O_589,N_49713,N_49423);
or UO_590 (O_590,N_49748,N_49207);
xnor UO_591 (O_591,N_49163,N_49644);
nor UO_592 (O_592,N_49762,N_49314);
xor UO_593 (O_593,N_49269,N_49769);
and UO_594 (O_594,N_49723,N_49563);
and UO_595 (O_595,N_49464,N_49440);
nor UO_596 (O_596,N_49127,N_49990);
or UO_597 (O_597,N_49002,N_49470);
nor UO_598 (O_598,N_49436,N_49126);
and UO_599 (O_599,N_49153,N_49128);
and UO_600 (O_600,N_49653,N_49279);
nand UO_601 (O_601,N_49797,N_49029);
xnor UO_602 (O_602,N_49114,N_49821);
xor UO_603 (O_603,N_49948,N_49779);
nand UO_604 (O_604,N_49548,N_49565);
xor UO_605 (O_605,N_49301,N_49535);
nor UO_606 (O_606,N_49590,N_49692);
xnor UO_607 (O_607,N_49043,N_49479);
nand UO_608 (O_608,N_49403,N_49487);
nor UO_609 (O_609,N_49536,N_49416);
xor UO_610 (O_610,N_49694,N_49404);
and UO_611 (O_611,N_49732,N_49468);
nand UO_612 (O_612,N_49651,N_49696);
or UO_613 (O_613,N_49878,N_49151);
nor UO_614 (O_614,N_49895,N_49111);
and UO_615 (O_615,N_49426,N_49847);
or UO_616 (O_616,N_49088,N_49016);
xor UO_617 (O_617,N_49228,N_49568);
or UO_618 (O_618,N_49987,N_49611);
nor UO_619 (O_619,N_49954,N_49846);
nor UO_620 (O_620,N_49407,N_49453);
nand UO_621 (O_621,N_49442,N_49304);
or UO_622 (O_622,N_49784,N_49687);
and UO_623 (O_623,N_49067,N_49781);
nand UO_624 (O_624,N_49621,N_49669);
and UO_625 (O_625,N_49652,N_49198);
nand UO_626 (O_626,N_49134,N_49084);
and UO_627 (O_627,N_49304,N_49807);
and UO_628 (O_628,N_49841,N_49604);
xnor UO_629 (O_629,N_49352,N_49248);
or UO_630 (O_630,N_49568,N_49756);
xnor UO_631 (O_631,N_49657,N_49971);
nand UO_632 (O_632,N_49963,N_49605);
nor UO_633 (O_633,N_49445,N_49063);
or UO_634 (O_634,N_49312,N_49987);
xor UO_635 (O_635,N_49737,N_49461);
xor UO_636 (O_636,N_49168,N_49476);
nand UO_637 (O_637,N_49595,N_49831);
xor UO_638 (O_638,N_49200,N_49226);
or UO_639 (O_639,N_49465,N_49619);
nor UO_640 (O_640,N_49617,N_49226);
nor UO_641 (O_641,N_49850,N_49306);
and UO_642 (O_642,N_49784,N_49201);
and UO_643 (O_643,N_49338,N_49914);
and UO_644 (O_644,N_49475,N_49418);
nand UO_645 (O_645,N_49927,N_49459);
nand UO_646 (O_646,N_49918,N_49840);
nor UO_647 (O_647,N_49053,N_49203);
and UO_648 (O_648,N_49203,N_49716);
and UO_649 (O_649,N_49962,N_49084);
xor UO_650 (O_650,N_49479,N_49181);
nand UO_651 (O_651,N_49517,N_49181);
and UO_652 (O_652,N_49926,N_49727);
xor UO_653 (O_653,N_49444,N_49421);
xnor UO_654 (O_654,N_49676,N_49813);
or UO_655 (O_655,N_49806,N_49395);
and UO_656 (O_656,N_49840,N_49299);
or UO_657 (O_657,N_49800,N_49503);
or UO_658 (O_658,N_49598,N_49197);
nor UO_659 (O_659,N_49896,N_49206);
or UO_660 (O_660,N_49964,N_49510);
and UO_661 (O_661,N_49316,N_49584);
and UO_662 (O_662,N_49737,N_49597);
nand UO_663 (O_663,N_49233,N_49002);
nand UO_664 (O_664,N_49020,N_49682);
or UO_665 (O_665,N_49320,N_49615);
or UO_666 (O_666,N_49898,N_49691);
nor UO_667 (O_667,N_49978,N_49946);
xor UO_668 (O_668,N_49860,N_49013);
or UO_669 (O_669,N_49863,N_49573);
nor UO_670 (O_670,N_49857,N_49370);
xor UO_671 (O_671,N_49699,N_49125);
nor UO_672 (O_672,N_49528,N_49940);
nand UO_673 (O_673,N_49125,N_49467);
xor UO_674 (O_674,N_49549,N_49678);
xnor UO_675 (O_675,N_49384,N_49504);
xnor UO_676 (O_676,N_49079,N_49882);
nand UO_677 (O_677,N_49667,N_49368);
and UO_678 (O_678,N_49520,N_49756);
nor UO_679 (O_679,N_49554,N_49662);
nor UO_680 (O_680,N_49941,N_49961);
nor UO_681 (O_681,N_49183,N_49033);
and UO_682 (O_682,N_49867,N_49400);
or UO_683 (O_683,N_49741,N_49181);
and UO_684 (O_684,N_49227,N_49526);
xnor UO_685 (O_685,N_49872,N_49187);
nand UO_686 (O_686,N_49451,N_49365);
or UO_687 (O_687,N_49765,N_49480);
nor UO_688 (O_688,N_49702,N_49890);
and UO_689 (O_689,N_49490,N_49134);
xnor UO_690 (O_690,N_49616,N_49571);
or UO_691 (O_691,N_49574,N_49942);
xor UO_692 (O_692,N_49085,N_49562);
and UO_693 (O_693,N_49792,N_49208);
xnor UO_694 (O_694,N_49132,N_49967);
nor UO_695 (O_695,N_49705,N_49175);
nor UO_696 (O_696,N_49490,N_49460);
xnor UO_697 (O_697,N_49796,N_49808);
nand UO_698 (O_698,N_49293,N_49629);
nor UO_699 (O_699,N_49589,N_49290);
or UO_700 (O_700,N_49097,N_49746);
or UO_701 (O_701,N_49511,N_49650);
nand UO_702 (O_702,N_49993,N_49421);
nor UO_703 (O_703,N_49466,N_49960);
nand UO_704 (O_704,N_49427,N_49885);
and UO_705 (O_705,N_49587,N_49648);
xnor UO_706 (O_706,N_49357,N_49687);
nor UO_707 (O_707,N_49870,N_49615);
or UO_708 (O_708,N_49880,N_49812);
and UO_709 (O_709,N_49291,N_49981);
nand UO_710 (O_710,N_49730,N_49429);
nor UO_711 (O_711,N_49269,N_49321);
nand UO_712 (O_712,N_49488,N_49640);
or UO_713 (O_713,N_49909,N_49231);
nor UO_714 (O_714,N_49335,N_49216);
and UO_715 (O_715,N_49611,N_49009);
nand UO_716 (O_716,N_49407,N_49034);
nand UO_717 (O_717,N_49621,N_49507);
and UO_718 (O_718,N_49445,N_49939);
nand UO_719 (O_719,N_49497,N_49891);
nand UO_720 (O_720,N_49141,N_49522);
or UO_721 (O_721,N_49363,N_49472);
nor UO_722 (O_722,N_49750,N_49598);
nor UO_723 (O_723,N_49673,N_49719);
or UO_724 (O_724,N_49478,N_49206);
xor UO_725 (O_725,N_49341,N_49053);
xnor UO_726 (O_726,N_49159,N_49054);
or UO_727 (O_727,N_49292,N_49684);
or UO_728 (O_728,N_49035,N_49271);
xor UO_729 (O_729,N_49197,N_49692);
or UO_730 (O_730,N_49025,N_49024);
nor UO_731 (O_731,N_49968,N_49999);
xnor UO_732 (O_732,N_49596,N_49366);
xnor UO_733 (O_733,N_49339,N_49380);
nor UO_734 (O_734,N_49362,N_49338);
or UO_735 (O_735,N_49055,N_49879);
xor UO_736 (O_736,N_49946,N_49405);
nor UO_737 (O_737,N_49086,N_49782);
or UO_738 (O_738,N_49604,N_49903);
or UO_739 (O_739,N_49666,N_49174);
xor UO_740 (O_740,N_49868,N_49810);
or UO_741 (O_741,N_49042,N_49155);
xnor UO_742 (O_742,N_49518,N_49054);
xnor UO_743 (O_743,N_49356,N_49925);
xor UO_744 (O_744,N_49098,N_49707);
and UO_745 (O_745,N_49199,N_49198);
nor UO_746 (O_746,N_49747,N_49979);
xnor UO_747 (O_747,N_49892,N_49832);
and UO_748 (O_748,N_49923,N_49645);
xor UO_749 (O_749,N_49731,N_49231);
xnor UO_750 (O_750,N_49170,N_49142);
xor UO_751 (O_751,N_49632,N_49569);
and UO_752 (O_752,N_49951,N_49075);
nor UO_753 (O_753,N_49578,N_49453);
xor UO_754 (O_754,N_49186,N_49372);
nor UO_755 (O_755,N_49632,N_49606);
nor UO_756 (O_756,N_49871,N_49132);
or UO_757 (O_757,N_49646,N_49505);
nand UO_758 (O_758,N_49036,N_49521);
nand UO_759 (O_759,N_49975,N_49532);
or UO_760 (O_760,N_49100,N_49538);
or UO_761 (O_761,N_49754,N_49010);
xnor UO_762 (O_762,N_49864,N_49481);
and UO_763 (O_763,N_49666,N_49125);
or UO_764 (O_764,N_49110,N_49109);
and UO_765 (O_765,N_49565,N_49292);
and UO_766 (O_766,N_49883,N_49754);
nand UO_767 (O_767,N_49990,N_49653);
and UO_768 (O_768,N_49780,N_49271);
and UO_769 (O_769,N_49349,N_49543);
nand UO_770 (O_770,N_49846,N_49790);
xor UO_771 (O_771,N_49596,N_49350);
nand UO_772 (O_772,N_49731,N_49978);
xnor UO_773 (O_773,N_49895,N_49041);
and UO_774 (O_774,N_49440,N_49025);
nand UO_775 (O_775,N_49257,N_49461);
nor UO_776 (O_776,N_49647,N_49757);
or UO_777 (O_777,N_49131,N_49663);
xor UO_778 (O_778,N_49091,N_49351);
nand UO_779 (O_779,N_49577,N_49260);
or UO_780 (O_780,N_49146,N_49560);
or UO_781 (O_781,N_49597,N_49714);
and UO_782 (O_782,N_49836,N_49198);
xnor UO_783 (O_783,N_49455,N_49081);
xnor UO_784 (O_784,N_49861,N_49312);
or UO_785 (O_785,N_49558,N_49712);
and UO_786 (O_786,N_49962,N_49406);
nand UO_787 (O_787,N_49617,N_49293);
and UO_788 (O_788,N_49229,N_49869);
or UO_789 (O_789,N_49467,N_49566);
xnor UO_790 (O_790,N_49507,N_49143);
and UO_791 (O_791,N_49730,N_49892);
nand UO_792 (O_792,N_49514,N_49437);
nand UO_793 (O_793,N_49754,N_49257);
or UO_794 (O_794,N_49796,N_49919);
xor UO_795 (O_795,N_49175,N_49682);
xor UO_796 (O_796,N_49547,N_49678);
nand UO_797 (O_797,N_49431,N_49121);
and UO_798 (O_798,N_49440,N_49240);
and UO_799 (O_799,N_49266,N_49782);
xnor UO_800 (O_800,N_49322,N_49223);
and UO_801 (O_801,N_49564,N_49108);
or UO_802 (O_802,N_49615,N_49929);
nand UO_803 (O_803,N_49280,N_49329);
and UO_804 (O_804,N_49143,N_49040);
or UO_805 (O_805,N_49527,N_49751);
or UO_806 (O_806,N_49528,N_49560);
xnor UO_807 (O_807,N_49813,N_49320);
or UO_808 (O_808,N_49981,N_49887);
xor UO_809 (O_809,N_49657,N_49634);
nor UO_810 (O_810,N_49665,N_49127);
nor UO_811 (O_811,N_49532,N_49669);
nand UO_812 (O_812,N_49436,N_49650);
nor UO_813 (O_813,N_49256,N_49763);
xnor UO_814 (O_814,N_49139,N_49323);
or UO_815 (O_815,N_49279,N_49206);
xnor UO_816 (O_816,N_49018,N_49468);
nor UO_817 (O_817,N_49907,N_49611);
xnor UO_818 (O_818,N_49770,N_49881);
nand UO_819 (O_819,N_49598,N_49825);
nor UO_820 (O_820,N_49566,N_49956);
xor UO_821 (O_821,N_49156,N_49713);
nor UO_822 (O_822,N_49096,N_49370);
nor UO_823 (O_823,N_49365,N_49251);
nand UO_824 (O_824,N_49995,N_49959);
and UO_825 (O_825,N_49691,N_49050);
nand UO_826 (O_826,N_49907,N_49131);
xnor UO_827 (O_827,N_49160,N_49398);
xnor UO_828 (O_828,N_49775,N_49424);
nor UO_829 (O_829,N_49387,N_49526);
nor UO_830 (O_830,N_49750,N_49881);
nor UO_831 (O_831,N_49105,N_49843);
and UO_832 (O_832,N_49790,N_49613);
xnor UO_833 (O_833,N_49492,N_49505);
or UO_834 (O_834,N_49970,N_49585);
and UO_835 (O_835,N_49078,N_49008);
and UO_836 (O_836,N_49099,N_49671);
nor UO_837 (O_837,N_49426,N_49892);
or UO_838 (O_838,N_49657,N_49085);
nor UO_839 (O_839,N_49190,N_49199);
xnor UO_840 (O_840,N_49540,N_49437);
or UO_841 (O_841,N_49366,N_49906);
xor UO_842 (O_842,N_49948,N_49639);
nor UO_843 (O_843,N_49281,N_49237);
nand UO_844 (O_844,N_49717,N_49333);
and UO_845 (O_845,N_49870,N_49320);
nand UO_846 (O_846,N_49561,N_49140);
nor UO_847 (O_847,N_49117,N_49102);
nor UO_848 (O_848,N_49127,N_49743);
and UO_849 (O_849,N_49842,N_49797);
nand UO_850 (O_850,N_49110,N_49480);
nand UO_851 (O_851,N_49954,N_49900);
or UO_852 (O_852,N_49991,N_49571);
and UO_853 (O_853,N_49056,N_49784);
nand UO_854 (O_854,N_49386,N_49824);
nand UO_855 (O_855,N_49731,N_49995);
xor UO_856 (O_856,N_49528,N_49733);
xor UO_857 (O_857,N_49938,N_49845);
or UO_858 (O_858,N_49279,N_49613);
and UO_859 (O_859,N_49269,N_49648);
nand UO_860 (O_860,N_49217,N_49925);
xnor UO_861 (O_861,N_49184,N_49949);
or UO_862 (O_862,N_49576,N_49939);
nor UO_863 (O_863,N_49513,N_49122);
or UO_864 (O_864,N_49134,N_49557);
nor UO_865 (O_865,N_49082,N_49437);
nand UO_866 (O_866,N_49548,N_49984);
xnor UO_867 (O_867,N_49663,N_49422);
nor UO_868 (O_868,N_49049,N_49857);
xor UO_869 (O_869,N_49572,N_49529);
xor UO_870 (O_870,N_49896,N_49462);
nand UO_871 (O_871,N_49732,N_49065);
or UO_872 (O_872,N_49261,N_49112);
nor UO_873 (O_873,N_49448,N_49313);
or UO_874 (O_874,N_49304,N_49572);
or UO_875 (O_875,N_49534,N_49020);
nor UO_876 (O_876,N_49089,N_49259);
and UO_877 (O_877,N_49935,N_49538);
nor UO_878 (O_878,N_49903,N_49467);
xnor UO_879 (O_879,N_49556,N_49078);
xnor UO_880 (O_880,N_49777,N_49547);
nand UO_881 (O_881,N_49278,N_49502);
nand UO_882 (O_882,N_49030,N_49257);
nand UO_883 (O_883,N_49241,N_49810);
xnor UO_884 (O_884,N_49599,N_49736);
nand UO_885 (O_885,N_49971,N_49160);
nor UO_886 (O_886,N_49221,N_49584);
or UO_887 (O_887,N_49452,N_49108);
xor UO_888 (O_888,N_49608,N_49115);
nor UO_889 (O_889,N_49908,N_49316);
nand UO_890 (O_890,N_49308,N_49900);
xor UO_891 (O_891,N_49106,N_49245);
and UO_892 (O_892,N_49375,N_49044);
xnor UO_893 (O_893,N_49025,N_49478);
xnor UO_894 (O_894,N_49428,N_49225);
nor UO_895 (O_895,N_49476,N_49671);
and UO_896 (O_896,N_49469,N_49156);
xnor UO_897 (O_897,N_49034,N_49755);
xor UO_898 (O_898,N_49447,N_49463);
and UO_899 (O_899,N_49365,N_49779);
nand UO_900 (O_900,N_49694,N_49092);
nor UO_901 (O_901,N_49700,N_49287);
or UO_902 (O_902,N_49975,N_49535);
or UO_903 (O_903,N_49419,N_49723);
nand UO_904 (O_904,N_49186,N_49739);
nand UO_905 (O_905,N_49406,N_49935);
nor UO_906 (O_906,N_49599,N_49816);
nor UO_907 (O_907,N_49730,N_49257);
nand UO_908 (O_908,N_49686,N_49349);
and UO_909 (O_909,N_49382,N_49322);
nand UO_910 (O_910,N_49404,N_49245);
xnor UO_911 (O_911,N_49382,N_49514);
and UO_912 (O_912,N_49339,N_49444);
or UO_913 (O_913,N_49594,N_49930);
nand UO_914 (O_914,N_49955,N_49219);
or UO_915 (O_915,N_49277,N_49995);
nand UO_916 (O_916,N_49049,N_49221);
or UO_917 (O_917,N_49023,N_49419);
or UO_918 (O_918,N_49631,N_49939);
and UO_919 (O_919,N_49575,N_49863);
and UO_920 (O_920,N_49068,N_49765);
nor UO_921 (O_921,N_49421,N_49415);
or UO_922 (O_922,N_49833,N_49176);
nand UO_923 (O_923,N_49763,N_49269);
and UO_924 (O_924,N_49471,N_49206);
nand UO_925 (O_925,N_49547,N_49291);
or UO_926 (O_926,N_49713,N_49700);
or UO_927 (O_927,N_49415,N_49163);
nand UO_928 (O_928,N_49867,N_49933);
or UO_929 (O_929,N_49474,N_49052);
xnor UO_930 (O_930,N_49245,N_49721);
or UO_931 (O_931,N_49670,N_49337);
and UO_932 (O_932,N_49653,N_49732);
or UO_933 (O_933,N_49609,N_49707);
xor UO_934 (O_934,N_49032,N_49104);
nand UO_935 (O_935,N_49824,N_49687);
or UO_936 (O_936,N_49665,N_49628);
and UO_937 (O_937,N_49227,N_49204);
nor UO_938 (O_938,N_49150,N_49072);
xor UO_939 (O_939,N_49476,N_49570);
xor UO_940 (O_940,N_49531,N_49158);
or UO_941 (O_941,N_49024,N_49580);
nand UO_942 (O_942,N_49147,N_49439);
nor UO_943 (O_943,N_49059,N_49595);
or UO_944 (O_944,N_49465,N_49615);
nor UO_945 (O_945,N_49784,N_49200);
and UO_946 (O_946,N_49198,N_49253);
nor UO_947 (O_947,N_49603,N_49043);
xor UO_948 (O_948,N_49322,N_49607);
xnor UO_949 (O_949,N_49150,N_49144);
nor UO_950 (O_950,N_49674,N_49251);
xnor UO_951 (O_951,N_49703,N_49310);
or UO_952 (O_952,N_49201,N_49731);
nor UO_953 (O_953,N_49564,N_49143);
or UO_954 (O_954,N_49586,N_49886);
xor UO_955 (O_955,N_49615,N_49014);
and UO_956 (O_956,N_49912,N_49083);
and UO_957 (O_957,N_49241,N_49134);
xnor UO_958 (O_958,N_49585,N_49020);
and UO_959 (O_959,N_49261,N_49779);
and UO_960 (O_960,N_49958,N_49545);
and UO_961 (O_961,N_49266,N_49140);
xor UO_962 (O_962,N_49116,N_49987);
nand UO_963 (O_963,N_49898,N_49074);
nand UO_964 (O_964,N_49306,N_49152);
or UO_965 (O_965,N_49395,N_49828);
or UO_966 (O_966,N_49141,N_49124);
or UO_967 (O_967,N_49575,N_49799);
or UO_968 (O_968,N_49773,N_49969);
or UO_969 (O_969,N_49499,N_49344);
xor UO_970 (O_970,N_49114,N_49611);
and UO_971 (O_971,N_49690,N_49123);
and UO_972 (O_972,N_49269,N_49429);
and UO_973 (O_973,N_49527,N_49800);
or UO_974 (O_974,N_49963,N_49209);
nand UO_975 (O_975,N_49394,N_49995);
or UO_976 (O_976,N_49900,N_49627);
nor UO_977 (O_977,N_49357,N_49545);
nor UO_978 (O_978,N_49947,N_49257);
and UO_979 (O_979,N_49463,N_49282);
or UO_980 (O_980,N_49280,N_49539);
or UO_981 (O_981,N_49725,N_49912);
nor UO_982 (O_982,N_49680,N_49789);
and UO_983 (O_983,N_49449,N_49795);
nand UO_984 (O_984,N_49006,N_49380);
nor UO_985 (O_985,N_49291,N_49540);
nand UO_986 (O_986,N_49434,N_49684);
and UO_987 (O_987,N_49121,N_49943);
xor UO_988 (O_988,N_49586,N_49344);
nor UO_989 (O_989,N_49374,N_49317);
or UO_990 (O_990,N_49382,N_49233);
nand UO_991 (O_991,N_49321,N_49015);
xor UO_992 (O_992,N_49541,N_49438);
nor UO_993 (O_993,N_49447,N_49677);
xor UO_994 (O_994,N_49083,N_49986);
or UO_995 (O_995,N_49631,N_49621);
xnor UO_996 (O_996,N_49756,N_49839);
and UO_997 (O_997,N_49752,N_49779);
nand UO_998 (O_998,N_49235,N_49710);
nor UO_999 (O_999,N_49647,N_49023);
nand UO_1000 (O_1000,N_49801,N_49218);
or UO_1001 (O_1001,N_49968,N_49465);
nor UO_1002 (O_1002,N_49719,N_49256);
and UO_1003 (O_1003,N_49935,N_49658);
xor UO_1004 (O_1004,N_49423,N_49066);
or UO_1005 (O_1005,N_49312,N_49791);
and UO_1006 (O_1006,N_49318,N_49367);
xor UO_1007 (O_1007,N_49527,N_49124);
xnor UO_1008 (O_1008,N_49412,N_49848);
nand UO_1009 (O_1009,N_49286,N_49777);
and UO_1010 (O_1010,N_49121,N_49212);
and UO_1011 (O_1011,N_49849,N_49282);
nor UO_1012 (O_1012,N_49551,N_49090);
or UO_1013 (O_1013,N_49435,N_49709);
nand UO_1014 (O_1014,N_49868,N_49804);
or UO_1015 (O_1015,N_49000,N_49959);
nand UO_1016 (O_1016,N_49831,N_49073);
and UO_1017 (O_1017,N_49999,N_49346);
or UO_1018 (O_1018,N_49359,N_49623);
and UO_1019 (O_1019,N_49092,N_49599);
xnor UO_1020 (O_1020,N_49541,N_49616);
and UO_1021 (O_1021,N_49452,N_49233);
nand UO_1022 (O_1022,N_49321,N_49115);
nand UO_1023 (O_1023,N_49141,N_49387);
xor UO_1024 (O_1024,N_49910,N_49354);
and UO_1025 (O_1025,N_49471,N_49656);
or UO_1026 (O_1026,N_49171,N_49183);
xor UO_1027 (O_1027,N_49060,N_49601);
xnor UO_1028 (O_1028,N_49940,N_49298);
or UO_1029 (O_1029,N_49356,N_49659);
xor UO_1030 (O_1030,N_49977,N_49040);
nor UO_1031 (O_1031,N_49975,N_49913);
xor UO_1032 (O_1032,N_49410,N_49736);
nor UO_1033 (O_1033,N_49884,N_49007);
or UO_1034 (O_1034,N_49132,N_49457);
nor UO_1035 (O_1035,N_49882,N_49383);
xnor UO_1036 (O_1036,N_49238,N_49083);
nor UO_1037 (O_1037,N_49798,N_49897);
nand UO_1038 (O_1038,N_49938,N_49784);
or UO_1039 (O_1039,N_49901,N_49770);
nand UO_1040 (O_1040,N_49149,N_49357);
xnor UO_1041 (O_1041,N_49587,N_49098);
and UO_1042 (O_1042,N_49250,N_49021);
nor UO_1043 (O_1043,N_49008,N_49791);
nor UO_1044 (O_1044,N_49658,N_49097);
and UO_1045 (O_1045,N_49380,N_49637);
or UO_1046 (O_1046,N_49189,N_49878);
xnor UO_1047 (O_1047,N_49454,N_49243);
or UO_1048 (O_1048,N_49497,N_49786);
nor UO_1049 (O_1049,N_49874,N_49452);
xnor UO_1050 (O_1050,N_49747,N_49140);
nand UO_1051 (O_1051,N_49818,N_49887);
or UO_1052 (O_1052,N_49816,N_49844);
and UO_1053 (O_1053,N_49714,N_49949);
and UO_1054 (O_1054,N_49137,N_49646);
nand UO_1055 (O_1055,N_49903,N_49845);
xor UO_1056 (O_1056,N_49063,N_49468);
nand UO_1057 (O_1057,N_49999,N_49881);
and UO_1058 (O_1058,N_49097,N_49127);
nand UO_1059 (O_1059,N_49356,N_49621);
xor UO_1060 (O_1060,N_49280,N_49925);
nor UO_1061 (O_1061,N_49146,N_49493);
and UO_1062 (O_1062,N_49195,N_49095);
xnor UO_1063 (O_1063,N_49745,N_49285);
xor UO_1064 (O_1064,N_49349,N_49467);
nand UO_1065 (O_1065,N_49595,N_49599);
and UO_1066 (O_1066,N_49383,N_49198);
xnor UO_1067 (O_1067,N_49648,N_49311);
nor UO_1068 (O_1068,N_49940,N_49789);
nand UO_1069 (O_1069,N_49571,N_49504);
or UO_1070 (O_1070,N_49489,N_49565);
nor UO_1071 (O_1071,N_49156,N_49695);
and UO_1072 (O_1072,N_49671,N_49738);
or UO_1073 (O_1073,N_49550,N_49284);
nor UO_1074 (O_1074,N_49857,N_49365);
nand UO_1075 (O_1075,N_49666,N_49508);
xnor UO_1076 (O_1076,N_49627,N_49674);
nand UO_1077 (O_1077,N_49134,N_49550);
nor UO_1078 (O_1078,N_49265,N_49022);
xor UO_1079 (O_1079,N_49413,N_49952);
nor UO_1080 (O_1080,N_49443,N_49005);
xnor UO_1081 (O_1081,N_49878,N_49064);
nor UO_1082 (O_1082,N_49322,N_49911);
xor UO_1083 (O_1083,N_49797,N_49354);
nor UO_1084 (O_1084,N_49001,N_49036);
xor UO_1085 (O_1085,N_49688,N_49591);
nor UO_1086 (O_1086,N_49198,N_49891);
or UO_1087 (O_1087,N_49434,N_49742);
nor UO_1088 (O_1088,N_49791,N_49016);
and UO_1089 (O_1089,N_49392,N_49246);
xor UO_1090 (O_1090,N_49226,N_49405);
or UO_1091 (O_1091,N_49337,N_49559);
and UO_1092 (O_1092,N_49769,N_49885);
or UO_1093 (O_1093,N_49388,N_49303);
and UO_1094 (O_1094,N_49716,N_49755);
and UO_1095 (O_1095,N_49316,N_49255);
nand UO_1096 (O_1096,N_49086,N_49741);
or UO_1097 (O_1097,N_49286,N_49926);
or UO_1098 (O_1098,N_49188,N_49503);
xor UO_1099 (O_1099,N_49610,N_49848);
nor UO_1100 (O_1100,N_49703,N_49777);
and UO_1101 (O_1101,N_49268,N_49170);
xor UO_1102 (O_1102,N_49687,N_49961);
and UO_1103 (O_1103,N_49430,N_49412);
nand UO_1104 (O_1104,N_49481,N_49977);
nand UO_1105 (O_1105,N_49654,N_49069);
or UO_1106 (O_1106,N_49943,N_49952);
and UO_1107 (O_1107,N_49691,N_49680);
nand UO_1108 (O_1108,N_49165,N_49800);
nand UO_1109 (O_1109,N_49066,N_49249);
or UO_1110 (O_1110,N_49874,N_49116);
or UO_1111 (O_1111,N_49041,N_49566);
and UO_1112 (O_1112,N_49883,N_49419);
nor UO_1113 (O_1113,N_49350,N_49816);
nor UO_1114 (O_1114,N_49738,N_49382);
and UO_1115 (O_1115,N_49649,N_49282);
xor UO_1116 (O_1116,N_49989,N_49786);
xnor UO_1117 (O_1117,N_49627,N_49227);
xor UO_1118 (O_1118,N_49008,N_49595);
nand UO_1119 (O_1119,N_49839,N_49179);
nand UO_1120 (O_1120,N_49295,N_49332);
nand UO_1121 (O_1121,N_49284,N_49115);
or UO_1122 (O_1122,N_49918,N_49792);
nor UO_1123 (O_1123,N_49658,N_49294);
and UO_1124 (O_1124,N_49768,N_49830);
and UO_1125 (O_1125,N_49437,N_49178);
nand UO_1126 (O_1126,N_49909,N_49327);
nand UO_1127 (O_1127,N_49688,N_49777);
or UO_1128 (O_1128,N_49970,N_49228);
or UO_1129 (O_1129,N_49004,N_49779);
and UO_1130 (O_1130,N_49292,N_49996);
nor UO_1131 (O_1131,N_49695,N_49654);
and UO_1132 (O_1132,N_49378,N_49072);
xnor UO_1133 (O_1133,N_49223,N_49133);
and UO_1134 (O_1134,N_49047,N_49111);
xnor UO_1135 (O_1135,N_49830,N_49422);
or UO_1136 (O_1136,N_49744,N_49461);
nand UO_1137 (O_1137,N_49155,N_49583);
nand UO_1138 (O_1138,N_49835,N_49693);
or UO_1139 (O_1139,N_49097,N_49154);
or UO_1140 (O_1140,N_49070,N_49227);
nor UO_1141 (O_1141,N_49850,N_49432);
nand UO_1142 (O_1142,N_49099,N_49119);
and UO_1143 (O_1143,N_49800,N_49575);
nand UO_1144 (O_1144,N_49404,N_49118);
and UO_1145 (O_1145,N_49911,N_49690);
xor UO_1146 (O_1146,N_49574,N_49433);
nand UO_1147 (O_1147,N_49879,N_49995);
xor UO_1148 (O_1148,N_49084,N_49335);
nor UO_1149 (O_1149,N_49670,N_49771);
nor UO_1150 (O_1150,N_49003,N_49037);
or UO_1151 (O_1151,N_49431,N_49703);
xnor UO_1152 (O_1152,N_49019,N_49699);
or UO_1153 (O_1153,N_49123,N_49086);
nor UO_1154 (O_1154,N_49613,N_49706);
xnor UO_1155 (O_1155,N_49794,N_49885);
and UO_1156 (O_1156,N_49723,N_49176);
or UO_1157 (O_1157,N_49556,N_49439);
or UO_1158 (O_1158,N_49472,N_49679);
nor UO_1159 (O_1159,N_49068,N_49713);
nand UO_1160 (O_1160,N_49163,N_49207);
or UO_1161 (O_1161,N_49751,N_49634);
nor UO_1162 (O_1162,N_49312,N_49169);
nor UO_1163 (O_1163,N_49032,N_49592);
or UO_1164 (O_1164,N_49690,N_49539);
nor UO_1165 (O_1165,N_49666,N_49882);
or UO_1166 (O_1166,N_49936,N_49502);
or UO_1167 (O_1167,N_49356,N_49624);
or UO_1168 (O_1168,N_49073,N_49769);
or UO_1169 (O_1169,N_49036,N_49598);
xor UO_1170 (O_1170,N_49689,N_49969);
or UO_1171 (O_1171,N_49465,N_49161);
nor UO_1172 (O_1172,N_49778,N_49038);
or UO_1173 (O_1173,N_49980,N_49850);
or UO_1174 (O_1174,N_49782,N_49806);
nor UO_1175 (O_1175,N_49955,N_49665);
and UO_1176 (O_1176,N_49749,N_49256);
nand UO_1177 (O_1177,N_49627,N_49176);
nor UO_1178 (O_1178,N_49969,N_49067);
xor UO_1179 (O_1179,N_49834,N_49818);
or UO_1180 (O_1180,N_49541,N_49308);
xnor UO_1181 (O_1181,N_49199,N_49273);
xor UO_1182 (O_1182,N_49584,N_49090);
or UO_1183 (O_1183,N_49011,N_49107);
and UO_1184 (O_1184,N_49966,N_49179);
xor UO_1185 (O_1185,N_49917,N_49093);
nor UO_1186 (O_1186,N_49361,N_49336);
nand UO_1187 (O_1187,N_49351,N_49957);
nand UO_1188 (O_1188,N_49833,N_49483);
or UO_1189 (O_1189,N_49504,N_49069);
xnor UO_1190 (O_1190,N_49018,N_49227);
or UO_1191 (O_1191,N_49588,N_49031);
and UO_1192 (O_1192,N_49374,N_49000);
and UO_1193 (O_1193,N_49812,N_49478);
nor UO_1194 (O_1194,N_49913,N_49963);
xnor UO_1195 (O_1195,N_49433,N_49317);
nand UO_1196 (O_1196,N_49061,N_49698);
xnor UO_1197 (O_1197,N_49753,N_49612);
and UO_1198 (O_1198,N_49168,N_49818);
nor UO_1199 (O_1199,N_49816,N_49845);
xor UO_1200 (O_1200,N_49565,N_49952);
xnor UO_1201 (O_1201,N_49487,N_49935);
nor UO_1202 (O_1202,N_49647,N_49496);
or UO_1203 (O_1203,N_49674,N_49660);
and UO_1204 (O_1204,N_49523,N_49121);
and UO_1205 (O_1205,N_49097,N_49036);
or UO_1206 (O_1206,N_49806,N_49595);
xor UO_1207 (O_1207,N_49250,N_49776);
nand UO_1208 (O_1208,N_49975,N_49020);
or UO_1209 (O_1209,N_49804,N_49793);
xnor UO_1210 (O_1210,N_49625,N_49294);
nand UO_1211 (O_1211,N_49116,N_49467);
or UO_1212 (O_1212,N_49373,N_49707);
and UO_1213 (O_1213,N_49130,N_49537);
or UO_1214 (O_1214,N_49291,N_49804);
nand UO_1215 (O_1215,N_49397,N_49060);
or UO_1216 (O_1216,N_49217,N_49876);
nor UO_1217 (O_1217,N_49206,N_49169);
and UO_1218 (O_1218,N_49684,N_49911);
nand UO_1219 (O_1219,N_49642,N_49489);
nor UO_1220 (O_1220,N_49789,N_49191);
and UO_1221 (O_1221,N_49925,N_49498);
and UO_1222 (O_1222,N_49173,N_49590);
xnor UO_1223 (O_1223,N_49254,N_49878);
or UO_1224 (O_1224,N_49815,N_49513);
nand UO_1225 (O_1225,N_49036,N_49300);
nor UO_1226 (O_1226,N_49167,N_49869);
nand UO_1227 (O_1227,N_49894,N_49306);
and UO_1228 (O_1228,N_49820,N_49103);
nand UO_1229 (O_1229,N_49071,N_49372);
xor UO_1230 (O_1230,N_49050,N_49976);
xor UO_1231 (O_1231,N_49990,N_49496);
nor UO_1232 (O_1232,N_49425,N_49347);
xnor UO_1233 (O_1233,N_49933,N_49215);
and UO_1234 (O_1234,N_49354,N_49080);
or UO_1235 (O_1235,N_49769,N_49683);
or UO_1236 (O_1236,N_49354,N_49485);
nor UO_1237 (O_1237,N_49655,N_49466);
and UO_1238 (O_1238,N_49107,N_49622);
nand UO_1239 (O_1239,N_49183,N_49122);
xor UO_1240 (O_1240,N_49793,N_49493);
nand UO_1241 (O_1241,N_49403,N_49809);
nor UO_1242 (O_1242,N_49707,N_49119);
xor UO_1243 (O_1243,N_49545,N_49169);
nor UO_1244 (O_1244,N_49651,N_49739);
or UO_1245 (O_1245,N_49741,N_49503);
nand UO_1246 (O_1246,N_49667,N_49606);
xnor UO_1247 (O_1247,N_49775,N_49554);
xor UO_1248 (O_1248,N_49604,N_49660);
or UO_1249 (O_1249,N_49057,N_49507);
or UO_1250 (O_1250,N_49013,N_49674);
and UO_1251 (O_1251,N_49364,N_49663);
and UO_1252 (O_1252,N_49168,N_49044);
and UO_1253 (O_1253,N_49196,N_49630);
nor UO_1254 (O_1254,N_49616,N_49907);
or UO_1255 (O_1255,N_49804,N_49110);
nor UO_1256 (O_1256,N_49380,N_49705);
or UO_1257 (O_1257,N_49215,N_49246);
nor UO_1258 (O_1258,N_49893,N_49833);
nand UO_1259 (O_1259,N_49266,N_49684);
nand UO_1260 (O_1260,N_49673,N_49024);
nand UO_1261 (O_1261,N_49903,N_49924);
xor UO_1262 (O_1262,N_49881,N_49268);
xnor UO_1263 (O_1263,N_49487,N_49949);
or UO_1264 (O_1264,N_49379,N_49818);
and UO_1265 (O_1265,N_49458,N_49733);
nor UO_1266 (O_1266,N_49221,N_49599);
nand UO_1267 (O_1267,N_49078,N_49429);
nand UO_1268 (O_1268,N_49387,N_49499);
nand UO_1269 (O_1269,N_49281,N_49233);
and UO_1270 (O_1270,N_49967,N_49081);
or UO_1271 (O_1271,N_49311,N_49494);
and UO_1272 (O_1272,N_49560,N_49558);
xnor UO_1273 (O_1273,N_49614,N_49385);
nand UO_1274 (O_1274,N_49758,N_49208);
xnor UO_1275 (O_1275,N_49043,N_49030);
nor UO_1276 (O_1276,N_49073,N_49535);
nor UO_1277 (O_1277,N_49325,N_49129);
nor UO_1278 (O_1278,N_49402,N_49570);
nor UO_1279 (O_1279,N_49693,N_49425);
nor UO_1280 (O_1280,N_49252,N_49044);
nor UO_1281 (O_1281,N_49469,N_49201);
nor UO_1282 (O_1282,N_49145,N_49303);
nand UO_1283 (O_1283,N_49947,N_49692);
nor UO_1284 (O_1284,N_49752,N_49320);
nor UO_1285 (O_1285,N_49890,N_49983);
or UO_1286 (O_1286,N_49476,N_49433);
nand UO_1287 (O_1287,N_49410,N_49072);
or UO_1288 (O_1288,N_49458,N_49286);
or UO_1289 (O_1289,N_49423,N_49277);
and UO_1290 (O_1290,N_49283,N_49953);
or UO_1291 (O_1291,N_49888,N_49554);
and UO_1292 (O_1292,N_49504,N_49005);
xor UO_1293 (O_1293,N_49582,N_49403);
and UO_1294 (O_1294,N_49506,N_49134);
or UO_1295 (O_1295,N_49519,N_49638);
xor UO_1296 (O_1296,N_49168,N_49067);
and UO_1297 (O_1297,N_49852,N_49019);
or UO_1298 (O_1298,N_49731,N_49249);
or UO_1299 (O_1299,N_49684,N_49160);
nor UO_1300 (O_1300,N_49976,N_49481);
or UO_1301 (O_1301,N_49803,N_49254);
xor UO_1302 (O_1302,N_49745,N_49435);
xor UO_1303 (O_1303,N_49057,N_49492);
nor UO_1304 (O_1304,N_49574,N_49108);
and UO_1305 (O_1305,N_49719,N_49570);
or UO_1306 (O_1306,N_49371,N_49195);
xnor UO_1307 (O_1307,N_49924,N_49571);
or UO_1308 (O_1308,N_49996,N_49266);
xnor UO_1309 (O_1309,N_49672,N_49826);
xor UO_1310 (O_1310,N_49150,N_49834);
and UO_1311 (O_1311,N_49328,N_49932);
or UO_1312 (O_1312,N_49398,N_49657);
nand UO_1313 (O_1313,N_49964,N_49680);
nor UO_1314 (O_1314,N_49445,N_49391);
and UO_1315 (O_1315,N_49408,N_49083);
nand UO_1316 (O_1316,N_49966,N_49019);
or UO_1317 (O_1317,N_49719,N_49281);
nor UO_1318 (O_1318,N_49786,N_49627);
and UO_1319 (O_1319,N_49976,N_49774);
nand UO_1320 (O_1320,N_49422,N_49217);
nand UO_1321 (O_1321,N_49210,N_49525);
nand UO_1322 (O_1322,N_49475,N_49694);
or UO_1323 (O_1323,N_49454,N_49341);
or UO_1324 (O_1324,N_49900,N_49181);
and UO_1325 (O_1325,N_49519,N_49618);
or UO_1326 (O_1326,N_49470,N_49557);
nand UO_1327 (O_1327,N_49984,N_49304);
nor UO_1328 (O_1328,N_49065,N_49071);
and UO_1329 (O_1329,N_49804,N_49674);
xnor UO_1330 (O_1330,N_49270,N_49232);
or UO_1331 (O_1331,N_49811,N_49840);
or UO_1332 (O_1332,N_49056,N_49212);
xnor UO_1333 (O_1333,N_49617,N_49596);
or UO_1334 (O_1334,N_49528,N_49572);
and UO_1335 (O_1335,N_49772,N_49090);
nand UO_1336 (O_1336,N_49152,N_49140);
nand UO_1337 (O_1337,N_49529,N_49370);
nand UO_1338 (O_1338,N_49579,N_49928);
xor UO_1339 (O_1339,N_49458,N_49083);
or UO_1340 (O_1340,N_49286,N_49102);
xnor UO_1341 (O_1341,N_49725,N_49481);
or UO_1342 (O_1342,N_49526,N_49515);
nor UO_1343 (O_1343,N_49364,N_49150);
and UO_1344 (O_1344,N_49322,N_49247);
nor UO_1345 (O_1345,N_49876,N_49053);
nand UO_1346 (O_1346,N_49894,N_49396);
and UO_1347 (O_1347,N_49785,N_49047);
or UO_1348 (O_1348,N_49473,N_49436);
and UO_1349 (O_1349,N_49968,N_49896);
or UO_1350 (O_1350,N_49666,N_49683);
nand UO_1351 (O_1351,N_49374,N_49179);
xnor UO_1352 (O_1352,N_49837,N_49833);
and UO_1353 (O_1353,N_49635,N_49511);
and UO_1354 (O_1354,N_49505,N_49836);
xor UO_1355 (O_1355,N_49174,N_49848);
nor UO_1356 (O_1356,N_49596,N_49882);
nor UO_1357 (O_1357,N_49867,N_49226);
and UO_1358 (O_1358,N_49970,N_49190);
or UO_1359 (O_1359,N_49637,N_49297);
and UO_1360 (O_1360,N_49202,N_49862);
nand UO_1361 (O_1361,N_49474,N_49404);
and UO_1362 (O_1362,N_49838,N_49819);
nand UO_1363 (O_1363,N_49033,N_49076);
or UO_1364 (O_1364,N_49138,N_49013);
nor UO_1365 (O_1365,N_49719,N_49564);
xor UO_1366 (O_1366,N_49051,N_49684);
and UO_1367 (O_1367,N_49139,N_49273);
nor UO_1368 (O_1368,N_49470,N_49294);
nor UO_1369 (O_1369,N_49049,N_49708);
and UO_1370 (O_1370,N_49097,N_49284);
xor UO_1371 (O_1371,N_49792,N_49564);
nor UO_1372 (O_1372,N_49015,N_49976);
nor UO_1373 (O_1373,N_49269,N_49073);
nand UO_1374 (O_1374,N_49582,N_49020);
and UO_1375 (O_1375,N_49692,N_49761);
nand UO_1376 (O_1376,N_49673,N_49465);
and UO_1377 (O_1377,N_49183,N_49733);
nor UO_1378 (O_1378,N_49196,N_49288);
and UO_1379 (O_1379,N_49129,N_49573);
xor UO_1380 (O_1380,N_49561,N_49100);
nand UO_1381 (O_1381,N_49801,N_49544);
nor UO_1382 (O_1382,N_49753,N_49411);
xnor UO_1383 (O_1383,N_49662,N_49598);
nand UO_1384 (O_1384,N_49565,N_49929);
xnor UO_1385 (O_1385,N_49600,N_49594);
or UO_1386 (O_1386,N_49415,N_49506);
and UO_1387 (O_1387,N_49428,N_49516);
or UO_1388 (O_1388,N_49447,N_49319);
and UO_1389 (O_1389,N_49763,N_49818);
and UO_1390 (O_1390,N_49257,N_49018);
nand UO_1391 (O_1391,N_49603,N_49312);
nand UO_1392 (O_1392,N_49662,N_49185);
nor UO_1393 (O_1393,N_49583,N_49788);
and UO_1394 (O_1394,N_49408,N_49004);
and UO_1395 (O_1395,N_49851,N_49212);
nor UO_1396 (O_1396,N_49707,N_49120);
xor UO_1397 (O_1397,N_49880,N_49925);
nor UO_1398 (O_1398,N_49226,N_49970);
xor UO_1399 (O_1399,N_49170,N_49119);
and UO_1400 (O_1400,N_49915,N_49584);
or UO_1401 (O_1401,N_49574,N_49829);
nor UO_1402 (O_1402,N_49495,N_49453);
nand UO_1403 (O_1403,N_49696,N_49138);
nand UO_1404 (O_1404,N_49673,N_49686);
nor UO_1405 (O_1405,N_49628,N_49322);
nand UO_1406 (O_1406,N_49465,N_49126);
and UO_1407 (O_1407,N_49444,N_49597);
nand UO_1408 (O_1408,N_49855,N_49396);
nand UO_1409 (O_1409,N_49613,N_49988);
nor UO_1410 (O_1410,N_49747,N_49955);
xor UO_1411 (O_1411,N_49529,N_49948);
xnor UO_1412 (O_1412,N_49631,N_49464);
or UO_1413 (O_1413,N_49731,N_49016);
xor UO_1414 (O_1414,N_49516,N_49509);
and UO_1415 (O_1415,N_49320,N_49773);
and UO_1416 (O_1416,N_49836,N_49730);
or UO_1417 (O_1417,N_49729,N_49000);
and UO_1418 (O_1418,N_49981,N_49998);
and UO_1419 (O_1419,N_49450,N_49571);
or UO_1420 (O_1420,N_49447,N_49725);
xor UO_1421 (O_1421,N_49800,N_49121);
nor UO_1422 (O_1422,N_49809,N_49505);
and UO_1423 (O_1423,N_49639,N_49331);
nor UO_1424 (O_1424,N_49239,N_49475);
xor UO_1425 (O_1425,N_49018,N_49362);
nor UO_1426 (O_1426,N_49265,N_49429);
or UO_1427 (O_1427,N_49035,N_49866);
or UO_1428 (O_1428,N_49126,N_49964);
or UO_1429 (O_1429,N_49711,N_49770);
or UO_1430 (O_1430,N_49525,N_49170);
and UO_1431 (O_1431,N_49605,N_49693);
nand UO_1432 (O_1432,N_49148,N_49018);
or UO_1433 (O_1433,N_49030,N_49535);
or UO_1434 (O_1434,N_49748,N_49869);
nor UO_1435 (O_1435,N_49555,N_49710);
nor UO_1436 (O_1436,N_49649,N_49775);
nand UO_1437 (O_1437,N_49746,N_49499);
or UO_1438 (O_1438,N_49838,N_49672);
or UO_1439 (O_1439,N_49874,N_49803);
or UO_1440 (O_1440,N_49262,N_49130);
and UO_1441 (O_1441,N_49587,N_49269);
or UO_1442 (O_1442,N_49113,N_49586);
xnor UO_1443 (O_1443,N_49246,N_49404);
or UO_1444 (O_1444,N_49402,N_49301);
or UO_1445 (O_1445,N_49731,N_49280);
nand UO_1446 (O_1446,N_49995,N_49737);
nand UO_1447 (O_1447,N_49905,N_49460);
nor UO_1448 (O_1448,N_49288,N_49697);
nor UO_1449 (O_1449,N_49280,N_49872);
and UO_1450 (O_1450,N_49319,N_49414);
and UO_1451 (O_1451,N_49481,N_49734);
nor UO_1452 (O_1452,N_49039,N_49623);
nand UO_1453 (O_1453,N_49938,N_49652);
xnor UO_1454 (O_1454,N_49319,N_49047);
nor UO_1455 (O_1455,N_49643,N_49677);
and UO_1456 (O_1456,N_49880,N_49782);
or UO_1457 (O_1457,N_49715,N_49075);
or UO_1458 (O_1458,N_49496,N_49669);
nand UO_1459 (O_1459,N_49092,N_49242);
and UO_1460 (O_1460,N_49821,N_49949);
or UO_1461 (O_1461,N_49973,N_49996);
xnor UO_1462 (O_1462,N_49572,N_49920);
and UO_1463 (O_1463,N_49209,N_49205);
nand UO_1464 (O_1464,N_49180,N_49949);
and UO_1465 (O_1465,N_49382,N_49412);
and UO_1466 (O_1466,N_49977,N_49466);
nor UO_1467 (O_1467,N_49397,N_49971);
nand UO_1468 (O_1468,N_49604,N_49718);
xor UO_1469 (O_1469,N_49400,N_49926);
nor UO_1470 (O_1470,N_49349,N_49062);
nand UO_1471 (O_1471,N_49248,N_49081);
xnor UO_1472 (O_1472,N_49744,N_49921);
nor UO_1473 (O_1473,N_49361,N_49788);
xnor UO_1474 (O_1474,N_49136,N_49344);
xnor UO_1475 (O_1475,N_49243,N_49758);
and UO_1476 (O_1476,N_49192,N_49971);
xnor UO_1477 (O_1477,N_49369,N_49316);
nor UO_1478 (O_1478,N_49964,N_49463);
xor UO_1479 (O_1479,N_49817,N_49595);
nand UO_1480 (O_1480,N_49857,N_49878);
xnor UO_1481 (O_1481,N_49317,N_49313);
and UO_1482 (O_1482,N_49578,N_49598);
and UO_1483 (O_1483,N_49381,N_49230);
or UO_1484 (O_1484,N_49848,N_49574);
xnor UO_1485 (O_1485,N_49734,N_49845);
and UO_1486 (O_1486,N_49803,N_49655);
xnor UO_1487 (O_1487,N_49259,N_49323);
nand UO_1488 (O_1488,N_49757,N_49129);
xnor UO_1489 (O_1489,N_49961,N_49501);
xnor UO_1490 (O_1490,N_49964,N_49452);
xnor UO_1491 (O_1491,N_49138,N_49799);
and UO_1492 (O_1492,N_49468,N_49535);
or UO_1493 (O_1493,N_49986,N_49786);
xor UO_1494 (O_1494,N_49314,N_49584);
xor UO_1495 (O_1495,N_49951,N_49417);
and UO_1496 (O_1496,N_49482,N_49021);
and UO_1497 (O_1497,N_49665,N_49177);
nand UO_1498 (O_1498,N_49640,N_49152);
nand UO_1499 (O_1499,N_49113,N_49004);
nor UO_1500 (O_1500,N_49249,N_49477);
and UO_1501 (O_1501,N_49097,N_49949);
or UO_1502 (O_1502,N_49736,N_49724);
and UO_1503 (O_1503,N_49239,N_49849);
and UO_1504 (O_1504,N_49294,N_49746);
and UO_1505 (O_1505,N_49247,N_49778);
or UO_1506 (O_1506,N_49431,N_49332);
nor UO_1507 (O_1507,N_49701,N_49586);
or UO_1508 (O_1508,N_49409,N_49598);
nor UO_1509 (O_1509,N_49545,N_49922);
xor UO_1510 (O_1510,N_49085,N_49089);
and UO_1511 (O_1511,N_49759,N_49748);
xor UO_1512 (O_1512,N_49660,N_49226);
and UO_1513 (O_1513,N_49266,N_49006);
nor UO_1514 (O_1514,N_49658,N_49469);
xnor UO_1515 (O_1515,N_49467,N_49298);
and UO_1516 (O_1516,N_49521,N_49562);
nor UO_1517 (O_1517,N_49745,N_49336);
and UO_1518 (O_1518,N_49989,N_49645);
nor UO_1519 (O_1519,N_49441,N_49398);
or UO_1520 (O_1520,N_49953,N_49081);
nor UO_1521 (O_1521,N_49151,N_49786);
xor UO_1522 (O_1522,N_49599,N_49086);
and UO_1523 (O_1523,N_49950,N_49703);
or UO_1524 (O_1524,N_49851,N_49014);
or UO_1525 (O_1525,N_49497,N_49850);
nor UO_1526 (O_1526,N_49833,N_49962);
or UO_1527 (O_1527,N_49904,N_49981);
xor UO_1528 (O_1528,N_49313,N_49965);
and UO_1529 (O_1529,N_49477,N_49928);
nand UO_1530 (O_1530,N_49957,N_49816);
nand UO_1531 (O_1531,N_49709,N_49882);
and UO_1532 (O_1532,N_49626,N_49667);
nand UO_1533 (O_1533,N_49882,N_49135);
nand UO_1534 (O_1534,N_49581,N_49255);
nand UO_1535 (O_1535,N_49145,N_49139);
nor UO_1536 (O_1536,N_49309,N_49263);
or UO_1537 (O_1537,N_49857,N_49487);
nand UO_1538 (O_1538,N_49987,N_49914);
nor UO_1539 (O_1539,N_49290,N_49993);
nand UO_1540 (O_1540,N_49435,N_49149);
nor UO_1541 (O_1541,N_49759,N_49989);
or UO_1542 (O_1542,N_49876,N_49348);
or UO_1543 (O_1543,N_49493,N_49350);
and UO_1544 (O_1544,N_49604,N_49922);
xor UO_1545 (O_1545,N_49448,N_49897);
and UO_1546 (O_1546,N_49875,N_49037);
nand UO_1547 (O_1547,N_49477,N_49561);
nor UO_1548 (O_1548,N_49435,N_49557);
nor UO_1549 (O_1549,N_49109,N_49850);
xnor UO_1550 (O_1550,N_49681,N_49425);
nand UO_1551 (O_1551,N_49831,N_49212);
nor UO_1552 (O_1552,N_49716,N_49880);
nor UO_1553 (O_1553,N_49576,N_49876);
nor UO_1554 (O_1554,N_49268,N_49365);
nand UO_1555 (O_1555,N_49363,N_49021);
and UO_1556 (O_1556,N_49796,N_49148);
nand UO_1557 (O_1557,N_49128,N_49609);
and UO_1558 (O_1558,N_49959,N_49364);
and UO_1559 (O_1559,N_49484,N_49662);
nor UO_1560 (O_1560,N_49939,N_49388);
and UO_1561 (O_1561,N_49357,N_49639);
nand UO_1562 (O_1562,N_49603,N_49563);
nand UO_1563 (O_1563,N_49380,N_49066);
nor UO_1564 (O_1564,N_49426,N_49053);
nor UO_1565 (O_1565,N_49100,N_49036);
xnor UO_1566 (O_1566,N_49717,N_49726);
nor UO_1567 (O_1567,N_49870,N_49734);
xor UO_1568 (O_1568,N_49615,N_49021);
or UO_1569 (O_1569,N_49224,N_49798);
nor UO_1570 (O_1570,N_49967,N_49649);
or UO_1571 (O_1571,N_49557,N_49988);
nor UO_1572 (O_1572,N_49939,N_49820);
and UO_1573 (O_1573,N_49540,N_49649);
and UO_1574 (O_1574,N_49482,N_49416);
nand UO_1575 (O_1575,N_49236,N_49115);
nor UO_1576 (O_1576,N_49776,N_49320);
xor UO_1577 (O_1577,N_49245,N_49415);
nor UO_1578 (O_1578,N_49767,N_49926);
or UO_1579 (O_1579,N_49970,N_49695);
nor UO_1580 (O_1580,N_49871,N_49348);
or UO_1581 (O_1581,N_49030,N_49120);
nor UO_1582 (O_1582,N_49994,N_49020);
nand UO_1583 (O_1583,N_49771,N_49731);
or UO_1584 (O_1584,N_49966,N_49882);
xnor UO_1585 (O_1585,N_49114,N_49776);
xnor UO_1586 (O_1586,N_49128,N_49005);
and UO_1587 (O_1587,N_49823,N_49572);
xnor UO_1588 (O_1588,N_49018,N_49803);
or UO_1589 (O_1589,N_49485,N_49523);
xnor UO_1590 (O_1590,N_49841,N_49308);
and UO_1591 (O_1591,N_49265,N_49561);
nor UO_1592 (O_1592,N_49052,N_49113);
or UO_1593 (O_1593,N_49874,N_49415);
and UO_1594 (O_1594,N_49468,N_49221);
xnor UO_1595 (O_1595,N_49690,N_49478);
or UO_1596 (O_1596,N_49470,N_49742);
nor UO_1597 (O_1597,N_49149,N_49926);
xor UO_1598 (O_1598,N_49999,N_49619);
nand UO_1599 (O_1599,N_49301,N_49178);
and UO_1600 (O_1600,N_49673,N_49691);
nor UO_1601 (O_1601,N_49801,N_49787);
xor UO_1602 (O_1602,N_49205,N_49937);
or UO_1603 (O_1603,N_49109,N_49684);
nand UO_1604 (O_1604,N_49789,N_49604);
nor UO_1605 (O_1605,N_49677,N_49475);
nand UO_1606 (O_1606,N_49437,N_49494);
and UO_1607 (O_1607,N_49069,N_49030);
nand UO_1608 (O_1608,N_49443,N_49631);
nor UO_1609 (O_1609,N_49945,N_49779);
nand UO_1610 (O_1610,N_49585,N_49750);
nor UO_1611 (O_1611,N_49460,N_49957);
nand UO_1612 (O_1612,N_49172,N_49953);
or UO_1613 (O_1613,N_49837,N_49187);
or UO_1614 (O_1614,N_49773,N_49425);
nor UO_1615 (O_1615,N_49052,N_49861);
xor UO_1616 (O_1616,N_49422,N_49262);
nor UO_1617 (O_1617,N_49056,N_49286);
xor UO_1618 (O_1618,N_49019,N_49666);
nand UO_1619 (O_1619,N_49458,N_49217);
or UO_1620 (O_1620,N_49914,N_49146);
xor UO_1621 (O_1621,N_49427,N_49853);
nand UO_1622 (O_1622,N_49871,N_49232);
xnor UO_1623 (O_1623,N_49037,N_49730);
or UO_1624 (O_1624,N_49144,N_49655);
or UO_1625 (O_1625,N_49164,N_49586);
and UO_1626 (O_1626,N_49776,N_49955);
or UO_1627 (O_1627,N_49628,N_49820);
or UO_1628 (O_1628,N_49505,N_49562);
or UO_1629 (O_1629,N_49475,N_49885);
or UO_1630 (O_1630,N_49852,N_49600);
xor UO_1631 (O_1631,N_49034,N_49170);
and UO_1632 (O_1632,N_49036,N_49246);
nand UO_1633 (O_1633,N_49138,N_49840);
and UO_1634 (O_1634,N_49376,N_49618);
and UO_1635 (O_1635,N_49112,N_49586);
xnor UO_1636 (O_1636,N_49743,N_49112);
or UO_1637 (O_1637,N_49495,N_49079);
or UO_1638 (O_1638,N_49587,N_49965);
and UO_1639 (O_1639,N_49905,N_49448);
or UO_1640 (O_1640,N_49664,N_49505);
and UO_1641 (O_1641,N_49173,N_49811);
nor UO_1642 (O_1642,N_49813,N_49865);
nand UO_1643 (O_1643,N_49754,N_49484);
nor UO_1644 (O_1644,N_49044,N_49967);
nor UO_1645 (O_1645,N_49560,N_49801);
and UO_1646 (O_1646,N_49510,N_49498);
or UO_1647 (O_1647,N_49922,N_49685);
xor UO_1648 (O_1648,N_49685,N_49693);
or UO_1649 (O_1649,N_49225,N_49335);
nand UO_1650 (O_1650,N_49751,N_49821);
or UO_1651 (O_1651,N_49604,N_49192);
nor UO_1652 (O_1652,N_49855,N_49335);
and UO_1653 (O_1653,N_49158,N_49020);
xnor UO_1654 (O_1654,N_49875,N_49074);
or UO_1655 (O_1655,N_49832,N_49961);
nand UO_1656 (O_1656,N_49086,N_49966);
nor UO_1657 (O_1657,N_49244,N_49224);
and UO_1658 (O_1658,N_49806,N_49343);
nand UO_1659 (O_1659,N_49323,N_49288);
nor UO_1660 (O_1660,N_49706,N_49195);
nand UO_1661 (O_1661,N_49595,N_49459);
xnor UO_1662 (O_1662,N_49167,N_49742);
or UO_1663 (O_1663,N_49692,N_49712);
xor UO_1664 (O_1664,N_49758,N_49560);
or UO_1665 (O_1665,N_49961,N_49304);
xnor UO_1666 (O_1666,N_49083,N_49581);
nand UO_1667 (O_1667,N_49893,N_49723);
nor UO_1668 (O_1668,N_49771,N_49559);
nand UO_1669 (O_1669,N_49861,N_49600);
nand UO_1670 (O_1670,N_49426,N_49944);
nand UO_1671 (O_1671,N_49459,N_49053);
and UO_1672 (O_1672,N_49741,N_49537);
nand UO_1673 (O_1673,N_49782,N_49645);
nor UO_1674 (O_1674,N_49312,N_49854);
and UO_1675 (O_1675,N_49049,N_49944);
and UO_1676 (O_1676,N_49396,N_49531);
or UO_1677 (O_1677,N_49544,N_49890);
xor UO_1678 (O_1678,N_49004,N_49338);
and UO_1679 (O_1679,N_49494,N_49518);
xor UO_1680 (O_1680,N_49830,N_49150);
xor UO_1681 (O_1681,N_49174,N_49661);
nand UO_1682 (O_1682,N_49001,N_49013);
nand UO_1683 (O_1683,N_49989,N_49285);
nand UO_1684 (O_1684,N_49258,N_49236);
xor UO_1685 (O_1685,N_49388,N_49889);
or UO_1686 (O_1686,N_49910,N_49158);
or UO_1687 (O_1687,N_49084,N_49020);
xor UO_1688 (O_1688,N_49816,N_49424);
and UO_1689 (O_1689,N_49073,N_49723);
and UO_1690 (O_1690,N_49058,N_49776);
xnor UO_1691 (O_1691,N_49462,N_49503);
and UO_1692 (O_1692,N_49941,N_49076);
xor UO_1693 (O_1693,N_49684,N_49371);
and UO_1694 (O_1694,N_49841,N_49218);
and UO_1695 (O_1695,N_49695,N_49257);
nor UO_1696 (O_1696,N_49694,N_49459);
or UO_1697 (O_1697,N_49119,N_49484);
xor UO_1698 (O_1698,N_49595,N_49109);
nand UO_1699 (O_1699,N_49015,N_49951);
or UO_1700 (O_1700,N_49601,N_49094);
nor UO_1701 (O_1701,N_49497,N_49366);
nand UO_1702 (O_1702,N_49364,N_49619);
nand UO_1703 (O_1703,N_49768,N_49825);
or UO_1704 (O_1704,N_49061,N_49350);
xor UO_1705 (O_1705,N_49500,N_49036);
or UO_1706 (O_1706,N_49092,N_49615);
or UO_1707 (O_1707,N_49007,N_49614);
nor UO_1708 (O_1708,N_49650,N_49891);
and UO_1709 (O_1709,N_49319,N_49535);
xnor UO_1710 (O_1710,N_49379,N_49744);
nor UO_1711 (O_1711,N_49451,N_49994);
or UO_1712 (O_1712,N_49276,N_49644);
xnor UO_1713 (O_1713,N_49274,N_49534);
xor UO_1714 (O_1714,N_49350,N_49974);
xor UO_1715 (O_1715,N_49241,N_49882);
xor UO_1716 (O_1716,N_49059,N_49429);
nand UO_1717 (O_1717,N_49023,N_49149);
nor UO_1718 (O_1718,N_49608,N_49316);
or UO_1719 (O_1719,N_49320,N_49463);
or UO_1720 (O_1720,N_49400,N_49164);
nor UO_1721 (O_1721,N_49190,N_49605);
xor UO_1722 (O_1722,N_49363,N_49550);
or UO_1723 (O_1723,N_49691,N_49855);
nor UO_1724 (O_1724,N_49799,N_49337);
xor UO_1725 (O_1725,N_49599,N_49171);
nor UO_1726 (O_1726,N_49014,N_49703);
nor UO_1727 (O_1727,N_49757,N_49417);
nand UO_1728 (O_1728,N_49734,N_49680);
and UO_1729 (O_1729,N_49832,N_49096);
xor UO_1730 (O_1730,N_49541,N_49095);
nand UO_1731 (O_1731,N_49163,N_49520);
or UO_1732 (O_1732,N_49081,N_49943);
nand UO_1733 (O_1733,N_49275,N_49354);
or UO_1734 (O_1734,N_49778,N_49447);
xnor UO_1735 (O_1735,N_49154,N_49094);
nor UO_1736 (O_1736,N_49383,N_49305);
xnor UO_1737 (O_1737,N_49013,N_49596);
or UO_1738 (O_1738,N_49364,N_49417);
xor UO_1739 (O_1739,N_49159,N_49232);
or UO_1740 (O_1740,N_49344,N_49972);
and UO_1741 (O_1741,N_49637,N_49386);
nand UO_1742 (O_1742,N_49402,N_49688);
or UO_1743 (O_1743,N_49053,N_49344);
or UO_1744 (O_1744,N_49530,N_49236);
nand UO_1745 (O_1745,N_49327,N_49318);
nor UO_1746 (O_1746,N_49340,N_49121);
xor UO_1747 (O_1747,N_49357,N_49123);
or UO_1748 (O_1748,N_49326,N_49283);
nand UO_1749 (O_1749,N_49362,N_49061);
xor UO_1750 (O_1750,N_49080,N_49023);
or UO_1751 (O_1751,N_49452,N_49949);
xor UO_1752 (O_1752,N_49746,N_49159);
or UO_1753 (O_1753,N_49882,N_49802);
or UO_1754 (O_1754,N_49346,N_49644);
nor UO_1755 (O_1755,N_49985,N_49885);
nand UO_1756 (O_1756,N_49858,N_49227);
xnor UO_1757 (O_1757,N_49820,N_49957);
xor UO_1758 (O_1758,N_49200,N_49317);
nand UO_1759 (O_1759,N_49169,N_49308);
nand UO_1760 (O_1760,N_49531,N_49957);
and UO_1761 (O_1761,N_49999,N_49062);
nor UO_1762 (O_1762,N_49030,N_49674);
or UO_1763 (O_1763,N_49460,N_49022);
and UO_1764 (O_1764,N_49411,N_49716);
nor UO_1765 (O_1765,N_49229,N_49337);
xnor UO_1766 (O_1766,N_49361,N_49906);
nor UO_1767 (O_1767,N_49342,N_49452);
or UO_1768 (O_1768,N_49297,N_49429);
or UO_1769 (O_1769,N_49081,N_49290);
nand UO_1770 (O_1770,N_49563,N_49621);
nand UO_1771 (O_1771,N_49963,N_49319);
xor UO_1772 (O_1772,N_49027,N_49298);
or UO_1773 (O_1773,N_49422,N_49829);
or UO_1774 (O_1774,N_49072,N_49325);
nand UO_1775 (O_1775,N_49110,N_49499);
or UO_1776 (O_1776,N_49404,N_49336);
nand UO_1777 (O_1777,N_49333,N_49798);
and UO_1778 (O_1778,N_49789,N_49779);
nand UO_1779 (O_1779,N_49090,N_49768);
nor UO_1780 (O_1780,N_49591,N_49430);
or UO_1781 (O_1781,N_49459,N_49290);
and UO_1782 (O_1782,N_49176,N_49396);
or UO_1783 (O_1783,N_49654,N_49232);
and UO_1784 (O_1784,N_49368,N_49455);
or UO_1785 (O_1785,N_49986,N_49380);
and UO_1786 (O_1786,N_49242,N_49750);
nand UO_1787 (O_1787,N_49514,N_49464);
xnor UO_1788 (O_1788,N_49536,N_49161);
nor UO_1789 (O_1789,N_49276,N_49330);
xnor UO_1790 (O_1790,N_49952,N_49378);
nand UO_1791 (O_1791,N_49210,N_49677);
xnor UO_1792 (O_1792,N_49870,N_49949);
nor UO_1793 (O_1793,N_49873,N_49912);
nor UO_1794 (O_1794,N_49196,N_49866);
nor UO_1795 (O_1795,N_49158,N_49625);
or UO_1796 (O_1796,N_49744,N_49493);
nand UO_1797 (O_1797,N_49049,N_49440);
nand UO_1798 (O_1798,N_49114,N_49775);
xor UO_1799 (O_1799,N_49222,N_49193);
or UO_1800 (O_1800,N_49551,N_49047);
nor UO_1801 (O_1801,N_49462,N_49530);
nand UO_1802 (O_1802,N_49266,N_49237);
xnor UO_1803 (O_1803,N_49445,N_49573);
xor UO_1804 (O_1804,N_49792,N_49090);
or UO_1805 (O_1805,N_49438,N_49895);
or UO_1806 (O_1806,N_49499,N_49268);
or UO_1807 (O_1807,N_49087,N_49788);
or UO_1808 (O_1808,N_49169,N_49591);
and UO_1809 (O_1809,N_49449,N_49446);
xor UO_1810 (O_1810,N_49388,N_49626);
nand UO_1811 (O_1811,N_49264,N_49681);
and UO_1812 (O_1812,N_49987,N_49230);
or UO_1813 (O_1813,N_49629,N_49633);
and UO_1814 (O_1814,N_49753,N_49277);
or UO_1815 (O_1815,N_49871,N_49765);
xnor UO_1816 (O_1816,N_49075,N_49673);
nor UO_1817 (O_1817,N_49397,N_49968);
nor UO_1818 (O_1818,N_49275,N_49696);
and UO_1819 (O_1819,N_49062,N_49902);
and UO_1820 (O_1820,N_49835,N_49324);
xor UO_1821 (O_1821,N_49112,N_49761);
xor UO_1822 (O_1822,N_49475,N_49992);
xnor UO_1823 (O_1823,N_49613,N_49877);
and UO_1824 (O_1824,N_49005,N_49424);
nand UO_1825 (O_1825,N_49957,N_49901);
nand UO_1826 (O_1826,N_49153,N_49089);
xor UO_1827 (O_1827,N_49804,N_49503);
or UO_1828 (O_1828,N_49435,N_49984);
nor UO_1829 (O_1829,N_49306,N_49511);
nand UO_1830 (O_1830,N_49239,N_49238);
nor UO_1831 (O_1831,N_49686,N_49448);
xor UO_1832 (O_1832,N_49901,N_49236);
nor UO_1833 (O_1833,N_49474,N_49090);
nand UO_1834 (O_1834,N_49193,N_49432);
or UO_1835 (O_1835,N_49898,N_49329);
xnor UO_1836 (O_1836,N_49599,N_49308);
xnor UO_1837 (O_1837,N_49479,N_49178);
or UO_1838 (O_1838,N_49875,N_49081);
and UO_1839 (O_1839,N_49355,N_49426);
or UO_1840 (O_1840,N_49754,N_49601);
xnor UO_1841 (O_1841,N_49399,N_49311);
or UO_1842 (O_1842,N_49760,N_49147);
nor UO_1843 (O_1843,N_49594,N_49083);
and UO_1844 (O_1844,N_49876,N_49829);
nand UO_1845 (O_1845,N_49609,N_49768);
or UO_1846 (O_1846,N_49913,N_49140);
nand UO_1847 (O_1847,N_49448,N_49906);
nand UO_1848 (O_1848,N_49479,N_49857);
nor UO_1849 (O_1849,N_49180,N_49719);
or UO_1850 (O_1850,N_49088,N_49242);
and UO_1851 (O_1851,N_49056,N_49552);
xnor UO_1852 (O_1852,N_49257,N_49600);
xnor UO_1853 (O_1853,N_49628,N_49007);
nor UO_1854 (O_1854,N_49788,N_49106);
or UO_1855 (O_1855,N_49834,N_49907);
or UO_1856 (O_1856,N_49406,N_49950);
nand UO_1857 (O_1857,N_49623,N_49414);
nor UO_1858 (O_1858,N_49641,N_49597);
or UO_1859 (O_1859,N_49050,N_49432);
and UO_1860 (O_1860,N_49502,N_49792);
nor UO_1861 (O_1861,N_49450,N_49115);
nor UO_1862 (O_1862,N_49031,N_49686);
and UO_1863 (O_1863,N_49119,N_49891);
nor UO_1864 (O_1864,N_49975,N_49843);
nor UO_1865 (O_1865,N_49992,N_49285);
xor UO_1866 (O_1866,N_49920,N_49506);
xnor UO_1867 (O_1867,N_49939,N_49549);
nand UO_1868 (O_1868,N_49556,N_49237);
xnor UO_1869 (O_1869,N_49682,N_49389);
nand UO_1870 (O_1870,N_49422,N_49929);
xor UO_1871 (O_1871,N_49516,N_49877);
and UO_1872 (O_1872,N_49981,N_49774);
xnor UO_1873 (O_1873,N_49784,N_49285);
nor UO_1874 (O_1874,N_49032,N_49188);
or UO_1875 (O_1875,N_49939,N_49299);
and UO_1876 (O_1876,N_49194,N_49368);
and UO_1877 (O_1877,N_49045,N_49352);
xnor UO_1878 (O_1878,N_49999,N_49827);
xnor UO_1879 (O_1879,N_49361,N_49074);
xnor UO_1880 (O_1880,N_49251,N_49762);
nand UO_1881 (O_1881,N_49454,N_49032);
xor UO_1882 (O_1882,N_49229,N_49471);
xnor UO_1883 (O_1883,N_49968,N_49158);
and UO_1884 (O_1884,N_49309,N_49770);
or UO_1885 (O_1885,N_49517,N_49406);
xnor UO_1886 (O_1886,N_49281,N_49877);
nor UO_1887 (O_1887,N_49147,N_49489);
or UO_1888 (O_1888,N_49734,N_49266);
nand UO_1889 (O_1889,N_49693,N_49022);
or UO_1890 (O_1890,N_49423,N_49188);
nand UO_1891 (O_1891,N_49430,N_49164);
and UO_1892 (O_1892,N_49362,N_49820);
nor UO_1893 (O_1893,N_49944,N_49537);
xnor UO_1894 (O_1894,N_49904,N_49594);
nor UO_1895 (O_1895,N_49753,N_49982);
and UO_1896 (O_1896,N_49520,N_49973);
and UO_1897 (O_1897,N_49708,N_49605);
xnor UO_1898 (O_1898,N_49517,N_49115);
nand UO_1899 (O_1899,N_49866,N_49362);
nor UO_1900 (O_1900,N_49620,N_49761);
nor UO_1901 (O_1901,N_49907,N_49394);
and UO_1902 (O_1902,N_49505,N_49297);
nor UO_1903 (O_1903,N_49271,N_49830);
xor UO_1904 (O_1904,N_49896,N_49725);
or UO_1905 (O_1905,N_49503,N_49235);
nand UO_1906 (O_1906,N_49122,N_49909);
or UO_1907 (O_1907,N_49036,N_49349);
or UO_1908 (O_1908,N_49758,N_49716);
or UO_1909 (O_1909,N_49642,N_49473);
and UO_1910 (O_1910,N_49339,N_49465);
or UO_1911 (O_1911,N_49104,N_49718);
or UO_1912 (O_1912,N_49609,N_49517);
nor UO_1913 (O_1913,N_49680,N_49995);
nand UO_1914 (O_1914,N_49975,N_49733);
nor UO_1915 (O_1915,N_49779,N_49220);
and UO_1916 (O_1916,N_49044,N_49488);
and UO_1917 (O_1917,N_49422,N_49725);
nor UO_1918 (O_1918,N_49861,N_49399);
nand UO_1919 (O_1919,N_49835,N_49641);
and UO_1920 (O_1920,N_49745,N_49390);
and UO_1921 (O_1921,N_49977,N_49604);
nor UO_1922 (O_1922,N_49021,N_49648);
xnor UO_1923 (O_1923,N_49740,N_49259);
xnor UO_1924 (O_1924,N_49134,N_49252);
and UO_1925 (O_1925,N_49443,N_49797);
or UO_1926 (O_1926,N_49708,N_49742);
xnor UO_1927 (O_1927,N_49610,N_49674);
xnor UO_1928 (O_1928,N_49749,N_49835);
nand UO_1929 (O_1929,N_49477,N_49086);
and UO_1930 (O_1930,N_49290,N_49759);
xor UO_1931 (O_1931,N_49943,N_49127);
nor UO_1932 (O_1932,N_49789,N_49718);
nor UO_1933 (O_1933,N_49167,N_49256);
and UO_1934 (O_1934,N_49010,N_49763);
xor UO_1935 (O_1935,N_49671,N_49683);
nor UO_1936 (O_1936,N_49140,N_49900);
or UO_1937 (O_1937,N_49787,N_49841);
or UO_1938 (O_1938,N_49247,N_49807);
nand UO_1939 (O_1939,N_49202,N_49112);
nand UO_1940 (O_1940,N_49171,N_49773);
nand UO_1941 (O_1941,N_49910,N_49923);
and UO_1942 (O_1942,N_49165,N_49863);
nand UO_1943 (O_1943,N_49631,N_49362);
nand UO_1944 (O_1944,N_49253,N_49772);
and UO_1945 (O_1945,N_49944,N_49706);
xor UO_1946 (O_1946,N_49072,N_49143);
and UO_1947 (O_1947,N_49562,N_49587);
nor UO_1948 (O_1948,N_49280,N_49011);
and UO_1949 (O_1949,N_49937,N_49068);
or UO_1950 (O_1950,N_49071,N_49484);
xor UO_1951 (O_1951,N_49880,N_49956);
and UO_1952 (O_1952,N_49388,N_49625);
nor UO_1953 (O_1953,N_49964,N_49176);
xnor UO_1954 (O_1954,N_49360,N_49145);
nor UO_1955 (O_1955,N_49292,N_49540);
nand UO_1956 (O_1956,N_49401,N_49927);
xnor UO_1957 (O_1957,N_49123,N_49215);
nand UO_1958 (O_1958,N_49573,N_49486);
nand UO_1959 (O_1959,N_49447,N_49613);
nand UO_1960 (O_1960,N_49266,N_49967);
or UO_1961 (O_1961,N_49631,N_49447);
nor UO_1962 (O_1962,N_49126,N_49532);
nor UO_1963 (O_1963,N_49019,N_49290);
or UO_1964 (O_1964,N_49342,N_49831);
xnor UO_1965 (O_1965,N_49824,N_49678);
and UO_1966 (O_1966,N_49180,N_49212);
nor UO_1967 (O_1967,N_49535,N_49002);
xor UO_1968 (O_1968,N_49910,N_49949);
and UO_1969 (O_1969,N_49393,N_49925);
or UO_1970 (O_1970,N_49465,N_49825);
xor UO_1971 (O_1971,N_49568,N_49794);
and UO_1972 (O_1972,N_49376,N_49284);
nand UO_1973 (O_1973,N_49589,N_49143);
nand UO_1974 (O_1974,N_49530,N_49317);
xor UO_1975 (O_1975,N_49557,N_49868);
nor UO_1976 (O_1976,N_49109,N_49466);
xnor UO_1977 (O_1977,N_49508,N_49784);
xor UO_1978 (O_1978,N_49589,N_49887);
nand UO_1979 (O_1979,N_49592,N_49849);
nor UO_1980 (O_1980,N_49757,N_49580);
xor UO_1981 (O_1981,N_49404,N_49676);
and UO_1982 (O_1982,N_49099,N_49680);
or UO_1983 (O_1983,N_49453,N_49926);
or UO_1984 (O_1984,N_49623,N_49467);
xnor UO_1985 (O_1985,N_49606,N_49377);
xor UO_1986 (O_1986,N_49747,N_49149);
or UO_1987 (O_1987,N_49677,N_49671);
or UO_1988 (O_1988,N_49117,N_49641);
nor UO_1989 (O_1989,N_49297,N_49605);
or UO_1990 (O_1990,N_49140,N_49672);
nand UO_1991 (O_1991,N_49314,N_49282);
nand UO_1992 (O_1992,N_49272,N_49781);
nor UO_1993 (O_1993,N_49340,N_49116);
xor UO_1994 (O_1994,N_49749,N_49309);
or UO_1995 (O_1995,N_49074,N_49628);
xor UO_1996 (O_1996,N_49547,N_49948);
nor UO_1997 (O_1997,N_49281,N_49001);
nor UO_1998 (O_1998,N_49748,N_49451);
and UO_1999 (O_1999,N_49098,N_49024);
nand UO_2000 (O_2000,N_49733,N_49014);
xnor UO_2001 (O_2001,N_49829,N_49995);
xor UO_2002 (O_2002,N_49603,N_49611);
and UO_2003 (O_2003,N_49084,N_49305);
xnor UO_2004 (O_2004,N_49770,N_49790);
and UO_2005 (O_2005,N_49847,N_49572);
or UO_2006 (O_2006,N_49750,N_49432);
xor UO_2007 (O_2007,N_49331,N_49240);
nand UO_2008 (O_2008,N_49008,N_49982);
xor UO_2009 (O_2009,N_49954,N_49384);
and UO_2010 (O_2010,N_49870,N_49619);
nand UO_2011 (O_2011,N_49468,N_49595);
nor UO_2012 (O_2012,N_49289,N_49144);
nand UO_2013 (O_2013,N_49887,N_49712);
and UO_2014 (O_2014,N_49105,N_49299);
nand UO_2015 (O_2015,N_49714,N_49281);
or UO_2016 (O_2016,N_49028,N_49768);
and UO_2017 (O_2017,N_49004,N_49544);
xor UO_2018 (O_2018,N_49597,N_49017);
nand UO_2019 (O_2019,N_49389,N_49790);
and UO_2020 (O_2020,N_49977,N_49336);
nor UO_2021 (O_2021,N_49017,N_49322);
nor UO_2022 (O_2022,N_49618,N_49194);
xnor UO_2023 (O_2023,N_49886,N_49145);
and UO_2024 (O_2024,N_49819,N_49159);
and UO_2025 (O_2025,N_49571,N_49223);
or UO_2026 (O_2026,N_49227,N_49650);
xor UO_2027 (O_2027,N_49579,N_49236);
or UO_2028 (O_2028,N_49109,N_49377);
and UO_2029 (O_2029,N_49654,N_49158);
and UO_2030 (O_2030,N_49698,N_49572);
xor UO_2031 (O_2031,N_49124,N_49664);
or UO_2032 (O_2032,N_49970,N_49078);
and UO_2033 (O_2033,N_49218,N_49731);
or UO_2034 (O_2034,N_49024,N_49695);
and UO_2035 (O_2035,N_49062,N_49938);
and UO_2036 (O_2036,N_49856,N_49189);
nand UO_2037 (O_2037,N_49562,N_49649);
nor UO_2038 (O_2038,N_49261,N_49023);
or UO_2039 (O_2039,N_49471,N_49043);
and UO_2040 (O_2040,N_49231,N_49830);
or UO_2041 (O_2041,N_49381,N_49829);
xnor UO_2042 (O_2042,N_49324,N_49999);
or UO_2043 (O_2043,N_49401,N_49147);
nand UO_2044 (O_2044,N_49212,N_49181);
or UO_2045 (O_2045,N_49508,N_49230);
nor UO_2046 (O_2046,N_49982,N_49708);
and UO_2047 (O_2047,N_49252,N_49906);
and UO_2048 (O_2048,N_49861,N_49005);
or UO_2049 (O_2049,N_49212,N_49855);
xnor UO_2050 (O_2050,N_49336,N_49243);
nor UO_2051 (O_2051,N_49027,N_49195);
xor UO_2052 (O_2052,N_49356,N_49670);
nor UO_2053 (O_2053,N_49805,N_49600);
nand UO_2054 (O_2054,N_49476,N_49348);
and UO_2055 (O_2055,N_49689,N_49977);
and UO_2056 (O_2056,N_49833,N_49670);
nor UO_2057 (O_2057,N_49867,N_49813);
nor UO_2058 (O_2058,N_49239,N_49811);
or UO_2059 (O_2059,N_49551,N_49337);
nor UO_2060 (O_2060,N_49069,N_49021);
or UO_2061 (O_2061,N_49843,N_49323);
xor UO_2062 (O_2062,N_49235,N_49919);
nand UO_2063 (O_2063,N_49987,N_49608);
nand UO_2064 (O_2064,N_49378,N_49268);
and UO_2065 (O_2065,N_49182,N_49461);
or UO_2066 (O_2066,N_49695,N_49567);
nand UO_2067 (O_2067,N_49562,N_49396);
or UO_2068 (O_2068,N_49618,N_49428);
and UO_2069 (O_2069,N_49869,N_49719);
nor UO_2070 (O_2070,N_49906,N_49279);
xor UO_2071 (O_2071,N_49091,N_49085);
or UO_2072 (O_2072,N_49569,N_49557);
and UO_2073 (O_2073,N_49422,N_49061);
or UO_2074 (O_2074,N_49014,N_49715);
xor UO_2075 (O_2075,N_49797,N_49866);
or UO_2076 (O_2076,N_49161,N_49804);
xor UO_2077 (O_2077,N_49069,N_49588);
nor UO_2078 (O_2078,N_49080,N_49821);
nor UO_2079 (O_2079,N_49738,N_49188);
xor UO_2080 (O_2080,N_49013,N_49929);
xor UO_2081 (O_2081,N_49465,N_49727);
xor UO_2082 (O_2082,N_49108,N_49166);
xor UO_2083 (O_2083,N_49626,N_49150);
nand UO_2084 (O_2084,N_49687,N_49380);
xnor UO_2085 (O_2085,N_49032,N_49389);
or UO_2086 (O_2086,N_49162,N_49446);
nand UO_2087 (O_2087,N_49987,N_49503);
and UO_2088 (O_2088,N_49961,N_49489);
xnor UO_2089 (O_2089,N_49359,N_49764);
or UO_2090 (O_2090,N_49232,N_49512);
or UO_2091 (O_2091,N_49640,N_49523);
nor UO_2092 (O_2092,N_49578,N_49839);
xnor UO_2093 (O_2093,N_49313,N_49941);
nor UO_2094 (O_2094,N_49006,N_49055);
nor UO_2095 (O_2095,N_49896,N_49514);
nor UO_2096 (O_2096,N_49760,N_49104);
xnor UO_2097 (O_2097,N_49978,N_49636);
and UO_2098 (O_2098,N_49997,N_49974);
xor UO_2099 (O_2099,N_49744,N_49134);
and UO_2100 (O_2100,N_49645,N_49737);
nand UO_2101 (O_2101,N_49764,N_49587);
or UO_2102 (O_2102,N_49466,N_49902);
and UO_2103 (O_2103,N_49494,N_49369);
xor UO_2104 (O_2104,N_49446,N_49066);
nand UO_2105 (O_2105,N_49389,N_49616);
or UO_2106 (O_2106,N_49573,N_49725);
and UO_2107 (O_2107,N_49918,N_49615);
xor UO_2108 (O_2108,N_49078,N_49900);
and UO_2109 (O_2109,N_49706,N_49398);
or UO_2110 (O_2110,N_49377,N_49256);
nand UO_2111 (O_2111,N_49798,N_49157);
or UO_2112 (O_2112,N_49036,N_49150);
and UO_2113 (O_2113,N_49492,N_49414);
nor UO_2114 (O_2114,N_49902,N_49236);
nand UO_2115 (O_2115,N_49647,N_49121);
and UO_2116 (O_2116,N_49708,N_49022);
and UO_2117 (O_2117,N_49550,N_49896);
nor UO_2118 (O_2118,N_49712,N_49756);
nand UO_2119 (O_2119,N_49841,N_49731);
nor UO_2120 (O_2120,N_49942,N_49507);
xor UO_2121 (O_2121,N_49430,N_49990);
or UO_2122 (O_2122,N_49246,N_49634);
and UO_2123 (O_2123,N_49521,N_49976);
or UO_2124 (O_2124,N_49555,N_49404);
nand UO_2125 (O_2125,N_49879,N_49977);
nor UO_2126 (O_2126,N_49868,N_49536);
xnor UO_2127 (O_2127,N_49667,N_49916);
or UO_2128 (O_2128,N_49519,N_49506);
or UO_2129 (O_2129,N_49082,N_49126);
xor UO_2130 (O_2130,N_49958,N_49378);
and UO_2131 (O_2131,N_49309,N_49280);
xnor UO_2132 (O_2132,N_49412,N_49543);
xor UO_2133 (O_2133,N_49178,N_49286);
nand UO_2134 (O_2134,N_49706,N_49182);
nor UO_2135 (O_2135,N_49963,N_49638);
and UO_2136 (O_2136,N_49560,N_49586);
nor UO_2137 (O_2137,N_49884,N_49021);
and UO_2138 (O_2138,N_49202,N_49706);
nor UO_2139 (O_2139,N_49391,N_49721);
nor UO_2140 (O_2140,N_49041,N_49684);
or UO_2141 (O_2141,N_49968,N_49431);
or UO_2142 (O_2142,N_49818,N_49420);
xnor UO_2143 (O_2143,N_49770,N_49137);
xnor UO_2144 (O_2144,N_49339,N_49483);
and UO_2145 (O_2145,N_49975,N_49277);
and UO_2146 (O_2146,N_49411,N_49118);
nand UO_2147 (O_2147,N_49154,N_49591);
and UO_2148 (O_2148,N_49054,N_49018);
xnor UO_2149 (O_2149,N_49803,N_49215);
or UO_2150 (O_2150,N_49659,N_49256);
and UO_2151 (O_2151,N_49209,N_49356);
or UO_2152 (O_2152,N_49095,N_49071);
or UO_2153 (O_2153,N_49155,N_49505);
nor UO_2154 (O_2154,N_49577,N_49851);
nor UO_2155 (O_2155,N_49585,N_49368);
nor UO_2156 (O_2156,N_49595,N_49158);
or UO_2157 (O_2157,N_49604,N_49646);
nor UO_2158 (O_2158,N_49450,N_49497);
nand UO_2159 (O_2159,N_49821,N_49314);
or UO_2160 (O_2160,N_49783,N_49735);
and UO_2161 (O_2161,N_49162,N_49984);
nand UO_2162 (O_2162,N_49552,N_49250);
nand UO_2163 (O_2163,N_49788,N_49899);
nor UO_2164 (O_2164,N_49813,N_49335);
nor UO_2165 (O_2165,N_49292,N_49706);
nor UO_2166 (O_2166,N_49300,N_49091);
nor UO_2167 (O_2167,N_49194,N_49903);
nand UO_2168 (O_2168,N_49780,N_49538);
nor UO_2169 (O_2169,N_49191,N_49430);
xnor UO_2170 (O_2170,N_49836,N_49957);
or UO_2171 (O_2171,N_49508,N_49999);
nand UO_2172 (O_2172,N_49404,N_49831);
nand UO_2173 (O_2173,N_49776,N_49138);
nor UO_2174 (O_2174,N_49332,N_49953);
xnor UO_2175 (O_2175,N_49307,N_49516);
xor UO_2176 (O_2176,N_49775,N_49804);
and UO_2177 (O_2177,N_49686,N_49490);
nand UO_2178 (O_2178,N_49662,N_49872);
or UO_2179 (O_2179,N_49595,N_49218);
nand UO_2180 (O_2180,N_49534,N_49745);
nor UO_2181 (O_2181,N_49459,N_49118);
xor UO_2182 (O_2182,N_49249,N_49467);
nor UO_2183 (O_2183,N_49803,N_49433);
and UO_2184 (O_2184,N_49399,N_49710);
nand UO_2185 (O_2185,N_49557,N_49537);
or UO_2186 (O_2186,N_49571,N_49095);
nor UO_2187 (O_2187,N_49671,N_49423);
and UO_2188 (O_2188,N_49391,N_49428);
xor UO_2189 (O_2189,N_49015,N_49684);
xor UO_2190 (O_2190,N_49723,N_49297);
nor UO_2191 (O_2191,N_49429,N_49727);
or UO_2192 (O_2192,N_49572,N_49962);
xor UO_2193 (O_2193,N_49630,N_49177);
nor UO_2194 (O_2194,N_49841,N_49999);
and UO_2195 (O_2195,N_49216,N_49921);
xor UO_2196 (O_2196,N_49545,N_49073);
xor UO_2197 (O_2197,N_49350,N_49007);
xor UO_2198 (O_2198,N_49304,N_49405);
or UO_2199 (O_2199,N_49218,N_49886);
and UO_2200 (O_2200,N_49978,N_49762);
or UO_2201 (O_2201,N_49429,N_49166);
nor UO_2202 (O_2202,N_49946,N_49919);
nor UO_2203 (O_2203,N_49301,N_49852);
xor UO_2204 (O_2204,N_49563,N_49920);
and UO_2205 (O_2205,N_49660,N_49250);
or UO_2206 (O_2206,N_49415,N_49626);
xnor UO_2207 (O_2207,N_49123,N_49266);
nor UO_2208 (O_2208,N_49622,N_49215);
nand UO_2209 (O_2209,N_49874,N_49406);
nor UO_2210 (O_2210,N_49035,N_49543);
and UO_2211 (O_2211,N_49769,N_49729);
xnor UO_2212 (O_2212,N_49923,N_49728);
and UO_2213 (O_2213,N_49441,N_49045);
nand UO_2214 (O_2214,N_49961,N_49781);
nand UO_2215 (O_2215,N_49427,N_49283);
nor UO_2216 (O_2216,N_49118,N_49795);
nor UO_2217 (O_2217,N_49414,N_49698);
nand UO_2218 (O_2218,N_49521,N_49174);
xnor UO_2219 (O_2219,N_49146,N_49660);
xnor UO_2220 (O_2220,N_49478,N_49835);
xnor UO_2221 (O_2221,N_49812,N_49268);
nor UO_2222 (O_2222,N_49586,N_49820);
xor UO_2223 (O_2223,N_49324,N_49146);
and UO_2224 (O_2224,N_49017,N_49018);
xnor UO_2225 (O_2225,N_49141,N_49330);
nand UO_2226 (O_2226,N_49086,N_49993);
nor UO_2227 (O_2227,N_49482,N_49903);
nor UO_2228 (O_2228,N_49526,N_49874);
or UO_2229 (O_2229,N_49337,N_49917);
nand UO_2230 (O_2230,N_49409,N_49487);
or UO_2231 (O_2231,N_49269,N_49804);
nand UO_2232 (O_2232,N_49538,N_49291);
nand UO_2233 (O_2233,N_49930,N_49452);
nand UO_2234 (O_2234,N_49936,N_49251);
and UO_2235 (O_2235,N_49959,N_49187);
xor UO_2236 (O_2236,N_49752,N_49209);
nor UO_2237 (O_2237,N_49275,N_49705);
nand UO_2238 (O_2238,N_49709,N_49105);
or UO_2239 (O_2239,N_49400,N_49987);
nor UO_2240 (O_2240,N_49704,N_49580);
and UO_2241 (O_2241,N_49356,N_49749);
nor UO_2242 (O_2242,N_49575,N_49297);
nor UO_2243 (O_2243,N_49704,N_49853);
xor UO_2244 (O_2244,N_49907,N_49879);
xor UO_2245 (O_2245,N_49791,N_49949);
nand UO_2246 (O_2246,N_49056,N_49191);
nor UO_2247 (O_2247,N_49495,N_49776);
xor UO_2248 (O_2248,N_49767,N_49944);
and UO_2249 (O_2249,N_49984,N_49497);
or UO_2250 (O_2250,N_49211,N_49818);
xor UO_2251 (O_2251,N_49501,N_49061);
and UO_2252 (O_2252,N_49790,N_49091);
nand UO_2253 (O_2253,N_49392,N_49402);
xnor UO_2254 (O_2254,N_49934,N_49025);
nor UO_2255 (O_2255,N_49324,N_49205);
xnor UO_2256 (O_2256,N_49565,N_49439);
nor UO_2257 (O_2257,N_49793,N_49751);
xor UO_2258 (O_2258,N_49960,N_49882);
nor UO_2259 (O_2259,N_49863,N_49402);
or UO_2260 (O_2260,N_49210,N_49918);
xor UO_2261 (O_2261,N_49761,N_49717);
and UO_2262 (O_2262,N_49340,N_49944);
or UO_2263 (O_2263,N_49484,N_49334);
nand UO_2264 (O_2264,N_49298,N_49214);
nand UO_2265 (O_2265,N_49759,N_49002);
nand UO_2266 (O_2266,N_49694,N_49510);
and UO_2267 (O_2267,N_49965,N_49277);
xnor UO_2268 (O_2268,N_49263,N_49876);
nor UO_2269 (O_2269,N_49116,N_49143);
nor UO_2270 (O_2270,N_49750,N_49263);
nand UO_2271 (O_2271,N_49637,N_49205);
nor UO_2272 (O_2272,N_49929,N_49900);
and UO_2273 (O_2273,N_49620,N_49254);
or UO_2274 (O_2274,N_49599,N_49708);
nor UO_2275 (O_2275,N_49207,N_49640);
nand UO_2276 (O_2276,N_49114,N_49479);
nor UO_2277 (O_2277,N_49722,N_49297);
xnor UO_2278 (O_2278,N_49257,N_49969);
and UO_2279 (O_2279,N_49430,N_49539);
nor UO_2280 (O_2280,N_49226,N_49787);
nand UO_2281 (O_2281,N_49887,N_49125);
nor UO_2282 (O_2282,N_49076,N_49519);
and UO_2283 (O_2283,N_49181,N_49240);
nor UO_2284 (O_2284,N_49059,N_49672);
and UO_2285 (O_2285,N_49793,N_49725);
nand UO_2286 (O_2286,N_49419,N_49343);
or UO_2287 (O_2287,N_49671,N_49541);
and UO_2288 (O_2288,N_49276,N_49945);
nand UO_2289 (O_2289,N_49099,N_49991);
nor UO_2290 (O_2290,N_49333,N_49713);
nand UO_2291 (O_2291,N_49511,N_49137);
and UO_2292 (O_2292,N_49378,N_49914);
xor UO_2293 (O_2293,N_49653,N_49447);
nand UO_2294 (O_2294,N_49971,N_49587);
xor UO_2295 (O_2295,N_49610,N_49093);
or UO_2296 (O_2296,N_49639,N_49805);
xor UO_2297 (O_2297,N_49562,N_49776);
nand UO_2298 (O_2298,N_49571,N_49843);
nor UO_2299 (O_2299,N_49683,N_49431);
nand UO_2300 (O_2300,N_49100,N_49814);
or UO_2301 (O_2301,N_49384,N_49073);
or UO_2302 (O_2302,N_49102,N_49401);
or UO_2303 (O_2303,N_49350,N_49288);
and UO_2304 (O_2304,N_49700,N_49886);
nand UO_2305 (O_2305,N_49831,N_49002);
xor UO_2306 (O_2306,N_49588,N_49281);
and UO_2307 (O_2307,N_49508,N_49727);
and UO_2308 (O_2308,N_49294,N_49240);
xor UO_2309 (O_2309,N_49557,N_49264);
nor UO_2310 (O_2310,N_49545,N_49219);
nor UO_2311 (O_2311,N_49335,N_49118);
or UO_2312 (O_2312,N_49140,N_49019);
and UO_2313 (O_2313,N_49451,N_49146);
nand UO_2314 (O_2314,N_49041,N_49403);
nand UO_2315 (O_2315,N_49285,N_49346);
and UO_2316 (O_2316,N_49748,N_49606);
or UO_2317 (O_2317,N_49897,N_49708);
and UO_2318 (O_2318,N_49466,N_49527);
nor UO_2319 (O_2319,N_49124,N_49938);
xnor UO_2320 (O_2320,N_49945,N_49450);
nor UO_2321 (O_2321,N_49353,N_49340);
nand UO_2322 (O_2322,N_49000,N_49389);
and UO_2323 (O_2323,N_49653,N_49401);
nor UO_2324 (O_2324,N_49521,N_49930);
and UO_2325 (O_2325,N_49102,N_49363);
and UO_2326 (O_2326,N_49149,N_49343);
nand UO_2327 (O_2327,N_49756,N_49548);
xnor UO_2328 (O_2328,N_49068,N_49312);
nand UO_2329 (O_2329,N_49425,N_49464);
nand UO_2330 (O_2330,N_49920,N_49671);
and UO_2331 (O_2331,N_49192,N_49534);
nand UO_2332 (O_2332,N_49948,N_49405);
or UO_2333 (O_2333,N_49814,N_49149);
nor UO_2334 (O_2334,N_49284,N_49440);
or UO_2335 (O_2335,N_49120,N_49460);
nor UO_2336 (O_2336,N_49759,N_49829);
nand UO_2337 (O_2337,N_49259,N_49632);
and UO_2338 (O_2338,N_49964,N_49817);
nor UO_2339 (O_2339,N_49785,N_49297);
and UO_2340 (O_2340,N_49268,N_49806);
nand UO_2341 (O_2341,N_49894,N_49224);
xnor UO_2342 (O_2342,N_49554,N_49543);
xor UO_2343 (O_2343,N_49692,N_49728);
nor UO_2344 (O_2344,N_49744,N_49410);
or UO_2345 (O_2345,N_49330,N_49725);
or UO_2346 (O_2346,N_49672,N_49489);
xor UO_2347 (O_2347,N_49770,N_49778);
or UO_2348 (O_2348,N_49767,N_49393);
xnor UO_2349 (O_2349,N_49380,N_49053);
and UO_2350 (O_2350,N_49919,N_49746);
nand UO_2351 (O_2351,N_49985,N_49326);
nor UO_2352 (O_2352,N_49817,N_49117);
or UO_2353 (O_2353,N_49970,N_49453);
nand UO_2354 (O_2354,N_49118,N_49597);
and UO_2355 (O_2355,N_49222,N_49562);
and UO_2356 (O_2356,N_49918,N_49602);
nand UO_2357 (O_2357,N_49412,N_49376);
nor UO_2358 (O_2358,N_49165,N_49587);
nand UO_2359 (O_2359,N_49792,N_49902);
and UO_2360 (O_2360,N_49538,N_49243);
nand UO_2361 (O_2361,N_49125,N_49401);
and UO_2362 (O_2362,N_49741,N_49872);
or UO_2363 (O_2363,N_49506,N_49906);
xor UO_2364 (O_2364,N_49975,N_49597);
or UO_2365 (O_2365,N_49503,N_49685);
nor UO_2366 (O_2366,N_49419,N_49605);
xor UO_2367 (O_2367,N_49273,N_49482);
or UO_2368 (O_2368,N_49788,N_49411);
nor UO_2369 (O_2369,N_49068,N_49924);
nor UO_2370 (O_2370,N_49163,N_49633);
nor UO_2371 (O_2371,N_49927,N_49717);
nand UO_2372 (O_2372,N_49472,N_49595);
xnor UO_2373 (O_2373,N_49962,N_49625);
and UO_2374 (O_2374,N_49646,N_49048);
xor UO_2375 (O_2375,N_49002,N_49153);
or UO_2376 (O_2376,N_49485,N_49665);
nand UO_2377 (O_2377,N_49871,N_49096);
xnor UO_2378 (O_2378,N_49535,N_49739);
and UO_2379 (O_2379,N_49131,N_49393);
nand UO_2380 (O_2380,N_49676,N_49127);
xor UO_2381 (O_2381,N_49517,N_49894);
and UO_2382 (O_2382,N_49358,N_49900);
nor UO_2383 (O_2383,N_49865,N_49886);
or UO_2384 (O_2384,N_49924,N_49077);
nand UO_2385 (O_2385,N_49619,N_49931);
and UO_2386 (O_2386,N_49095,N_49788);
xor UO_2387 (O_2387,N_49655,N_49918);
nand UO_2388 (O_2388,N_49541,N_49504);
and UO_2389 (O_2389,N_49873,N_49120);
and UO_2390 (O_2390,N_49397,N_49691);
or UO_2391 (O_2391,N_49849,N_49343);
nand UO_2392 (O_2392,N_49583,N_49393);
nor UO_2393 (O_2393,N_49919,N_49144);
xor UO_2394 (O_2394,N_49418,N_49637);
xor UO_2395 (O_2395,N_49337,N_49320);
or UO_2396 (O_2396,N_49977,N_49851);
and UO_2397 (O_2397,N_49137,N_49554);
or UO_2398 (O_2398,N_49503,N_49972);
xnor UO_2399 (O_2399,N_49922,N_49184);
nand UO_2400 (O_2400,N_49191,N_49875);
or UO_2401 (O_2401,N_49594,N_49897);
nor UO_2402 (O_2402,N_49512,N_49595);
xnor UO_2403 (O_2403,N_49676,N_49106);
xor UO_2404 (O_2404,N_49619,N_49438);
nor UO_2405 (O_2405,N_49584,N_49893);
or UO_2406 (O_2406,N_49173,N_49361);
or UO_2407 (O_2407,N_49820,N_49305);
nor UO_2408 (O_2408,N_49064,N_49095);
xor UO_2409 (O_2409,N_49013,N_49852);
nand UO_2410 (O_2410,N_49888,N_49542);
or UO_2411 (O_2411,N_49010,N_49935);
and UO_2412 (O_2412,N_49562,N_49268);
nand UO_2413 (O_2413,N_49332,N_49185);
and UO_2414 (O_2414,N_49230,N_49172);
and UO_2415 (O_2415,N_49516,N_49355);
or UO_2416 (O_2416,N_49098,N_49786);
or UO_2417 (O_2417,N_49499,N_49751);
and UO_2418 (O_2418,N_49815,N_49070);
nand UO_2419 (O_2419,N_49399,N_49462);
xor UO_2420 (O_2420,N_49433,N_49718);
or UO_2421 (O_2421,N_49474,N_49074);
nor UO_2422 (O_2422,N_49668,N_49660);
and UO_2423 (O_2423,N_49919,N_49873);
nor UO_2424 (O_2424,N_49864,N_49925);
nor UO_2425 (O_2425,N_49124,N_49593);
nor UO_2426 (O_2426,N_49756,N_49713);
and UO_2427 (O_2427,N_49402,N_49864);
or UO_2428 (O_2428,N_49550,N_49775);
nand UO_2429 (O_2429,N_49809,N_49421);
and UO_2430 (O_2430,N_49642,N_49533);
nor UO_2431 (O_2431,N_49994,N_49570);
xnor UO_2432 (O_2432,N_49403,N_49610);
and UO_2433 (O_2433,N_49774,N_49563);
nand UO_2434 (O_2434,N_49255,N_49888);
xnor UO_2435 (O_2435,N_49031,N_49158);
or UO_2436 (O_2436,N_49391,N_49537);
nand UO_2437 (O_2437,N_49413,N_49678);
nand UO_2438 (O_2438,N_49563,N_49387);
or UO_2439 (O_2439,N_49392,N_49269);
and UO_2440 (O_2440,N_49301,N_49039);
nor UO_2441 (O_2441,N_49670,N_49686);
nand UO_2442 (O_2442,N_49732,N_49586);
or UO_2443 (O_2443,N_49411,N_49196);
nor UO_2444 (O_2444,N_49905,N_49491);
nor UO_2445 (O_2445,N_49689,N_49718);
nand UO_2446 (O_2446,N_49168,N_49058);
nand UO_2447 (O_2447,N_49728,N_49976);
xnor UO_2448 (O_2448,N_49908,N_49954);
xor UO_2449 (O_2449,N_49472,N_49368);
nand UO_2450 (O_2450,N_49212,N_49274);
and UO_2451 (O_2451,N_49821,N_49421);
or UO_2452 (O_2452,N_49447,N_49874);
and UO_2453 (O_2453,N_49727,N_49870);
xnor UO_2454 (O_2454,N_49077,N_49232);
xnor UO_2455 (O_2455,N_49932,N_49452);
nor UO_2456 (O_2456,N_49166,N_49985);
nor UO_2457 (O_2457,N_49361,N_49737);
xor UO_2458 (O_2458,N_49578,N_49621);
or UO_2459 (O_2459,N_49197,N_49540);
and UO_2460 (O_2460,N_49282,N_49388);
xnor UO_2461 (O_2461,N_49368,N_49852);
nor UO_2462 (O_2462,N_49726,N_49834);
nor UO_2463 (O_2463,N_49956,N_49399);
or UO_2464 (O_2464,N_49316,N_49376);
nand UO_2465 (O_2465,N_49437,N_49956);
xor UO_2466 (O_2466,N_49161,N_49104);
xor UO_2467 (O_2467,N_49175,N_49240);
or UO_2468 (O_2468,N_49719,N_49280);
nor UO_2469 (O_2469,N_49928,N_49835);
or UO_2470 (O_2470,N_49182,N_49575);
nand UO_2471 (O_2471,N_49593,N_49892);
nor UO_2472 (O_2472,N_49199,N_49375);
xnor UO_2473 (O_2473,N_49126,N_49775);
or UO_2474 (O_2474,N_49640,N_49750);
nor UO_2475 (O_2475,N_49455,N_49468);
nand UO_2476 (O_2476,N_49733,N_49640);
nand UO_2477 (O_2477,N_49262,N_49472);
and UO_2478 (O_2478,N_49687,N_49757);
xnor UO_2479 (O_2479,N_49656,N_49173);
xor UO_2480 (O_2480,N_49248,N_49939);
or UO_2481 (O_2481,N_49697,N_49115);
or UO_2482 (O_2482,N_49739,N_49106);
or UO_2483 (O_2483,N_49963,N_49574);
and UO_2484 (O_2484,N_49085,N_49147);
and UO_2485 (O_2485,N_49690,N_49522);
xor UO_2486 (O_2486,N_49099,N_49776);
nand UO_2487 (O_2487,N_49278,N_49438);
or UO_2488 (O_2488,N_49455,N_49930);
nand UO_2489 (O_2489,N_49533,N_49496);
xor UO_2490 (O_2490,N_49890,N_49839);
or UO_2491 (O_2491,N_49318,N_49294);
and UO_2492 (O_2492,N_49001,N_49205);
xor UO_2493 (O_2493,N_49417,N_49745);
nor UO_2494 (O_2494,N_49506,N_49505);
or UO_2495 (O_2495,N_49449,N_49084);
and UO_2496 (O_2496,N_49028,N_49901);
nand UO_2497 (O_2497,N_49882,N_49245);
and UO_2498 (O_2498,N_49809,N_49361);
nand UO_2499 (O_2499,N_49564,N_49920);
and UO_2500 (O_2500,N_49976,N_49914);
and UO_2501 (O_2501,N_49367,N_49649);
xor UO_2502 (O_2502,N_49998,N_49727);
or UO_2503 (O_2503,N_49813,N_49482);
nor UO_2504 (O_2504,N_49850,N_49177);
nand UO_2505 (O_2505,N_49322,N_49431);
xnor UO_2506 (O_2506,N_49552,N_49537);
xnor UO_2507 (O_2507,N_49258,N_49143);
or UO_2508 (O_2508,N_49343,N_49990);
xnor UO_2509 (O_2509,N_49090,N_49391);
nand UO_2510 (O_2510,N_49614,N_49716);
and UO_2511 (O_2511,N_49917,N_49064);
and UO_2512 (O_2512,N_49517,N_49058);
xnor UO_2513 (O_2513,N_49281,N_49750);
or UO_2514 (O_2514,N_49619,N_49475);
nor UO_2515 (O_2515,N_49474,N_49680);
and UO_2516 (O_2516,N_49421,N_49110);
nand UO_2517 (O_2517,N_49032,N_49987);
xor UO_2518 (O_2518,N_49206,N_49180);
or UO_2519 (O_2519,N_49262,N_49250);
and UO_2520 (O_2520,N_49704,N_49978);
xor UO_2521 (O_2521,N_49361,N_49089);
or UO_2522 (O_2522,N_49106,N_49965);
xor UO_2523 (O_2523,N_49809,N_49100);
or UO_2524 (O_2524,N_49498,N_49040);
nor UO_2525 (O_2525,N_49585,N_49696);
xor UO_2526 (O_2526,N_49830,N_49994);
or UO_2527 (O_2527,N_49920,N_49743);
or UO_2528 (O_2528,N_49598,N_49925);
nor UO_2529 (O_2529,N_49056,N_49986);
or UO_2530 (O_2530,N_49514,N_49115);
xnor UO_2531 (O_2531,N_49342,N_49238);
nand UO_2532 (O_2532,N_49505,N_49743);
xor UO_2533 (O_2533,N_49915,N_49886);
xor UO_2534 (O_2534,N_49078,N_49941);
and UO_2535 (O_2535,N_49844,N_49789);
and UO_2536 (O_2536,N_49549,N_49133);
nand UO_2537 (O_2537,N_49504,N_49154);
nand UO_2538 (O_2538,N_49174,N_49398);
nor UO_2539 (O_2539,N_49306,N_49321);
xnor UO_2540 (O_2540,N_49418,N_49110);
nand UO_2541 (O_2541,N_49706,N_49523);
xor UO_2542 (O_2542,N_49316,N_49872);
or UO_2543 (O_2543,N_49800,N_49500);
xnor UO_2544 (O_2544,N_49809,N_49729);
and UO_2545 (O_2545,N_49449,N_49305);
and UO_2546 (O_2546,N_49053,N_49058);
and UO_2547 (O_2547,N_49826,N_49382);
or UO_2548 (O_2548,N_49234,N_49470);
or UO_2549 (O_2549,N_49459,N_49467);
xor UO_2550 (O_2550,N_49713,N_49289);
and UO_2551 (O_2551,N_49308,N_49243);
nand UO_2552 (O_2552,N_49542,N_49116);
nor UO_2553 (O_2553,N_49859,N_49080);
nor UO_2554 (O_2554,N_49950,N_49351);
nor UO_2555 (O_2555,N_49997,N_49658);
xnor UO_2556 (O_2556,N_49819,N_49847);
xnor UO_2557 (O_2557,N_49439,N_49295);
xnor UO_2558 (O_2558,N_49143,N_49997);
and UO_2559 (O_2559,N_49122,N_49799);
xnor UO_2560 (O_2560,N_49683,N_49484);
nor UO_2561 (O_2561,N_49504,N_49010);
nand UO_2562 (O_2562,N_49057,N_49175);
xor UO_2563 (O_2563,N_49798,N_49095);
nor UO_2564 (O_2564,N_49003,N_49124);
xnor UO_2565 (O_2565,N_49565,N_49228);
xnor UO_2566 (O_2566,N_49378,N_49350);
nand UO_2567 (O_2567,N_49473,N_49724);
nand UO_2568 (O_2568,N_49288,N_49311);
xnor UO_2569 (O_2569,N_49854,N_49736);
or UO_2570 (O_2570,N_49389,N_49657);
and UO_2571 (O_2571,N_49867,N_49327);
and UO_2572 (O_2572,N_49273,N_49695);
nand UO_2573 (O_2573,N_49329,N_49160);
nand UO_2574 (O_2574,N_49052,N_49015);
nor UO_2575 (O_2575,N_49963,N_49987);
nand UO_2576 (O_2576,N_49991,N_49121);
and UO_2577 (O_2577,N_49903,N_49533);
xor UO_2578 (O_2578,N_49310,N_49850);
and UO_2579 (O_2579,N_49287,N_49270);
xnor UO_2580 (O_2580,N_49446,N_49611);
nand UO_2581 (O_2581,N_49366,N_49084);
or UO_2582 (O_2582,N_49783,N_49471);
nor UO_2583 (O_2583,N_49772,N_49695);
or UO_2584 (O_2584,N_49716,N_49125);
nand UO_2585 (O_2585,N_49727,N_49132);
or UO_2586 (O_2586,N_49001,N_49132);
or UO_2587 (O_2587,N_49768,N_49166);
xor UO_2588 (O_2588,N_49360,N_49600);
nand UO_2589 (O_2589,N_49179,N_49382);
xor UO_2590 (O_2590,N_49387,N_49438);
xor UO_2591 (O_2591,N_49905,N_49167);
or UO_2592 (O_2592,N_49601,N_49398);
or UO_2593 (O_2593,N_49535,N_49129);
nand UO_2594 (O_2594,N_49629,N_49329);
or UO_2595 (O_2595,N_49530,N_49267);
or UO_2596 (O_2596,N_49730,N_49336);
xnor UO_2597 (O_2597,N_49085,N_49063);
nor UO_2598 (O_2598,N_49712,N_49854);
or UO_2599 (O_2599,N_49774,N_49038);
and UO_2600 (O_2600,N_49455,N_49217);
and UO_2601 (O_2601,N_49934,N_49070);
nor UO_2602 (O_2602,N_49395,N_49548);
nand UO_2603 (O_2603,N_49021,N_49805);
or UO_2604 (O_2604,N_49518,N_49480);
xor UO_2605 (O_2605,N_49626,N_49551);
or UO_2606 (O_2606,N_49455,N_49372);
and UO_2607 (O_2607,N_49485,N_49903);
or UO_2608 (O_2608,N_49073,N_49469);
or UO_2609 (O_2609,N_49211,N_49571);
nor UO_2610 (O_2610,N_49320,N_49548);
nand UO_2611 (O_2611,N_49659,N_49372);
or UO_2612 (O_2612,N_49977,N_49937);
nor UO_2613 (O_2613,N_49466,N_49100);
nand UO_2614 (O_2614,N_49438,N_49352);
nor UO_2615 (O_2615,N_49717,N_49697);
nand UO_2616 (O_2616,N_49739,N_49515);
xnor UO_2617 (O_2617,N_49511,N_49113);
and UO_2618 (O_2618,N_49577,N_49079);
and UO_2619 (O_2619,N_49808,N_49936);
nor UO_2620 (O_2620,N_49442,N_49799);
nand UO_2621 (O_2621,N_49575,N_49051);
or UO_2622 (O_2622,N_49747,N_49454);
xor UO_2623 (O_2623,N_49269,N_49520);
and UO_2624 (O_2624,N_49888,N_49025);
and UO_2625 (O_2625,N_49327,N_49163);
or UO_2626 (O_2626,N_49697,N_49845);
nor UO_2627 (O_2627,N_49889,N_49317);
or UO_2628 (O_2628,N_49679,N_49718);
xnor UO_2629 (O_2629,N_49691,N_49416);
nor UO_2630 (O_2630,N_49733,N_49925);
xnor UO_2631 (O_2631,N_49094,N_49146);
nand UO_2632 (O_2632,N_49188,N_49145);
and UO_2633 (O_2633,N_49638,N_49603);
nand UO_2634 (O_2634,N_49551,N_49938);
nand UO_2635 (O_2635,N_49983,N_49393);
and UO_2636 (O_2636,N_49764,N_49653);
and UO_2637 (O_2637,N_49182,N_49977);
nor UO_2638 (O_2638,N_49342,N_49462);
or UO_2639 (O_2639,N_49255,N_49043);
or UO_2640 (O_2640,N_49094,N_49258);
xnor UO_2641 (O_2641,N_49722,N_49821);
nand UO_2642 (O_2642,N_49283,N_49246);
xor UO_2643 (O_2643,N_49988,N_49666);
and UO_2644 (O_2644,N_49996,N_49004);
or UO_2645 (O_2645,N_49102,N_49369);
and UO_2646 (O_2646,N_49054,N_49036);
or UO_2647 (O_2647,N_49547,N_49664);
nand UO_2648 (O_2648,N_49526,N_49922);
nor UO_2649 (O_2649,N_49107,N_49679);
or UO_2650 (O_2650,N_49855,N_49718);
xnor UO_2651 (O_2651,N_49112,N_49901);
nor UO_2652 (O_2652,N_49207,N_49729);
xnor UO_2653 (O_2653,N_49066,N_49788);
nand UO_2654 (O_2654,N_49334,N_49181);
and UO_2655 (O_2655,N_49763,N_49457);
nor UO_2656 (O_2656,N_49037,N_49113);
xor UO_2657 (O_2657,N_49043,N_49001);
and UO_2658 (O_2658,N_49077,N_49698);
xnor UO_2659 (O_2659,N_49561,N_49716);
or UO_2660 (O_2660,N_49991,N_49290);
nand UO_2661 (O_2661,N_49987,N_49706);
nor UO_2662 (O_2662,N_49076,N_49648);
and UO_2663 (O_2663,N_49935,N_49451);
xor UO_2664 (O_2664,N_49381,N_49119);
nand UO_2665 (O_2665,N_49125,N_49807);
or UO_2666 (O_2666,N_49804,N_49988);
or UO_2667 (O_2667,N_49117,N_49698);
or UO_2668 (O_2668,N_49229,N_49248);
and UO_2669 (O_2669,N_49645,N_49536);
or UO_2670 (O_2670,N_49044,N_49407);
or UO_2671 (O_2671,N_49462,N_49723);
or UO_2672 (O_2672,N_49386,N_49487);
and UO_2673 (O_2673,N_49413,N_49286);
xnor UO_2674 (O_2674,N_49887,N_49298);
nand UO_2675 (O_2675,N_49875,N_49230);
and UO_2676 (O_2676,N_49057,N_49030);
nand UO_2677 (O_2677,N_49328,N_49727);
nand UO_2678 (O_2678,N_49690,N_49204);
nand UO_2679 (O_2679,N_49159,N_49270);
and UO_2680 (O_2680,N_49747,N_49419);
or UO_2681 (O_2681,N_49414,N_49650);
nand UO_2682 (O_2682,N_49557,N_49866);
xnor UO_2683 (O_2683,N_49842,N_49113);
xor UO_2684 (O_2684,N_49192,N_49356);
or UO_2685 (O_2685,N_49218,N_49001);
xor UO_2686 (O_2686,N_49978,N_49435);
nand UO_2687 (O_2687,N_49150,N_49011);
nand UO_2688 (O_2688,N_49176,N_49406);
or UO_2689 (O_2689,N_49164,N_49709);
nor UO_2690 (O_2690,N_49418,N_49502);
or UO_2691 (O_2691,N_49647,N_49718);
nand UO_2692 (O_2692,N_49039,N_49497);
nand UO_2693 (O_2693,N_49237,N_49527);
or UO_2694 (O_2694,N_49319,N_49871);
or UO_2695 (O_2695,N_49657,N_49521);
or UO_2696 (O_2696,N_49217,N_49007);
nand UO_2697 (O_2697,N_49349,N_49817);
xor UO_2698 (O_2698,N_49292,N_49265);
and UO_2699 (O_2699,N_49097,N_49401);
nor UO_2700 (O_2700,N_49163,N_49374);
and UO_2701 (O_2701,N_49409,N_49749);
nor UO_2702 (O_2702,N_49954,N_49133);
nand UO_2703 (O_2703,N_49010,N_49866);
or UO_2704 (O_2704,N_49898,N_49246);
and UO_2705 (O_2705,N_49057,N_49169);
nor UO_2706 (O_2706,N_49492,N_49869);
and UO_2707 (O_2707,N_49175,N_49973);
nor UO_2708 (O_2708,N_49905,N_49380);
and UO_2709 (O_2709,N_49466,N_49457);
and UO_2710 (O_2710,N_49234,N_49775);
nor UO_2711 (O_2711,N_49883,N_49819);
xor UO_2712 (O_2712,N_49704,N_49602);
or UO_2713 (O_2713,N_49983,N_49022);
nor UO_2714 (O_2714,N_49193,N_49261);
nand UO_2715 (O_2715,N_49595,N_49047);
xnor UO_2716 (O_2716,N_49983,N_49871);
nand UO_2717 (O_2717,N_49249,N_49139);
nor UO_2718 (O_2718,N_49864,N_49171);
nand UO_2719 (O_2719,N_49214,N_49765);
and UO_2720 (O_2720,N_49982,N_49847);
xor UO_2721 (O_2721,N_49407,N_49824);
and UO_2722 (O_2722,N_49219,N_49914);
xnor UO_2723 (O_2723,N_49513,N_49287);
or UO_2724 (O_2724,N_49962,N_49832);
and UO_2725 (O_2725,N_49960,N_49711);
nor UO_2726 (O_2726,N_49484,N_49452);
or UO_2727 (O_2727,N_49526,N_49048);
and UO_2728 (O_2728,N_49641,N_49312);
and UO_2729 (O_2729,N_49958,N_49306);
and UO_2730 (O_2730,N_49444,N_49386);
nand UO_2731 (O_2731,N_49876,N_49636);
nand UO_2732 (O_2732,N_49611,N_49623);
and UO_2733 (O_2733,N_49901,N_49195);
xnor UO_2734 (O_2734,N_49148,N_49691);
nand UO_2735 (O_2735,N_49952,N_49099);
nor UO_2736 (O_2736,N_49223,N_49921);
nor UO_2737 (O_2737,N_49867,N_49399);
nor UO_2738 (O_2738,N_49720,N_49534);
or UO_2739 (O_2739,N_49072,N_49204);
nand UO_2740 (O_2740,N_49298,N_49282);
nor UO_2741 (O_2741,N_49550,N_49141);
xor UO_2742 (O_2742,N_49939,N_49162);
nor UO_2743 (O_2743,N_49348,N_49342);
or UO_2744 (O_2744,N_49437,N_49657);
and UO_2745 (O_2745,N_49759,N_49485);
or UO_2746 (O_2746,N_49786,N_49845);
xor UO_2747 (O_2747,N_49197,N_49925);
or UO_2748 (O_2748,N_49311,N_49242);
nor UO_2749 (O_2749,N_49997,N_49854);
nand UO_2750 (O_2750,N_49397,N_49488);
xor UO_2751 (O_2751,N_49785,N_49320);
nand UO_2752 (O_2752,N_49782,N_49124);
and UO_2753 (O_2753,N_49406,N_49368);
and UO_2754 (O_2754,N_49168,N_49013);
and UO_2755 (O_2755,N_49036,N_49180);
and UO_2756 (O_2756,N_49392,N_49114);
or UO_2757 (O_2757,N_49149,N_49806);
and UO_2758 (O_2758,N_49588,N_49327);
xnor UO_2759 (O_2759,N_49208,N_49218);
nand UO_2760 (O_2760,N_49597,N_49526);
nand UO_2761 (O_2761,N_49190,N_49916);
or UO_2762 (O_2762,N_49372,N_49600);
or UO_2763 (O_2763,N_49224,N_49184);
nand UO_2764 (O_2764,N_49128,N_49252);
nand UO_2765 (O_2765,N_49348,N_49300);
or UO_2766 (O_2766,N_49239,N_49501);
or UO_2767 (O_2767,N_49848,N_49365);
nor UO_2768 (O_2768,N_49653,N_49405);
nor UO_2769 (O_2769,N_49199,N_49914);
nor UO_2770 (O_2770,N_49512,N_49270);
nor UO_2771 (O_2771,N_49824,N_49164);
or UO_2772 (O_2772,N_49621,N_49229);
nand UO_2773 (O_2773,N_49627,N_49834);
nand UO_2774 (O_2774,N_49764,N_49208);
xor UO_2775 (O_2775,N_49996,N_49446);
and UO_2776 (O_2776,N_49516,N_49697);
nor UO_2777 (O_2777,N_49652,N_49241);
or UO_2778 (O_2778,N_49190,N_49893);
and UO_2779 (O_2779,N_49800,N_49847);
xnor UO_2780 (O_2780,N_49107,N_49489);
nand UO_2781 (O_2781,N_49734,N_49177);
nor UO_2782 (O_2782,N_49095,N_49080);
nor UO_2783 (O_2783,N_49857,N_49920);
and UO_2784 (O_2784,N_49129,N_49760);
nand UO_2785 (O_2785,N_49701,N_49175);
nand UO_2786 (O_2786,N_49577,N_49945);
nor UO_2787 (O_2787,N_49716,N_49341);
and UO_2788 (O_2788,N_49082,N_49859);
or UO_2789 (O_2789,N_49222,N_49411);
xnor UO_2790 (O_2790,N_49039,N_49338);
and UO_2791 (O_2791,N_49487,N_49224);
nand UO_2792 (O_2792,N_49959,N_49328);
nand UO_2793 (O_2793,N_49515,N_49561);
and UO_2794 (O_2794,N_49678,N_49233);
or UO_2795 (O_2795,N_49071,N_49170);
xnor UO_2796 (O_2796,N_49153,N_49228);
xor UO_2797 (O_2797,N_49616,N_49396);
nor UO_2798 (O_2798,N_49146,N_49976);
and UO_2799 (O_2799,N_49475,N_49457);
or UO_2800 (O_2800,N_49894,N_49557);
nor UO_2801 (O_2801,N_49449,N_49215);
or UO_2802 (O_2802,N_49253,N_49899);
and UO_2803 (O_2803,N_49943,N_49101);
nor UO_2804 (O_2804,N_49100,N_49859);
nand UO_2805 (O_2805,N_49938,N_49546);
or UO_2806 (O_2806,N_49160,N_49078);
nor UO_2807 (O_2807,N_49740,N_49683);
and UO_2808 (O_2808,N_49383,N_49381);
nand UO_2809 (O_2809,N_49307,N_49788);
xor UO_2810 (O_2810,N_49811,N_49425);
nor UO_2811 (O_2811,N_49664,N_49003);
xor UO_2812 (O_2812,N_49140,N_49529);
or UO_2813 (O_2813,N_49377,N_49345);
xnor UO_2814 (O_2814,N_49107,N_49798);
xnor UO_2815 (O_2815,N_49966,N_49716);
xnor UO_2816 (O_2816,N_49294,N_49351);
xnor UO_2817 (O_2817,N_49117,N_49583);
xor UO_2818 (O_2818,N_49249,N_49527);
or UO_2819 (O_2819,N_49849,N_49095);
nor UO_2820 (O_2820,N_49499,N_49319);
nand UO_2821 (O_2821,N_49994,N_49343);
nor UO_2822 (O_2822,N_49343,N_49378);
nand UO_2823 (O_2823,N_49503,N_49314);
or UO_2824 (O_2824,N_49962,N_49523);
and UO_2825 (O_2825,N_49461,N_49644);
nor UO_2826 (O_2826,N_49174,N_49186);
or UO_2827 (O_2827,N_49990,N_49252);
xnor UO_2828 (O_2828,N_49850,N_49108);
and UO_2829 (O_2829,N_49743,N_49911);
nor UO_2830 (O_2830,N_49179,N_49116);
and UO_2831 (O_2831,N_49097,N_49623);
nand UO_2832 (O_2832,N_49713,N_49194);
or UO_2833 (O_2833,N_49437,N_49376);
nand UO_2834 (O_2834,N_49545,N_49666);
xnor UO_2835 (O_2835,N_49072,N_49287);
or UO_2836 (O_2836,N_49637,N_49794);
nor UO_2837 (O_2837,N_49724,N_49097);
and UO_2838 (O_2838,N_49620,N_49025);
nand UO_2839 (O_2839,N_49486,N_49870);
nand UO_2840 (O_2840,N_49462,N_49381);
nand UO_2841 (O_2841,N_49056,N_49285);
nor UO_2842 (O_2842,N_49731,N_49031);
nand UO_2843 (O_2843,N_49451,N_49502);
and UO_2844 (O_2844,N_49963,N_49447);
or UO_2845 (O_2845,N_49595,N_49531);
nor UO_2846 (O_2846,N_49038,N_49429);
xor UO_2847 (O_2847,N_49083,N_49975);
and UO_2848 (O_2848,N_49775,N_49975);
or UO_2849 (O_2849,N_49511,N_49848);
and UO_2850 (O_2850,N_49350,N_49735);
xnor UO_2851 (O_2851,N_49835,N_49269);
nand UO_2852 (O_2852,N_49019,N_49598);
xnor UO_2853 (O_2853,N_49501,N_49110);
and UO_2854 (O_2854,N_49490,N_49777);
nand UO_2855 (O_2855,N_49693,N_49757);
xor UO_2856 (O_2856,N_49898,N_49941);
xor UO_2857 (O_2857,N_49945,N_49117);
or UO_2858 (O_2858,N_49391,N_49475);
nor UO_2859 (O_2859,N_49645,N_49614);
nor UO_2860 (O_2860,N_49801,N_49215);
xor UO_2861 (O_2861,N_49588,N_49632);
xnor UO_2862 (O_2862,N_49261,N_49594);
or UO_2863 (O_2863,N_49769,N_49293);
or UO_2864 (O_2864,N_49430,N_49420);
and UO_2865 (O_2865,N_49223,N_49609);
or UO_2866 (O_2866,N_49147,N_49667);
nand UO_2867 (O_2867,N_49264,N_49316);
xor UO_2868 (O_2868,N_49490,N_49331);
nand UO_2869 (O_2869,N_49151,N_49872);
and UO_2870 (O_2870,N_49548,N_49784);
and UO_2871 (O_2871,N_49731,N_49907);
nor UO_2872 (O_2872,N_49129,N_49213);
nand UO_2873 (O_2873,N_49856,N_49605);
and UO_2874 (O_2874,N_49925,N_49741);
and UO_2875 (O_2875,N_49708,N_49890);
nor UO_2876 (O_2876,N_49655,N_49936);
nor UO_2877 (O_2877,N_49779,N_49469);
or UO_2878 (O_2878,N_49919,N_49202);
or UO_2879 (O_2879,N_49831,N_49761);
nor UO_2880 (O_2880,N_49546,N_49828);
nand UO_2881 (O_2881,N_49852,N_49107);
nor UO_2882 (O_2882,N_49132,N_49863);
or UO_2883 (O_2883,N_49813,N_49807);
xnor UO_2884 (O_2884,N_49810,N_49395);
and UO_2885 (O_2885,N_49087,N_49331);
xnor UO_2886 (O_2886,N_49843,N_49565);
xnor UO_2887 (O_2887,N_49210,N_49383);
and UO_2888 (O_2888,N_49296,N_49967);
or UO_2889 (O_2889,N_49846,N_49635);
nor UO_2890 (O_2890,N_49612,N_49466);
or UO_2891 (O_2891,N_49337,N_49406);
or UO_2892 (O_2892,N_49595,N_49562);
and UO_2893 (O_2893,N_49450,N_49524);
nand UO_2894 (O_2894,N_49430,N_49410);
nor UO_2895 (O_2895,N_49252,N_49694);
nand UO_2896 (O_2896,N_49639,N_49125);
or UO_2897 (O_2897,N_49189,N_49009);
and UO_2898 (O_2898,N_49069,N_49025);
nor UO_2899 (O_2899,N_49774,N_49171);
nor UO_2900 (O_2900,N_49280,N_49770);
xor UO_2901 (O_2901,N_49853,N_49642);
nand UO_2902 (O_2902,N_49497,N_49013);
or UO_2903 (O_2903,N_49691,N_49128);
nor UO_2904 (O_2904,N_49270,N_49878);
nor UO_2905 (O_2905,N_49041,N_49086);
nand UO_2906 (O_2906,N_49275,N_49254);
or UO_2907 (O_2907,N_49061,N_49118);
nand UO_2908 (O_2908,N_49790,N_49775);
nor UO_2909 (O_2909,N_49061,N_49669);
xnor UO_2910 (O_2910,N_49424,N_49300);
xor UO_2911 (O_2911,N_49538,N_49161);
xor UO_2912 (O_2912,N_49229,N_49117);
nand UO_2913 (O_2913,N_49093,N_49718);
nor UO_2914 (O_2914,N_49207,N_49377);
and UO_2915 (O_2915,N_49782,N_49546);
nand UO_2916 (O_2916,N_49805,N_49679);
or UO_2917 (O_2917,N_49369,N_49344);
or UO_2918 (O_2918,N_49104,N_49079);
nand UO_2919 (O_2919,N_49445,N_49284);
or UO_2920 (O_2920,N_49707,N_49540);
nand UO_2921 (O_2921,N_49128,N_49227);
xnor UO_2922 (O_2922,N_49552,N_49882);
nor UO_2923 (O_2923,N_49471,N_49923);
and UO_2924 (O_2924,N_49790,N_49823);
and UO_2925 (O_2925,N_49301,N_49022);
nor UO_2926 (O_2926,N_49159,N_49642);
nor UO_2927 (O_2927,N_49557,N_49586);
nand UO_2928 (O_2928,N_49615,N_49097);
xor UO_2929 (O_2929,N_49314,N_49543);
nand UO_2930 (O_2930,N_49997,N_49911);
nand UO_2931 (O_2931,N_49309,N_49023);
nand UO_2932 (O_2932,N_49408,N_49015);
nor UO_2933 (O_2933,N_49109,N_49094);
or UO_2934 (O_2934,N_49821,N_49173);
nand UO_2935 (O_2935,N_49976,N_49758);
and UO_2936 (O_2936,N_49458,N_49385);
and UO_2937 (O_2937,N_49102,N_49475);
and UO_2938 (O_2938,N_49928,N_49436);
nand UO_2939 (O_2939,N_49126,N_49500);
or UO_2940 (O_2940,N_49782,N_49284);
or UO_2941 (O_2941,N_49642,N_49762);
nand UO_2942 (O_2942,N_49416,N_49699);
nand UO_2943 (O_2943,N_49400,N_49383);
xor UO_2944 (O_2944,N_49180,N_49913);
nor UO_2945 (O_2945,N_49907,N_49290);
xnor UO_2946 (O_2946,N_49092,N_49548);
xnor UO_2947 (O_2947,N_49688,N_49153);
or UO_2948 (O_2948,N_49851,N_49980);
nor UO_2949 (O_2949,N_49405,N_49714);
and UO_2950 (O_2950,N_49906,N_49207);
nor UO_2951 (O_2951,N_49268,N_49091);
xor UO_2952 (O_2952,N_49469,N_49525);
nand UO_2953 (O_2953,N_49642,N_49726);
xor UO_2954 (O_2954,N_49831,N_49540);
xor UO_2955 (O_2955,N_49105,N_49165);
or UO_2956 (O_2956,N_49850,N_49944);
nand UO_2957 (O_2957,N_49328,N_49571);
nand UO_2958 (O_2958,N_49736,N_49277);
and UO_2959 (O_2959,N_49340,N_49831);
nor UO_2960 (O_2960,N_49100,N_49030);
nand UO_2961 (O_2961,N_49580,N_49061);
nand UO_2962 (O_2962,N_49072,N_49789);
or UO_2963 (O_2963,N_49223,N_49660);
nand UO_2964 (O_2964,N_49489,N_49811);
xnor UO_2965 (O_2965,N_49524,N_49090);
nor UO_2966 (O_2966,N_49228,N_49307);
nor UO_2967 (O_2967,N_49964,N_49118);
or UO_2968 (O_2968,N_49083,N_49876);
and UO_2969 (O_2969,N_49854,N_49940);
and UO_2970 (O_2970,N_49945,N_49097);
and UO_2971 (O_2971,N_49889,N_49791);
and UO_2972 (O_2972,N_49030,N_49472);
xor UO_2973 (O_2973,N_49671,N_49947);
nand UO_2974 (O_2974,N_49797,N_49932);
and UO_2975 (O_2975,N_49598,N_49145);
nand UO_2976 (O_2976,N_49023,N_49642);
or UO_2977 (O_2977,N_49198,N_49350);
and UO_2978 (O_2978,N_49260,N_49798);
or UO_2979 (O_2979,N_49200,N_49248);
xnor UO_2980 (O_2980,N_49154,N_49061);
or UO_2981 (O_2981,N_49515,N_49450);
or UO_2982 (O_2982,N_49329,N_49504);
xnor UO_2983 (O_2983,N_49366,N_49240);
and UO_2984 (O_2984,N_49534,N_49700);
and UO_2985 (O_2985,N_49937,N_49393);
xnor UO_2986 (O_2986,N_49392,N_49112);
and UO_2987 (O_2987,N_49329,N_49848);
nand UO_2988 (O_2988,N_49713,N_49547);
nand UO_2989 (O_2989,N_49896,N_49049);
xnor UO_2990 (O_2990,N_49594,N_49383);
nand UO_2991 (O_2991,N_49031,N_49521);
and UO_2992 (O_2992,N_49751,N_49272);
xnor UO_2993 (O_2993,N_49237,N_49268);
nor UO_2994 (O_2994,N_49044,N_49963);
nand UO_2995 (O_2995,N_49443,N_49538);
xor UO_2996 (O_2996,N_49649,N_49563);
and UO_2997 (O_2997,N_49364,N_49010);
or UO_2998 (O_2998,N_49524,N_49347);
nand UO_2999 (O_2999,N_49335,N_49415);
nand UO_3000 (O_3000,N_49980,N_49524);
and UO_3001 (O_3001,N_49017,N_49135);
or UO_3002 (O_3002,N_49372,N_49781);
nand UO_3003 (O_3003,N_49079,N_49876);
or UO_3004 (O_3004,N_49666,N_49137);
nand UO_3005 (O_3005,N_49339,N_49726);
xnor UO_3006 (O_3006,N_49349,N_49396);
nor UO_3007 (O_3007,N_49658,N_49143);
xnor UO_3008 (O_3008,N_49238,N_49882);
and UO_3009 (O_3009,N_49805,N_49872);
xor UO_3010 (O_3010,N_49447,N_49848);
nand UO_3011 (O_3011,N_49752,N_49442);
and UO_3012 (O_3012,N_49466,N_49668);
nor UO_3013 (O_3013,N_49379,N_49772);
xor UO_3014 (O_3014,N_49028,N_49146);
xor UO_3015 (O_3015,N_49522,N_49614);
or UO_3016 (O_3016,N_49859,N_49669);
or UO_3017 (O_3017,N_49890,N_49562);
xnor UO_3018 (O_3018,N_49987,N_49115);
xor UO_3019 (O_3019,N_49151,N_49789);
nand UO_3020 (O_3020,N_49881,N_49600);
nor UO_3021 (O_3021,N_49535,N_49499);
or UO_3022 (O_3022,N_49159,N_49524);
xor UO_3023 (O_3023,N_49689,N_49829);
nand UO_3024 (O_3024,N_49336,N_49605);
xor UO_3025 (O_3025,N_49254,N_49956);
and UO_3026 (O_3026,N_49453,N_49433);
xor UO_3027 (O_3027,N_49815,N_49915);
nand UO_3028 (O_3028,N_49319,N_49708);
xor UO_3029 (O_3029,N_49056,N_49591);
nand UO_3030 (O_3030,N_49315,N_49861);
nor UO_3031 (O_3031,N_49898,N_49117);
xor UO_3032 (O_3032,N_49662,N_49045);
nor UO_3033 (O_3033,N_49498,N_49031);
and UO_3034 (O_3034,N_49683,N_49142);
nor UO_3035 (O_3035,N_49584,N_49673);
and UO_3036 (O_3036,N_49075,N_49900);
nor UO_3037 (O_3037,N_49452,N_49923);
and UO_3038 (O_3038,N_49621,N_49647);
nand UO_3039 (O_3039,N_49494,N_49440);
and UO_3040 (O_3040,N_49556,N_49888);
or UO_3041 (O_3041,N_49644,N_49580);
and UO_3042 (O_3042,N_49403,N_49434);
or UO_3043 (O_3043,N_49004,N_49720);
nor UO_3044 (O_3044,N_49249,N_49096);
and UO_3045 (O_3045,N_49399,N_49753);
xor UO_3046 (O_3046,N_49789,N_49471);
nor UO_3047 (O_3047,N_49492,N_49622);
xnor UO_3048 (O_3048,N_49044,N_49025);
or UO_3049 (O_3049,N_49506,N_49402);
and UO_3050 (O_3050,N_49001,N_49223);
nor UO_3051 (O_3051,N_49582,N_49481);
nor UO_3052 (O_3052,N_49167,N_49301);
or UO_3053 (O_3053,N_49488,N_49807);
or UO_3054 (O_3054,N_49734,N_49075);
and UO_3055 (O_3055,N_49534,N_49198);
nor UO_3056 (O_3056,N_49777,N_49717);
nand UO_3057 (O_3057,N_49864,N_49197);
xor UO_3058 (O_3058,N_49512,N_49384);
xor UO_3059 (O_3059,N_49747,N_49411);
nor UO_3060 (O_3060,N_49373,N_49516);
xor UO_3061 (O_3061,N_49535,N_49285);
xor UO_3062 (O_3062,N_49838,N_49048);
or UO_3063 (O_3063,N_49942,N_49261);
nor UO_3064 (O_3064,N_49818,N_49060);
nand UO_3065 (O_3065,N_49598,N_49583);
nor UO_3066 (O_3066,N_49240,N_49284);
nor UO_3067 (O_3067,N_49119,N_49038);
or UO_3068 (O_3068,N_49540,N_49395);
and UO_3069 (O_3069,N_49585,N_49545);
and UO_3070 (O_3070,N_49396,N_49134);
nor UO_3071 (O_3071,N_49038,N_49925);
xor UO_3072 (O_3072,N_49379,N_49629);
and UO_3073 (O_3073,N_49295,N_49016);
and UO_3074 (O_3074,N_49884,N_49080);
nor UO_3075 (O_3075,N_49412,N_49154);
nor UO_3076 (O_3076,N_49936,N_49326);
and UO_3077 (O_3077,N_49547,N_49868);
and UO_3078 (O_3078,N_49172,N_49401);
and UO_3079 (O_3079,N_49333,N_49793);
nor UO_3080 (O_3080,N_49223,N_49129);
xnor UO_3081 (O_3081,N_49433,N_49198);
or UO_3082 (O_3082,N_49614,N_49151);
nand UO_3083 (O_3083,N_49886,N_49259);
xor UO_3084 (O_3084,N_49758,N_49582);
nor UO_3085 (O_3085,N_49995,N_49083);
nand UO_3086 (O_3086,N_49316,N_49543);
nor UO_3087 (O_3087,N_49816,N_49917);
nor UO_3088 (O_3088,N_49147,N_49703);
nand UO_3089 (O_3089,N_49304,N_49977);
nand UO_3090 (O_3090,N_49157,N_49900);
xor UO_3091 (O_3091,N_49956,N_49628);
nor UO_3092 (O_3092,N_49867,N_49390);
xnor UO_3093 (O_3093,N_49529,N_49141);
or UO_3094 (O_3094,N_49543,N_49199);
or UO_3095 (O_3095,N_49132,N_49478);
nand UO_3096 (O_3096,N_49415,N_49294);
or UO_3097 (O_3097,N_49872,N_49300);
nand UO_3098 (O_3098,N_49245,N_49099);
or UO_3099 (O_3099,N_49824,N_49854);
and UO_3100 (O_3100,N_49603,N_49187);
nand UO_3101 (O_3101,N_49561,N_49371);
nand UO_3102 (O_3102,N_49210,N_49096);
xnor UO_3103 (O_3103,N_49227,N_49653);
xnor UO_3104 (O_3104,N_49686,N_49278);
nor UO_3105 (O_3105,N_49368,N_49995);
or UO_3106 (O_3106,N_49836,N_49698);
and UO_3107 (O_3107,N_49338,N_49675);
nor UO_3108 (O_3108,N_49112,N_49148);
xor UO_3109 (O_3109,N_49746,N_49343);
and UO_3110 (O_3110,N_49264,N_49686);
xnor UO_3111 (O_3111,N_49028,N_49301);
and UO_3112 (O_3112,N_49966,N_49286);
nor UO_3113 (O_3113,N_49173,N_49579);
nor UO_3114 (O_3114,N_49715,N_49648);
or UO_3115 (O_3115,N_49627,N_49004);
nor UO_3116 (O_3116,N_49727,N_49077);
xor UO_3117 (O_3117,N_49695,N_49391);
nor UO_3118 (O_3118,N_49378,N_49985);
nor UO_3119 (O_3119,N_49305,N_49493);
and UO_3120 (O_3120,N_49420,N_49573);
xnor UO_3121 (O_3121,N_49262,N_49272);
nor UO_3122 (O_3122,N_49802,N_49244);
nor UO_3123 (O_3123,N_49423,N_49694);
and UO_3124 (O_3124,N_49612,N_49677);
or UO_3125 (O_3125,N_49710,N_49587);
and UO_3126 (O_3126,N_49472,N_49412);
and UO_3127 (O_3127,N_49583,N_49476);
nand UO_3128 (O_3128,N_49911,N_49746);
nand UO_3129 (O_3129,N_49973,N_49771);
and UO_3130 (O_3130,N_49106,N_49042);
nand UO_3131 (O_3131,N_49870,N_49771);
or UO_3132 (O_3132,N_49874,N_49393);
xor UO_3133 (O_3133,N_49922,N_49200);
nand UO_3134 (O_3134,N_49295,N_49379);
nand UO_3135 (O_3135,N_49068,N_49693);
and UO_3136 (O_3136,N_49949,N_49798);
or UO_3137 (O_3137,N_49383,N_49457);
or UO_3138 (O_3138,N_49375,N_49505);
nand UO_3139 (O_3139,N_49150,N_49311);
xnor UO_3140 (O_3140,N_49484,N_49542);
or UO_3141 (O_3141,N_49597,N_49710);
nand UO_3142 (O_3142,N_49928,N_49159);
nor UO_3143 (O_3143,N_49272,N_49600);
or UO_3144 (O_3144,N_49899,N_49573);
nor UO_3145 (O_3145,N_49598,N_49946);
xor UO_3146 (O_3146,N_49811,N_49625);
xnor UO_3147 (O_3147,N_49299,N_49003);
nor UO_3148 (O_3148,N_49868,N_49939);
xor UO_3149 (O_3149,N_49551,N_49215);
xor UO_3150 (O_3150,N_49160,N_49506);
nor UO_3151 (O_3151,N_49724,N_49671);
or UO_3152 (O_3152,N_49724,N_49393);
nor UO_3153 (O_3153,N_49812,N_49796);
xnor UO_3154 (O_3154,N_49061,N_49902);
xnor UO_3155 (O_3155,N_49365,N_49723);
xnor UO_3156 (O_3156,N_49421,N_49879);
or UO_3157 (O_3157,N_49725,N_49921);
nand UO_3158 (O_3158,N_49076,N_49077);
xor UO_3159 (O_3159,N_49377,N_49148);
or UO_3160 (O_3160,N_49909,N_49839);
nor UO_3161 (O_3161,N_49407,N_49631);
or UO_3162 (O_3162,N_49805,N_49687);
xnor UO_3163 (O_3163,N_49258,N_49646);
xor UO_3164 (O_3164,N_49014,N_49967);
and UO_3165 (O_3165,N_49419,N_49515);
or UO_3166 (O_3166,N_49835,N_49741);
or UO_3167 (O_3167,N_49752,N_49519);
nor UO_3168 (O_3168,N_49031,N_49707);
and UO_3169 (O_3169,N_49338,N_49943);
or UO_3170 (O_3170,N_49047,N_49469);
nand UO_3171 (O_3171,N_49439,N_49238);
xnor UO_3172 (O_3172,N_49801,N_49901);
nor UO_3173 (O_3173,N_49989,N_49258);
nand UO_3174 (O_3174,N_49353,N_49200);
nor UO_3175 (O_3175,N_49538,N_49790);
nand UO_3176 (O_3176,N_49911,N_49326);
nand UO_3177 (O_3177,N_49999,N_49895);
xnor UO_3178 (O_3178,N_49114,N_49404);
nor UO_3179 (O_3179,N_49945,N_49640);
or UO_3180 (O_3180,N_49638,N_49699);
or UO_3181 (O_3181,N_49762,N_49196);
and UO_3182 (O_3182,N_49741,N_49492);
xnor UO_3183 (O_3183,N_49010,N_49996);
nor UO_3184 (O_3184,N_49974,N_49880);
nand UO_3185 (O_3185,N_49348,N_49121);
or UO_3186 (O_3186,N_49737,N_49119);
nand UO_3187 (O_3187,N_49601,N_49355);
nor UO_3188 (O_3188,N_49465,N_49910);
nor UO_3189 (O_3189,N_49927,N_49011);
and UO_3190 (O_3190,N_49239,N_49974);
and UO_3191 (O_3191,N_49434,N_49903);
or UO_3192 (O_3192,N_49036,N_49606);
nor UO_3193 (O_3193,N_49062,N_49857);
and UO_3194 (O_3194,N_49102,N_49242);
nor UO_3195 (O_3195,N_49940,N_49508);
nor UO_3196 (O_3196,N_49401,N_49269);
or UO_3197 (O_3197,N_49732,N_49313);
nand UO_3198 (O_3198,N_49029,N_49396);
xor UO_3199 (O_3199,N_49511,N_49024);
nand UO_3200 (O_3200,N_49870,N_49671);
nor UO_3201 (O_3201,N_49475,N_49405);
and UO_3202 (O_3202,N_49961,N_49306);
and UO_3203 (O_3203,N_49972,N_49778);
nand UO_3204 (O_3204,N_49843,N_49689);
and UO_3205 (O_3205,N_49318,N_49255);
nor UO_3206 (O_3206,N_49547,N_49612);
or UO_3207 (O_3207,N_49398,N_49593);
or UO_3208 (O_3208,N_49795,N_49065);
nand UO_3209 (O_3209,N_49137,N_49156);
xnor UO_3210 (O_3210,N_49651,N_49661);
xnor UO_3211 (O_3211,N_49284,N_49491);
and UO_3212 (O_3212,N_49698,N_49222);
and UO_3213 (O_3213,N_49877,N_49478);
xor UO_3214 (O_3214,N_49422,N_49245);
nand UO_3215 (O_3215,N_49162,N_49156);
nor UO_3216 (O_3216,N_49172,N_49560);
and UO_3217 (O_3217,N_49017,N_49118);
nand UO_3218 (O_3218,N_49023,N_49051);
or UO_3219 (O_3219,N_49103,N_49173);
nand UO_3220 (O_3220,N_49572,N_49492);
nand UO_3221 (O_3221,N_49802,N_49258);
and UO_3222 (O_3222,N_49639,N_49673);
nand UO_3223 (O_3223,N_49004,N_49040);
nand UO_3224 (O_3224,N_49922,N_49097);
xnor UO_3225 (O_3225,N_49629,N_49852);
and UO_3226 (O_3226,N_49051,N_49845);
xnor UO_3227 (O_3227,N_49504,N_49926);
nor UO_3228 (O_3228,N_49350,N_49319);
nor UO_3229 (O_3229,N_49093,N_49629);
or UO_3230 (O_3230,N_49102,N_49381);
or UO_3231 (O_3231,N_49509,N_49764);
nand UO_3232 (O_3232,N_49557,N_49693);
xnor UO_3233 (O_3233,N_49513,N_49742);
or UO_3234 (O_3234,N_49137,N_49604);
xnor UO_3235 (O_3235,N_49572,N_49496);
xor UO_3236 (O_3236,N_49201,N_49747);
or UO_3237 (O_3237,N_49840,N_49206);
xnor UO_3238 (O_3238,N_49125,N_49192);
xnor UO_3239 (O_3239,N_49074,N_49823);
and UO_3240 (O_3240,N_49757,N_49412);
and UO_3241 (O_3241,N_49223,N_49144);
or UO_3242 (O_3242,N_49924,N_49520);
xnor UO_3243 (O_3243,N_49965,N_49577);
nand UO_3244 (O_3244,N_49211,N_49262);
or UO_3245 (O_3245,N_49716,N_49474);
nand UO_3246 (O_3246,N_49226,N_49786);
and UO_3247 (O_3247,N_49213,N_49253);
or UO_3248 (O_3248,N_49534,N_49705);
or UO_3249 (O_3249,N_49139,N_49090);
nor UO_3250 (O_3250,N_49899,N_49544);
nand UO_3251 (O_3251,N_49905,N_49666);
and UO_3252 (O_3252,N_49126,N_49930);
nor UO_3253 (O_3253,N_49999,N_49127);
nor UO_3254 (O_3254,N_49256,N_49860);
xnor UO_3255 (O_3255,N_49791,N_49471);
and UO_3256 (O_3256,N_49924,N_49158);
and UO_3257 (O_3257,N_49971,N_49992);
or UO_3258 (O_3258,N_49573,N_49770);
nor UO_3259 (O_3259,N_49000,N_49678);
or UO_3260 (O_3260,N_49349,N_49758);
or UO_3261 (O_3261,N_49812,N_49911);
xnor UO_3262 (O_3262,N_49805,N_49065);
nor UO_3263 (O_3263,N_49710,N_49703);
nand UO_3264 (O_3264,N_49226,N_49664);
or UO_3265 (O_3265,N_49731,N_49469);
and UO_3266 (O_3266,N_49038,N_49767);
nand UO_3267 (O_3267,N_49269,N_49172);
or UO_3268 (O_3268,N_49430,N_49732);
and UO_3269 (O_3269,N_49192,N_49498);
and UO_3270 (O_3270,N_49161,N_49785);
xnor UO_3271 (O_3271,N_49612,N_49131);
or UO_3272 (O_3272,N_49842,N_49445);
xor UO_3273 (O_3273,N_49129,N_49331);
nor UO_3274 (O_3274,N_49837,N_49509);
or UO_3275 (O_3275,N_49522,N_49556);
and UO_3276 (O_3276,N_49550,N_49378);
nand UO_3277 (O_3277,N_49437,N_49067);
and UO_3278 (O_3278,N_49383,N_49960);
and UO_3279 (O_3279,N_49991,N_49616);
or UO_3280 (O_3280,N_49470,N_49256);
nor UO_3281 (O_3281,N_49748,N_49552);
nand UO_3282 (O_3282,N_49470,N_49968);
or UO_3283 (O_3283,N_49369,N_49509);
nand UO_3284 (O_3284,N_49027,N_49940);
nor UO_3285 (O_3285,N_49492,N_49901);
or UO_3286 (O_3286,N_49208,N_49106);
nand UO_3287 (O_3287,N_49028,N_49261);
nand UO_3288 (O_3288,N_49506,N_49794);
nand UO_3289 (O_3289,N_49903,N_49072);
and UO_3290 (O_3290,N_49427,N_49266);
or UO_3291 (O_3291,N_49468,N_49907);
nor UO_3292 (O_3292,N_49512,N_49593);
nand UO_3293 (O_3293,N_49096,N_49802);
and UO_3294 (O_3294,N_49971,N_49002);
xnor UO_3295 (O_3295,N_49081,N_49222);
nand UO_3296 (O_3296,N_49420,N_49485);
nor UO_3297 (O_3297,N_49605,N_49528);
and UO_3298 (O_3298,N_49417,N_49776);
or UO_3299 (O_3299,N_49221,N_49932);
xor UO_3300 (O_3300,N_49543,N_49799);
nand UO_3301 (O_3301,N_49499,N_49386);
or UO_3302 (O_3302,N_49760,N_49610);
nand UO_3303 (O_3303,N_49406,N_49207);
or UO_3304 (O_3304,N_49605,N_49622);
nor UO_3305 (O_3305,N_49316,N_49840);
nand UO_3306 (O_3306,N_49284,N_49111);
xnor UO_3307 (O_3307,N_49602,N_49964);
nand UO_3308 (O_3308,N_49612,N_49199);
xor UO_3309 (O_3309,N_49023,N_49844);
xnor UO_3310 (O_3310,N_49512,N_49636);
nor UO_3311 (O_3311,N_49338,N_49855);
nand UO_3312 (O_3312,N_49044,N_49285);
and UO_3313 (O_3313,N_49381,N_49653);
xnor UO_3314 (O_3314,N_49291,N_49987);
xnor UO_3315 (O_3315,N_49263,N_49622);
nor UO_3316 (O_3316,N_49553,N_49750);
and UO_3317 (O_3317,N_49011,N_49180);
xor UO_3318 (O_3318,N_49530,N_49540);
or UO_3319 (O_3319,N_49776,N_49493);
nand UO_3320 (O_3320,N_49840,N_49386);
and UO_3321 (O_3321,N_49449,N_49266);
xnor UO_3322 (O_3322,N_49554,N_49719);
or UO_3323 (O_3323,N_49408,N_49049);
and UO_3324 (O_3324,N_49241,N_49025);
xor UO_3325 (O_3325,N_49934,N_49886);
nand UO_3326 (O_3326,N_49251,N_49427);
and UO_3327 (O_3327,N_49310,N_49200);
nor UO_3328 (O_3328,N_49122,N_49657);
or UO_3329 (O_3329,N_49336,N_49758);
xnor UO_3330 (O_3330,N_49921,N_49814);
xor UO_3331 (O_3331,N_49505,N_49045);
nand UO_3332 (O_3332,N_49471,N_49880);
or UO_3333 (O_3333,N_49924,N_49791);
xor UO_3334 (O_3334,N_49361,N_49851);
nand UO_3335 (O_3335,N_49265,N_49688);
or UO_3336 (O_3336,N_49676,N_49003);
nor UO_3337 (O_3337,N_49645,N_49033);
or UO_3338 (O_3338,N_49836,N_49886);
nor UO_3339 (O_3339,N_49360,N_49613);
and UO_3340 (O_3340,N_49901,N_49270);
nand UO_3341 (O_3341,N_49871,N_49414);
nor UO_3342 (O_3342,N_49502,N_49523);
nand UO_3343 (O_3343,N_49431,N_49715);
or UO_3344 (O_3344,N_49872,N_49395);
xnor UO_3345 (O_3345,N_49641,N_49058);
nand UO_3346 (O_3346,N_49598,N_49720);
nor UO_3347 (O_3347,N_49418,N_49676);
xnor UO_3348 (O_3348,N_49876,N_49412);
xor UO_3349 (O_3349,N_49619,N_49772);
xor UO_3350 (O_3350,N_49145,N_49736);
and UO_3351 (O_3351,N_49184,N_49778);
or UO_3352 (O_3352,N_49836,N_49693);
nand UO_3353 (O_3353,N_49221,N_49913);
and UO_3354 (O_3354,N_49176,N_49743);
or UO_3355 (O_3355,N_49299,N_49785);
xnor UO_3356 (O_3356,N_49342,N_49350);
nand UO_3357 (O_3357,N_49814,N_49068);
xnor UO_3358 (O_3358,N_49912,N_49894);
xnor UO_3359 (O_3359,N_49245,N_49154);
or UO_3360 (O_3360,N_49011,N_49608);
or UO_3361 (O_3361,N_49875,N_49260);
or UO_3362 (O_3362,N_49475,N_49738);
or UO_3363 (O_3363,N_49565,N_49699);
or UO_3364 (O_3364,N_49357,N_49071);
and UO_3365 (O_3365,N_49816,N_49719);
nor UO_3366 (O_3366,N_49669,N_49964);
xor UO_3367 (O_3367,N_49014,N_49160);
or UO_3368 (O_3368,N_49119,N_49540);
xnor UO_3369 (O_3369,N_49127,N_49599);
or UO_3370 (O_3370,N_49445,N_49549);
or UO_3371 (O_3371,N_49377,N_49673);
xor UO_3372 (O_3372,N_49830,N_49879);
xor UO_3373 (O_3373,N_49639,N_49871);
nand UO_3374 (O_3374,N_49264,N_49621);
and UO_3375 (O_3375,N_49054,N_49736);
xnor UO_3376 (O_3376,N_49904,N_49691);
nor UO_3377 (O_3377,N_49859,N_49532);
nor UO_3378 (O_3378,N_49285,N_49166);
nand UO_3379 (O_3379,N_49430,N_49627);
xnor UO_3380 (O_3380,N_49578,N_49743);
xor UO_3381 (O_3381,N_49063,N_49726);
nand UO_3382 (O_3382,N_49544,N_49881);
or UO_3383 (O_3383,N_49674,N_49979);
xor UO_3384 (O_3384,N_49918,N_49885);
nand UO_3385 (O_3385,N_49527,N_49674);
or UO_3386 (O_3386,N_49662,N_49968);
nor UO_3387 (O_3387,N_49597,N_49677);
and UO_3388 (O_3388,N_49761,N_49301);
nand UO_3389 (O_3389,N_49395,N_49464);
xnor UO_3390 (O_3390,N_49151,N_49455);
and UO_3391 (O_3391,N_49981,N_49952);
nor UO_3392 (O_3392,N_49895,N_49313);
nand UO_3393 (O_3393,N_49560,N_49257);
and UO_3394 (O_3394,N_49748,N_49307);
or UO_3395 (O_3395,N_49797,N_49226);
nor UO_3396 (O_3396,N_49788,N_49904);
and UO_3397 (O_3397,N_49490,N_49675);
xor UO_3398 (O_3398,N_49723,N_49924);
nor UO_3399 (O_3399,N_49258,N_49515);
xor UO_3400 (O_3400,N_49177,N_49014);
xnor UO_3401 (O_3401,N_49710,N_49147);
and UO_3402 (O_3402,N_49726,N_49423);
nor UO_3403 (O_3403,N_49973,N_49596);
nand UO_3404 (O_3404,N_49265,N_49169);
xor UO_3405 (O_3405,N_49007,N_49632);
xor UO_3406 (O_3406,N_49278,N_49513);
or UO_3407 (O_3407,N_49420,N_49816);
or UO_3408 (O_3408,N_49323,N_49201);
nand UO_3409 (O_3409,N_49743,N_49329);
or UO_3410 (O_3410,N_49359,N_49722);
or UO_3411 (O_3411,N_49009,N_49801);
nand UO_3412 (O_3412,N_49458,N_49335);
nor UO_3413 (O_3413,N_49240,N_49658);
nand UO_3414 (O_3414,N_49771,N_49636);
nand UO_3415 (O_3415,N_49970,N_49502);
nor UO_3416 (O_3416,N_49697,N_49049);
or UO_3417 (O_3417,N_49415,N_49244);
or UO_3418 (O_3418,N_49809,N_49786);
xor UO_3419 (O_3419,N_49820,N_49250);
or UO_3420 (O_3420,N_49396,N_49566);
and UO_3421 (O_3421,N_49543,N_49458);
and UO_3422 (O_3422,N_49139,N_49750);
and UO_3423 (O_3423,N_49954,N_49893);
or UO_3424 (O_3424,N_49598,N_49259);
or UO_3425 (O_3425,N_49823,N_49821);
nand UO_3426 (O_3426,N_49071,N_49329);
nor UO_3427 (O_3427,N_49617,N_49161);
and UO_3428 (O_3428,N_49618,N_49197);
and UO_3429 (O_3429,N_49709,N_49601);
or UO_3430 (O_3430,N_49109,N_49883);
nor UO_3431 (O_3431,N_49585,N_49726);
or UO_3432 (O_3432,N_49598,N_49475);
and UO_3433 (O_3433,N_49248,N_49553);
nor UO_3434 (O_3434,N_49285,N_49573);
or UO_3435 (O_3435,N_49174,N_49462);
nand UO_3436 (O_3436,N_49181,N_49265);
and UO_3437 (O_3437,N_49572,N_49177);
and UO_3438 (O_3438,N_49914,N_49741);
or UO_3439 (O_3439,N_49270,N_49994);
nand UO_3440 (O_3440,N_49070,N_49828);
or UO_3441 (O_3441,N_49259,N_49441);
and UO_3442 (O_3442,N_49827,N_49861);
xor UO_3443 (O_3443,N_49793,N_49442);
and UO_3444 (O_3444,N_49660,N_49145);
nor UO_3445 (O_3445,N_49238,N_49737);
nand UO_3446 (O_3446,N_49803,N_49542);
xnor UO_3447 (O_3447,N_49189,N_49860);
nand UO_3448 (O_3448,N_49862,N_49623);
nor UO_3449 (O_3449,N_49268,N_49382);
and UO_3450 (O_3450,N_49147,N_49033);
or UO_3451 (O_3451,N_49401,N_49760);
xnor UO_3452 (O_3452,N_49198,N_49098);
nand UO_3453 (O_3453,N_49220,N_49540);
xnor UO_3454 (O_3454,N_49877,N_49006);
or UO_3455 (O_3455,N_49893,N_49901);
nor UO_3456 (O_3456,N_49073,N_49559);
or UO_3457 (O_3457,N_49990,N_49222);
nand UO_3458 (O_3458,N_49515,N_49355);
or UO_3459 (O_3459,N_49831,N_49429);
nor UO_3460 (O_3460,N_49077,N_49127);
xnor UO_3461 (O_3461,N_49865,N_49890);
or UO_3462 (O_3462,N_49063,N_49388);
or UO_3463 (O_3463,N_49839,N_49306);
nor UO_3464 (O_3464,N_49917,N_49979);
nand UO_3465 (O_3465,N_49161,N_49884);
nand UO_3466 (O_3466,N_49649,N_49138);
or UO_3467 (O_3467,N_49536,N_49668);
xor UO_3468 (O_3468,N_49960,N_49683);
nand UO_3469 (O_3469,N_49474,N_49075);
nand UO_3470 (O_3470,N_49301,N_49500);
xnor UO_3471 (O_3471,N_49497,N_49596);
or UO_3472 (O_3472,N_49195,N_49405);
nor UO_3473 (O_3473,N_49471,N_49018);
or UO_3474 (O_3474,N_49559,N_49358);
nand UO_3475 (O_3475,N_49195,N_49317);
nor UO_3476 (O_3476,N_49368,N_49716);
nand UO_3477 (O_3477,N_49693,N_49690);
and UO_3478 (O_3478,N_49778,N_49746);
xor UO_3479 (O_3479,N_49990,N_49646);
or UO_3480 (O_3480,N_49342,N_49071);
and UO_3481 (O_3481,N_49639,N_49615);
or UO_3482 (O_3482,N_49204,N_49513);
and UO_3483 (O_3483,N_49471,N_49732);
xnor UO_3484 (O_3484,N_49537,N_49348);
or UO_3485 (O_3485,N_49155,N_49397);
or UO_3486 (O_3486,N_49378,N_49332);
and UO_3487 (O_3487,N_49841,N_49962);
nand UO_3488 (O_3488,N_49191,N_49553);
and UO_3489 (O_3489,N_49904,N_49042);
or UO_3490 (O_3490,N_49637,N_49788);
and UO_3491 (O_3491,N_49071,N_49827);
and UO_3492 (O_3492,N_49709,N_49581);
nor UO_3493 (O_3493,N_49442,N_49487);
xnor UO_3494 (O_3494,N_49075,N_49564);
and UO_3495 (O_3495,N_49468,N_49356);
nand UO_3496 (O_3496,N_49938,N_49176);
and UO_3497 (O_3497,N_49836,N_49229);
nand UO_3498 (O_3498,N_49524,N_49848);
nand UO_3499 (O_3499,N_49203,N_49837);
or UO_3500 (O_3500,N_49517,N_49285);
or UO_3501 (O_3501,N_49062,N_49534);
nor UO_3502 (O_3502,N_49559,N_49018);
and UO_3503 (O_3503,N_49909,N_49997);
nand UO_3504 (O_3504,N_49458,N_49447);
nand UO_3505 (O_3505,N_49165,N_49569);
nand UO_3506 (O_3506,N_49896,N_49439);
or UO_3507 (O_3507,N_49451,N_49231);
nand UO_3508 (O_3508,N_49394,N_49568);
and UO_3509 (O_3509,N_49348,N_49632);
and UO_3510 (O_3510,N_49397,N_49307);
or UO_3511 (O_3511,N_49791,N_49535);
and UO_3512 (O_3512,N_49105,N_49529);
nor UO_3513 (O_3513,N_49088,N_49587);
nand UO_3514 (O_3514,N_49846,N_49693);
and UO_3515 (O_3515,N_49787,N_49691);
and UO_3516 (O_3516,N_49798,N_49287);
and UO_3517 (O_3517,N_49337,N_49270);
nand UO_3518 (O_3518,N_49540,N_49934);
xnor UO_3519 (O_3519,N_49087,N_49275);
nand UO_3520 (O_3520,N_49329,N_49742);
nand UO_3521 (O_3521,N_49158,N_49145);
nand UO_3522 (O_3522,N_49216,N_49655);
xor UO_3523 (O_3523,N_49411,N_49477);
or UO_3524 (O_3524,N_49955,N_49941);
nand UO_3525 (O_3525,N_49874,N_49183);
nand UO_3526 (O_3526,N_49904,N_49575);
and UO_3527 (O_3527,N_49372,N_49419);
nor UO_3528 (O_3528,N_49397,N_49329);
nor UO_3529 (O_3529,N_49307,N_49704);
nor UO_3530 (O_3530,N_49598,N_49457);
nand UO_3531 (O_3531,N_49221,N_49335);
xor UO_3532 (O_3532,N_49086,N_49561);
and UO_3533 (O_3533,N_49832,N_49979);
nor UO_3534 (O_3534,N_49791,N_49114);
nand UO_3535 (O_3535,N_49255,N_49605);
xnor UO_3536 (O_3536,N_49113,N_49800);
or UO_3537 (O_3537,N_49036,N_49006);
or UO_3538 (O_3538,N_49872,N_49956);
nand UO_3539 (O_3539,N_49199,N_49145);
nand UO_3540 (O_3540,N_49096,N_49085);
nor UO_3541 (O_3541,N_49721,N_49229);
and UO_3542 (O_3542,N_49693,N_49967);
nand UO_3543 (O_3543,N_49518,N_49866);
nor UO_3544 (O_3544,N_49830,N_49675);
xnor UO_3545 (O_3545,N_49557,N_49488);
nor UO_3546 (O_3546,N_49924,N_49601);
nand UO_3547 (O_3547,N_49989,N_49085);
or UO_3548 (O_3548,N_49279,N_49394);
or UO_3549 (O_3549,N_49909,N_49272);
nor UO_3550 (O_3550,N_49498,N_49490);
or UO_3551 (O_3551,N_49695,N_49733);
nand UO_3552 (O_3552,N_49767,N_49396);
xor UO_3553 (O_3553,N_49001,N_49175);
or UO_3554 (O_3554,N_49172,N_49786);
nand UO_3555 (O_3555,N_49837,N_49213);
nor UO_3556 (O_3556,N_49901,N_49774);
and UO_3557 (O_3557,N_49248,N_49849);
and UO_3558 (O_3558,N_49286,N_49313);
nand UO_3559 (O_3559,N_49644,N_49319);
nor UO_3560 (O_3560,N_49985,N_49576);
nor UO_3561 (O_3561,N_49859,N_49890);
and UO_3562 (O_3562,N_49831,N_49182);
nand UO_3563 (O_3563,N_49919,N_49964);
nor UO_3564 (O_3564,N_49089,N_49910);
nand UO_3565 (O_3565,N_49037,N_49061);
xor UO_3566 (O_3566,N_49682,N_49411);
and UO_3567 (O_3567,N_49233,N_49228);
nand UO_3568 (O_3568,N_49601,N_49506);
or UO_3569 (O_3569,N_49114,N_49842);
nor UO_3570 (O_3570,N_49073,N_49646);
and UO_3571 (O_3571,N_49253,N_49695);
xor UO_3572 (O_3572,N_49848,N_49533);
nand UO_3573 (O_3573,N_49051,N_49474);
nand UO_3574 (O_3574,N_49340,N_49811);
and UO_3575 (O_3575,N_49809,N_49194);
and UO_3576 (O_3576,N_49394,N_49377);
or UO_3577 (O_3577,N_49224,N_49633);
nor UO_3578 (O_3578,N_49247,N_49568);
nand UO_3579 (O_3579,N_49136,N_49976);
nand UO_3580 (O_3580,N_49454,N_49024);
and UO_3581 (O_3581,N_49579,N_49612);
xnor UO_3582 (O_3582,N_49355,N_49811);
nor UO_3583 (O_3583,N_49800,N_49043);
and UO_3584 (O_3584,N_49780,N_49822);
nor UO_3585 (O_3585,N_49059,N_49872);
nand UO_3586 (O_3586,N_49244,N_49595);
xor UO_3587 (O_3587,N_49550,N_49968);
and UO_3588 (O_3588,N_49545,N_49795);
xnor UO_3589 (O_3589,N_49064,N_49035);
nand UO_3590 (O_3590,N_49755,N_49636);
nor UO_3591 (O_3591,N_49971,N_49429);
and UO_3592 (O_3592,N_49453,N_49936);
nand UO_3593 (O_3593,N_49585,N_49969);
nor UO_3594 (O_3594,N_49950,N_49094);
and UO_3595 (O_3595,N_49922,N_49691);
xor UO_3596 (O_3596,N_49468,N_49895);
or UO_3597 (O_3597,N_49299,N_49676);
xor UO_3598 (O_3598,N_49963,N_49351);
and UO_3599 (O_3599,N_49491,N_49930);
xnor UO_3600 (O_3600,N_49876,N_49836);
or UO_3601 (O_3601,N_49910,N_49496);
xor UO_3602 (O_3602,N_49632,N_49364);
nor UO_3603 (O_3603,N_49083,N_49863);
xnor UO_3604 (O_3604,N_49804,N_49898);
and UO_3605 (O_3605,N_49949,N_49546);
nand UO_3606 (O_3606,N_49071,N_49197);
nand UO_3607 (O_3607,N_49632,N_49965);
and UO_3608 (O_3608,N_49389,N_49893);
and UO_3609 (O_3609,N_49803,N_49409);
or UO_3610 (O_3610,N_49040,N_49808);
nor UO_3611 (O_3611,N_49217,N_49580);
or UO_3612 (O_3612,N_49481,N_49542);
or UO_3613 (O_3613,N_49832,N_49271);
or UO_3614 (O_3614,N_49674,N_49848);
and UO_3615 (O_3615,N_49831,N_49413);
nor UO_3616 (O_3616,N_49383,N_49881);
nor UO_3617 (O_3617,N_49770,N_49380);
nor UO_3618 (O_3618,N_49545,N_49168);
and UO_3619 (O_3619,N_49214,N_49926);
nor UO_3620 (O_3620,N_49767,N_49830);
and UO_3621 (O_3621,N_49796,N_49126);
and UO_3622 (O_3622,N_49084,N_49057);
xnor UO_3623 (O_3623,N_49971,N_49994);
xor UO_3624 (O_3624,N_49735,N_49954);
and UO_3625 (O_3625,N_49827,N_49531);
and UO_3626 (O_3626,N_49548,N_49243);
xnor UO_3627 (O_3627,N_49569,N_49598);
nand UO_3628 (O_3628,N_49811,N_49279);
and UO_3629 (O_3629,N_49776,N_49914);
nor UO_3630 (O_3630,N_49773,N_49772);
or UO_3631 (O_3631,N_49356,N_49956);
nor UO_3632 (O_3632,N_49050,N_49202);
nor UO_3633 (O_3633,N_49152,N_49361);
nand UO_3634 (O_3634,N_49250,N_49311);
xor UO_3635 (O_3635,N_49457,N_49910);
xnor UO_3636 (O_3636,N_49294,N_49360);
nor UO_3637 (O_3637,N_49540,N_49721);
nand UO_3638 (O_3638,N_49346,N_49665);
nand UO_3639 (O_3639,N_49022,N_49609);
nor UO_3640 (O_3640,N_49869,N_49853);
and UO_3641 (O_3641,N_49053,N_49699);
or UO_3642 (O_3642,N_49976,N_49417);
and UO_3643 (O_3643,N_49004,N_49177);
or UO_3644 (O_3644,N_49168,N_49872);
or UO_3645 (O_3645,N_49925,N_49719);
nand UO_3646 (O_3646,N_49408,N_49343);
and UO_3647 (O_3647,N_49578,N_49186);
xnor UO_3648 (O_3648,N_49150,N_49232);
xnor UO_3649 (O_3649,N_49251,N_49363);
and UO_3650 (O_3650,N_49457,N_49169);
or UO_3651 (O_3651,N_49071,N_49454);
xor UO_3652 (O_3652,N_49595,N_49825);
or UO_3653 (O_3653,N_49994,N_49779);
nor UO_3654 (O_3654,N_49272,N_49819);
or UO_3655 (O_3655,N_49722,N_49934);
xor UO_3656 (O_3656,N_49980,N_49506);
or UO_3657 (O_3657,N_49638,N_49734);
xor UO_3658 (O_3658,N_49767,N_49466);
nor UO_3659 (O_3659,N_49074,N_49742);
or UO_3660 (O_3660,N_49328,N_49849);
nand UO_3661 (O_3661,N_49490,N_49485);
or UO_3662 (O_3662,N_49779,N_49235);
nor UO_3663 (O_3663,N_49142,N_49999);
nor UO_3664 (O_3664,N_49084,N_49119);
nand UO_3665 (O_3665,N_49231,N_49056);
xor UO_3666 (O_3666,N_49952,N_49900);
xor UO_3667 (O_3667,N_49885,N_49836);
and UO_3668 (O_3668,N_49072,N_49358);
xor UO_3669 (O_3669,N_49555,N_49605);
nor UO_3670 (O_3670,N_49964,N_49508);
nor UO_3671 (O_3671,N_49286,N_49648);
and UO_3672 (O_3672,N_49773,N_49726);
and UO_3673 (O_3673,N_49263,N_49982);
or UO_3674 (O_3674,N_49556,N_49071);
and UO_3675 (O_3675,N_49299,N_49571);
nand UO_3676 (O_3676,N_49720,N_49904);
nor UO_3677 (O_3677,N_49427,N_49714);
nand UO_3678 (O_3678,N_49766,N_49927);
xor UO_3679 (O_3679,N_49619,N_49908);
and UO_3680 (O_3680,N_49887,N_49583);
and UO_3681 (O_3681,N_49731,N_49542);
xnor UO_3682 (O_3682,N_49749,N_49636);
or UO_3683 (O_3683,N_49147,N_49848);
xnor UO_3684 (O_3684,N_49431,N_49584);
nor UO_3685 (O_3685,N_49722,N_49981);
and UO_3686 (O_3686,N_49790,N_49578);
and UO_3687 (O_3687,N_49763,N_49914);
and UO_3688 (O_3688,N_49777,N_49423);
or UO_3689 (O_3689,N_49169,N_49069);
or UO_3690 (O_3690,N_49502,N_49400);
nand UO_3691 (O_3691,N_49390,N_49405);
xor UO_3692 (O_3692,N_49671,N_49331);
nor UO_3693 (O_3693,N_49122,N_49049);
or UO_3694 (O_3694,N_49801,N_49625);
and UO_3695 (O_3695,N_49931,N_49527);
xnor UO_3696 (O_3696,N_49154,N_49345);
or UO_3697 (O_3697,N_49742,N_49581);
nand UO_3698 (O_3698,N_49887,N_49461);
xnor UO_3699 (O_3699,N_49893,N_49335);
or UO_3700 (O_3700,N_49691,N_49566);
xnor UO_3701 (O_3701,N_49826,N_49698);
xnor UO_3702 (O_3702,N_49824,N_49598);
nand UO_3703 (O_3703,N_49541,N_49037);
or UO_3704 (O_3704,N_49552,N_49014);
or UO_3705 (O_3705,N_49488,N_49116);
nor UO_3706 (O_3706,N_49507,N_49121);
nor UO_3707 (O_3707,N_49010,N_49392);
xnor UO_3708 (O_3708,N_49038,N_49584);
nand UO_3709 (O_3709,N_49960,N_49268);
nand UO_3710 (O_3710,N_49551,N_49131);
xor UO_3711 (O_3711,N_49854,N_49199);
nand UO_3712 (O_3712,N_49339,N_49714);
and UO_3713 (O_3713,N_49780,N_49779);
nor UO_3714 (O_3714,N_49203,N_49420);
xor UO_3715 (O_3715,N_49483,N_49071);
xnor UO_3716 (O_3716,N_49228,N_49286);
or UO_3717 (O_3717,N_49307,N_49440);
xnor UO_3718 (O_3718,N_49056,N_49297);
nand UO_3719 (O_3719,N_49838,N_49934);
or UO_3720 (O_3720,N_49744,N_49681);
xnor UO_3721 (O_3721,N_49589,N_49536);
or UO_3722 (O_3722,N_49478,N_49926);
xnor UO_3723 (O_3723,N_49674,N_49167);
xor UO_3724 (O_3724,N_49097,N_49470);
nor UO_3725 (O_3725,N_49811,N_49408);
nand UO_3726 (O_3726,N_49417,N_49718);
or UO_3727 (O_3727,N_49905,N_49465);
or UO_3728 (O_3728,N_49155,N_49498);
nor UO_3729 (O_3729,N_49238,N_49331);
nand UO_3730 (O_3730,N_49950,N_49070);
or UO_3731 (O_3731,N_49850,N_49762);
or UO_3732 (O_3732,N_49387,N_49645);
nor UO_3733 (O_3733,N_49558,N_49194);
and UO_3734 (O_3734,N_49352,N_49967);
nor UO_3735 (O_3735,N_49494,N_49948);
xnor UO_3736 (O_3736,N_49193,N_49789);
nor UO_3737 (O_3737,N_49704,N_49231);
and UO_3738 (O_3738,N_49976,N_49342);
xor UO_3739 (O_3739,N_49817,N_49920);
nor UO_3740 (O_3740,N_49451,N_49780);
or UO_3741 (O_3741,N_49207,N_49561);
nor UO_3742 (O_3742,N_49720,N_49614);
nand UO_3743 (O_3743,N_49069,N_49621);
nor UO_3744 (O_3744,N_49193,N_49438);
and UO_3745 (O_3745,N_49431,N_49350);
xor UO_3746 (O_3746,N_49709,N_49489);
or UO_3747 (O_3747,N_49247,N_49780);
xnor UO_3748 (O_3748,N_49012,N_49301);
nand UO_3749 (O_3749,N_49476,N_49529);
nor UO_3750 (O_3750,N_49355,N_49737);
nor UO_3751 (O_3751,N_49615,N_49917);
and UO_3752 (O_3752,N_49845,N_49001);
nor UO_3753 (O_3753,N_49650,N_49379);
nand UO_3754 (O_3754,N_49304,N_49066);
nand UO_3755 (O_3755,N_49969,N_49771);
or UO_3756 (O_3756,N_49098,N_49618);
xnor UO_3757 (O_3757,N_49704,N_49312);
nor UO_3758 (O_3758,N_49566,N_49569);
nand UO_3759 (O_3759,N_49871,N_49236);
and UO_3760 (O_3760,N_49995,N_49728);
or UO_3761 (O_3761,N_49228,N_49276);
nand UO_3762 (O_3762,N_49395,N_49933);
or UO_3763 (O_3763,N_49419,N_49873);
and UO_3764 (O_3764,N_49702,N_49117);
nor UO_3765 (O_3765,N_49693,N_49827);
xor UO_3766 (O_3766,N_49018,N_49454);
xor UO_3767 (O_3767,N_49723,N_49309);
xnor UO_3768 (O_3768,N_49900,N_49310);
nand UO_3769 (O_3769,N_49434,N_49768);
nand UO_3770 (O_3770,N_49743,N_49434);
and UO_3771 (O_3771,N_49616,N_49368);
and UO_3772 (O_3772,N_49484,N_49241);
nor UO_3773 (O_3773,N_49455,N_49023);
and UO_3774 (O_3774,N_49490,N_49564);
nor UO_3775 (O_3775,N_49940,N_49548);
or UO_3776 (O_3776,N_49337,N_49384);
xor UO_3777 (O_3777,N_49428,N_49688);
or UO_3778 (O_3778,N_49519,N_49214);
nor UO_3779 (O_3779,N_49559,N_49873);
xnor UO_3780 (O_3780,N_49517,N_49238);
nand UO_3781 (O_3781,N_49826,N_49571);
and UO_3782 (O_3782,N_49587,N_49571);
or UO_3783 (O_3783,N_49897,N_49380);
xnor UO_3784 (O_3784,N_49413,N_49971);
and UO_3785 (O_3785,N_49786,N_49587);
xnor UO_3786 (O_3786,N_49042,N_49579);
and UO_3787 (O_3787,N_49930,N_49236);
or UO_3788 (O_3788,N_49693,N_49583);
xor UO_3789 (O_3789,N_49002,N_49793);
nand UO_3790 (O_3790,N_49466,N_49658);
nor UO_3791 (O_3791,N_49079,N_49451);
xor UO_3792 (O_3792,N_49540,N_49634);
and UO_3793 (O_3793,N_49578,N_49113);
nand UO_3794 (O_3794,N_49525,N_49269);
or UO_3795 (O_3795,N_49545,N_49732);
xnor UO_3796 (O_3796,N_49856,N_49762);
nor UO_3797 (O_3797,N_49583,N_49370);
or UO_3798 (O_3798,N_49363,N_49240);
and UO_3799 (O_3799,N_49028,N_49806);
xor UO_3800 (O_3800,N_49875,N_49048);
nor UO_3801 (O_3801,N_49595,N_49815);
nand UO_3802 (O_3802,N_49738,N_49416);
nor UO_3803 (O_3803,N_49412,N_49056);
xnor UO_3804 (O_3804,N_49634,N_49609);
nor UO_3805 (O_3805,N_49976,N_49589);
nand UO_3806 (O_3806,N_49271,N_49055);
nor UO_3807 (O_3807,N_49233,N_49880);
nor UO_3808 (O_3808,N_49242,N_49098);
and UO_3809 (O_3809,N_49721,N_49974);
xor UO_3810 (O_3810,N_49260,N_49831);
nor UO_3811 (O_3811,N_49544,N_49826);
nand UO_3812 (O_3812,N_49146,N_49262);
xor UO_3813 (O_3813,N_49589,N_49443);
and UO_3814 (O_3814,N_49405,N_49626);
or UO_3815 (O_3815,N_49792,N_49585);
nand UO_3816 (O_3816,N_49432,N_49698);
nand UO_3817 (O_3817,N_49514,N_49674);
nor UO_3818 (O_3818,N_49115,N_49125);
xnor UO_3819 (O_3819,N_49593,N_49858);
xor UO_3820 (O_3820,N_49009,N_49271);
nand UO_3821 (O_3821,N_49070,N_49203);
and UO_3822 (O_3822,N_49526,N_49327);
nand UO_3823 (O_3823,N_49690,N_49458);
or UO_3824 (O_3824,N_49723,N_49194);
or UO_3825 (O_3825,N_49537,N_49985);
xor UO_3826 (O_3826,N_49183,N_49763);
or UO_3827 (O_3827,N_49583,N_49849);
nand UO_3828 (O_3828,N_49514,N_49570);
nand UO_3829 (O_3829,N_49061,N_49793);
xor UO_3830 (O_3830,N_49689,N_49991);
and UO_3831 (O_3831,N_49429,N_49579);
nor UO_3832 (O_3832,N_49829,N_49933);
and UO_3833 (O_3833,N_49305,N_49189);
nand UO_3834 (O_3834,N_49166,N_49471);
nor UO_3835 (O_3835,N_49559,N_49369);
nor UO_3836 (O_3836,N_49758,N_49814);
xnor UO_3837 (O_3837,N_49663,N_49159);
nor UO_3838 (O_3838,N_49328,N_49063);
or UO_3839 (O_3839,N_49947,N_49732);
xnor UO_3840 (O_3840,N_49717,N_49945);
nor UO_3841 (O_3841,N_49889,N_49733);
xnor UO_3842 (O_3842,N_49107,N_49129);
nor UO_3843 (O_3843,N_49514,N_49101);
and UO_3844 (O_3844,N_49582,N_49630);
or UO_3845 (O_3845,N_49839,N_49979);
and UO_3846 (O_3846,N_49077,N_49057);
nand UO_3847 (O_3847,N_49390,N_49384);
or UO_3848 (O_3848,N_49888,N_49628);
or UO_3849 (O_3849,N_49319,N_49089);
nand UO_3850 (O_3850,N_49142,N_49210);
and UO_3851 (O_3851,N_49704,N_49050);
nand UO_3852 (O_3852,N_49041,N_49323);
nand UO_3853 (O_3853,N_49951,N_49801);
or UO_3854 (O_3854,N_49626,N_49298);
xnor UO_3855 (O_3855,N_49314,N_49681);
and UO_3856 (O_3856,N_49420,N_49224);
or UO_3857 (O_3857,N_49919,N_49179);
xnor UO_3858 (O_3858,N_49696,N_49557);
and UO_3859 (O_3859,N_49922,N_49261);
or UO_3860 (O_3860,N_49623,N_49541);
and UO_3861 (O_3861,N_49455,N_49327);
nand UO_3862 (O_3862,N_49708,N_49686);
or UO_3863 (O_3863,N_49518,N_49512);
and UO_3864 (O_3864,N_49572,N_49347);
and UO_3865 (O_3865,N_49967,N_49479);
nand UO_3866 (O_3866,N_49758,N_49726);
nand UO_3867 (O_3867,N_49855,N_49960);
nor UO_3868 (O_3868,N_49670,N_49960);
nor UO_3869 (O_3869,N_49523,N_49794);
or UO_3870 (O_3870,N_49523,N_49859);
nand UO_3871 (O_3871,N_49711,N_49835);
nand UO_3872 (O_3872,N_49781,N_49301);
or UO_3873 (O_3873,N_49056,N_49271);
nand UO_3874 (O_3874,N_49238,N_49786);
or UO_3875 (O_3875,N_49665,N_49364);
xor UO_3876 (O_3876,N_49227,N_49493);
or UO_3877 (O_3877,N_49822,N_49884);
and UO_3878 (O_3878,N_49976,N_49897);
or UO_3879 (O_3879,N_49485,N_49103);
or UO_3880 (O_3880,N_49920,N_49803);
nand UO_3881 (O_3881,N_49714,N_49167);
or UO_3882 (O_3882,N_49173,N_49608);
xnor UO_3883 (O_3883,N_49363,N_49605);
and UO_3884 (O_3884,N_49999,N_49073);
nor UO_3885 (O_3885,N_49161,N_49114);
xnor UO_3886 (O_3886,N_49555,N_49513);
xnor UO_3887 (O_3887,N_49551,N_49372);
or UO_3888 (O_3888,N_49456,N_49178);
xor UO_3889 (O_3889,N_49857,N_49177);
xnor UO_3890 (O_3890,N_49946,N_49980);
and UO_3891 (O_3891,N_49141,N_49176);
nor UO_3892 (O_3892,N_49447,N_49455);
xnor UO_3893 (O_3893,N_49815,N_49024);
or UO_3894 (O_3894,N_49715,N_49371);
and UO_3895 (O_3895,N_49528,N_49783);
and UO_3896 (O_3896,N_49680,N_49632);
xnor UO_3897 (O_3897,N_49261,N_49174);
and UO_3898 (O_3898,N_49883,N_49523);
nand UO_3899 (O_3899,N_49832,N_49265);
nor UO_3900 (O_3900,N_49952,N_49644);
and UO_3901 (O_3901,N_49950,N_49060);
xnor UO_3902 (O_3902,N_49425,N_49061);
nand UO_3903 (O_3903,N_49240,N_49494);
nor UO_3904 (O_3904,N_49095,N_49469);
nor UO_3905 (O_3905,N_49759,N_49225);
or UO_3906 (O_3906,N_49809,N_49327);
nor UO_3907 (O_3907,N_49525,N_49160);
nor UO_3908 (O_3908,N_49746,N_49359);
xnor UO_3909 (O_3909,N_49781,N_49126);
xnor UO_3910 (O_3910,N_49639,N_49710);
and UO_3911 (O_3911,N_49250,N_49017);
nand UO_3912 (O_3912,N_49093,N_49366);
nand UO_3913 (O_3913,N_49683,N_49408);
and UO_3914 (O_3914,N_49932,N_49442);
or UO_3915 (O_3915,N_49860,N_49563);
xor UO_3916 (O_3916,N_49453,N_49305);
or UO_3917 (O_3917,N_49164,N_49764);
nand UO_3918 (O_3918,N_49445,N_49393);
nand UO_3919 (O_3919,N_49381,N_49828);
nor UO_3920 (O_3920,N_49465,N_49010);
xnor UO_3921 (O_3921,N_49087,N_49762);
nor UO_3922 (O_3922,N_49640,N_49237);
nand UO_3923 (O_3923,N_49792,N_49026);
nand UO_3924 (O_3924,N_49605,N_49967);
nor UO_3925 (O_3925,N_49969,N_49529);
and UO_3926 (O_3926,N_49660,N_49482);
xor UO_3927 (O_3927,N_49823,N_49004);
and UO_3928 (O_3928,N_49101,N_49474);
or UO_3929 (O_3929,N_49107,N_49578);
nor UO_3930 (O_3930,N_49103,N_49254);
and UO_3931 (O_3931,N_49210,N_49766);
nor UO_3932 (O_3932,N_49476,N_49642);
and UO_3933 (O_3933,N_49401,N_49135);
nand UO_3934 (O_3934,N_49519,N_49528);
nor UO_3935 (O_3935,N_49816,N_49409);
and UO_3936 (O_3936,N_49371,N_49012);
nand UO_3937 (O_3937,N_49979,N_49829);
xor UO_3938 (O_3938,N_49866,N_49730);
and UO_3939 (O_3939,N_49153,N_49202);
nand UO_3940 (O_3940,N_49897,N_49693);
nor UO_3941 (O_3941,N_49392,N_49618);
nand UO_3942 (O_3942,N_49335,N_49887);
xor UO_3943 (O_3943,N_49794,N_49745);
xnor UO_3944 (O_3944,N_49945,N_49558);
or UO_3945 (O_3945,N_49209,N_49958);
and UO_3946 (O_3946,N_49595,N_49411);
and UO_3947 (O_3947,N_49853,N_49777);
xnor UO_3948 (O_3948,N_49571,N_49244);
xnor UO_3949 (O_3949,N_49480,N_49721);
xnor UO_3950 (O_3950,N_49818,N_49258);
nand UO_3951 (O_3951,N_49262,N_49507);
nand UO_3952 (O_3952,N_49574,N_49557);
nor UO_3953 (O_3953,N_49561,N_49066);
nand UO_3954 (O_3954,N_49605,N_49001);
nor UO_3955 (O_3955,N_49177,N_49385);
or UO_3956 (O_3956,N_49721,N_49340);
or UO_3957 (O_3957,N_49420,N_49980);
nand UO_3958 (O_3958,N_49203,N_49533);
xnor UO_3959 (O_3959,N_49488,N_49102);
and UO_3960 (O_3960,N_49455,N_49677);
nor UO_3961 (O_3961,N_49281,N_49850);
nor UO_3962 (O_3962,N_49549,N_49244);
and UO_3963 (O_3963,N_49770,N_49482);
and UO_3964 (O_3964,N_49845,N_49898);
nand UO_3965 (O_3965,N_49886,N_49007);
and UO_3966 (O_3966,N_49911,N_49831);
nor UO_3967 (O_3967,N_49951,N_49898);
xnor UO_3968 (O_3968,N_49919,N_49278);
xor UO_3969 (O_3969,N_49545,N_49584);
nor UO_3970 (O_3970,N_49602,N_49654);
xnor UO_3971 (O_3971,N_49167,N_49733);
and UO_3972 (O_3972,N_49214,N_49614);
nor UO_3973 (O_3973,N_49781,N_49293);
xnor UO_3974 (O_3974,N_49662,N_49476);
nand UO_3975 (O_3975,N_49968,N_49167);
xor UO_3976 (O_3976,N_49155,N_49114);
nand UO_3977 (O_3977,N_49945,N_49871);
or UO_3978 (O_3978,N_49716,N_49882);
nor UO_3979 (O_3979,N_49848,N_49521);
and UO_3980 (O_3980,N_49925,N_49613);
nand UO_3981 (O_3981,N_49377,N_49536);
xnor UO_3982 (O_3982,N_49267,N_49397);
and UO_3983 (O_3983,N_49302,N_49156);
xnor UO_3984 (O_3984,N_49740,N_49644);
nor UO_3985 (O_3985,N_49294,N_49199);
or UO_3986 (O_3986,N_49594,N_49577);
nand UO_3987 (O_3987,N_49831,N_49054);
or UO_3988 (O_3988,N_49687,N_49494);
nand UO_3989 (O_3989,N_49249,N_49602);
and UO_3990 (O_3990,N_49926,N_49904);
and UO_3991 (O_3991,N_49283,N_49123);
or UO_3992 (O_3992,N_49724,N_49355);
or UO_3993 (O_3993,N_49506,N_49535);
nand UO_3994 (O_3994,N_49161,N_49265);
nand UO_3995 (O_3995,N_49833,N_49671);
nor UO_3996 (O_3996,N_49723,N_49712);
or UO_3997 (O_3997,N_49958,N_49361);
nand UO_3998 (O_3998,N_49236,N_49842);
and UO_3999 (O_3999,N_49381,N_49916);
nor UO_4000 (O_4000,N_49622,N_49811);
or UO_4001 (O_4001,N_49794,N_49641);
nand UO_4002 (O_4002,N_49588,N_49510);
or UO_4003 (O_4003,N_49066,N_49179);
nor UO_4004 (O_4004,N_49162,N_49858);
or UO_4005 (O_4005,N_49241,N_49495);
or UO_4006 (O_4006,N_49122,N_49646);
and UO_4007 (O_4007,N_49694,N_49744);
and UO_4008 (O_4008,N_49216,N_49364);
nand UO_4009 (O_4009,N_49837,N_49902);
nand UO_4010 (O_4010,N_49462,N_49271);
nor UO_4011 (O_4011,N_49507,N_49079);
or UO_4012 (O_4012,N_49408,N_49288);
nor UO_4013 (O_4013,N_49880,N_49614);
nor UO_4014 (O_4014,N_49560,N_49400);
nor UO_4015 (O_4015,N_49417,N_49621);
and UO_4016 (O_4016,N_49704,N_49712);
and UO_4017 (O_4017,N_49105,N_49704);
nor UO_4018 (O_4018,N_49917,N_49230);
and UO_4019 (O_4019,N_49277,N_49713);
xor UO_4020 (O_4020,N_49447,N_49474);
nand UO_4021 (O_4021,N_49980,N_49930);
and UO_4022 (O_4022,N_49794,N_49640);
nand UO_4023 (O_4023,N_49201,N_49138);
xor UO_4024 (O_4024,N_49234,N_49460);
nand UO_4025 (O_4025,N_49886,N_49588);
nand UO_4026 (O_4026,N_49550,N_49737);
xnor UO_4027 (O_4027,N_49170,N_49586);
or UO_4028 (O_4028,N_49900,N_49675);
nor UO_4029 (O_4029,N_49813,N_49420);
xor UO_4030 (O_4030,N_49999,N_49608);
or UO_4031 (O_4031,N_49881,N_49266);
or UO_4032 (O_4032,N_49661,N_49111);
nand UO_4033 (O_4033,N_49385,N_49421);
or UO_4034 (O_4034,N_49841,N_49214);
nor UO_4035 (O_4035,N_49491,N_49099);
or UO_4036 (O_4036,N_49210,N_49569);
nor UO_4037 (O_4037,N_49857,N_49548);
and UO_4038 (O_4038,N_49969,N_49591);
and UO_4039 (O_4039,N_49855,N_49997);
and UO_4040 (O_4040,N_49984,N_49677);
nor UO_4041 (O_4041,N_49186,N_49753);
or UO_4042 (O_4042,N_49113,N_49608);
or UO_4043 (O_4043,N_49597,N_49589);
nand UO_4044 (O_4044,N_49941,N_49585);
or UO_4045 (O_4045,N_49720,N_49238);
nor UO_4046 (O_4046,N_49901,N_49970);
nor UO_4047 (O_4047,N_49631,N_49119);
nor UO_4048 (O_4048,N_49436,N_49981);
nor UO_4049 (O_4049,N_49098,N_49938);
nor UO_4050 (O_4050,N_49236,N_49571);
nor UO_4051 (O_4051,N_49867,N_49346);
nor UO_4052 (O_4052,N_49114,N_49009);
nor UO_4053 (O_4053,N_49916,N_49332);
or UO_4054 (O_4054,N_49099,N_49727);
nand UO_4055 (O_4055,N_49744,N_49955);
and UO_4056 (O_4056,N_49357,N_49506);
nand UO_4057 (O_4057,N_49086,N_49444);
xnor UO_4058 (O_4058,N_49866,N_49855);
nor UO_4059 (O_4059,N_49111,N_49062);
and UO_4060 (O_4060,N_49117,N_49620);
nand UO_4061 (O_4061,N_49331,N_49893);
nand UO_4062 (O_4062,N_49331,N_49397);
nand UO_4063 (O_4063,N_49493,N_49005);
xnor UO_4064 (O_4064,N_49236,N_49605);
nor UO_4065 (O_4065,N_49734,N_49725);
xor UO_4066 (O_4066,N_49929,N_49446);
and UO_4067 (O_4067,N_49527,N_49011);
and UO_4068 (O_4068,N_49042,N_49773);
xor UO_4069 (O_4069,N_49464,N_49975);
xnor UO_4070 (O_4070,N_49967,N_49094);
xnor UO_4071 (O_4071,N_49293,N_49543);
nor UO_4072 (O_4072,N_49420,N_49973);
and UO_4073 (O_4073,N_49632,N_49474);
nand UO_4074 (O_4074,N_49103,N_49847);
or UO_4075 (O_4075,N_49834,N_49527);
nand UO_4076 (O_4076,N_49376,N_49998);
xnor UO_4077 (O_4077,N_49247,N_49695);
or UO_4078 (O_4078,N_49529,N_49135);
nor UO_4079 (O_4079,N_49254,N_49978);
or UO_4080 (O_4080,N_49506,N_49460);
nor UO_4081 (O_4081,N_49640,N_49706);
xor UO_4082 (O_4082,N_49809,N_49034);
and UO_4083 (O_4083,N_49481,N_49945);
xnor UO_4084 (O_4084,N_49496,N_49175);
nand UO_4085 (O_4085,N_49859,N_49188);
nor UO_4086 (O_4086,N_49253,N_49736);
nand UO_4087 (O_4087,N_49802,N_49202);
or UO_4088 (O_4088,N_49490,N_49461);
nand UO_4089 (O_4089,N_49953,N_49782);
and UO_4090 (O_4090,N_49069,N_49483);
or UO_4091 (O_4091,N_49539,N_49660);
and UO_4092 (O_4092,N_49049,N_49587);
or UO_4093 (O_4093,N_49298,N_49018);
and UO_4094 (O_4094,N_49095,N_49152);
or UO_4095 (O_4095,N_49318,N_49789);
nor UO_4096 (O_4096,N_49293,N_49297);
and UO_4097 (O_4097,N_49024,N_49216);
and UO_4098 (O_4098,N_49607,N_49832);
and UO_4099 (O_4099,N_49027,N_49412);
nor UO_4100 (O_4100,N_49358,N_49971);
and UO_4101 (O_4101,N_49105,N_49241);
or UO_4102 (O_4102,N_49576,N_49971);
xor UO_4103 (O_4103,N_49999,N_49331);
and UO_4104 (O_4104,N_49143,N_49076);
xor UO_4105 (O_4105,N_49761,N_49213);
and UO_4106 (O_4106,N_49894,N_49057);
nand UO_4107 (O_4107,N_49919,N_49092);
or UO_4108 (O_4108,N_49725,N_49873);
and UO_4109 (O_4109,N_49729,N_49952);
nand UO_4110 (O_4110,N_49126,N_49899);
or UO_4111 (O_4111,N_49233,N_49180);
and UO_4112 (O_4112,N_49670,N_49424);
nor UO_4113 (O_4113,N_49643,N_49959);
or UO_4114 (O_4114,N_49477,N_49509);
xnor UO_4115 (O_4115,N_49204,N_49322);
or UO_4116 (O_4116,N_49150,N_49497);
nor UO_4117 (O_4117,N_49659,N_49987);
nand UO_4118 (O_4118,N_49716,N_49320);
nor UO_4119 (O_4119,N_49852,N_49200);
nor UO_4120 (O_4120,N_49806,N_49214);
or UO_4121 (O_4121,N_49523,N_49617);
or UO_4122 (O_4122,N_49281,N_49382);
or UO_4123 (O_4123,N_49168,N_49488);
or UO_4124 (O_4124,N_49535,N_49903);
or UO_4125 (O_4125,N_49283,N_49006);
nand UO_4126 (O_4126,N_49409,N_49127);
nand UO_4127 (O_4127,N_49537,N_49410);
or UO_4128 (O_4128,N_49131,N_49662);
nand UO_4129 (O_4129,N_49101,N_49395);
and UO_4130 (O_4130,N_49024,N_49523);
nor UO_4131 (O_4131,N_49017,N_49057);
nor UO_4132 (O_4132,N_49465,N_49652);
xor UO_4133 (O_4133,N_49742,N_49245);
xnor UO_4134 (O_4134,N_49036,N_49803);
nand UO_4135 (O_4135,N_49013,N_49833);
nand UO_4136 (O_4136,N_49712,N_49763);
nor UO_4137 (O_4137,N_49434,N_49624);
nor UO_4138 (O_4138,N_49695,N_49415);
or UO_4139 (O_4139,N_49388,N_49190);
nor UO_4140 (O_4140,N_49314,N_49248);
nor UO_4141 (O_4141,N_49475,N_49333);
nor UO_4142 (O_4142,N_49881,N_49142);
nand UO_4143 (O_4143,N_49969,N_49826);
nor UO_4144 (O_4144,N_49093,N_49535);
or UO_4145 (O_4145,N_49956,N_49037);
or UO_4146 (O_4146,N_49731,N_49315);
nand UO_4147 (O_4147,N_49234,N_49336);
and UO_4148 (O_4148,N_49863,N_49203);
nor UO_4149 (O_4149,N_49782,N_49210);
or UO_4150 (O_4150,N_49684,N_49231);
nand UO_4151 (O_4151,N_49775,N_49273);
and UO_4152 (O_4152,N_49828,N_49583);
nand UO_4153 (O_4153,N_49818,N_49200);
nor UO_4154 (O_4154,N_49083,N_49232);
nor UO_4155 (O_4155,N_49651,N_49191);
nor UO_4156 (O_4156,N_49652,N_49925);
or UO_4157 (O_4157,N_49980,N_49826);
or UO_4158 (O_4158,N_49107,N_49672);
and UO_4159 (O_4159,N_49893,N_49781);
nand UO_4160 (O_4160,N_49794,N_49324);
xor UO_4161 (O_4161,N_49730,N_49076);
and UO_4162 (O_4162,N_49124,N_49886);
or UO_4163 (O_4163,N_49895,N_49583);
nand UO_4164 (O_4164,N_49435,N_49009);
xor UO_4165 (O_4165,N_49298,N_49863);
nor UO_4166 (O_4166,N_49037,N_49213);
and UO_4167 (O_4167,N_49069,N_49808);
nand UO_4168 (O_4168,N_49939,N_49183);
or UO_4169 (O_4169,N_49157,N_49070);
or UO_4170 (O_4170,N_49837,N_49982);
nand UO_4171 (O_4171,N_49773,N_49771);
nor UO_4172 (O_4172,N_49063,N_49324);
and UO_4173 (O_4173,N_49252,N_49686);
xnor UO_4174 (O_4174,N_49127,N_49096);
and UO_4175 (O_4175,N_49792,N_49014);
and UO_4176 (O_4176,N_49141,N_49996);
and UO_4177 (O_4177,N_49226,N_49841);
or UO_4178 (O_4178,N_49542,N_49600);
or UO_4179 (O_4179,N_49212,N_49963);
or UO_4180 (O_4180,N_49089,N_49997);
nand UO_4181 (O_4181,N_49934,N_49539);
and UO_4182 (O_4182,N_49205,N_49280);
xnor UO_4183 (O_4183,N_49984,N_49571);
or UO_4184 (O_4184,N_49569,N_49572);
xor UO_4185 (O_4185,N_49664,N_49731);
or UO_4186 (O_4186,N_49691,N_49785);
or UO_4187 (O_4187,N_49547,N_49350);
or UO_4188 (O_4188,N_49268,N_49450);
nor UO_4189 (O_4189,N_49578,N_49659);
xnor UO_4190 (O_4190,N_49098,N_49769);
nor UO_4191 (O_4191,N_49980,N_49924);
and UO_4192 (O_4192,N_49171,N_49110);
xor UO_4193 (O_4193,N_49967,N_49385);
or UO_4194 (O_4194,N_49043,N_49264);
xor UO_4195 (O_4195,N_49365,N_49919);
or UO_4196 (O_4196,N_49094,N_49070);
or UO_4197 (O_4197,N_49679,N_49070);
or UO_4198 (O_4198,N_49133,N_49389);
xor UO_4199 (O_4199,N_49164,N_49456);
or UO_4200 (O_4200,N_49062,N_49779);
and UO_4201 (O_4201,N_49840,N_49515);
nor UO_4202 (O_4202,N_49248,N_49828);
or UO_4203 (O_4203,N_49429,N_49828);
or UO_4204 (O_4204,N_49579,N_49250);
xor UO_4205 (O_4205,N_49940,N_49657);
and UO_4206 (O_4206,N_49338,N_49488);
nand UO_4207 (O_4207,N_49473,N_49738);
and UO_4208 (O_4208,N_49468,N_49867);
and UO_4209 (O_4209,N_49544,N_49604);
or UO_4210 (O_4210,N_49095,N_49485);
and UO_4211 (O_4211,N_49789,N_49307);
or UO_4212 (O_4212,N_49703,N_49364);
or UO_4213 (O_4213,N_49182,N_49688);
xor UO_4214 (O_4214,N_49157,N_49847);
nand UO_4215 (O_4215,N_49736,N_49291);
xnor UO_4216 (O_4216,N_49271,N_49231);
or UO_4217 (O_4217,N_49683,N_49110);
nor UO_4218 (O_4218,N_49707,N_49502);
nor UO_4219 (O_4219,N_49399,N_49569);
nand UO_4220 (O_4220,N_49016,N_49265);
xor UO_4221 (O_4221,N_49293,N_49382);
nand UO_4222 (O_4222,N_49542,N_49852);
nand UO_4223 (O_4223,N_49712,N_49934);
nor UO_4224 (O_4224,N_49178,N_49628);
xor UO_4225 (O_4225,N_49997,N_49550);
and UO_4226 (O_4226,N_49131,N_49952);
nor UO_4227 (O_4227,N_49024,N_49362);
nand UO_4228 (O_4228,N_49235,N_49461);
nand UO_4229 (O_4229,N_49997,N_49820);
xor UO_4230 (O_4230,N_49347,N_49808);
nand UO_4231 (O_4231,N_49305,N_49708);
and UO_4232 (O_4232,N_49039,N_49033);
xor UO_4233 (O_4233,N_49174,N_49026);
and UO_4234 (O_4234,N_49691,N_49391);
and UO_4235 (O_4235,N_49750,N_49866);
nand UO_4236 (O_4236,N_49865,N_49626);
nand UO_4237 (O_4237,N_49064,N_49220);
xnor UO_4238 (O_4238,N_49071,N_49859);
nand UO_4239 (O_4239,N_49835,N_49521);
xor UO_4240 (O_4240,N_49871,N_49576);
nor UO_4241 (O_4241,N_49418,N_49651);
nand UO_4242 (O_4242,N_49963,N_49458);
nor UO_4243 (O_4243,N_49953,N_49807);
xnor UO_4244 (O_4244,N_49192,N_49695);
xnor UO_4245 (O_4245,N_49868,N_49629);
or UO_4246 (O_4246,N_49587,N_49272);
xnor UO_4247 (O_4247,N_49116,N_49990);
xnor UO_4248 (O_4248,N_49954,N_49213);
nand UO_4249 (O_4249,N_49364,N_49333);
or UO_4250 (O_4250,N_49146,N_49713);
xnor UO_4251 (O_4251,N_49522,N_49069);
nor UO_4252 (O_4252,N_49991,N_49187);
nor UO_4253 (O_4253,N_49239,N_49756);
or UO_4254 (O_4254,N_49287,N_49648);
and UO_4255 (O_4255,N_49436,N_49686);
or UO_4256 (O_4256,N_49347,N_49224);
nand UO_4257 (O_4257,N_49643,N_49949);
nand UO_4258 (O_4258,N_49818,N_49583);
xnor UO_4259 (O_4259,N_49683,N_49396);
and UO_4260 (O_4260,N_49547,N_49670);
and UO_4261 (O_4261,N_49231,N_49177);
and UO_4262 (O_4262,N_49764,N_49317);
nor UO_4263 (O_4263,N_49127,N_49576);
nor UO_4264 (O_4264,N_49473,N_49644);
xnor UO_4265 (O_4265,N_49770,N_49843);
or UO_4266 (O_4266,N_49582,N_49922);
or UO_4267 (O_4267,N_49673,N_49533);
xnor UO_4268 (O_4268,N_49478,N_49611);
nand UO_4269 (O_4269,N_49355,N_49685);
and UO_4270 (O_4270,N_49351,N_49656);
nor UO_4271 (O_4271,N_49808,N_49486);
or UO_4272 (O_4272,N_49119,N_49642);
and UO_4273 (O_4273,N_49020,N_49843);
nor UO_4274 (O_4274,N_49182,N_49971);
xor UO_4275 (O_4275,N_49628,N_49423);
or UO_4276 (O_4276,N_49701,N_49703);
and UO_4277 (O_4277,N_49509,N_49812);
or UO_4278 (O_4278,N_49656,N_49795);
xnor UO_4279 (O_4279,N_49199,N_49023);
nor UO_4280 (O_4280,N_49921,N_49911);
or UO_4281 (O_4281,N_49279,N_49692);
nor UO_4282 (O_4282,N_49820,N_49942);
nor UO_4283 (O_4283,N_49727,N_49100);
nor UO_4284 (O_4284,N_49246,N_49136);
xnor UO_4285 (O_4285,N_49292,N_49059);
and UO_4286 (O_4286,N_49170,N_49116);
and UO_4287 (O_4287,N_49684,N_49868);
nand UO_4288 (O_4288,N_49731,N_49811);
and UO_4289 (O_4289,N_49755,N_49697);
nor UO_4290 (O_4290,N_49075,N_49649);
nand UO_4291 (O_4291,N_49596,N_49948);
or UO_4292 (O_4292,N_49392,N_49152);
nor UO_4293 (O_4293,N_49337,N_49747);
nor UO_4294 (O_4294,N_49715,N_49570);
or UO_4295 (O_4295,N_49628,N_49691);
xnor UO_4296 (O_4296,N_49336,N_49818);
xnor UO_4297 (O_4297,N_49563,N_49832);
xor UO_4298 (O_4298,N_49312,N_49667);
nand UO_4299 (O_4299,N_49407,N_49646);
nand UO_4300 (O_4300,N_49108,N_49695);
nor UO_4301 (O_4301,N_49388,N_49689);
nor UO_4302 (O_4302,N_49627,N_49629);
nor UO_4303 (O_4303,N_49089,N_49626);
or UO_4304 (O_4304,N_49405,N_49321);
and UO_4305 (O_4305,N_49860,N_49816);
or UO_4306 (O_4306,N_49300,N_49533);
xor UO_4307 (O_4307,N_49636,N_49474);
nand UO_4308 (O_4308,N_49682,N_49198);
nor UO_4309 (O_4309,N_49670,N_49727);
nand UO_4310 (O_4310,N_49122,N_49628);
xor UO_4311 (O_4311,N_49652,N_49182);
and UO_4312 (O_4312,N_49596,N_49845);
and UO_4313 (O_4313,N_49431,N_49288);
xor UO_4314 (O_4314,N_49427,N_49990);
nand UO_4315 (O_4315,N_49451,N_49383);
xor UO_4316 (O_4316,N_49270,N_49396);
and UO_4317 (O_4317,N_49091,N_49811);
or UO_4318 (O_4318,N_49789,N_49900);
nor UO_4319 (O_4319,N_49027,N_49069);
and UO_4320 (O_4320,N_49859,N_49529);
and UO_4321 (O_4321,N_49728,N_49213);
xor UO_4322 (O_4322,N_49023,N_49315);
nor UO_4323 (O_4323,N_49502,N_49226);
and UO_4324 (O_4324,N_49754,N_49190);
and UO_4325 (O_4325,N_49156,N_49823);
nand UO_4326 (O_4326,N_49726,N_49618);
nor UO_4327 (O_4327,N_49241,N_49446);
or UO_4328 (O_4328,N_49276,N_49119);
and UO_4329 (O_4329,N_49288,N_49584);
nor UO_4330 (O_4330,N_49200,N_49173);
nand UO_4331 (O_4331,N_49375,N_49207);
or UO_4332 (O_4332,N_49807,N_49752);
xnor UO_4333 (O_4333,N_49506,N_49637);
or UO_4334 (O_4334,N_49207,N_49799);
and UO_4335 (O_4335,N_49541,N_49203);
and UO_4336 (O_4336,N_49097,N_49430);
nand UO_4337 (O_4337,N_49414,N_49064);
or UO_4338 (O_4338,N_49999,N_49845);
or UO_4339 (O_4339,N_49128,N_49480);
nor UO_4340 (O_4340,N_49627,N_49287);
or UO_4341 (O_4341,N_49633,N_49989);
nor UO_4342 (O_4342,N_49054,N_49377);
and UO_4343 (O_4343,N_49126,N_49701);
nand UO_4344 (O_4344,N_49776,N_49343);
nor UO_4345 (O_4345,N_49164,N_49167);
or UO_4346 (O_4346,N_49003,N_49324);
or UO_4347 (O_4347,N_49515,N_49909);
nor UO_4348 (O_4348,N_49899,N_49698);
or UO_4349 (O_4349,N_49937,N_49110);
or UO_4350 (O_4350,N_49392,N_49670);
xor UO_4351 (O_4351,N_49086,N_49357);
nor UO_4352 (O_4352,N_49721,N_49522);
or UO_4353 (O_4353,N_49889,N_49036);
xnor UO_4354 (O_4354,N_49147,N_49698);
or UO_4355 (O_4355,N_49911,N_49466);
xor UO_4356 (O_4356,N_49271,N_49539);
and UO_4357 (O_4357,N_49966,N_49035);
nor UO_4358 (O_4358,N_49755,N_49447);
or UO_4359 (O_4359,N_49678,N_49209);
xnor UO_4360 (O_4360,N_49942,N_49092);
nor UO_4361 (O_4361,N_49611,N_49884);
or UO_4362 (O_4362,N_49408,N_49946);
and UO_4363 (O_4363,N_49094,N_49000);
nand UO_4364 (O_4364,N_49555,N_49479);
nor UO_4365 (O_4365,N_49784,N_49894);
and UO_4366 (O_4366,N_49985,N_49032);
nor UO_4367 (O_4367,N_49333,N_49397);
and UO_4368 (O_4368,N_49852,N_49046);
nand UO_4369 (O_4369,N_49688,N_49074);
nor UO_4370 (O_4370,N_49178,N_49140);
or UO_4371 (O_4371,N_49018,N_49916);
nor UO_4372 (O_4372,N_49020,N_49776);
or UO_4373 (O_4373,N_49857,N_49482);
nor UO_4374 (O_4374,N_49750,N_49683);
and UO_4375 (O_4375,N_49640,N_49205);
or UO_4376 (O_4376,N_49157,N_49896);
nor UO_4377 (O_4377,N_49369,N_49868);
xnor UO_4378 (O_4378,N_49789,N_49005);
nand UO_4379 (O_4379,N_49267,N_49878);
and UO_4380 (O_4380,N_49815,N_49515);
or UO_4381 (O_4381,N_49536,N_49599);
nand UO_4382 (O_4382,N_49647,N_49341);
and UO_4383 (O_4383,N_49296,N_49923);
and UO_4384 (O_4384,N_49090,N_49272);
or UO_4385 (O_4385,N_49928,N_49426);
or UO_4386 (O_4386,N_49855,N_49893);
nand UO_4387 (O_4387,N_49190,N_49597);
and UO_4388 (O_4388,N_49275,N_49198);
and UO_4389 (O_4389,N_49174,N_49084);
nand UO_4390 (O_4390,N_49012,N_49198);
or UO_4391 (O_4391,N_49301,N_49790);
nand UO_4392 (O_4392,N_49138,N_49636);
nand UO_4393 (O_4393,N_49168,N_49819);
nor UO_4394 (O_4394,N_49888,N_49950);
or UO_4395 (O_4395,N_49316,N_49900);
nand UO_4396 (O_4396,N_49870,N_49318);
nor UO_4397 (O_4397,N_49407,N_49415);
or UO_4398 (O_4398,N_49438,N_49892);
nor UO_4399 (O_4399,N_49814,N_49613);
and UO_4400 (O_4400,N_49163,N_49850);
nand UO_4401 (O_4401,N_49915,N_49796);
and UO_4402 (O_4402,N_49570,N_49592);
or UO_4403 (O_4403,N_49645,N_49071);
xnor UO_4404 (O_4404,N_49466,N_49029);
xor UO_4405 (O_4405,N_49776,N_49912);
nor UO_4406 (O_4406,N_49255,N_49733);
nor UO_4407 (O_4407,N_49303,N_49191);
nor UO_4408 (O_4408,N_49698,N_49980);
and UO_4409 (O_4409,N_49997,N_49043);
nor UO_4410 (O_4410,N_49670,N_49520);
or UO_4411 (O_4411,N_49437,N_49312);
nand UO_4412 (O_4412,N_49690,N_49328);
nand UO_4413 (O_4413,N_49578,N_49182);
or UO_4414 (O_4414,N_49692,N_49158);
nor UO_4415 (O_4415,N_49597,N_49702);
nor UO_4416 (O_4416,N_49715,N_49812);
xor UO_4417 (O_4417,N_49591,N_49434);
nor UO_4418 (O_4418,N_49962,N_49101);
or UO_4419 (O_4419,N_49613,N_49391);
or UO_4420 (O_4420,N_49210,N_49163);
nor UO_4421 (O_4421,N_49817,N_49228);
and UO_4422 (O_4422,N_49937,N_49686);
or UO_4423 (O_4423,N_49006,N_49409);
and UO_4424 (O_4424,N_49628,N_49817);
and UO_4425 (O_4425,N_49549,N_49576);
or UO_4426 (O_4426,N_49905,N_49499);
nor UO_4427 (O_4427,N_49938,N_49320);
xor UO_4428 (O_4428,N_49723,N_49883);
and UO_4429 (O_4429,N_49580,N_49495);
and UO_4430 (O_4430,N_49315,N_49254);
xnor UO_4431 (O_4431,N_49564,N_49969);
xor UO_4432 (O_4432,N_49960,N_49725);
nor UO_4433 (O_4433,N_49580,N_49354);
and UO_4434 (O_4434,N_49190,N_49253);
or UO_4435 (O_4435,N_49110,N_49282);
xnor UO_4436 (O_4436,N_49347,N_49326);
and UO_4437 (O_4437,N_49516,N_49320);
and UO_4438 (O_4438,N_49771,N_49664);
or UO_4439 (O_4439,N_49326,N_49654);
or UO_4440 (O_4440,N_49921,N_49695);
nor UO_4441 (O_4441,N_49596,N_49481);
nand UO_4442 (O_4442,N_49629,N_49752);
and UO_4443 (O_4443,N_49641,N_49629);
and UO_4444 (O_4444,N_49184,N_49984);
or UO_4445 (O_4445,N_49242,N_49587);
nand UO_4446 (O_4446,N_49366,N_49148);
nor UO_4447 (O_4447,N_49844,N_49780);
and UO_4448 (O_4448,N_49020,N_49939);
or UO_4449 (O_4449,N_49263,N_49991);
nand UO_4450 (O_4450,N_49960,N_49662);
nor UO_4451 (O_4451,N_49575,N_49215);
and UO_4452 (O_4452,N_49582,N_49229);
and UO_4453 (O_4453,N_49968,N_49627);
or UO_4454 (O_4454,N_49797,N_49783);
or UO_4455 (O_4455,N_49067,N_49970);
nor UO_4456 (O_4456,N_49764,N_49939);
nand UO_4457 (O_4457,N_49665,N_49976);
nand UO_4458 (O_4458,N_49331,N_49769);
xnor UO_4459 (O_4459,N_49954,N_49274);
nand UO_4460 (O_4460,N_49753,N_49741);
or UO_4461 (O_4461,N_49234,N_49197);
and UO_4462 (O_4462,N_49330,N_49551);
xor UO_4463 (O_4463,N_49861,N_49813);
xnor UO_4464 (O_4464,N_49134,N_49368);
nand UO_4465 (O_4465,N_49165,N_49366);
or UO_4466 (O_4466,N_49729,N_49862);
or UO_4467 (O_4467,N_49184,N_49686);
nand UO_4468 (O_4468,N_49947,N_49731);
and UO_4469 (O_4469,N_49558,N_49856);
and UO_4470 (O_4470,N_49767,N_49728);
and UO_4471 (O_4471,N_49312,N_49265);
nor UO_4472 (O_4472,N_49497,N_49026);
nand UO_4473 (O_4473,N_49021,N_49284);
nand UO_4474 (O_4474,N_49780,N_49541);
nor UO_4475 (O_4475,N_49543,N_49203);
xor UO_4476 (O_4476,N_49799,N_49287);
xor UO_4477 (O_4477,N_49593,N_49086);
xor UO_4478 (O_4478,N_49858,N_49584);
xor UO_4479 (O_4479,N_49751,N_49650);
xnor UO_4480 (O_4480,N_49006,N_49277);
and UO_4481 (O_4481,N_49069,N_49619);
and UO_4482 (O_4482,N_49909,N_49815);
or UO_4483 (O_4483,N_49871,N_49617);
nand UO_4484 (O_4484,N_49149,N_49170);
and UO_4485 (O_4485,N_49258,N_49381);
and UO_4486 (O_4486,N_49283,N_49385);
or UO_4487 (O_4487,N_49862,N_49490);
nand UO_4488 (O_4488,N_49776,N_49228);
and UO_4489 (O_4489,N_49651,N_49774);
nor UO_4490 (O_4490,N_49260,N_49670);
xnor UO_4491 (O_4491,N_49038,N_49010);
or UO_4492 (O_4492,N_49503,N_49959);
nand UO_4493 (O_4493,N_49720,N_49557);
nor UO_4494 (O_4494,N_49794,N_49890);
nand UO_4495 (O_4495,N_49515,N_49485);
or UO_4496 (O_4496,N_49677,N_49360);
nor UO_4497 (O_4497,N_49458,N_49928);
xor UO_4498 (O_4498,N_49298,N_49927);
nor UO_4499 (O_4499,N_49581,N_49818);
nand UO_4500 (O_4500,N_49258,N_49943);
nand UO_4501 (O_4501,N_49445,N_49171);
xor UO_4502 (O_4502,N_49427,N_49912);
nor UO_4503 (O_4503,N_49117,N_49256);
and UO_4504 (O_4504,N_49222,N_49583);
nand UO_4505 (O_4505,N_49180,N_49758);
and UO_4506 (O_4506,N_49592,N_49168);
nand UO_4507 (O_4507,N_49727,N_49957);
nand UO_4508 (O_4508,N_49415,N_49046);
and UO_4509 (O_4509,N_49636,N_49018);
and UO_4510 (O_4510,N_49619,N_49580);
nor UO_4511 (O_4511,N_49306,N_49456);
nor UO_4512 (O_4512,N_49334,N_49319);
nor UO_4513 (O_4513,N_49106,N_49781);
xnor UO_4514 (O_4514,N_49497,N_49819);
xor UO_4515 (O_4515,N_49328,N_49687);
nor UO_4516 (O_4516,N_49010,N_49328);
or UO_4517 (O_4517,N_49399,N_49850);
and UO_4518 (O_4518,N_49179,N_49113);
or UO_4519 (O_4519,N_49221,N_49718);
xnor UO_4520 (O_4520,N_49397,N_49425);
and UO_4521 (O_4521,N_49284,N_49082);
nor UO_4522 (O_4522,N_49771,N_49456);
nor UO_4523 (O_4523,N_49631,N_49252);
nand UO_4524 (O_4524,N_49525,N_49834);
or UO_4525 (O_4525,N_49055,N_49889);
xnor UO_4526 (O_4526,N_49529,N_49080);
nor UO_4527 (O_4527,N_49402,N_49854);
xnor UO_4528 (O_4528,N_49891,N_49019);
xnor UO_4529 (O_4529,N_49977,N_49379);
nor UO_4530 (O_4530,N_49896,N_49342);
nor UO_4531 (O_4531,N_49661,N_49198);
xnor UO_4532 (O_4532,N_49099,N_49716);
or UO_4533 (O_4533,N_49138,N_49876);
or UO_4534 (O_4534,N_49374,N_49283);
xnor UO_4535 (O_4535,N_49509,N_49729);
and UO_4536 (O_4536,N_49964,N_49097);
xor UO_4537 (O_4537,N_49636,N_49837);
xnor UO_4538 (O_4538,N_49745,N_49644);
and UO_4539 (O_4539,N_49549,N_49432);
nand UO_4540 (O_4540,N_49887,N_49176);
xnor UO_4541 (O_4541,N_49655,N_49269);
and UO_4542 (O_4542,N_49697,N_49850);
nor UO_4543 (O_4543,N_49567,N_49595);
and UO_4544 (O_4544,N_49769,N_49896);
and UO_4545 (O_4545,N_49726,N_49540);
xor UO_4546 (O_4546,N_49564,N_49926);
nand UO_4547 (O_4547,N_49379,N_49286);
xor UO_4548 (O_4548,N_49080,N_49447);
xor UO_4549 (O_4549,N_49236,N_49801);
nor UO_4550 (O_4550,N_49192,N_49588);
nor UO_4551 (O_4551,N_49071,N_49699);
and UO_4552 (O_4552,N_49906,N_49240);
nor UO_4553 (O_4553,N_49763,N_49796);
xor UO_4554 (O_4554,N_49499,N_49102);
or UO_4555 (O_4555,N_49576,N_49438);
or UO_4556 (O_4556,N_49578,N_49988);
or UO_4557 (O_4557,N_49305,N_49883);
and UO_4558 (O_4558,N_49726,N_49435);
nor UO_4559 (O_4559,N_49038,N_49969);
nor UO_4560 (O_4560,N_49203,N_49624);
nand UO_4561 (O_4561,N_49397,N_49152);
nand UO_4562 (O_4562,N_49078,N_49275);
xnor UO_4563 (O_4563,N_49558,N_49748);
xor UO_4564 (O_4564,N_49746,N_49446);
nor UO_4565 (O_4565,N_49039,N_49105);
and UO_4566 (O_4566,N_49647,N_49222);
nand UO_4567 (O_4567,N_49680,N_49169);
nand UO_4568 (O_4568,N_49146,N_49615);
or UO_4569 (O_4569,N_49368,N_49706);
xor UO_4570 (O_4570,N_49581,N_49247);
nor UO_4571 (O_4571,N_49307,N_49580);
nor UO_4572 (O_4572,N_49408,N_49798);
nor UO_4573 (O_4573,N_49288,N_49341);
nand UO_4574 (O_4574,N_49906,N_49305);
and UO_4575 (O_4575,N_49827,N_49559);
and UO_4576 (O_4576,N_49295,N_49743);
xnor UO_4577 (O_4577,N_49806,N_49753);
and UO_4578 (O_4578,N_49882,N_49236);
nand UO_4579 (O_4579,N_49951,N_49762);
and UO_4580 (O_4580,N_49481,N_49882);
nand UO_4581 (O_4581,N_49263,N_49772);
nand UO_4582 (O_4582,N_49325,N_49696);
nor UO_4583 (O_4583,N_49987,N_49558);
nand UO_4584 (O_4584,N_49985,N_49711);
nand UO_4585 (O_4585,N_49125,N_49219);
nor UO_4586 (O_4586,N_49960,N_49338);
or UO_4587 (O_4587,N_49007,N_49293);
xor UO_4588 (O_4588,N_49687,N_49685);
or UO_4589 (O_4589,N_49237,N_49467);
xnor UO_4590 (O_4590,N_49506,N_49560);
and UO_4591 (O_4591,N_49627,N_49621);
or UO_4592 (O_4592,N_49556,N_49627);
xnor UO_4593 (O_4593,N_49143,N_49419);
or UO_4594 (O_4594,N_49447,N_49194);
xor UO_4595 (O_4595,N_49883,N_49856);
nor UO_4596 (O_4596,N_49330,N_49065);
nor UO_4597 (O_4597,N_49521,N_49273);
nand UO_4598 (O_4598,N_49586,N_49288);
or UO_4599 (O_4599,N_49168,N_49840);
nand UO_4600 (O_4600,N_49028,N_49573);
and UO_4601 (O_4601,N_49263,N_49959);
nor UO_4602 (O_4602,N_49989,N_49586);
nor UO_4603 (O_4603,N_49591,N_49740);
and UO_4604 (O_4604,N_49881,N_49534);
and UO_4605 (O_4605,N_49623,N_49672);
xor UO_4606 (O_4606,N_49987,N_49548);
or UO_4607 (O_4607,N_49935,N_49617);
xor UO_4608 (O_4608,N_49996,N_49880);
xor UO_4609 (O_4609,N_49941,N_49042);
nor UO_4610 (O_4610,N_49225,N_49579);
nand UO_4611 (O_4611,N_49019,N_49925);
and UO_4612 (O_4612,N_49826,N_49138);
nor UO_4613 (O_4613,N_49846,N_49339);
nand UO_4614 (O_4614,N_49999,N_49300);
or UO_4615 (O_4615,N_49005,N_49008);
nor UO_4616 (O_4616,N_49569,N_49490);
xor UO_4617 (O_4617,N_49368,N_49103);
nand UO_4618 (O_4618,N_49907,N_49316);
nor UO_4619 (O_4619,N_49418,N_49890);
xnor UO_4620 (O_4620,N_49759,N_49038);
xor UO_4621 (O_4621,N_49932,N_49082);
nor UO_4622 (O_4622,N_49555,N_49522);
or UO_4623 (O_4623,N_49151,N_49291);
or UO_4624 (O_4624,N_49682,N_49115);
nand UO_4625 (O_4625,N_49820,N_49340);
nor UO_4626 (O_4626,N_49041,N_49982);
nand UO_4627 (O_4627,N_49280,N_49733);
nor UO_4628 (O_4628,N_49137,N_49654);
nand UO_4629 (O_4629,N_49716,N_49148);
nand UO_4630 (O_4630,N_49913,N_49500);
xor UO_4631 (O_4631,N_49153,N_49551);
or UO_4632 (O_4632,N_49904,N_49467);
nand UO_4633 (O_4633,N_49582,N_49417);
nand UO_4634 (O_4634,N_49033,N_49488);
nor UO_4635 (O_4635,N_49817,N_49099);
xor UO_4636 (O_4636,N_49099,N_49334);
xor UO_4637 (O_4637,N_49308,N_49778);
xnor UO_4638 (O_4638,N_49386,N_49294);
and UO_4639 (O_4639,N_49622,N_49674);
xor UO_4640 (O_4640,N_49083,N_49000);
xnor UO_4641 (O_4641,N_49237,N_49611);
nor UO_4642 (O_4642,N_49980,N_49124);
and UO_4643 (O_4643,N_49301,N_49141);
and UO_4644 (O_4644,N_49737,N_49755);
nand UO_4645 (O_4645,N_49871,N_49550);
nor UO_4646 (O_4646,N_49480,N_49420);
and UO_4647 (O_4647,N_49121,N_49799);
or UO_4648 (O_4648,N_49784,N_49109);
or UO_4649 (O_4649,N_49307,N_49049);
xnor UO_4650 (O_4650,N_49230,N_49680);
nor UO_4651 (O_4651,N_49709,N_49512);
or UO_4652 (O_4652,N_49568,N_49475);
xor UO_4653 (O_4653,N_49532,N_49022);
or UO_4654 (O_4654,N_49502,N_49003);
xnor UO_4655 (O_4655,N_49825,N_49744);
nor UO_4656 (O_4656,N_49415,N_49056);
xnor UO_4657 (O_4657,N_49106,N_49842);
nand UO_4658 (O_4658,N_49663,N_49915);
or UO_4659 (O_4659,N_49511,N_49302);
nand UO_4660 (O_4660,N_49043,N_49521);
xor UO_4661 (O_4661,N_49979,N_49698);
or UO_4662 (O_4662,N_49171,N_49098);
xor UO_4663 (O_4663,N_49335,N_49301);
xnor UO_4664 (O_4664,N_49498,N_49889);
and UO_4665 (O_4665,N_49860,N_49666);
or UO_4666 (O_4666,N_49153,N_49381);
xor UO_4667 (O_4667,N_49693,N_49468);
nand UO_4668 (O_4668,N_49730,N_49085);
and UO_4669 (O_4669,N_49511,N_49500);
xnor UO_4670 (O_4670,N_49720,N_49630);
or UO_4671 (O_4671,N_49734,N_49478);
nor UO_4672 (O_4672,N_49854,N_49774);
nor UO_4673 (O_4673,N_49731,N_49385);
or UO_4674 (O_4674,N_49463,N_49247);
or UO_4675 (O_4675,N_49364,N_49818);
nand UO_4676 (O_4676,N_49165,N_49138);
and UO_4677 (O_4677,N_49617,N_49894);
and UO_4678 (O_4678,N_49563,N_49902);
and UO_4679 (O_4679,N_49018,N_49297);
and UO_4680 (O_4680,N_49697,N_49581);
nor UO_4681 (O_4681,N_49793,N_49608);
and UO_4682 (O_4682,N_49803,N_49736);
and UO_4683 (O_4683,N_49530,N_49041);
xnor UO_4684 (O_4684,N_49905,N_49217);
nor UO_4685 (O_4685,N_49211,N_49556);
nor UO_4686 (O_4686,N_49574,N_49553);
and UO_4687 (O_4687,N_49585,N_49197);
xor UO_4688 (O_4688,N_49400,N_49067);
or UO_4689 (O_4689,N_49605,N_49171);
nor UO_4690 (O_4690,N_49467,N_49826);
nand UO_4691 (O_4691,N_49091,N_49189);
nor UO_4692 (O_4692,N_49302,N_49190);
or UO_4693 (O_4693,N_49131,N_49991);
and UO_4694 (O_4694,N_49273,N_49892);
or UO_4695 (O_4695,N_49794,N_49710);
xnor UO_4696 (O_4696,N_49832,N_49873);
xor UO_4697 (O_4697,N_49150,N_49886);
and UO_4698 (O_4698,N_49739,N_49339);
nor UO_4699 (O_4699,N_49091,N_49286);
nand UO_4700 (O_4700,N_49039,N_49606);
xnor UO_4701 (O_4701,N_49798,N_49371);
or UO_4702 (O_4702,N_49996,N_49773);
or UO_4703 (O_4703,N_49527,N_49510);
nand UO_4704 (O_4704,N_49179,N_49176);
nor UO_4705 (O_4705,N_49910,N_49748);
and UO_4706 (O_4706,N_49694,N_49438);
nor UO_4707 (O_4707,N_49677,N_49650);
nor UO_4708 (O_4708,N_49613,N_49208);
nand UO_4709 (O_4709,N_49049,N_49083);
or UO_4710 (O_4710,N_49993,N_49316);
nor UO_4711 (O_4711,N_49236,N_49863);
nor UO_4712 (O_4712,N_49397,N_49801);
xor UO_4713 (O_4713,N_49066,N_49943);
nand UO_4714 (O_4714,N_49816,N_49094);
xnor UO_4715 (O_4715,N_49363,N_49662);
or UO_4716 (O_4716,N_49504,N_49659);
and UO_4717 (O_4717,N_49415,N_49212);
or UO_4718 (O_4718,N_49996,N_49865);
and UO_4719 (O_4719,N_49227,N_49158);
nand UO_4720 (O_4720,N_49070,N_49730);
or UO_4721 (O_4721,N_49945,N_49735);
nor UO_4722 (O_4722,N_49162,N_49547);
or UO_4723 (O_4723,N_49002,N_49280);
nor UO_4724 (O_4724,N_49258,N_49146);
and UO_4725 (O_4725,N_49042,N_49593);
nand UO_4726 (O_4726,N_49148,N_49612);
nand UO_4727 (O_4727,N_49259,N_49508);
nor UO_4728 (O_4728,N_49646,N_49550);
nor UO_4729 (O_4729,N_49780,N_49078);
and UO_4730 (O_4730,N_49414,N_49953);
nor UO_4731 (O_4731,N_49168,N_49196);
nor UO_4732 (O_4732,N_49456,N_49288);
nand UO_4733 (O_4733,N_49142,N_49558);
xor UO_4734 (O_4734,N_49324,N_49972);
nor UO_4735 (O_4735,N_49978,N_49198);
xor UO_4736 (O_4736,N_49751,N_49243);
nor UO_4737 (O_4737,N_49690,N_49862);
nand UO_4738 (O_4738,N_49744,N_49251);
nand UO_4739 (O_4739,N_49517,N_49742);
or UO_4740 (O_4740,N_49678,N_49265);
nor UO_4741 (O_4741,N_49741,N_49822);
nor UO_4742 (O_4742,N_49598,N_49797);
nand UO_4743 (O_4743,N_49208,N_49465);
nand UO_4744 (O_4744,N_49541,N_49834);
nand UO_4745 (O_4745,N_49180,N_49622);
nor UO_4746 (O_4746,N_49522,N_49327);
xnor UO_4747 (O_4747,N_49312,N_49485);
or UO_4748 (O_4748,N_49199,N_49470);
or UO_4749 (O_4749,N_49026,N_49427);
xnor UO_4750 (O_4750,N_49537,N_49917);
nand UO_4751 (O_4751,N_49926,N_49217);
and UO_4752 (O_4752,N_49907,N_49032);
xor UO_4753 (O_4753,N_49163,N_49412);
nor UO_4754 (O_4754,N_49035,N_49545);
nand UO_4755 (O_4755,N_49815,N_49543);
xor UO_4756 (O_4756,N_49917,N_49359);
xnor UO_4757 (O_4757,N_49309,N_49586);
nor UO_4758 (O_4758,N_49684,N_49807);
or UO_4759 (O_4759,N_49412,N_49012);
and UO_4760 (O_4760,N_49714,N_49145);
and UO_4761 (O_4761,N_49061,N_49741);
xor UO_4762 (O_4762,N_49874,N_49578);
or UO_4763 (O_4763,N_49418,N_49663);
and UO_4764 (O_4764,N_49443,N_49188);
or UO_4765 (O_4765,N_49198,N_49001);
nand UO_4766 (O_4766,N_49885,N_49879);
and UO_4767 (O_4767,N_49549,N_49181);
and UO_4768 (O_4768,N_49847,N_49140);
and UO_4769 (O_4769,N_49400,N_49056);
xnor UO_4770 (O_4770,N_49565,N_49001);
nand UO_4771 (O_4771,N_49092,N_49429);
nand UO_4772 (O_4772,N_49721,N_49663);
nand UO_4773 (O_4773,N_49364,N_49759);
nor UO_4774 (O_4774,N_49667,N_49036);
nand UO_4775 (O_4775,N_49234,N_49816);
xor UO_4776 (O_4776,N_49137,N_49437);
nor UO_4777 (O_4777,N_49816,N_49589);
nand UO_4778 (O_4778,N_49597,N_49547);
or UO_4779 (O_4779,N_49849,N_49700);
or UO_4780 (O_4780,N_49805,N_49921);
or UO_4781 (O_4781,N_49918,N_49562);
xnor UO_4782 (O_4782,N_49062,N_49615);
and UO_4783 (O_4783,N_49519,N_49259);
or UO_4784 (O_4784,N_49364,N_49722);
and UO_4785 (O_4785,N_49367,N_49241);
xor UO_4786 (O_4786,N_49980,N_49357);
or UO_4787 (O_4787,N_49920,N_49357);
and UO_4788 (O_4788,N_49654,N_49121);
nor UO_4789 (O_4789,N_49459,N_49181);
nand UO_4790 (O_4790,N_49714,N_49252);
nor UO_4791 (O_4791,N_49317,N_49018);
nor UO_4792 (O_4792,N_49540,N_49745);
nor UO_4793 (O_4793,N_49597,N_49538);
xor UO_4794 (O_4794,N_49084,N_49786);
nand UO_4795 (O_4795,N_49834,N_49994);
xnor UO_4796 (O_4796,N_49209,N_49319);
xnor UO_4797 (O_4797,N_49269,N_49750);
or UO_4798 (O_4798,N_49314,N_49876);
nor UO_4799 (O_4799,N_49822,N_49889);
nor UO_4800 (O_4800,N_49475,N_49077);
xor UO_4801 (O_4801,N_49701,N_49592);
and UO_4802 (O_4802,N_49522,N_49456);
xnor UO_4803 (O_4803,N_49342,N_49570);
nor UO_4804 (O_4804,N_49949,N_49717);
nand UO_4805 (O_4805,N_49661,N_49136);
or UO_4806 (O_4806,N_49240,N_49995);
nor UO_4807 (O_4807,N_49362,N_49065);
xor UO_4808 (O_4808,N_49678,N_49281);
or UO_4809 (O_4809,N_49947,N_49313);
or UO_4810 (O_4810,N_49323,N_49135);
or UO_4811 (O_4811,N_49125,N_49814);
nand UO_4812 (O_4812,N_49171,N_49260);
or UO_4813 (O_4813,N_49437,N_49648);
and UO_4814 (O_4814,N_49977,N_49186);
nand UO_4815 (O_4815,N_49330,N_49119);
and UO_4816 (O_4816,N_49298,N_49050);
xor UO_4817 (O_4817,N_49201,N_49606);
and UO_4818 (O_4818,N_49979,N_49713);
or UO_4819 (O_4819,N_49197,N_49667);
nand UO_4820 (O_4820,N_49258,N_49368);
nor UO_4821 (O_4821,N_49623,N_49332);
nor UO_4822 (O_4822,N_49074,N_49001);
or UO_4823 (O_4823,N_49466,N_49722);
xor UO_4824 (O_4824,N_49297,N_49979);
nand UO_4825 (O_4825,N_49617,N_49330);
xor UO_4826 (O_4826,N_49124,N_49177);
and UO_4827 (O_4827,N_49467,N_49111);
nand UO_4828 (O_4828,N_49264,N_49263);
and UO_4829 (O_4829,N_49552,N_49230);
or UO_4830 (O_4830,N_49021,N_49097);
and UO_4831 (O_4831,N_49741,N_49542);
and UO_4832 (O_4832,N_49281,N_49246);
nor UO_4833 (O_4833,N_49269,N_49424);
xnor UO_4834 (O_4834,N_49863,N_49906);
nor UO_4835 (O_4835,N_49843,N_49722);
or UO_4836 (O_4836,N_49486,N_49935);
xnor UO_4837 (O_4837,N_49655,N_49914);
or UO_4838 (O_4838,N_49222,N_49376);
xnor UO_4839 (O_4839,N_49094,N_49058);
and UO_4840 (O_4840,N_49328,N_49646);
nor UO_4841 (O_4841,N_49655,N_49092);
nand UO_4842 (O_4842,N_49416,N_49266);
nor UO_4843 (O_4843,N_49632,N_49940);
nand UO_4844 (O_4844,N_49862,N_49215);
nand UO_4845 (O_4845,N_49934,N_49708);
nand UO_4846 (O_4846,N_49984,N_49365);
and UO_4847 (O_4847,N_49047,N_49232);
xor UO_4848 (O_4848,N_49980,N_49254);
and UO_4849 (O_4849,N_49347,N_49424);
and UO_4850 (O_4850,N_49141,N_49822);
and UO_4851 (O_4851,N_49610,N_49109);
nor UO_4852 (O_4852,N_49730,N_49438);
nand UO_4853 (O_4853,N_49853,N_49057);
nor UO_4854 (O_4854,N_49314,N_49809);
nor UO_4855 (O_4855,N_49125,N_49616);
xnor UO_4856 (O_4856,N_49044,N_49944);
or UO_4857 (O_4857,N_49764,N_49977);
or UO_4858 (O_4858,N_49238,N_49192);
or UO_4859 (O_4859,N_49458,N_49388);
nand UO_4860 (O_4860,N_49523,N_49018);
nor UO_4861 (O_4861,N_49778,N_49685);
or UO_4862 (O_4862,N_49383,N_49589);
xnor UO_4863 (O_4863,N_49424,N_49167);
and UO_4864 (O_4864,N_49131,N_49230);
or UO_4865 (O_4865,N_49060,N_49235);
nor UO_4866 (O_4866,N_49073,N_49416);
xnor UO_4867 (O_4867,N_49158,N_49299);
nand UO_4868 (O_4868,N_49085,N_49627);
and UO_4869 (O_4869,N_49294,N_49609);
or UO_4870 (O_4870,N_49017,N_49139);
xor UO_4871 (O_4871,N_49821,N_49958);
nor UO_4872 (O_4872,N_49063,N_49077);
and UO_4873 (O_4873,N_49298,N_49651);
or UO_4874 (O_4874,N_49440,N_49698);
or UO_4875 (O_4875,N_49716,N_49480);
nor UO_4876 (O_4876,N_49112,N_49462);
xor UO_4877 (O_4877,N_49781,N_49856);
nand UO_4878 (O_4878,N_49854,N_49273);
xor UO_4879 (O_4879,N_49088,N_49389);
and UO_4880 (O_4880,N_49746,N_49075);
and UO_4881 (O_4881,N_49043,N_49153);
or UO_4882 (O_4882,N_49964,N_49209);
xnor UO_4883 (O_4883,N_49057,N_49387);
nand UO_4884 (O_4884,N_49890,N_49350);
nand UO_4885 (O_4885,N_49397,N_49106);
or UO_4886 (O_4886,N_49432,N_49989);
and UO_4887 (O_4887,N_49277,N_49243);
xnor UO_4888 (O_4888,N_49945,N_49170);
and UO_4889 (O_4889,N_49203,N_49951);
and UO_4890 (O_4890,N_49667,N_49764);
xnor UO_4891 (O_4891,N_49435,N_49640);
nor UO_4892 (O_4892,N_49122,N_49348);
xor UO_4893 (O_4893,N_49360,N_49350);
nand UO_4894 (O_4894,N_49060,N_49799);
nor UO_4895 (O_4895,N_49474,N_49323);
nor UO_4896 (O_4896,N_49772,N_49060);
and UO_4897 (O_4897,N_49643,N_49435);
and UO_4898 (O_4898,N_49133,N_49773);
xor UO_4899 (O_4899,N_49350,N_49841);
and UO_4900 (O_4900,N_49378,N_49172);
xnor UO_4901 (O_4901,N_49957,N_49890);
nor UO_4902 (O_4902,N_49992,N_49069);
or UO_4903 (O_4903,N_49475,N_49294);
or UO_4904 (O_4904,N_49179,N_49587);
and UO_4905 (O_4905,N_49747,N_49902);
nor UO_4906 (O_4906,N_49240,N_49752);
nor UO_4907 (O_4907,N_49965,N_49554);
nand UO_4908 (O_4908,N_49420,N_49409);
xnor UO_4909 (O_4909,N_49098,N_49982);
and UO_4910 (O_4910,N_49421,N_49507);
nor UO_4911 (O_4911,N_49546,N_49435);
nand UO_4912 (O_4912,N_49458,N_49721);
xor UO_4913 (O_4913,N_49167,N_49589);
and UO_4914 (O_4914,N_49595,N_49749);
xor UO_4915 (O_4915,N_49103,N_49692);
nor UO_4916 (O_4916,N_49376,N_49154);
nand UO_4917 (O_4917,N_49940,N_49935);
xnor UO_4918 (O_4918,N_49198,N_49523);
nor UO_4919 (O_4919,N_49967,N_49289);
nor UO_4920 (O_4920,N_49488,N_49273);
nor UO_4921 (O_4921,N_49888,N_49314);
and UO_4922 (O_4922,N_49336,N_49040);
or UO_4923 (O_4923,N_49249,N_49263);
nand UO_4924 (O_4924,N_49565,N_49695);
nand UO_4925 (O_4925,N_49122,N_49477);
nor UO_4926 (O_4926,N_49430,N_49536);
nor UO_4927 (O_4927,N_49697,N_49767);
nand UO_4928 (O_4928,N_49056,N_49697);
nand UO_4929 (O_4929,N_49404,N_49492);
or UO_4930 (O_4930,N_49785,N_49762);
nand UO_4931 (O_4931,N_49824,N_49482);
nand UO_4932 (O_4932,N_49871,N_49471);
xor UO_4933 (O_4933,N_49659,N_49785);
and UO_4934 (O_4934,N_49026,N_49071);
and UO_4935 (O_4935,N_49359,N_49420);
nor UO_4936 (O_4936,N_49917,N_49886);
nand UO_4937 (O_4937,N_49709,N_49337);
xnor UO_4938 (O_4938,N_49225,N_49561);
nor UO_4939 (O_4939,N_49984,N_49722);
or UO_4940 (O_4940,N_49970,N_49487);
or UO_4941 (O_4941,N_49042,N_49412);
xnor UO_4942 (O_4942,N_49765,N_49017);
nor UO_4943 (O_4943,N_49722,N_49758);
nand UO_4944 (O_4944,N_49214,N_49581);
or UO_4945 (O_4945,N_49245,N_49061);
and UO_4946 (O_4946,N_49206,N_49884);
or UO_4947 (O_4947,N_49642,N_49419);
xor UO_4948 (O_4948,N_49116,N_49566);
and UO_4949 (O_4949,N_49950,N_49331);
nand UO_4950 (O_4950,N_49772,N_49630);
or UO_4951 (O_4951,N_49900,N_49688);
nor UO_4952 (O_4952,N_49089,N_49571);
xnor UO_4953 (O_4953,N_49446,N_49144);
and UO_4954 (O_4954,N_49856,N_49901);
nand UO_4955 (O_4955,N_49652,N_49387);
and UO_4956 (O_4956,N_49875,N_49756);
nor UO_4957 (O_4957,N_49658,N_49585);
or UO_4958 (O_4958,N_49188,N_49391);
xor UO_4959 (O_4959,N_49024,N_49657);
nor UO_4960 (O_4960,N_49165,N_49014);
or UO_4961 (O_4961,N_49111,N_49312);
nand UO_4962 (O_4962,N_49172,N_49475);
or UO_4963 (O_4963,N_49590,N_49847);
nand UO_4964 (O_4964,N_49079,N_49579);
nand UO_4965 (O_4965,N_49148,N_49486);
or UO_4966 (O_4966,N_49359,N_49781);
xnor UO_4967 (O_4967,N_49597,N_49635);
nand UO_4968 (O_4968,N_49973,N_49765);
nor UO_4969 (O_4969,N_49494,N_49444);
and UO_4970 (O_4970,N_49685,N_49924);
and UO_4971 (O_4971,N_49547,N_49705);
or UO_4972 (O_4972,N_49002,N_49267);
xor UO_4973 (O_4973,N_49742,N_49823);
nand UO_4974 (O_4974,N_49921,N_49077);
and UO_4975 (O_4975,N_49801,N_49841);
and UO_4976 (O_4976,N_49347,N_49992);
nand UO_4977 (O_4977,N_49449,N_49281);
or UO_4978 (O_4978,N_49609,N_49420);
xnor UO_4979 (O_4979,N_49211,N_49371);
nand UO_4980 (O_4980,N_49380,N_49500);
nor UO_4981 (O_4981,N_49463,N_49178);
or UO_4982 (O_4982,N_49087,N_49856);
nand UO_4983 (O_4983,N_49530,N_49279);
or UO_4984 (O_4984,N_49352,N_49792);
nand UO_4985 (O_4985,N_49330,N_49288);
or UO_4986 (O_4986,N_49738,N_49548);
and UO_4987 (O_4987,N_49955,N_49158);
and UO_4988 (O_4988,N_49606,N_49197);
xor UO_4989 (O_4989,N_49267,N_49909);
nor UO_4990 (O_4990,N_49228,N_49095);
xor UO_4991 (O_4991,N_49223,N_49163);
and UO_4992 (O_4992,N_49416,N_49588);
nand UO_4993 (O_4993,N_49983,N_49783);
or UO_4994 (O_4994,N_49511,N_49891);
nor UO_4995 (O_4995,N_49883,N_49645);
nor UO_4996 (O_4996,N_49081,N_49564);
nor UO_4997 (O_4997,N_49737,N_49129);
nor UO_4998 (O_4998,N_49653,N_49563);
or UO_4999 (O_4999,N_49478,N_49619);
endmodule