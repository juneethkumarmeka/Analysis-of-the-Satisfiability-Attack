module basic_750_5000_1000_10_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_359,In_630);
and U1 (N_1,In_733,In_634);
or U2 (N_2,In_111,In_233);
and U3 (N_3,In_223,In_641);
nand U4 (N_4,In_149,In_110);
nor U5 (N_5,In_382,In_441);
and U6 (N_6,In_131,In_188);
and U7 (N_7,In_406,In_332);
nor U8 (N_8,In_374,In_513);
nor U9 (N_9,In_372,In_124);
nor U10 (N_10,In_338,In_708);
or U11 (N_11,In_38,In_690);
nand U12 (N_12,In_646,In_526);
and U13 (N_13,In_468,In_366);
nand U14 (N_14,In_368,In_572);
and U15 (N_15,In_317,In_410);
nand U16 (N_16,In_55,In_23);
and U17 (N_17,In_325,In_692);
and U18 (N_18,In_621,In_527);
nand U19 (N_19,In_628,In_439);
nor U20 (N_20,In_531,In_252);
and U21 (N_21,In_369,In_289);
or U22 (N_22,In_578,In_389);
nor U23 (N_23,In_106,In_243);
nor U24 (N_24,In_134,In_503);
nor U25 (N_25,In_58,In_493);
nor U26 (N_26,In_525,In_228);
nor U27 (N_27,In_377,In_213);
or U28 (N_28,In_658,In_509);
and U29 (N_29,In_267,In_734);
nor U30 (N_30,In_222,In_484);
nor U31 (N_31,In_554,In_590);
or U32 (N_32,In_667,In_5);
nor U33 (N_33,In_595,In_284);
and U34 (N_34,In_73,In_594);
or U35 (N_35,In_492,In_523);
and U36 (N_36,In_614,In_730);
and U37 (N_37,In_120,In_370);
nor U38 (N_38,In_97,In_448);
and U39 (N_39,In_564,In_376);
and U40 (N_40,In_313,In_601);
xor U41 (N_41,In_547,In_112);
nand U42 (N_42,In_697,In_597);
nand U43 (N_43,In_13,In_447);
and U44 (N_44,In_424,In_123);
or U45 (N_45,In_113,In_655);
or U46 (N_46,In_218,In_612);
and U47 (N_47,In_463,In_203);
and U48 (N_48,In_155,In_105);
nand U49 (N_49,In_585,In_619);
nand U50 (N_50,In_748,In_82);
nor U51 (N_51,In_540,In_714);
or U52 (N_52,In_420,In_242);
nor U53 (N_53,In_170,In_573);
nor U54 (N_54,In_486,In_345);
and U55 (N_55,In_742,In_109);
nand U56 (N_56,In_225,In_268);
or U57 (N_57,In_740,In_732);
and U58 (N_58,In_373,In_207);
and U59 (N_59,In_434,In_545);
nand U60 (N_60,In_76,In_19);
nor U61 (N_61,In_472,In_495);
nor U62 (N_62,In_505,In_181);
and U63 (N_63,In_659,In_603);
or U64 (N_64,In_127,In_42);
and U65 (N_65,In_588,In_411);
or U66 (N_66,In_502,In_611);
nor U67 (N_67,In_549,In_744);
nand U68 (N_68,In_262,In_148);
or U69 (N_69,In_153,In_45);
and U70 (N_70,In_276,In_553);
nand U71 (N_71,In_602,In_164);
and U72 (N_72,In_536,In_670);
nor U73 (N_73,In_577,In_64);
and U74 (N_74,In_261,In_586);
or U75 (N_75,In_237,In_186);
or U76 (N_76,In_280,In_562);
or U77 (N_77,In_197,In_147);
nor U78 (N_78,In_741,In_168);
nor U79 (N_79,In_644,In_520);
or U80 (N_80,In_44,In_558);
or U81 (N_81,In_632,In_108);
nand U82 (N_82,In_639,In_299);
nor U83 (N_83,In_57,In_461);
and U84 (N_84,In_182,In_727);
and U85 (N_85,In_673,In_99);
nor U86 (N_86,In_446,In_140);
nor U87 (N_87,In_548,In_532);
and U88 (N_88,In_357,In_167);
xor U89 (N_89,In_189,In_426);
nand U90 (N_90,In_239,In_592);
and U91 (N_91,In_542,In_178);
or U92 (N_92,In_93,In_378);
or U93 (N_93,In_269,In_214);
and U94 (N_94,In_138,In_21);
or U95 (N_95,In_337,In_693);
and U96 (N_96,In_204,In_386);
or U97 (N_97,In_398,In_666);
nand U98 (N_98,In_622,In_83);
and U99 (N_99,In_437,In_724);
and U100 (N_100,In_662,In_226);
or U101 (N_101,In_24,In_653);
nand U102 (N_102,In_100,In_467);
nor U103 (N_103,In_422,In_728);
nor U104 (N_104,In_84,In_176);
and U105 (N_105,In_647,In_43);
and U106 (N_106,In_184,In_416);
and U107 (N_107,In_629,In_321);
nand U108 (N_108,In_241,In_414);
or U109 (N_109,In_118,In_388);
xnor U110 (N_110,In_60,In_713);
and U111 (N_111,In_198,In_75);
nand U112 (N_112,In_668,In_444);
and U113 (N_113,In_432,In_31);
nor U114 (N_114,In_557,In_343);
nand U115 (N_115,In_428,In_185);
or U116 (N_116,In_627,In_654);
and U117 (N_117,In_354,In_179);
or U118 (N_118,In_273,In_695);
nand U119 (N_119,In_353,In_92);
or U120 (N_120,In_687,In_686);
nand U121 (N_121,In_143,In_66);
nor U122 (N_122,In_429,In_624);
nor U123 (N_123,In_555,In_535);
or U124 (N_124,In_6,In_649);
nand U125 (N_125,In_291,In_516);
nor U126 (N_126,In_180,In_52);
nand U127 (N_127,In_550,In_236);
nor U128 (N_128,In_606,In_580);
and U129 (N_129,In_682,In_599);
and U130 (N_130,In_618,In_401);
or U131 (N_131,In_174,In_521);
or U132 (N_132,In_0,In_165);
nand U133 (N_133,In_596,In_16);
or U134 (N_134,In_543,In_150);
nand U135 (N_135,In_7,In_479);
or U136 (N_136,In_77,In_567);
or U137 (N_137,In_196,In_254);
nor U138 (N_138,In_315,In_613);
nor U139 (N_139,In_14,In_583);
nor U140 (N_140,In_417,In_605);
nand U141 (N_141,In_617,In_623);
nand U142 (N_142,In_249,In_669);
or U143 (N_143,In_304,In_663);
and U144 (N_144,In_729,In_508);
and U145 (N_145,In_642,In_735);
nor U146 (N_146,In_90,In_114);
nor U147 (N_147,In_286,In_344);
nand U148 (N_148,In_465,In_308);
nor U149 (N_149,In_559,In_419);
nor U150 (N_150,In_171,In_173);
and U151 (N_151,In_296,In_327);
and U152 (N_152,In_674,In_475);
or U153 (N_153,In_541,In_538);
or U154 (N_154,In_330,In_183);
or U155 (N_155,In_200,In_247);
or U156 (N_156,In_231,In_3);
nor U157 (N_157,In_498,In_470);
nor U158 (N_158,In_25,In_476);
and U159 (N_159,In_528,In_709);
and U160 (N_160,In_648,In_89);
nand U161 (N_161,In_85,In_442);
nor U162 (N_162,In_340,In_529);
nor U163 (N_163,In_88,In_240);
or U164 (N_164,In_347,In_719);
and U165 (N_165,In_193,In_440);
or U166 (N_166,In_318,In_506);
nand U167 (N_167,In_568,In_86);
nor U168 (N_168,In_297,In_229);
nand U169 (N_169,In_457,In_11);
nor U170 (N_170,In_404,In_309);
or U171 (N_171,In_556,In_339);
nor U172 (N_172,In_175,In_636);
and U173 (N_173,In_571,In_8);
nand U174 (N_174,In_40,In_707);
nor U175 (N_175,In_409,In_352);
or U176 (N_176,In_537,In_511);
nand U177 (N_177,In_1,In_598);
or U178 (N_178,In_563,In_546);
nand U179 (N_179,In_80,In_219);
nand U180 (N_180,In_435,In_22);
or U181 (N_181,In_530,In_518);
nand U182 (N_182,In_620,In_427);
or U183 (N_183,In_128,In_294);
or U184 (N_184,In_702,In_117);
and U185 (N_185,In_326,In_320);
nor U186 (N_186,In_177,In_122);
nand U187 (N_187,In_626,In_681);
nand U188 (N_188,In_350,In_358);
and U189 (N_189,In_224,In_95);
and U190 (N_190,In_699,In_41);
nor U191 (N_191,In_711,In_746);
or U192 (N_192,In_361,In_433);
and U193 (N_193,In_397,In_251);
and U194 (N_194,In_519,In_683);
nor U195 (N_195,In_387,In_657);
and U196 (N_196,In_221,In_15);
or U197 (N_197,In_608,In_49);
nor U198 (N_198,In_290,In_696);
nand U199 (N_199,In_72,In_474);
nand U200 (N_200,In_34,In_718);
and U201 (N_201,In_96,In_582);
or U202 (N_202,In_544,In_383);
and U203 (N_203,In_480,In_302);
or U204 (N_204,In_438,In_487);
or U205 (N_205,In_266,In_285);
nand U206 (N_206,In_379,In_314);
or U207 (N_207,In_640,In_270);
nand U208 (N_208,In_485,In_121);
and U209 (N_209,In_385,In_2);
and U210 (N_210,In_48,In_355);
nor U211 (N_211,In_551,In_561);
nor U212 (N_212,In_295,In_604);
and U213 (N_213,In_287,In_56);
nand U214 (N_214,In_698,In_232);
nand U215 (N_215,In_381,In_125);
or U216 (N_216,In_610,In_609);
nor U217 (N_217,In_584,In_201);
or U218 (N_218,In_736,In_104);
and U219 (N_219,In_160,In_615);
and U220 (N_220,In_635,In_216);
nor U221 (N_221,In_129,In_452);
nor U222 (N_222,In_334,In_625);
and U223 (N_223,In_208,In_192);
nor U224 (N_224,In_282,In_688);
nor U225 (N_225,In_703,In_685);
nand U226 (N_226,In_54,In_704);
nor U227 (N_227,In_691,In_616);
or U228 (N_228,In_26,In_749);
or U229 (N_229,In_271,In_489);
nor U230 (N_230,In_514,In_281);
and U231 (N_231,In_74,In_473);
or U232 (N_232,In_245,In_10);
and U233 (N_233,In_154,In_575);
nor U234 (N_234,In_20,In_510);
and U235 (N_235,In_471,In_399);
or U236 (N_236,In_211,In_70);
nor U237 (N_237,In_607,In_293);
or U238 (N_238,In_591,In_278);
nor U239 (N_239,In_190,In_29);
nand U240 (N_240,In_589,In_497);
nand U241 (N_241,In_569,In_600);
and U242 (N_242,In_35,In_68);
xnor U243 (N_243,In_483,In_715);
nand U244 (N_244,In_37,In_394);
and U245 (N_245,In_660,In_464);
nand U246 (N_246,In_720,In_362);
and U247 (N_247,In_512,In_212);
nor U248 (N_248,In_39,In_491);
nor U249 (N_249,In_552,In_135);
or U250 (N_250,In_169,In_81);
or U251 (N_251,In_316,In_283);
nand U252 (N_252,In_210,In_722);
and U253 (N_253,In_51,In_69);
nand U254 (N_254,In_126,In_94);
and U255 (N_255,In_33,In_712);
and U256 (N_256,In_425,In_462);
or U257 (N_257,In_671,In_507);
nor U258 (N_258,In_676,In_28);
and U259 (N_259,In_162,In_402);
and U260 (N_260,In_407,In_53);
or U261 (N_261,In_454,In_737);
nor U262 (N_262,In_253,In_408);
nor U263 (N_263,In_672,In_159);
nand U264 (N_264,In_494,In_431);
nor U265 (N_265,In_705,In_141);
or U266 (N_266,In_132,In_445);
nor U267 (N_267,In_460,In_328);
and U268 (N_268,In_264,In_499);
nor U269 (N_269,In_329,In_215);
nor U270 (N_270,In_65,In_59);
nor U271 (N_271,In_684,In_195);
and U272 (N_272,In_263,In_348);
xnor U273 (N_273,In_534,In_365);
or U274 (N_274,In_101,In_87);
or U275 (N_275,In_451,In_194);
and U276 (N_276,In_423,In_560);
nor U277 (N_277,In_393,In_675);
and U278 (N_278,In_488,In_139);
or U279 (N_279,In_103,In_166);
or U280 (N_280,In_115,In_651);
and U281 (N_281,In_650,In_300);
or U282 (N_282,In_107,In_119);
nand U283 (N_283,In_288,In_466);
nor U284 (N_284,In_701,In_477);
nor U285 (N_285,In_12,In_258);
or U286 (N_286,In_716,In_360);
nand U287 (N_287,In_9,In_205);
nand U288 (N_288,In_312,In_694);
nor U289 (N_289,In_230,In_581);
or U290 (N_290,In_136,In_371);
and U291 (N_291,In_310,In_656);
and U292 (N_292,In_335,In_305);
nand U293 (N_293,In_633,In_71);
or U294 (N_294,In_579,In_116);
nor U295 (N_295,In_652,In_391);
and U296 (N_296,In_248,In_430);
and U297 (N_297,In_206,In_78);
nor U298 (N_298,In_478,In_721);
nand U299 (N_299,In_375,In_235);
nor U300 (N_300,In_587,In_47);
or U301 (N_301,In_517,In_458);
nand U302 (N_302,In_333,In_346);
nand U303 (N_303,In_400,In_710);
or U304 (N_304,In_172,In_227);
or U305 (N_305,In_456,In_565);
and U306 (N_306,In_645,In_133);
or U307 (N_307,In_396,In_36);
nand U308 (N_308,In_678,In_323);
nand U309 (N_309,In_706,In_217);
or U310 (N_310,In_449,In_4);
nor U311 (N_311,In_256,In_380);
nor U312 (N_312,In_234,In_574);
nand U313 (N_313,In_331,In_700);
or U314 (N_314,In_46,In_161);
and U315 (N_315,In_303,In_539);
nor U316 (N_316,In_443,In_307);
and U317 (N_317,In_342,In_500);
or U318 (N_318,In_412,In_367);
nand U319 (N_319,In_341,In_50);
nor U320 (N_320,In_336,In_490);
nand U321 (N_321,In_91,In_726);
nand U322 (N_322,In_743,In_504);
or U323 (N_323,In_279,In_392);
or U324 (N_324,In_717,In_257);
and U325 (N_325,In_319,In_725);
or U326 (N_326,In_274,In_364);
or U327 (N_327,In_566,In_481);
or U328 (N_328,In_524,In_723);
nor U329 (N_329,In_418,In_144);
nor U330 (N_330,In_661,In_453);
or U331 (N_331,In_405,In_158);
nand U332 (N_332,In_260,In_18);
or U333 (N_333,In_311,In_356);
or U334 (N_334,In_67,In_250);
xnor U335 (N_335,In_515,In_259);
or U336 (N_336,In_30,In_421);
nand U337 (N_337,In_677,In_17);
or U338 (N_338,In_137,In_63);
nor U339 (N_339,In_27,In_32);
and U340 (N_340,In_631,In_415);
or U341 (N_341,In_152,In_220);
or U342 (N_342,In_277,In_98);
nand U343 (N_343,In_747,In_469);
nor U344 (N_344,In_151,In_322);
or U345 (N_345,In_238,In_665);
nor U346 (N_346,In_306,In_363);
and U347 (N_347,In_501,In_163);
nand U348 (N_348,In_413,In_202);
and U349 (N_349,In_255,In_637);
nand U350 (N_350,In_157,In_209);
nand U351 (N_351,In_533,In_244);
or U352 (N_352,In_496,In_146);
or U353 (N_353,In_301,In_731);
nor U354 (N_354,In_275,In_680);
and U355 (N_355,In_265,In_156);
or U356 (N_356,In_384,In_199);
and U357 (N_357,In_62,In_745);
or U358 (N_358,In_570,In_191);
and U359 (N_359,In_436,In_292);
or U360 (N_360,In_145,In_324);
and U361 (N_361,In_664,In_459);
or U362 (N_362,In_455,In_403);
or U363 (N_363,In_689,In_272);
nand U364 (N_364,In_576,In_395);
and U365 (N_365,In_246,In_522);
and U366 (N_366,In_643,In_79);
and U367 (N_367,In_130,In_390);
nor U368 (N_368,In_349,In_102);
nor U369 (N_369,In_187,In_298);
or U370 (N_370,In_679,In_482);
nand U371 (N_371,In_739,In_738);
nand U372 (N_372,In_351,In_450);
nor U373 (N_373,In_61,In_593);
nand U374 (N_374,In_142,In_638);
or U375 (N_375,In_258,In_632);
and U376 (N_376,In_60,In_223);
and U377 (N_377,In_312,In_3);
and U378 (N_378,In_507,In_292);
nor U379 (N_379,In_604,In_690);
nand U380 (N_380,In_413,In_389);
and U381 (N_381,In_144,In_485);
and U382 (N_382,In_130,In_33);
or U383 (N_383,In_271,In_272);
nor U384 (N_384,In_305,In_25);
nand U385 (N_385,In_318,In_397);
nand U386 (N_386,In_2,In_143);
or U387 (N_387,In_417,In_240);
or U388 (N_388,In_479,In_444);
nor U389 (N_389,In_434,In_93);
and U390 (N_390,In_215,In_703);
and U391 (N_391,In_681,In_285);
nand U392 (N_392,In_140,In_194);
xnor U393 (N_393,In_158,In_390);
nor U394 (N_394,In_578,In_522);
and U395 (N_395,In_466,In_588);
or U396 (N_396,In_463,In_24);
and U397 (N_397,In_343,In_391);
nor U398 (N_398,In_401,In_644);
nand U399 (N_399,In_386,In_28);
nand U400 (N_400,In_28,In_205);
and U401 (N_401,In_416,In_222);
and U402 (N_402,In_191,In_410);
or U403 (N_403,In_407,In_312);
nand U404 (N_404,In_347,In_368);
nor U405 (N_405,In_311,In_113);
xnor U406 (N_406,In_584,In_421);
or U407 (N_407,In_526,In_423);
nand U408 (N_408,In_720,In_278);
nor U409 (N_409,In_43,In_84);
or U410 (N_410,In_495,In_377);
or U411 (N_411,In_303,In_8);
nand U412 (N_412,In_691,In_621);
xor U413 (N_413,In_114,In_227);
or U414 (N_414,In_658,In_255);
nor U415 (N_415,In_33,In_684);
and U416 (N_416,In_542,In_155);
or U417 (N_417,In_596,In_227);
and U418 (N_418,In_680,In_258);
or U419 (N_419,In_70,In_364);
nor U420 (N_420,In_135,In_419);
nor U421 (N_421,In_373,In_554);
or U422 (N_422,In_704,In_588);
nor U423 (N_423,In_629,In_619);
nand U424 (N_424,In_702,In_457);
or U425 (N_425,In_547,In_442);
xnor U426 (N_426,In_668,In_611);
xnor U427 (N_427,In_303,In_16);
nand U428 (N_428,In_365,In_37);
or U429 (N_429,In_311,In_709);
nor U430 (N_430,In_318,In_252);
nand U431 (N_431,In_741,In_309);
or U432 (N_432,In_58,In_325);
nand U433 (N_433,In_727,In_523);
and U434 (N_434,In_663,In_30);
and U435 (N_435,In_372,In_18);
nor U436 (N_436,In_214,In_84);
and U437 (N_437,In_748,In_58);
or U438 (N_438,In_53,In_417);
nor U439 (N_439,In_31,In_643);
and U440 (N_440,In_571,In_227);
nand U441 (N_441,In_677,In_722);
nor U442 (N_442,In_720,In_482);
nor U443 (N_443,In_86,In_410);
or U444 (N_444,In_254,In_293);
nand U445 (N_445,In_493,In_483);
nor U446 (N_446,In_289,In_54);
nand U447 (N_447,In_422,In_447);
and U448 (N_448,In_714,In_602);
and U449 (N_449,In_108,In_106);
and U450 (N_450,In_250,In_526);
or U451 (N_451,In_582,In_309);
or U452 (N_452,In_247,In_288);
and U453 (N_453,In_83,In_462);
and U454 (N_454,In_571,In_35);
nand U455 (N_455,In_170,In_109);
nand U456 (N_456,In_337,In_681);
nand U457 (N_457,In_537,In_475);
nor U458 (N_458,In_103,In_38);
nor U459 (N_459,In_58,In_386);
nor U460 (N_460,In_113,In_732);
and U461 (N_461,In_296,In_31);
or U462 (N_462,In_611,In_685);
nor U463 (N_463,In_618,In_680);
nand U464 (N_464,In_208,In_448);
and U465 (N_465,In_393,In_343);
nor U466 (N_466,In_646,In_400);
nor U467 (N_467,In_493,In_120);
or U468 (N_468,In_372,In_444);
nor U469 (N_469,In_198,In_337);
or U470 (N_470,In_172,In_698);
nand U471 (N_471,In_449,In_93);
or U472 (N_472,In_442,In_288);
nand U473 (N_473,In_588,In_525);
nor U474 (N_474,In_722,In_659);
nand U475 (N_475,In_162,In_56);
and U476 (N_476,In_379,In_95);
nand U477 (N_477,In_534,In_370);
nor U478 (N_478,In_186,In_601);
nor U479 (N_479,In_623,In_412);
and U480 (N_480,In_126,In_270);
nor U481 (N_481,In_51,In_684);
nor U482 (N_482,In_217,In_408);
xnor U483 (N_483,In_10,In_668);
or U484 (N_484,In_620,In_695);
or U485 (N_485,In_691,In_459);
nand U486 (N_486,In_229,In_215);
nand U487 (N_487,In_566,In_59);
and U488 (N_488,In_362,In_394);
and U489 (N_489,In_569,In_560);
nand U490 (N_490,In_465,In_478);
and U491 (N_491,In_632,In_330);
or U492 (N_492,In_217,In_643);
nand U493 (N_493,In_140,In_252);
and U494 (N_494,In_103,In_195);
or U495 (N_495,In_697,In_114);
nor U496 (N_496,In_456,In_528);
nand U497 (N_497,In_493,In_454);
nor U498 (N_498,In_620,In_605);
and U499 (N_499,In_219,In_128);
nor U500 (N_500,N_384,N_493);
or U501 (N_501,N_491,N_119);
or U502 (N_502,N_0,N_74);
nand U503 (N_503,N_34,N_390);
nor U504 (N_504,N_197,N_355);
nand U505 (N_505,N_262,N_461);
nand U506 (N_506,N_454,N_372);
nand U507 (N_507,N_125,N_349);
nor U508 (N_508,N_367,N_344);
or U509 (N_509,N_183,N_200);
and U510 (N_510,N_171,N_7);
or U511 (N_511,N_338,N_305);
or U512 (N_512,N_20,N_335);
or U513 (N_513,N_45,N_463);
nor U514 (N_514,N_421,N_253);
and U515 (N_515,N_292,N_66);
nand U516 (N_516,N_481,N_206);
nand U517 (N_517,N_269,N_356);
or U518 (N_518,N_361,N_170);
and U519 (N_519,N_208,N_113);
nand U520 (N_520,N_209,N_373);
nand U521 (N_521,N_64,N_59);
nor U522 (N_522,N_212,N_179);
and U523 (N_523,N_231,N_8);
or U524 (N_524,N_464,N_260);
or U525 (N_525,N_104,N_385);
and U526 (N_526,N_340,N_342);
or U527 (N_527,N_453,N_249);
or U528 (N_528,N_75,N_409);
nand U529 (N_529,N_275,N_380);
nand U530 (N_530,N_479,N_279);
nor U531 (N_531,N_163,N_194);
and U532 (N_532,N_118,N_255);
and U533 (N_533,N_254,N_416);
or U534 (N_534,N_16,N_6);
nand U535 (N_535,N_304,N_175);
or U536 (N_536,N_314,N_432);
and U537 (N_537,N_233,N_497);
nand U538 (N_538,N_450,N_230);
nand U539 (N_539,N_474,N_297);
and U540 (N_540,N_401,N_376);
or U541 (N_541,N_382,N_40);
nand U542 (N_542,N_133,N_307);
and U543 (N_543,N_404,N_121);
nor U544 (N_544,N_465,N_17);
nand U545 (N_545,N_167,N_186);
and U546 (N_546,N_131,N_389);
or U547 (N_547,N_190,N_144);
or U548 (N_548,N_318,N_41);
or U549 (N_549,N_429,N_483);
nand U550 (N_550,N_63,N_241);
nand U551 (N_551,N_21,N_30);
or U552 (N_552,N_236,N_298);
nand U553 (N_553,N_224,N_283);
or U554 (N_554,N_132,N_343);
nand U555 (N_555,N_383,N_152);
nor U556 (N_556,N_61,N_245);
nand U557 (N_557,N_123,N_29);
or U558 (N_558,N_146,N_55);
nand U559 (N_559,N_265,N_435);
nand U560 (N_560,N_378,N_4);
and U561 (N_561,N_311,N_109);
nand U562 (N_562,N_138,N_181);
nand U563 (N_563,N_237,N_334);
and U564 (N_564,N_227,N_428);
and U565 (N_565,N_191,N_103);
or U566 (N_566,N_422,N_106);
nand U567 (N_567,N_440,N_470);
or U568 (N_568,N_351,N_370);
or U569 (N_569,N_168,N_290);
and U570 (N_570,N_176,N_221);
and U571 (N_571,N_90,N_177);
or U572 (N_572,N_281,N_51);
and U573 (N_573,N_219,N_486);
nand U574 (N_574,N_19,N_160);
or U575 (N_575,N_328,N_252);
or U576 (N_576,N_295,N_434);
nor U577 (N_577,N_431,N_316);
nand U578 (N_578,N_353,N_69);
nor U579 (N_579,N_216,N_98);
nand U580 (N_580,N_50,N_325);
and U581 (N_581,N_229,N_47);
nand U582 (N_582,N_388,N_495);
and U583 (N_583,N_57,N_204);
or U584 (N_584,N_226,N_419);
and U585 (N_585,N_195,N_79);
or U586 (N_586,N_360,N_306);
nand U587 (N_587,N_358,N_15);
nand U588 (N_588,N_25,N_484);
and U589 (N_589,N_95,N_80);
nand U590 (N_590,N_157,N_331);
nand U591 (N_591,N_174,N_150);
or U592 (N_592,N_143,N_257);
or U593 (N_593,N_151,N_140);
and U594 (N_594,N_147,N_498);
and U595 (N_595,N_345,N_217);
nor U596 (N_596,N_72,N_202);
and U597 (N_597,N_359,N_398);
nand U598 (N_598,N_412,N_366);
and U599 (N_599,N_251,N_38);
nor U600 (N_600,N_134,N_472);
or U601 (N_601,N_101,N_270);
nor U602 (N_602,N_264,N_299);
or U603 (N_603,N_426,N_112);
and U604 (N_604,N_324,N_452);
nand U605 (N_605,N_87,N_84);
and U606 (N_606,N_271,N_399);
nor U607 (N_607,N_27,N_89);
nor U608 (N_608,N_33,N_102);
and U609 (N_609,N_192,N_363);
nand U610 (N_610,N_142,N_267);
and U611 (N_611,N_415,N_213);
or U612 (N_612,N_327,N_128);
nand U613 (N_613,N_165,N_261);
nand U614 (N_614,N_396,N_365);
and U615 (N_615,N_291,N_184);
nand U616 (N_616,N_433,N_185);
nor U617 (N_617,N_162,N_395);
nand U618 (N_618,N_43,N_78);
nand U619 (N_619,N_466,N_81);
and U620 (N_620,N_456,N_336);
or U621 (N_621,N_12,N_468);
nand U622 (N_622,N_469,N_259);
nand U623 (N_623,N_476,N_490);
nor U624 (N_624,N_26,N_294);
nand U625 (N_625,N_284,N_228);
or U626 (N_626,N_499,N_148);
or U627 (N_627,N_203,N_56);
nand U628 (N_628,N_321,N_341);
nor U629 (N_629,N_193,N_444);
or U630 (N_630,N_449,N_53);
nor U631 (N_631,N_127,N_489);
nand U632 (N_632,N_392,N_52);
nor U633 (N_633,N_94,N_408);
and U634 (N_634,N_242,N_480);
and U635 (N_635,N_166,N_425);
xor U636 (N_636,N_477,N_446);
nand U637 (N_637,N_473,N_110);
nor U638 (N_638,N_354,N_445);
or U639 (N_639,N_207,N_39);
nor U640 (N_640,N_350,N_418);
nor U641 (N_641,N_402,N_240);
and U642 (N_642,N_139,N_149);
nor U643 (N_643,N_141,N_386);
nor U644 (N_644,N_315,N_459);
and U645 (N_645,N_405,N_215);
or U646 (N_646,N_250,N_169);
or U647 (N_647,N_88,N_234);
nor U648 (N_648,N_13,N_263);
nor U649 (N_649,N_205,N_130);
and U650 (N_650,N_492,N_218);
or U651 (N_651,N_457,N_210);
nand U652 (N_652,N_96,N_180);
nand U653 (N_653,N_332,N_277);
or U654 (N_654,N_309,N_485);
nor U655 (N_655,N_420,N_49);
or U656 (N_656,N_46,N_124);
or U657 (N_657,N_153,N_154);
nor U658 (N_658,N_278,N_317);
and U659 (N_659,N_482,N_312);
and U660 (N_660,N_10,N_442);
nor U661 (N_661,N_164,N_310);
nor U662 (N_662,N_268,N_313);
or U663 (N_663,N_379,N_320);
or U664 (N_664,N_77,N_411);
nor U665 (N_665,N_375,N_400);
or U666 (N_666,N_467,N_282);
nor U667 (N_667,N_371,N_68);
and U668 (N_668,N_48,N_3);
nor U669 (N_669,N_9,N_54);
nand U670 (N_670,N_460,N_451);
nand U671 (N_671,N_222,N_182);
or U672 (N_672,N_329,N_289);
nand U673 (N_673,N_394,N_173);
or U674 (N_674,N_447,N_397);
and U675 (N_675,N_246,N_407);
nor U676 (N_676,N_410,N_301);
nand U677 (N_677,N_274,N_145);
nand U678 (N_678,N_238,N_427);
nand U679 (N_679,N_302,N_232);
and U680 (N_680,N_424,N_114);
and U681 (N_681,N_462,N_1);
nand U682 (N_682,N_136,N_478);
and U683 (N_683,N_28,N_187);
nor U684 (N_684,N_116,N_158);
or U685 (N_685,N_35,N_188);
nor U686 (N_686,N_235,N_296);
nor U687 (N_687,N_487,N_5);
and U688 (N_688,N_137,N_248);
nor U689 (N_689,N_417,N_196);
nor U690 (N_690,N_172,N_239);
nand U691 (N_691,N_36,N_11);
and U692 (N_692,N_377,N_494);
nor U693 (N_693,N_42,N_330);
nand U694 (N_694,N_266,N_326);
or U695 (N_695,N_91,N_244);
or U696 (N_696,N_437,N_67);
and U697 (N_697,N_111,N_243);
and U698 (N_698,N_70,N_293);
nand U699 (N_699,N_413,N_100);
and U700 (N_700,N_117,N_120);
nor U701 (N_701,N_308,N_272);
nand U702 (N_702,N_155,N_135);
and U703 (N_703,N_438,N_107);
nor U704 (N_704,N_288,N_86);
and U705 (N_705,N_280,N_76);
nor U706 (N_706,N_333,N_256);
nand U707 (N_707,N_73,N_475);
nand U708 (N_708,N_225,N_441);
nand U709 (N_709,N_31,N_339);
nand U710 (N_710,N_414,N_71);
or U711 (N_711,N_362,N_93);
and U712 (N_712,N_37,N_448);
nand U713 (N_713,N_82,N_108);
nand U714 (N_714,N_273,N_423);
or U715 (N_715,N_60,N_223);
and U716 (N_716,N_85,N_22);
and U717 (N_717,N_44,N_247);
nor U718 (N_718,N_496,N_115);
and U719 (N_719,N_322,N_348);
or U720 (N_720,N_23,N_287);
nand U721 (N_721,N_65,N_97);
nand U722 (N_722,N_14,N_99);
nor U723 (N_723,N_156,N_488);
nor U724 (N_724,N_126,N_347);
or U725 (N_725,N_276,N_58);
nor U726 (N_726,N_357,N_211);
nand U727 (N_727,N_436,N_430);
nor U728 (N_728,N_285,N_300);
nand U729 (N_729,N_381,N_323);
nand U730 (N_730,N_364,N_319);
or U731 (N_731,N_443,N_406);
or U732 (N_732,N_286,N_199);
nor U733 (N_733,N_122,N_214);
and U734 (N_734,N_201,N_337);
nor U735 (N_735,N_393,N_198);
or U736 (N_736,N_105,N_178);
and U737 (N_737,N_303,N_24);
nand U738 (N_738,N_83,N_2);
nand U739 (N_739,N_18,N_258);
and U740 (N_740,N_458,N_439);
nand U741 (N_741,N_161,N_62);
nor U742 (N_742,N_92,N_189);
and U743 (N_743,N_403,N_391);
nor U744 (N_744,N_220,N_346);
or U745 (N_745,N_352,N_455);
nand U746 (N_746,N_159,N_129);
or U747 (N_747,N_32,N_471);
and U748 (N_748,N_368,N_369);
nor U749 (N_749,N_374,N_387);
and U750 (N_750,N_432,N_398);
or U751 (N_751,N_303,N_499);
nand U752 (N_752,N_70,N_187);
and U753 (N_753,N_46,N_383);
and U754 (N_754,N_255,N_176);
or U755 (N_755,N_40,N_261);
nand U756 (N_756,N_369,N_127);
or U757 (N_757,N_185,N_285);
nor U758 (N_758,N_96,N_188);
nor U759 (N_759,N_411,N_275);
or U760 (N_760,N_185,N_265);
and U761 (N_761,N_324,N_137);
nor U762 (N_762,N_465,N_279);
nor U763 (N_763,N_97,N_464);
nand U764 (N_764,N_248,N_24);
or U765 (N_765,N_403,N_284);
nand U766 (N_766,N_155,N_236);
nand U767 (N_767,N_96,N_182);
nor U768 (N_768,N_255,N_291);
nand U769 (N_769,N_276,N_113);
nor U770 (N_770,N_398,N_448);
or U771 (N_771,N_299,N_438);
nor U772 (N_772,N_282,N_34);
and U773 (N_773,N_8,N_112);
nor U774 (N_774,N_136,N_336);
nand U775 (N_775,N_443,N_323);
nand U776 (N_776,N_258,N_113);
or U777 (N_777,N_16,N_73);
nor U778 (N_778,N_306,N_177);
nor U779 (N_779,N_470,N_279);
nor U780 (N_780,N_337,N_32);
and U781 (N_781,N_422,N_207);
and U782 (N_782,N_97,N_132);
nand U783 (N_783,N_206,N_104);
nor U784 (N_784,N_31,N_103);
nand U785 (N_785,N_449,N_392);
nor U786 (N_786,N_52,N_396);
and U787 (N_787,N_399,N_238);
or U788 (N_788,N_325,N_99);
or U789 (N_789,N_116,N_289);
nand U790 (N_790,N_309,N_188);
and U791 (N_791,N_95,N_108);
nor U792 (N_792,N_134,N_308);
nand U793 (N_793,N_199,N_438);
nand U794 (N_794,N_309,N_354);
and U795 (N_795,N_434,N_80);
or U796 (N_796,N_244,N_266);
nor U797 (N_797,N_386,N_121);
and U798 (N_798,N_209,N_1);
nor U799 (N_799,N_0,N_139);
and U800 (N_800,N_133,N_13);
nand U801 (N_801,N_58,N_354);
or U802 (N_802,N_492,N_67);
or U803 (N_803,N_200,N_176);
nand U804 (N_804,N_235,N_153);
or U805 (N_805,N_446,N_245);
nand U806 (N_806,N_139,N_274);
nor U807 (N_807,N_188,N_443);
nor U808 (N_808,N_75,N_240);
or U809 (N_809,N_65,N_292);
nor U810 (N_810,N_96,N_216);
nor U811 (N_811,N_110,N_25);
nor U812 (N_812,N_342,N_59);
and U813 (N_813,N_60,N_470);
nand U814 (N_814,N_343,N_454);
or U815 (N_815,N_471,N_247);
and U816 (N_816,N_375,N_402);
nand U817 (N_817,N_232,N_245);
or U818 (N_818,N_370,N_329);
nand U819 (N_819,N_139,N_410);
nand U820 (N_820,N_259,N_217);
nand U821 (N_821,N_0,N_443);
nor U822 (N_822,N_18,N_189);
nand U823 (N_823,N_37,N_41);
nand U824 (N_824,N_326,N_497);
nand U825 (N_825,N_478,N_97);
or U826 (N_826,N_244,N_184);
or U827 (N_827,N_354,N_92);
or U828 (N_828,N_200,N_383);
nand U829 (N_829,N_145,N_178);
or U830 (N_830,N_398,N_60);
nor U831 (N_831,N_185,N_466);
and U832 (N_832,N_364,N_247);
or U833 (N_833,N_419,N_258);
or U834 (N_834,N_225,N_435);
or U835 (N_835,N_287,N_0);
nand U836 (N_836,N_247,N_165);
and U837 (N_837,N_276,N_306);
nor U838 (N_838,N_114,N_418);
nand U839 (N_839,N_128,N_41);
and U840 (N_840,N_352,N_12);
nand U841 (N_841,N_492,N_184);
nand U842 (N_842,N_368,N_394);
nand U843 (N_843,N_4,N_73);
nor U844 (N_844,N_49,N_296);
and U845 (N_845,N_291,N_313);
and U846 (N_846,N_120,N_17);
or U847 (N_847,N_290,N_90);
or U848 (N_848,N_49,N_413);
and U849 (N_849,N_35,N_28);
or U850 (N_850,N_298,N_16);
nor U851 (N_851,N_352,N_257);
xor U852 (N_852,N_299,N_237);
and U853 (N_853,N_292,N_351);
nand U854 (N_854,N_243,N_279);
nor U855 (N_855,N_368,N_286);
or U856 (N_856,N_199,N_468);
or U857 (N_857,N_141,N_370);
nor U858 (N_858,N_50,N_331);
nand U859 (N_859,N_377,N_452);
nand U860 (N_860,N_429,N_466);
nand U861 (N_861,N_177,N_498);
and U862 (N_862,N_387,N_382);
or U863 (N_863,N_25,N_3);
nand U864 (N_864,N_219,N_353);
nor U865 (N_865,N_218,N_322);
nor U866 (N_866,N_495,N_265);
and U867 (N_867,N_78,N_411);
nand U868 (N_868,N_169,N_43);
nand U869 (N_869,N_7,N_189);
xnor U870 (N_870,N_498,N_148);
or U871 (N_871,N_100,N_326);
nor U872 (N_872,N_249,N_110);
or U873 (N_873,N_426,N_473);
or U874 (N_874,N_328,N_341);
nand U875 (N_875,N_245,N_241);
nand U876 (N_876,N_443,N_23);
or U877 (N_877,N_367,N_212);
nand U878 (N_878,N_449,N_97);
nor U879 (N_879,N_441,N_331);
nand U880 (N_880,N_494,N_277);
and U881 (N_881,N_148,N_59);
nand U882 (N_882,N_56,N_132);
or U883 (N_883,N_167,N_321);
nand U884 (N_884,N_423,N_292);
nor U885 (N_885,N_401,N_186);
or U886 (N_886,N_387,N_286);
nand U887 (N_887,N_140,N_216);
nand U888 (N_888,N_55,N_412);
nor U889 (N_889,N_277,N_38);
and U890 (N_890,N_379,N_337);
nor U891 (N_891,N_25,N_48);
nand U892 (N_892,N_212,N_361);
nand U893 (N_893,N_309,N_247);
or U894 (N_894,N_50,N_7);
nand U895 (N_895,N_434,N_424);
or U896 (N_896,N_107,N_103);
nor U897 (N_897,N_223,N_227);
or U898 (N_898,N_147,N_63);
and U899 (N_899,N_238,N_178);
and U900 (N_900,N_158,N_135);
nor U901 (N_901,N_420,N_81);
or U902 (N_902,N_103,N_330);
nor U903 (N_903,N_280,N_395);
or U904 (N_904,N_390,N_272);
or U905 (N_905,N_246,N_238);
or U906 (N_906,N_185,N_121);
nand U907 (N_907,N_158,N_237);
or U908 (N_908,N_154,N_204);
or U909 (N_909,N_429,N_373);
nand U910 (N_910,N_8,N_470);
or U911 (N_911,N_97,N_121);
and U912 (N_912,N_121,N_235);
or U913 (N_913,N_368,N_268);
nor U914 (N_914,N_441,N_446);
nand U915 (N_915,N_20,N_458);
or U916 (N_916,N_62,N_216);
nand U917 (N_917,N_338,N_282);
and U918 (N_918,N_60,N_386);
or U919 (N_919,N_154,N_70);
and U920 (N_920,N_46,N_93);
or U921 (N_921,N_219,N_277);
or U922 (N_922,N_48,N_475);
nand U923 (N_923,N_227,N_470);
or U924 (N_924,N_239,N_140);
nand U925 (N_925,N_30,N_442);
and U926 (N_926,N_311,N_342);
xnor U927 (N_927,N_170,N_429);
or U928 (N_928,N_300,N_281);
nor U929 (N_929,N_209,N_196);
and U930 (N_930,N_388,N_169);
and U931 (N_931,N_45,N_170);
nor U932 (N_932,N_327,N_26);
and U933 (N_933,N_45,N_370);
nor U934 (N_934,N_373,N_8);
nand U935 (N_935,N_296,N_319);
nor U936 (N_936,N_86,N_317);
and U937 (N_937,N_482,N_207);
nand U938 (N_938,N_313,N_426);
and U939 (N_939,N_257,N_153);
nand U940 (N_940,N_245,N_40);
and U941 (N_941,N_173,N_141);
or U942 (N_942,N_32,N_28);
nand U943 (N_943,N_98,N_241);
or U944 (N_944,N_273,N_223);
nand U945 (N_945,N_6,N_354);
nand U946 (N_946,N_321,N_492);
and U947 (N_947,N_472,N_341);
and U948 (N_948,N_73,N_115);
nor U949 (N_949,N_86,N_343);
and U950 (N_950,N_442,N_432);
and U951 (N_951,N_109,N_227);
nand U952 (N_952,N_187,N_455);
or U953 (N_953,N_147,N_397);
nand U954 (N_954,N_272,N_476);
nand U955 (N_955,N_89,N_117);
or U956 (N_956,N_160,N_405);
or U957 (N_957,N_481,N_491);
and U958 (N_958,N_240,N_411);
nor U959 (N_959,N_29,N_35);
nor U960 (N_960,N_446,N_232);
or U961 (N_961,N_475,N_320);
nor U962 (N_962,N_180,N_2);
and U963 (N_963,N_79,N_141);
or U964 (N_964,N_245,N_74);
and U965 (N_965,N_180,N_318);
nand U966 (N_966,N_374,N_178);
or U967 (N_967,N_27,N_245);
nor U968 (N_968,N_471,N_222);
nor U969 (N_969,N_263,N_222);
nand U970 (N_970,N_384,N_130);
or U971 (N_971,N_179,N_467);
nand U972 (N_972,N_339,N_106);
or U973 (N_973,N_481,N_289);
nand U974 (N_974,N_359,N_95);
nand U975 (N_975,N_225,N_4);
nand U976 (N_976,N_341,N_98);
nand U977 (N_977,N_465,N_491);
or U978 (N_978,N_110,N_177);
or U979 (N_979,N_307,N_210);
and U980 (N_980,N_194,N_156);
nor U981 (N_981,N_305,N_366);
nor U982 (N_982,N_218,N_420);
nor U983 (N_983,N_229,N_140);
or U984 (N_984,N_207,N_252);
or U985 (N_985,N_114,N_137);
and U986 (N_986,N_69,N_478);
nor U987 (N_987,N_81,N_456);
nand U988 (N_988,N_177,N_493);
and U989 (N_989,N_346,N_16);
nand U990 (N_990,N_287,N_389);
or U991 (N_991,N_420,N_262);
and U992 (N_992,N_248,N_424);
and U993 (N_993,N_473,N_9);
nand U994 (N_994,N_269,N_255);
nand U995 (N_995,N_315,N_20);
nand U996 (N_996,N_430,N_110);
xor U997 (N_997,N_305,N_83);
nand U998 (N_998,N_306,N_2);
nand U999 (N_999,N_375,N_205);
and U1000 (N_1000,N_943,N_692);
or U1001 (N_1001,N_578,N_851);
and U1002 (N_1002,N_574,N_678);
or U1003 (N_1003,N_765,N_741);
or U1004 (N_1004,N_637,N_800);
nand U1005 (N_1005,N_534,N_909);
nor U1006 (N_1006,N_702,N_693);
or U1007 (N_1007,N_840,N_973);
and U1008 (N_1008,N_616,N_756);
and U1009 (N_1009,N_597,N_661);
or U1010 (N_1010,N_872,N_532);
nor U1011 (N_1011,N_594,N_876);
or U1012 (N_1012,N_729,N_914);
nand U1013 (N_1013,N_605,N_975);
or U1014 (N_1014,N_844,N_648);
nor U1015 (N_1015,N_548,N_832);
and U1016 (N_1016,N_948,N_962);
nand U1017 (N_1017,N_697,N_645);
nor U1018 (N_1018,N_923,N_894);
nand U1019 (N_1019,N_576,N_720);
and U1020 (N_1020,N_768,N_682);
nand U1021 (N_1021,N_836,N_513);
nor U1022 (N_1022,N_989,N_842);
or U1023 (N_1023,N_683,N_618);
nor U1024 (N_1024,N_599,N_620);
nor U1025 (N_1025,N_520,N_514);
xor U1026 (N_1026,N_655,N_971);
nor U1027 (N_1027,N_603,N_503);
nor U1028 (N_1028,N_721,N_934);
or U1029 (N_1029,N_865,N_572);
nor U1030 (N_1030,N_992,N_788);
and U1031 (N_1031,N_970,N_560);
nor U1032 (N_1032,N_527,N_843);
and U1033 (N_1033,N_783,N_808);
and U1034 (N_1034,N_759,N_984);
or U1035 (N_1035,N_910,N_707);
nor U1036 (N_1036,N_554,N_859);
nor U1037 (N_1037,N_680,N_883);
xor U1038 (N_1038,N_536,N_977);
nand U1039 (N_1039,N_623,N_922);
nor U1040 (N_1040,N_807,N_966);
and U1041 (N_1041,N_608,N_588);
nand U1042 (N_1042,N_586,N_595);
or U1043 (N_1043,N_557,N_856);
or U1044 (N_1044,N_607,N_744);
nand U1045 (N_1045,N_545,N_521);
and U1046 (N_1046,N_695,N_945);
or U1047 (N_1047,N_619,N_689);
nor U1048 (N_1048,N_657,N_612);
or U1049 (N_1049,N_921,N_541);
nand U1050 (N_1050,N_562,N_946);
nand U1051 (N_1051,N_954,N_858);
or U1052 (N_1052,N_801,N_860);
nand U1053 (N_1053,N_906,N_955);
and U1054 (N_1054,N_979,N_627);
or U1055 (N_1055,N_867,N_929);
nand U1056 (N_1056,N_990,N_714);
nand U1057 (N_1057,N_863,N_820);
or U1058 (N_1058,N_677,N_630);
or U1059 (N_1059,N_877,N_811);
nor U1060 (N_1060,N_500,N_584);
nand U1061 (N_1061,N_747,N_804);
nand U1062 (N_1062,N_559,N_717);
nand U1063 (N_1063,N_512,N_806);
and U1064 (N_1064,N_932,N_999);
nand U1065 (N_1065,N_930,N_543);
or U1066 (N_1066,N_882,N_571);
or U1067 (N_1067,N_972,N_861);
nand U1068 (N_1068,N_901,N_838);
nand U1069 (N_1069,N_740,N_902);
and U1070 (N_1070,N_722,N_937);
nand U1071 (N_1071,N_666,N_896);
nor U1072 (N_1072,N_868,N_596);
and U1073 (N_1073,N_665,N_508);
nand U1074 (N_1074,N_862,N_736);
or U1075 (N_1075,N_748,N_938);
nand U1076 (N_1076,N_815,N_501);
nor U1077 (N_1077,N_950,N_887);
nor U1078 (N_1078,N_542,N_924);
nand U1079 (N_1079,N_685,N_864);
nand U1080 (N_1080,N_684,N_530);
nor U1081 (N_1081,N_763,N_725);
or U1082 (N_1082,N_647,N_994);
nor U1083 (N_1083,N_825,N_770);
nor U1084 (N_1084,N_715,N_538);
nand U1085 (N_1085,N_517,N_790);
nand U1086 (N_1086,N_651,N_964);
or U1087 (N_1087,N_944,N_587);
or U1088 (N_1088,N_591,N_658);
nand U1089 (N_1089,N_733,N_749);
or U1090 (N_1090,N_564,N_762);
and U1091 (N_1091,N_956,N_886);
nand U1092 (N_1092,N_731,N_670);
nor U1093 (N_1093,N_789,N_505);
nor U1094 (N_1094,N_598,N_660);
nor U1095 (N_1095,N_617,N_573);
nor U1096 (N_1096,N_813,N_656);
nor U1097 (N_1097,N_539,N_986);
and U1098 (N_1098,N_752,N_643);
nor U1099 (N_1099,N_734,N_687);
or U1100 (N_1100,N_965,N_775);
nand U1101 (N_1101,N_787,N_719);
nor U1102 (N_1102,N_751,N_933);
nand U1103 (N_1103,N_679,N_766);
and U1104 (N_1104,N_526,N_590);
and U1105 (N_1105,N_985,N_976);
nor U1106 (N_1106,N_614,N_940);
or U1107 (N_1107,N_515,N_609);
nor U1108 (N_1108,N_926,N_919);
and U1109 (N_1109,N_593,N_529);
and U1110 (N_1110,N_848,N_502);
nor U1111 (N_1111,N_793,N_908);
or U1112 (N_1112,N_925,N_604);
nor U1113 (N_1113,N_664,N_662);
or U1114 (N_1114,N_738,N_935);
nor U1115 (N_1115,N_897,N_852);
nand U1116 (N_1116,N_889,N_646);
xnor U1117 (N_1117,N_668,N_761);
nand U1118 (N_1118,N_869,N_960);
nand U1119 (N_1119,N_931,N_803);
nor U1120 (N_1120,N_784,N_785);
and U1121 (N_1121,N_633,N_703);
and U1122 (N_1122,N_780,N_892);
nand U1123 (N_1123,N_760,N_581);
and U1124 (N_1124,N_525,N_589);
and U1125 (N_1125,N_511,N_899);
nand U1126 (N_1126,N_575,N_953);
and U1127 (N_1127,N_639,N_621);
nand U1128 (N_1128,N_917,N_568);
nor U1129 (N_1129,N_654,N_839);
nand U1130 (N_1130,N_528,N_735);
and U1131 (N_1131,N_730,N_957);
and U1132 (N_1132,N_822,N_750);
or U1133 (N_1133,N_905,N_968);
and U1134 (N_1134,N_516,N_847);
and U1135 (N_1135,N_628,N_712);
and U1136 (N_1136,N_846,N_629);
and U1137 (N_1137,N_533,N_767);
and U1138 (N_1138,N_831,N_890);
nor U1139 (N_1139,N_509,N_708);
or U1140 (N_1140,N_546,N_879);
nand U1141 (N_1141,N_757,N_563);
nand U1142 (N_1142,N_829,N_833);
nand U1143 (N_1143,N_998,N_995);
nor U1144 (N_1144,N_540,N_510);
or U1145 (N_1145,N_958,N_911);
or U1146 (N_1146,N_531,N_981);
nand U1147 (N_1147,N_853,N_936);
nor U1148 (N_1148,N_795,N_653);
and U1149 (N_1149,N_522,N_781);
nor U1150 (N_1150,N_786,N_916);
or U1151 (N_1151,N_942,N_737);
nor U1152 (N_1152,N_898,N_710);
nand U1153 (N_1153,N_828,N_772);
nand U1154 (N_1154,N_967,N_812);
nor U1155 (N_1155,N_506,N_728);
or U1156 (N_1156,N_727,N_773);
nor U1157 (N_1157,N_570,N_724);
and U1158 (N_1158,N_866,N_821);
or U1159 (N_1159,N_652,N_997);
nor U1160 (N_1160,N_732,N_739);
nor U1161 (N_1161,N_798,N_993);
nor U1162 (N_1162,N_547,N_706);
and U1163 (N_1163,N_817,N_939);
nor U1164 (N_1164,N_704,N_947);
nand U1165 (N_1165,N_871,N_686);
or U1166 (N_1166,N_927,N_711);
or U1167 (N_1167,N_602,N_814);
or U1168 (N_1168,N_754,N_850);
and U1169 (N_1169,N_673,N_777);
nor U1170 (N_1170,N_636,N_907);
nand U1171 (N_1171,N_555,N_941);
nand U1172 (N_1172,N_870,N_726);
nand U1173 (N_1173,N_561,N_891);
or U1174 (N_1174,N_663,N_782);
or U1175 (N_1175,N_791,N_904);
nand U1176 (N_1176,N_745,N_582);
nand U1177 (N_1177,N_794,N_600);
or U1178 (N_1178,N_885,N_895);
and U1179 (N_1179,N_649,N_606);
xor U1180 (N_1180,N_792,N_912);
nand U1181 (N_1181,N_857,N_524);
nand U1182 (N_1182,N_699,N_718);
or U1183 (N_1183,N_830,N_688);
or U1184 (N_1184,N_552,N_625);
nand U1185 (N_1185,N_816,N_613);
or U1186 (N_1186,N_996,N_746);
nor U1187 (N_1187,N_713,N_928);
and U1188 (N_1188,N_963,N_802);
or U1189 (N_1189,N_796,N_676);
and U1190 (N_1190,N_799,N_983);
and U1191 (N_1191,N_974,N_881);
and U1192 (N_1192,N_826,N_626);
nor U1193 (N_1193,N_553,N_631);
nor U1194 (N_1194,N_650,N_583);
nor U1195 (N_1195,N_674,N_615);
nor U1196 (N_1196,N_638,N_873);
or U1197 (N_1197,N_837,N_519);
or U1198 (N_1198,N_982,N_961);
and U1199 (N_1199,N_959,N_819);
nor U1200 (N_1200,N_742,N_690);
and U1201 (N_1201,N_698,N_888);
and U1202 (N_1202,N_507,N_980);
nor U1203 (N_1203,N_949,N_523);
nor U1204 (N_1204,N_878,N_827);
nand U1205 (N_1205,N_567,N_755);
nor U1206 (N_1206,N_854,N_743);
or U1207 (N_1207,N_709,N_841);
xnor U1208 (N_1208,N_913,N_566);
or U1209 (N_1209,N_809,N_810);
nor U1210 (N_1210,N_544,N_805);
and U1211 (N_1211,N_558,N_622);
or U1212 (N_1212,N_978,N_644);
or U1213 (N_1213,N_969,N_705);
nor U1214 (N_1214,N_556,N_580);
nor U1215 (N_1215,N_610,N_669);
nor U1216 (N_1216,N_701,N_642);
or U1217 (N_1217,N_504,N_880);
nand U1218 (N_1218,N_824,N_634);
and U1219 (N_1219,N_845,N_797);
xor U1220 (N_1220,N_550,N_835);
or U1221 (N_1221,N_641,N_700);
nand U1222 (N_1222,N_691,N_640);
nor U1223 (N_1223,N_535,N_778);
nand U1224 (N_1224,N_549,N_551);
nand U1225 (N_1225,N_694,N_987);
nand U1226 (N_1226,N_771,N_834);
nand U1227 (N_1227,N_874,N_758);
or U1228 (N_1228,N_723,N_875);
or U1229 (N_1229,N_920,N_818);
nor U1230 (N_1230,N_681,N_624);
nand U1231 (N_1231,N_915,N_672);
nor U1232 (N_1232,N_537,N_779);
nor U1233 (N_1233,N_764,N_952);
nor U1234 (N_1234,N_823,N_585);
nor U1235 (N_1235,N_577,N_855);
and U1236 (N_1236,N_918,N_776);
nand U1237 (N_1237,N_659,N_579);
or U1238 (N_1238,N_716,N_667);
or U1239 (N_1239,N_671,N_601);
and U1240 (N_1240,N_753,N_903);
nor U1241 (N_1241,N_592,N_696);
nor U1242 (N_1242,N_569,N_884);
nor U1243 (N_1243,N_951,N_991);
or U1244 (N_1244,N_988,N_518);
or U1245 (N_1245,N_675,N_611);
or U1246 (N_1246,N_849,N_893);
or U1247 (N_1247,N_900,N_565);
or U1248 (N_1248,N_635,N_769);
nand U1249 (N_1249,N_774,N_632);
nor U1250 (N_1250,N_588,N_688);
nand U1251 (N_1251,N_886,N_537);
nand U1252 (N_1252,N_601,N_626);
and U1253 (N_1253,N_865,N_634);
or U1254 (N_1254,N_673,N_771);
nand U1255 (N_1255,N_881,N_859);
or U1256 (N_1256,N_850,N_941);
nor U1257 (N_1257,N_638,N_634);
and U1258 (N_1258,N_644,N_805);
xnor U1259 (N_1259,N_977,N_553);
nor U1260 (N_1260,N_928,N_740);
or U1261 (N_1261,N_736,N_987);
nand U1262 (N_1262,N_786,N_562);
nand U1263 (N_1263,N_896,N_980);
nand U1264 (N_1264,N_895,N_508);
and U1265 (N_1265,N_554,N_991);
and U1266 (N_1266,N_810,N_844);
and U1267 (N_1267,N_668,N_502);
or U1268 (N_1268,N_518,N_810);
nor U1269 (N_1269,N_661,N_888);
and U1270 (N_1270,N_748,N_644);
nor U1271 (N_1271,N_994,N_851);
or U1272 (N_1272,N_545,N_705);
and U1273 (N_1273,N_925,N_626);
nor U1274 (N_1274,N_846,N_698);
nand U1275 (N_1275,N_838,N_703);
nand U1276 (N_1276,N_977,N_974);
or U1277 (N_1277,N_508,N_877);
or U1278 (N_1278,N_771,N_691);
nor U1279 (N_1279,N_828,N_762);
nand U1280 (N_1280,N_874,N_811);
nor U1281 (N_1281,N_615,N_809);
or U1282 (N_1282,N_804,N_512);
and U1283 (N_1283,N_632,N_976);
nand U1284 (N_1284,N_816,N_622);
or U1285 (N_1285,N_739,N_553);
and U1286 (N_1286,N_752,N_571);
or U1287 (N_1287,N_527,N_592);
or U1288 (N_1288,N_620,N_724);
nor U1289 (N_1289,N_711,N_760);
nor U1290 (N_1290,N_758,N_998);
and U1291 (N_1291,N_948,N_513);
nor U1292 (N_1292,N_821,N_891);
nor U1293 (N_1293,N_946,N_880);
or U1294 (N_1294,N_730,N_603);
nand U1295 (N_1295,N_712,N_964);
nor U1296 (N_1296,N_696,N_787);
nor U1297 (N_1297,N_853,N_509);
or U1298 (N_1298,N_997,N_841);
nand U1299 (N_1299,N_634,N_775);
nor U1300 (N_1300,N_806,N_902);
or U1301 (N_1301,N_723,N_705);
and U1302 (N_1302,N_960,N_741);
and U1303 (N_1303,N_736,N_630);
nand U1304 (N_1304,N_793,N_843);
nand U1305 (N_1305,N_619,N_573);
or U1306 (N_1306,N_727,N_956);
nand U1307 (N_1307,N_865,N_543);
nand U1308 (N_1308,N_770,N_913);
nand U1309 (N_1309,N_726,N_565);
nand U1310 (N_1310,N_604,N_576);
or U1311 (N_1311,N_822,N_574);
nor U1312 (N_1312,N_914,N_980);
and U1313 (N_1313,N_720,N_617);
and U1314 (N_1314,N_576,N_848);
nand U1315 (N_1315,N_692,N_823);
and U1316 (N_1316,N_688,N_617);
or U1317 (N_1317,N_985,N_559);
nor U1318 (N_1318,N_903,N_625);
and U1319 (N_1319,N_664,N_959);
or U1320 (N_1320,N_637,N_680);
nor U1321 (N_1321,N_581,N_997);
or U1322 (N_1322,N_880,N_839);
and U1323 (N_1323,N_516,N_594);
nand U1324 (N_1324,N_696,N_861);
nand U1325 (N_1325,N_889,N_987);
nor U1326 (N_1326,N_780,N_717);
or U1327 (N_1327,N_759,N_617);
or U1328 (N_1328,N_552,N_528);
nand U1329 (N_1329,N_539,N_975);
or U1330 (N_1330,N_918,N_739);
and U1331 (N_1331,N_777,N_596);
nand U1332 (N_1332,N_772,N_524);
nand U1333 (N_1333,N_759,N_640);
nor U1334 (N_1334,N_620,N_574);
nor U1335 (N_1335,N_652,N_694);
or U1336 (N_1336,N_952,N_664);
and U1337 (N_1337,N_728,N_757);
and U1338 (N_1338,N_888,N_997);
or U1339 (N_1339,N_632,N_734);
and U1340 (N_1340,N_829,N_970);
xor U1341 (N_1341,N_701,N_685);
or U1342 (N_1342,N_947,N_970);
nand U1343 (N_1343,N_566,N_552);
nand U1344 (N_1344,N_576,N_842);
nor U1345 (N_1345,N_954,N_673);
and U1346 (N_1346,N_938,N_981);
nand U1347 (N_1347,N_936,N_901);
nand U1348 (N_1348,N_966,N_727);
and U1349 (N_1349,N_584,N_517);
nand U1350 (N_1350,N_945,N_561);
or U1351 (N_1351,N_597,N_523);
or U1352 (N_1352,N_681,N_762);
xnor U1353 (N_1353,N_603,N_936);
nor U1354 (N_1354,N_984,N_603);
or U1355 (N_1355,N_562,N_882);
or U1356 (N_1356,N_868,N_912);
and U1357 (N_1357,N_748,N_856);
nor U1358 (N_1358,N_854,N_800);
nor U1359 (N_1359,N_792,N_984);
and U1360 (N_1360,N_771,N_660);
nor U1361 (N_1361,N_967,N_902);
or U1362 (N_1362,N_959,N_928);
nor U1363 (N_1363,N_525,N_625);
and U1364 (N_1364,N_662,N_943);
and U1365 (N_1365,N_719,N_888);
nand U1366 (N_1366,N_606,N_926);
nor U1367 (N_1367,N_633,N_852);
nor U1368 (N_1368,N_699,N_856);
or U1369 (N_1369,N_572,N_712);
and U1370 (N_1370,N_654,N_619);
nor U1371 (N_1371,N_548,N_860);
or U1372 (N_1372,N_569,N_860);
and U1373 (N_1373,N_685,N_729);
nand U1374 (N_1374,N_731,N_513);
or U1375 (N_1375,N_704,N_745);
and U1376 (N_1376,N_639,N_997);
or U1377 (N_1377,N_722,N_591);
nand U1378 (N_1378,N_864,N_840);
nand U1379 (N_1379,N_852,N_862);
nand U1380 (N_1380,N_677,N_610);
and U1381 (N_1381,N_867,N_574);
nor U1382 (N_1382,N_788,N_566);
nand U1383 (N_1383,N_908,N_844);
and U1384 (N_1384,N_953,N_577);
or U1385 (N_1385,N_669,N_784);
nor U1386 (N_1386,N_774,N_924);
or U1387 (N_1387,N_567,N_728);
nand U1388 (N_1388,N_751,N_871);
and U1389 (N_1389,N_525,N_730);
nor U1390 (N_1390,N_694,N_692);
nand U1391 (N_1391,N_915,N_963);
nand U1392 (N_1392,N_723,N_623);
and U1393 (N_1393,N_697,N_859);
or U1394 (N_1394,N_539,N_812);
nor U1395 (N_1395,N_646,N_680);
or U1396 (N_1396,N_914,N_678);
nand U1397 (N_1397,N_866,N_621);
or U1398 (N_1398,N_531,N_859);
nor U1399 (N_1399,N_947,N_628);
nor U1400 (N_1400,N_694,N_586);
or U1401 (N_1401,N_799,N_989);
and U1402 (N_1402,N_717,N_612);
nand U1403 (N_1403,N_552,N_610);
nor U1404 (N_1404,N_841,N_666);
and U1405 (N_1405,N_505,N_868);
or U1406 (N_1406,N_973,N_827);
or U1407 (N_1407,N_950,N_569);
nor U1408 (N_1408,N_872,N_701);
and U1409 (N_1409,N_665,N_869);
nand U1410 (N_1410,N_986,N_938);
nor U1411 (N_1411,N_507,N_993);
nand U1412 (N_1412,N_929,N_944);
nand U1413 (N_1413,N_661,N_939);
or U1414 (N_1414,N_525,N_964);
or U1415 (N_1415,N_576,N_668);
or U1416 (N_1416,N_658,N_726);
and U1417 (N_1417,N_886,N_599);
nor U1418 (N_1418,N_725,N_864);
or U1419 (N_1419,N_710,N_560);
or U1420 (N_1420,N_915,N_577);
and U1421 (N_1421,N_592,N_732);
nand U1422 (N_1422,N_972,N_771);
and U1423 (N_1423,N_678,N_949);
and U1424 (N_1424,N_837,N_679);
nand U1425 (N_1425,N_629,N_808);
and U1426 (N_1426,N_731,N_869);
nor U1427 (N_1427,N_873,N_785);
or U1428 (N_1428,N_954,N_500);
and U1429 (N_1429,N_908,N_942);
or U1430 (N_1430,N_506,N_842);
nor U1431 (N_1431,N_670,N_546);
and U1432 (N_1432,N_634,N_845);
and U1433 (N_1433,N_981,N_831);
nand U1434 (N_1434,N_875,N_656);
nor U1435 (N_1435,N_743,N_542);
and U1436 (N_1436,N_672,N_515);
or U1437 (N_1437,N_558,N_510);
and U1438 (N_1438,N_645,N_922);
and U1439 (N_1439,N_798,N_503);
and U1440 (N_1440,N_964,N_935);
and U1441 (N_1441,N_834,N_505);
or U1442 (N_1442,N_629,N_828);
and U1443 (N_1443,N_984,N_736);
nand U1444 (N_1444,N_540,N_770);
and U1445 (N_1445,N_838,N_663);
nor U1446 (N_1446,N_536,N_696);
and U1447 (N_1447,N_857,N_635);
nor U1448 (N_1448,N_865,N_870);
xor U1449 (N_1449,N_501,N_620);
nor U1450 (N_1450,N_875,N_516);
or U1451 (N_1451,N_609,N_809);
and U1452 (N_1452,N_931,N_701);
and U1453 (N_1453,N_590,N_735);
and U1454 (N_1454,N_507,N_835);
nor U1455 (N_1455,N_871,N_729);
nor U1456 (N_1456,N_781,N_697);
nor U1457 (N_1457,N_600,N_675);
or U1458 (N_1458,N_802,N_584);
or U1459 (N_1459,N_869,N_835);
nand U1460 (N_1460,N_512,N_552);
and U1461 (N_1461,N_793,N_730);
and U1462 (N_1462,N_686,N_602);
and U1463 (N_1463,N_997,N_847);
or U1464 (N_1464,N_810,N_788);
nand U1465 (N_1465,N_917,N_644);
nor U1466 (N_1466,N_768,N_950);
nand U1467 (N_1467,N_901,N_734);
nand U1468 (N_1468,N_901,N_849);
and U1469 (N_1469,N_788,N_653);
nor U1470 (N_1470,N_865,N_755);
or U1471 (N_1471,N_542,N_555);
xor U1472 (N_1472,N_813,N_629);
nand U1473 (N_1473,N_557,N_764);
or U1474 (N_1474,N_666,N_969);
or U1475 (N_1475,N_578,N_919);
nor U1476 (N_1476,N_710,N_816);
nor U1477 (N_1477,N_674,N_633);
or U1478 (N_1478,N_516,N_651);
and U1479 (N_1479,N_528,N_602);
xnor U1480 (N_1480,N_810,N_531);
nand U1481 (N_1481,N_878,N_805);
or U1482 (N_1482,N_828,N_616);
and U1483 (N_1483,N_821,N_714);
nor U1484 (N_1484,N_691,N_774);
or U1485 (N_1485,N_979,N_701);
or U1486 (N_1486,N_720,N_851);
and U1487 (N_1487,N_875,N_789);
nor U1488 (N_1488,N_594,N_591);
nor U1489 (N_1489,N_534,N_613);
nor U1490 (N_1490,N_986,N_712);
nand U1491 (N_1491,N_915,N_779);
nand U1492 (N_1492,N_786,N_972);
and U1493 (N_1493,N_734,N_761);
nand U1494 (N_1494,N_633,N_988);
nand U1495 (N_1495,N_963,N_546);
nand U1496 (N_1496,N_965,N_581);
or U1497 (N_1497,N_733,N_731);
nand U1498 (N_1498,N_863,N_990);
and U1499 (N_1499,N_934,N_557);
and U1500 (N_1500,N_1194,N_1346);
nand U1501 (N_1501,N_1487,N_1328);
nor U1502 (N_1502,N_1127,N_1455);
and U1503 (N_1503,N_1089,N_1313);
nand U1504 (N_1504,N_1415,N_1104);
nor U1505 (N_1505,N_1460,N_1097);
and U1506 (N_1506,N_1279,N_1249);
nor U1507 (N_1507,N_1491,N_1014);
or U1508 (N_1508,N_1190,N_1137);
nand U1509 (N_1509,N_1217,N_1065);
or U1510 (N_1510,N_1475,N_1253);
and U1511 (N_1511,N_1111,N_1292);
or U1512 (N_1512,N_1411,N_1446);
or U1513 (N_1513,N_1096,N_1403);
nor U1514 (N_1514,N_1418,N_1353);
and U1515 (N_1515,N_1086,N_1185);
or U1516 (N_1516,N_1236,N_1494);
nand U1517 (N_1517,N_1126,N_1219);
nand U1518 (N_1518,N_1216,N_1283);
nor U1519 (N_1519,N_1492,N_1113);
and U1520 (N_1520,N_1360,N_1020);
nor U1521 (N_1521,N_1343,N_1178);
nor U1522 (N_1522,N_1076,N_1291);
nand U1523 (N_1523,N_1234,N_1183);
nor U1524 (N_1524,N_1468,N_1390);
nor U1525 (N_1525,N_1430,N_1409);
nor U1526 (N_1526,N_1429,N_1392);
nor U1527 (N_1527,N_1401,N_1123);
nor U1528 (N_1528,N_1196,N_1386);
and U1529 (N_1529,N_1237,N_1444);
nor U1530 (N_1530,N_1277,N_1458);
nor U1531 (N_1531,N_1477,N_1296);
nand U1532 (N_1532,N_1042,N_1263);
nor U1533 (N_1533,N_1110,N_1044);
nor U1534 (N_1534,N_1079,N_1136);
nor U1535 (N_1535,N_1266,N_1301);
or U1536 (N_1536,N_1319,N_1267);
and U1537 (N_1537,N_1469,N_1378);
nor U1538 (N_1538,N_1356,N_1214);
nor U1539 (N_1539,N_1471,N_1115);
or U1540 (N_1540,N_1256,N_1311);
nor U1541 (N_1541,N_1281,N_1348);
nand U1542 (N_1542,N_1399,N_1054);
nand U1543 (N_1543,N_1481,N_1226);
nand U1544 (N_1544,N_1410,N_1336);
and U1545 (N_1545,N_1149,N_1305);
and U1546 (N_1546,N_1182,N_1359);
or U1547 (N_1547,N_1252,N_1337);
nand U1548 (N_1548,N_1275,N_1206);
and U1549 (N_1549,N_1333,N_1048);
or U1550 (N_1550,N_1037,N_1141);
or U1551 (N_1551,N_1280,N_1327);
and U1552 (N_1552,N_1165,N_1445);
or U1553 (N_1553,N_1201,N_1091);
nor U1554 (N_1554,N_1131,N_1015);
and U1555 (N_1555,N_1187,N_1486);
or U1556 (N_1556,N_1189,N_1312);
or U1557 (N_1557,N_1405,N_1464);
nor U1558 (N_1558,N_1225,N_1254);
nand U1559 (N_1559,N_1140,N_1284);
nand U1560 (N_1560,N_1320,N_1240);
nor U1561 (N_1561,N_1478,N_1423);
nor U1562 (N_1562,N_1218,N_1022);
nand U1563 (N_1563,N_1151,N_1310);
nor U1564 (N_1564,N_1130,N_1035);
nor U1565 (N_1565,N_1422,N_1109);
and U1566 (N_1566,N_1294,N_1160);
nor U1567 (N_1567,N_1176,N_1461);
nand U1568 (N_1568,N_1424,N_1043);
nor U1569 (N_1569,N_1358,N_1023);
and U1570 (N_1570,N_1306,N_1457);
nand U1571 (N_1571,N_1456,N_1069);
nor U1572 (N_1572,N_1416,N_1102);
and U1573 (N_1573,N_1062,N_1395);
nand U1574 (N_1574,N_1350,N_1302);
or U1575 (N_1575,N_1146,N_1215);
nand U1576 (N_1576,N_1011,N_1125);
and U1577 (N_1577,N_1288,N_1352);
or U1578 (N_1578,N_1195,N_1051);
nand U1579 (N_1579,N_1078,N_1421);
nand U1580 (N_1580,N_1332,N_1036);
and U1581 (N_1581,N_1060,N_1384);
nor U1582 (N_1582,N_1393,N_1066);
and U1583 (N_1583,N_1150,N_1070);
nor U1584 (N_1584,N_1479,N_1171);
nor U1585 (N_1585,N_1370,N_1056);
or U1586 (N_1586,N_1166,N_1309);
and U1587 (N_1587,N_1064,N_1412);
nor U1588 (N_1588,N_1221,N_1318);
and U1589 (N_1589,N_1453,N_1307);
nor U1590 (N_1590,N_1139,N_1326);
nor U1591 (N_1591,N_1483,N_1147);
nand U1592 (N_1592,N_1268,N_1255);
and U1593 (N_1593,N_1003,N_1324);
and U1594 (N_1594,N_1466,N_1321);
or U1595 (N_1595,N_1260,N_1282);
nor U1596 (N_1596,N_1028,N_1055);
nor U1597 (N_1597,N_1013,N_1278);
nand U1598 (N_1598,N_1114,N_1442);
or U1599 (N_1599,N_1230,N_1400);
and U1600 (N_1600,N_1335,N_1007);
nor U1601 (N_1601,N_1026,N_1357);
nand U1602 (N_1602,N_1027,N_1362);
nand U1603 (N_1603,N_1205,N_1168);
and U1604 (N_1604,N_1454,N_1375);
or U1605 (N_1605,N_1372,N_1222);
and U1606 (N_1606,N_1046,N_1231);
or U1607 (N_1607,N_1059,N_1385);
nand U1608 (N_1608,N_1024,N_1116);
nand U1609 (N_1609,N_1239,N_1315);
or U1610 (N_1610,N_1404,N_1298);
and U1611 (N_1611,N_1068,N_1467);
and U1612 (N_1612,N_1001,N_1170);
nor U1613 (N_1613,N_1261,N_1413);
and U1614 (N_1614,N_1379,N_1241);
or U1615 (N_1615,N_1476,N_1490);
nand U1616 (N_1616,N_1163,N_1374);
and U1617 (N_1617,N_1145,N_1247);
nand U1618 (N_1618,N_1016,N_1088);
nand U1619 (N_1619,N_1224,N_1355);
or U1620 (N_1620,N_1197,N_1174);
and U1621 (N_1621,N_1159,N_1387);
or U1622 (N_1622,N_1199,N_1331);
and U1623 (N_1623,N_1200,N_1019);
or U1624 (N_1624,N_1175,N_1057);
and U1625 (N_1625,N_1484,N_1351);
nand U1626 (N_1626,N_1329,N_1128);
or U1627 (N_1627,N_1269,N_1153);
or U1628 (N_1628,N_1244,N_1246);
nor U1629 (N_1629,N_1106,N_1207);
and U1630 (N_1630,N_1155,N_1427);
nand U1631 (N_1631,N_1010,N_1039);
nand U1632 (N_1632,N_1095,N_1245);
or U1633 (N_1633,N_1052,N_1432);
nor U1634 (N_1634,N_1474,N_1090);
nor U1635 (N_1635,N_1154,N_1377);
nor U1636 (N_1636,N_1167,N_1496);
and U1637 (N_1637,N_1080,N_1450);
nand U1638 (N_1638,N_1488,N_1363);
and U1639 (N_1639,N_1323,N_1041);
or U1640 (N_1640,N_1220,N_1050);
nand U1641 (N_1641,N_1135,N_1193);
or U1642 (N_1642,N_1138,N_1472);
nor U1643 (N_1643,N_1436,N_1417);
or U1644 (N_1644,N_1349,N_1152);
and U1645 (N_1645,N_1473,N_1124);
and U1646 (N_1646,N_1021,N_1162);
nand U1647 (N_1647,N_1232,N_1173);
nand U1648 (N_1648,N_1265,N_1184);
and U1649 (N_1649,N_1045,N_1361);
nor U1650 (N_1650,N_1286,N_1434);
or U1651 (N_1651,N_1148,N_1383);
nand U1652 (N_1652,N_1463,N_1177);
or U1653 (N_1653,N_1497,N_1293);
and U1654 (N_1654,N_1408,N_1388);
and U1655 (N_1655,N_1025,N_1227);
nand U1656 (N_1656,N_1164,N_1376);
and U1657 (N_1657,N_1299,N_1002);
and U1658 (N_1658,N_1258,N_1105);
xnor U1659 (N_1659,N_1061,N_1264);
and U1660 (N_1660,N_1158,N_1420);
nor U1661 (N_1661,N_1005,N_1017);
nor U1662 (N_1662,N_1303,N_1493);
nor U1663 (N_1663,N_1325,N_1081);
nor U1664 (N_1664,N_1047,N_1276);
nand U1665 (N_1665,N_1074,N_1391);
nand U1666 (N_1666,N_1287,N_1233);
or U1667 (N_1667,N_1439,N_1438);
and U1668 (N_1668,N_1181,N_1248);
and U1669 (N_1669,N_1431,N_1203);
nor U1670 (N_1670,N_1489,N_1314);
or U1671 (N_1671,N_1373,N_1053);
or U1672 (N_1672,N_1270,N_1228);
nand U1673 (N_1673,N_1364,N_1397);
and U1674 (N_1674,N_1103,N_1330);
nand U1675 (N_1675,N_1202,N_1449);
nor U1676 (N_1676,N_1122,N_1440);
or U1677 (N_1677,N_1212,N_1414);
nand U1678 (N_1678,N_1188,N_1006);
and U1679 (N_1679,N_1441,N_1425);
nor U1680 (N_1680,N_1443,N_1129);
or U1681 (N_1681,N_1134,N_1008);
or U1682 (N_1682,N_1398,N_1304);
and U1683 (N_1683,N_1000,N_1119);
and U1684 (N_1684,N_1480,N_1085);
nand U1685 (N_1685,N_1100,N_1034);
nor U1686 (N_1686,N_1428,N_1342);
nor U1687 (N_1687,N_1345,N_1300);
or U1688 (N_1688,N_1251,N_1334);
nand U1689 (N_1689,N_1208,N_1009);
nor U1690 (N_1690,N_1067,N_1072);
nor U1691 (N_1691,N_1098,N_1108);
nand U1692 (N_1692,N_1213,N_1250);
nor U1693 (N_1693,N_1172,N_1368);
xnor U1694 (N_1694,N_1465,N_1344);
nor U1695 (N_1695,N_1426,N_1262);
nor U1696 (N_1696,N_1031,N_1093);
or U1697 (N_1697,N_1406,N_1180);
and U1698 (N_1698,N_1243,N_1082);
and U1699 (N_1699,N_1448,N_1144);
nor U1700 (N_1700,N_1257,N_1308);
and U1701 (N_1701,N_1075,N_1101);
nand U1702 (N_1702,N_1092,N_1118);
nor U1703 (N_1703,N_1132,N_1317);
nor U1704 (N_1704,N_1340,N_1133);
nor U1705 (N_1705,N_1143,N_1482);
and U1706 (N_1706,N_1402,N_1198);
nand U1707 (N_1707,N_1462,N_1419);
xor U1708 (N_1708,N_1030,N_1107);
and U1709 (N_1709,N_1459,N_1367);
and U1710 (N_1710,N_1380,N_1274);
nand U1711 (N_1711,N_1338,N_1447);
and U1712 (N_1712,N_1433,N_1087);
and U1713 (N_1713,N_1407,N_1499);
nand U1714 (N_1714,N_1366,N_1238);
nand U1715 (N_1715,N_1211,N_1396);
or U1716 (N_1716,N_1365,N_1322);
nor U1717 (N_1717,N_1120,N_1077);
nor U1718 (N_1718,N_1084,N_1142);
nor U1719 (N_1719,N_1049,N_1371);
nand U1720 (N_1720,N_1316,N_1192);
nand U1721 (N_1721,N_1495,N_1191);
nor U1722 (N_1722,N_1210,N_1223);
and U1723 (N_1723,N_1381,N_1354);
nand U1724 (N_1724,N_1169,N_1451);
and U1725 (N_1725,N_1290,N_1485);
nor U1726 (N_1726,N_1112,N_1121);
nand U1727 (N_1727,N_1285,N_1452);
and U1728 (N_1728,N_1229,N_1038);
nor U1729 (N_1729,N_1209,N_1063);
nor U1730 (N_1730,N_1179,N_1339);
nand U1731 (N_1731,N_1437,N_1004);
nand U1732 (N_1732,N_1295,N_1094);
or U1733 (N_1733,N_1341,N_1271);
or U1734 (N_1734,N_1156,N_1117);
or U1735 (N_1735,N_1297,N_1204);
nand U1736 (N_1736,N_1032,N_1498);
nor U1737 (N_1737,N_1040,N_1369);
nand U1738 (N_1738,N_1289,N_1029);
nand U1739 (N_1739,N_1012,N_1235);
nor U1740 (N_1740,N_1099,N_1259);
and U1741 (N_1741,N_1033,N_1347);
and U1742 (N_1742,N_1161,N_1058);
and U1743 (N_1743,N_1389,N_1073);
or U1744 (N_1744,N_1083,N_1242);
xnor U1745 (N_1745,N_1157,N_1273);
nand U1746 (N_1746,N_1272,N_1470);
nor U1747 (N_1747,N_1394,N_1435);
and U1748 (N_1748,N_1382,N_1018);
nand U1749 (N_1749,N_1186,N_1071);
or U1750 (N_1750,N_1058,N_1276);
and U1751 (N_1751,N_1165,N_1461);
and U1752 (N_1752,N_1478,N_1029);
nand U1753 (N_1753,N_1216,N_1096);
and U1754 (N_1754,N_1384,N_1429);
or U1755 (N_1755,N_1474,N_1222);
nand U1756 (N_1756,N_1158,N_1173);
nor U1757 (N_1757,N_1295,N_1451);
nor U1758 (N_1758,N_1178,N_1220);
nor U1759 (N_1759,N_1150,N_1196);
nand U1760 (N_1760,N_1441,N_1448);
nand U1761 (N_1761,N_1253,N_1299);
nand U1762 (N_1762,N_1008,N_1193);
nand U1763 (N_1763,N_1281,N_1162);
nand U1764 (N_1764,N_1066,N_1315);
nand U1765 (N_1765,N_1404,N_1286);
nand U1766 (N_1766,N_1157,N_1147);
nand U1767 (N_1767,N_1210,N_1043);
nor U1768 (N_1768,N_1307,N_1368);
and U1769 (N_1769,N_1489,N_1026);
nor U1770 (N_1770,N_1016,N_1498);
nor U1771 (N_1771,N_1290,N_1021);
nor U1772 (N_1772,N_1337,N_1113);
nor U1773 (N_1773,N_1221,N_1414);
and U1774 (N_1774,N_1459,N_1113);
or U1775 (N_1775,N_1142,N_1292);
and U1776 (N_1776,N_1082,N_1406);
nand U1777 (N_1777,N_1405,N_1121);
and U1778 (N_1778,N_1237,N_1396);
and U1779 (N_1779,N_1388,N_1447);
nand U1780 (N_1780,N_1487,N_1258);
nand U1781 (N_1781,N_1314,N_1317);
nand U1782 (N_1782,N_1125,N_1220);
nor U1783 (N_1783,N_1005,N_1343);
nand U1784 (N_1784,N_1308,N_1231);
nand U1785 (N_1785,N_1166,N_1213);
and U1786 (N_1786,N_1363,N_1151);
nand U1787 (N_1787,N_1221,N_1350);
nand U1788 (N_1788,N_1110,N_1273);
and U1789 (N_1789,N_1429,N_1368);
or U1790 (N_1790,N_1067,N_1236);
nor U1791 (N_1791,N_1441,N_1239);
and U1792 (N_1792,N_1258,N_1337);
or U1793 (N_1793,N_1498,N_1345);
or U1794 (N_1794,N_1247,N_1466);
or U1795 (N_1795,N_1047,N_1004);
nor U1796 (N_1796,N_1028,N_1470);
nand U1797 (N_1797,N_1399,N_1329);
nor U1798 (N_1798,N_1254,N_1296);
and U1799 (N_1799,N_1267,N_1111);
nand U1800 (N_1800,N_1021,N_1042);
and U1801 (N_1801,N_1275,N_1154);
and U1802 (N_1802,N_1140,N_1384);
or U1803 (N_1803,N_1201,N_1372);
and U1804 (N_1804,N_1080,N_1019);
nand U1805 (N_1805,N_1108,N_1186);
nor U1806 (N_1806,N_1308,N_1394);
or U1807 (N_1807,N_1349,N_1305);
nand U1808 (N_1808,N_1397,N_1360);
or U1809 (N_1809,N_1044,N_1116);
xnor U1810 (N_1810,N_1327,N_1256);
nand U1811 (N_1811,N_1042,N_1009);
or U1812 (N_1812,N_1018,N_1194);
or U1813 (N_1813,N_1345,N_1476);
nand U1814 (N_1814,N_1296,N_1475);
xor U1815 (N_1815,N_1124,N_1260);
or U1816 (N_1816,N_1345,N_1354);
xor U1817 (N_1817,N_1246,N_1201);
and U1818 (N_1818,N_1377,N_1172);
nand U1819 (N_1819,N_1152,N_1388);
and U1820 (N_1820,N_1217,N_1295);
and U1821 (N_1821,N_1183,N_1240);
nor U1822 (N_1822,N_1153,N_1353);
nand U1823 (N_1823,N_1389,N_1067);
nor U1824 (N_1824,N_1408,N_1267);
or U1825 (N_1825,N_1253,N_1474);
nand U1826 (N_1826,N_1179,N_1004);
nand U1827 (N_1827,N_1012,N_1129);
nor U1828 (N_1828,N_1383,N_1394);
or U1829 (N_1829,N_1407,N_1130);
nand U1830 (N_1830,N_1446,N_1205);
nor U1831 (N_1831,N_1300,N_1413);
nand U1832 (N_1832,N_1219,N_1265);
nand U1833 (N_1833,N_1149,N_1142);
nand U1834 (N_1834,N_1047,N_1052);
nand U1835 (N_1835,N_1346,N_1018);
nor U1836 (N_1836,N_1376,N_1408);
nor U1837 (N_1837,N_1347,N_1373);
and U1838 (N_1838,N_1088,N_1058);
and U1839 (N_1839,N_1368,N_1147);
and U1840 (N_1840,N_1417,N_1406);
or U1841 (N_1841,N_1116,N_1495);
and U1842 (N_1842,N_1133,N_1400);
or U1843 (N_1843,N_1125,N_1341);
nand U1844 (N_1844,N_1441,N_1265);
nand U1845 (N_1845,N_1493,N_1294);
or U1846 (N_1846,N_1131,N_1381);
nor U1847 (N_1847,N_1224,N_1274);
and U1848 (N_1848,N_1077,N_1494);
nor U1849 (N_1849,N_1346,N_1307);
nand U1850 (N_1850,N_1025,N_1206);
nand U1851 (N_1851,N_1160,N_1244);
nand U1852 (N_1852,N_1125,N_1359);
and U1853 (N_1853,N_1239,N_1229);
nand U1854 (N_1854,N_1166,N_1319);
nand U1855 (N_1855,N_1446,N_1123);
and U1856 (N_1856,N_1038,N_1230);
or U1857 (N_1857,N_1049,N_1041);
nand U1858 (N_1858,N_1070,N_1170);
and U1859 (N_1859,N_1232,N_1322);
and U1860 (N_1860,N_1387,N_1115);
nor U1861 (N_1861,N_1352,N_1024);
nor U1862 (N_1862,N_1428,N_1373);
and U1863 (N_1863,N_1214,N_1038);
and U1864 (N_1864,N_1001,N_1408);
nand U1865 (N_1865,N_1413,N_1390);
and U1866 (N_1866,N_1379,N_1454);
and U1867 (N_1867,N_1479,N_1397);
or U1868 (N_1868,N_1195,N_1268);
nor U1869 (N_1869,N_1007,N_1357);
and U1870 (N_1870,N_1319,N_1088);
nand U1871 (N_1871,N_1018,N_1057);
nand U1872 (N_1872,N_1325,N_1204);
xor U1873 (N_1873,N_1161,N_1229);
and U1874 (N_1874,N_1179,N_1151);
and U1875 (N_1875,N_1113,N_1433);
or U1876 (N_1876,N_1363,N_1236);
and U1877 (N_1877,N_1165,N_1464);
nand U1878 (N_1878,N_1097,N_1304);
or U1879 (N_1879,N_1215,N_1035);
and U1880 (N_1880,N_1375,N_1263);
or U1881 (N_1881,N_1271,N_1252);
and U1882 (N_1882,N_1488,N_1208);
nor U1883 (N_1883,N_1013,N_1162);
nand U1884 (N_1884,N_1090,N_1499);
and U1885 (N_1885,N_1332,N_1030);
nand U1886 (N_1886,N_1319,N_1089);
nor U1887 (N_1887,N_1461,N_1230);
nor U1888 (N_1888,N_1022,N_1392);
and U1889 (N_1889,N_1170,N_1186);
nand U1890 (N_1890,N_1496,N_1437);
and U1891 (N_1891,N_1244,N_1055);
and U1892 (N_1892,N_1225,N_1068);
nor U1893 (N_1893,N_1264,N_1312);
nand U1894 (N_1894,N_1465,N_1171);
nand U1895 (N_1895,N_1496,N_1066);
nor U1896 (N_1896,N_1459,N_1432);
and U1897 (N_1897,N_1060,N_1177);
or U1898 (N_1898,N_1383,N_1131);
and U1899 (N_1899,N_1345,N_1102);
nor U1900 (N_1900,N_1030,N_1329);
and U1901 (N_1901,N_1024,N_1484);
nor U1902 (N_1902,N_1078,N_1056);
nand U1903 (N_1903,N_1252,N_1110);
or U1904 (N_1904,N_1143,N_1320);
or U1905 (N_1905,N_1478,N_1002);
or U1906 (N_1906,N_1184,N_1107);
nand U1907 (N_1907,N_1137,N_1305);
nor U1908 (N_1908,N_1261,N_1149);
and U1909 (N_1909,N_1441,N_1302);
and U1910 (N_1910,N_1159,N_1082);
or U1911 (N_1911,N_1491,N_1313);
nand U1912 (N_1912,N_1149,N_1451);
nand U1913 (N_1913,N_1178,N_1307);
or U1914 (N_1914,N_1271,N_1488);
nand U1915 (N_1915,N_1094,N_1134);
nand U1916 (N_1916,N_1024,N_1004);
nor U1917 (N_1917,N_1172,N_1008);
nor U1918 (N_1918,N_1477,N_1073);
or U1919 (N_1919,N_1358,N_1046);
and U1920 (N_1920,N_1013,N_1202);
nand U1921 (N_1921,N_1300,N_1258);
nor U1922 (N_1922,N_1125,N_1204);
nor U1923 (N_1923,N_1247,N_1069);
nand U1924 (N_1924,N_1182,N_1144);
and U1925 (N_1925,N_1159,N_1439);
nor U1926 (N_1926,N_1071,N_1259);
nor U1927 (N_1927,N_1384,N_1181);
nand U1928 (N_1928,N_1107,N_1210);
nor U1929 (N_1929,N_1235,N_1283);
and U1930 (N_1930,N_1415,N_1245);
nor U1931 (N_1931,N_1248,N_1183);
nor U1932 (N_1932,N_1047,N_1421);
and U1933 (N_1933,N_1250,N_1194);
or U1934 (N_1934,N_1172,N_1020);
nand U1935 (N_1935,N_1381,N_1105);
nor U1936 (N_1936,N_1248,N_1043);
nor U1937 (N_1937,N_1200,N_1348);
nand U1938 (N_1938,N_1007,N_1241);
nor U1939 (N_1939,N_1448,N_1492);
nand U1940 (N_1940,N_1431,N_1126);
nor U1941 (N_1941,N_1245,N_1324);
nand U1942 (N_1942,N_1067,N_1279);
xor U1943 (N_1943,N_1339,N_1479);
and U1944 (N_1944,N_1260,N_1133);
and U1945 (N_1945,N_1142,N_1057);
nand U1946 (N_1946,N_1136,N_1375);
nand U1947 (N_1947,N_1291,N_1412);
or U1948 (N_1948,N_1221,N_1171);
and U1949 (N_1949,N_1487,N_1090);
nor U1950 (N_1950,N_1459,N_1131);
nor U1951 (N_1951,N_1019,N_1091);
nor U1952 (N_1952,N_1237,N_1306);
or U1953 (N_1953,N_1199,N_1212);
nor U1954 (N_1954,N_1142,N_1424);
nor U1955 (N_1955,N_1267,N_1373);
nand U1956 (N_1956,N_1371,N_1075);
nor U1957 (N_1957,N_1291,N_1316);
nand U1958 (N_1958,N_1481,N_1319);
nand U1959 (N_1959,N_1467,N_1028);
nand U1960 (N_1960,N_1253,N_1372);
nor U1961 (N_1961,N_1164,N_1395);
and U1962 (N_1962,N_1040,N_1144);
or U1963 (N_1963,N_1055,N_1219);
nor U1964 (N_1964,N_1359,N_1477);
or U1965 (N_1965,N_1274,N_1402);
or U1966 (N_1966,N_1357,N_1054);
or U1967 (N_1967,N_1227,N_1343);
nor U1968 (N_1968,N_1453,N_1458);
xnor U1969 (N_1969,N_1126,N_1466);
or U1970 (N_1970,N_1083,N_1273);
nand U1971 (N_1971,N_1017,N_1401);
nor U1972 (N_1972,N_1010,N_1186);
and U1973 (N_1973,N_1241,N_1318);
nand U1974 (N_1974,N_1224,N_1469);
nand U1975 (N_1975,N_1320,N_1024);
nand U1976 (N_1976,N_1486,N_1485);
nor U1977 (N_1977,N_1074,N_1245);
nor U1978 (N_1978,N_1182,N_1023);
nand U1979 (N_1979,N_1392,N_1437);
nand U1980 (N_1980,N_1050,N_1069);
and U1981 (N_1981,N_1078,N_1476);
nand U1982 (N_1982,N_1395,N_1128);
and U1983 (N_1983,N_1466,N_1365);
or U1984 (N_1984,N_1469,N_1417);
nand U1985 (N_1985,N_1464,N_1315);
nand U1986 (N_1986,N_1377,N_1318);
nor U1987 (N_1987,N_1317,N_1044);
and U1988 (N_1988,N_1489,N_1180);
nor U1989 (N_1989,N_1415,N_1257);
nor U1990 (N_1990,N_1280,N_1483);
nand U1991 (N_1991,N_1261,N_1390);
and U1992 (N_1992,N_1046,N_1406);
nor U1993 (N_1993,N_1469,N_1246);
or U1994 (N_1994,N_1225,N_1248);
nand U1995 (N_1995,N_1093,N_1433);
nor U1996 (N_1996,N_1152,N_1439);
nand U1997 (N_1997,N_1338,N_1217);
nor U1998 (N_1998,N_1155,N_1039);
and U1999 (N_1999,N_1017,N_1127);
and U2000 (N_2000,N_1645,N_1913);
or U2001 (N_2001,N_1651,N_1742);
and U2002 (N_2002,N_1515,N_1667);
nor U2003 (N_2003,N_1860,N_1665);
nand U2004 (N_2004,N_1600,N_1863);
and U2005 (N_2005,N_1516,N_1743);
nor U2006 (N_2006,N_1748,N_1893);
or U2007 (N_2007,N_1880,N_1935);
nand U2008 (N_2008,N_1703,N_1779);
or U2009 (N_2009,N_1841,N_1585);
and U2010 (N_2010,N_1956,N_1560);
or U2011 (N_2011,N_1686,N_1986);
or U2012 (N_2012,N_1720,N_1506);
nor U2013 (N_2013,N_1750,N_1662);
nand U2014 (N_2014,N_1640,N_1993);
and U2015 (N_2015,N_1701,N_1940);
and U2016 (N_2016,N_1998,N_1961);
nand U2017 (N_2017,N_1788,N_1738);
nand U2018 (N_2018,N_1710,N_1796);
or U2019 (N_2019,N_1866,N_1716);
nor U2020 (N_2020,N_1916,N_1555);
and U2021 (N_2021,N_1890,N_1769);
or U2022 (N_2022,N_1569,N_1904);
and U2023 (N_2023,N_1994,N_1632);
and U2024 (N_2024,N_1839,N_1643);
nor U2025 (N_2025,N_1894,N_1753);
nor U2026 (N_2026,N_1931,N_1543);
nor U2027 (N_2027,N_1759,N_1656);
or U2028 (N_2028,N_1781,N_1694);
and U2029 (N_2029,N_1576,N_1617);
nor U2030 (N_2030,N_1652,N_1887);
nor U2031 (N_2031,N_1991,N_1877);
nand U2032 (N_2032,N_1823,N_1731);
or U2033 (N_2033,N_1535,N_1911);
nand U2034 (N_2034,N_1666,N_1875);
and U2035 (N_2035,N_1618,N_1886);
xnor U2036 (N_2036,N_1815,N_1970);
or U2037 (N_2037,N_1708,N_1533);
nor U2038 (N_2038,N_1974,N_1871);
nor U2039 (N_2039,N_1592,N_1587);
and U2040 (N_2040,N_1719,N_1715);
nand U2041 (N_2041,N_1704,N_1628);
nor U2042 (N_2042,N_1534,N_1761);
and U2043 (N_2043,N_1567,N_1709);
nor U2044 (N_2044,N_1786,N_1514);
nand U2045 (N_2045,N_1510,N_1959);
or U2046 (N_2046,N_1607,N_1845);
nor U2047 (N_2047,N_1827,N_1856);
nand U2048 (N_2048,N_1676,N_1598);
nand U2049 (N_2049,N_1990,N_1816);
nor U2050 (N_2050,N_1835,N_1732);
and U2051 (N_2051,N_1783,N_1895);
or U2052 (N_2052,N_1699,N_1647);
or U2053 (N_2053,N_1879,N_1995);
or U2054 (N_2054,N_1541,N_1517);
or U2055 (N_2055,N_1899,N_1603);
nor U2056 (N_2056,N_1767,N_1957);
nand U2057 (N_2057,N_1644,N_1696);
nor U2058 (N_2058,N_1649,N_1824);
or U2059 (N_2059,N_1523,N_1967);
nor U2060 (N_2060,N_1776,N_1648);
nor U2061 (N_2061,N_1881,N_1745);
nor U2062 (N_2062,N_1669,N_1758);
and U2063 (N_2063,N_1684,N_1718);
nand U2064 (N_2064,N_1829,N_1646);
or U2065 (N_2065,N_1905,N_1733);
nor U2066 (N_2066,N_1789,N_1528);
nor U2067 (N_2067,N_1689,N_1948);
nand U2068 (N_2068,N_1629,N_1818);
nor U2069 (N_2069,N_1817,N_1942);
nor U2070 (N_2070,N_1688,N_1853);
nor U2071 (N_2071,N_1724,N_1826);
nor U2072 (N_2072,N_1971,N_1531);
and U2073 (N_2073,N_1945,N_1691);
or U2074 (N_2074,N_1932,N_1925);
or U2075 (N_2075,N_1770,N_1568);
or U2076 (N_2076,N_1988,N_1982);
or U2077 (N_2077,N_1946,N_1864);
or U2078 (N_2078,N_1583,N_1519);
and U2079 (N_2079,N_1849,N_1918);
nor U2080 (N_2080,N_1638,N_1921);
nand U2081 (N_2081,N_1819,N_1615);
or U2082 (N_2082,N_1804,N_1828);
or U2083 (N_2083,N_1854,N_1884);
or U2084 (N_2084,N_1682,N_1698);
and U2085 (N_2085,N_1685,N_1923);
and U2086 (N_2086,N_1654,N_1504);
nand U2087 (N_2087,N_1591,N_1520);
nor U2088 (N_2088,N_1883,N_1604);
nor U2089 (N_2089,N_1821,N_1680);
or U2090 (N_2090,N_1540,N_1909);
and U2091 (N_2091,N_1888,N_1848);
nor U2092 (N_2092,N_1589,N_1869);
or U2093 (N_2093,N_1919,N_1976);
and U2094 (N_2094,N_1536,N_1772);
nand U2095 (N_2095,N_1842,N_1642);
nor U2096 (N_2096,N_1798,N_1822);
nand U2097 (N_2097,N_1787,N_1952);
nor U2098 (N_2098,N_1814,N_1502);
or U2099 (N_2099,N_1930,N_1511);
nand U2100 (N_2100,N_1725,N_1601);
or U2101 (N_2101,N_1668,N_1717);
or U2102 (N_2102,N_1693,N_1914);
and U2103 (N_2103,N_1800,N_1855);
nor U2104 (N_2104,N_1846,N_1868);
nand U2105 (N_2105,N_1559,N_1627);
nand U2106 (N_2106,N_1663,N_1527);
and U2107 (N_2107,N_1726,N_1985);
or U2108 (N_2108,N_1766,N_1978);
or U2109 (N_2109,N_1941,N_1746);
and U2110 (N_2110,N_1579,N_1737);
and U2111 (N_2111,N_1874,N_1915);
and U2112 (N_2112,N_1577,N_1962);
and U2113 (N_2113,N_1679,N_1833);
or U2114 (N_2114,N_1987,N_1512);
and U2115 (N_2115,N_1505,N_1508);
nand U2116 (N_2116,N_1614,N_1675);
and U2117 (N_2117,N_1657,N_1844);
nand U2118 (N_2118,N_1713,N_1972);
or U2119 (N_2119,N_1963,N_1530);
nand U2120 (N_2120,N_1714,N_1609);
and U2121 (N_2121,N_1729,N_1736);
and U2122 (N_2122,N_1562,N_1912);
and U2123 (N_2123,N_1859,N_1795);
and U2124 (N_2124,N_1934,N_1660);
nor U2125 (N_2125,N_1581,N_1850);
and U2126 (N_2126,N_1605,N_1805);
nor U2127 (N_2127,N_1791,N_1723);
nor U2128 (N_2128,N_1621,N_1712);
and U2129 (N_2129,N_1898,N_1586);
or U2130 (N_2130,N_1619,N_1794);
and U2131 (N_2131,N_1760,N_1861);
or U2132 (N_2132,N_1922,N_1782);
nand U2133 (N_2133,N_1658,N_1545);
nand U2134 (N_2134,N_1539,N_1937);
nand U2135 (N_2135,N_1885,N_1705);
nor U2136 (N_2136,N_1938,N_1650);
and U2137 (N_2137,N_1683,N_1901);
and U2138 (N_2138,N_1672,N_1843);
or U2139 (N_2139,N_1551,N_1752);
xor U2140 (N_2140,N_1616,N_1953);
nand U2141 (N_2141,N_1623,N_1852);
and U2142 (N_2142,N_1557,N_1588);
nor U2143 (N_2143,N_1754,N_1613);
or U2144 (N_2144,N_1521,N_1566);
nand U2145 (N_2145,N_1548,N_1639);
xnor U2146 (N_2146,N_1744,N_1801);
or U2147 (N_2147,N_1837,N_1740);
or U2148 (N_2148,N_1996,N_1981);
and U2149 (N_2149,N_1602,N_1739);
nor U2150 (N_2150,N_1634,N_1550);
nor U2151 (N_2151,N_1624,N_1812);
and U2152 (N_2152,N_1858,N_1687);
and U2153 (N_2153,N_1674,N_1778);
and U2154 (N_2154,N_1813,N_1870);
nor U2155 (N_2155,N_1896,N_1573);
and U2156 (N_2156,N_1630,N_1608);
and U2157 (N_2157,N_1965,N_1906);
and U2158 (N_2158,N_1622,N_1582);
and U2159 (N_2159,N_1764,N_1825);
and U2160 (N_2160,N_1873,N_1867);
and U2161 (N_2161,N_1721,N_1999);
or U2162 (N_2162,N_1626,N_1917);
and U2163 (N_2163,N_1792,N_1572);
or U2164 (N_2164,N_1964,N_1785);
nor U2165 (N_2165,N_1574,N_1524);
or U2166 (N_2166,N_1851,N_1809);
nor U2167 (N_2167,N_1728,N_1553);
or U2168 (N_2168,N_1525,N_1635);
nor U2169 (N_2169,N_1969,N_1507);
nor U2170 (N_2170,N_1671,N_1831);
or U2171 (N_2171,N_1975,N_1926);
xor U2172 (N_2172,N_1730,N_1878);
nor U2173 (N_2173,N_1735,N_1933);
and U2174 (N_2174,N_1857,N_1538);
or U2175 (N_2175,N_1907,N_1774);
xnor U2176 (N_2176,N_1811,N_1872);
and U2177 (N_2177,N_1775,N_1697);
and U2178 (N_2178,N_1980,N_1768);
nand U2179 (N_2179,N_1659,N_1947);
and U2180 (N_2180,N_1762,N_1711);
and U2181 (N_2181,N_1780,N_1908);
and U2182 (N_2182,N_1678,N_1611);
and U2183 (N_2183,N_1832,N_1700);
nor U2184 (N_2184,N_1722,N_1847);
nand U2185 (N_2185,N_1977,N_1803);
nand U2186 (N_2186,N_1876,N_1771);
or U2187 (N_2187,N_1690,N_1897);
nor U2188 (N_2188,N_1902,N_1564);
nand U2189 (N_2189,N_1653,N_1554);
nand U2190 (N_2190,N_1500,N_1992);
and U2191 (N_2191,N_1862,N_1997);
and U2192 (N_2192,N_1664,N_1612);
and U2193 (N_2193,N_1563,N_1636);
nor U2194 (N_2194,N_1599,N_1637);
nand U2195 (N_2195,N_1891,N_1900);
nor U2196 (N_2196,N_1633,N_1943);
nor U2197 (N_2197,N_1747,N_1802);
nor U2198 (N_2198,N_1677,N_1692);
or U2199 (N_2199,N_1840,N_1751);
and U2200 (N_2200,N_1797,N_1532);
nor U2201 (N_2201,N_1570,N_1892);
nor U2202 (N_2202,N_1928,N_1620);
nor U2203 (N_2203,N_1954,N_1673);
or U2204 (N_2204,N_1596,N_1889);
nand U2205 (N_2205,N_1777,N_1966);
or U2206 (N_2206,N_1641,N_1522);
or U2207 (N_2207,N_1989,N_1707);
nand U2208 (N_2208,N_1513,N_1910);
nand U2209 (N_2209,N_1575,N_1610);
or U2210 (N_2210,N_1939,N_1830);
nor U2211 (N_2211,N_1790,N_1749);
nor U2212 (N_2212,N_1625,N_1756);
or U2213 (N_2213,N_1979,N_1734);
nor U2214 (N_2214,N_1549,N_1501);
nor U2215 (N_2215,N_1951,N_1593);
nand U2216 (N_2216,N_1983,N_1838);
or U2217 (N_2217,N_1544,N_1565);
or U2218 (N_2218,N_1509,N_1537);
nand U2219 (N_2219,N_1773,N_1924);
and U2220 (N_2220,N_1556,N_1706);
or U2221 (N_2221,N_1882,N_1558);
nand U2222 (N_2222,N_1806,N_1807);
and U2223 (N_2223,N_1973,N_1580);
or U2224 (N_2224,N_1763,N_1552);
nor U2225 (N_2225,N_1808,N_1865);
and U2226 (N_2226,N_1526,N_1944);
and U2227 (N_2227,N_1757,N_1584);
nand U2228 (N_2228,N_1793,N_1547);
or U2229 (N_2229,N_1571,N_1542);
nor U2230 (N_2230,N_1727,N_1836);
nor U2231 (N_2231,N_1799,N_1518);
or U2232 (N_2232,N_1631,N_1960);
or U2233 (N_2233,N_1597,N_1949);
nand U2234 (N_2234,N_1834,N_1929);
and U2235 (N_2235,N_1741,N_1784);
or U2236 (N_2236,N_1590,N_1670);
nand U2237 (N_2237,N_1820,N_1958);
nand U2238 (N_2238,N_1578,N_1936);
nor U2239 (N_2239,N_1955,N_1546);
or U2240 (N_2240,N_1503,N_1529);
nand U2241 (N_2241,N_1661,N_1681);
or U2242 (N_2242,N_1903,N_1655);
nand U2243 (N_2243,N_1765,N_1920);
and U2244 (N_2244,N_1561,N_1968);
or U2245 (N_2245,N_1984,N_1755);
or U2246 (N_2246,N_1595,N_1695);
or U2247 (N_2247,N_1594,N_1950);
nand U2248 (N_2248,N_1810,N_1702);
or U2249 (N_2249,N_1927,N_1606);
nor U2250 (N_2250,N_1507,N_1874);
nand U2251 (N_2251,N_1822,N_1563);
or U2252 (N_2252,N_1648,N_1674);
nor U2253 (N_2253,N_1557,N_1555);
and U2254 (N_2254,N_1554,N_1855);
or U2255 (N_2255,N_1718,N_1883);
nor U2256 (N_2256,N_1848,N_1804);
nor U2257 (N_2257,N_1711,N_1738);
nor U2258 (N_2258,N_1656,N_1967);
and U2259 (N_2259,N_1656,N_1973);
nor U2260 (N_2260,N_1660,N_1915);
and U2261 (N_2261,N_1923,N_1546);
and U2262 (N_2262,N_1696,N_1584);
nor U2263 (N_2263,N_1702,N_1940);
nand U2264 (N_2264,N_1781,N_1644);
and U2265 (N_2265,N_1649,N_1534);
nand U2266 (N_2266,N_1781,N_1700);
or U2267 (N_2267,N_1606,N_1729);
nand U2268 (N_2268,N_1784,N_1992);
and U2269 (N_2269,N_1975,N_1553);
and U2270 (N_2270,N_1600,N_1531);
and U2271 (N_2271,N_1890,N_1771);
and U2272 (N_2272,N_1941,N_1966);
and U2273 (N_2273,N_1943,N_1881);
or U2274 (N_2274,N_1852,N_1949);
and U2275 (N_2275,N_1769,N_1768);
nand U2276 (N_2276,N_1766,N_1964);
nor U2277 (N_2277,N_1799,N_1656);
nor U2278 (N_2278,N_1547,N_1684);
or U2279 (N_2279,N_1689,N_1558);
nand U2280 (N_2280,N_1570,N_1994);
and U2281 (N_2281,N_1931,N_1822);
or U2282 (N_2282,N_1778,N_1567);
xnor U2283 (N_2283,N_1889,N_1932);
or U2284 (N_2284,N_1786,N_1831);
or U2285 (N_2285,N_1813,N_1679);
xor U2286 (N_2286,N_1764,N_1736);
nand U2287 (N_2287,N_1521,N_1535);
nor U2288 (N_2288,N_1615,N_1837);
nor U2289 (N_2289,N_1614,N_1788);
and U2290 (N_2290,N_1824,N_1908);
nand U2291 (N_2291,N_1620,N_1829);
nand U2292 (N_2292,N_1682,N_1512);
or U2293 (N_2293,N_1769,N_1915);
nand U2294 (N_2294,N_1651,N_1795);
and U2295 (N_2295,N_1520,N_1756);
and U2296 (N_2296,N_1984,N_1691);
nand U2297 (N_2297,N_1993,N_1611);
and U2298 (N_2298,N_1523,N_1507);
and U2299 (N_2299,N_1623,N_1578);
nand U2300 (N_2300,N_1868,N_1874);
nor U2301 (N_2301,N_1902,N_1527);
and U2302 (N_2302,N_1784,N_1593);
nand U2303 (N_2303,N_1674,N_1914);
nand U2304 (N_2304,N_1990,N_1958);
and U2305 (N_2305,N_1625,N_1821);
nor U2306 (N_2306,N_1975,N_1987);
or U2307 (N_2307,N_1942,N_1513);
or U2308 (N_2308,N_1942,N_1805);
nor U2309 (N_2309,N_1884,N_1579);
nor U2310 (N_2310,N_1731,N_1957);
or U2311 (N_2311,N_1696,N_1769);
nor U2312 (N_2312,N_1961,N_1667);
and U2313 (N_2313,N_1964,N_1869);
nand U2314 (N_2314,N_1801,N_1946);
nand U2315 (N_2315,N_1748,N_1823);
nand U2316 (N_2316,N_1641,N_1501);
or U2317 (N_2317,N_1973,N_1691);
and U2318 (N_2318,N_1556,N_1538);
nor U2319 (N_2319,N_1708,N_1753);
and U2320 (N_2320,N_1566,N_1978);
and U2321 (N_2321,N_1924,N_1605);
nand U2322 (N_2322,N_1793,N_1686);
xnor U2323 (N_2323,N_1516,N_1643);
nand U2324 (N_2324,N_1751,N_1824);
nor U2325 (N_2325,N_1945,N_1690);
or U2326 (N_2326,N_1525,N_1958);
and U2327 (N_2327,N_1851,N_1500);
nand U2328 (N_2328,N_1936,N_1645);
and U2329 (N_2329,N_1936,N_1626);
nand U2330 (N_2330,N_1795,N_1666);
or U2331 (N_2331,N_1870,N_1954);
or U2332 (N_2332,N_1948,N_1842);
nor U2333 (N_2333,N_1712,N_1860);
and U2334 (N_2334,N_1750,N_1903);
nor U2335 (N_2335,N_1786,N_1861);
nand U2336 (N_2336,N_1685,N_1510);
nand U2337 (N_2337,N_1559,N_1651);
and U2338 (N_2338,N_1937,N_1685);
or U2339 (N_2339,N_1512,N_1654);
and U2340 (N_2340,N_1589,N_1738);
or U2341 (N_2341,N_1999,N_1993);
nand U2342 (N_2342,N_1754,N_1773);
nand U2343 (N_2343,N_1541,N_1969);
or U2344 (N_2344,N_1689,N_1903);
nand U2345 (N_2345,N_1591,N_1547);
nand U2346 (N_2346,N_1514,N_1854);
or U2347 (N_2347,N_1760,N_1647);
nand U2348 (N_2348,N_1763,N_1904);
or U2349 (N_2349,N_1611,N_1813);
nand U2350 (N_2350,N_1968,N_1812);
xnor U2351 (N_2351,N_1917,N_1885);
or U2352 (N_2352,N_1855,N_1919);
and U2353 (N_2353,N_1632,N_1951);
or U2354 (N_2354,N_1682,N_1817);
and U2355 (N_2355,N_1886,N_1610);
nand U2356 (N_2356,N_1633,N_1779);
nand U2357 (N_2357,N_1931,N_1751);
nor U2358 (N_2358,N_1569,N_1945);
or U2359 (N_2359,N_1811,N_1777);
nor U2360 (N_2360,N_1951,N_1510);
and U2361 (N_2361,N_1946,N_1877);
nor U2362 (N_2362,N_1856,N_1551);
and U2363 (N_2363,N_1827,N_1876);
or U2364 (N_2364,N_1780,N_1852);
and U2365 (N_2365,N_1937,N_1909);
or U2366 (N_2366,N_1647,N_1704);
nor U2367 (N_2367,N_1814,N_1759);
nand U2368 (N_2368,N_1641,N_1690);
nand U2369 (N_2369,N_1556,N_1539);
or U2370 (N_2370,N_1938,N_1652);
or U2371 (N_2371,N_1785,N_1827);
and U2372 (N_2372,N_1833,N_1985);
or U2373 (N_2373,N_1686,N_1816);
nor U2374 (N_2374,N_1696,N_1898);
or U2375 (N_2375,N_1609,N_1916);
and U2376 (N_2376,N_1793,N_1955);
nand U2377 (N_2377,N_1771,N_1602);
or U2378 (N_2378,N_1544,N_1722);
or U2379 (N_2379,N_1602,N_1634);
nor U2380 (N_2380,N_1935,N_1896);
nand U2381 (N_2381,N_1979,N_1930);
nor U2382 (N_2382,N_1705,N_1731);
nand U2383 (N_2383,N_1987,N_1608);
or U2384 (N_2384,N_1590,N_1560);
and U2385 (N_2385,N_1595,N_1607);
nor U2386 (N_2386,N_1830,N_1975);
nand U2387 (N_2387,N_1692,N_1805);
nor U2388 (N_2388,N_1816,N_1579);
or U2389 (N_2389,N_1531,N_1682);
or U2390 (N_2390,N_1933,N_1575);
or U2391 (N_2391,N_1620,N_1636);
and U2392 (N_2392,N_1893,N_1642);
or U2393 (N_2393,N_1713,N_1664);
nor U2394 (N_2394,N_1784,N_1589);
and U2395 (N_2395,N_1543,N_1708);
or U2396 (N_2396,N_1772,N_1854);
or U2397 (N_2397,N_1796,N_1914);
and U2398 (N_2398,N_1886,N_1731);
nand U2399 (N_2399,N_1585,N_1746);
and U2400 (N_2400,N_1860,N_1882);
nor U2401 (N_2401,N_1828,N_1738);
nor U2402 (N_2402,N_1967,N_1798);
nand U2403 (N_2403,N_1686,N_1593);
nor U2404 (N_2404,N_1596,N_1940);
nand U2405 (N_2405,N_1589,N_1588);
nor U2406 (N_2406,N_1505,N_1552);
nor U2407 (N_2407,N_1963,N_1788);
and U2408 (N_2408,N_1976,N_1991);
and U2409 (N_2409,N_1935,N_1609);
nor U2410 (N_2410,N_1535,N_1759);
or U2411 (N_2411,N_1734,N_1552);
or U2412 (N_2412,N_1634,N_1594);
or U2413 (N_2413,N_1916,N_1867);
nor U2414 (N_2414,N_1579,N_1504);
and U2415 (N_2415,N_1919,N_1646);
and U2416 (N_2416,N_1655,N_1692);
nor U2417 (N_2417,N_1672,N_1754);
and U2418 (N_2418,N_1796,N_1844);
and U2419 (N_2419,N_1529,N_1958);
or U2420 (N_2420,N_1734,N_1661);
and U2421 (N_2421,N_1857,N_1792);
nand U2422 (N_2422,N_1995,N_1679);
or U2423 (N_2423,N_1619,N_1510);
xnor U2424 (N_2424,N_1603,N_1605);
nor U2425 (N_2425,N_1599,N_1566);
nand U2426 (N_2426,N_1750,N_1521);
nor U2427 (N_2427,N_1680,N_1770);
nand U2428 (N_2428,N_1999,N_1759);
nor U2429 (N_2429,N_1889,N_1906);
nor U2430 (N_2430,N_1914,N_1554);
nor U2431 (N_2431,N_1899,N_1949);
and U2432 (N_2432,N_1780,N_1988);
nand U2433 (N_2433,N_1551,N_1543);
and U2434 (N_2434,N_1915,N_1529);
nand U2435 (N_2435,N_1832,N_1504);
and U2436 (N_2436,N_1725,N_1911);
or U2437 (N_2437,N_1759,N_1688);
or U2438 (N_2438,N_1999,N_1905);
and U2439 (N_2439,N_1839,N_1914);
and U2440 (N_2440,N_1927,N_1857);
nand U2441 (N_2441,N_1887,N_1709);
and U2442 (N_2442,N_1914,N_1788);
or U2443 (N_2443,N_1866,N_1933);
and U2444 (N_2444,N_1699,N_1613);
xnor U2445 (N_2445,N_1762,N_1566);
or U2446 (N_2446,N_1980,N_1796);
and U2447 (N_2447,N_1650,N_1533);
and U2448 (N_2448,N_1815,N_1834);
or U2449 (N_2449,N_1733,N_1836);
or U2450 (N_2450,N_1595,N_1939);
nor U2451 (N_2451,N_1718,N_1895);
nor U2452 (N_2452,N_1504,N_1613);
nand U2453 (N_2453,N_1541,N_1503);
nand U2454 (N_2454,N_1592,N_1894);
nor U2455 (N_2455,N_1940,N_1714);
nor U2456 (N_2456,N_1504,N_1577);
and U2457 (N_2457,N_1884,N_1720);
nand U2458 (N_2458,N_1504,N_1866);
or U2459 (N_2459,N_1505,N_1754);
or U2460 (N_2460,N_1550,N_1809);
nor U2461 (N_2461,N_1639,N_1713);
and U2462 (N_2462,N_1911,N_1939);
nor U2463 (N_2463,N_1629,N_1528);
nand U2464 (N_2464,N_1583,N_1846);
nand U2465 (N_2465,N_1584,N_1773);
or U2466 (N_2466,N_1613,N_1806);
xor U2467 (N_2467,N_1993,N_1525);
or U2468 (N_2468,N_1518,N_1545);
and U2469 (N_2469,N_1973,N_1649);
nor U2470 (N_2470,N_1709,N_1857);
nand U2471 (N_2471,N_1618,N_1984);
and U2472 (N_2472,N_1620,N_1907);
and U2473 (N_2473,N_1816,N_1994);
and U2474 (N_2474,N_1817,N_1571);
and U2475 (N_2475,N_1574,N_1657);
nor U2476 (N_2476,N_1958,N_1916);
nor U2477 (N_2477,N_1837,N_1512);
xor U2478 (N_2478,N_1600,N_1858);
nand U2479 (N_2479,N_1503,N_1598);
or U2480 (N_2480,N_1751,N_1838);
nor U2481 (N_2481,N_1834,N_1575);
and U2482 (N_2482,N_1708,N_1645);
and U2483 (N_2483,N_1870,N_1735);
or U2484 (N_2484,N_1974,N_1909);
or U2485 (N_2485,N_1721,N_1977);
and U2486 (N_2486,N_1999,N_1832);
nor U2487 (N_2487,N_1997,N_1791);
or U2488 (N_2488,N_1920,N_1973);
nand U2489 (N_2489,N_1649,N_1720);
or U2490 (N_2490,N_1588,N_1683);
and U2491 (N_2491,N_1741,N_1753);
or U2492 (N_2492,N_1867,N_1748);
or U2493 (N_2493,N_1943,N_1719);
and U2494 (N_2494,N_1586,N_1886);
or U2495 (N_2495,N_1734,N_1692);
and U2496 (N_2496,N_1855,N_1816);
nor U2497 (N_2497,N_1855,N_1633);
or U2498 (N_2498,N_1842,N_1954);
and U2499 (N_2499,N_1830,N_1752);
and U2500 (N_2500,N_2140,N_2425);
or U2501 (N_2501,N_2241,N_2077);
nor U2502 (N_2502,N_2417,N_2052);
and U2503 (N_2503,N_2161,N_2202);
nor U2504 (N_2504,N_2245,N_2451);
and U2505 (N_2505,N_2251,N_2012);
and U2506 (N_2506,N_2483,N_2356);
nor U2507 (N_2507,N_2058,N_2133);
nor U2508 (N_2508,N_2281,N_2086);
and U2509 (N_2509,N_2351,N_2034);
and U2510 (N_2510,N_2230,N_2346);
nor U2511 (N_2511,N_2238,N_2313);
nand U2512 (N_2512,N_2082,N_2211);
nor U2513 (N_2513,N_2299,N_2395);
and U2514 (N_2514,N_2322,N_2329);
nand U2515 (N_2515,N_2009,N_2272);
and U2516 (N_2516,N_2099,N_2427);
and U2517 (N_2517,N_2048,N_2057);
nand U2518 (N_2518,N_2167,N_2355);
nor U2519 (N_2519,N_2364,N_2162);
nor U2520 (N_2520,N_2114,N_2145);
xor U2521 (N_2521,N_2401,N_2404);
nor U2522 (N_2522,N_2337,N_2340);
nor U2523 (N_2523,N_2187,N_2498);
nor U2524 (N_2524,N_2343,N_2460);
nor U2525 (N_2525,N_2113,N_2370);
and U2526 (N_2526,N_2260,N_2361);
nor U2527 (N_2527,N_2111,N_2358);
or U2528 (N_2528,N_2492,N_2029);
or U2529 (N_2529,N_2488,N_2160);
and U2530 (N_2530,N_2352,N_2378);
and U2531 (N_2531,N_2333,N_2231);
and U2532 (N_2532,N_2342,N_2375);
nor U2533 (N_2533,N_2206,N_2153);
or U2534 (N_2534,N_2221,N_2156);
nor U2535 (N_2535,N_2386,N_2440);
nand U2536 (N_2536,N_2495,N_2219);
nor U2537 (N_2537,N_2345,N_2257);
nor U2538 (N_2538,N_2096,N_2213);
nor U2539 (N_2539,N_2317,N_2262);
and U2540 (N_2540,N_2115,N_2007);
nor U2541 (N_2541,N_2042,N_2142);
or U2542 (N_2542,N_2423,N_2470);
nor U2543 (N_2543,N_2429,N_2028);
nor U2544 (N_2544,N_2419,N_2217);
or U2545 (N_2545,N_2189,N_2319);
nand U2546 (N_2546,N_2149,N_2316);
or U2547 (N_2547,N_2023,N_2478);
nor U2548 (N_2548,N_2258,N_2192);
and U2549 (N_2549,N_2475,N_2323);
xor U2550 (N_2550,N_2409,N_2093);
or U2551 (N_2551,N_2239,N_2068);
and U2552 (N_2552,N_2122,N_2128);
and U2553 (N_2553,N_2341,N_2050);
and U2554 (N_2554,N_2216,N_2198);
nand U2555 (N_2555,N_2391,N_2067);
and U2556 (N_2556,N_2416,N_2001);
nand U2557 (N_2557,N_2325,N_2166);
and U2558 (N_2558,N_2083,N_2264);
nor U2559 (N_2559,N_2092,N_2462);
nand U2560 (N_2560,N_2490,N_2004);
or U2561 (N_2561,N_2038,N_2013);
nor U2562 (N_2562,N_2053,N_2434);
and U2563 (N_2563,N_2410,N_2399);
nor U2564 (N_2564,N_2256,N_2125);
or U2565 (N_2565,N_2232,N_2396);
and U2566 (N_2566,N_2458,N_2357);
and U2567 (N_2567,N_2110,N_2151);
nor U2568 (N_2568,N_2267,N_2467);
nand U2569 (N_2569,N_2392,N_2019);
or U2570 (N_2570,N_2307,N_2180);
and U2571 (N_2571,N_2199,N_2225);
nor U2572 (N_2572,N_2081,N_2365);
nand U2573 (N_2573,N_2095,N_2273);
or U2574 (N_2574,N_2044,N_2308);
nand U2575 (N_2575,N_2465,N_2484);
and U2576 (N_2576,N_2105,N_2320);
nand U2577 (N_2577,N_2301,N_2218);
and U2578 (N_2578,N_2448,N_2466);
and U2579 (N_2579,N_2335,N_2190);
and U2580 (N_2580,N_2306,N_2398);
or U2581 (N_2581,N_2049,N_2062);
or U2582 (N_2582,N_2107,N_2336);
or U2583 (N_2583,N_2443,N_2129);
nand U2584 (N_2584,N_2304,N_2477);
and U2585 (N_2585,N_2246,N_2065);
or U2586 (N_2586,N_2175,N_2168);
and U2587 (N_2587,N_2100,N_2310);
nand U2588 (N_2588,N_2247,N_2282);
or U2589 (N_2589,N_2430,N_2303);
and U2590 (N_2590,N_2205,N_2233);
or U2591 (N_2591,N_2384,N_2075);
and U2592 (N_2592,N_2182,N_2033);
and U2593 (N_2593,N_2387,N_2445);
and U2594 (N_2594,N_2152,N_2089);
or U2595 (N_2595,N_2418,N_2084);
nor U2596 (N_2596,N_2131,N_2056);
and U2597 (N_2597,N_2031,N_2453);
nand U2598 (N_2598,N_2435,N_2135);
or U2599 (N_2599,N_2132,N_2286);
nor U2600 (N_2600,N_2324,N_2103);
and U2601 (N_2601,N_2177,N_2176);
and U2602 (N_2602,N_2002,N_2220);
nor U2603 (N_2603,N_2390,N_2097);
nor U2604 (N_2604,N_2312,N_2071);
or U2605 (N_2605,N_2347,N_2380);
or U2606 (N_2606,N_2431,N_2108);
or U2607 (N_2607,N_2382,N_2452);
nand U2608 (N_2608,N_2268,N_2393);
nand U2609 (N_2609,N_2373,N_2250);
nor U2610 (N_2610,N_2274,N_2080);
nand U2611 (N_2611,N_2188,N_2291);
nor U2612 (N_2612,N_2036,N_2191);
nand U2613 (N_2613,N_2457,N_2041);
nor U2614 (N_2614,N_2179,N_2332);
or U2615 (N_2615,N_2172,N_2374);
and U2616 (N_2616,N_2385,N_2094);
and U2617 (N_2617,N_2208,N_2428);
nand U2618 (N_2618,N_2328,N_2234);
nand U2619 (N_2619,N_2116,N_2405);
and U2620 (N_2620,N_2339,N_2447);
and U2621 (N_2621,N_2456,N_2400);
or U2622 (N_2622,N_2330,N_2064);
or U2623 (N_2623,N_2117,N_2059);
nor U2624 (N_2624,N_2441,N_2224);
nand U2625 (N_2625,N_2302,N_2124);
nand U2626 (N_2626,N_2368,N_2076);
nand U2627 (N_2627,N_2214,N_2047);
nor U2628 (N_2628,N_2287,N_2063);
or U2629 (N_2629,N_2388,N_2223);
xnor U2630 (N_2630,N_2020,N_2482);
or U2631 (N_2631,N_2338,N_2464);
and U2632 (N_2632,N_2439,N_2376);
and U2633 (N_2633,N_2253,N_2178);
nor U2634 (N_2634,N_2265,N_2035);
and U2635 (N_2635,N_2136,N_2204);
or U2636 (N_2636,N_2102,N_2315);
and U2637 (N_2637,N_2421,N_2203);
and U2638 (N_2638,N_2266,N_2163);
or U2639 (N_2639,N_2018,N_2277);
nand U2640 (N_2640,N_2344,N_2349);
and U2641 (N_2641,N_2354,N_2109);
or U2642 (N_2642,N_2454,N_2164);
nor U2643 (N_2643,N_2046,N_2173);
nand U2644 (N_2644,N_2106,N_2061);
nor U2645 (N_2645,N_2437,N_2289);
and U2646 (N_2646,N_2074,N_2359);
or U2647 (N_2647,N_2237,N_2037);
or U2648 (N_2648,N_2016,N_2280);
nor U2649 (N_2649,N_2367,N_2181);
or U2650 (N_2650,N_2010,N_2139);
nand U2651 (N_2651,N_2121,N_2331);
nand U2652 (N_2652,N_2024,N_2011);
nor U2653 (N_2653,N_2284,N_2207);
or U2654 (N_2654,N_2126,N_2450);
nand U2655 (N_2655,N_2079,N_2496);
nand U2656 (N_2656,N_2039,N_2120);
and U2657 (N_2657,N_2436,N_2027);
or U2658 (N_2658,N_2150,N_2006);
and U2659 (N_2659,N_2295,N_2311);
nand U2660 (N_2660,N_2292,N_2479);
nand U2661 (N_2661,N_2297,N_2293);
nand U2662 (N_2662,N_2472,N_2446);
nand U2663 (N_2663,N_2269,N_2073);
and U2664 (N_2664,N_2271,N_2169);
and U2665 (N_2665,N_2334,N_2473);
nor U2666 (N_2666,N_2085,N_2438);
or U2667 (N_2667,N_2014,N_2489);
or U2668 (N_2668,N_2305,N_2363);
nand U2669 (N_2669,N_2123,N_2165);
and U2670 (N_2670,N_2261,N_2461);
or U2671 (N_2671,N_2078,N_2055);
nand U2672 (N_2672,N_2459,N_2413);
and U2673 (N_2673,N_2314,N_2248);
nand U2674 (N_2674,N_2285,N_2090);
or U2675 (N_2675,N_2426,N_2383);
or U2676 (N_2676,N_2487,N_2130);
and U2677 (N_2677,N_2411,N_2184);
nand U2678 (N_2678,N_2194,N_2088);
nor U2679 (N_2679,N_2252,N_2101);
or U2680 (N_2680,N_2432,N_2069);
and U2681 (N_2681,N_2379,N_2275);
nor U2682 (N_2682,N_2406,N_2158);
or U2683 (N_2683,N_2300,N_2433);
or U2684 (N_2684,N_2497,N_2104);
nand U2685 (N_2685,N_2159,N_2227);
or U2686 (N_2686,N_2283,N_2212);
nand U2687 (N_2687,N_2259,N_2424);
or U2688 (N_2688,N_2493,N_2228);
nor U2689 (N_2689,N_2141,N_2022);
nor U2690 (N_2690,N_2134,N_2209);
or U2691 (N_2691,N_2449,N_2494);
nor U2692 (N_2692,N_2394,N_2455);
or U2693 (N_2693,N_2112,N_2087);
nor U2694 (N_2694,N_2442,N_2402);
nand U2695 (N_2695,N_2174,N_2254);
nor U2696 (N_2696,N_2279,N_2348);
nor U2697 (N_2697,N_2371,N_2408);
or U2698 (N_2698,N_2154,N_2362);
or U2699 (N_2699,N_2066,N_2235);
nand U2700 (N_2700,N_2025,N_2118);
nor U2701 (N_2701,N_2499,N_2236);
or U2702 (N_2702,N_2389,N_2127);
and U2703 (N_2703,N_2485,N_2326);
nor U2704 (N_2704,N_2444,N_2296);
nor U2705 (N_2705,N_2360,N_2119);
or U2706 (N_2706,N_2407,N_2040);
and U2707 (N_2707,N_2193,N_2215);
xor U2708 (N_2708,N_2185,N_2369);
or U2709 (N_2709,N_2210,N_2353);
nand U2710 (N_2710,N_2294,N_2196);
and U2711 (N_2711,N_2298,N_2143);
nand U2712 (N_2712,N_2422,N_2201);
and U2713 (N_2713,N_2469,N_2397);
and U2714 (N_2714,N_2186,N_2008);
nand U2715 (N_2715,N_2054,N_2278);
nor U2716 (N_2716,N_2015,N_2468);
nor U2717 (N_2717,N_2486,N_2030);
nor U2718 (N_2718,N_2327,N_2412);
and U2719 (N_2719,N_2032,N_2276);
or U2720 (N_2720,N_2491,N_2000);
or U2721 (N_2721,N_2144,N_2060);
nor U2722 (N_2722,N_2420,N_2415);
nor U2723 (N_2723,N_2366,N_2157);
nand U2724 (N_2724,N_2017,N_2463);
and U2725 (N_2725,N_2350,N_2197);
nor U2726 (N_2726,N_2045,N_2098);
nor U2727 (N_2727,N_2243,N_2321);
nand U2728 (N_2728,N_2222,N_2240);
and U2729 (N_2729,N_2255,N_2072);
nor U2730 (N_2730,N_2148,N_2318);
or U2731 (N_2731,N_2471,N_2414);
nand U2732 (N_2732,N_2137,N_2005);
nand U2733 (N_2733,N_2309,N_2043);
and U2734 (N_2734,N_2270,N_2403);
and U2735 (N_2735,N_2026,N_2249);
and U2736 (N_2736,N_2377,N_2480);
nand U2737 (N_2737,N_2372,N_2290);
nor U2738 (N_2738,N_2381,N_2229);
and U2739 (N_2739,N_2070,N_2021);
nor U2740 (N_2740,N_2091,N_2244);
or U2741 (N_2741,N_2226,N_2051);
nand U2742 (N_2742,N_2200,N_2170);
or U2743 (N_2743,N_2195,N_2171);
and U2744 (N_2744,N_2242,N_2474);
or U2745 (N_2745,N_2288,N_2003);
nand U2746 (N_2746,N_2263,N_2138);
nand U2747 (N_2747,N_2147,N_2146);
nand U2748 (N_2748,N_2183,N_2476);
and U2749 (N_2749,N_2481,N_2155);
nand U2750 (N_2750,N_2228,N_2042);
or U2751 (N_2751,N_2271,N_2017);
and U2752 (N_2752,N_2414,N_2236);
nand U2753 (N_2753,N_2144,N_2140);
and U2754 (N_2754,N_2456,N_2027);
nand U2755 (N_2755,N_2084,N_2014);
nand U2756 (N_2756,N_2084,N_2036);
or U2757 (N_2757,N_2296,N_2454);
nand U2758 (N_2758,N_2172,N_2107);
nand U2759 (N_2759,N_2310,N_2378);
nor U2760 (N_2760,N_2027,N_2320);
nand U2761 (N_2761,N_2497,N_2014);
and U2762 (N_2762,N_2361,N_2252);
and U2763 (N_2763,N_2358,N_2336);
or U2764 (N_2764,N_2384,N_2089);
nand U2765 (N_2765,N_2190,N_2171);
or U2766 (N_2766,N_2044,N_2484);
nand U2767 (N_2767,N_2108,N_2445);
and U2768 (N_2768,N_2485,N_2339);
nor U2769 (N_2769,N_2065,N_2276);
nor U2770 (N_2770,N_2164,N_2342);
or U2771 (N_2771,N_2155,N_2079);
and U2772 (N_2772,N_2324,N_2366);
or U2773 (N_2773,N_2388,N_2330);
nor U2774 (N_2774,N_2344,N_2188);
nor U2775 (N_2775,N_2438,N_2400);
nor U2776 (N_2776,N_2185,N_2412);
nor U2777 (N_2777,N_2334,N_2423);
or U2778 (N_2778,N_2493,N_2243);
and U2779 (N_2779,N_2029,N_2302);
nor U2780 (N_2780,N_2157,N_2378);
nand U2781 (N_2781,N_2014,N_2453);
nor U2782 (N_2782,N_2411,N_2226);
or U2783 (N_2783,N_2074,N_2479);
nor U2784 (N_2784,N_2480,N_2005);
nor U2785 (N_2785,N_2469,N_2135);
nand U2786 (N_2786,N_2133,N_2040);
nor U2787 (N_2787,N_2308,N_2264);
or U2788 (N_2788,N_2053,N_2261);
nor U2789 (N_2789,N_2275,N_2172);
nor U2790 (N_2790,N_2390,N_2170);
or U2791 (N_2791,N_2428,N_2117);
nor U2792 (N_2792,N_2298,N_2152);
or U2793 (N_2793,N_2075,N_2091);
nor U2794 (N_2794,N_2319,N_2051);
or U2795 (N_2795,N_2323,N_2443);
and U2796 (N_2796,N_2461,N_2001);
or U2797 (N_2797,N_2054,N_2032);
nand U2798 (N_2798,N_2282,N_2031);
and U2799 (N_2799,N_2231,N_2297);
nand U2800 (N_2800,N_2214,N_2160);
xor U2801 (N_2801,N_2470,N_2026);
nor U2802 (N_2802,N_2103,N_2283);
or U2803 (N_2803,N_2178,N_2330);
and U2804 (N_2804,N_2148,N_2305);
and U2805 (N_2805,N_2183,N_2356);
or U2806 (N_2806,N_2387,N_2239);
nand U2807 (N_2807,N_2072,N_2390);
and U2808 (N_2808,N_2179,N_2303);
or U2809 (N_2809,N_2488,N_2184);
nor U2810 (N_2810,N_2327,N_2310);
and U2811 (N_2811,N_2096,N_2427);
nor U2812 (N_2812,N_2050,N_2037);
and U2813 (N_2813,N_2094,N_2319);
or U2814 (N_2814,N_2314,N_2412);
and U2815 (N_2815,N_2003,N_2350);
and U2816 (N_2816,N_2494,N_2237);
nor U2817 (N_2817,N_2426,N_2467);
nor U2818 (N_2818,N_2339,N_2315);
or U2819 (N_2819,N_2259,N_2461);
nand U2820 (N_2820,N_2425,N_2434);
and U2821 (N_2821,N_2185,N_2260);
nand U2822 (N_2822,N_2164,N_2067);
nor U2823 (N_2823,N_2454,N_2009);
xor U2824 (N_2824,N_2153,N_2013);
nand U2825 (N_2825,N_2326,N_2289);
xor U2826 (N_2826,N_2471,N_2258);
and U2827 (N_2827,N_2333,N_2010);
nor U2828 (N_2828,N_2067,N_2065);
or U2829 (N_2829,N_2361,N_2031);
nand U2830 (N_2830,N_2036,N_2316);
nor U2831 (N_2831,N_2087,N_2201);
or U2832 (N_2832,N_2408,N_2186);
nor U2833 (N_2833,N_2106,N_2199);
nor U2834 (N_2834,N_2377,N_2423);
nand U2835 (N_2835,N_2457,N_2265);
or U2836 (N_2836,N_2373,N_2226);
xor U2837 (N_2837,N_2331,N_2295);
and U2838 (N_2838,N_2059,N_2290);
and U2839 (N_2839,N_2321,N_2213);
or U2840 (N_2840,N_2117,N_2131);
or U2841 (N_2841,N_2471,N_2372);
nor U2842 (N_2842,N_2435,N_2090);
nand U2843 (N_2843,N_2131,N_2155);
and U2844 (N_2844,N_2343,N_2350);
or U2845 (N_2845,N_2243,N_2305);
nor U2846 (N_2846,N_2118,N_2324);
nor U2847 (N_2847,N_2032,N_2291);
nor U2848 (N_2848,N_2104,N_2174);
nor U2849 (N_2849,N_2026,N_2081);
nand U2850 (N_2850,N_2324,N_2015);
or U2851 (N_2851,N_2319,N_2317);
nor U2852 (N_2852,N_2123,N_2351);
nand U2853 (N_2853,N_2117,N_2415);
nor U2854 (N_2854,N_2313,N_2446);
nor U2855 (N_2855,N_2209,N_2107);
or U2856 (N_2856,N_2339,N_2272);
and U2857 (N_2857,N_2104,N_2353);
nor U2858 (N_2858,N_2173,N_2255);
and U2859 (N_2859,N_2100,N_2099);
and U2860 (N_2860,N_2331,N_2116);
or U2861 (N_2861,N_2229,N_2096);
nand U2862 (N_2862,N_2395,N_2052);
and U2863 (N_2863,N_2417,N_2030);
nor U2864 (N_2864,N_2145,N_2085);
nor U2865 (N_2865,N_2079,N_2223);
or U2866 (N_2866,N_2170,N_2147);
nor U2867 (N_2867,N_2268,N_2183);
or U2868 (N_2868,N_2294,N_2342);
and U2869 (N_2869,N_2136,N_2301);
nor U2870 (N_2870,N_2082,N_2429);
and U2871 (N_2871,N_2071,N_2381);
nand U2872 (N_2872,N_2446,N_2398);
and U2873 (N_2873,N_2155,N_2088);
nor U2874 (N_2874,N_2030,N_2078);
nor U2875 (N_2875,N_2409,N_2008);
nor U2876 (N_2876,N_2025,N_2459);
nor U2877 (N_2877,N_2402,N_2178);
nor U2878 (N_2878,N_2134,N_2007);
nor U2879 (N_2879,N_2043,N_2348);
nor U2880 (N_2880,N_2099,N_2098);
and U2881 (N_2881,N_2495,N_2006);
or U2882 (N_2882,N_2447,N_2009);
or U2883 (N_2883,N_2402,N_2279);
or U2884 (N_2884,N_2288,N_2078);
nor U2885 (N_2885,N_2202,N_2010);
and U2886 (N_2886,N_2285,N_2472);
or U2887 (N_2887,N_2256,N_2137);
or U2888 (N_2888,N_2299,N_2377);
nor U2889 (N_2889,N_2194,N_2069);
and U2890 (N_2890,N_2357,N_2179);
nand U2891 (N_2891,N_2005,N_2049);
nor U2892 (N_2892,N_2151,N_2270);
nor U2893 (N_2893,N_2277,N_2286);
or U2894 (N_2894,N_2112,N_2339);
or U2895 (N_2895,N_2013,N_2454);
nand U2896 (N_2896,N_2456,N_2341);
or U2897 (N_2897,N_2354,N_2022);
and U2898 (N_2898,N_2099,N_2256);
and U2899 (N_2899,N_2362,N_2374);
nor U2900 (N_2900,N_2272,N_2373);
nor U2901 (N_2901,N_2133,N_2286);
nor U2902 (N_2902,N_2212,N_2385);
or U2903 (N_2903,N_2339,N_2217);
nand U2904 (N_2904,N_2054,N_2281);
and U2905 (N_2905,N_2191,N_2402);
or U2906 (N_2906,N_2314,N_2379);
and U2907 (N_2907,N_2405,N_2109);
or U2908 (N_2908,N_2468,N_2431);
and U2909 (N_2909,N_2090,N_2057);
or U2910 (N_2910,N_2196,N_2230);
nor U2911 (N_2911,N_2165,N_2461);
or U2912 (N_2912,N_2326,N_2170);
or U2913 (N_2913,N_2350,N_2415);
and U2914 (N_2914,N_2070,N_2230);
and U2915 (N_2915,N_2113,N_2041);
nand U2916 (N_2916,N_2328,N_2175);
and U2917 (N_2917,N_2179,N_2163);
nand U2918 (N_2918,N_2439,N_2430);
or U2919 (N_2919,N_2216,N_2386);
nor U2920 (N_2920,N_2214,N_2055);
nor U2921 (N_2921,N_2461,N_2481);
nor U2922 (N_2922,N_2243,N_2071);
and U2923 (N_2923,N_2440,N_2241);
and U2924 (N_2924,N_2018,N_2351);
and U2925 (N_2925,N_2350,N_2335);
nand U2926 (N_2926,N_2297,N_2105);
and U2927 (N_2927,N_2422,N_2260);
or U2928 (N_2928,N_2435,N_2490);
or U2929 (N_2929,N_2021,N_2489);
or U2930 (N_2930,N_2053,N_2448);
and U2931 (N_2931,N_2450,N_2187);
nand U2932 (N_2932,N_2369,N_2434);
nand U2933 (N_2933,N_2268,N_2360);
nor U2934 (N_2934,N_2084,N_2425);
and U2935 (N_2935,N_2291,N_2488);
and U2936 (N_2936,N_2071,N_2472);
and U2937 (N_2937,N_2057,N_2276);
xnor U2938 (N_2938,N_2010,N_2445);
or U2939 (N_2939,N_2326,N_2108);
and U2940 (N_2940,N_2262,N_2419);
nor U2941 (N_2941,N_2097,N_2116);
nand U2942 (N_2942,N_2062,N_2347);
or U2943 (N_2943,N_2044,N_2445);
and U2944 (N_2944,N_2146,N_2251);
or U2945 (N_2945,N_2146,N_2071);
nor U2946 (N_2946,N_2145,N_2004);
and U2947 (N_2947,N_2017,N_2319);
nor U2948 (N_2948,N_2064,N_2100);
and U2949 (N_2949,N_2287,N_2165);
nor U2950 (N_2950,N_2211,N_2181);
and U2951 (N_2951,N_2472,N_2445);
or U2952 (N_2952,N_2225,N_2283);
and U2953 (N_2953,N_2366,N_2180);
and U2954 (N_2954,N_2302,N_2253);
and U2955 (N_2955,N_2178,N_2064);
nor U2956 (N_2956,N_2268,N_2447);
and U2957 (N_2957,N_2006,N_2268);
nand U2958 (N_2958,N_2010,N_2385);
nor U2959 (N_2959,N_2238,N_2105);
or U2960 (N_2960,N_2021,N_2202);
and U2961 (N_2961,N_2315,N_2091);
xnor U2962 (N_2962,N_2213,N_2146);
nand U2963 (N_2963,N_2201,N_2304);
nor U2964 (N_2964,N_2199,N_2485);
and U2965 (N_2965,N_2180,N_2241);
nor U2966 (N_2966,N_2334,N_2176);
xnor U2967 (N_2967,N_2039,N_2187);
and U2968 (N_2968,N_2009,N_2055);
nor U2969 (N_2969,N_2100,N_2301);
nand U2970 (N_2970,N_2062,N_2458);
or U2971 (N_2971,N_2178,N_2494);
and U2972 (N_2972,N_2048,N_2473);
nor U2973 (N_2973,N_2162,N_2427);
nor U2974 (N_2974,N_2364,N_2397);
nor U2975 (N_2975,N_2163,N_2059);
nor U2976 (N_2976,N_2161,N_2341);
or U2977 (N_2977,N_2339,N_2020);
or U2978 (N_2978,N_2208,N_2106);
or U2979 (N_2979,N_2016,N_2480);
nand U2980 (N_2980,N_2356,N_2042);
or U2981 (N_2981,N_2092,N_2317);
nor U2982 (N_2982,N_2139,N_2253);
or U2983 (N_2983,N_2301,N_2325);
or U2984 (N_2984,N_2401,N_2315);
nor U2985 (N_2985,N_2425,N_2219);
nor U2986 (N_2986,N_2299,N_2454);
nand U2987 (N_2987,N_2018,N_2133);
and U2988 (N_2988,N_2486,N_2090);
or U2989 (N_2989,N_2117,N_2199);
and U2990 (N_2990,N_2254,N_2385);
nand U2991 (N_2991,N_2459,N_2464);
and U2992 (N_2992,N_2388,N_2429);
nor U2993 (N_2993,N_2361,N_2359);
nand U2994 (N_2994,N_2102,N_2241);
or U2995 (N_2995,N_2321,N_2383);
and U2996 (N_2996,N_2169,N_2125);
and U2997 (N_2997,N_2321,N_2051);
nor U2998 (N_2998,N_2159,N_2234);
or U2999 (N_2999,N_2485,N_2463);
nand U3000 (N_3000,N_2658,N_2564);
or U3001 (N_3001,N_2595,N_2747);
nand U3002 (N_3002,N_2851,N_2729);
and U3003 (N_3003,N_2930,N_2645);
xnor U3004 (N_3004,N_2966,N_2889);
and U3005 (N_3005,N_2810,N_2788);
or U3006 (N_3006,N_2840,N_2994);
nor U3007 (N_3007,N_2869,N_2519);
nand U3008 (N_3008,N_2937,N_2524);
or U3009 (N_3009,N_2567,N_2861);
nor U3010 (N_3010,N_2902,N_2804);
and U3011 (N_3011,N_2728,N_2936);
and U3012 (N_3012,N_2617,N_2976);
nor U3013 (N_3013,N_2980,N_2755);
or U3014 (N_3014,N_2708,N_2673);
and U3015 (N_3015,N_2569,N_2856);
nor U3016 (N_3016,N_2963,N_2648);
nand U3017 (N_3017,N_2894,N_2985);
or U3018 (N_3018,N_2609,N_2814);
nor U3019 (N_3019,N_2642,N_2874);
nor U3020 (N_3020,N_2765,N_2596);
nand U3021 (N_3021,N_2749,N_2721);
or U3022 (N_3022,N_2694,N_2759);
or U3023 (N_3023,N_2972,N_2982);
nor U3024 (N_3024,N_2657,N_2723);
and U3025 (N_3025,N_2919,N_2960);
nor U3026 (N_3026,N_2622,N_2614);
or U3027 (N_3027,N_2616,N_2741);
or U3028 (N_3028,N_2999,N_2654);
nand U3029 (N_3029,N_2732,N_2568);
nor U3030 (N_3030,N_2899,N_2775);
nand U3031 (N_3031,N_2895,N_2761);
and U3032 (N_3032,N_2929,N_2957);
nand U3033 (N_3033,N_2961,N_2865);
nor U3034 (N_3034,N_2707,N_2954);
and U3035 (N_3035,N_2717,N_2688);
or U3036 (N_3036,N_2964,N_2668);
nand U3037 (N_3037,N_2752,N_2795);
nor U3038 (N_3038,N_2867,N_2855);
nand U3039 (N_3039,N_2881,N_2698);
and U3040 (N_3040,N_2720,N_2998);
or U3041 (N_3041,N_2634,N_2534);
nor U3042 (N_3042,N_2639,N_2904);
nor U3043 (N_3043,N_2535,N_2968);
or U3044 (N_3044,N_2823,N_2763);
and U3045 (N_3045,N_2510,N_2913);
xnor U3046 (N_3046,N_2934,N_2638);
and U3047 (N_3047,N_2692,N_2809);
or U3048 (N_3048,N_2532,N_2601);
or U3049 (N_3049,N_2852,N_2676);
nand U3050 (N_3050,N_2602,N_2892);
nor U3051 (N_3051,N_2822,N_2635);
nand U3052 (N_3052,N_2562,N_2826);
nand U3053 (N_3053,N_2770,N_2608);
or U3054 (N_3054,N_2613,N_2610);
nor U3055 (N_3055,N_2706,N_2956);
nand U3056 (N_3056,N_2912,N_2592);
nand U3057 (N_3057,N_2883,N_2719);
and U3058 (N_3058,N_2644,N_2695);
nand U3059 (N_3059,N_2838,N_2818);
nand U3060 (N_3060,N_2570,N_2783);
and U3061 (N_3061,N_2647,N_2864);
nand U3062 (N_3062,N_2983,N_2683);
nand U3063 (N_3063,N_2819,N_2841);
and U3064 (N_3064,N_2882,N_2834);
nor U3065 (N_3065,N_2915,N_2751);
and U3066 (N_3066,N_2884,N_2900);
or U3067 (N_3067,N_2794,N_2790);
nand U3068 (N_3068,N_2766,N_2726);
nor U3069 (N_3069,N_2559,N_2646);
or U3070 (N_3070,N_2828,N_2573);
or U3071 (N_3071,N_2932,N_2544);
nand U3072 (N_3072,N_2606,N_2757);
and U3073 (N_3073,N_2538,N_2798);
and U3074 (N_3074,N_2944,N_2947);
and U3075 (N_3075,N_2537,N_2878);
nand U3076 (N_3076,N_2962,N_2722);
nand U3077 (N_3077,N_2560,N_2886);
nor U3078 (N_3078,N_2923,N_2628);
nor U3079 (N_3079,N_2920,N_2687);
nor U3080 (N_3080,N_2862,N_2603);
nor U3081 (N_3081,N_2807,N_2522);
or U3082 (N_3082,N_2517,N_2927);
nand U3083 (N_3083,N_2933,N_2831);
nor U3084 (N_3084,N_2565,N_2710);
nor U3085 (N_3085,N_2580,N_2776);
and U3086 (N_3086,N_2997,N_2597);
and U3087 (N_3087,N_2636,N_2820);
nand U3088 (N_3088,N_2989,N_2619);
or U3089 (N_3089,N_2812,N_2725);
nor U3090 (N_3090,N_2750,N_2712);
or U3091 (N_3091,N_2896,N_2854);
and U3092 (N_3092,N_2718,N_2802);
nand U3093 (N_3093,N_2769,N_2660);
nand U3094 (N_3094,N_2590,N_2772);
nor U3095 (N_3095,N_2743,N_2662);
nand U3096 (N_3096,N_2873,N_2815);
or U3097 (N_3097,N_2625,N_2893);
nor U3098 (N_3098,N_2779,N_2939);
nor U3099 (N_3099,N_2691,N_2835);
nor U3100 (N_3100,N_2500,N_2605);
nor U3101 (N_3101,N_2531,N_2552);
and U3102 (N_3102,N_2724,N_2686);
and U3103 (N_3103,N_2702,N_2700);
nor U3104 (N_3104,N_2846,N_2773);
or U3105 (N_3105,N_2548,N_2951);
or U3106 (N_3106,N_2604,N_2787);
and U3107 (N_3107,N_2526,N_2670);
or U3108 (N_3108,N_2576,N_2914);
and U3109 (N_3109,N_2921,N_2857);
or U3110 (N_3110,N_2512,N_2827);
nor U3111 (N_3111,N_2950,N_2906);
nor U3112 (N_3112,N_2860,N_2736);
nor U3113 (N_3113,N_2905,N_2916);
nor U3114 (N_3114,N_2942,N_2641);
or U3115 (N_3115,N_2618,N_2612);
nor U3116 (N_3116,N_2653,N_2539);
nand U3117 (N_3117,N_2629,N_2542);
nor U3118 (N_3118,N_2599,N_2554);
or U3119 (N_3119,N_2786,N_2829);
nor U3120 (N_3120,N_2816,N_2656);
and U3121 (N_3121,N_2533,N_2756);
nor U3122 (N_3122,N_2571,N_2824);
and U3123 (N_3123,N_2825,N_2516);
nor U3124 (N_3124,N_2931,N_2711);
and U3125 (N_3125,N_2973,N_2515);
or U3126 (N_3126,N_2620,N_2696);
nand U3127 (N_3127,N_2587,N_2777);
and U3128 (N_3128,N_2607,N_2940);
nor U3129 (N_3129,N_2563,N_2955);
or U3130 (N_3130,N_2746,N_2655);
nand U3131 (N_3131,N_2995,N_2979);
nor U3132 (N_3132,N_2556,N_2791);
and U3133 (N_3133,N_2774,N_2745);
nor U3134 (N_3134,N_2730,N_2967);
or U3135 (N_3135,N_2768,N_2672);
nand U3136 (N_3136,N_2561,N_2782);
or U3137 (N_3137,N_2551,N_2850);
and U3138 (N_3138,N_2843,N_2546);
nor U3139 (N_3139,N_2922,N_2758);
nand U3140 (N_3140,N_2527,N_2611);
nor U3141 (N_3141,N_2689,N_2987);
or U3142 (N_3142,N_2523,N_2945);
nor U3143 (N_3143,N_2764,N_2671);
nand U3144 (N_3144,N_2853,N_2891);
nor U3145 (N_3145,N_2742,N_2970);
nor U3146 (N_3146,N_2615,N_2566);
and U3147 (N_3147,N_2778,N_2578);
nand U3148 (N_3148,N_2858,N_2977);
nor U3149 (N_3149,N_2792,N_2924);
nand U3150 (N_3150,N_2935,N_2953);
or U3151 (N_3151,N_2907,N_2594);
nor U3152 (N_3152,N_2502,N_2507);
and U3153 (N_3153,N_2514,N_2627);
or U3154 (N_3154,N_2577,N_2740);
or U3155 (N_3155,N_2553,N_2842);
nand U3156 (N_3156,N_2591,N_2697);
nand U3157 (N_3157,N_2789,N_2793);
nand U3158 (N_3158,N_2879,N_2784);
nand U3159 (N_3159,N_2897,N_2701);
or U3160 (N_3160,N_2880,N_2704);
and U3161 (N_3161,N_2928,N_2811);
nor U3162 (N_3162,N_2941,N_2659);
nand U3163 (N_3163,N_2529,N_2525);
nor U3164 (N_3164,N_2991,N_2543);
nor U3165 (N_3165,N_2589,N_2665);
or U3166 (N_3166,N_2583,N_2925);
nor U3167 (N_3167,N_2875,N_2518);
nor U3168 (N_3168,N_2572,N_2969);
nand U3169 (N_3169,N_2859,N_2753);
or U3170 (N_3170,N_2909,N_2682);
or U3171 (N_3171,N_2677,N_2585);
or U3172 (N_3172,N_2744,N_2830);
nor U3173 (N_3173,N_2974,N_2650);
and U3174 (N_3174,N_2986,N_2958);
and U3175 (N_3175,N_2870,N_2505);
and U3176 (N_3176,N_2513,N_2716);
and U3177 (N_3177,N_2681,N_2643);
and U3178 (N_3178,N_2959,N_2952);
nor U3179 (N_3179,N_2801,N_2817);
and U3180 (N_3180,N_2806,N_2888);
nor U3181 (N_3181,N_2651,N_2549);
and U3182 (N_3182,N_2637,N_2690);
or U3183 (N_3183,N_2738,N_2675);
or U3184 (N_3184,N_2624,N_2547);
nand U3185 (N_3185,N_2581,N_2984);
and U3186 (N_3186,N_2988,N_2876);
xor U3187 (N_3187,N_2785,N_2661);
and U3188 (N_3188,N_2848,N_2832);
nand U3189 (N_3189,N_2993,N_2714);
nand U3190 (N_3190,N_2530,N_2508);
nor U3191 (N_3191,N_2975,N_2623);
and U3192 (N_3192,N_2803,N_2990);
or U3193 (N_3193,N_2621,N_2693);
and U3194 (N_3194,N_2938,N_2703);
and U3195 (N_3195,N_2946,N_2911);
nor U3196 (N_3196,N_2713,N_2917);
and U3197 (N_3197,N_2511,N_2632);
or U3198 (N_3198,N_2981,N_2890);
nor U3199 (N_3199,N_2805,N_2735);
nor U3200 (N_3200,N_2885,N_2705);
and U3201 (N_3201,N_2575,N_2593);
or U3202 (N_3202,N_2948,N_2833);
nor U3203 (N_3203,N_2908,N_2536);
nor U3204 (N_3204,N_2579,N_2540);
xnor U3205 (N_3205,N_2845,N_2521);
or U3206 (N_3206,N_2978,N_2898);
nor U3207 (N_3207,N_2748,N_2754);
nand U3208 (N_3208,N_2506,N_2630);
or U3209 (N_3209,N_2734,N_2877);
and U3210 (N_3210,N_2965,N_2910);
nor U3211 (N_3211,N_2781,N_2797);
and U3212 (N_3212,N_2586,N_2664);
nor U3213 (N_3213,N_2762,N_2588);
or U3214 (N_3214,N_2631,N_2780);
nor U3215 (N_3215,N_2715,N_2584);
nand U3216 (N_3216,N_2739,N_2863);
nor U3217 (N_3217,N_2847,N_2598);
or U3218 (N_3218,N_2680,N_2872);
nor U3219 (N_3219,N_2550,N_2582);
nor U3220 (N_3220,N_2545,N_2868);
or U3221 (N_3221,N_2992,N_2558);
nand U3222 (N_3222,N_2767,N_2737);
nand U3223 (N_3223,N_2685,N_2557);
or U3224 (N_3224,N_2666,N_2800);
xor U3225 (N_3225,N_2799,N_2771);
and U3226 (N_3226,N_2731,N_2836);
nand U3227 (N_3227,N_2813,N_2679);
and U3228 (N_3228,N_2943,N_2663);
and U3229 (N_3229,N_2520,N_2808);
nand U3230 (N_3230,N_2678,N_2669);
nor U3231 (N_3231,N_2839,N_2509);
or U3232 (N_3232,N_2849,N_2709);
or U3233 (N_3233,N_2684,N_2667);
nand U3234 (N_3234,N_2640,N_2887);
and U3235 (N_3235,N_2626,N_2837);
or U3236 (N_3236,N_2844,N_2528);
and U3237 (N_3237,N_2633,N_2649);
or U3238 (N_3238,N_2903,N_2574);
or U3239 (N_3239,N_2901,N_2727);
or U3240 (N_3240,N_2926,N_2504);
and U3241 (N_3241,N_2699,N_2600);
nand U3242 (N_3242,N_2996,N_2674);
or U3243 (N_3243,N_2541,N_2796);
nand U3244 (N_3244,N_2652,N_2971);
nand U3245 (N_3245,N_2760,N_2949);
nand U3246 (N_3246,N_2501,N_2821);
or U3247 (N_3247,N_2866,N_2918);
and U3248 (N_3248,N_2871,N_2733);
nor U3249 (N_3249,N_2555,N_2503);
nand U3250 (N_3250,N_2582,N_2889);
nand U3251 (N_3251,N_2687,N_2995);
or U3252 (N_3252,N_2645,N_2923);
and U3253 (N_3253,N_2516,N_2633);
and U3254 (N_3254,N_2906,N_2754);
and U3255 (N_3255,N_2687,N_2597);
or U3256 (N_3256,N_2836,N_2937);
or U3257 (N_3257,N_2957,N_2519);
nand U3258 (N_3258,N_2927,N_2808);
nand U3259 (N_3259,N_2953,N_2969);
and U3260 (N_3260,N_2895,N_2625);
nand U3261 (N_3261,N_2519,N_2852);
and U3262 (N_3262,N_2548,N_2512);
nor U3263 (N_3263,N_2713,N_2797);
and U3264 (N_3264,N_2984,N_2706);
and U3265 (N_3265,N_2650,N_2903);
nor U3266 (N_3266,N_2980,N_2777);
nor U3267 (N_3267,N_2812,N_2715);
nor U3268 (N_3268,N_2691,N_2769);
and U3269 (N_3269,N_2532,N_2913);
nand U3270 (N_3270,N_2819,N_2790);
or U3271 (N_3271,N_2644,N_2579);
or U3272 (N_3272,N_2760,N_2651);
or U3273 (N_3273,N_2941,N_2856);
and U3274 (N_3274,N_2671,N_2772);
nand U3275 (N_3275,N_2575,N_2842);
or U3276 (N_3276,N_2798,N_2605);
and U3277 (N_3277,N_2769,N_2899);
and U3278 (N_3278,N_2869,N_2864);
or U3279 (N_3279,N_2537,N_2581);
and U3280 (N_3280,N_2854,N_2876);
nand U3281 (N_3281,N_2913,N_2938);
or U3282 (N_3282,N_2562,N_2730);
or U3283 (N_3283,N_2625,N_2632);
and U3284 (N_3284,N_2878,N_2921);
and U3285 (N_3285,N_2967,N_2841);
and U3286 (N_3286,N_2609,N_2711);
nor U3287 (N_3287,N_2952,N_2799);
nor U3288 (N_3288,N_2575,N_2716);
nand U3289 (N_3289,N_2820,N_2764);
nor U3290 (N_3290,N_2989,N_2651);
nand U3291 (N_3291,N_2697,N_2607);
nand U3292 (N_3292,N_2853,N_2684);
and U3293 (N_3293,N_2950,N_2693);
nor U3294 (N_3294,N_2533,N_2877);
or U3295 (N_3295,N_2746,N_2667);
nand U3296 (N_3296,N_2502,N_2755);
nand U3297 (N_3297,N_2987,N_2612);
nor U3298 (N_3298,N_2734,N_2996);
or U3299 (N_3299,N_2580,N_2798);
nand U3300 (N_3300,N_2943,N_2999);
nor U3301 (N_3301,N_2731,N_2855);
nand U3302 (N_3302,N_2777,N_2669);
or U3303 (N_3303,N_2729,N_2728);
nand U3304 (N_3304,N_2951,N_2913);
nand U3305 (N_3305,N_2878,N_2678);
or U3306 (N_3306,N_2947,N_2653);
nor U3307 (N_3307,N_2772,N_2505);
nand U3308 (N_3308,N_2706,N_2902);
nand U3309 (N_3309,N_2753,N_2990);
or U3310 (N_3310,N_2584,N_2986);
and U3311 (N_3311,N_2745,N_2913);
nand U3312 (N_3312,N_2501,N_2934);
and U3313 (N_3313,N_2859,N_2957);
and U3314 (N_3314,N_2700,N_2996);
nand U3315 (N_3315,N_2920,N_2646);
and U3316 (N_3316,N_2649,N_2504);
nor U3317 (N_3317,N_2520,N_2555);
or U3318 (N_3318,N_2900,N_2944);
nor U3319 (N_3319,N_2793,N_2720);
nand U3320 (N_3320,N_2886,N_2811);
nor U3321 (N_3321,N_2563,N_2863);
or U3322 (N_3322,N_2882,N_2955);
and U3323 (N_3323,N_2576,N_2606);
or U3324 (N_3324,N_2517,N_2657);
or U3325 (N_3325,N_2635,N_2548);
or U3326 (N_3326,N_2501,N_2722);
and U3327 (N_3327,N_2886,N_2571);
nand U3328 (N_3328,N_2625,N_2744);
and U3329 (N_3329,N_2786,N_2621);
and U3330 (N_3330,N_2817,N_2761);
xor U3331 (N_3331,N_2533,N_2740);
and U3332 (N_3332,N_2832,N_2780);
and U3333 (N_3333,N_2850,N_2535);
nand U3334 (N_3334,N_2768,N_2973);
or U3335 (N_3335,N_2816,N_2750);
or U3336 (N_3336,N_2737,N_2733);
nor U3337 (N_3337,N_2562,N_2831);
nor U3338 (N_3338,N_2509,N_2743);
nor U3339 (N_3339,N_2971,N_2948);
nor U3340 (N_3340,N_2831,N_2876);
or U3341 (N_3341,N_2844,N_2567);
nand U3342 (N_3342,N_2658,N_2518);
nand U3343 (N_3343,N_2628,N_2782);
and U3344 (N_3344,N_2691,N_2527);
and U3345 (N_3345,N_2901,N_2843);
nand U3346 (N_3346,N_2852,N_2632);
or U3347 (N_3347,N_2947,N_2567);
nand U3348 (N_3348,N_2720,N_2702);
or U3349 (N_3349,N_2917,N_2916);
and U3350 (N_3350,N_2674,N_2747);
nor U3351 (N_3351,N_2841,N_2662);
and U3352 (N_3352,N_2597,N_2899);
and U3353 (N_3353,N_2873,N_2578);
nand U3354 (N_3354,N_2975,N_2631);
or U3355 (N_3355,N_2793,N_2968);
or U3356 (N_3356,N_2829,N_2894);
nor U3357 (N_3357,N_2967,N_2904);
nand U3358 (N_3358,N_2962,N_2568);
or U3359 (N_3359,N_2646,N_2649);
or U3360 (N_3360,N_2826,N_2867);
nand U3361 (N_3361,N_2877,N_2570);
or U3362 (N_3362,N_2884,N_2507);
or U3363 (N_3363,N_2956,N_2568);
nand U3364 (N_3364,N_2677,N_2823);
nor U3365 (N_3365,N_2868,N_2730);
nor U3366 (N_3366,N_2521,N_2632);
nor U3367 (N_3367,N_2892,N_2648);
nor U3368 (N_3368,N_2739,N_2673);
nor U3369 (N_3369,N_2810,N_2831);
or U3370 (N_3370,N_2504,N_2906);
nor U3371 (N_3371,N_2753,N_2770);
or U3372 (N_3372,N_2961,N_2712);
nor U3373 (N_3373,N_2876,N_2970);
nor U3374 (N_3374,N_2871,N_2678);
nand U3375 (N_3375,N_2997,N_2594);
nor U3376 (N_3376,N_2833,N_2899);
nand U3377 (N_3377,N_2892,N_2503);
nor U3378 (N_3378,N_2722,N_2593);
or U3379 (N_3379,N_2770,N_2869);
and U3380 (N_3380,N_2656,N_2861);
and U3381 (N_3381,N_2753,N_2993);
nor U3382 (N_3382,N_2516,N_2959);
nor U3383 (N_3383,N_2782,N_2565);
and U3384 (N_3384,N_2648,N_2866);
nor U3385 (N_3385,N_2973,N_2773);
and U3386 (N_3386,N_2778,N_2958);
nor U3387 (N_3387,N_2926,N_2537);
nand U3388 (N_3388,N_2902,N_2774);
nand U3389 (N_3389,N_2659,N_2729);
and U3390 (N_3390,N_2626,N_2994);
or U3391 (N_3391,N_2657,N_2796);
or U3392 (N_3392,N_2598,N_2885);
nand U3393 (N_3393,N_2820,N_2987);
or U3394 (N_3394,N_2959,N_2798);
nor U3395 (N_3395,N_2692,N_2542);
or U3396 (N_3396,N_2748,N_2830);
nand U3397 (N_3397,N_2836,N_2934);
or U3398 (N_3398,N_2511,N_2629);
xnor U3399 (N_3399,N_2834,N_2898);
and U3400 (N_3400,N_2625,N_2508);
xnor U3401 (N_3401,N_2594,N_2544);
nor U3402 (N_3402,N_2548,N_2826);
or U3403 (N_3403,N_2883,N_2528);
or U3404 (N_3404,N_2867,N_2696);
nor U3405 (N_3405,N_2672,N_2581);
and U3406 (N_3406,N_2767,N_2779);
and U3407 (N_3407,N_2891,N_2571);
nor U3408 (N_3408,N_2530,N_2692);
and U3409 (N_3409,N_2893,N_2626);
nand U3410 (N_3410,N_2653,N_2542);
nor U3411 (N_3411,N_2553,N_2981);
nor U3412 (N_3412,N_2677,N_2907);
or U3413 (N_3413,N_2742,N_2648);
or U3414 (N_3414,N_2593,N_2837);
and U3415 (N_3415,N_2855,N_2906);
nand U3416 (N_3416,N_2926,N_2828);
and U3417 (N_3417,N_2829,N_2722);
or U3418 (N_3418,N_2794,N_2574);
and U3419 (N_3419,N_2779,N_2827);
or U3420 (N_3420,N_2916,N_2605);
and U3421 (N_3421,N_2738,N_2811);
nor U3422 (N_3422,N_2832,N_2776);
nand U3423 (N_3423,N_2682,N_2735);
nor U3424 (N_3424,N_2622,N_2518);
and U3425 (N_3425,N_2553,N_2625);
nand U3426 (N_3426,N_2914,N_2940);
or U3427 (N_3427,N_2711,N_2532);
or U3428 (N_3428,N_2658,N_2524);
and U3429 (N_3429,N_2633,N_2932);
nand U3430 (N_3430,N_2917,N_2875);
or U3431 (N_3431,N_2617,N_2969);
nor U3432 (N_3432,N_2809,N_2922);
and U3433 (N_3433,N_2798,N_2552);
and U3434 (N_3434,N_2842,N_2601);
nor U3435 (N_3435,N_2811,N_2777);
and U3436 (N_3436,N_2587,N_2970);
and U3437 (N_3437,N_2925,N_2658);
nor U3438 (N_3438,N_2543,N_2768);
or U3439 (N_3439,N_2751,N_2750);
nand U3440 (N_3440,N_2958,N_2557);
and U3441 (N_3441,N_2758,N_2567);
and U3442 (N_3442,N_2650,N_2870);
nand U3443 (N_3443,N_2797,N_2571);
nand U3444 (N_3444,N_2559,N_2531);
or U3445 (N_3445,N_2541,N_2600);
nand U3446 (N_3446,N_2806,N_2501);
or U3447 (N_3447,N_2752,N_2849);
nand U3448 (N_3448,N_2675,N_2729);
and U3449 (N_3449,N_2506,N_2985);
or U3450 (N_3450,N_2592,N_2591);
or U3451 (N_3451,N_2920,N_2694);
and U3452 (N_3452,N_2944,N_2747);
nand U3453 (N_3453,N_2743,N_2947);
and U3454 (N_3454,N_2815,N_2614);
nor U3455 (N_3455,N_2788,N_2978);
nor U3456 (N_3456,N_2768,N_2846);
or U3457 (N_3457,N_2745,N_2984);
nand U3458 (N_3458,N_2613,N_2763);
or U3459 (N_3459,N_2966,N_2671);
nor U3460 (N_3460,N_2895,N_2610);
or U3461 (N_3461,N_2609,N_2726);
or U3462 (N_3462,N_2911,N_2969);
and U3463 (N_3463,N_2996,N_2701);
or U3464 (N_3464,N_2653,N_2782);
nand U3465 (N_3465,N_2663,N_2640);
nand U3466 (N_3466,N_2878,N_2933);
or U3467 (N_3467,N_2642,N_2961);
nand U3468 (N_3468,N_2833,N_2669);
nand U3469 (N_3469,N_2548,N_2704);
nor U3470 (N_3470,N_2840,N_2799);
or U3471 (N_3471,N_2804,N_2879);
nand U3472 (N_3472,N_2655,N_2645);
and U3473 (N_3473,N_2606,N_2741);
nand U3474 (N_3474,N_2785,N_2622);
nor U3475 (N_3475,N_2824,N_2597);
xor U3476 (N_3476,N_2786,N_2684);
nand U3477 (N_3477,N_2609,N_2549);
and U3478 (N_3478,N_2740,N_2693);
nor U3479 (N_3479,N_2595,N_2870);
nor U3480 (N_3480,N_2951,N_2914);
nor U3481 (N_3481,N_2525,N_2543);
or U3482 (N_3482,N_2740,N_2945);
nand U3483 (N_3483,N_2639,N_2898);
and U3484 (N_3484,N_2951,N_2660);
and U3485 (N_3485,N_2736,N_2932);
or U3486 (N_3486,N_2953,N_2832);
or U3487 (N_3487,N_2631,N_2932);
nand U3488 (N_3488,N_2997,N_2549);
nor U3489 (N_3489,N_2579,N_2810);
nand U3490 (N_3490,N_2603,N_2672);
nand U3491 (N_3491,N_2907,N_2642);
or U3492 (N_3492,N_2993,N_2750);
nor U3493 (N_3493,N_2928,N_2836);
or U3494 (N_3494,N_2847,N_2875);
nand U3495 (N_3495,N_2718,N_2702);
or U3496 (N_3496,N_2791,N_2546);
nand U3497 (N_3497,N_2828,N_2776);
nand U3498 (N_3498,N_2512,N_2941);
or U3499 (N_3499,N_2888,N_2900);
or U3500 (N_3500,N_3280,N_3398);
nor U3501 (N_3501,N_3170,N_3117);
and U3502 (N_3502,N_3295,N_3340);
or U3503 (N_3503,N_3099,N_3252);
nand U3504 (N_3504,N_3347,N_3000);
nor U3505 (N_3505,N_3088,N_3459);
nor U3506 (N_3506,N_3351,N_3037);
nor U3507 (N_3507,N_3349,N_3255);
nand U3508 (N_3508,N_3372,N_3231);
and U3509 (N_3509,N_3011,N_3472);
nor U3510 (N_3510,N_3393,N_3498);
or U3511 (N_3511,N_3499,N_3067);
and U3512 (N_3512,N_3019,N_3222);
nand U3513 (N_3513,N_3003,N_3208);
nor U3514 (N_3514,N_3091,N_3266);
or U3515 (N_3515,N_3029,N_3188);
nor U3516 (N_3516,N_3048,N_3150);
nor U3517 (N_3517,N_3213,N_3131);
and U3518 (N_3518,N_3490,N_3310);
and U3519 (N_3519,N_3444,N_3203);
nor U3520 (N_3520,N_3425,N_3427);
xnor U3521 (N_3521,N_3385,N_3350);
and U3522 (N_3522,N_3405,N_3027);
nand U3523 (N_3523,N_3047,N_3026);
nor U3524 (N_3524,N_3002,N_3078);
and U3525 (N_3525,N_3141,N_3030);
and U3526 (N_3526,N_3288,N_3487);
and U3527 (N_3527,N_3390,N_3173);
nand U3528 (N_3528,N_3068,N_3101);
nand U3529 (N_3529,N_3040,N_3479);
or U3530 (N_3530,N_3440,N_3371);
nand U3531 (N_3531,N_3367,N_3057);
nor U3532 (N_3532,N_3332,N_3066);
and U3533 (N_3533,N_3275,N_3401);
nand U3534 (N_3534,N_3442,N_3120);
or U3535 (N_3535,N_3061,N_3361);
and U3536 (N_3536,N_3481,N_3122);
and U3537 (N_3537,N_3060,N_3248);
nand U3538 (N_3538,N_3077,N_3053);
or U3539 (N_3539,N_3100,N_3297);
and U3540 (N_3540,N_3449,N_3278);
nor U3541 (N_3541,N_3375,N_3056);
nand U3542 (N_3542,N_3238,N_3291);
and U3543 (N_3543,N_3197,N_3191);
nand U3544 (N_3544,N_3308,N_3407);
or U3545 (N_3545,N_3109,N_3158);
or U3546 (N_3546,N_3012,N_3443);
nand U3547 (N_3547,N_3098,N_3301);
nand U3548 (N_3548,N_3335,N_3123);
or U3549 (N_3549,N_3286,N_3177);
and U3550 (N_3550,N_3155,N_3320);
nand U3551 (N_3551,N_3148,N_3475);
or U3552 (N_3552,N_3273,N_3272);
nor U3553 (N_3553,N_3355,N_3160);
and U3554 (N_3554,N_3014,N_3467);
nand U3555 (N_3555,N_3094,N_3154);
or U3556 (N_3556,N_3435,N_3179);
nor U3557 (N_3557,N_3492,N_3031);
and U3558 (N_3558,N_3161,N_3083);
nand U3559 (N_3559,N_3451,N_3189);
and U3560 (N_3560,N_3457,N_3129);
and U3561 (N_3561,N_3313,N_3009);
or U3562 (N_3562,N_3192,N_3366);
and U3563 (N_3563,N_3035,N_3309);
nor U3564 (N_3564,N_3430,N_3424);
nand U3565 (N_3565,N_3110,N_3130);
nand U3566 (N_3566,N_3193,N_3403);
nor U3567 (N_3567,N_3384,N_3196);
nor U3568 (N_3568,N_3111,N_3233);
nor U3569 (N_3569,N_3169,N_3043);
nor U3570 (N_3570,N_3071,N_3132);
nand U3571 (N_3571,N_3113,N_3338);
and U3572 (N_3572,N_3432,N_3257);
nand U3573 (N_3573,N_3337,N_3015);
nand U3574 (N_3574,N_3413,N_3339);
or U3575 (N_3575,N_3034,N_3059);
and U3576 (N_3576,N_3323,N_3209);
and U3577 (N_3577,N_3325,N_3382);
nand U3578 (N_3578,N_3477,N_3051);
and U3579 (N_3579,N_3454,N_3108);
and U3580 (N_3580,N_3423,N_3023);
nor U3581 (N_3581,N_3360,N_3317);
nor U3582 (N_3582,N_3227,N_3281);
and U3583 (N_3583,N_3241,N_3473);
nor U3584 (N_3584,N_3041,N_3303);
nor U3585 (N_3585,N_3363,N_3033);
or U3586 (N_3586,N_3396,N_3207);
nor U3587 (N_3587,N_3307,N_3431);
or U3588 (N_3588,N_3290,N_3146);
nand U3589 (N_3589,N_3497,N_3005);
or U3590 (N_3590,N_3462,N_3107);
or U3591 (N_3591,N_3190,N_3089);
xnor U3592 (N_3592,N_3260,N_3478);
or U3593 (N_3593,N_3453,N_3416);
and U3594 (N_3594,N_3326,N_3226);
nand U3595 (N_3595,N_3330,N_3391);
nor U3596 (N_3596,N_3495,N_3439);
or U3597 (N_3597,N_3420,N_3183);
or U3598 (N_3598,N_3400,N_3311);
nand U3599 (N_3599,N_3097,N_3235);
and U3600 (N_3600,N_3247,N_3345);
nor U3601 (N_3601,N_3218,N_3489);
nand U3602 (N_3602,N_3465,N_3239);
or U3603 (N_3603,N_3464,N_3446);
nand U3604 (N_3604,N_3044,N_3016);
and U3605 (N_3605,N_3484,N_3073);
and U3606 (N_3606,N_3463,N_3152);
or U3607 (N_3607,N_3085,N_3333);
nor U3608 (N_3608,N_3368,N_3025);
or U3609 (N_3609,N_3104,N_3352);
nor U3610 (N_3610,N_3164,N_3379);
nor U3611 (N_3611,N_3181,N_3017);
or U3612 (N_3612,N_3476,N_3292);
nor U3613 (N_3613,N_3046,N_3175);
nand U3614 (N_3614,N_3269,N_3039);
nor U3615 (N_3615,N_3377,N_3293);
nor U3616 (N_3616,N_3232,N_3024);
xnor U3617 (N_3617,N_3204,N_3185);
and U3618 (N_3618,N_3329,N_3112);
nand U3619 (N_3619,N_3282,N_3210);
or U3620 (N_3620,N_3187,N_3386);
nor U3621 (N_3621,N_3328,N_3450);
and U3622 (N_3622,N_3483,N_3318);
nand U3623 (N_3623,N_3052,N_3080);
and U3624 (N_3624,N_3397,N_3277);
or U3625 (N_3625,N_3171,N_3010);
or U3626 (N_3626,N_3186,N_3054);
nor U3627 (N_3627,N_3402,N_3229);
or U3628 (N_3628,N_3434,N_3032);
nor U3629 (N_3629,N_3470,N_3182);
nand U3630 (N_3630,N_3394,N_3006);
and U3631 (N_3631,N_3143,N_3139);
or U3632 (N_3632,N_3283,N_3373);
or U3633 (N_3633,N_3460,N_3075);
nand U3634 (N_3634,N_3008,N_3331);
nor U3635 (N_3635,N_3334,N_3485);
xnor U3636 (N_3636,N_3096,N_3421);
nor U3637 (N_3637,N_3092,N_3474);
and U3638 (N_3638,N_3162,N_3168);
nor U3639 (N_3639,N_3215,N_3426);
nand U3640 (N_3640,N_3422,N_3221);
or U3641 (N_3641,N_3365,N_3312);
nand U3642 (N_3642,N_3357,N_3412);
or U3643 (N_3643,N_3176,N_3064);
or U3644 (N_3644,N_3126,N_3270);
or U3645 (N_3645,N_3408,N_3279);
or U3646 (N_3646,N_3072,N_3488);
nor U3647 (N_3647,N_3156,N_3294);
nand U3648 (N_3648,N_3202,N_3315);
or U3649 (N_3649,N_3265,N_3167);
and U3650 (N_3650,N_3262,N_3268);
and U3651 (N_3651,N_3105,N_3086);
nor U3652 (N_3652,N_3304,N_3458);
and U3653 (N_3653,N_3261,N_3151);
nor U3654 (N_3654,N_3429,N_3389);
nor U3655 (N_3655,N_3256,N_3242);
nor U3656 (N_3656,N_3418,N_3127);
nand U3657 (N_3657,N_3259,N_3493);
or U3658 (N_3658,N_3081,N_3198);
nor U3659 (N_3659,N_3336,N_3145);
and U3660 (N_3660,N_3230,N_3195);
or U3661 (N_3661,N_3165,N_3285);
nand U3662 (N_3662,N_3178,N_3321);
nor U3663 (N_3663,N_3201,N_3219);
nor U3664 (N_3664,N_3021,N_3249);
nand U3665 (N_3665,N_3199,N_3433);
and U3666 (N_3666,N_3007,N_3211);
or U3667 (N_3667,N_3095,N_3417);
and U3668 (N_3668,N_3243,N_3228);
nor U3669 (N_3669,N_3159,N_3074);
nor U3670 (N_3670,N_3387,N_3314);
nand U3671 (N_3671,N_3172,N_3376);
or U3672 (N_3672,N_3494,N_3264);
or U3673 (N_3673,N_3374,N_3049);
nand U3674 (N_3674,N_3448,N_3084);
nand U3675 (N_3675,N_3322,N_3267);
nor U3676 (N_3676,N_3036,N_3236);
and U3677 (N_3677,N_3496,N_3468);
or U3678 (N_3678,N_3217,N_3456);
nand U3679 (N_3679,N_3038,N_3020);
nor U3680 (N_3680,N_3106,N_3364);
nand U3681 (N_3681,N_3022,N_3409);
or U3682 (N_3682,N_3380,N_3436);
nor U3683 (N_3683,N_3319,N_3234);
and U3684 (N_3684,N_3245,N_3244);
nand U3685 (N_3685,N_3471,N_3486);
nand U3686 (N_3686,N_3346,N_3466);
and U3687 (N_3687,N_3118,N_3018);
nor U3688 (N_3688,N_3289,N_3306);
and U3689 (N_3689,N_3469,N_3406);
and U3690 (N_3690,N_3258,N_3119);
nand U3691 (N_3691,N_3103,N_3028);
and U3692 (N_3692,N_3237,N_3296);
nor U3693 (N_3693,N_3224,N_3410);
or U3694 (N_3694,N_3153,N_3001);
or U3695 (N_3695,N_3042,N_3205);
or U3696 (N_3696,N_3399,N_3136);
nand U3697 (N_3697,N_3194,N_3452);
nand U3698 (N_3698,N_3287,N_3276);
and U3699 (N_3699,N_3147,N_3263);
or U3700 (N_3700,N_3299,N_3137);
nor U3701 (N_3701,N_3013,N_3220);
or U3702 (N_3702,N_3370,N_3174);
and U3703 (N_3703,N_3133,N_3225);
or U3704 (N_3704,N_3157,N_3004);
nor U3705 (N_3705,N_3271,N_3206);
nor U3706 (N_3706,N_3445,N_3180);
and U3707 (N_3707,N_3302,N_3216);
xnor U3708 (N_3708,N_3362,N_3342);
nor U3709 (N_3709,N_3115,N_3087);
or U3710 (N_3710,N_3461,N_3070);
and U3711 (N_3711,N_3327,N_3447);
xnor U3712 (N_3712,N_3144,N_3438);
and U3713 (N_3713,N_3065,N_3114);
nor U3714 (N_3714,N_3316,N_3093);
nor U3715 (N_3715,N_3140,N_3344);
nand U3716 (N_3716,N_3254,N_3356);
nand U3717 (N_3717,N_3354,N_3480);
nor U3718 (N_3718,N_3284,N_3125);
or U3719 (N_3719,N_3079,N_3274);
or U3720 (N_3720,N_3341,N_3102);
or U3721 (N_3721,N_3240,N_3482);
nor U3722 (N_3722,N_3135,N_3411);
nand U3723 (N_3723,N_3124,N_3149);
nand U3724 (N_3724,N_3166,N_3058);
nor U3725 (N_3725,N_3343,N_3414);
and U3726 (N_3726,N_3383,N_3121);
and U3727 (N_3727,N_3298,N_3395);
nand U3728 (N_3728,N_3348,N_3082);
and U3729 (N_3729,N_3305,N_3223);
or U3730 (N_3730,N_3253,N_3128);
or U3731 (N_3731,N_3076,N_3090);
or U3732 (N_3732,N_3063,N_3491);
nor U3733 (N_3733,N_3050,N_3045);
nor U3734 (N_3734,N_3392,N_3062);
nor U3735 (N_3735,N_3359,N_3069);
or U3736 (N_3736,N_3134,N_3415);
xnor U3737 (N_3737,N_3358,N_3419);
and U3738 (N_3738,N_3184,N_3324);
nor U3739 (N_3739,N_3163,N_3404);
nand U3740 (N_3740,N_3200,N_3353);
nand U3741 (N_3741,N_3116,N_3251);
nor U3742 (N_3742,N_3250,N_3428);
xor U3743 (N_3743,N_3369,N_3441);
nand U3744 (N_3744,N_3300,N_3388);
or U3745 (N_3745,N_3381,N_3437);
or U3746 (N_3746,N_3212,N_3142);
or U3747 (N_3747,N_3378,N_3246);
nand U3748 (N_3748,N_3214,N_3138);
nor U3749 (N_3749,N_3455,N_3055);
nand U3750 (N_3750,N_3124,N_3469);
or U3751 (N_3751,N_3485,N_3441);
nor U3752 (N_3752,N_3056,N_3261);
and U3753 (N_3753,N_3290,N_3387);
and U3754 (N_3754,N_3276,N_3337);
nor U3755 (N_3755,N_3410,N_3247);
or U3756 (N_3756,N_3283,N_3282);
and U3757 (N_3757,N_3257,N_3327);
nor U3758 (N_3758,N_3175,N_3044);
or U3759 (N_3759,N_3438,N_3128);
and U3760 (N_3760,N_3119,N_3050);
or U3761 (N_3761,N_3366,N_3231);
nor U3762 (N_3762,N_3192,N_3476);
and U3763 (N_3763,N_3416,N_3016);
or U3764 (N_3764,N_3197,N_3422);
nor U3765 (N_3765,N_3396,N_3157);
nand U3766 (N_3766,N_3211,N_3091);
or U3767 (N_3767,N_3234,N_3390);
nor U3768 (N_3768,N_3373,N_3028);
nand U3769 (N_3769,N_3092,N_3104);
nand U3770 (N_3770,N_3251,N_3289);
nand U3771 (N_3771,N_3215,N_3121);
and U3772 (N_3772,N_3443,N_3194);
nand U3773 (N_3773,N_3318,N_3403);
or U3774 (N_3774,N_3131,N_3035);
and U3775 (N_3775,N_3055,N_3005);
nand U3776 (N_3776,N_3020,N_3195);
and U3777 (N_3777,N_3447,N_3467);
or U3778 (N_3778,N_3390,N_3490);
or U3779 (N_3779,N_3122,N_3331);
or U3780 (N_3780,N_3186,N_3120);
nand U3781 (N_3781,N_3216,N_3102);
nor U3782 (N_3782,N_3395,N_3436);
or U3783 (N_3783,N_3241,N_3021);
or U3784 (N_3784,N_3453,N_3081);
nor U3785 (N_3785,N_3066,N_3328);
or U3786 (N_3786,N_3458,N_3216);
or U3787 (N_3787,N_3336,N_3473);
nand U3788 (N_3788,N_3183,N_3237);
or U3789 (N_3789,N_3065,N_3465);
nor U3790 (N_3790,N_3169,N_3185);
nand U3791 (N_3791,N_3037,N_3244);
and U3792 (N_3792,N_3434,N_3198);
nand U3793 (N_3793,N_3240,N_3311);
or U3794 (N_3794,N_3000,N_3425);
nand U3795 (N_3795,N_3067,N_3172);
nor U3796 (N_3796,N_3025,N_3223);
and U3797 (N_3797,N_3391,N_3474);
nor U3798 (N_3798,N_3240,N_3399);
nor U3799 (N_3799,N_3120,N_3022);
nand U3800 (N_3800,N_3484,N_3091);
nor U3801 (N_3801,N_3141,N_3332);
and U3802 (N_3802,N_3080,N_3271);
nor U3803 (N_3803,N_3263,N_3412);
nor U3804 (N_3804,N_3458,N_3267);
or U3805 (N_3805,N_3225,N_3373);
nand U3806 (N_3806,N_3362,N_3198);
or U3807 (N_3807,N_3291,N_3436);
or U3808 (N_3808,N_3391,N_3065);
or U3809 (N_3809,N_3031,N_3111);
and U3810 (N_3810,N_3449,N_3368);
or U3811 (N_3811,N_3143,N_3011);
nor U3812 (N_3812,N_3381,N_3082);
or U3813 (N_3813,N_3054,N_3105);
nor U3814 (N_3814,N_3209,N_3003);
nor U3815 (N_3815,N_3049,N_3184);
or U3816 (N_3816,N_3158,N_3405);
nor U3817 (N_3817,N_3245,N_3057);
and U3818 (N_3818,N_3375,N_3239);
or U3819 (N_3819,N_3422,N_3418);
nor U3820 (N_3820,N_3220,N_3430);
and U3821 (N_3821,N_3497,N_3499);
nand U3822 (N_3822,N_3367,N_3162);
and U3823 (N_3823,N_3053,N_3003);
nor U3824 (N_3824,N_3481,N_3119);
nor U3825 (N_3825,N_3164,N_3374);
and U3826 (N_3826,N_3071,N_3238);
and U3827 (N_3827,N_3102,N_3199);
nor U3828 (N_3828,N_3199,N_3209);
and U3829 (N_3829,N_3345,N_3476);
or U3830 (N_3830,N_3480,N_3027);
nand U3831 (N_3831,N_3457,N_3446);
nor U3832 (N_3832,N_3120,N_3322);
nor U3833 (N_3833,N_3202,N_3112);
or U3834 (N_3834,N_3220,N_3182);
nand U3835 (N_3835,N_3041,N_3120);
nor U3836 (N_3836,N_3499,N_3043);
and U3837 (N_3837,N_3262,N_3385);
nand U3838 (N_3838,N_3125,N_3163);
and U3839 (N_3839,N_3022,N_3220);
nand U3840 (N_3840,N_3118,N_3298);
nor U3841 (N_3841,N_3230,N_3055);
and U3842 (N_3842,N_3082,N_3071);
nor U3843 (N_3843,N_3425,N_3319);
nor U3844 (N_3844,N_3287,N_3488);
nand U3845 (N_3845,N_3420,N_3457);
nor U3846 (N_3846,N_3174,N_3397);
or U3847 (N_3847,N_3144,N_3290);
nor U3848 (N_3848,N_3074,N_3204);
nor U3849 (N_3849,N_3280,N_3040);
and U3850 (N_3850,N_3274,N_3149);
nand U3851 (N_3851,N_3129,N_3050);
and U3852 (N_3852,N_3029,N_3272);
nand U3853 (N_3853,N_3283,N_3240);
nor U3854 (N_3854,N_3346,N_3168);
or U3855 (N_3855,N_3297,N_3238);
nor U3856 (N_3856,N_3264,N_3355);
nand U3857 (N_3857,N_3449,N_3426);
nand U3858 (N_3858,N_3303,N_3265);
nor U3859 (N_3859,N_3019,N_3229);
or U3860 (N_3860,N_3190,N_3469);
and U3861 (N_3861,N_3385,N_3229);
nand U3862 (N_3862,N_3426,N_3483);
and U3863 (N_3863,N_3000,N_3031);
nor U3864 (N_3864,N_3454,N_3094);
and U3865 (N_3865,N_3120,N_3297);
and U3866 (N_3866,N_3471,N_3208);
nand U3867 (N_3867,N_3463,N_3432);
or U3868 (N_3868,N_3311,N_3364);
and U3869 (N_3869,N_3483,N_3314);
or U3870 (N_3870,N_3244,N_3398);
nand U3871 (N_3871,N_3001,N_3294);
and U3872 (N_3872,N_3043,N_3055);
nand U3873 (N_3873,N_3163,N_3352);
nand U3874 (N_3874,N_3126,N_3092);
nor U3875 (N_3875,N_3377,N_3455);
or U3876 (N_3876,N_3418,N_3085);
or U3877 (N_3877,N_3031,N_3175);
nor U3878 (N_3878,N_3256,N_3234);
and U3879 (N_3879,N_3441,N_3194);
or U3880 (N_3880,N_3209,N_3443);
nand U3881 (N_3881,N_3420,N_3050);
and U3882 (N_3882,N_3482,N_3195);
nor U3883 (N_3883,N_3457,N_3437);
nand U3884 (N_3884,N_3176,N_3251);
and U3885 (N_3885,N_3281,N_3255);
or U3886 (N_3886,N_3498,N_3218);
or U3887 (N_3887,N_3431,N_3410);
nand U3888 (N_3888,N_3086,N_3343);
nand U3889 (N_3889,N_3071,N_3360);
nor U3890 (N_3890,N_3182,N_3442);
nor U3891 (N_3891,N_3313,N_3232);
nand U3892 (N_3892,N_3011,N_3213);
nand U3893 (N_3893,N_3263,N_3485);
and U3894 (N_3894,N_3465,N_3190);
and U3895 (N_3895,N_3087,N_3226);
nor U3896 (N_3896,N_3445,N_3488);
nor U3897 (N_3897,N_3101,N_3147);
and U3898 (N_3898,N_3377,N_3204);
or U3899 (N_3899,N_3138,N_3457);
and U3900 (N_3900,N_3259,N_3495);
or U3901 (N_3901,N_3084,N_3139);
nand U3902 (N_3902,N_3295,N_3140);
or U3903 (N_3903,N_3331,N_3001);
nor U3904 (N_3904,N_3025,N_3091);
and U3905 (N_3905,N_3219,N_3403);
nand U3906 (N_3906,N_3467,N_3278);
nand U3907 (N_3907,N_3328,N_3299);
nor U3908 (N_3908,N_3080,N_3267);
or U3909 (N_3909,N_3346,N_3417);
nor U3910 (N_3910,N_3440,N_3064);
xnor U3911 (N_3911,N_3113,N_3281);
nand U3912 (N_3912,N_3017,N_3359);
and U3913 (N_3913,N_3259,N_3191);
and U3914 (N_3914,N_3416,N_3280);
and U3915 (N_3915,N_3037,N_3423);
nor U3916 (N_3916,N_3411,N_3323);
and U3917 (N_3917,N_3015,N_3173);
nand U3918 (N_3918,N_3306,N_3483);
and U3919 (N_3919,N_3268,N_3366);
nand U3920 (N_3920,N_3000,N_3417);
and U3921 (N_3921,N_3460,N_3229);
or U3922 (N_3922,N_3437,N_3241);
or U3923 (N_3923,N_3387,N_3338);
nor U3924 (N_3924,N_3371,N_3119);
nor U3925 (N_3925,N_3331,N_3250);
and U3926 (N_3926,N_3082,N_3205);
or U3927 (N_3927,N_3313,N_3200);
or U3928 (N_3928,N_3054,N_3262);
nand U3929 (N_3929,N_3316,N_3262);
nor U3930 (N_3930,N_3257,N_3106);
or U3931 (N_3931,N_3483,N_3444);
nor U3932 (N_3932,N_3337,N_3489);
nor U3933 (N_3933,N_3131,N_3423);
and U3934 (N_3934,N_3220,N_3063);
nand U3935 (N_3935,N_3467,N_3283);
or U3936 (N_3936,N_3441,N_3087);
and U3937 (N_3937,N_3016,N_3127);
nand U3938 (N_3938,N_3483,N_3178);
or U3939 (N_3939,N_3332,N_3408);
and U3940 (N_3940,N_3383,N_3313);
nor U3941 (N_3941,N_3374,N_3246);
nand U3942 (N_3942,N_3446,N_3452);
nand U3943 (N_3943,N_3292,N_3069);
nand U3944 (N_3944,N_3029,N_3105);
and U3945 (N_3945,N_3454,N_3341);
or U3946 (N_3946,N_3092,N_3182);
or U3947 (N_3947,N_3461,N_3029);
nand U3948 (N_3948,N_3013,N_3265);
or U3949 (N_3949,N_3462,N_3165);
and U3950 (N_3950,N_3245,N_3107);
or U3951 (N_3951,N_3368,N_3007);
nor U3952 (N_3952,N_3284,N_3069);
nor U3953 (N_3953,N_3431,N_3271);
or U3954 (N_3954,N_3180,N_3209);
or U3955 (N_3955,N_3096,N_3403);
and U3956 (N_3956,N_3119,N_3395);
nor U3957 (N_3957,N_3327,N_3105);
and U3958 (N_3958,N_3459,N_3213);
or U3959 (N_3959,N_3010,N_3009);
nor U3960 (N_3960,N_3091,N_3190);
nand U3961 (N_3961,N_3090,N_3498);
or U3962 (N_3962,N_3172,N_3174);
nand U3963 (N_3963,N_3096,N_3315);
and U3964 (N_3964,N_3468,N_3409);
nor U3965 (N_3965,N_3328,N_3353);
or U3966 (N_3966,N_3379,N_3279);
or U3967 (N_3967,N_3495,N_3327);
nor U3968 (N_3968,N_3165,N_3048);
nand U3969 (N_3969,N_3178,N_3382);
or U3970 (N_3970,N_3214,N_3165);
and U3971 (N_3971,N_3349,N_3410);
nor U3972 (N_3972,N_3201,N_3007);
and U3973 (N_3973,N_3222,N_3480);
nand U3974 (N_3974,N_3450,N_3155);
nor U3975 (N_3975,N_3177,N_3095);
or U3976 (N_3976,N_3270,N_3016);
nor U3977 (N_3977,N_3182,N_3469);
or U3978 (N_3978,N_3062,N_3441);
or U3979 (N_3979,N_3160,N_3278);
or U3980 (N_3980,N_3370,N_3069);
nor U3981 (N_3981,N_3212,N_3420);
nor U3982 (N_3982,N_3025,N_3379);
xor U3983 (N_3983,N_3354,N_3438);
or U3984 (N_3984,N_3148,N_3095);
nor U3985 (N_3985,N_3412,N_3087);
nor U3986 (N_3986,N_3357,N_3058);
nand U3987 (N_3987,N_3140,N_3059);
and U3988 (N_3988,N_3317,N_3347);
and U3989 (N_3989,N_3390,N_3283);
and U3990 (N_3990,N_3207,N_3450);
nor U3991 (N_3991,N_3415,N_3345);
and U3992 (N_3992,N_3186,N_3304);
nand U3993 (N_3993,N_3391,N_3061);
nor U3994 (N_3994,N_3487,N_3411);
or U3995 (N_3995,N_3002,N_3157);
nand U3996 (N_3996,N_3026,N_3211);
nor U3997 (N_3997,N_3034,N_3102);
nor U3998 (N_3998,N_3426,N_3428);
nor U3999 (N_3999,N_3083,N_3279);
or U4000 (N_4000,N_3613,N_3828);
and U4001 (N_4001,N_3797,N_3693);
and U4002 (N_4002,N_3782,N_3692);
and U4003 (N_4003,N_3686,N_3629);
nor U4004 (N_4004,N_3829,N_3976);
nand U4005 (N_4005,N_3521,N_3823);
nor U4006 (N_4006,N_3665,N_3537);
nor U4007 (N_4007,N_3622,N_3577);
nor U4008 (N_4008,N_3887,N_3790);
nand U4009 (N_4009,N_3516,N_3940);
nand U4010 (N_4010,N_3851,N_3654);
or U4011 (N_4011,N_3554,N_3758);
or U4012 (N_4012,N_3566,N_3941);
nor U4013 (N_4013,N_3747,N_3750);
and U4014 (N_4014,N_3520,N_3694);
nand U4015 (N_4015,N_3727,N_3717);
nand U4016 (N_4016,N_3548,N_3738);
nor U4017 (N_4017,N_3610,N_3531);
nor U4018 (N_4018,N_3651,N_3589);
and U4019 (N_4019,N_3700,N_3999);
and U4020 (N_4020,N_3964,N_3988);
nor U4021 (N_4021,N_3615,N_3706);
and U4022 (N_4022,N_3752,N_3663);
nand U4023 (N_4023,N_3619,N_3906);
and U4024 (N_4024,N_3506,N_3594);
xor U4025 (N_4025,N_3898,N_3779);
nand U4026 (N_4026,N_3691,N_3908);
nand U4027 (N_4027,N_3867,N_3839);
and U4028 (N_4028,N_3860,N_3844);
nand U4029 (N_4029,N_3904,N_3592);
and U4030 (N_4030,N_3564,N_3813);
nor U4031 (N_4031,N_3842,N_3715);
and U4032 (N_4032,N_3796,N_3677);
and U4033 (N_4033,N_3518,N_3511);
nor U4034 (N_4034,N_3788,N_3959);
nor U4035 (N_4035,N_3581,N_3659);
nand U4036 (N_4036,N_3556,N_3895);
and U4037 (N_4037,N_3673,N_3640);
nor U4038 (N_4038,N_3504,N_3939);
nor U4039 (N_4039,N_3534,N_3626);
or U4040 (N_4040,N_3536,N_3837);
nand U4041 (N_4041,N_3970,N_3580);
and U4042 (N_4042,N_3757,N_3645);
or U4043 (N_4043,N_3984,N_3962);
or U4044 (N_4044,N_3967,N_3523);
and U4045 (N_4045,N_3890,N_3910);
nand U4046 (N_4046,N_3668,N_3666);
nor U4047 (N_4047,N_3912,N_3740);
or U4048 (N_4048,N_3869,N_3771);
nand U4049 (N_4049,N_3990,N_3917);
nand U4050 (N_4050,N_3925,N_3816);
or U4051 (N_4051,N_3878,N_3558);
or U4052 (N_4052,N_3835,N_3633);
nand U4053 (N_4053,N_3948,N_3679);
nor U4054 (N_4054,N_3944,N_3896);
nand U4055 (N_4055,N_3606,N_3625);
and U4056 (N_4056,N_3932,N_3923);
or U4057 (N_4057,N_3689,N_3522);
nor U4058 (N_4058,N_3563,N_3934);
or U4059 (N_4059,N_3911,N_3726);
nor U4060 (N_4060,N_3876,N_3731);
nand U4061 (N_4061,N_3593,N_3525);
or U4062 (N_4062,N_3517,N_3781);
nor U4063 (N_4063,N_3817,N_3560);
or U4064 (N_4064,N_3831,N_3724);
nor U4065 (N_4065,N_3818,N_3950);
or U4066 (N_4066,N_3682,N_3996);
or U4067 (N_4067,N_3840,N_3968);
nor U4068 (N_4068,N_3672,N_3985);
or U4069 (N_4069,N_3576,N_3685);
or U4070 (N_4070,N_3684,N_3500);
or U4071 (N_4071,N_3883,N_3768);
nand U4072 (N_4072,N_3922,N_3725);
nand U4073 (N_4073,N_3528,N_3765);
or U4074 (N_4074,N_3667,N_3637);
nor U4075 (N_4075,N_3688,N_3756);
nand U4076 (N_4076,N_3703,N_3600);
nand U4077 (N_4077,N_3760,N_3822);
and U4078 (N_4078,N_3671,N_3928);
and U4079 (N_4079,N_3572,N_3872);
and U4080 (N_4080,N_3643,N_3845);
nor U4081 (N_4081,N_3529,N_3841);
nand U4082 (N_4082,N_3924,N_3893);
and U4083 (N_4083,N_3949,N_3761);
xnor U4084 (N_4084,N_3510,N_3854);
nand U4085 (N_4085,N_3656,N_3705);
or U4086 (N_4086,N_3798,N_3561);
nand U4087 (N_4087,N_3855,N_3743);
or U4088 (N_4088,N_3834,N_3826);
nor U4089 (N_4089,N_3609,N_3721);
or U4090 (N_4090,N_3591,N_3951);
and U4091 (N_4091,N_3824,N_3960);
and U4092 (N_4092,N_3929,N_3870);
or U4093 (N_4093,N_3909,N_3644);
or U4094 (N_4094,N_3859,N_3567);
or U4095 (N_4095,N_3555,N_3601);
or U4096 (N_4096,N_3545,N_3992);
nand U4097 (N_4097,N_3966,N_3995);
nand U4098 (N_4098,N_3612,N_3819);
nand U4099 (N_4099,N_3736,N_3820);
nand U4100 (N_4100,N_3713,N_3806);
and U4101 (N_4101,N_3695,N_3604);
or U4102 (N_4102,N_3739,N_3975);
or U4103 (N_4103,N_3920,N_3642);
nor U4104 (N_4104,N_3772,N_3596);
or U4105 (N_4105,N_3954,N_3579);
nand U4106 (N_4106,N_3956,N_3857);
nand U4107 (N_4107,N_3569,N_3546);
nand U4108 (N_4108,N_3681,N_3658);
and U4109 (N_4109,N_3570,N_3778);
and U4110 (N_4110,N_3568,N_3864);
or U4111 (N_4111,N_3884,N_3707);
or U4112 (N_4112,N_3852,N_3661);
or U4113 (N_4113,N_3955,N_3942);
or U4114 (N_4114,N_3755,N_3540);
nor U4115 (N_4115,N_3698,N_3833);
and U4116 (N_4116,N_3542,N_3557);
or U4117 (N_4117,N_3914,N_3611);
nor U4118 (N_4118,N_3512,N_3926);
and U4119 (N_4119,N_3730,N_3897);
or U4120 (N_4120,N_3605,N_3565);
or U4121 (N_4121,N_3571,N_3935);
nor U4122 (N_4122,N_3623,N_3957);
nor U4123 (N_4123,N_3735,N_3550);
nand U4124 (N_4124,N_3802,N_3662);
and U4125 (N_4125,N_3687,N_3972);
nor U4126 (N_4126,N_3903,N_3649);
and U4127 (N_4127,N_3608,N_3745);
and U4128 (N_4128,N_3514,N_3748);
nand U4129 (N_4129,N_3559,N_3858);
nor U4130 (N_4130,N_3582,N_3916);
nor U4131 (N_4131,N_3775,N_3921);
or U4132 (N_4132,N_3762,N_3809);
or U4133 (N_4133,N_3991,N_3902);
and U4134 (N_4134,N_3888,N_3751);
nand U4135 (N_4135,N_3795,N_3807);
nand U4136 (N_4136,N_3746,N_3527);
or U4137 (N_4137,N_3821,N_3657);
and U4138 (N_4138,N_3804,N_3501);
nor U4139 (N_4139,N_3803,N_3543);
and U4140 (N_4140,N_3843,N_3513);
and U4141 (N_4141,N_3614,N_3899);
and U4142 (N_4142,N_3936,N_3862);
xor U4143 (N_4143,N_3575,N_3590);
nand U4144 (N_4144,N_3723,N_3764);
nand U4145 (N_4145,N_3616,N_3709);
xor U4146 (N_4146,N_3509,N_3598);
or U4147 (N_4147,N_3719,N_3793);
or U4148 (N_4148,N_3722,N_3907);
nand U4149 (N_4149,N_3552,N_3982);
nor U4150 (N_4150,N_3507,N_3763);
nor U4151 (N_4151,N_3749,N_3850);
or U4152 (N_4152,N_3866,N_3676);
and U4153 (N_4153,N_3786,N_3639);
and U4154 (N_4154,N_3573,N_3635);
and U4155 (N_4155,N_3885,N_3986);
nand U4156 (N_4156,N_3503,N_3958);
nand U4157 (N_4157,N_3541,N_3508);
and U4158 (N_4158,N_3838,N_3718);
and U4159 (N_4159,N_3627,N_3690);
and U4160 (N_4160,N_3787,N_3947);
nor U4161 (N_4161,N_3800,N_3825);
or U4162 (N_4162,N_3767,N_3773);
nor U4163 (N_4163,N_3994,N_3776);
or U4164 (N_4164,N_3953,N_3544);
or U4165 (N_4165,N_3938,N_3987);
and U4166 (N_4166,N_3997,N_3785);
nor U4167 (N_4167,N_3549,N_3993);
or U4168 (N_4168,N_3524,N_3946);
and U4169 (N_4169,N_3965,N_3647);
xor U4170 (N_4170,N_3583,N_3653);
or U4171 (N_4171,N_3810,N_3780);
nor U4172 (N_4172,N_3728,N_3894);
nand U4173 (N_4173,N_3704,N_3539);
nand U4174 (N_4174,N_3905,N_3562);
or U4175 (N_4175,N_3979,N_3634);
nand U4176 (N_4176,N_3930,N_3770);
and U4177 (N_4177,N_3597,N_3865);
and U4178 (N_4178,N_3853,N_3660);
nand U4179 (N_4179,N_3879,N_3836);
nor U4180 (N_4180,N_3849,N_3900);
and U4181 (N_4181,N_3873,N_3814);
nor U4182 (N_4182,N_3599,N_3961);
nand U4183 (N_4183,N_3710,N_3526);
nor U4184 (N_4184,N_3641,N_3714);
and U4185 (N_4185,N_3670,N_3505);
nand U4186 (N_4186,N_3980,N_3655);
or U4187 (N_4187,N_3981,N_3766);
nor U4188 (N_4188,N_3875,N_3880);
nor U4189 (N_4189,N_3532,N_3881);
nor U4190 (N_4190,N_3618,N_3812);
nor U4191 (N_4191,N_3733,N_3978);
and U4192 (N_4192,N_3886,N_3919);
or U4193 (N_4193,N_3547,N_3551);
and U4194 (N_4194,N_3784,N_3701);
and U4195 (N_4195,N_3650,N_3732);
and U4196 (N_4196,N_3753,N_3519);
and U4197 (N_4197,N_3848,N_3933);
nor U4198 (N_4198,N_3617,N_3533);
nor U4199 (N_4199,N_3502,N_3832);
nand U4200 (N_4200,N_3791,N_3977);
nor U4201 (N_4201,N_3607,N_3553);
nor U4202 (N_4202,N_3774,N_3595);
and U4203 (N_4203,N_3631,N_3963);
nor U4204 (N_4204,N_3587,N_3892);
nor U4205 (N_4205,N_3603,N_3734);
nor U4206 (N_4206,N_3801,N_3901);
nand U4207 (N_4207,N_3874,N_3863);
nor U4208 (N_4208,N_3696,N_3877);
nand U4209 (N_4209,N_3646,N_3846);
xnor U4210 (N_4210,N_3669,N_3871);
nand U4211 (N_4211,N_3769,N_3530);
nand U4212 (N_4212,N_3983,N_3868);
or U4213 (N_4213,N_3811,N_3712);
or U4214 (N_4214,N_3973,N_3620);
nand U4215 (N_4215,N_3621,N_3711);
and U4216 (N_4216,N_3638,N_3515);
and U4217 (N_4217,N_3585,N_3808);
or U4218 (N_4218,N_3927,N_3989);
nor U4219 (N_4219,N_3754,N_3856);
nor U4220 (N_4220,N_3974,N_3729);
nand U4221 (N_4221,N_3584,N_3943);
nor U4222 (N_4222,N_3759,N_3624);
or U4223 (N_4223,N_3588,N_3716);
nor U4224 (N_4224,N_3889,N_3815);
and U4225 (N_4225,N_3799,N_3805);
nor U4226 (N_4226,N_3697,N_3737);
or U4227 (N_4227,N_3702,N_3648);
or U4228 (N_4228,N_3792,N_3783);
nand U4229 (N_4229,N_3861,N_3952);
and U4230 (N_4230,N_3636,N_3538);
and U4231 (N_4231,N_3891,N_3602);
and U4232 (N_4232,N_3586,N_3789);
nor U4233 (N_4233,N_3674,N_3915);
or U4234 (N_4234,N_3741,N_3777);
nand U4235 (N_4235,N_3630,N_3913);
nor U4236 (N_4236,N_3998,N_3742);
and U4237 (N_4237,N_3937,N_3664);
nand U4238 (N_4238,N_3720,N_3971);
and U4239 (N_4239,N_3628,N_3847);
and U4240 (N_4240,N_3931,N_3683);
nand U4241 (N_4241,N_3830,N_3632);
and U4242 (N_4242,N_3969,N_3574);
nor U4243 (N_4243,N_3794,N_3678);
or U4244 (N_4244,N_3680,N_3578);
nand U4245 (N_4245,N_3652,N_3699);
or U4246 (N_4246,N_3535,N_3708);
or U4247 (N_4247,N_3827,N_3675);
nor U4248 (N_4248,N_3882,N_3744);
and U4249 (N_4249,N_3918,N_3945);
and U4250 (N_4250,N_3657,N_3570);
or U4251 (N_4251,N_3558,N_3542);
nor U4252 (N_4252,N_3630,N_3932);
and U4253 (N_4253,N_3581,N_3809);
xnor U4254 (N_4254,N_3588,N_3755);
nor U4255 (N_4255,N_3938,N_3546);
nand U4256 (N_4256,N_3698,N_3790);
nor U4257 (N_4257,N_3905,N_3637);
or U4258 (N_4258,N_3880,N_3537);
and U4259 (N_4259,N_3709,N_3634);
and U4260 (N_4260,N_3685,N_3643);
xor U4261 (N_4261,N_3800,N_3730);
nor U4262 (N_4262,N_3613,N_3713);
nor U4263 (N_4263,N_3623,N_3874);
nand U4264 (N_4264,N_3914,N_3643);
and U4265 (N_4265,N_3906,N_3716);
nand U4266 (N_4266,N_3623,N_3678);
or U4267 (N_4267,N_3885,N_3936);
nor U4268 (N_4268,N_3533,N_3952);
nor U4269 (N_4269,N_3556,N_3546);
nor U4270 (N_4270,N_3986,N_3948);
nand U4271 (N_4271,N_3623,N_3538);
nand U4272 (N_4272,N_3984,N_3881);
nand U4273 (N_4273,N_3595,N_3865);
nor U4274 (N_4274,N_3804,N_3891);
nand U4275 (N_4275,N_3836,N_3568);
nor U4276 (N_4276,N_3854,N_3895);
nand U4277 (N_4277,N_3500,N_3870);
or U4278 (N_4278,N_3759,N_3807);
nor U4279 (N_4279,N_3864,N_3855);
nor U4280 (N_4280,N_3993,N_3971);
or U4281 (N_4281,N_3712,N_3827);
nor U4282 (N_4282,N_3656,N_3608);
and U4283 (N_4283,N_3974,N_3804);
or U4284 (N_4284,N_3751,N_3537);
or U4285 (N_4285,N_3683,N_3885);
xor U4286 (N_4286,N_3912,N_3738);
nor U4287 (N_4287,N_3881,N_3768);
and U4288 (N_4288,N_3979,N_3724);
and U4289 (N_4289,N_3615,N_3651);
nor U4290 (N_4290,N_3605,N_3688);
nand U4291 (N_4291,N_3852,N_3928);
nor U4292 (N_4292,N_3917,N_3532);
or U4293 (N_4293,N_3734,N_3978);
nor U4294 (N_4294,N_3517,N_3629);
nor U4295 (N_4295,N_3843,N_3784);
nand U4296 (N_4296,N_3860,N_3576);
nor U4297 (N_4297,N_3663,N_3697);
and U4298 (N_4298,N_3516,N_3655);
nor U4299 (N_4299,N_3542,N_3733);
or U4300 (N_4300,N_3735,N_3996);
nand U4301 (N_4301,N_3573,N_3792);
or U4302 (N_4302,N_3968,N_3786);
nor U4303 (N_4303,N_3763,N_3521);
nand U4304 (N_4304,N_3759,N_3984);
and U4305 (N_4305,N_3819,N_3789);
or U4306 (N_4306,N_3586,N_3702);
and U4307 (N_4307,N_3836,N_3690);
nor U4308 (N_4308,N_3918,N_3511);
nand U4309 (N_4309,N_3851,N_3539);
or U4310 (N_4310,N_3587,N_3696);
nor U4311 (N_4311,N_3843,N_3737);
nor U4312 (N_4312,N_3946,N_3862);
nor U4313 (N_4313,N_3979,N_3534);
or U4314 (N_4314,N_3545,N_3865);
or U4315 (N_4315,N_3683,N_3966);
nand U4316 (N_4316,N_3669,N_3881);
or U4317 (N_4317,N_3706,N_3502);
or U4318 (N_4318,N_3677,N_3888);
and U4319 (N_4319,N_3610,N_3659);
and U4320 (N_4320,N_3985,N_3993);
or U4321 (N_4321,N_3625,N_3577);
and U4322 (N_4322,N_3502,N_3587);
nand U4323 (N_4323,N_3571,N_3517);
nor U4324 (N_4324,N_3596,N_3578);
nand U4325 (N_4325,N_3880,N_3994);
or U4326 (N_4326,N_3910,N_3501);
and U4327 (N_4327,N_3973,N_3660);
and U4328 (N_4328,N_3700,N_3575);
nor U4329 (N_4329,N_3865,N_3660);
nand U4330 (N_4330,N_3703,N_3572);
nor U4331 (N_4331,N_3540,N_3990);
nand U4332 (N_4332,N_3695,N_3968);
nor U4333 (N_4333,N_3735,N_3513);
nand U4334 (N_4334,N_3757,N_3822);
nor U4335 (N_4335,N_3604,N_3932);
nor U4336 (N_4336,N_3504,N_3544);
and U4337 (N_4337,N_3849,N_3650);
and U4338 (N_4338,N_3621,N_3692);
and U4339 (N_4339,N_3899,N_3633);
or U4340 (N_4340,N_3928,N_3947);
or U4341 (N_4341,N_3516,N_3737);
nor U4342 (N_4342,N_3753,N_3585);
nand U4343 (N_4343,N_3538,N_3612);
or U4344 (N_4344,N_3646,N_3771);
nand U4345 (N_4345,N_3883,N_3525);
nand U4346 (N_4346,N_3686,N_3595);
nor U4347 (N_4347,N_3955,N_3649);
nor U4348 (N_4348,N_3538,N_3586);
and U4349 (N_4349,N_3978,N_3987);
or U4350 (N_4350,N_3772,N_3696);
nand U4351 (N_4351,N_3576,N_3839);
or U4352 (N_4352,N_3806,N_3776);
or U4353 (N_4353,N_3591,N_3703);
nand U4354 (N_4354,N_3511,N_3957);
or U4355 (N_4355,N_3719,N_3966);
or U4356 (N_4356,N_3747,N_3826);
nand U4357 (N_4357,N_3680,N_3601);
nor U4358 (N_4358,N_3800,N_3799);
or U4359 (N_4359,N_3884,N_3987);
and U4360 (N_4360,N_3520,N_3945);
nand U4361 (N_4361,N_3998,N_3997);
nor U4362 (N_4362,N_3855,N_3825);
and U4363 (N_4363,N_3610,N_3804);
nand U4364 (N_4364,N_3718,N_3756);
nor U4365 (N_4365,N_3800,N_3624);
and U4366 (N_4366,N_3996,N_3597);
nor U4367 (N_4367,N_3946,N_3581);
or U4368 (N_4368,N_3796,N_3940);
or U4369 (N_4369,N_3585,N_3809);
or U4370 (N_4370,N_3540,N_3756);
and U4371 (N_4371,N_3805,N_3993);
or U4372 (N_4372,N_3807,N_3705);
nand U4373 (N_4373,N_3877,N_3873);
nor U4374 (N_4374,N_3819,N_3513);
and U4375 (N_4375,N_3601,N_3578);
nand U4376 (N_4376,N_3952,N_3523);
and U4377 (N_4377,N_3910,N_3824);
nor U4378 (N_4378,N_3814,N_3588);
nor U4379 (N_4379,N_3680,N_3644);
nor U4380 (N_4380,N_3921,N_3553);
nand U4381 (N_4381,N_3981,N_3824);
nor U4382 (N_4382,N_3513,N_3979);
nor U4383 (N_4383,N_3656,N_3939);
and U4384 (N_4384,N_3877,N_3579);
and U4385 (N_4385,N_3715,N_3654);
or U4386 (N_4386,N_3658,N_3892);
nand U4387 (N_4387,N_3944,N_3568);
nor U4388 (N_4388,N_3610,N_3598);
and U4389 (N_4389,N_3855,N_3845);
or U4390 (N_4390,N_3994,N_3795);
and U4391 (N_4391,N_3732,N_3991);
nand U4392 (N_4392,N_3589,N_3715);
nor U4393 (N_4393,N_3989,N_3706);
nor U4394 (N_4394,N_3682,N_3799);
or U4395 (N_4395,N_3826,N_3995);
and U4396 (N_4396,N_3648,N_3563);
nand U4397 (N_4397,N_3605,N_3967);
and U4398 (N_4398,N_3618,N_3891);
and U4399 (N_4399,N_3734,N_3558);
and U4400 (N_4400,N_3843,N_3635);
nor U4401 (N_4401,N_3733,N_3614);
nand U4402 (N_4402,N_3774,N_3841);
or U4403 (N_4403,N_3905,N_3877);
nor U4404 (N_4404,N_3698,N_3787);
or U4405 (N_4405,N_3612,N_3948);
nand U4406 (N_4406,N_3680,N_3751);
nor U4407 (N_4407,N_3896,N_3681);
nor U4408 (N_4408,N_3922,N_3890);
or U4409 (N_4409,N_3941,N_3998);
nand U4410 (N_4410,N_3869,N_3648);
nand U4411 (N_4411,N_3692,N_3877);
and U4412 (N_4412,N_3546,N_3832);
or U4413 (N_4413,N_3913,N_3747);
nand U4414 (N_4414,N_3622,N_3832);
or U4415 (N_4415,N_3967,N_3543);
or U4416 (N_4416,N_3586,N_3613);
xor U4417 (N_4417,N_3636,N_3988);
nor U4418 (N_4418,N_3984,N_3514);
and U4419 (N_4419,N_3768,N_3844);
and U4420 (N_4420,N_3964,N_3797);
nor U4421 (N_4421,N_3964,N_3528);
and U4422 (N_4422,N_3522,N_3644);
or U4423 (N_4423,N_3783,N_3595);
nand U4424 (N_4424,N_3959,N_3732);
and U4425 (N_4425,N_3693,N_3989);
or U4426 (N_4426,N_3926,N_3762);
nor U4427 (N_4427,N_3764,N_3961);
or U4428 (N_4428,N_3681,N_3902);
and U4429 (N_4429,N_3641,N_3868);
nand U4430 (N_4430,N_3569,N_3829);
or U4431 (N_4431,N_3922,N_3777);
or U4432 (N_4432,N_3852,N_3916);
nor U4433 (N_4433,N_3844,N_3549);
or U4434 (N_4434,N_3572,N_3674);
and U4435 (N_4435,N_3940,N_3630);
nor U4436 (N_4436,N_3976,N_3900);
nand U4437 (N_4437,N_3565,N_3952);
nor U4438 (N_4438,N_3664,N_3548);
or U4439 (N_4439,N_3955,N_3944);
nor U4440 (N_4440,N_3868,N_3668);
nand U4441 (N_4441,N_3668,N_3550);
nand U4442 (N_4442,N_3537,N_3980);
nor U4443 (N_4443,N_3783,N_3768);
and U4444 (N_4444,N_3565,N_3621);
or U4445 (N_4445,N_3924,N_3683);
and U4446 (N_4446,N_3834,N_3858);
nor U4447 (N_4447,N_3808,N_3662);
nand U4448 (N_4448,N_3756,N_3788);
or U4449 (N_4449,N_3579,N_3928);
or U4450 (N_4450,N_3991,N_3584);
nor U4451 (N_4451,N_3887,N_3676);
nand U4452 (N_4452,N_3500,N_3566);
and U4453 (N_4453,N_3654,N_3977);
or U4454 (N_4454,N_3604,N_3979);
and U4455 (N_4455,N_3776,N_3983);
nor U4456 (N_4456,N_3735,N_3945);
nand U4457 (N_4457,N_3551,N_3548);
or U4458 (N_4458,N_3686,N_3844);
nor U4459 (N_4459,N_3981,N_3857);
nor U4460 (N_4460,N_3660,N_3774);
nor U4461 (N_4461,N_3603,N_3598);
and U4462 (N_4462,N_3845,N_3997);
nand U4463 (N_4463,N_3744,N_3654);
and U4464 (N_4464,N_3573,N_3577);
nand U4465 (N_4465,N_3605,N_3734);
nand U4466 (N_4466,N_3728,N_3786);
and U4467 (N_4467,N_3723,N_3998);
or U4468 (N_4468,N_3910,N_3636);
and U4469 (N_4469,N_3960,N_3859);
nor U4470 (N_4470,N_3583,N_3723);
or U4471 (N_4471,N_3547,N_3898);
nor U4472 (N_4472,N_3637,N_3776);
or U4473 (N_4473,N_3654,N_3926);
nand U4474 (N_4474,N_3648,N_3502);
nand U4475 (N_4475,N_3940,N_3809);
or U4476 (N_4476,N_3785,N_3664);
nor U4477 (N_4477,N_3770,N_3829);
and U4478 (N_4478,N_3820,N_3976);
nor U4479 (N_4479,N_3507,N_3742);
and U4480 (N_4480,N_3551,N_3812);
nand U4481 (N_4481,N_3890,N_3982);
nor U4482 (N_4482,N_3884,N_3650);
nor U4483 (N_4483,N_3504,N_3552);
and U4484 (N_4484,N_3524,N_3917);
nand U4485 (N_4485,N_3910,N_3723);
nand U4486 (N_4486,N_3956,N_3755);
nor U4487 (N_4487,N_3955,N_3572);
nand U4488 (N_4488,N_3955,N_3620);
and U4489 (N_4489,N_3872,N_3603);
and U4490 (N_4490,N_3783,N_3517);
nand U4491 (N_4491,N_3568,N_3650);
nor U4492 (N_4492,N_3526,N_3889);
and U4493 (N_4493,N_3522,N_3637);
nand U4494 (N_4494,N_3585,N_3806);
or U4495 (N_4495,N_3779,N_3962);
and U4496 (N_4496,N_3869,N_3794);
and U4497 (N_4497,N_3691,N_3874);
nor U4498 (N_4498,N_3897,N_3959);
nand U4499 (N_4499,N_3588,N_3511);
or U4500 (N_4500,N_4351,N_4137);
and U4501 (N_4501,N_4101,N_4222);
nand U4502 (N_4502,N_4205,N_4200);
or U4503 (N_4503,N_4343,N_4053);
and U4504 (N_4504,N_4006,N_4297);
xor U4505 (N_4505,N_4023,N_4198);
nand U4506 (N_4506,N_4376,N_4044);
nor U4507 (N_4507,N_4307,N_4031);
nand U4508 (N_4508,N_4496,N_4319);
nor U4509 (N_4509,N_4258,N_4158);
nor U4510 (N_4510,N_4471,N_4194);
or U4511 (N_4511,N_4466,N_4163);
nor U4512 (N_4512,N_4264,N_4040);
and U4513 (N_4513,N_4089,N_4227);
nand U4514 (N_4514,N_4456,N_4396);
or U4515 (N_4515,N_4363,N_4488);
or U4516 (N_4516,N_4132,N_4027);
nand U4517 (N_4517,N_4094,N_4315);
or U4518 (N_4518,N_4393,N_4398);
and U4519 (N_4519,N_4468,N_4131);
or U4520 (N_4520,N_4026,N_4388);
nand U4521 (N_4521,N_4331,N_4152);
and U4522 (N_4522,N_4417,N_4107);
or U4523 (N_4523,N_4123,N_4165);
or U4524 (N_4524,N_4216,N_4430);
and U4525 (N_4525,N_4408,N_4321);
nor U4526 (N_4526,N_4234,N_4074);
nor U4527 (N_4527,N_4223,N_4025);
and U4528 (N_4528,N_4405,N_4486);
or U4529 (N_4529,N_4374,N_4356);
nor U4530 (N_4530,N_4231,N_4141);
nand U4531 (N_4531,N_4279,N_4059);
and U4532 (N_4532,N_4220,N_4497);
nand U4533 (N_4533,N_4328,N_4483);
and U4534 (N_4534,N_4291,N_4447);
nor U4535 (N_4535,N_4326,N_4047);
nand U4536 (N_4536,N_4353,N_4125);
nand U4537 (N_4537,N_4282,N_4359);
nor U4538 (N_4538,N_4357,N_4401);
and U4539 (N_4539,N_4117,N_4365);
and U4540 (N_4540,N_4247,N_4176);
nand U4541 (N_4541,N_4085,N_4358);
or U4542 (N_4542,N_4428,N_4229);
nand U4543 (N_4543,N_4270,N_4219);
and U4544 (N_4544,N_4453,N_4492);
nor U4545 (N_4545,N_4221,N_4450);
nor U4546 (N_4546,N_4467,N_4436);
and U4547 (N_4547,N_4314,N_4173);
nand U4548 (N_4548,N_4061,N_4160);
nand U4549 (N_4549,N_4201,N_4440);
or U4550 (N_4550,N_4364,N_4338);
nor U4551 (N_4551,N_4480,N_4341);
nand U4552 (N_4552,N_4278,N_4499);
or U4553 (N_4553,N_4369,N_4469);
nand U4554 (N_4554,N_4087,N_4170);
nand U4555 (N_4555,N_4057,N_4442);
nand U4556 (N_4556,N_4213,N_4275);
nor U4557 (N_4557,N_4241,N_4427);
and U4558 (N_4558,N_4254,N_4419);
and U4559 (N_4559,N_4106,N_4460);
and U4560 (N_4560,N_4204,N_4407);
or U4561 (N_4561,N_4140,N_4082);
nand U4562 (N_4562,N_4009,N_4235);
or U4563 (N_4563,N_4086,N_4049);
nor U4564 (N_4564,N_4293,N_4155);
and U4565 (N_4565,N_4064,N_4373);
or U4566 (N_4566,N_4146,N_4084);
or U4567 (N_4567,N_4120,N_4295);
nor U4568 (N_4568,N_4413,N_4102);
and U4569 (N_4569,N_4475,N_4304);
nor U4570 (N_4570,N_4178,N_4001);
nand U4571 (N_4571,N_4323,N_4362);
xor U4572 (N_4572,N_4072,N_4010);
nor U4573 (N_4573,N_4179,N_4016);
nor U4574 (N_4574,N_4199,N_4210);
nor U4575 (N_4575,N_4252,N_4150);
and U4576 (N_4576,N_4193,N_4237);
or U4577 (N_4577,N_4069,N_4448);
and U4578 (N_4578,N_4281,N_4415);
and U4579 (N_4579,N_4112,N_4077);
or U4580 (N_4580,N_4138,N_4144);
nor U4581 (N_4581,N_4133,N_4259);
or U4582 (N_4582,N_4156,N_4246);
and U4583 (N_4583,N_4286,N_4379);
or U4584 (N_4584,N_4352,N_4377);
or U4585 (N_4585,N_4294,N_4498);
nor U4586 (N_4586,N_4402,N_4230);
and U4587 (N_4587,N_4113,N_4370);
nand U4588 (N_4588,N_4105,N_4142);
nor U4589 (N_4589,N_4092,N_4301);
and U4590 (N_4590,N_4147,N_4269);
nand U4591 (N_4591,N_4476,N_4285);
nor U4592 (N_4592,N_4245,N_4439);
nor U4593 (N_4593,N_4096,N_4070);
nor U4594 (N_4594,N_4477,N_4065);
nor U4595 (N_4595,N_4090,N_4083);
nor U4596 (N_4596,N_4330,N_4325);
and U4597 (N_4597,N_4148,N_4349);
nor U4598 (N_4598,N_4055,N_4303);
or U4599 (N_4599,N_4067,N_4244);
and U4600 (N_4600,N_4175,N_4122);
nor U4601 (N_4601,N_4197,N_4078);
or U4602 (N_4602,N_4076,N_4186);
and U4603 (N_4603,N_4190,N_4028);
or U4604 (N_4604,N_4214,N_4313);
or U4605 (N_4605,N_4350,N_4260);
nand U4606 (N_4606,N_4273,N_4161);
or U4607 (N_4607,N_4397,N_4038);
and U4608 (N_4608,N_4015,N_4143);
nor U4609 (N_4609,N_4494,N_4491);
nor U4610 (N_4610,N_4149,N_4042);
xor U4611 (N_4611,N_4058,N_4110);
nor U4612 (N_4612,N_4354,N_4322);
or U4613 (N_4613,N_4207,N_4139);
or U4614 (N_4614,N_4045,N_4075);
nor U4615 (N_4615,N_4262,N_4462);
nand U4616 (N_4616,N_4103,N_4212);
nand U4617 (N_4617,N_4167,N_4181);
nand U4618 (N_4618,N_4274,N_4024);
and U4619 (N_4619,N_4288,N_4432);
nor U4620 (N_4620,N_4030,N_4206);
nand U4621 (N_4621,N_4154,N_4451);
nand U4622 (N_4622,N_4290,N_4080);
and U4623 (N_4623,N_4253,N_4433);
nor U4624 (N_4624,N_4097,N_4337);
and U4625 (N_4625,N_4126,N_4265);
nor U4626 (N_4626,N_4479,N_4118);
nor U4627 (N_4627,N_4127,N_4162);
and U4628 (N_4628,N_4386,N_4056);
nor U4629 (N_4629,N_4021,N_4403);
nor U4630 (N_4630,N_4425,N_4151);
nor U4631 (N_4631,N_4159,N_4284);
or U4632 (N_4632,N_4052,N_4478);
or U4633 (N_4633,N_4355,N_4302);
nand U4634 (N_4634,N_4007,N_4366);
nor U4635 (N_4635,N_4130,N_4164);
nor U4636 (N_4636,N_4215,N_4093);
nor U4637 (N_4637,N_4342,N_4283);
and U4638 (N_4638,N_4232,N_4458);
and U4639 (N_4639,N_4005,N_4088);
and U4640 (N_4640,N_4012,N_4261);
nor U4641 (N_4641,N_4431,N_4412);
and U4642 (N_4642,N_4034,N_4449);
nand U4643 (N_4643,N_4404,N_4188);
nor U4644 (N_4644,N_4424,N_4043);
and U4645 (N_4645,N_4111,N_4224);
and U4646 (N_4646,N_4387,N_4312);
or U4647 (N_4647,N_4276,N_4367);
nor U4648 (N_4648,N_4251,N_4166);
or U4649 (N_4649,N_4004,N_4305);
or U4650 (N_4650,N_4172,N_4384);
nor U4651 (N_4651,N_4310,N_4033);
nand U4652 (N_4652,N_4320,N_4309);
or U4653 (N_4653,N_4203,N_4434);
or U4654 (N_4654,N_4184,N_4060);
or U4655 (N_4655,N_4375,N_4240);
or U4656 (N_4656,N_4036,N_4109);
nand U4657 (N_4657,N_4192,N_4134);
and U4658 (N_4658,N_4124,N_4311);
nand U4659 (N_4659,N_4287,N_4421);
and U4660 (N_4660,N_4062,N_4454);
or U4661 (N_4661,N_4266,N_4068);
nor U4662 (N_4662,N_4243,N_4029);
and U4663 (N_4663,N_4298,N_4187);
xnor U4664 (N_4664,N_4063,N_4228);
nand U4665 (N_4665,N_4332,N_4128);
nor U4666 (N_4666,N_4100,N_4344);
nand U4667 (N_4667,N_4002,N_4390);
and U4668 (N_4668,N_4169,N_4463);
xnor U4669 (N_4669,N_4493,N_4054);
nand U4670 (N_4670,N_4416,N_4255);
and U4671 (N_4671,N_4037,N_4180);
or U4672 (N_4672,N_4014,N_4066);
nand U4673 (N_4673,N_4019,N_4098);
nor U4674 (N_4674,N_4115,N_4385);
or U4675 (N_4675,N_4108,N_4008);
nand U4676 (N_4676,N_4300,N_4153);
nor U4677 (N_4677,N_4202,N_4461);
nand U4678 (N_4678,N_4383,N_4095);
nand U4679 (N_4679,N_4423,N_4104);
and U4680 (N_4680,N_4368,N_4011);
or U4681 (N_4681,N_4444,N_4272);
nand U4682 (N_4682,N_4437,N_4168);
nor U4683 (N_4683,N_4073,N_4081);
nand U4684 (N_4684,N_4429,N_4211);
nand U4685 (N_4685,N_4399,N_4372);
nor U4686 (N_4686,N_4474,N_4316);
or U4687 (N_4687,N_4348,N_4380);
and U4688 (N_4688,N_4324,N_4459);
nor U4689 (N_4689,N_4361,N_4490);
nor U4690 (N_4690,N_4329,N_4406);
or U4691 (N_4691,N_4400,N_4487);
or U4692 (N_4692,N_4017,N_4418);
and U4693 (N_4693,N_4182,N_4345);
nand U4694 (N_4694,N_4336,N_4422);
nand U4695 (N_4695,N_4195,N_4157);
nand U4696 (N_4696,N_4382,N_4208);
or U4697 (N_4697,N_4389,N_4420);
and U4698 (N_4698,N_4317,N_4267);
xnor U4699 (N_4699,N_4177,N_4039);
and U4700 (N_4700,N_4051,N_4013);
or U4701 (N_4701,N_4472,N_4189);
and U4702 (N_4702,N_4046,N_4116);
nor U4703 (N_4703,N_4426,N_4174);
nand U4704 (N_4704,N_4292,N_4409);
nor U4705 (N_4705,N_4018,N_4308);
and U4706 (N_4706,N_4340,N_4257);
or U4707 (N_4707,N_4091,N_4136);
and U4708 (N_4708,N_4000,N_4035);
nand U4709 (N_4709,N_4347,N_4470);
or U4710 (N_4710,N_4296,N_4183);
and U4711 (N_4711,N_4452,N_4414);
and U4712 (N_4712,N_4495,N_4289);
nand U4713 (N_4713,N_4489,N_4242);
nand U4714 (N_4714,N_4263,N_4022);
and U4715 (N_4715,N_4248,N_4339);
nor U4716 (N_4716,N_4438,N_4225);
nand U4717 (N_4717,N_4135,N_4238);
nor U4718 (N_4718,N_4482,N_4171);
nand U4719 (N_4719,N_4119,N_4020);
or U4720 (N_4720,N_4334,N_4129);
or U4721 (N_4721,N_4327,N_4236);
or U4722 (N_4722,N_4455,N_4071);
nand U4723 (N_4723,N_4465,N_4485);
nor U4724 (N_4724,N_4209,N_4391);
and U4725 (N_4725,N_4277,N_4395);
nand U4726 (N_4726,N_4185,N_4280);
nand U4727 (N_4727,N_4333,N_4239);
nand U4728 (N_4728,N_4464,N_4360);
nand U4729 (N_4729,N_4218,N_4256);
nor U4730 (N_4730,N_4378,N_4445);
or U4731 (N_4731,N_4003,N_4196);
or U4732 (N_4732,N_4217,N_4032);
and U4733 (N_4733,N_4233,N_4318);
or U4734 (N_4734,N_4145,N_4048);
or U4735 (N_4735,N_4441,N_4457);
or U4736 (N_4736,N_4121,N_4099);
nand U4737 (N_4737,N_4446,N_4481);
nor U4738 (N_4738,N_4271,N_4411);
nor U4739 (N_4739,N_4249,N_4473);
and U4740 (N_4740,N_4191,N_4114);
nand U4741 (N_4741,N_4050,N_4410);
nor U4742 (N_4742,N_4268,N_4250);
nor U4743 (N_4743,N_4346,N_4394);
nand U4744 (N_4744,N_4392,N_4381);
and U4745 (N_4745,N_4443,N_4226);
nor U4746 (N_4746,N_4335,N_4306);
or U4747 (N_4747,N_4435,N_4079);
nor U4748 (N_4748,N_4371,N_4484);
and U4749 (N_4749,N_4299,N_4041);
nand U4750 (N_4750,N_4213,N_4393);
nand U4751 (N_4751,N_4357,N_4468);
and U4752 (N_4752,N_4349,N_4060);
and U4753 (N_4753,N_4299,N_4264);
and U4754 (N_4754,N_4248,N_4438);
nand U4755 (N_4755,N_4292,N_4238);
nor U4756 (N_4756,N_4343,N_4419);
nand U4757 (N_4757,N_4068,N_4082);
and U4758 (N_4758,N_4482,N_4017);
and U4759 (N_4759,N_4420,N_4332);
nand U4760 (N_4760,N_4496,N_4072);
nor U4761 (N_4761,N_4136,N_4180);
or U4762 (N_4762,N_4467,N_4248);
or U4763 (N_4763,N_4279,N_4465);
xor U4764 (N_4764,N_4117,N_4024);
nor U4765 (N_4765,N_4454,N_4084);
or U4766 (N_4766,N_4140,N_4374);
and U4767 (N_4767,N_4367,N_4150);
and U4768 (N_4768,N_4123,N_4367);
nor U4769 (N_4769,N_4345,N_4346);
or U4770 (N_4770,N_4030,N_4183);
nor U4771 (N_4771,N_4440,N_4248);
nor U4772 (N_4772,N_4496,N_4297);
nand U4773 (N_4773,N_4479,N_4463);
nor U4774 (N_4774,N_4168,N_4281);
and U4775 (N_4775,N_4317,N_4233);
or U4776 (N_4776,N_4346,N_4108);
or U4777 (N_4777,N_4185,N_4456);
and U4778 (N_4778,N_4144,N_4414);
nor U4779 (N_4779,N_4024,N_4139);
or U4780 (N_4780,N_4132,N_4269);
and U4781 (N_4781,N_4283,N_4149);
nand U4782 (N_4782,N_4383,N_4246);
nor U4783 (N_4783,N_4214,N_4006);
nand U4784 (N_4784,N_4494,N_4053);
and U4785 (N_4785,N_4101,N_4227);
nand U4786 (N_4786,N_4034,N_4299);
or U4787 (N_4787,N_4394,N_4242);
and U4788 (N_4788,N_4145,N_4028);
and U4789 (N_4789,N_4381,N_4345);
and U4790 (N_4790,N_4248,N_4245);
nand U4791 (N_4791,N_4361,N_4325);
or U4792 (N_4792,N_4330,N_4100);
or U4793 (N_4793,N_4116,N_4492);
and U4794 (N_4794,N_4234,N_4405);
nand U4795 (N_4795,N_4330,N_4192);
nand U4796 (N_4796,N_4422,N_4412);
nor U4797 (N_4797,N_4273,N_4153);
or U4798 (N_4798,N_4409,N_4252);
nor U4799 (N_4799,N_4192,N_4017);
nor U4800 (N_4800,N_4261,N_4284);
or U4801 (N_4801,N_4327,N_4421);
and U4802 (N_4802,N_4293,N_4454);
nand U4803 (N_4803,N_4066,N_4082);
and U4804 (N_4804,N_4187,N_4485);
nand U4805 (N_4805,N_4203,N_4487);
nor U4806 (N_4806,N_4228,N_4439);
nor U4807 (N_4807,N_4349,N_4008);
nor U4808 (N_4808,N_4223,N_4458);
nor U4809 (N_4809,N_4272,N_4248);
nor U4810 (N_4810,N_4414,N_4482);
nor U4811 (N_4811,N_4024,N_4044);
and U4812 (N_4812,N_4091,N_4382);
nor U4813 (N_4813,N_4230,N_4204);
nor U4814 (N_4814,N_4342,N_4281);
and U4815 (N_4815,N_4391,N_4203);
or U4816 (N_4816,N_4202,N_4001);
nor U4817 (N_4817,N_4459,N_4102);
or U4818 (N_4818,N_4020,N_4081);
or U4819 (N_4819,N_4397,N_4118);
and U4820 (N_4820,N_4229,N_4271);
or U4821 (N_4821,N_4222,N_4177);
nor U4822 (N_4822,N_4458,N_4076);
nor U4823 (N_4823,N_4189,N_4299);
nor U4824 (N_4824,N_4330,N_4019);
and U4825 (N_4825,N_4326,N_4188);
and U4826 (N_4826,N_4353,N_4004);
and U4827 (N_4827,N_4411,N_4204);
nor U4828 (N_4828,N_4466,N_4481);
nor U4829 (N_4829,N_4037,N_4092);
and U4830 (N_4830,N_4192,N_4402);
nand U4831 (N_4831,N_4221,N_4011);
nor U4832 (N_4832,N_4061,N_4441);
or U4833 (N_4833,N_4160,N_4398);
nor U4834 (N_4834,N_4152,N_4185);
or U4835 (N_4835,N_4254,N_4112);
nand U4836 (N_4836,N_4111,N_4186);
or U4837 (N_4837,N_4254,N_4423);
nor U4838 (N_4838,N_4077,N_4488);
or U4839 (N_4839,N_4455,N_4014);
and U4840 (N_4840,N_4302,N_4417);
nor U4841 (N_4841,N_4275,N_4416);
nor U4842 (N_4842,N_4474,N_4084);
or U4843 (N_4843,N_4375,N_4138);
and U4844 (N_4844,N_4428,N_4167);
and U4845 (N_4845,N_4195,N_4419);
and U4846 (N_4846,N_4087,N_4031);
nand U4847 (N_4847,N_4072,N_4036);
and U4848 (N_4848,N_4416,N_4367);
and U4849 (N_4849,N_4034,N_4332);
or U4850 (N_4850,N_4092,N_4036);
and U4851 (N_4851,N_4321,N_4204);
nor U4852 (N_4852,N_4283,N_4393);
nand U4853 (N_4853,N_4460,N_4220);
nand U4854 (N_4854,N_4439,N_4145);
and U4855 (N_4855,N_4179,N_4474);
nand U4856 (N_4856,N_4216,N_4304);
nor U4857 (N_4857,N_4012,N_4008);
nand U4858 (N_4858,N_4018,N_4143);
nor U4859 (N_4859,N_4275,N_4457);
or U4860 (N_4860,N_4497,N_4050);
and U4861 (N_4861,N_4135,N_4378);
or U4862 (N_4862,N_4402,N_4138);
and U4863 (N_4863,N_4094,N_4419);
or U4864 (N_4864,N_4228,N_4404);
and U4865 (N_4865,N_4008,N_4297);
or U4866 (N_4866,N_4378,N_4196);
or U4867 (N_4867,N_4007,N_4054);
and U4868 (N_4868,N_4327,N_4331);
nor U4869 (N_4869,N_4327,N_4450);
nor U4870 (N_4870,N_4465,N_4067);
nor U4871 (N_4871,N_4035,N_4384);
and U4872 (N_4872,N_4198,N_4008);
or U4873 (N_4873,N_4286,N_4189);
or U4874 (N_4874,N_4237,N_4053);
and U4875 (N_4875,N_4033,N_4271);
or U4876 (N_4876,N_4443,N_4417);
nor U4877 (N_4877,N_4207,N_4164);
or U4878 (N_4878,N_4280,N_4470);
or U4879 (N_4879,N_4285,N_4094);
nand U4880 (N_4880,N_4263,N_4157);
or U4881 (N_4881,N_4322,N_4393);
and U4882 (N_4882,N_4300,N_4190);
nand U4883 (N_4883,N_4179,N_4283);
nand U4884 (N_4884,N_4362,N_4159);
nand U4885 (N_4885,N_4284,N_4134);
nand U4886 (N_4886,N_4231,N_4310);
nor U4887 (N_4887,N_4282,N_4052);
nand U4888 (N_4888,N_4427,N_4376);
or U4889 (N_4889,N_4456,N_4086);
or U4890 (N_4890,N_4206,N_4356);
nor U4891 (N_4891,N_4055,N_4240);
nand U4892 (N_4892,N_4065,N_4030);
and U4893 (N_4893,N_4456,N_4429);
or U4894 (N_4894,N_4498,N_4277);
or U4895 (N_4895,N_4287,N_4126);
nor U4896 (N_4896,N_4135,N_4105);
or U4897 (N_4897,N_4124,N_4004);
nor U4898 (N_4898,N_4395,N_4407);
nor U4899 (N_4899,N_4318,N_4137);
nor U4900 (N_4900,N_4130,N_4354);
or U4901 (N_4901,N_4283,N_4203);
nand U4902 (N_4902,N_4304,N_4492);
or U4903 (N_4903,N_4187,N_4025);
nand U4904 (N_4904,N_4055,N_4237);
and U4905 (N_4905,N_4213,N_4361);
nand U4906 (N_4906,N_4295,N_4249);
and U4907 (N_4907,N_4133,N_4382);
nor U4908 (N_4908,N_4394,N_4000);
and U4909 (N_4909,N_4097,N_4323);
or U4910 (N_4910,N_4051,N_4338);
and U4911 (N_4911,N_4389,N_4032);
and U4912 (N_4912,N_4258,N_4205);
or U4913 (N_4913,N_4484,N_4475);
or U4914 (N_4914,N_4384,N_4430);
or U4915 (N_4915,N_4021,N_4388);
or U4916 (N_4916,N_4350,N_4030);
nand U4917 (N_4917,N_4043,N_4068);
and U4918 (N_4918,N_4255,N_4440);
nor U4919 (N_4919,N_4122,N_4282);
or U4920 (N_4920,N_4099,N_4107);
nor U4921 (N_4921,N_4338,N_4116);
nor U4922 (N_4922,N_4255,N_4290);
and U4923 (N_4923,N_4270,N_4104);
nor U4924 (N_4924,N_4399,N_4274);
nor U4925 (N_4925,N_4337,N_4351);
and U4926 (N_4926,N_4348,N_4285);
or U4927 (N_4927,N_4403,N_4283);
nor U4928 (N_4928,N_4022,N_4026);
nand U4929 (N_4929,N_4132,N_4379);
nand U4930 (N_4930,N_4452,N_4069);
nand U4931 (N_4931,N_4172,N_4040);
nand U4932 (N_4932,N_4439,N_4411);
or U4933 (N_4933,N_4168,N_4154);
or U4934 (N_4934,N_4370,N_4287);
nand U4935 (N_4935,N_4003,N_4039);
xor U4936 (N_4936,N_4489,N_4323);
or U4937 (N_4937,N_4371,N_4232);
nand U4938 (N_4938,N_4106,N_4356);
and U4939 (N_4939,N_4113,N_4306);
nor U4940 (N_4940,N_4456,N_4065);
nor U4941 (N_4941,N_4375,N_4446);
nor U4942 (N_4942,N_4417,N_4160);
nand U4943 (N_4943,N_4378,N_4455);
nand U4944 (N_4944,N_4385,N_4063);
and U4945 (N_4945,N_4213,N_4387);
and U4946 (N_4946,N_4031,N_4188);
and U4947 (N_4947,N_4293,N_4219);
or U4948 (N_4948,N_4465,N_4369);
nor U4949 (N_4949,N_4463,N_4115);
or U4950 (N_4950,N_4451,N_4183);
nand U4951 (N_4951,N_4115,N_4425);
and U4952 (N_4952,N_4305,N_4323);
xor U4953 (N_4953,N_4483,N_4204);
nand U4954 (N_4954,N_4215,N_4094);
and U4955 (N_4955,N_4005,N_4291);
or U4956 (N_4956,N_4483,N_4065);
or U4957 (N_4957,N_4486,N_4458);
or U4958 (N_4958,N_4368,N_4460);
nand U4959 (N_4959,N_4129,N_4309);
and U4960 (N_4960,N_4184,N_4114);
nor U4961 (N_4961,N_4389,N_4136);
nor U4962 (N_4962,N_4417,N_4128);
nor U4963 (N_4963,N_4007,N_4468);
nand U4964 (N_4964,N_4279,N_4266);
nand U4965 (N_4965,N_4312,N_4437);
nor U4966 (N_4966,N_4487,N_4239);
and U4967 (N_4967,N_4410,N_4317);
and U4968 (N_4968,N_4101,N_4357);
or U4969 (N_4969,N_4428,N_4272);
and U4970 (N_4970,N_4049,N_4485);
nand U4971 (N_4971,N_4489,N_4069);
nor U4972 (N_4972,N_4293,N_4077);
or U4973 (N_4973,N_4139,N_4489);
nand U4974 (N_4974,N_4436,N_4463);
nor U4975 (N_4975,N_4276,N_4369);
and U4976 (N_4976,N_4048,N_4015);
nand U4977 (N_4977,N_4284,N_4098);
nor U4978 (N_4978,N_4217,N_4431);
nor U4979 (N_4979,N_4097,N_4186);
nor U4980 (N_4980,N_4293,N_4493);
and U4981 (N_4981,N_4071,N_4317);
nor U4982 (N_4982,N_4032,N_4123);
nor U4983 (N_4983,N_4162,N_4292);
and U4984 (N_4984,N_4070,N_4033);
and U4985 (N_4985,N_4303,N_4357);
nor U4986 (N_4986,N_4043,N_4216);
nor U4987 (N_4987,N_4102,N_4161);
and U4988 (N_4988,N_4441,N_4460);
nor U4989 (N_4989,N_4109,N_4016);
nand U4990 (N_4990,N_4060,N_4436);
and U4991 (N_4991,N_4199,N_4224);
nand U4992 (N_4992,N_4463,N_4226);
or U4993 (N_4993,N_4462,N_4488);
nand U4994 (N_4994,N_4043,N_4137);
nand U4995 (N_4995,N_4103,N_4268);
or U4996 (N_4996,N_4437,N_4191);
and U4997 (N_4997,N_4448,N_4262);
nor U4998 (N_4998,N_4167,N_4340);
nand U4999 (N_4999,N_4477,N_4253);
and UO_0 (O_0,N_4868,N_4627);
nand UO_1 (O_1,N_4935,N_4521);
and UO_2 (O_2,N_4602,N_4604);
nor UO_3 (O_3,N_4708,N_4832);
and UO_4 (O_4,N_4502,N_4750);
or UO_5 (O_5,N_4505,N_4683);
and UO_6 (O_6,N_4624,N_4967);
nand UO_7 (O_7,N_4993,N_4518);
nor UO_8 (O_8,N_4830,N_4836);
and UO_9 (O_9,N_4648,N_4882);
and UO_10 (O_10,N_4654,N_4721);
nor UO_11 (O_11,N_4735,N_4684);
or UO_12 (O_12,N_4664,N_4906);
nand UO_13 (O_13,N_4810,N_4558);
nand UO_14 (O_14,N_4957,N_4831);
and UO_15 (O_15,N_4710,N_4771);
nor UO_16 (O_16,N_4519,N_4788);
nand UO_17 (O_17,N_4525,N_4951);
nor UO_18 (O_18,N_4839,N_4621);
nor UO_19 (O_19,N_4887,N_4506);
nor UO_20 (O_20,N_4755,N_4989);
or UO_21 (O_21,N_4612,N_4799);
or UO_22 (O_22,N_4819,N_4659);
nand UO_23 (O_23,N_4855,N_4509);
and UO_24 (O_24,N_4939,N_4741);
xor UO_25 (O_25,N_4965,N_4784);
nand UO_26 (O_26,N_4572,N_4707);
or UO_27 (O_27,N_4941,N_4813);
nor UO_28 (O_28,N_4926,N_4875);
and UO_29 (O_29,N_4542,N_4745);
nor UO_30 (O_30,N_4733,N_4879);
nor UO_31 (O_31,N_4652,N_4711);
nor UO_32 (O_32,N_4559,N_4662);
nand UO_33 (O_33,N_4988,N_4686);
nor UO_34 (O_34,N_4985,N_4562);
and UO_35 (O_35,N_4590,N_4553);
and UO_36 (O_36,N_4829,N_4962);
nor UO_37 (O_37,N_4774,N_4514);
and UO_38 (O_38,N_4673,N_4880);
and UO_39 (O_39,N_4675,N_4805);
nand UO_40 (O_40,N_4874,N_4797);
and UO_41 (O_41,N_4751,N_4640);
and UO_42 (O_42,N_4690,N_4615);
nand UO_43 (O_43,N_4959,N_4762);
and UO_44 (O_44,N_4802,N_4894);
nand UO_45 (O_45,N_4948,N_4807);
nand UO_46 (O_46,N_4945,N_4703);
nand UO_47 (O_47,N_4983,N_4942);
or UO_48 (O_48,N_4950,N_4680);
or UO_49 (O_49,N_4717,N_4936);
and UO_50 (O_50,N_4638,N_4793);
and UO_51 (O_51,N_4619,N_4757);
nor UO_52 (O_52,N_4840,N_4593);
nand UO_53 (O_53,N_4713,N_4731);
or UO_54 (O_54,N_4556,N_4865);
or UO_55 (O_55,N_4920,N_4599);
nor UO_56 (O_56,N_4584,N_4543);
nand UO_57 (O_57,N_4603,N_4552);
nand UO_58 (O_58,N_4607,N_4586);
nand UO_59 (O_59,N_4977,N_4761);
or UO_60 (O_60,N_4528,N_4620);
nor UO_61 (O_61,N_4611,N_4642);
nand UO_62 (O_62,N_4958,N_4651);
nand UO_63 (O_63,N_4925,N_4682);
and UO_64 (O_64,N_4693,N_4606);
or UO_65 (O_65,N_4854,N_4554);
or UO_66 (O_66,N_4698,N_4576);
or UO_67 (O_67,N_4695,N_4567);
nand UO_68 (O_68,N_4522,N_4823);
or UO_69 (O_69,N_4706,N_4971);
nor UO_70 (O_70,N_4808,N_4669);
and UO_71 (O_71,N_4623,N_4534);
nor UO_72 (O_72,N_4952,N_4895);
or UO_73 (O_73,N_4786,N_4866);
nand UO_74 (O_74,N_4881,N_4550);
or UO_75 (O_75,N_4591,N_4500);
or UO_76 (O_76,N_4828,N_4595);
nand UO_77 (O_77,N_4845,N_4859);
or UO_78 (O_78,N_4949,N_4561);
or UO_79 (O_79,N_4566,N_4943);
nor UO_80 (O_80,N_4577,N_4626);
or UO_81 (O_81,N_4650,N_4516);
nand UO_82 (O_82,N_4876,N_4955);
or UO_83 (O_83,N_4582,N_4512);
and UO_84 (O_84,N_4665,N_4589);
nor UO_85 (O_85,N_4547,N_4800);
nand UO_86 (O_86,N_4990,N_4563);
nand UO_87 (O_87,N_4764,N_4700);
or UO_88 (O_88,N_4885,N_4724);
nor UO_89 (O_89,N_4523,N_4631);
or UO_90 (O_90,N_4794,N_4574);
or UO_91 (O_91,N_4656,N_4646);
and UO_92 (O_92,N_4816,N_4727);
nand UO_93 (O_93,N_4934,N_4918);
nand UO_94 (O_94,N_4692,N_4780);
and UO_95 (O_95,N_4746,N_4548);
nand UO_96 (O_96,N_4744,N_4928);
nor UO_97 (O_97,N_4919,N_4610);
nor UO_98 (O_98,N_4573,N_4995);
and UO_99 (O_99,N_4791,N_4981);
nor UO_100 (O_100,N_4898,N_4689);
or UO_101 (O_101,N_4725,N_4817);
nand UO_102 (O_102,N_4888,N_4782);
or UO_103 (O_103,N_4601,N_4598);
nand UO_104 (O_104,N_4777,N_4637);
nor UO_105 (O_105,N_4860,N_4511);
or UO_106 (O_106,N_4583,N_4766);
nor UO_107 (O_107,N_4527,N_4768);
nand UO_108 (O_108,N_4825,N_4685);
and UO_109 (O_109,N_4886,N_4809);
and UO_110 (O_110,N_4901,N_4778);
nor UO_111 (O_111,N_4975,N_4565);
xor UO_112 (O_112,N_4931,N_4676);
and UO_113 (O_113,N_4767,N_4740);
and UO_114 (O_114,N_4564,N_4785);
or UO_115 (O_115,N_4663,N_4980);
nand UO_116 (O_116,N_4944,N_4504);
nand UO_117 (O_117,N_4629,N_4917);
or UO_118 (O_118,N_4691,N_4914);
or UO_119 (O_119,N_4847,N_4739);
or UO_120 (O_120,N_4668,N_4862);
or UO_121 (O_121,N_4608,N_4963);
or UO_122 (O_122,N_4578,N_4570);
and UO_123 (O_123,N_4970,N_4661);
and UO_124 (O_124,N_4753,N_4770);
and UO_125 (O_125,N_4848,N_4940);
and UO_126 (O_126,N_4575,N_4537);
and UO_127 (O_127,N_4737,N_4699);
and UO_128 (O_128,N_4643,N_4723);
and UO_129 (O_129,N_4787,N_4776);
or UO_130 (O_130,N_4890,N_4987);
nor UO_131 (O_131,N_4658,N_4947);
nand UO_132 (O_132,N_4927,N_4670);
and UO_133 (O_133,N_4545,N_4969);
and UO_134 (O_134,N_4588,N_4858);
nand UO_135 (O_135,N_4672,N_4529);
or UO_136 (O_136,N_4709,N_4869);
nor UO_137 (O_137,N_4758,N_4933);
and UO_138 (O_138,N_4968,N_4540);
or UO_139 (O_139,N_4671,N_4846);
and UO_140 (O_140,N_4795,N_4736);
nand UO_141 (O_141,N_4551,N_4946);
nand UO_142 (O_142,N_4715,N_4634);
nand UO_143 (O_143,N_4982,N_4687);
and UO_144 (O_144,N_4870,N_4913);
and UO_145 (O_145,N_4956,N_4826);
or UO_146 (O_146,N_4597,N_4763);
and UO_147 (O_147,N_4580,N_4877);
or UO_148 (O_148,N_4806,N_4726);
and UO_149 (O_149,N_4867,N_4824);
or UO_150 (O_150,N_4961,N_4924);
or UO_151 (O_151,N_4533,N_4722);
nor UO_152 (O_152,N_4660,N_4732);
and UO_153 (O_153,N_4701,N_4520);
nor UO_154 (O_154,N_4748,N_4850);
nor UO_155 (O_155,N_4702,N_4738);
nor UO_156 (O_156,N_4605,N_4508);
nand UO_157 (O_157,N_4953,N_4716);
nand UO_158 (O_158,N_4842,N_4843);
nor UO_159 (O_159,N_4600,N_4835);
nor UO_160 (O_160,N_4635,N_4891);
nand UO_161 (O_161,N_4754,N_4636);
or UO_162 (O_162,N_4694,N_4530);
nand UO_163 (O_163,N_4954,N_4639);
nor UO_164 (O_164,N_4790,N_4697);
nand UO_165 (O_165,N_4932,N_4938);
nor UO_166 (O_166,N_4728,N_4861);
and UO_167 (O_167,N_4812,N_4811);
and UO_168 (O_168,N_4515,N_4789);
or UO_169 (O_169,N_4966,N_4999);
nor UO_170 (O_170,N_4674,N_4622);
or UO_171 (O_171,N_4837,N_4994);
and UO_172 (O_172,N_4613,N_4792);
nor UO_173 (O_173,N_4507,N_4517);
nand UO_174 (O_174,N_4546,N_4992);
nand UO_175 (O_175,N_4531,N_4900);
or UO_176 (O_176,N_4844,N_4827);
nand UO_177 (O_177,N_4743,N_4772);
and UO_178 (O_178,N_4922,N_4779);
nor UO_179 (O_179,N_4899,N_4625);
and UO_180 (O_180,N_4557,N_4781);
nand UO_181 (O_181,N_4617,N_4976);
nand UO_182 (O_182,N_4614,N_4814);
or UO_183 (O_183,N_4863,N_4657);
nor UO_184 (O_184,N_4719,N_4585);
nand UO_185 (O_185,N_4749,N_4532);
nand UO_186 (O_186,N_4747,N_4972);
or UO_187 (O_187,N_4857,N_4873);
nand UO_188 (O_188,N_4775,N_4524);
and UO_189 (O_189,N_4594,N_4718);
nor UO_190 (O_190,N_4923,N_4915);
nand UO_191 (O_191,N_4756,N_4804);
or UO_192 (O_192,N_4618,N_4632);
nand UO_193 (O_193,N_4596,N_4752);
or UO_194 (O_194,N_4641,N_4760);
or UO_195 (O_195,N_4503,N_4974);
nand UO_196 (O_196,N_4679,N_4921);
nand UO_197 (O_197,N_4730,N_4960);
or UO_198 (O_198,N_4526,N_4783);
nor UO_199 (O_199,N_4904,N_4910);
and UO_200 (O_200,N_4649,N_4849);
nand UO_201 (O_201,N_4609,N_4838);
nor UO_202 (O_202,N_4688,N_4883);
nand UO_203 (O_203,N_4677,N_4912);
or UO_204 (O_204,N_4705,N_4630);
and UO_205 (O_205,N_4538,N_4964);
or UO_206 (O_206,N_4905,N_4571);
and UO_207 (O_207,N_4513,N_4852);
nor UO_208 (O_208,N_4544,N_4916);
nor UO_209 (O_209,N_4773,N_4893);
nor UO_210 (O_210,N_4841,N_4569);
or UO_211 (O_211,N_4796,N_4579);
xnor UO_212 (O_212,N_4896,N_4549);
and UO_213 (O_213,N_4729,N_4510);
nor UO_214 (O_214,N_4555,N_4889);
or UO_215 (O_215,N_4984,N_4678);
nand UO_216 (O_216,N_4734,N_4929);
nand UO_217 (O_217,N_4803,N_4653);
nand UO_218 (O_218,N_4986,N_4560);
nor UO_219 (O_219,N_4645,N_4535);
or UO_220 (O_220,N_4655,N_4878);
nor UO_221 (O_221,N_4979,N_4801);
nand UO_222 (O_222,N_4712,N_4798);
nor UO_223 (O_223,N_4667,N_4536);
nor UO_224 (O_224,N_4991,N_4908);
nand UO_225 (O_225,N_4834,N_4907);
nand UO_226 (O_226,N_4937,N_4903);
or UO_227 (O_227,N_4892,N_4996);
or UO_228 (O_228,N_4820,N_4853);
nand UO_229 (O_229,N_4714,N_4633);
and UO_230 (O_230,N_4997,N_4587);
and UO_231 (O_231,N_4851,N_4884);
or UO_232 (O_232,N_4902,N_4856);
and UO_233 (O_233,N_4765,N_4616);
nor UO_234 (O_234,N_4930,N_4973);
nand UO_235 (O_235,N_4720,N_4978);
and UO_236 (O_236,N_4818,N_4897);
and UO_237 (O_237,N_4833,N_4998);
or UO_238 (O_238,N_4592,N_4647);
and UO_239 (O_239,N_4872,N_4911);
nand UO_240 (O_240,N_4822,N_4815);
nand UO_241 (O_241,N_4628,N_4681);
and UO_242 (O_242,N_4501,N_4704);
nor UO_243 (O_243,N_4759,N_4909);
nand UO_244 (O_244,N_4769,N_4541);
and UO_245 (O_245,N_4821,N_4696);
and UO_246 (O_246,N_4581,N_4864);
xnor UO_247 (O_247,N_4539,N_4742);
nand UO_248 (O_248,N_4666,N_4871);
or UO_249 (O_249,N_4644,N_4568);
and UO_250 (O_250,N_4644,N_4646);
xnor UO_251 (O_251,N_4691,N_4594);
nand UO_252 (O_252,N_4550,N_4608);
nor UO_253 (O_253,N_4970,N_4967);
nor UO_254 (O_254,N_4936,N_4775);
nor UO_255 (O_255,N_4904,N_4728);
nand UO_256 (O_256,N_4524,N_4961);
nor UO_257 (O_257,N_4931,N_4576);
nand UO_258 (O_258,N_4696,N_4857);
and UO_259 (O_259,N_4603,N_4514);
nor UO_260 (O_260,N_4951,N_4852);
nand UO_261 (O_261,N_4716,N_4663);
and UO_262 (O_262,N_4565,N_4674);
nand UO_263 (O_263,N_4678,N_4880);
nand UO_264 (O_264,N_4849,N_4531);
nor UO_265 (O_265,N_4655,N_4841);
nor UO_266 (O_266,N_4733,N_4947);
or UO_267 (O_267,N_4558,N_4685);
or UO_268 (O_268,N_4857,N_4894);
or UO_269 (O_269,N_4856,N_4819);
and UO_270 (O_270,N_4955,N_4866);
nand UO_271 (O_271,N_4824,N_4724);
nor UO_272 (O_272,N_4530,N_4522);
nor UO_273 (O_273,N_4684,N_4976);
nand UO_274 (O_274,N_4641,N_4549);
nand UO_275 (O_275,N_4700,N_4849);
and UO_276 (O_276,N_4623,N_4573);
or UO_277 (O_277,N_4964,N_4935);
and UO_278 (O_278,N_4918,N_4774);
nand UO_279 (O_279,N_4581,N_4627);
and UO_280 (O_280,N_4820,N_4801);
nand UO_281 (O_281,N_4542,N_4512);
nand UO_282 (O_282,N_4645,N_4883);
nor UO_283 (O_283,N_4892,N_4679);
and UO_284 (O_284,N_4666,N_4841);
nand UO_285 (O_285,N_4888,N_4968);
or UO_286 (O_286,N_4713,N_4725);
nor UO_287 (O_287,N_4504,N_4917);
nor UO_288 (O_288,N_4848,N_4801);
or UO_289 (O_289,N_4995,N_4552);
or UO_290 (O_290,N_4754,N_4874);
nand UO_291 (O_291,N_4915,N_4801);
nand UO_292 (O_292,N_4976,N_4963);
nand UO_293 (O_293,N_4941,N_4518);
nand UO_294 (O_294,N_4698,N_4646);
and UO_295 (O_295,N_4994,N_4864);
and UO_296 (O_296,N_4608,N_4630);
nand UO_297 (O_297,N_4662,N_4891);
or UO_298 (O_298,N_4504,N_4523);
or UO_299 (O_299,N_4702,N_4913);
or UO_300 (O_300,N_4603,N_4763);
nor UO_301 (O_301,N_4603,N_4973);
nand UO_302 (O_302,N_4778,N_4683);
and UO_303 (O_303,N_4579,N_4697);
or UO_304 (O_304,N_4552,N_4926);
nor UO_305 (O_305,N_4880,N_4774);
nor UO_306 (O_306,N_4962,N_4500);
or UO_307 (O_307,N_4859,N_4713);
nor UO_308 (O_308,N_4805,N_4519);
nor UO_309 (O_309,N_4772,N_4708);
or UO_310 (O_310,N_4864,N_4735);
nand UO_311 (O_311,N_4738,N_4981);
nor UO_312 (O_312,N_4908,N_4712);
nand UO_313 (O_313,N_4575,N_4751);
or UO_314 (O_314,N_4815,N_4921);
or UO_315 (O_315,N_4615,N_4649);
nor UO_316 (O_316,N_4523,N_4990);
and UO_317 (O_317,N_4502,N_4854);
nor UO_318 (O_318,N_4914,N_4606);
or UO_319 (O_319,N_4796,N_4790);
nand UO_320 (O_320,N_4681,N_4535);
or UO_321 (O_321,N_4561,N_4614);
nand UO_322 (O_322,N_4906,N_4985);
nand UO_323 (O_323,N_4644,N_4924);
and UO_324 (O_324,N_4859,N_4925);
and UO_325 (O_325,N_4574,N_4617);
and UO_326 (O_326,N_4803,N_4536);
nand UO_327 (O_327,N_4507,N_4780);
nor UO_328 (O_328,N_4593,N_4819);
nor UO_329 (O_329,N_4690,N_4932);
xnor UO_330 (O_330,N_4717,N_4537);
and UO_331 (O_331,N_4748,N_4896);
nor UO_332 (O_332,N_4731,N_4512);
or UO_333 (O_333,N_4972,N_4687);
and UO_334 (O_334,N_4895,N_4625);
and UO_335 (O_335,N_4892,N_4854);
nor UO_336 (O_336,N_4934,N_4899);
nand UO_337 (O_337,N_4598,N_4500);
or UO_338 (O_338,N_4706,N_4778);
and UO_339 (O_339,N_4674,N_4606);
nor UO_340 (O_340,N_4838,N_4572);
nor UO_341 (O_341,N_4617,N_4950);
nor UO_342 (O_342,N_4567,N_4795);
or UO_343 (O_343,N_4646,N_4760);
and UO_344 (O_344,N_4938,N_4862);
nor UO_345 (O_345,N_4517,N_4976);
nand UO_346 (O_346,N_4605,N_4708);
nor UO_347 (O_347,N_4595,N_4991);
and UO_348 (O_348,N_4828,N_4616);
or UO_349 (O_349,N_4778,N_4676);
nand UO_350 (O_350,N_4912,N_4932);
and UO_351 (O_351,N_4696,N_4732);
and UO_352 (O_352,N_4545,N_4908);
xnor UO_353 (O_353,N_4644,N_4507);
and UO_354 (O_354,N_4800,N_4519);
and UO_355 (O_355,N_4937,N_4546);
nand UO_356 (O_356,N_4940,N_4941);
nand UO_357 (O_357,N_4737,N_4515);
or UO_358 (O_358,N_4780,N_4785);
and UO_359 (O_359,N_4787,N_4638);
or UO_360 (O_360,N_4537,N_4668);
and UO_361 (O_361,N_4528,N_4974);
or UO_362 (O_362,N_4857,N_4921);
and UO_363 (O_363,N_4646,N_4692);
nor UO_364 (O_364,N_4633,N_4549);
or UO_365 (O_365,N_4855,N_4945);
or UO_366 (O_366,N_4623,N_4935);
xnor UO_367 (O_367,N_4798,N_4583);
nand UO_368 (O_368,N_4557,N_4690);
and UO_369 (O_369,N_4597,N_4835);
or UO_370 (O_370,N_4979,N_4681);
and UO_371 (O_371,N_4660,N_4639);
nor UO_372 (O_372,N_4546,N_4586);
and UO_373 (O_373,N_4956,N_4615);
nand UO_374 (O_374,N_4952,N_4613);
xor UO_375 (O_375,N_4677,N_4883);
and UO_376 (O_376,N_4589,N_4906);
nand UO_377 (O_377,N_4959,N_4807);
or UO_378 (O_378,N_4552,N_4978);
or UO_379 (O_379,N_4712,N_4819);
and UO_380 (O_380,N_4994,N_4936);
and UO_381 (O_381,N_4908,N_4828);
and UO_382 (O_382,N_4732,N_4993);
and UO_383 (O_383,N_4889,N_4780);
nor UO_384 (O_384,N_4938,N_4709);
nand UO_385 (O_385,N_4704,N_4982);
nand UO_386 (O_386,N_4985,N_4679);
and UO_387 (O_387,N_4963,N_4732);
and UO_388 (O_388,N_4568,N_4738);
nor UO_389 (O_389,N_4833,N_4793);
or UO_390 (O_390,N_4693,N_4949);
and UO_391 (O_391,N_4697,N_4857);
nor UO_392 (O_392,N_4991,N_4593);
and UO_393 (O_393,N_4660,N_4640);
and UO_394 (O_394,N_4758,N_4972);
and UO_395 (O_395,N_4504,N_4612);
nand UO_396 (O_396,N_4635,N_4934);
or UO_397 (O_397,N_4862,N_4673);
nor UO_398 (O_398,N_4930,N_4929);
and UO_399 (O_399,N_4625,N_4612);
or UO_400 (O_400,N_4687,N_4748);
nand UO_401 (O_401,N_4750,N_4696);
and UO_402 (O_402,N_4781,N_4640);
nand UO_403 (O_403,N_4635,N_4940);
and UO_404 (O_404,N_4556,N_4676);
nor UO_405 (O_405,N_4960,N_4966);
nor UO_406 (O_406,N_4670,N_4544);
and UO_407 (O_407,N_4664,N_4985);
or UO_408 (O_408,N_4753,N_4747);
and UO_409 (O_409,N_4952,N_4810);
and UO_410 (O_410,N_4875,N_4541);
and UO_411 (O_411,N_4578,N_4560);
or UO_412 (O_412,N_4922,N_4896);
and UO_413 (O_413,N_4800,N_4744);
and UO_414 (O_414,N_4639,N_4738);
or UO_415 (O_415,N_4571,N_4710);
nand UO_416 (O_416,N_4741,N_4959);
nand UO_417 (O_417,N_4793,N_4697);
nor UO_418 (O_418,N_4708,N_4854);
nand UO_419 (O_419,N_4966,N_4673);
and UO_420 (O_420,N_4786,N_4776);
nor UO_421 (O_421,N_4986,N_4987);
nor UO_422 (O_422,N_4624,N_4770);
nand UO_423 (O_423,N_4809,N_4567);
and UO_424 (O_424,N_4756,N_4805);
nor UO_425 (O_425,N_4740,N_4874);
nor UO_426 (O_426,N_4905,N_4867);
nor UO_427 (O_427,N_4717,N_4771);
and UO_428 (O_428,N_4691,N_4835);
and UO_429 (O_429,N_4614,N_4693);
or UO_430 (O_430,N_4950,N_4830);
or UO_431 (O_431,N_4595,N_4809);
nor UO_432 (O_432,N_4702,N_4699);
or UO_433 (O_433,N_4986,N_4925);
or UO_434 (O_434,N_4912,N_4606);
nand UO_435 (O_435,N_4906,N_4768);
or UO_436 (O_436,N_4908,N_4803);
and UO_437 (O_437,N_4758,N_4660);
nor UO_438 (O_438,N_4971,N_4690);
or UO_439 (O_439,N_4642,N_4878);
nor UO_440 (O_440,N_4792,N_4577);
nand UO_441 (O_441,N_4884,N_4794);
nor UO_442 (O_442,N_4551,N_4672);
nand UO_443 (O_443,N_4731,N_4808);
nor UO_444 (O_444,N_4989,N_4879);
and UO_445 (O_445,N_4648,N_4998);
and UO_446 (O_446,N_4613,N_4750);
nor UO_447 (O_447,N_4960,N_4946);
or UO_448 (O_448,N_4724,N_4608);
nand UO_449 (O_449,N_4692,N_4898);
nand UO_450 (O_450,N_4991,N_4936);
nand UO_451 (O_451,N_4894,N_4916);
or UO_452 (O_452,N_4789,N_4685);
nand UO_453 (O_453,N_4935,N_4527);
or UO_454 (O_454,N_4524,N_4620);
or UO_455 (O_455,N_4709,N_4578);
nand UO_456 (O_456,N_4946,N_4937);
and UO_457 (O_457,N_4672,N_4710);
or UO_458 (O_458,N_4572,N_4524);
nand UO_459 (O_459,N_4675,N_4901);
nand UO_460 (O_460,N_4742,N_4875);
nor UO_461 (O_461,N_4715,N_4547);
nand UO_462 (O_462,N_4888,N_4923);
or UO_463 (O_463,N_4637,N_4645);
nand UO_464 (O_464,N_4622,N_4512);
and UO_465 (O_465,N_4718,N_4696);
nand UO_466 (O_466,N_4635,N_4501);
and UO_467 (O_467,N_4581,N_4899);
nand UO_468 (O_468,N_4714,N_4760);
xor UO_469 (O_469,N_4624,N_4754);
nand UO_470 (O_470,N_4983,N_4566);
and UO_471 (O_471,N_4721,N_4507);
nand UO_472 (O_472,N_4531,N_4693);
and UO_473 (O_473,N_4780,N_4972);
or UO_474 (O_474,N_4880,N_4995);
or UO_475 (O_475,N_4608,N_4775);
and UO_476 (O_476,N_4721,N_4697);
or UO_477 (O_477,N_4577,N_4604);
nor UO_478 (O_478,N_4946,N_4710);
nand UO_479 (O_479,N_4691,N_4894);
or UO_480 (O_480,N_4954,N_4853);
and UO_481 (O_481,N_4589,N_4986);
and UO_482 (O_482,N_4659,N_4609);
nand UO_483 (O_483,N_4698,N_4571);
or UO_484 (O_484,N_4571,N_4520);
nand UO_485 (O_485,N_4636,N_4891);
xnor UO_486 (O_486,N_4697,N_4561);
or UO_487 (O_487,N_4826,N_4570);
and UO_488 (O_488,N_4547,N_4886);
and UO_489 (O_489,N_4977,N_4674);
and UO_490 (O_490,N_4544,N_4527);
or UO_491 (O_491,N_4826,N_4711);
or UO_492 (O_492,N_4942,N_4501);
nor UO_493 (O_493,N_4620,N_4535);
and UO_494 (O_494,N_4675,N_4783);
nand UO_495 (O_495,N_4995,N_4825);
nor UO_496 (O_496,N_4592,N_4842);
nand UO_497 (O_497,N_4708,N_4697);
or UO_498 (O_498,N_4633,N_4891);
nand UO_499 (O_499,N_4793,N_4799);
nand UO_500 (O_500,N_4944,N_4926);
nor UO_501 (O_501,N_4552,N_4921);
nand UO_502 (O_502,N_4755,N_4974);
and UO_503 (O_503,N_4656,N_4544);
or UO_504 (O_504,N_4565,N_4633);
and UO_505 (O_505,N_4713,N_4917);
and UO_506 (O_506,N_4510,N_4711);
nand UO_507 (O_507,N_4500,N_4929);
and UO_508 (O_508,N_4813,N_4718);
nand UO_509 (O_509,N_4500,N_4680);
nor UO_510 (O_510,N_4712,N_4773);
nand UO_511 (O_511,N_4704,N_4794);
nor UO_512 (O_512,N_4602,N_4626);
or UO_513 (O_513,N_4665,N_4818);
nand UO_514 (O_514,N_4722,N_4518);
nand UO_515 (O_515,N_4851,N_4907);
or UO_516 (O_516,N_4738,N_4662);
and UO_517 (O_517,N_4908,N_4974);
nor UO_518 (O_518,N_4982,N_4842);
and UO_519 (O_519,N_4746,N_4807);
nor UO_520 (O_520,N_4867,N_4549);
nor UO_521 (O_521,N_4707,N_4716);
or UO_522 (O_522,N_4891,N_4834);
and UO_523 (O_523,N_4656,N_4748);
and UO_524 (O_524,N_4623,N_4739);
nand UO_525 (O_525,N_4506,N_4923);
nor UO_526 (O_526,N_4896,N_4516);
or UO_527 (O_527,N_4557,N_4792);
and UO_528 (O_528,N_4923,N_4503);
or UO_529 (O_529,N_4994,N_4922);
or UO_530 (O_530,N_4587,N_4900);
and UO_531 (O_531,N_4641,N_4934);
and UO_532 (O_532,N_4531,N_4605);
and UO_533 (O_533,N_4778,N_4691);
nor UO_534 (O_534,N_4638,N_4726);
nor UO_535 (O_535,N_4820,N_4510);
nor UO_536 (O_536,N_4866,N_4908);
nor UO_537 (O_537,N_4562,N_4998);
or UO_538 (O_538,N_4912,N_4985);
and UO_539 (O_539,N_4583,N_4717);
xnor UO_540 (O_540,N_4591,N_4897);
or UO_541 (O_541,N_4940,N_4750);
and UO_542 (O_542,N_4973,N_4710);
nor UO_543 (O_543,N_4536,N_4776);
nor UO_544 (O_544,N_4976,N_4941);
nor UO_545 (O_545,N_4922,N_4787);
xor UO_546 (O_546,N_4801,N_4923);
nor UO_547 (O_547,N_4545,N_4850);
or UO_548 (O_548,N_4863,N_4637);
nand UO_549 (O_549,N_4530,N_4897);
xnor UO_550 (O_550,N_4743,N_4976);
and UO_551 (O_551,N_4599,N_4602);
and UO_552 (O_552,N_4833,N_4613);
nor UO_553 (O_553,N_4819,N_4756);
nand UO_554 (O_554,N_4741,N_4962);
nand UO_555 (O_555,N_4732,N_4874);
nor UO_556 (O_556,N_4515,N_4658);
nor UO_557 (O_557,N_4636,N_4771);
nand UO_558 (O_558,N_4521,N_4813);
or UO_559 (O_559,N_4612,N_4871);
or UO_560 (O_560,N_4616,N_4854);
nand UO_561 (O_561,N_4964,N_4960);
nand UO_562 (O_562,N_4926,N_4550);
xor UO_563 (O_563,N_4540,N_4500);
nand UO_564 (O_564,N_4754,N_4873);
nor UO_565 (O_565,N_4681,N_4677);
or UO_566 (O_566,N_4952,N_4647);
nand UO_567 (O_567,N_4632,N_4981);
or UO_568 (O_568,N_4959,N_4743);
or UO_569 (O_569,N_4506,N_4636);
nand UO_570 (O_570,N_4966,N_4648);
nand UO_571 (O_571,N_4717,N_4670);
and UO_572 (O_572,N_4521,N_4724);
or UO_573 (O_573,N_4841,N_4825);
nor UO_574 (O_574,N_4647,N_4767);
nand UO_575 (O_575,N_4564,N_4580);
and UO_576 (O_576,N_4942,N_4696);
and UO_577 (O_577,N_4824,N_4728);
nor UO_578 (O_578,N_4772,N_4630);
nand UO_579 (O_579,N_4555,N_4904);
and UO_580 (O_580,N_4755,N_4754);
nor UO_581 (O_581,N_4851,N_4641);
and UO_582 (O_582,N_4728,N_4607);
nand UO_583 (O_583,N_4931,N_4967);
or UO_584 (O_584,N_4993,N_4994);
and UO_585 (O_585,N_4794,N_4579);
or UO_586 (O_586,N_4655,N_4865);
and UO_587 (O_587,N_4739,N_4795);
and UO_588 (O_588,N_4881,N_4689);
nor UO_589 (O_589,N_4747,N_4530);
or UO_590 (O_590,N_4605,N_4843);
and UO_591 (O_591,N_4814,N_4788);
nor UO_592 (O_592,N_4866,N_4627);
or UO_593 (O_593,N_4683,N_4944);
or UO_594 (O_594,N_4540,N_4790);
and UO_595 (O_595,N_4898,N_4876);
or UO_596 (O_596,N_4938,N_4634);
or UO_597 (O_597,N_4865,N_4792);
and UO_598 (O_598,N_4791,N_4952);
and UO_599 (O_599,N_4751,N_4658);
nor UO_600 (O_600,N_4558,N_4717);
nor UO_601 (O_601,N_4767,N_4721);
or UO_602 (O_602,N_4674,N_4612);
or UO_603 (O_603,N_4818,N_4706);
nor UO_604 (O_604,N_4550,N_4559);
nand UO_605 (O_605,N_4734,N_4509);
or UO_606 (O_606,N_4734,N_4695);
and UO_607 (O_607,N_4671,N_4998);
xnor UO_608 (O_608,N_4780,N_4648);
or UO_609 (O_609,N_4501,N_4695);
nor UO_610 (O_610,N_4563,N_4601);
nand UO_611 (O_611,N_4947,N_4565);
or UO_612 (O_612,N_4693,N_4539);
nor UO_613 (O_613,N_4867,N_4785);
nand UO_614 (O_614,N_4800,N_4581);
nand UO_615 (O_615,N_4603,N_4697);
or UO_616 (O_616,N_4563,N_4655);
nand UO_617 (O_617,N_4562,N_4921);
nor UO_618 (O_618,N_4823,N_4851);
nand UO_619 (O_619,N_4711,N_4722);
nor UO_620 (O_620,N_4958,N_4881);
or UO_621 (O_621,N_4965,N_4695);
or UO_622 (O_622,N_4580,N_4958);
nor UO_623 (O_623,N_4998,N_4997);
nor UO_624 (O_624,N_4989,N_4986);
or UO_625 (O_625,N_4624,N_4939);
nand UO_626 (O_626,N_4555,N_4982);
or UO_627 (O_627,N_4985,N_4601);
nand UO_628 (O_628,N_4853,N_4959);
and UO_629 (O_629,N_4503,N_4728);
nand UO_630 (O_630,N_4584,N_4526);
or UO_631 (O_631,N_4959,N_4808);
nor UO_632 (O_632,N_4726,N_4775);
and UO_633 (O_633,N_4705,N_4590);
nand UO_634 (O_634,N_4746,N_4841);
nor UO_635 (O_635,N_4742,N_4502);
nand UO_636 (O_636,N_4970,N_4575);
nand UO_637 (O_637,N_4979,N_4630);
and UO_638 (O_638,N_4709,N_4851);
or UO_639 (O_639,N_4809,N_4734);
or UO_640 (O_640,N_4501,N_4726);
and UO_641 (O_641,N_4743,N_4747);
nor UO_642 (O_642,N_4906,N_4629);
nor UO_643 (O_643,N_4864,N_4558);
and UO_644 (O_644,N_4511,N_4987);
and UO_645 (O_645,N_4767,N_4639);
or UO_646 (O_646,N_4873,N_4880);
nor UO_647 (O_647,N_4697,N_4774);
nor UO_648 (O_648,N_4551,N_4516);
and UO_649 (O_649,N_4801,N_4973);
nor UO_650 (O_650,N_4694,N_4732);
and UO_651 (O_651,N_4707,N_4883);
and UO_652 (O_652,N_4750,N_4682);
or UO_653 (O_653,N_4828,N_4625);
or UO_654 (O_654,N_4742,N_4931);
nor UO_655 (O_655,N_4518,N_4637);
nor UO_656 (O_656,N_4766,N_4579);
and UO_657 (O_657,N_4612,N_4993);
and UO_658 (O_658,N_4603,N_4851);
and UO_659 (O_659,N_4986,N_4882);
and UO_660 (O_660,N_4934,N_4862);
nand UO_661 (O_661,N_4704,N_4594);
nand UO_662 (O_662,N_4517,N_4860);
or UO_663 (O_663,N_4745,N_4806);
and UO_664 (O_664,N_4777,N_4743);
xnor UO_665 (O_665,N_4704,N_4900);
nor UO_666 (O_666,N_4543,N_4876);
and UO_667 (O_667,N_4813,N_4755);
nor UO_668 (O_668,N_4995,N_4801);
nand UO_669 (O_669,N_4940,N_4715);
nor UO_670 (O_670,N_4666,N_4693);
or UO_671 (O_671,N_4718,N_4814);
nand UO_672 (O_672,N_4793,N_4910);
or UO_673 (O_673,N_4902,N_4679);
and UO_674 (O_674,N_4963,N_4650);
and UO_675 (O_675,N_4765,N_4678);
nand UO_676 (O_676,N_4500,N_4607);
or UO_677 (O_677,N_4729,N_4711);
or UO_678 (O_678,N_4505,N_4752);
and UO_679 (O_679,N_4717,N_4847);
or UO_680 (O_680,N_4790,N_4907);
nor UO_681 (O_681,N_4502,N_4692);
nand UO_682 (O_682,N_4998,N_4735);
and UO_683 (O_683,N_4551,N_4923);
nor UO_684 (O_684,N_4722,N_4678);
nand UO_685 (O_685,N_4593,N_4984);
nand UO_686 (O_686,N_4578,N_4731);
nor UO_687 (O_687,N_4893,N_4953);
or UO_688 (O_688,N_4901,N_4978);
or UO_689 (O_689,N_4982,N_4843);
nor UO_690 (O_690,N_4679,N_4846);
and UO_691 (O_691,N_4948,N_4846);
nand UO_692 (O_692,N_4624,N_4896);
nand UO_693 (O_693,N_4738,N_4555);
or UO_694 (O_694,N_4780,N_4995);
nand UO_695 (O_695,N_4786,N_4676);
nand UO_696 (O_696,N_4636,N_4742);
nand UO_697 (O_697,N_4684,N_4886);
or UO_698 (O_698,N_4923,N_4897);
and UO_699 (O_699,N_4831,N_4749);
nor UO_700 (O_700,N_4960,N_4789);
nor UO_701 (O_701,N_4813,N_4612);
nand UO_702 (O_702,N_4782,N_4811);
or UO_703 (O_703,N_4768,N_4546);
or UO_704 (O_704,N_4883,N_4998);
or UO_705 (O_705,N_4832,N_4824);
nand UO_706 (O_706,N_4838,N_4869);
and UO_707 (O_707,N_4994,N_4971);
nand UO_708 (O_708,N_4813,N_4893);
nand UO_709 (O_709,N_4545,N_4844);
and UO_710 (O_710,N_4962,N_4783);
nor UO_711 (O_711,N_4810,N_4626);
or UO_712 (O_712,N_4548,N_4915);
and UO_713 (O_713,N_4565,N_4834);
or UO_714 (O_714,N_4850,N_4644);
or UO_715 (O_715,N_4731,N_4901);
nand UO_716 (O_716,N_4614,N_4878);
nor UO_717 (O_717,N_4953,N_4510);
and UO_718 (O_718,N_4717,N_4956);
and UO_719 (O_719,N_4640,N_4731);
or UO_720 (O_720,N_4861,N_4594);
nor UO_721 (O_721,N_4714,N_4712);
and UO_722 (O_722,N_4763,N_4970);
or UO_723 (O_723,N_4900,N_4625);
and UO_724 (O_724,N_4932,N_4999);
nor UO_725 (O_725,N_4562,N_4639);
nor UO_726 (O_726,N_4822,N_4817);
nor UO_727 (O_727,N_4665,N_4805);
nand UO_728 (O_728,N_4580,N_4894);
nor UO_729 (O_729,N_4706,N_4789);
nor UO_730 (O_730,N_4880,N_4912);
nand UO_731 (O_731,N_4828,N_4709);
nor UO_732 (O_732,N_4990,N_4861);
or UO_733 (O_733,N_4579,N_4590);
nand UO_734 (O_734,N_4909,N_4687);
nand UO_735 (O_735,N_4643,N_4744);
or UO_736 (O_736,N_4681,N_4867);
and UO_737 (O_737,N_4802,N_4763);
nand UO_738 (O_738,N_4811,N_4606);
and UO_739 (O_739,N_4553,N_4589);
and UO_740 (O_740,N_4510,N_4885);
and UO_741 (O_741,N_4639,N_4908);
nor UO_742 (O_742,N_4909,N_4815);
and UO_743 (O_743,N_4900,N_4567);
nand UO_744 (O_744,N_4865,N_4987);
or UO_745 (O_745,N_4913,N_4936);
nand UO_746 (O_746,N_4572,N_4876);
and UO_747 (O_747,N_4713,N_4912);
or UO_748 (O_748,N_4798,N_4969);
nand UO_749 (O_749,N_4508,N_4584);
nor UO_750 (O_750,N_4877,N_4645);
and UO_751 (O_751,N_4522,N_4694);
nand UO_752 (O_752,N_4637,N_4571);
or UO_753 (O_753,N_4884,N_4635);
nor UO_754 (O_754,N_4671,N_4994);
nor UO_755 (O_755,N_4840,N_4818);
nand UO_756 (O_756,N_4689,N_4563);
and UO_757 (O_757,N_4950,N_4555);
or UO_758 (O_758,N_4552,N_4608);
nand UO_759 (O_759,N_4801,N_4529);
and UO_760 (O_760,N_4923,N_4772);
and UO_761 (O_761,N_4674,N_4916);
nor UO_762 (O_762,N_4887,N_4663);
and UO_763 (O_763,N_4767,N_4916);
nor UO_764 (O_764,N_4928,N_4960);
nand UO_765 (O_765,N_4820,N_4836);
and UO_766 (O_766,N_4510,N_4781);
nor UO_767 (O_767,N_4991,N_4810);
nor UO_768 (O_768,N_4855,N_4902);
or UO_769 (O_769,N_4534,N_4605);
nor UO_770 (O_770,N_4937,N_4928);
nand UO_771 (O_771,N_4820,N_4810);
and UO_772 (O_772,N_4966,N_4521);
nor UO_773 (O_773,N_4802,N_4661);
nor UO_774 (O_774,N_4649,N_4509);
nand UO_775 (O_775,N_4510,N_4793);
or UO_776 (O_776,N_4627,N_4595);
nor UO_777 (O_777,N_4922,N_4950);
or UO_778 (O_778,N_4845,N_4936);
and UO_779 (O_779,N_4637,N_4952);
nor UO_780 (O_780,N_4676,N_4898);
nor UO_781 (O_781,N_4683,N_4659);
or UO_782 (O_782,N_4599,N_4590);
or UO_783 (O_783,N_4748,N_4852);
nor UO_784 (O_784,N_4530,N_4823);
and UO_785 (O_785,N_4540,N_4712);
nand UO_786 (O_786,N_4562,N_4529);
and UO_787 (O_787,N_4988,N_4790);
and UO_788 (O_788,N_4939,N_4869);
and UO_789 (O_789,N_4811,N_4947);
nor UO_790 (O_790,N_4842,N_4563);
and UO_791 (O_791,N_4540,N_4627);
and UO_792 (O_792,N_4759,N_4679);
and UO_793 (O_793,N_4734,N_4593);
and UO_794 (O_794,N_4933,N_4775);
and UO_795 (O_795,N_4584,N_4588);
nand UO_796 (O_796,N_4749,N_4842);
xnor UO_797 (O_797,N_4523,N_4627);
nor UO_798 (O_798,N_4523,N_4594);
nand UO_799 (O_799,N_4522,N_4620);
nor UO_800 (O_800,N_4907,N_4674);
nor UO_801 (O_801,N_4576,N_4619);
nor UO_802 (O_802,N_4606,N_4563);
and UO_803 (O_803,N_4858,N_4964);
nand UO_804 (O_804,N_4669,N_4660);
and UO_805 (O_805,N_4865,N_4940);
and UO_806 (O_806,N_4755,N_4923);
nor UO_807 (O_807,N_4844,N_4901);
nor UO_808 (O_808,N_4785,N_4737);
and UO_809 (O_809,N_4550,N_4675);
nand UO_810 (O_810,N_4661,N_4969);
xnor UO_811 (O_811,N_4651,N_4944);
and UO_812 (O_812,N_4798,N_4898);
nand UO_813 (O_813,N_4551,N_4829);
nand UO_814 (O_814,N_4886,N_4767);
and UO_815 (O_815,N_4975,N_4639);
or UO_816 (O_816,N_4700,N_4684);
and UO_817 (O_817,N_4644,N_4594);
nor UO_818 (O_818,N_4621,N_4755);
nand UO_819 (O_819,N_4679,N_4898);
nand UO_820 (O_820,N_4708,N_4882);
nor UO_821 (O_821,N_4796,N_4754);
nand UO_822 (O_822,N_4607,N_4881);
nor UO_823 (O_823,N_4897,N_4747);
nand UO_824 (O_824,N_4943,N_4533);
or UO_825 (O_825,N_4974,N_4894);
nand UO_826 (O_826,N_4508,N_4663);
or UO_827 (O_827,N_4640,N_4755);
and UO_828 (O_828,N_4716,N_4531);
and UO_829 (O_829,N_4928,N_4687);
and UO_830 (O_830,N_4523,N_4591);
or UO_831 (O_831,N_4666,N_4925);
and UO_832 (O_832,N_4853,N_4539);
nand UO_833 (O_833,N_4531,N_4940);
and UO_834 (O_834,N_4798,N_4811);
nor UO_835 (O_835,N_4728,N_4759);
or UO_836 (O_836,N_4931,N_4610);
nor UO_837 (O_837,N_4896,N_4635);
and UO_838 (O_838,N_4530,N_4920);
or UO_839 (O_839,N_4517,N_4651);
nor UO_840 (O_840,N_4829,N_4719);
nor UO_841 (O_841,N_4705,N_4681);
nand UO_842 (O_842,N_4706,N_4928);
or UO_843 (O_843,N_4990,N_4905);
nor UO_844 (O_844,N_4706,N_4745);
and UO_845 (O_845,N_4735,N_4872);
or UO_846 (O_846,N_4910,N_4852);
and UO_847 (O_847,N_4556,N_4554);
and UO_848 (O_848,N_4508,N_4745);
or UO_849 (O_849,N_4727,N_4923);
nand UO_850 (O_850,N_4984,N_4625);
or UO_851 (O_851,N_4580,N_4876);
or UO_852 (O_852,N_4886,N_4683);
or UO_853 (O_853,N_4723,N_4798);
or UO_854 (O_854,N_4977,N_4523);
nand UO_855 (O_855,N_4698,N_4810);
nor UO_856 (O_856,N_4891,N_4990);
nor UO_857 (O_857,N_4711,N_4599);
and UO_858 (O_858,N_4920,N_4554);
and UO_859 (O_859,N_4731,N_4542);
nor UO_860 (O_860,N_4885,N_4974);
nand UO_861 (O_861,N_4916,N_4877);
and UO_862 (O_862,N_4601,N_4862);
and UO_863 (O_863,N_4740,N_4967);
and UO_864 (O_864,N_4966,N_4793);
nor UO_865 (O_865,N_4797,N_4904);
or UO_866 (O_866,N_4918,N_4768);
or UO_867 (O_867,N_4953,N_4561);
or UO_868 (O_868,N_4996,N_4727);
or UO_869 (O_869,N_4970,N_4535);
and UO_870 (O_870,N_4635,N_4849);
nand UO_871 (O_871,N_4922,N_4839);
and UO_872 (O_872,N_4608,N_4598);
nand UO_873 (O_873,N_4809,N_4706);
or UO_874 (O_874,N_4560,N_4601);
nor UO_875 (O_875,N_4896,N_4743);
nand UO_876 (O_876,N_4699,N_4973);
and UO_877 (O_877,N_4755,N_4774);
and UO_878 (O_878,N_4607,N_4984);
nor UO_879 (O_879,N_4677,N_4861);
or UO_880 (O_880,N_4691,N_4909);
nand UO_881 (O_881,N_4526,N_4592);
nor UO_882 (O_882,N_4978,N_4858);
and UO_883 (O_883,N_4620,N_4539);
nand UO_884 (O_884,N_4708,N_4540);
nor UO_885 (O_885,N_4561,N_4619);
nor UO_886 (O_886,N_4891,N_4790);
nand UO_887 (O_887,N_4701,N_4967);
nand UO_888 (O_888,N_4756,N_4617);
nand UO_889 (O_889,N_4650,N_4744);
or UO_890 (O_890,N_4557,N_4822);
and UO_891 (O_891,N_4543,N_4732);
nor UO_892 (O_892,N_4607,N_4510);
xor UO_893 (O_893,N_4619,N_4732);
nand UO_894 (O_894,N_4703,N_4887);
nand UO_895 (O_895,N_4984,N_4995);
and UO_896 (O_896,N_4728,N_4790);
nor UO_897 (O_897,N_4955,N_4735);
nor UO_898 (O_898,N_4565,N_4965);
or UO_899 (O_899,N_4626,N_4900);
or UO_900 (O_900,N_4638,N_4724);
and UO_901 (O_901,N_4721,N_4853);
nor UO_902 (O_902,N_4932,N_4814);
nor UO_903 (O_903,N_4781,N_4990);
nor UO_904 (O_904,N_4772,N_4674);
nand UO_905 (O_905,N_4650,N_4718);
nand UO_906 (O_906,N_4824,N_4626);
nand UO_907 (O_907,N_4623,N_4767);
nor UO_908 (O_908,N_4672,N_4664);
nor UO_909 (O_909,N_4792,N_4764);
nor UO_910 (O_910,N_4529,N_4976);
xnor UO_911 (O_911,N_4711,N_4752);
or UO_912 (O_912,N_4985,N_4757);
and UO_913 (O_913,N_4567,N_4973);
nand UO_914 (O_914,N_4591,N_4567);
nor UO_915 (O_915,N_4854,N_4615);
or UO_916 (O_916,N_4566,N_4671);
nor UO_917 (O_917,N_4563,N_4514);
or UO_918 (O_918,N_4938,N_4751);
and UO_919 (O_919,N_4938,N_4817);
nor UO_920 (O_920,N_4962,N_4846);
or UO_921 (O_921,N_4943,N_4564);
nand UO_922 (O_922,N_4983,N_4684);
and UO_923 (O_923,N_4981,N_4668);
xnor UO_924 (O_924,N_4685,N_4831);
nand UO_925 (O_925,N_4828,N_4650);
nand UO_926 (O_926,N_4749,N_4991);
nor UO_927 (O_927,N_4692,N_4617);
or UO_928 (O_928,N_4536,N_4546);
or UO_929 (O_929,N_4535,N_4597);
or UO_930 (O_930,N_4755,N_4854);
and UO_931 (O_931,N_4710,N_4978);
nor UO_932 (O_932,N_4956,N_4687);
and UO_933 (O_933,N_4697,N_4983);
nor UO_934 (O_934,N_4971,N_4948);
nor UO_935 (O_935,N_4899,N_4875);
and UO_936 (O_936,N_4756,N_4812);
nor UO_937 (O_937,N_4682,N_4891);
and UO_938 (O_938,N_4588,N_4523);
nor UO_939 (O_939,N_4569,N_4980);
or UO_940 (O_940,N_4532,N_4641);
or UO_941 (O_941,N_4889,N_4578);
nand UO_942 (O_942,N_4790,N_4917);
nand UO_943 (O_943,N_4869,N_4959);
and UO_944 (O_944,N_4515,N_4657);
nor UO_945 (O_945,N_4743,N_4685);
nor UO_946 (O_946,N_4758,N_4633);
nor UO_947 (O_947,N_4965,N_4813);
nor UO_948 (O_948,N_4907,N_4882);
and UO_949 (O_949,N_4741,N_4500);
nor UO_950 (O_950,N_4793,N_4915);
nor UO_951 (O_951,N_4997,N_4877);
or UO_952 (O_952,N_4852,N_4656);
nand UO_953 (O_953,N_4607,N_4606);
nor UO_954 (O_954,N_4990,N_4966);
and UO_955 (O_955,N_4931,N_4771);
nand UO_956 (O_956,N_4879,N_4611);
nand UO_957 (O_957,N_4682,N_4822);
or UO_958 (O_958,N_4654,N_4909);
nand UO_959 (O_959,N_4982,N_4533);
nand UO_960 (O_960,N_4550,N_4950);
or UO_961 (O_961,N_4866,N_4878);
nor UO_962 (O_962,N_4863,N_4832);
nand UO_963 (O_963,N_4739,N_4710);
or UO_964 (O_964,N_4747,N_4819);
or UO_965 (O_965,N_4734,N_4851);
and UO_966 (O_966,N_4848,N_4774);
and UO_967 (O_967,N_4995,N_4722);
or UO_968 (O_968,N_4664,N_4602);
nand UO_969 (O_969,N_4926,N_4951);
and UO_970 (O_970,N_4952,N_4756);
or UO_971 (O_971,N_4585,N_4632);
and UO_972 (O_972,N_4902,N_4991);
nand UO_973 (O_973,N_4719,N_4592);
or UO_974 (O_974,N_4608,N_4939);
nand UO_975 (O_975,N_4807,N_4541);
and UO_976 (O_976,N_4920,N_4563);
nor UO_977 (O_977,N_4888,N_4502);
nor UO_978 (O_978,N_4672,N_4560);
nor UO_979 (O_979,N_4560,N_4540);
nor UO_980 (O_980,N_4852,N_4702);
or UO_981 (O_981,N_4596,N_4501);
nor UO_982 (O_982,N_4803,N_4929);
and UO_983 (O_983,N_4968,N_4875);
and UO_984 (O_984,N_4645,N_4757);
nor UO_985 (O_985,N_4591,N_4876);
nor UO_986 (O_986,N_4689,N_4511);
and UO_987 (O_987,N_4784,N_4886);
and UO_988 (O_988,N_4787,N_4856);
or UO_989 (O_989,N_4711,N_4869);
and UO_990 (O_990,N_4832,N_4930);
nor UO_991 (O_991,N_4964,N_4571);
nand UO_992 (O_992,N_4732,N_4727);
nor UO_993 (O_993,N_4721,N_4757);
nand UO_994 (O_994,N_4556,N_4970);
and UO_995 (O_995,N_4843,N_4682);
or UO_996 (O_996,N_4750,N_4879);
nor UO_997 (O_997,N_4865,N_4626);
or UO_998 (O_998,N_4607,N_4904);
nand UO_999 (O_999,N_4592,N_4921);
endmodule