module basic_1000_10000_1500_20_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_978,In_326);
and U1 (N_1,In_426,In_351);
nor U2 (N_2,In_303,In_700);
or U3 (N_3,In_840,In_831);
or U4 (N_4,In_730,In_21);
xor U5 (N_5,In_740,In_844);
nand U6 (N_6,In_176,In_557);
or U7 (N_7,In_886,In_569);
nor U8 (N_8,In_735,In_500);
and U9 (N_9,In_245,In_954);
and U10 (N_10,In_698,In_935);
or U11 (N_11,In_342,In_533);
or U12 (N_12,In_504,In_145);
xor U13 (N_13,In_617,In_763);
nand U14 (N_14,In_593,In_339);
or U15 (N_15,In_572,In_251);
nand U16 (N_16,In_933,In_919);
nand U17 (N_17,In_911,In_729);
xor U18 (N_18,In_415,In_109);
nor U19 (N_19,In_794,In_389);
nand U20 (N_20,In_937,In_237);
or U21 (N_21,In_535,In_129);
and U22 (N_22,In_489,In_51);
and U23 (N_23,In_548,In_728);
nor U24 (N_24,In_519,In_272);
xnor U25 (N_25,In_90,In_287);
and U26 (N_26,In_475,In_545);
or U27 (N_27,In_638,In_725);
nand U28 (N_28,In_770,In_95);
xor U29 (N_29,In_715,In_455);
or U30 (N_30,In_456,In_396);
and U31 (N_31,In_521,In_139);
nor U32 (N_32,In_822,In_970);
xor U33 (N_33,In_880,In_12);
nor U34 (N_34,In_589,In_927);
or U35 (N_35,In_819,In_391);
and U36 (N_36,In_946,In_57);
and U37 (N_37,In_513,In_140);
or U38 (N_38,In_321,In_163);
nor U39 (N_39,In_741,In_515);
and U40 (N_40,In_767,In_153);
xor U41 (N_41,In_848,In_25);
xnor U42 (N_42,In_923,In_590);
or U43 (N_43,In_731,In_874);
or U44 (N_44,In_266,In_601);
nand U45 (N_45,In_256,In_657);
and U46 (N_46,In_616,In_688);
nor U47 (N_47,In_639,In_812);
nand U48 (N_48,In_713,In_422);
xnor U49 (N_49,In_193,In_520);
nand U50 (N_50,In_184,In_828);
or U51 (N_51,In_486,In_746);
and U52 (N_52,In_214,In_296);
or U53 (N_53,In_580,In_119);
or U54 (N_54,In_663,In_79);
xor U55 (N_55,In_733,In_228);
nor U56 (N_56,In_753,In_567);
nor U57 (N_57,In_853,In_654);
nand U58 (N_58,In_563,In_642);
nand U59 (N_59,In_449,In_434);
and U60 (N_60,In_641,In_527);
nor U61 (N_61,In_181,In_706);
nand U62 (N_62,In_464,In_39);
and U63 (N_63,In_634,In_30);
and U64 (N_64,In_373,In_930);
nor U65 (N_65,In_273,In_277);
xor U66 (N_66,In_877,In_755);
and U67 (N_67,In_405,In_227);
nor U68 (N_68,In_661,In_483);
nand U69 (N_69,In_438,In_268);
nand U70 (N_70,In_439,In_827);
xor U71 (N_71,In_627,In_28);
nand U72 (N_72,In_726,In_155);
nand U73 (N_73,In_189,In_673);
and U74 (N_74,In_292,In_487);
and U75 (N_75,In_843,In_143);
or U76 (N_76,In_530,In_727);
xor U77 (N_77,In_84,In_141);
nor U78 (N_78,In_187,In_879);
xnor U79 (N_79,In_311,In_855);
nand U80 (N_80,In_103,In_199);
or U81 (N_81,In_402,In_1);
nand U82 (N_82,In_918,In_959);
and U83 (N_83,In_159,In_156);
nand U84 (N_84,In_85,In_556);
nor U85 (N_85,In_404,In_512);
and U86 (N_86,In_470,In_818);
and U87 (N_87,In_117,In_416);
or U88 (N_88,In_33,In_86);
and U89 (N_89,In_357,In_480);
nand U90 (N_90,In_604,In_742);
or U91 (N_91,In_795,In_197);
and U92 (N_92,In_211,In_766);
and U93 (N_93,In_826,In_99);
nand U94 (N_94,In_329,In_297);
or U95 (N_95,In_150,In_349);
and U96 (N_96,In_757,In_429);
nand U97 (N_97,In_413,In_88);
nand U98 (N_98,In_288,In_125);
nor U99 (N_99,In_101,In_204);
nor U100 (N_100,In_255,In_330);
nor U101 (N_101,In_111,In_104);
nor U102 (N_102,In_932,In_680);
and U103 (N_103,In_909,In_461);
or U104 (N_104,In_369,In_687);
or U105 (N_105,In_550,In_575);
or U106 (N_106,In_11,In_246);
nand U107 (N_107,In_171,In_465);
and U108 (N_108,In_518,In_242);
or U109 (N_109,In_577,In_793);
and U110 (N_110,In_136,In_560);
or U111 (N_111,In_825,In_234);
or U112 (N_112,In_397,In_218);
xor U113 (N_113,In_913,In_867);
or U114 (N_114,In_714,In_154);
nor U115 (N_115,In_683,In_46);
and U116 (N_116,In_360,In_705);
xnor U117 (N_117,In_35,In_985);
or U118 (N_118,In_926,In_137);
nor U119 (N_119,In_953,In_161);
or U120 (N_120,In_442,In_398);
xnor U121 (N_121,In_230,In_80);
xnor U122 (N_122,In_23,In_865);
xor U123 (N_123,In_325,In_942);
nand U124 (N_124,In_903,In_192);
nand U125 (N_125,In_804,In_891);
and U126 (N_126,In_578,In_356);
nand U127 (N_127,In_463,In_717);
or U128 (N_128,In_291,In_643);
or U129 (N_129,In_447,In_586);
and U130 (N_130,In_681,In_710);
nand U131 (N_131,In_510,In_365);
nor U132 (N_132,In_36,In_957);
and U133 (N_133,In_83,In_724);
xor U134 (N_134,In_559,In_162);
and U135 (N_135,In_89,In_528);
nor U136 (N_136,In_996,In_372);
nor U137 (N_137,In_183,In_40);
and U138 (N_138,In_829,In_780);
xor U139 (N_139,In_409,In_453);
xnor U140 (N_140,In_363,In_249);
and U141 (N_141,In_212,In_987);
or U142 (N_142,In_802,In_784);
xnor U143 (N_143,In_789,In_202);
nor U144 (N_144,In_179,In_842);
or U145 (N_145,In_158,In_252);
and U146 (N_146,In_536,In_947);
or U147 (N_147,In_364,In_446);
nand U148 (N_148,In_846,In_223);
or U149 (N_149,In_400,In_629);
or U150 (N_150,In_54,In_595);
nand U151 (N_151,In_979,In_152);
nand U152 (N_152,In_116,In_368);
or U153 (N_153,In_293,In_613);
or U154 (N_154,In_259,In_34);
nand U155 (N_155,In_379,In_597);
nor U156 (N_156,In_221,In_612);
nor U157 (N_157,In_554,In_943);
nand U158 (N_158,In_602,In_749);
nand U159 (N_159,In_824,In_10);
nand U160 (N_160,In_336,In_8);
and U161 (N_161,In_546,In_838);
nor U162 (N_162,In_587,In_649);
nor U163 (N_163,In_509,In_474);
and U164 (N_164,In_219,In_123);
and U165 (N_165,In_241,In_931);
xor U166 (N_166,In_526,In_236);
or U167 (N_167,In_902,In_581);
xor U168 (N_168,In_722,In_801);
or U169 (N_169,In_60,In_320);
nor U170 (N_170,In_543,In_863);
or U171 (N_171,In_823,In_561);
xnor U172 (N_172,In_693,In_149);
nor U173 (N_173,In_186,In_315);
or U174 (N_174,In_967,In_873);
or U175 (N_175,In_185,In_70);
nand U176 (N_176,In_854,In_458);
or U177 (N_177,In_542,In_977);
nor U178 (N_178,In_924,In_883);
nand U179 (N_179,In_424,In_170);
xnor U180 (N_180,In_45,In_870);
nor U181 (N_181,In_66,In_997);
nor U182 (N_182,In_275,In_188);
nand U183 (N_183,In_989,In_382);
xnor U184 (N_184,In_632,In_395);
nor U185 (N_185,In_748,In_490);
and U186 (N_186,In_477,In_875);
nor U187 (N_187,In_645,In_745);
and U188 (N_188,In_696,In_882);
nor U189 (N_189,In_852,In_91);
xnor U190 (N_190,In_380,In_956);
and U191 (N_191,In_232,In_42);
and U192 (N_192,In_999,In_459);
or U193 (N_193,In_872,In_410);
xor U194 (N_194,In_492,In_841);
and U195 (N_195,In_899,In_0);
nand U196 (N_196,In_318,In_427);
xor U197 (N_197,In_120,In_418);
or U198 (N_198,In_984,In_226);
and U199 (N_199,In_55,In_102);
and U200 (N_200,In_350,In_113);
nand U201 (N_201,In_760,In_386);
nand U202 (N_202,In_553,In_220);
nor U203 (N_203,In_114,In_274);
nand U204 (N_204,In_614,In_355);
nor U205 (N_205,In_282,In_544);
nor U206 (N_206,In_790,In_235);
nor U207 (N_207,In_37,In_626);
nand U208 (N_208,In_945,In_267);
nand U209 (N_209,In_132,In_988);
or U210 (N_210,In_312,In_169);
or U211 (N_211,In_408,In_962);
nor U212 (N_212,In_276,In_63);
xnor U213 (N_213,In_306,In_15);
nor U214 (N_214,In_343,In_96);
nor U215 (N_215,In_478,In_624);
xnor U216 (N_216,In_885,In_920);
or U217 (N_217,In_87,In_704);
nand U218 (N_218,In_914,In_271);
and U219 (N_219,In_625,In_534);
and U220 (N_220,In_417,In_743);
or U221 (N_221,In_777,In_805);
nand U222 (N_222,In_836,In_44);
nand U223 (N_223,In_655,In_720);
and U224 (N_224,In_280,In_635);
and U225 (N_225,In_32,In_866);
nor U226 (N_226,In_283,In_603);
nor U227 (N_227,In_662,In_319);
and U228 (N_228,In_623,In_340);
xnor U229 (N_229,In_305,In_423);
nand U230 (N_230,In_570,In_507);
xnor U231 (N_231,In_253,In_61);
nor U232 (N_232,In_332,In_172);
nor U233 (N_233,In_195,In_890);
or U234 (N_234,In_532,In_815);
nor U235 (N_235,In_868,In_205);
nor U236 (N_236,In_367,In_168);
nand U237 (N_237,In_936,In_958);
or U238 (N_238,In_494,In_495);
and U239 (N_239,In_975,In_652);
or U240 (N_240,In_265,In_961);
and U241 (N_241,In_76,In_19);
nor U242 (N_242,In_750,In_778);
nor U243 (N_243,In_56,In_301);
and U244 (N_244,In_980,In_191);
or U245 (N_245,In_651,In_26);
nand U246 (N_246,In_862,In_881);
nand U247 (N_247,In_765,In_327);
xor U248 (N_248,In_732,In_991);
nor U249 (N_249,In_524,In_194);
xnor U250 (N_250,In_74,In_75);
xor U251 (N_251,In_562,In_501);
xor U252 (N_252,In_4,In_243);
nand U253 (N_253,In_498,In_290);
nor U254 (N_254,In_531,In_514);
xnor U255 (N_255,In_122,In_224);
and U256 (N_256,In_52,In_16);
nor U257 (N_257,In_250,In_529);
nor U258 (N_258,In_506,In_262);
xor U259 (N_259,In_460,In_738);
and U260 (N_260,In_497,In_403);
and U261 (N_261,In_38,In_485);
nand U262 (N_262,In_960,In_547);
nor U263 (N_263,In_7,In_166);
nor U264 (N_264,In_915,In_678);
xor U265 (N_265,In_257,In_739);
or U266 (N_266,In_47,In_371);
nor U267 (N_267,In_381,In_261);
xor U268 (N_268,In_322,In_686);
nand U269 (N_269,In_955,In_517);
or U270 (N_270,In_944,In_647);
nor U271 (N_271,In_650,In_279);
xnor U272 (N_272,In_43,In_345);
nand U273 (N_273,In_938,In_664);
xnor U274 (N_274,In_974,In_433);
xnor U275 (N_275,In_631,In_414);
nand U276 (N_276,In_736,In_177);
or U277 (N_277,In_289,In_965);
and U278 (N_278,In_338,In_94);
nor U279 (N_279,In_708,In_799);
and U280 (N_280,In_685,In_203);
nand U281 (N_281,In_49,In_448);
nor U282 (N_282,In_800,In_806);
nand U283 (N_283,In_734,In_896);
and U284 (N_284,In_180,In_467);
and U285 (N_285,In_344,In_860);
or U286 (N_286,In_796,In_737);
or U287 (N_287,In_348,In_648);
nor U288 (N_288,In_248,In_399);
nor U289 (N_289,In_952,In_718);
or U290 (N_290,In_674,In_670);
xnor U291 (N_291,In_951,In_508);
nor U292 (N_292,In_59,In_582);
xor U293 (N_293,In_759,In_24);
and U294 (N_294,In_555,In_637);
xnor U295 (N_295,In_69,In_479);
nor U296 (N_296,In_392,In_768);
or U297 (N_297,In_353,In_549);
xnor U298 (N_298,In_845,In_895);
or U299 (N_299,In_949,In_393);
nor U300 (N_300,In_747,In_901);
xor U301 (N_301,In_928,In_995);
nand U302 (N_302,In_756,In_209);
or U303 (N_303,In_107,In_67);
nand U304 (N_304,In_317,In_68);
xor U305 (N_305,In_13,In_201);
or U306 (N_306,In_27,In_151);
nand U307 (N_307,In_869,In_50);
nand U308 (N_308,In_254,In_898);
nor U309 (N_309,In_31,In_551);
nor U310 (N_310,In_144,In_900);
or U311 (N_311,In_752,In_502);
nand U312 (N_312,In_659,In_973);
and U313 (N_313,In_665,In_208);
nand U314 (N_314,In_105,In_803);
xnor U315 (N_315,In_244,In_771);
and U316 (N_316,In_964,In_335);
or U317 (N_317,In_976,In_830);
and U318 (N_318,In_668,In_309);
or U319 (N_319,In_981,In_912);
nor U320 (N_320,In_231,In_892);
and U321 (N_321,In_934,In_878);
xnor U322 (N_322,In_761,In_849);
xnor U323 (N_323,In_412,In_676);
nand U324 (N_324,In_834,In_993);
nor U325 (N_325,In_904,In_764);
nor U326 (N_326,In_217,In_247);
nor U327 (N_327,In_14,In_142);
nor U328 (N_328,In_295,In_482);
nand U329 (N_329,In_376,In_440);
or U330 (N_330,In_505,In_971);
and U331 (N_331,In_472,In_260);
xnor U332 (N_332,In_797,In_135);
nor U333 (N_333,In_695,In_488);
and U334 (N_334,In_270,In_916);
or U335 (N_335,In_798,In_432);
and U336 (N_336,In_388,In_471);
xnor U337 (N_337,In_175,In_22);
nor U338 (N_338,In_640,In_697);
xor U339 (N_339,In_711,In_894);
or U340 (N_340,In_112,In_889);
or U341 (N_341,In_78,In_907);
and U342 (N_342,In_299,In_887);
nor U343 (N_343,In_691,In_876);
xor U344 (N_344,In_628,In_240);
nand U345 (N_345,In_592,In_484);
or U346 (N_346,In_791,In_630);
and U347 (N_347,In_857,In_174);
or U348 (N_348,In_584,In_128);
and U349 (N_349,In_127,In_775);
nor U350 (N_350,In_148,In_307);
or U351 (N_351,In_782,In_98);
nor U352 (N_352,In_374,In_682);
and U353 (N_353,In_552,In_82);
xnor U354 (N_354,In_222,In_390);
xnor U355 (N_355,In_281,In_333);
nor U356 (N_356,In_476,In_182);
nand U357 (N_357,In_607,In_690);
nor U358 (N_358,In_523,In_354);
or U359 (N_359,In_566,In_576);
nor U360 (N_360,In_646,In_568);
or U361 (N_361,In_383,In_701);
and U362 (N_362,In_92,In_58);
or U363 (N_363,In_888,In_998);
or U364 (N_364,In_164,In_821);
or U365 (N_365,In_787,In_384);
or U366 (N_366,In_337,In_751);
and U367 (N_367,In_198,In_20);
and U368 (N_368,In_675,In_130);
nor U369 (N_369,In_776,In_658);
and U370 (N_370,In_666,In_864);
and U371 (N_371,In_377,In_917);
or U372 (N_372,In_361,In_493);
and U373 (N_373,In_769,In_983);
or U374 (N_374,In_200,In_859);
or U375 (N_375,In_157,In_407);
and U376 (N_376,In_48,In_81);
and U377 (N_377,In_788,In_18);
nand U378 (N_378,In_814,In_540);
nand U379 (N_379,In_516,In_709);
and U380 (N_380,In_622,In_839);
nand U381 (N_381,In_394,In_147);
nand U382 (N_382,In_263,In_950);
nor U383 (N_383,In_167,In_366);
or U384 (N_384,In_437,In_660);
and U385 (N_385,In_615,In_452);
xor U386 (N_386,In_385,In_588);
nor U387 (N_387,In_445,In_565);
or U388 (N_388,In_62,In_963);
or U389 (N_389,In_5,In_611);
or U390 (N_390,In_454,In_994);
and U391 (N_391,In_608,In_126);
and U392 (N_392,In_115,In_605);
or U393 (N_393,In_972,In_421);
and U394 (N_394,In_851,In_284);
and U395 (N_395,In_419,In_832);
nand U396 (N_396,In_905,In_702);
nor U397 (N_397,In_431,In_100);
xnor U398 (N_398,In_134,In_178);
and U399 (N_399,In_481,In_539);
and U400 (N_400,In_897,In_810);
nor U401 (N_401,In_346,In_466);
or U402 (N_402,In_165,In_196);
or U403 (N_403,In_990,In_334);
nor U404 (N_404,In_893,In_302);
xor U405 (N_405,In_537,In_636);
or U406 (N_406,In_310,In_451);
nor U407 (N_407,In_966,In_286);
nor U408 (N_408,In_331,In_411);
and U409 (N_409,In_656,In_378);
or U410 (N_410,In_375,In_571);
nand U411 (N_411,In_758,In_968);
nand U412 (N_412,In_807,In_77);
nor U413 (N_413,In_689,In_406);
xor U414 (N_414,In_837,In_712);
or U415 (N_415,In_856,In_131);
nand U416 (N_416,In_430,In_969);
nand U417 (N_417,In_992,In_352);
or U418 (N_418,In_583,In_744);
nand U419 (N_419,In_817,In_925);
and U420 (N_420,In_621,In_72);
xnor U421 (N_421,In_591,In_285);
or U422 (N_422,In_216,In_847);
nand U423 (N_423,In_772,In_239);
xnor U424 (N_424,In_347,In_215);
nor U425 (N_425,In_564,In_473);
nor U426 (N_426,In_206,In_316);
xor U427 (N_427,In_370,In_618);
nand U428 (N_428,In_229,In_816);
or U429 (N_429,In_619,In_6);
nand U430 (N_430,In_213,In_41);
nand U431 (N_431,In_792,In_541);
xnor U432 (N_432,In_762,In_667);
or U433 (N_433,In_341,In_820);
and U434 (N_434,In_65,In_594);
nand U435 (N_435,In_677,In_225);
or U436 (N_436,In_754,In_986);
nand U437 (N_437,In_190,In_17);
nand U438 (N_438,In_133,In_358);
xor U439 (N_439,In_558,In_929);
or U440 (N_440,In_278,In_684);
xor U441 (N_441,In_138,In_585);
nand U442 (N_442,In_910,In_644);
or U443 (N_443,In_450,In_64);
nor U444 (N_444,In_721,In_359);
or U445 (N_445,In_443,In_941);
or U446 (N_446,In_323,In_29);
or U447 (N_447,In_146,In_97);
nand U448 (N_448,In_922,In_574);
nand U449 (N_449,In_858,In_939);
nor U450 (N_450,In_719,In_948);
and U451 (N_451,In_811,In_813);
nor U452 (N_452,In_457,In_884);
nand U453 (N_453,In_210,In_362);
or U454 (N_454,In_420,In_633);
or U455 (N_455,In_600,In_462);
nand U456 (N_456,In_982,In_444);
nor U457 (N_457,In_786,In_850);
xor U458 (N_458,In_469,In_703);
or U459 (N_459,In_833,In_671);
nand U460 (N_460,In_707,In_921);
xnor U461 (N_461,In_783,In_436);
xor U462 (N_462,In_596,In_908);
nor U463 (N_463,In_672,In_906);
or U464 (N_464,In_579,In_233);
and U465 (N_465,In_106,In_2);
xnor U466 (N_466,In_108,In_499);
and U467 (N_467,In_328,In_9);
xnor U468 (N_468,In_781,In_606);
nand U469 (N_469,In_298,In_468);
and U470 (N_470,In_53,In_238);
xnor U471 (N_471,In_522,In_491);
xor U472 (N_472,In_679,In_773);
and U473 (N_473,In_428,In_653);
nand U474 (N_474,In_313,In_861);
nor U475 (N_475,In_324,In_610);
or U476 (N_476,In_314,In_496);
and U477 (N_477,In_809,In_264);
xor U478 (N_478,In_503,In_425);
and U479 (N_479,In_835,In_620);
xor U480 (N_480,In_173,In_93);
nand U481 (N_481,In_387,In_124);
and U482 (N_482,In_207,In_808);
nor U483 (N_483,In_692,In_716);
nor U484 (N_484,In_118,In_669);
xnor U485 (N_485,In_511,In_785);
or U486 (N_486,In_308,In_940);
nand U487 (N_487,In_525,In_779);
nand U488 (N_488,In_598,In_723);
nand U489 (N_489,In_435,In_699);
or U490 (N_490,In_71,In_401);
xor U491 (N_491,In_294,In_694);
nor U492 (N_492,In_160,In_3);
nor U493 (N_493,In_871,In_121);
or U494 (N_494,In_110,In_258);
and U495 (N_495,In_599,In_304);
xor U496 (N_496,In_73,In_269);
and U497 (N_497,In_573,In_774);
nor U498 (N_498,In_441,In_300);
nor U499 (N_499,In_538,In_609);
xor U500 (N_500,N_458,N_119);
and U501 (N_501,N_141,N_483);
and U502 (N_502,N_152,N_164);
nor U503 (N_503,N_475,N_111);
nor U504 (N_504,N_175,N_27);
or U505 (N_505,N_12,N_346);
xnor U506 (N_506,N_138,N_278);
or U507 (N_507,N_373,N_344);
xnor U508 (N_508,N_364,N_279);
xor U509 (N_509,N_95,N_424);
and U510 (N_510,N_441,N_15);
nand U511 (N_511,N_228,N_133);
or U512 (N_512,N_492,N_7);
or U513 (N_513,N_24,N_480);
nand U514 (N_514,N_334,N_67);
xnor U515 (N_515,N_137,N_429);
and U516 (N_516,N_491,N_333);
xnor U517 (N_517,N_257,N_470);
and U518 (N_518,N_244,N_230);
or U519 (N_519,N_390,N_19);
or U520 (N_520,N_265,N_487);
xnor U521 (N_521,N_339,N_394);
nor U522 (N_522,N_358,N_253);
nand U523 (N_523,N_497,N_303);
xnor U524 (N_524,N_290,N_146);
and U525 (N_525,N_467,N_147);
or U526 (N_526,N_326,N_255);
nor U527 (N_527,N_311,N_272);
nor U528 (N_528,N_476,N_362);
nor U529 (N_529,N_204,N_238);
and U530 (N_530,N_50,N_430);
xnor U531 (N_531,N_347,N_450);
nand U532 (N_532,N_182,N_155);
nand U533 (N_533,N_374,N_348);
and U534 (N_534,N_325,N_336);
nand U535 (N_535,N_163,N_337);
and U536 (N_536,N_454,N_335);
nand U537 (N_537,N_8,N_360);
nand U538 (N_538,N_150,N_74);
nor U539 (N_539,N_332,N_202);
nor U540 (N_540,N_384,N_271);
or U541 (N_541,N_187,N_256);
or U542 (N_542,N_401,N_149);
or U543 (N_543,N_183,N_40);
and U544 (N_544,N_295,N_59);
and U545 (N_545,N_100,N_197);
nand U546 (N_546,N_203,N_341);
nor U547 (N_547,N_157,N_165);
and U548 (N_548,N_105,N_75);
and U549 (N_549,N_453,N_456);
and U550 (N_550,N_222,N_385);
xor U551 (N_551,N_215,N_386);
and U552 (N_552,N_220,N_324);
and U553 (N_553,N_35,N_103);
or U554 (N_554,N_414,N_52);
xor U555 (N_555,N_304,N_323);
or U556 (N_556,N_134,N_104);
nor U557 (N_557,N_299,N_393);
xnor U558 (N_558,N_315,N_32);
and U559 (N_559,N_208,N_353);
nand U560 (N_560,N_479,N_387);
xor U561 (N_561,N_76,N_248);
nor U562 (N_562,N_190,N_411);
nor U563 (N_563,N_34,N_468);
or U564 (N_564,N_116,N_498);
nand U565 (N_565,N_107,N_41);
and U566 (N_566,N_136,N_478);
and U567 (N_567,N_170,N_158);
and U568 (N_568,N_367,N_345);
xnor U569 (N_569,N_375,N_53);
nand U570 (N_570,N_406,N_145);
xor U571 (N_571,N_285,N_433);
and U572 (N_572,N_57,N_397);
nor U573 (N_573,N_263,N_51);
nand U574 (N_574,N_122,N_378);
nand U575 (N_575,N_437,N_457);
xor U576 (N_576,N_464,N_440);
or U577 (N_577,N_366,N_110);
nor U578 (N_578,N_319,N_160);
nor U579 (N_579,N_260,N_308);
and U580 (N_580,N_317,N_232);
nand U581 (N_581,N_269,N_445);
or U582 (N_582,N_28,N_338);
or U583 (N_583,N_350,N_313);
nor U584 (N_584,N_184,N_188);
nor U585 (N_585,N_365,N_417);
nand U586 (N_586,N_212,N_143);
nor U587 (N_587,N_247,N_493);
or U588 (N_588,N_6,N_206);
and U589 (N_589,N_114,N_77);
xor U590 (N_590,N_473,N_224);
nand U591 (N_591,N_415,N_148);
or U592 (N_592,N_455,N_259);
or U593 (N_593,N_0,N_402);
and U594 (N_594,N_249,N_472);
or U595 (N_595,N_490,N_210);
nand U596 (N_596,N_274,N_11);
nor U597 (N_597,N_217,N_398);
xor U598 (N_598,N_29,N_356);
xor U599 (N_599,N_139,N_292);
and U600 (N_600,N_55,N_70);
xnor U601 (N_601,N_426,N_185);
and U602 (N_602,N_460,N_209);
nand U603 (N_603,N_245,N_236);
xnor U604 (N_604,N_132,N_276);
and U605 (N_605,N_83,N_49);
nor U606 (N_606,N_250,N_225);
nand U607 (N_607,N_93,N_471);
or U608 (N_608,N_258,N_286);
nand U609 (N_609,N_38,N_156);
nand U610 (N_610,N_72,N_180);
nor U611 (N_611,N_425,N_316);
nand U612 (N_612,N_444,N_408);
or U613 (N_613,N_307,N_305);
xnor U614 (N_614,N_294,N_101);
nand U615 (N_615,N_314,N_30);
xnor U616 (N_616,N_115,N_89);
xor U617 (N_617,N_465,N_399);
nor U618 (N_618,N_283,N_140);
xnor U619 (N_619,N_173,N_25);
or U620 (N_620,N_392,N_466);
xor U621 (N_621,N_351,N_439);
or U622 (N_622,N_126,N_17);
xnor U623 (N_623,N_131,N_376);
nor U624 (N_624,N_291,N_79);
and U625 (N_625,N_391,N_484);
nand U626 (N_626,N_380,N_186);
and U627 (N_627,N_62,N_127);
or U628 (N_628,N_481,N_112);
and U629 (N_629,N_43,N_462);
xor U630 (N_630,N_297,N_58);
and U631 (N_631,N_166,N_64);
or U632 (N_632,N_428,N_80);
nor U633 (N_633,N_71,N_306);
nor U634 (N_634,N_194,N_388);
or U635 (N_635,N_69,N_289);
nor U636 (N_636,N_85,N_177);
nand U637 (N_637,N_407,N_342);
and U638 (N_638,N_423,N_461);
nand U639 (N_639,N_495,N_205);
and U640 (N_640,N_310,N_239);
and U641 (N_641,N_192,N_45);
xnor U642 (N_642,N_68,N_262);
and U643 (N_643,N_370,N_14);
nor U644 (N_644,N_161,N_409);
or U645 (N_645,N_389,N_92);
xnor U646 (N_646,N_125,N_113);
and U647 (N_647,N_447,N_412);
xnor U648 (N_648,N_355,N_296);
or U649 (N_649,N_178,N_282);
nor U650 (N_650,N_3,N_382);
or U651 (N_651,N_494,N_97);
xor U652 (N_652,N_168,N_486);
xnor U653 (N_653,N_331,N_432);
nor U654 (N_654,N_434,N_328);
nor U655 (N_655,N_78,N_96);
xnor U656 (N_656,N_267,N_176);
nand U657 (N_657,N_442,N_237);
and U658 (N_658,N_88,N_416);
and U659 (N_659,N_159,N_54);
xor U660 (N_660,N_82,N_31);
nor U661 (N_661,N_363,N_223);
or U662 (N_662,N_233,N_235);
nand U663 (N_663,N_443,N_354);
nand U664 (N_664,N_56,N_422);
xnor U665 (N_665,N_18,N_129);
and U666 (N_666,N_193,N_118);
nor U667 (N_667,N_329,N_266);
and U668 (N_668,N_372,N_469);
xor U669 (N_669,N_153,N_66);
nand U670 (N_670,N_9,N_270);
and U671 (N_671,N_10,N_26);
nor U672 (N_672,N_128,N_448);
xnor U673 (N_673,N_154,N_195);
nor U674 (N_674,N_214,N_162);
xor U675 (N_675,N_418,N_94);
nor U676 (N_676,N_48,N_167);
nor U677 (N_677,N_106,N_327);
and U678 (N_678,N_5,N_300);
nor U679 (N_679,N_117,N_254);
nor U680 (N_680,N_171,N_231);
nor U681 (N_681,N_144,N_135);
nand U682 (N_682,N_65,N_400);
or U683 (N_683,N_488,N_298);
nor U684 (N_684,N_446,N_102);
or U685 (N_685,N_301,N_37);
xor U686 (N_686,N_368,N_179);
nand U687 (N_687,N_361,N_169);
or U688 (N_688,N_280,N_309);
or U689 (N_689,N_436,N_482);
or U690 (N_690,N_485,N_451);
nand U691 (N_691,N_318,N_22);
or U692 (N_692,N_42,N_477);
or U693 (N_693,N_21,N_463);
nand U694 (N_694,N_381,N_90);
nor U695 (N_695,N_379,N_86);
and U696 (N_696,N_199,N_268);
and U697 (N_697,N_340,N_349);
nand U698 (N_698,N_13,N_275);
and U699 (N_699,N_4,N_405);
nor U700 (N_700,N_39,N_121);
nor U701 (N_701,N_63,N_449);
xor U702 (N_702,N_2,N_264);
xnor U703 (N_703,N_427,N_221);
xor U704 (N_704,N_240,N_383);
or U705 (N_705,N_73,N_284);
or U706 (N_706,N_142,N_420);
nor U707 (N_707,N_241,N_60);
nand U708 (N_708,N_281,N_343);
or U709 (N_709,N_20,N_251);
or U710 (N_710,N_352,N_229);
nor U711 (N_711,N_61,N_99);
or U712 (N_712,N_109,N_218);
nand U713 (N_713,N_261,N_452);
xor U714 (N_714,N_84,N_181);
and U715 (N_715,N_293,N_322);
nand U716 (N_716,N_211,N_321);
nor U717 (N_717,N_243,N_252);
or U718 (N_718,N_234,N_98);
and U719 (N_719,N_174,N_36);
nand U720 (N_720,N_46,N_16);
nor U721 (N_721,N_287,N_496);
nand U722 (N_722,N_312,N_23);
xnor U723 (N_723,N_273,N_87);
or U724 (N_724,N_120,N_302);
nand U725 (N_725,N_196,N_151);
nor U726 (N_726,N_44,N_216);
and U727 (N_727,N_219,N_499);
and U728 (N_728,N_213,N_320);
or U729 (N_729,N_201,N_459);
and U730 (N_730,N_191,N_371);
xnor U731 (N_731,N_47,N_123);
xnor U732 (N_732,N_130,N_489);
and U733 (N_733,N_200,N_357);
nand U734 (N_734,N_81,N_108);
xor U735 (N_735,N_377,N_438);
xnor U736 (N_736,N_359,N_421);
and U737 (N_737,N_288,N_474);
and U738 (N_738,N_435,N_403);
nor U739 (N_739,N_413,N_246);
xnor U740 (N_740,N_172,N_396);
nand U741 (N_741,N_124,N_226);
nand U742 (N_742,N_395,N_207);
nor U743 (N_743,N_404,N_227);
xnor U744 (N_744,N_419,N_1);
or U745 (N_745,N_369,N_242);
nand U746 (N_746,N_410,N_189);
and U747 (N_747,N_198,N_277);
xor U748 (N_748,N_91,N_33);
nor U749 (N_749,N_431,N_330);
nand U750 (N_750,N_321,N_312);
xor U751 (N_751,N_302,N_347);
nand U752 (N_752,N_445,N_411);
and U753 (N_753,N_302,N_349);
or U754 (N_754,N_410,N_227);
or U755 (N_755,N_209,N_112);
and U756 (N_756,N_247,N_38);
or U757 (N_757,N_164,N_310);
and U758 (N_758,N_411,N_25);
xnor U759 (N_759,N_415,N_121);
nor U760 (N_760,N_149,N_261);
and U761 (N_761,N_97,N_449);
or U762 (N_762,N_153,N_121);
nand U763 (N_763,N_31,N_395);
nand U764 (N_764,N_421,N_490);
nor U765 (N_765,N_415,N_96);
nor U766 (N_766,N_369,N_489);
xor U767 (N_767,N_364,N_467);
nand U768 (N_768,N_89,N_107);
and U769 (N_769,N_63,N_331);
or U770 (N_770,N_338,N_303);
nor U771 (N_771,N_84,N_22);
or U772 (N_772,N_323,N_276);
nor U773 (N_773,N_168,N_413);
and U774 (N_774,N_128,N_276);
or U775 (N_775,N_309,N_30);
nand U776 (N_776,N_136,N_116);
and U777 (N_777,N_181,N_236);
and U778 (N_778,N_349,N_137);
and U779 (N_779,N_391,N_186);
nand U780 (N_780,N_319,N_423);
and U781 (N_781,N_401,N_377);
nand U782 (N_782,N_255,N_474);
nor U783 (N_783,N_392,N_496);
nand U784 (N_784,N_75,N_7);
nor U785 (N_785,N_115,N_272);
nor U786 (N_786,N_11,N_227);
and U787 (N_787,N_491,N_59);
nand U788 (N_788,N_166,N_406);
or U789 (N_789,N_448,N_273);
xor U790 (N_790,N_284,N_445);
nand U791 (N_791,N_224,N_209);
and U792 (N_792,N_70,N_468);
nor U793 (N_793,N_35,N_357);
and U794 (N_794,N_484,N_301);
nand U795 (N_795,N_76,N_453);
xnor U796 (N_796,N_388,N_190);
nor U797 (N_797,N_439,N_95);
xnor U798 (N_798,N_17,N_74);
nor U799 (N_799,N_406,N_220);
and U800 (N_800,N_499,N_368);
nor U801 (N_801,N_377,N_95);
or U802 (N_802,N_185,N_14);
and U803 (N_803,N_159,N_363);
nor U804 (N_804,N_31,N_23);
or U805 (N_805,N_192,N_228);
xnor U806 (N_806,N_35,N_169);
xnor U807 (N_807,N_52,N_492);
and U808 (N_808,N_92,N_75);
and U809 (N_809,N_359,N_446);
xor U810 (N_810,N_151,N_416);
xnor U811 (N_811,N_315,N_215);
or U812 (N_812,N_404,N_123);
and U813 (N_813,N_267,N_327);
xor U814 (N_814,N_181,N_10);
nand U815 (N_815,N_305,N_266);
nor U816 (N_816,N_191,N_223);
or U817 (N_817,N_305,N_451);
xor U818 (N_818,N_290,N_84);
or U819 (N_819,N_285,N_38);
nor U820 (N_820,N_308,N_245);
and U821 (N_821,N_418,N_487);
or U822 (N_822,N_133,N_214);
nor U823 (N_823,N_52,N_27);
and U824 (N_824,N_469,N_70);
and U825 (N_825,N_269,N_325);
nand U826 (N_826,N_227,N_255);
nor U827 (N_827,N_87,N_421);
or U828 (N_828,N_157,N_40);
and U829 (N_829,N_36,N_399);
xor U830 (N_830,N_72,N_36);
nor U831 (N_831,N_64,N_181);
nand U832 (N_832,N_119,N_317);
nand U833 (N_833,N_448,N_490);
nand U834 (N_834,N_447,N_128);
and U835 (N_835,N_270,N_370);
xnor U836 (N_836,N_288,N_165);
or U837 (N_837,N_70,N_166);
and U838 (N_838,N_131,N_103);
nand U839 (N_839,N_168,N_222);
nand U840 (N_840,N_408,N_383);
and U841 (N_841,N_431,N_198);
nand U842 (N_842,N_374,N_450);
nand U843 (N_843,N_294,N_260);
and U844 (N_844,N_402,N_325);
nor U845 (N_845,N_263,N_460);
or U846 (N_846,N_490,N_191);
nor U847 (N_847,N_195,N_442);
xnor U848 (N_848,N_251,N_198);
nor U849 (N_849,N_338,N_158);
or U850 (N_850,N_206,N_228);
and U851 (N_851,N_373,N_247);
or U852 (N_852,N_466,N_43);
nand U853 (N_853,N_73,N_366);
xnor U854 (N_854,N_441,N_3);
xor U855 (N_855,N_41,N_213);
xnor U856 (N_856,N_281,N_394);
nor U857 (N_857,N_47,N_55);
nor U858 (N_858,N_133,N_391);
xor U859 (N_859,N_283,N_204);
nand U860 (N_860,N_184,N_33);
xnor U861 (N_861,N_442,N_338);
nand U862 (N_862,N_86,N_147);
nor U863 (N_863,N_82,N_67);
and U864 (N_864,N_477,N_362);
nor U865 (N_865,N_419,N_171);
xnor U866 (N_866,N_398,N_117);
nor U867 (N_867,N_309,N_378);
and U868 (N_868,N_352,N_96);
nor U869 (N_869,N_191,N_148);
and U870 (N_870,N_410,N_472);
or U871 (N_871,N_281,N_267);
and U872 (N_872,N_428,N_448);
nor U873 (N_873,N_43,N_247);
nor U874 (N_874,N_236,N_22);
nand U875 (N_875,N_404,N_357);
xnor U876 (N_876,N_131,N_277);
and U877 (N_877,N_14,N_422);
nand U878 (N_878,N_340,N_32);
and U879 (N_879,N_479,N_378);
nand U880 (N_880,N_149,N_359);
and U881 (N_881,N_209,N_240);
and U882 (N_882,N_109,N_237);
nor U883 (N_883,N_45,N_300);
or U884 (N_884,N_105,N_123);
nand U885 (N_885,N_456,N_220);
and U886 (N_886,N_224,N_36);
xor U887 (N_887,N_121,N_129);
nor U888 (N_888,N_222,N_481);
xnor U889 (N_889,N_182,N_412);
nor U890 (N_890,N_294,N_414);
xnor U891 (N_891,N_163,N_453);
and U892 (N_892,N_60,N_312);
or U893 (N_893,N_142,N_340);
or U894 (N_894,N_50,N_342);
and U895 (N_895,N_473,N_203);
and U896 (N_896,N_491,N_461);
xnor U897 (N_897,N_315,N_433);
or U898 (N_898,N_91,N_304);
or U899 (N_899,N_10,N_162);
or U900 (N_900,N_484,N_434);
and U901 (N_901,N_461,N_307);
nor U902 (N_902,N_349,N_63);
or U903 (N_903,N_288,N_289);
nand U904 (N_904,N_285,N_227);
xnor U905 (N_905,N_343,N_171);
and U906 (N_906,N_158,N_195);
nand U907 (N_907,N_27,N_28);
nor U908 (N_908,N_424,N_434);
nand U909 (N_909,N_406,N_173);
and U910 (N_910,N_449,N_461);
nand U911 (N_911,N_361,N_75);
nand U912 (N_912,N_386,N_259);
or U913 (N_913,N_402,N_389);
xnor U914 (N_914,N_37,N_408);
nand U915 (N_915,N_282,N_68);
nand U916 (N_916,N_436,N_128);
xor U917 (N_917,N_44,N_443);
nand U918 (N_918,N_156,N_197);
nand U919 (N_919,N_402,N_464);
xnor U920 (N_920,N_256,N_25);
nor U921 (N_921,N_429,N_31);
xnor U922 (N_922,N_164,N_484);
xnor U923 (N_923,N_49,N_354);
nor U924 (N_924,N_180,N_359);
and U925 (N_925,N_179,N_385);
nand U926 (N_926,N_435,N_449);
nor U927 (N_927,N_128,N_206);
nor U928 (N_928,N_285,N_257);
or U929 (N_929,N_347,N_431);
xnor U930 (N_930,N_499,N_282);
xnor U931 (N_931,N_249,N_397);
nand U932 (N_932,N_322,N_76);
xnor U933 (N_933,N_372,N_8);
and U934 (N_934,N_86,N_143);
and U935 (N_935,N_407,N_38);
and U936 (N_936,N_44,N_60);
nor U937 (N_937,N_444,N_455);
nand U938 (N_938,N_333,N_154);
nor U939 (N_939,N_469,N_433);
and U940 (N_940,N_431,N_477);
nor U941 (N_941,N_403,N_148);
or U942 (N_942,N_287,N_161);
and U943 (N_943,N_55,N_135);
xnor U944 (N_944,N_122,N_57);
or U945 (N_945,N_391,N_82);
nor U946 (N_946,N_238,N_294);
and U947 (N_947,N_445,N_281);
or U948 (N_948,N_445,N_263);
and U949 (N_949,N_264,N_306);
nor U950 (N_950,N_38,N_1);
or U951 (N_951,N_451,N_64);
nor U952 (N_952,N_13,N_230);
xnor U953 (N_953,N_115,N_403);
xor U954 (N_954,N_348,N_21);
and U955 (N_955,N_306,N_362);
and U956 (N_956,N_256,N_453);
nand U957 (N_957,N_21,N_313);
nand U958 (N_958,N_126,N_164);
nor U959 (N_959,N_48,N_440);
nand U960 (N_960,N_497,N_81);
xnor U961 (N_961,N_317,N_70);
xnor U962 (N_962,N_245,N_329);
nand U963 (N_963,N_20,N_370);
and U964 (N_964,N_310,N_371);
xnor U965 (N_965,N_92,N_406);
or U966 (N_966,N_397,N_44);
xor U967 (N_967,N_431,N_437);
or U968 (N_968,N_440,N_406);
or U969 (N_969,N_355,N_128);
xnor U970 (N_970,N_467,N_154);
nand U971 (N_971,N_218,N_3);
and U972 (N_972,N_393,N_407);
and U973 (N_973,N_436,N_340);
nor U974 (N_974,N_316,N_125);
nand U975 (N_975,N_52,N_334);
nand U976 (N_976,N_291,N_44);
or U977 (N_977,N_231,N_77);
nor U978 (N_978,N_146,N_3);
nor U979 (N_979,N_406,N_318);
or U980 (N_980,N_386,N_1);
xor U981 (N_981,N_364,N_13);
and U982 (N_982,N_21,N_440);
xnor U983 (N_983,N_344,N_140);
or U984 (N_984,N_8,N_315);
and U985 (N_985,N_359,N_240);
and U986 (N_986,N_272,N_414);
or U987 (N_987,N_256,N_378);
nand U988 (N_988,N_220,N_171);
and U989 (N_989,N_41,N_77);
or U990 (N_990,N_230,N_411);
nand U991 (N_991,N_251,N_178);
and U992 (N_992,N_133,N_428);
xor U993 (N_993,N_492,N_195);
nand U994 (N_994,N_152,N_381);
and U995 (N_995,N_69,N_404);
nor U996 (N_996,N_106,N_176);
and U997 (N_997,N_12,N_462);
xor U998 (N_998,N_307,N_304);
and U999 (N_999,N_10,N_106);
or U1000 (N_1000,N_928,N_975);
nor U1001 (N_1001,N_702,N_534);
nand U1002 (N_1002,N_869,N_575);
and U1003 (N_1003,N_859,N_662);
nor U1004 (N_1004,N_592,N_586);
nor U1005 (N_1005,N_627,N_503);
xnor U1006 (N_1006,N_800,N_915);
or U1007 (N_1007,N_533,N_753);
or U1008 (N_1008,N_687,N_861);
nand U1009 (N_1009,N_585,N_581);
nand U1010 (N_1010,N_544,N_748);
nand U1011 (N_1011,N_628,N_953);
nand U1012 (N_1012,N_538,N_736);
or U1013 (N_1013,N_689,N_738);
and U1014 (N_1014,N_996,N_770);
xnor U1015 (N_1015,N_910,N_519);
xnor U1016 (N_1016,N_542,N_630);
or U1017 (N_1017,N_709,N_973);
nand U1018 (N_1018,N_725,N_768);
nand U1019 (N_1019,N_781,N_918);
and U1020 (N_1020,N_956,N_909);
or U1021 (N_1021,N_563,N_941);
nand U1022 (N_1022,N_512,N_990);
and U1023 (N_1023,N_500,N_774);
nor U1024 (N_1024,N_857,N_751);
and U1025 (N_1025,N_670,N_693);
nand U1026 (N_1026,N_742,N_783);
or U1027 (N_1027,N_819,N_714);
xnor U1028 (N_1028,N_710,N_816);
nand U1029 (N_1029,N_858,N_605);
and U1030 (N_1030,N_808,N_949);
xnor U1031 (N_1031,N_588,N_691);
nand U1032 (N_1032,N_527,N_947);
nand U1033 (N_1033,N_663,N_815);
xnor U1034 (N_1034,N_986,N_580);
nor U1035 (N_1035,N_578,N_922);
nor U1036 (N_1036,N_923,N_607);
xor U1037 (N_1037,N_591,N_963);
and U1038 (N_1038,N_719,N_900);
nor U1039 (N_1039,N_878,N_549);
xor U1040 (N_1040,N_883,N_690);
and U1041 (N_1041,N_934,N_658);
and U1042 (N_1042,N_638,N_769);
and U1043 (N_1043,N_631,N_896);
or U1044 (N_1044,N_801,N_921);
or U1045 (N_1045,N_643,N_571);
or U1046 (N_1046,N_672,N_969);
nor U1047 (N_1047,N_757,N_884);
or U1048 (N_1048,N_699,N_582);
nand U1049 (N_1049,N_705,N_706);
nor U1050 (N_1050,N_860,N_741);
nor U1051 (N_1051,N_756,N_532);
and U1052 (N_1052,N_752,N_807);
nand U1053 (N_1053,N_961,N_895);
or U1054 (N_1054,N_782,N_565);
nor U1055 (N_1055,N_708,N_914);
nand U1056 (N_1056,N_601,N_676);
nor U1057 (N_1057,N_526,N_573);
xnor U1058 (N_1058,N_604,N_556);
or U1059 (N_1059,N_991,N_642);
nand U1060 (N_1060,N_911,N_727);
or U1061 (N_1061,N_987,N_570);
nand U1062 (N_1062,N_576,N_822);
and U1063 (N_1063,N_614,N_793);
and U1064 (N_1064,N_721,N_632);
nor U1065 (N_1065,N_537,N_868);
nand U1066 (N_1066,N_660,N_810);
xor U1067 (N_1067,N_718,N_787);
nor U1068 (N_1068,N_707,N_794);
and U1069 (N_1069,N_515,N_776);
nor U1070 (N_1070,N_907,N_558);
xor U1071 (N_1071,N_671,N_650);
or U1072 (N_1072,N_729,N_885);
or U1073 (N_1073,N_716,N_624);
or U1074 (N_1074,N_698,N_731);
nand U1075 (N_1075,N_572,N_964);
nand U1076 (N_1076,N_970,N_775);
and U1077 (N_1077,N_971,N_593);
or U1078 (N_1078,N_539,N_695);
and U1079 (N_1079,N_674,N_746);
or U1080 (N_1080,N_880,N_636);
nand U1081 (N_1081,N_951,N_613);
or U1082 (N_1082,N_639,N_750);
nand U1083 (N_1083,N_616,N_891);
nor U1084 (N_1084,N_762,N_546);
nand U1085 (N_1085,N_802,N_826);
xnor U1086 (N_1086,N_930,N_755);
and U1087 (N_1087,N_747,N_608);
and U1088 (N_1088,N_579,N_720);
nor U1089 (N_1089,N_870,N_893);
xnor U1090 (N_1090,N_505,N_871);
xor U1091 (N_1091,N_559,N_897);
xnor U1092 (N_1092,N_550,N_506);
xnor U1093 (N_1093,N_933,N_817);
and U1094 (N_1094,N_540,N_844);
nor U1095 (N_1095,N_739,N_993);
xnor U1096 (N_1096,N_865,N_645);
nor U1097 (N_1097,N_637,N_812);
nor U1098 (N_1098,N_851,N_843);
nor U1099 (N_1099,N_945,N_959);
nor U1100 (N_1100,N_668,N_879);
xnor U1101 (N_1101,N_875,N_978);
nor U1102 (N_1102,N_543,N_912);
nor U1103 (N_1103,N_984,N_764);
xor U1104 (N_1104,N_678,N_696);
and U1105 (N_1105,N_590,N_566);
xnor U1106 (N_1106,N_905,N_979);
nor U1107 (N_1107,N_866,N_656);
nand U1108 (N_1108,N_595,N_618);
nand U1109 (N_1109,N_514,N_925);
and U1110 (N_1110,N_771,N_846);
or U1111 (N_1111,N_936,N_659);
nand U1112 (N_1112,N_856,N_823);
nor U1113 (N_1113,N_838,N_640);
and U1114 (N_1114,N_862,N_745);
and U1115 (N_1115,N_943,N_908);
nand U1116 (N_1116,N_655,N_902);
and U1117 (N_1117,N_913,N_901);
nand U1118 (N_1118,N_615,N_799);
nand U1119 (N_1119,N_806,N_597);
nor U1120 (N_1120,N_726,N_818);
nand U1121 (N_1121,N_744,N_966);
nor U1122 (N_1122,N_648,N_832);
nor U1123 (N_1123,N_686,N_560);
nand U1124 (N_1124,N_621,N_767);
or U1125 (N_1125,N_958,N_797);
and U1126 (N_1126,N_661,N_829);
nand U1127 (N_1127,N_513,N_634);
nand U1128 (N_1128,N_939,N_723);
and U1129 (N_1129,N_531,N_647);
and U1130 (N_1130,N_536,N_853);
nor U1131 (N_1131,N_619,N_825);
xor U1132 (N_1132,N_623,N_522);
xor U1133 (N_1133,N_836,N_955);
nor U1134 (N_1134,N_541,N_790);
nor U1135 (N_1135,N_960,N_665);
nand U1136 (N_1136,N_803,N_840);
nor U1137 (N_1137,N_681,N_873);
or U1138 (N_1138,N_610,N_917);
xnor U1139 (N_1139,N_552,N_938);
or U1140 (N_1140,N_511,N_679);
nand U1141 (N_1141,N_555,N_694);
or U1142 (N_1142,N_811,N_730);
nor U1143 (N_1143,N_927,N_646);
xnor U1144 (N_1144,N_667,N_942);
and U1145 (N_1145,N_703,N_952);
nor U1146 (N_1146,N_983,N_521);
nor U1147 (N_1147,N_995,N_564);
nand U1148 (N_1148,N_666,N_772);
xor U1149 (N_1149,N_965,N_898);
or U1150 (N_1150,N_805,N_830);
and U1151 (N_1151,N_673,N_664);
xnor U1152 (N_1152,N_598,N_889);
or U1153 (N_1153,N_849,N_734);
and U1154 (N_1154,N_735,N_904);
nand U1155 (N_1155,N_848,N_976);
nand U1156 (N_1156,N_946,N_795);
nand U1157 (N_1157,N_626,N_528);
nor U1158 (N_1158,N_997,N_937);
xor U1159 (N_1159,N_692,N_791);
nand U1160 (N_1160,N_989,N_599);
nand U1161 (N_1161,N_924,N_688);
nand U1162 (N_1162,N_920,N_777);
xnor U1163 (N_1163,N_728,N_711);
xor U1164 (N_1164,N_675,N_557);
nand U1165 (N_1165,N_821,N_715);
xnor U1166 (N_1166,N_874,N_722);
nor U1167 (N_1167,N_929,N_653);
xnor U1168 (N_1168,N_523,N_881);
nand U1169 (N_1169,N_831,N_654);
xor U1170 (N_1170,N_568,N_888);
nand U1171 (N_1171,N_785,N_784);
or U1172 (N_1172,N_834,N_733);
nor U1173 (N_1173,N_780,N_779);
and U1174 (N_1174,N_839,N_548);
or U1175 (N_1175,N_743,N_847);
xor U1176 (N_1176,N_510,N_789);
and U1177 (N_1177,N_809,N_890);
nor U1178 (N_1178,N_887,N_824);
or U1179 (N_1179,N_957,N_697);
or U1180 (N_1180,N_855,N_649);
xor U1181 (N_1181,N_886,N_758);
or U1182 (N_1182,N_931,N_919);
nand U1183 (N_1183,N_798,N_792);
nand U1184 (N_1184,N_583,N_551);
and U1185 (N_1185,N_863,N_517);
nand U1186 (N_1186,N_545,N_788);
xnor U1187 (N_1187,N_737,N_606);
xor U1188 (N_1188,N_704,N_754);
nand U1189 (N_1189,N_916,N_980);
nand U1190 (N_1190,N_684,N_981);
nand U1191 (N_1191,N_948,N_828);
nor U1192 (N_1192,N_520,N_852);
xor U1193 (N_1193,N_877,N_972);
xnor U1194 (N_1194,N_504,N_932);
and U1195 (N_1195,N_600,N_713);
or U1196 (N_1196,N_562,N_760);
xor U1197 (N_1197,N_633,N_587);
xor U1198 (N_1198,N_589,N_535);
and U1199 (N_1199,N_561,N_827);
nor U1200 (N_1200,N_892,N_651);
nand U1201 (N_1201,N_501,N_554);
nor U1202 (N_1202,N_529,N_509);
xor U1203 (N_1203,N_525,N_954);
or U1204 (N_1204,N_837,N_569);
and U1205 (N_1205,N_611,N_603);
or U1206 (N_1206,N_724,N_872);
and U1207 (N_1207,N_982,N_749);
nor U1208 (N_1208,N_712,N_967);
nand U1209 (N_1209,N_962,N_899);
nand U1210 (N_1210,N_577,N_629);
or U1211 (N_1211,N_974,N_502);
or U1212 (N_1212,N_804,N_524);
or U1213 (N_1213,N_507,N_682);
nand U1214 (N_1214,N_820,N_657);
xnor U1215 (N_1215,N_635,N_850);
xnor U1216 (N_1216,N_814,N_567);
nand U1217 (N_1217,N_584,N_622);
and U1218 (N_1218,N_845,N_683);
and U1219 (N_1219,N_574,N_669);
and U1220 (N_1220,N_841,N_701);
nand U1221 (N_1221,N_944,N_763);
nand U1222 (N_1222,N_761,N_903);
and U1223 (N_1223,N_732,N_894);
or U1224 (N_1224,N_620,N_765);
nor U1225 (N_1225,N_596,N_652);
and U1226 (N_1226,N_547,N_786);
nand U1227 (N_1227,N_935,N_602);
nor U1228 (N_1228,N_625,N_977);
xnor U1229 (N_1229,N_641,N_876);
xor U1230 (N_1230,N_685,N_842);
nor U1231 (N_1231,N_609,N_700);
or U1232 (N_1232,N_833,N_612);
xor U1233 (N_1233,N_988,N_867);
xnor U1234 (N_1234,N_516,N_677);
nand U1235 (N_1235,N_773,N_994);
or U1236 (N_1236,N_882,N_926);
or U1237 (N_1237,N_518,N_508);
nor U1238 (N_1238,N_680,N_985);
nor U1239 (N_1239,N_940,N_950);
nand U1240 (N_1240,N_813,N_854);
and U1241 (N_1241,N_778,N_992);
nor U1242 (N_1242,N_530,N_594);
nand U1243 (N_1243,N_766,N_998);
and U1244 (N_1244,N_553,N_644);
nand U1245 (N_1245,N_617,N_864);
nor U1246 (N_1246,N_835,N_796);
or U1247 (N_1247,N_999,N_740);
or U1248 (N_1248,N_968,N_717);
or U1249 (N_1249,N_906,N_759);
or U1250 (N_1250,N_829,N_613);
xor U1251 (N_1251,N_826,N_759);
nand U1252 (N_1252,N_854,N_591);
and U1253 (N_1253,N_600,N_740);
nor U1254 (N_1254,N_813,N_739);
nor U1255 (N_1255,N_915,N_532);
nand U1256 (N_1256,N_595,N_519);
or U1257 (N_1257,N_542,N_718);
xnor U1258 (N_1258,N_772,N_760);
and U1259 (N_1259,N_962,N_846);
xor U1260 (N_1260,N_503,N_900);
or U1261 (N_1261,N_597,N_922);
nor U1262 (N_1262,N_579,N_840);
nor U1263 (N_1263,N_984,N_688);
nand U1264 (N_1264,N_907,N_557);
xnor U1265 (N_1265,N_595,N_746);
or U1266 (N_1266,N_518,N_812);
nor U1267 (N_1267,N_501,N_953);
or U1268 (N_1268,N_665,N_577);
xor U1269 (N_1269,N_712,N_702);
xor U1270 (N_1270,N_545,N_783);
xor U1271 (N_1271,N_860,N_935);
nor U1272 (N_1272,N_806,N_566);
nor U1273 (N_1273,N_961,N_500);
xnor U1274 (N_1274,N_956,N_503);
and U1275 (N_1275,N_845,N_725);
or U1276 (N_1276,N_730,N_867);
xnor U1277 (N_1277,N_616,N_868);
nand U1278 (N_1278,N_906,N_965);
xor U1279 (N_1279,N_780,N_574);
nand U1280 (N_1280,N_613,N_812);
nor U1281 (N_1281,N_951,N_622);
or U1282 (N_1282,N_754,N_568);
and U1283 (N_1283,N_973,N_923);
xor U1284 (N_1284,N_830,N_602);
or U1285 (N_1285,N_540,N_535);
nor U1286 (N_1286,N_619,N_870);
nand U1287 (N_1287,N_815,N_973);
or U1288 (N_1288,N_914,N_797);
or U1289 (N_1289,N_751,N_987);
xnor U1290 (N_1290,N_560,N_742);
nor U1291 (N_1291,N_570,N_612);
or U1292 (N_1292,N_897,N_738);
and U1293 (N_1293,N_905,N_807);
xnor U1294 (N_1294,N_535,N_513);
xnor U1295 (N_1295,N_864,N_553);
and U1296 (N_1296,N_653,N_594);
nand U1297 (N_1297,N_871,N_869);
xnor U1298 (N_1298,N_571,N_500);
or U1299 (N_1299,N_550,N_788);
nand U1300 (N_1300,N_973,N_512);
xnor U1301 (N_1301,N_856,N_869);
nor U1302 (N_1302,N_979,N_711);
or U1303 (N_1303,N_983,N_869);
xnor U1304 (N_1304,N_825,N_706);
nor U1305 (N_1305,N_852,N_655);
or U1306 (N_1306,N_550,N_778);
nor U1307 (N_1307,N_986,N_644);
xor U1308 (N_1308,N_702,N_627);
xnor U1309 (N_1309,N_951,N_549);
or U1310 (N_1310,N_510,N_728);
or U1311 (N_1311,N_520,N_920);
and U1312 (N_1312,N_992,N_688);
or U1313 (N_1313,N_835,N_929);
nand U1314 (N_1314,N_672,N_988);
nor U1315 (N_1315,N_674,N_894);
xnor U1316 (N_1316,N_914,N_858);
xnor U1317 (N_1317,N_616,N_772);
and U1318 (N_1318,N_742,N_872);
nand U1319 (N_1319,N_602,N_909);
and U1320 (N_1320,N_700,N_848);
nor U1321 (N_1321,N_952,N_589);
nand U1322 (N_1322,N_666,N_575);
and U1323 (N_1323,N_922,N_975);
or U1324 (N_1324,N_990,N_917);
xnor U1325 (N_1325,N_796,N_816);
nor U1326 (N_1326,N_857,N_735);
xnor U1327 (N_1327,N_972,N_816);
xnor U1328 (N_1328,N_764,N_926);
and U1329 (N_1329,N_679,N_879);
xnor U1330 (N_1330,N_607,N_804);
xnor U1331 (N_1331,N_901,N_591);
or U1332 (N_1332,N_540,N_807);
xor U1333 (N_1333,N_957,N_608);
and U1334 (N_1334,N_758,N_625);
xor U1335 (N_1335,N_702,N_715);
nor U1336 (N_1336,N_718,N_529);
or U1337 (N_1337,N_660,N_695);
nor U1338 (N_1338,N_820,N_609);
or U1339 (N_1339,N_986,N_586);
and U1340 (N_1340,N_560,N_885);
and U1341 (N_1341,N_716,N_833);
nand U1342 (N_1342,N_707,N_604);
and U1343 (N_1343,N_599,N_870);
xor U1344 (N_1344,N_661,N_536);
and U1345 (N_1345,N_867,N_778);
or U1346 (N_1346,N_766,N_993);
or U1347 (N_1347,N_590,N_717);
and U1348 (N_1348,N_544,N_729);
and U1349 (N_1349,N_711,N_947);
and U1350 (N_1350,N_838,N_780);
or U1351 (N_1351,N_893,N_972);
nor U1352 (N_1352,N_603,N_749);
nor U1353 (N_1353,N_864,N_823);
or U1354 (N_1354,N_860,N_989);
nand U1355 (N_1355,N_944,N_929);
and U1356 (N_1356,N_579,N_878);
xor U1357 (N_1357,N_984,N_610);
xnor U1358 (N_1358,N_501,N_741);
xnor U1359 (N_1359,N_767,N_560);
and U1360 (N_1360,N_868,N_656);
and U1361 (N_1361,N_741,N_913);
and U1362 (N_1362,N_898,N_897);
nand U1363 (N_1363,N_757,N_639);
xnor U1364 (N_1364,N_937,N_828);
or U1365 (N_1365,N_509,N_991);
nand U1366 (N_1366,N_590,N_779);
xor U1367 (N_1367,N_509,N_654);
xor U1368 (N_1368,N_526,N_736);
and U1369 (N_1369,N_695,N_533);
xnor U1370 (N_1370,N_963,N_566);
nand U1371 (N_1371,N_504,N_988);
nor U1372 (N_1372,N_941,N_802);
nor U1373 (N_1373,N_938,N_935);
nand U1374 (N_1374,N_680,N_642);
nand U1375 (N_1375,N_929,N_586);
xnor U1376 (N_1376,N_545,N_970);
and U1377 (N_1377,N_985,N_649);
or U1378 (N_1378,N_910,N_506);
or U1379 (N_1379,N_500,N_687);
xor U1380 (N_1380,N_518,N_858);
and U1381 (N_1381,N_863,N_901);
nor U1382 (N_1382,N_723,N_995);
nand U1383 (N_1383,N_912,N_897);
nand U1384 (N_1384,N_657,N_611);
or U1385 (N_1385,N_899,N_765);
or U1386 (N_1386,N_635,N_525);
nand U1387 (N_1387,N_817,N_594);
nand U1388 (N_1388,N_746,N_551);
and U1389 (N_1389,N_647,N_785);
xor U1390 (N_1390,N_986,N_574);
xor U1391 (N_1391,N_861,N_941);
nor U1392 (N_1392,N_655,N_843);
or U1393 (N_1393,N_563,N_928);
or U1394 (N_1394,N_616,N_745);
nand U1395 (N_1395,N_948,N_667);
or U1396 (N_1396,N_528,N_561);
nand U1397 (N_1397,N_991,N_840);
and U1398 (N_1398,N_845,N_865);
xnor U1399 (N_1399,N_875,N_772);
nor U1400 (N_1400,N_583,N_556);
or U1401 (N_1401,N_834,N_656);
nor U1402 (N_1402,N_602,N_635);
nand U1403 (N_1403,N_892,N_582);
or U1404 (N_1404,N_530,N_997);
or U1405 (N_1405,N_518,N_838);
and U1406 (N_1406,N_966,N_864);
xnor U1407 (N_1407,N_911,N_933);
nand U1408 (N_1408,N_942,N_929);
nor U1409 (N_1409,N_552,N_509);
nand U1410 (N_1410,N_949,N_856);
or U1411 (N_1411,N_866,N_677);
nor U1412 (N_1412,N_706,N_668);
nor U1413 (N_1413,N_860,N_638);
or U1414 (N_1414,N_971,N_619);
or U1415 (N_1415,N_931,N_563);
or U1416 (N_1416,N_994,N_720);
xnor U1417 (N_1417,N_757,N_985);
nor U1418 (N_1418,N_563,N_553);
nand U1419 (N_1419,N_726,N_952);
xnor U1420 (N_1420,N_990,N_734);
xnor U1421 (N_1421,N_548,N_767);
nor U1422 (N_1422,N_747,N_552);
and U1423 (N_1423,N_927,N_740);
xor U1424 (N_1424,N_924,N_545);
and U1425 (N_1425,N_580,N_757);
nor U1426 (N_1426,N_604,N_761);
or U1427 (N_1427,N_803,N_533);
nand U1428 (N_1428,N_733,N_663);
and U1429 (N_1429,N_700,N_965);
nand U1430 (N_1430,N_644,N_759);
or U1431 (N_1431,N_907,N_724);
nand U1432 (N_1432,N_797,N_810);
and U1433 (N_1433,N_841,N_600);
and U1434 (N_1434,N_687,N_820);
nor U1435 (N_1435,N_849,N_590);
nand U1436 (N_1436,N_721,N_540);
or U1437 (N_1437,N_930,N_507);
nand U1438 (N_1438,N_503,N_881);
xor U1439 (N_1439,N_680,N_547);
nand U1440 (N_1440,N_763,N_608);
xnor U1441 (N_1441,N_576,N_764);
xnor U1442 (N_1442,N_509,N_857);
nor U1443 (N_1443,N_934,N_947);
nand U1444 (N_1444,N_666,N_992);
and U1445 (N_1445,N_558,N_655);
nand U1446 (N_1446,N_569,N_684);
and U1447 (N_1447,N_813,N_914);
xnor U1448 (N_1448,N_509,N_830);
and U1449 (N_1449,N_572,N_857);
or U1450 (N_1450,N_784,N_517);
and U1451 (N_1451,N_577,N_984);
nand U1452 (N_1452,N_650,N_684);
and U1453 (N_1453,N_508,N_770);
xor U1454 (N_1454,N_774,N_765);
nand U1455 (N_1455,N_979,N_690);
and U1456 (N_1456,N_885,N_522);
or U1457 (N_1457,N_509,N_879);
or U1458 (N_1458,N_627,N_933);
or U1459 (N_1459,N_821,N_626);
or U1460 (N_1460,N_553,N_622);
nand U1461 (N_1461,N_832,N_800);
nand U1462 (N_1462,N_707,N_891);
and U1463 (N_1463,N_740,N_846);
nor U1464 (N_1464,N_832,N_679);
nor U1465 (N_1465,N_574,N_702);
or U1466 (N_1466,N_630,N_769);
or U1467 (N_1467,N_723,N_542);
nor U1468 (N_1468,N_953,N_580);
nor U1469 (N_1469,N_787,N_744);
xnor U1470 (N_1470,N_954,N_702);
xnor U1471 (N_1471,N_996,N_629);
nor U1472 (N_1472,N_811,N_814);
nor U1473 (N_1473,N_596,N_751);
xnor U1474 (N_1474,N_989,N_773);
nor U1475 (N_1475,N_828,N_611);
and U1476 (N_1476,N_952,N_752);
nand U1477 (N_1477,N_854,N_902);
xor U1478 (N_1478,N_800,N_568);
nand U1479 (N_1479,N_985,N_660);
or U1480 (N_1480,N_560,N_709);
or U1481 (N_1481,N_662,N_773);
nand U1482 (N_1482,N_753,N_693);
xor U1483 (N_1483,N_811,N_596);
and U1484 (N_1484,N_705,N_732);
xor U1485 (N_1485,N_880,N_802);
nor U1486 (N_1486,N_867,N_678);
or U1487 (N_1487,N_700,N_804);
xnor U1488 (N_1488,N_682,N_841);
xor U1489 (N_1489,N_657,N_801);
and U1490 (N_1490,N_507,N_863);
nor U1491 (N_1491,N_552,N_961);
nor U1492 (N_1492,N_518,N_826);
and U1493 (N_1493,N_937,N_762);
or U1494 (N_1494,N_662,N_996);
nand U1495 (N_1495,N_703,N_863);
nand U1496 (N_1496,N_798,N_718);
nand U1497 (N_1497,N_882,N_774);
nand U1498 (N_1498,N_847,N_657);
nand U1499 (N_1499,N_738,N_891);
xnor U1500 (N_1500,N_1267,N_1411);
and U1501 (N_1501,N_1038,N_1288);
or U1502 (N_1502,N_1496,N_1010);
nor U1503 (N_1503,N_1189,N_1112);
or U1504 (N_1504,N_1223,N_1212);
xor U1505 (N_1505,N_1269,N_1428);
xor U1506 (N_1506,N_1181,N_1484);
or U1507 (N_1507,N_1215,N_1356);
nor U1508 (N_1508,N_1338,N_1433);
and U1509 (N_1509,N_1253,N_1244);
nor U1510 (N_1510,N_1236,N_1095);
xnor U1511 (N_1511,N_1418,N_1254);
nor U1512 (N_1512,N_1314,N_1372);
nand U1513 (N_1513,N_1022,N_1376);
xnor U1514 (N_1514,N_1284,N_1447);
nor U1515 (N_1515,N_1238,N_1343);
xor U1516 (N_1516,N_1091,N_1319);
xor U1517 (N_1517,N_1102,N_1043);
and U1518 (N_1518,N_1193,N_1082);
nor U1519 (N_1519,N_1436,N_1390);
and U1520 (N_1520,N_1282,N_1074);
nand U1521 (N_1521,N_1161,N_1008);
nand U1522 (N_1522,N_1046,N_1339);
xnor U1523 (N_1523,N_1031,N_1086);
nor U1524 (N_1524,N_1332,N_1287);
nor U1525 (N_1525,N_1029,N_1308);
xor U1526 (N_1526,N_1385,N_1173);
or U1527 (N_1527,N_1266,N_1312);
or U1528 (N_1528,N_1408,N_1256);
nor U1529 (N_1529,N_1291,N_1130);
or U1530 (N_1530,N_1456,N_1042);
and U1531 (N_1531,N_1018,N_1076);
xnor U1532 (N_1532,N_1063,N_1220);
xor U1533 (N_1533,N_1019,N_1242);
or U1534 (N_1534,N_1011,N_1151);
or U1535 (N_1535,N_1003,N_1213);
nand U1536 (N_1536,N_1283,N_1286);
or U1537 (N_1537,N_1106,N_1261);
xnor U1538 (N_1538,N_1405,N_1497);
nand U1539 (N_1539,N_1157,N_1237);
and U1540 (N_1540,N_1363,N_1264);
nor U1541 (N_1541,N_1426,N_1085);
or U1542 (N_1542,N_1443,N_1285);
and U1543 (N_1543,N_1201,N_1369);
or U1544 (N_1544,N_1446,N_1167);
and U1545 (N_1545,N_1122,N_1057);
nand U1546 (N_1546,N_1333,N_1227);
and U1547 (N_1547,N_1410,N_1134);
xnor U1548 (N_1548,N_1358,N_1054);
and U1549 (N_1549,N_1421,N_1050);
and U1550 (N_1550,N_1216,N_1274);
nor U1551 (N_1551,N_1462,N_1171);
and U1552 (N_1552,N_1473,N_1103);
nor U1553 (N_1553,N_1056,N_1163);
nor U1554 (N_1554,N_1077,N_1360);
and U1555 (N_1555,N_1115,N_1118);
and U1556 (N_1556,N_1222,N_1335);
xor U1557 (N_1557,N_1487,N_1359);
and U1558 (N_1558,N_1302,N_1326);
or U1559 (N_1559,N_1420,N_1039);
nand U1560 (N_1560,N_1384,N_1402);
xnor U1561 (N_1561,N_1133,N_1191);
nand U1562 (N_1562,N_1355,N_1431);
and U1563 (N_1563,N_1178,N_1255);
and U1564 (N_1564,N_1015,N_1025);
nand U1565 (N_1565,N_1272,N_1262);
nor U1566 (N_1566,N_1455,N_1467);
and U1567 (N_1567,N_1107,N_1217);
nand U1568 (N_1568,N_1305,N_1395);
nor U1569 (N_1569,N_1224,N_1105);
nand U1570 (N_1570,N_1318,N_1186);
and U1571 (N_1571,N_1126,N_1035);
nand U1572 (N_1572,N_1407,N_1012);
xnor U1573 (N_1573,N_1329,N_1202);
xor U1574 (N_1574,N_1069,N_1048);
or U1575 (N_1575,N_1239,N_1422);
and U1576 (N_1576,N_1474,N_1044);
xor U1577 (N_1577,N_1009,N_1014);
or U1578 (N_1578,N_1463,N_1321);
and U1579 (N_1579,N_1245,N_1336);
and U1580 (N_1580,N_1393,N_1158);
or U1581 (N_1581,N_1001,N_1445);
xor U1582 (N_1582,N_1041,N_1226);
xnor U1583 (N_1583,N_1243,N_1209);
xor U1584 (N_1584,N_1442,N_1415);
nor U1585 (N_1585,N_1028,N_1437);
nor U1586 (N_1586,N_1240,N_1362);
xor U1587 (N_1587,N_1067,N_1300);
nor U1588 (N_1588,N_1294,N_1465);
xor U1589 (N_1589,N_1229,N_1049);
nor U1590 (N_1590,N_1346,N_1398);
and U1591 (N_1591,N_1386,N_1169);
or U1592 (N_1592,N_1155,N_1290);
nor U1593 (N_1593,N_1109,N_1352);
nor U1594 (N_1594,N_1354,N_1108);
nor U1595 (N_1595,N_1208,N_1205);
and U1596 (N_1596,N_1366,N_1160);
nand U1597 (N_1597,N_1148,N_1486);
nand U1598 (N_1598,N_1174,N_1053);
nor U1599 (N_1599,N_1060,N_1068);
xnor U1600 (N_1600,N_1016,N_1476);
or U1601 (N_1601,N_1460,N_1493);
and U1602 (N_1602,N_1198,N_1006);
nor U1603 (N_1603,N_1152,N_1021);
or U1604 (N_1604,N_1268,N_1187);
nor U1605 (N_1605,N_1111,N_1197);
nor U1606 (N_1606,N_1051,N_1119);
and U1607 (N_1607,N_1124,N_1150);
nor U1608 (N_1608,N_1489,N_1438);
or U1609 (N_1609,N_1005,N_1383);
xor U1610 (N_1610,N_1481,N_1092);
and U1611 (N_1611,N_1013,N_1277);
or U1612 (N_1612,N_1417,N_1088);
and U1613 (N_1613,N_1147,N_1221);
nor U1614 (N_1614,N_1032,N_1328);
or U1615 (N_1615,N_1348,N_1425);
xor U1616 (N_1616,N_1342,N_1062);
xnor U1617 (N_1617,N_1026,N_1081);
and U1618 (N_1618,N_1172,N_1475);
nor U1619 (N_1619,N_1128,N_1298);
nand U1620 (N_1620,N_1164,N_1113);
nor U1621 (N_1621,N_1457,N_1144);
nand U1622 (N_1622,N_1492,N_1353);
and U1623 (N_1623,N_1203,N_1278);
nor U1624 (N_1624,N_1034,N_1233);
and U1625 (N_1625,N_1414,N_1271);
nor U1626 (N_1626,N_1132,N_1146);
xnor U1627 (N_1627,N_1154,N_1066);
nand U1628 (N_1628,N_1194,N_1490);
or U1629 (N_1629,N_1120,N_1380);
nor U1630 (N_1630,N_1488,N_1270);
nor U1631 (N_1631,N_1024,N_1000);
nor U1632 (N_1632,N_1072,N_1337);
nand U1633 (N_1633,N_1450,N_1378);
or U1634 (N_1634,N_1491,N_1280);
nor U1635 (N_1635,N_1257,N_1177);
nand U1636 (N_1636,N_1180,N_1104);
xor U1637 (N_1637,N_1002,N_1145);
nand U1638 (N_1638,N_1131,N_1089);
nand U1639 (N_1639,N_1235,N_1419);
and U1640 (N_1640,N_1023,N_1045);
nor U1641 (N_1641,N_1030,N_1248);
or U1642 (N_1642,N_1073,N_1070);
or U1643 (N_1643,N_1211,N_1192);
or U1644 (N_1644,N_1219,N_1303);
nand U1645 (N_1645,N_1281,N_1061);
and U1646 (N_1646,N_1409,N_1260);
nor U1647 (N_1647,N_1483,N_1495);
xnor U1648 (N_1648,N_1293,N_1470);
xnor U1649 (N_1649,N_1389,N_1176);
xnor U1650 (N_1650,N_1004,N_1199);
or U1651 (N_1651,N_1365,N_1065);
or U1652 (N_1652,N_1183,N_1079);
xnor U1653 (N_1653,N_1184,N_1188);
xor U1654 (N_1654,N_1439,N_1114);
or U1655 (N_1655,N_1448,N_1454);
and U1656 (N_1656,N_1100,N_1400);
and U1657 (N_1657,N_1230,N_1361);
and U1658 (N_1658,N_1432,N_1382);
nand U1659 (N_1659,N_1391,N_1273);
or U1660 (N_1660,N_1416,N_1033);
nor U1661 (N_1661,N_1047,N_1471);
nor U1662 (N_1662,N_1207,N_1196);
and U1663 (N_1663,N_1121,N_1017);
nand U1664 (N_1664,N_1096,N_1175);
or U1665 (N_1665,N_1251,N_1055);
xnor U1666 (N_1666,N_1345,N_1330);
xor U1667 (N_1667,N_1064,N_1093);
nor U1668 (N_1668,N_1214,N_1451);
xnor U1669 (N_1669,N_1485,N_1137);
nand U1670 (N_1670,N_1040,N_1397);
nor U1671 (N_1671,N_1263,N_1292);
xnor U1672 (N_1672,N_1482,N_1441);
or U1673 (N_1673,N_1480,N_1401);
xor U1674 (N_1674,N_1166,N_1058);
or U1675 (N_1675,N_1138,N_1429);
or U1676 (N_1676,N_1306,N_1206);
and U1677 (N_1677,N_1097,N_1071);
nor U1678 (N_1678,N_1478,N_1427);
and U1679 (N_1679,N_1347,N_1084);
nor U1680 (N_1680,N_1494,N_1379);
and U1681 (N_1681,N_1116,N_1083);
nor U1682 (N_1682,N_1394,N_1052);
and U1683 (N_1683,N_1125,N_1466);
and U1684 (N_1684,N_1170,N_1351);
and U1685 (N_1685,N_1368,N_1204);
and U1686 (N_1686,N_1444,N_1252);
xnor U1687 (N_1687,N_1179,N_1453);
xnor U1688 (N_1688,N_1499,N_1404);
xnor U1689 (N_1689,N_1373,N_1249);
nor U1690 (N_1690,N_1094,N_1344);
and U1691 (N_1691,N_1357,N_1440);
xnor U1692 (N_1692,N_1090,N_1129);
and U1693 (N_1693,N_1258,N_1101);
nor U1694 (N_1694,N_1424,N_1375);
nor U1695 (N_1695,N_1078,N_1110);
nor U1696 (N_1696,N_1316,N_1477);
and U1697 (N_1697,N_1430,N_1231);
or U1698 (N_1698,N_1377,N_1310);
and U1699 (N_1699,N_1200,N_1452);
nor U1700 (N_1700,N_1364,N_1246);
and U1701 (N_1701,N_1479,N_1210);
xor U1702 (N_1702,N_1461,N_1472);
nand U1703 (N_1703,N_1295,N_1317);
nand U1704 (N_1704,N_1127,N_1140);
or U1705 (N_1705,N_1334,N_1315);
or U1706 (N_1706,N_1098,N_1406);
nand U1707 (N_1707,N_1468,N_1322);
xor U1708 (N_1708,N_1396,N_1123);
xnor U1709 (N_1709,N_1371,N_1323);
and U1710 (N_1710,N_1099,N_1182);
or U1711 (N_1711,N_1250,N_1080);
nand U1712 (N_1712,N_1307,N_1301);
and U1713 (N_1713,N_1087,N_1399);
nand U1714 (N_1714,N_1392,N_1225);
nand U1715 (N_1715,N_1218,N_1075);
nand U1716 (N_1716,N_1403,N_1136);
xnor U1717 (N_1717,N_1279,N_1412);
xor U1718 (N_1718,N_1340,N_1434);
and U1719 (N_1719,N_1387,N_1141);
or U1720 (N_1720,N_1143,N_1367);
or U1721 (N_1721,N_1325,N_1027);
nand U1722 (N_1722,N_1275,N_1149);
xor U1723 (N_1723,N_1168,N_1327);
and U1724 (N_1724,N_1374,N_1413);
and U1725 (N_1725,N_1036,N_1142);
xnor U1726 (N_1726,N_1247,N_1388);
nand U1727 (N_1727,N_1153,N_1165);
or U1728 (N_1728,N_1331,N_1304);
nand U1729 (N_1729,N_1349,N_1469);
xor U1730 (N_1730,N_1297,N_1299);
nand U1731 (N_1731,N_1313,N_1435);
nor U1732 (N_1732,N_1162,N_1498);
xnor U1733 (N_1733,N_1296,N_1449);
nor U1734 (N_1734,N_1381,N_1458);
nor U1735 (N_1735,N_1020,N_1309);
nor U1736 (N_1736,N_1324,N_1259);
or U1737 (N_1737,N_1228,N_1289);
and U1738 (N_1738,N_1350,N_1341);
and U1739 (N_1739,N_1464,N_1265);
and U1740 (N_1740,N_1311,N_1117);
xnor U1741 (N_1741,N_1241,N_1037);
nand U1742 (N_1742,N_1423,N_1190);
nand U1743 (N_1743,N_1156,N_1185);
and U1744 (N_1744,N_1370,N_1059);
xnor U1745 (N_1745,N_1320,N_1135);
or U1746 (N_1746,N_1139,N_1234);
nor U1747 (N_1747,N_1195,N_1007);
and U1748 (N_1748,N_1232,N_1276);
or U1749 (N_1749,N_1159,N_1459);
xnor U1750 (N_1750,N_1059,N_1172);
or U1751 (N_1751,N_1307,N_1020);
and U1752 (N_1752,N_1028,N_1464);
nand U1753 (N_1753,N_1249,N_1251);
nor U1754 (N_1754,N_1363,N_1190);
nand U1755 (N_1755,N_1373,N_1123);
xnor U1756 (N_1756,N_1037,N_1417);
or U1757 (N_1757,N_1313,N_1350);
nor U1758 (N_1758,N_1471,N_1145);
or U1759 (N_1759,N_1177,N_1173);
or U1760 (N_1760,N_1402,N_1060);
xnor U1761 (N_1761,N_1364,N_1322);
xnor U1762 (N_1762,N_1245,N_1170);
nand U1763 (N_1763,N_1176,N_1054);
and U1764 (N_1764,N_1273,N_1055);
or U1765 (N_1765,N_1431,N_1016);
xor U1766 (N_1766,N_1198,N_1343);
and U1767 (N_1767,N_1263,N_1347);
nand U1768 (N_1768,N_1380,N_1072);
or U1769 (N_1769,N_1337,N_1046);
or U1770 (N_1770,N_1385,N_1255);
nor U1771 (N_1771,N_1464,N_1004);
nor U1772 (N_1772,N_1154,N_1233);
and U1773 (N_1773,N_1268,N_1152);
xor U1774 (N_1774,N_1338,N_1163);
nor U1775 (N_1775,N_1397,N_1330);
or U1776 (N_1776,N_1421,N_1263);
nand U1777 (N_1777,N_1169,N_1166);
or U1778 (N_1778,N_1112,N_1468);
or U1779 (N_1779,N_1078,N_1322);
and U1780 (N_1780,N_1392,N_1155);
nand U1781 (N_1781,N_1085,N_1436);
nor U1782 (N_1782,N_1319,N_1455);
nand U1783 (N_1783,N_1418,N_1249);
nand U1784 (N_1784,N_1136,N_1057);
and U1785 (N_1785,N_1210,N_1271);
xnor U1786 (N_1786,N_1450,N_1193);
or U1787 (N_1787,N_1097,N_1297);
or U1788 (N_1788,N_1309,N_1140);
or U1789 (N_1789,N_1378,N_1121);
and U1790 (N_1790,N_1040,N_1497);
or U1791 (N_1791,N_1277,N_1381);
or U1792 (N_1792,N_1402,N_1241);
or U1793 (N_1793,N_1462,N_1090);
nand U1794 (N_1794,N_1185,N_1175);
nand U1795 (N_1795,N_1200,N_1250);
xor U1796 (N_1796,N_1369,N_1207);
nand U1797 (N_1797,N_1251,N_1422);
and U1798 (N_1798,N_1020,N_1156);
nand U1799 (N_1799,N_1365,N_1040);
nor U1800 (N_1800,N_1173,N_1122);
nor U1801 (N_1801,N_1261,N_1145);
and U1802 (N_1802,N_1464,N_1351);
nand U1803 (N_1803,N_1160,N_1041);
nand U1804 (N_1804,N_1457,N_1220);
or U1805 (N_1805,N_1303,N_1379);
nor U1806 (N_1806,N_1124,N_1202);
and U1807 (N_1807,N_1361,N_1019);
xor U1808 (N_1808,N_1494,N_1144);
nor U1809 (N_1809,N_1327,N_1129);
xnor U1810 (N_1810,N_1380,N_1044);
xnor U1811 (N_1811,N_1325,N_1343);
and U1812 (N_1812,N_1220,N_1192);
and U1813 (N_1813,N_1476,N_1032);
nor U1814 (N_1814,N_1342,N_1334);
or U1815 (N_1815,N_1161,N_1258);
or U1816 (N_1816,N_1168,N_1247);
nand U1817 (N_1817,N_1233,N_1204);
or U1818 (N_1818,N_1224,N_1278);
and U1819 (N_1819,N_1346,N_1290);
nand U1820 (N_1820,N_1098,N_1298);
nor U1821 (N_1821,N_1249,N_1139);
nand U1822 (N_1822,N_1190,N_1346);
nor U1823 (N_1823,N_1450,N_1417);
nor U1824 (N_1824,N_1280,N_1016);
or U1825 (N_1825,N_1364,N_1245);
xor U1826 (N_1826,N_1449,N_1293);
xor U1827 (N_1827,N_1021,N_1197);
and U1828 (N_1828,N_1115,N_1075);
xor U1829 (N_1829,N_1227,N_1318);
nor U1830 (N_1830,N_1178,N_1470);
xor U1831 (N_1831,N_1266,N_1478);
nor U1832 (N_1832,N_1382,N_1444);
nor U1833 (N_1833,N_1491,N_1099);
or U1834 (N_1834,N_1229,N_1481);
and U1835 (N_1835,N_1336,N_1094);
and U1836 (N_1836,N_1068,N_1400);
or U1837 (N_1837,N_1422,N_1399);
nor U1838 (N_1838,N_1189,N_1323);
xor U1839 (N_1839,N_1419,N_1152);
and U1840 (N_1840,N_1001,N_1119);
and U1841 (N_1841,N_1345,N_1111);
nor U1842 (N_1842,N_1238,N_1316);
nand U1843 (N_1843,N_1301,N_1319);
and U1844 (N_1844,N_1139,N_1141);
nand U1845 (N_1845,N_1343,N_1056);
xnor U1846 (N_1846,N_1201,N_1326);
nand U1847 (N_1847,N_1429,N_1287);
and U1848 (N_1848,N_1407,N_1129);
and U1849 (N_1849,N_1244,N_1067);
nor U1850 (N_1850,N_1357,N_1214);
or U1851 (N_1851,N_1030,N_1015);
nand U1852 (N_1852,N_1389,N_1258);
nor U1853 (N_1853,N_1401,N_1246);
or U1854 (N_1854,N_1001,N_1324);
nor U1855 (N_1855,N_1010,N_1348);
nand U1856 (N_1856,N_1286,N_1144);
nor U1857 (N_1857,N_1165,N_1341);
and U1858 (N_1858,N_1493,N_1300);
nand U1859 (N_1859,N_1237,N_1247);
nor U1860 (N_1860,N_1351,N_1254);
or U1861 (N_1861,N_1169,N_1449);
nand U1862 (N_1862,N_1499,N_1169);
nand U1863 (N_1863,N_1313,N_1431);
or U1864 (N_1864,N_1125,N_1177);
xnor U1865 (N_1865,N_1052,N_1093);
nor U1866 (N_1866,N_1125,N_1397);
nand U1867 (N_1867,N_1374,N_1471);
and U1868 (N_1868,N_1003,N_1033);
nor U1869 (N_1869,N_1194,N_1208);
xnor U1870 (N_1870,N_1144,N_1304);
or U1871 (N_1871,N_1429,N_1458);
or U1872 (N_1872,N_1215,N_1312);
or U1873 (N_1873,N_1313,N_1330);
xnor U1874 (N_1874,N_1067,N_1304);
or U1875 (N_1875,N_1350,N_1416);
nand U1876 (N_1876,N_1266,N_1138);
nor U1877 (N_1877,N_1098,N_1454);
nand U1878 (N_1878,N_1216,N_1452);
nand U1879 (N_1879,N_1206,N_1183);
nand U1880 (N_1880,N_1259,N_1005);
nor U1881 (N_1881,N_1167,N_1213);
xor U1882 (N_1882,N_1337,N_1135);
or U1883 (N_1883,N_1322,N_1262);
xor U1884 (N_1884,N_1361,N_1107);
or U1885 (N_1885,N_1164,N_1294);
or U1886 (N_1886,N_1156,N_1024);
xnor U1887 (N_1887,N_1179,N_1303);
and U1888 (N_1888,N_1335,N_1263);
and U1889 (N_1889,N_1359,N_1375);
and U1890 (N_1890,N_1458,N_1159);
nand U1891 (N_1891,N_1274,N_1054);
xnor U1892 (N_1892,N_1134,N_1120);
and U1893 (N_1893,N_1441,N_1417);
or U1894 (N_1894,N_1495,N_1150);
xor U1895 (N_1895,N_1412,N_1338);
nor U1896 (N_1896,N_1196,N_1100);
or U1897 (N_1897,N_1114,N_1477);
or U1898 (N_1898,N_1362,N_1460);
and U1899 (N_1899,N_1377,N_1194);
or U1900 (N_1900,N_1101,N_1432);
xor U1901 (N_1901,N_1352,N_1191);
xnor U1902 (N_1902,N_1442,N_1473);
or U1903 (N_1903,N_1080,N_1363);
or U1904 (N_1904,N_1148,N_1165);
and U1905 (N_1905,N_1085,N_1475);
and U1906 (N_1906,N_1259,N_1256);
or U1907 (N_1907,N_1184,N_1054);
nor U1908 (N_1908,N_1067,N_1217);
nand U1909 (N_1909,N_1267,N_1429);
and U1910 (N_1910,N_1241,N_1450);
and U1911 (N_1911,N_1071,N_1012);
xor U1912 (N_1912,N_1479,N_1040);
nor U1913 (N_1913,N_1362,N_1432);
or U1914 (N_1914,N_1488,N_1382);
xor U1915 (N_1915,N_1306,N_1208);
or U1916 (N_1916,N_1006,N_1342);
and U1917 (N_1917,N_1383,N_1318);
or U1918 (N_1918,N_1324,N_1450);
xor U1919 (N_1919,N_1425,N_1295);
nand U1920 (N_1920,N_1080,N_1169);
nand U1921 (N_1921,N_1148,N_1331);
and U1922 (N_1922,N_1419,N_1136);
xnor U1923 (N_1923,N_1375,N_1454);
or U1924 (N_1924,N_1052,N_1036);
nor U1925 (N_1925,N_1310,N_1000);
nor U1926 (N_1926,N_1475,N_1203);
xor U1927 (N_1927,N_1276,N_1453);
or U1928 (N_1928,N_1177,N_1269);
nor U1929 (N_1929,N_1111,N_1432);
nand U1930 (N_1930,N_1152,N_1148);
nand U1931 (N_1931,N_1300,N_1128);
and U1932 (N_1932,N_1175,N_1397);
nor U1933 (N_1933,N_1428,N_1493);
xor U1934 (N_1934,N_1338,N_1388);
xor U1935 (N_1935,N_1038,N_1297);
and U1936 (N_1936,N_1313,N_1056);
and U1937 (N_1937,N_1236,N_1311);
nand U1938 (N_1938,N_1313,N_1034);
and U1939 (N_1939,N_1038,N_1458);
nor U1940 (N_1940,N_1243,N_1450);
and U1941 (N_1941,N_1216,N_1053);
and U1942 (N_1942,N_1197,N_1273);
or U1943 (N_1943,N_1452,N_1364);
and U1944 (N_1944,N_1078,N_1437);
nor U1945 (N_1945,N_1157,N_1067);
xnor U1946 (N_1946,N_1098,N_1483);
nor U1947 (N_1947,N_1201,N_1454);
and U1948 (N_1948,N_1480,N_1212);
and U1949 (N_1949,N_1106,N_1068);
xor U1950 (N_1950,N_1385,N_1207);
or U1951 (N_1951,N_1419,N_1433);
or U1952 (N_1952,N_1411,N_1005);
and U1953 (N_1953,N_1051,N_1358);
nand U1954 (N_1954,N_1343,N_1414);
xor U1955 (N_1955,N_1125,N_1291);
or U1956 (N_1956,N_1022,N_1246);
xnor U1957 (N_1957,N_1032,N_1492);
and U1958 (N_1958,N_1424,N_1453);
or U1959 (N_1959,N_1398,N_1262);
nand U1960 (N_1960,N_1281,N_1052);
xor U1961 (N_1961,N_1266,N_1127);
nand U1962 (N_1962,N_1434,N_1279);
xnor U1963 (N_1963,N_1081,N_1433);
nor U1964 (N_1964,N_1365,N_1217);
nand U1965 (N_1965,N_1168,N_1289);
xor U1966 (N_1966,N_1038,N_1359);
and U1967 (N_1967,N_1370,N_1062);
nor U1968 (N_1968,N_1190,N_1078);
nor U1969 (N_1969,N_1077,N_1428);
or U1970 (N_1970,N_1084,N_1197);
nand U1971 (N_1971,N_1230,N_1151);
and U1972 (N_1972,N_1055,N_1327);
and U1973 (N_1973,N_1370,N_1377);
nor U1974 (N_1974,N_1397,N_1237);
nand U1975 (N_1975,N_1189,N_1080);
nor U1976 (N_1976,N_1402,N_1258);
nor U1977 (N_1977,N_1113,N_1294);
or U1978 (N_1978,N_1473,N_1202);
and U1979 (N_1979,N_1294,N_1193);
nand U1980 (N_1980,N_1325,N_1359);
or U1981 (N_1981,N_1171,N_1187);
xor U1982 (N_1982,N_1102,N_1431);
nand U1983 (N_1983,N_1347,N_1316);
xnor U1984 (N_1984,N_1054,N_1418);
or U1985 (N_1985,N_1208,N_1449);
or U1986 (N_1986,N_1099,N_1085);
xor U1987 (N_1987,N_1484,N_1291);
xor U1988 (N_1988,N_1026,N_1331);
nand U1989 (N_1989,N_1006,N_1217);
nand U1990 (N_1990,N_1327,N_1486);
nor U1991 (N_1991,N_1342,N_1362);
nand U1992 (N_1992,N_1030,N_1183);
nand U1993 (N_1993,N_1411,N_1114);
xnor U1994 (N_1994,N_1072,N_1041);
nand U1995 (N_1995,N_1025,N_1221);
nor U1996 (N_1996,N_1270,N_1130);
nor U1997 (N_1997,N_1114,N_1424);
or U1998 (N_1998,N_1311,N_1479);
xor U1999 (N_1999,N_1314,N_1427);
or U2000 (N_2000,N_1776,N_1997);
nor U2001 (N_2001,N_1599,N_1533);
or U2002 (N_2002,N_1936,N_1931);
nor U2003 (N_2003,N_1510,N_1993);
and U2004 (N_2004,N_1565,N_1544);
and U2005 (N_2005,N_1849,N_1625);
nor U2006 (N_2006,N_1793,N_1698);
nor U2007 (N_2007,N_1669,N_1885);
xnor U2008 (N_2008,N_1954,N_1588);
xnor U2009 (N_2009,N_1674,N_1632);
or U2010 (N_2010,N_1508,N_1883);
or U2011 (N_2011,N_1903,N_1548);
or U2012 (N_2012,N_1767,N_1760);
nand U2013 (N_2013,N_1937,N_1904);
or U2014 (N_2014,N_1745,N_1718);
and U2015 (N_2015,N_1724,N_1703);
nand U2016 (N_2016,N_1956,N_1863);
xnor U2017 (N_2017,N_1605,N_1817);
nand U2018 (N_2018,N_1556,N_1946);
and U2019 (N_2019,N_1731,N_1733);
nor U2020 (N_2020,N_1995,N_1860);
or U2021 (N_2021,N_1546,N_1511);
or U2022 (N_2022,N_1716,N_1920);
nand U2023 (N_2023,N_1870,N_1528);
and U2024 (N_2024,N_1873,N_1626);
nand U2025 (N_2025,N_1827,N_1671);
or U2026 (N_2026,N_1816,N_1747);
or U2027 (N_2027,N_1711,N_1557);
nor U2028 (N_2028,N_1818,N_1868);
xnor U2029 (N_2029,N_1710,N_1551);
xor U2030 (N_2030,N_1647,N_1813);
xnor U2031 (N_2031,N_1771,N_1953);
or U2032 (N_2032,N_1730,N_1962);
xnor U2033 (N_2033,N_1622,N_1823);
nand U2034 (N_2034,N_1738,N_1694);
nand U2035 (N_2035,N_1643,N_1828);
nand U2036 (N_2036,N_1998,N_1811);
and U2037 (N_2037,N_1705,N_1968);
xor U2038 (N_2038,N_1985,N_1950);
xor U2039 (N_2039,N_1829,N_1838);
nor U2040 (N_2040,N_1629,N_1963);
and U2041 (N_2041,N_1875,N_1843);
nor U2042 (N_2042,N_1668,N_1642);
xnor U2043 (N_2043,N_1539,N_1696);
xnor U2044 (N_2044,N_1879,N_1513);
nand U2045 (N_2045,N_1725,N_1559);
nor U2046 (N_2046,N_1666,N_1803);
nand U2047 (N_2047,N_1789,N_1790);
and U2048 (N_2048,N_1919,N_1871);
nand U2049 (N_2049,N_1680,N_1742);
or U2050 (N_2050,N_1924,N_1939);
nor U2051 (N_2051,N_1825,N_1713);
xnor U2052 (N_2052,N_1646,N_1683);
and U2053 (N_2053,N_1639,N_1656);
xor U2054 (N_2054,N_1990,N_1612);
and U2055 (N_2055,N_1748,N_1610);
nand U2056 (N_2056,N_1844,N_1890);
nor U2057 (N_2057,N_1925,N_1787);
nor U2058 (N_2058,N_1611,N_1678);
xor U2059 (N_2059,N_1690,N_1603);
xor U2060 (N_2060,N_1580,N_1977);
nand U2061 (N_2061,N_1577,N_1504);
nand U2062 (N_2062,N_1943,N_1567);
or U2063 (N_2063,N_1799,N_1882);
xnor U2064 (N_2064,N_1571,N_1675);
or U2065 (N_2065,N_1880,N_1765);
nand U2066 (N_2066,N_1732,N_1630);
nand U2067 (N_2067,N_1794,N_1709);
nor U2068 (N_2068,N_1547,N_1653);
and U2069 (N_2069,N_1769,N_1992);
nor U2070 (N_2070,N_1948,N_1833);
or U2071 (N_2071,N_1581,N_1673);
xor U2072 (N_2072,N_1966,N_1706);
xnor U2073 (N_2073,N_1807,N_1652);
nor U2074 (N_2074,N_1561,N_1558);
nand U2075 (N_2075,N_1988,N_1623);
xor U2076 (N_2076,N_1785,N_1552);
nor U2077 (N_2077,N_1874,N_1714);
nand U2078 (N_2078,N_1834,N_1568);
nor U2079 (N_2079,N_1687,N_1695);
nor U2080 (N_2080,N_1831,N_1648);
nor U2081 (N_2081,N_1859,N_1501);
or U2082 (N_2082,N_1665,N_1543);
or U2083 (N_2083,N_1654,N_1979);
xnor U2084 (N_2084,N_1820,N_1999);
nor U2085 (N_2085,N_1585,N_1762);
xnor U2086 (N_2086,N_1633,N_1826);
nor U2087 (N_2087,N_1685,N_1505);
xnor U2088 (N_2088,N_1788,N_1726);
xnor U2089 (N_2089,N_1525,N_1965);
xor U2090 (N_2090,N_1692,N_1715);
nand U2091 (N_2091,N_1810,N_1905);
nor U2092 (N_2092,N_1851,N_1911);
xor U2093 (N_2093,N_1945,N_1894);
nand U2094 (N_2094,N_1514,N_1644);
nand U2095 (N_2095,N_1867,N_1524);
xor U2096 (N_2096,N_1969,N_1518);
or U2097 (N_2097,N_1502,N_1753);
nand U2098 (N_2098,N_1899,N_1516);
nor U2099 (N_2099,N_1907,N_1560);
xnor U2100 (N_2100,N_1822,N_1627);
or U2101 (N_2101,N_1841,N_1930);
or U2102 (N_2102,N_1881,N_1637);
and U2103 (N_2103,N_1719,N_1717);
nor U2104 (N_2104,N_1708,N_1529);
and U2105 (N_2105,N_1620,N_1846);
and U2106 (N_2106,N_1602,N_1888);
nor U2107 (N_2107,N_1676,N_1847);
xor U2108 (N_2108,N_1865,N_1951);
and U2109 (N_2109,N_1806,N_1645);
xnor U2110 (N_2110,N_1686,N_1712);
xnor U2111 (N_2111,N_1579,N_1592);
or U2112 (N_2112,N_1751,N_1781);
and U2113 (N_2113,N_1955,N_1815);
or U2114 (N_2114,N_1743,N_1667);
and U2115 (N_2115,N_1933,N_1621);
or U2116 (N_2116,N_1739,N_1512);
nand U2117 (N_2117,N_1857,N_1532);
and U2118 (N_2118,N_1897,N_1809);
and U2119 (N_2119,N_1974,N_1636);
or U2120 (N_2120,N_1624,N_1594);
xor U2121 (N_2121,N_1677,N_1606);
xor U2122 (N_2122,N_1596,N_1864);
or U2123 (N_2123,N_1804,N_1766);
xor U2124 (N_2124,N_1854,N_1728);
xnor U2125 (N_2125,N_1850,N_1791);
and U2126 (N_2126,N_1663,N_1910);
nand U2127 (N_2127,N_1964,N_1856);
nor U2128 (N_2128,N_1942,N_1978);
or U2129 (N_2129,N_1540,N_1835);
or U2130 (N_2130,N_1893,N_1901);
xor U2131 (N_2131,N_1613,N_1832);
nand U2132 (N_2132,N_1758,N_1536);
nand U2133 (N_2133,N_1628,N_1957);
xor U2134 (N_2134,N_1961,N_1898);
or U2135 (N_2135,N_1763,N_1682);
nand U2136 (N_2136,N_1576,N_1554);
and U2137 (N_2137,N_1520,N_1616);
or U2138 (N_2138,N_1757,N_1784);
xor U2139 (N_2139,N_1534,N_1651);
or U2140 (N_2140,N_1734,N_1858);
or U2141 (N_2141,N_1808,N_1770);
or U2142 (N_2142,N_1889,N_1779);
xor U2143 (N_2143,N_1506,N_1615);
and U2144 (N_2144,N_1658,N_1562);
xnor U2145 (N_2145,N_1523,N_1740);
nor U2146 (N_2146,N_1821,N_1775);
nand U2147 (N_2147,N_1866,N_1878);
and U2148 (N_2148,N_1641,N_1921);
nor U2149 (N_2149,N_1908,N_1564);
xnor U2150 (N_2150,N_1952,N_1575);
nor U2151 (N_2151,N_1940,N_1737);
xor U2152 (N_2152,N_1617,N_1563);
xor U2153 (N_2153,N_1587,N_1573);
nand U2154 (N_2154,N_1805,N_1824);
nor U2155 (N_2155,N_1507,N_1773);
nor U2156 (N_2156,N_1614,N_1600);
nand U2157 (N_2157,N_1782,N_1689);
xor U2158 (N_2158,N_1852,N_1982);
or U2159 (N_2159,N_1699,N_1601);
nor U2160 (N_2160,N_1700,N_1635);
or U2161 (N_2161,N_1991,N_1877);
or U2162 (N_2162,N_1792,N_1727);
and U2163 (N_2163,N_1721,N_1538);
nor U2164 (N_2164,N_1842,N_1927);
nor U2165 (N_2165,N_1741,N_1780);
or U2166 (N_2166,N_1526,N_1913);
nor U2167 (N_2167,N_1631,N_1723);
nand U2168 (N_2168,N_1944,N_1521);
nor U2169 (N_2169,N_1746,N_1752);
nand U2170 (N_2170,N_1574,N_1688);
and U2171 (N_2171,N_1607,N_1691);
nor U2172 (N_2172,N_1609,N_1959);
nand U2173 (N_2173,N_1650,N_1802);
nor U2174 (N_2174,N_1917,N_1972);
or U2175 (N_2175,N_1928,N_1918);
and U2176 (N_2176,N_1527,N_1996);
nor U2177 (N_2177,N_1778,N_1598);
or U2178 (N_2178,N_1976,N_1555);
and U2179 (N_2179,N_1915,N_1693);
and U2180 (N_2180,N_1761,N_1566);
xor U2181 (N_2181,N_1681,N_1736);
nand U2182 (N_2182,N_1500,N_1923);
xor U2183 (N_2183,N_1986,N_1672);
nor U2184 (N_2184,N_1720,N_1934);
nor U2185 (N_2185,N_1662,N_1589);
nor U2186 (N_2186,N_1941,N_1595);
nand U2187 (N_2187,N_1900,N_1970);
nand U2188 (N_2188,N_1545,N_1947);
and U2189 (N_2189,N_1649,N_1798);
and U2190 (N_2190,N_1553,N_1814);
nor U2191 (N_2191,N_1768,N_1517);
or U2192 (N_2192,N_1722,N_1619);
nand U2193 (N_2193,N_1584,N_1812);
nor U2194 (N_2194,N_1604,N_1801);
nand U2195 (N_2195,N_1912,N_1980);
and U2196 (N_2196,N_1896,N_1994);
xnor U2197 (N_2197,N_1892,N_1783);
nor U2198 (N_2198,N_1702,N_1704);
and U2199 (N_2199,N_1749,N_1519);
nand U2200 (N_2200,N_1891,N_1697);
xnor U2201 (N_2201,N_1759,N_1593);
nor U2202 (N_2202,N_1531,N_1530);
nand U2203 (N_2203,N_1906,N_1664);
and U2204 (N_2204,N_1922,N_1655);
nor U2205 (N_2205,N_1569,N_1729);
or U2206 (N_2206,N_1914,N_1884);
xnor U2207 (N_2207,N_1684,N_1861);
nor U2208 (N_2208,N_1756,N_1597);
xor U2209 (N_2209,N_1661,N_1967);
and U2210 (N_2210,N_1855,N_1872);
xor U2211 (N_2211,N_1935,N_1503);
xnor U2212 (N_2212,N_1679,N_1591);
nor U2213 (N_2213,N_1848,N_1839);
nand U2214 (N_2214,N_1670,N_1984);
xor U2215 (N_2215,N_1796,N_1583);
nor U2216 (N_2216,N_1657,N_1707);
nor U2217 (N_2217,N_1550,N_1640);
nand U2218 (N_2218,N_1537,N_1701);
and U2219 (N_2219,N_1830,N_1772);
xor U2220 (N_2220,N_1862,N_1960);
and U2221 (N_2221,N_1958,N_1618);
nor U2222 (N_2222,N_1975,N_1582);
or U2223 (N_2223,N_1515,N_1578);
xnor U2224 (N_2224,N_1837,N_1542);
nor U2225 (N_2225,N_1949,N_1886);
nor U2226 (N_2226,N_1754,N_1853);
or U2227 (N_2227,N_1797,N_1938);
nor U2228 (N_2228,N_1586,N_1869);
nand U2229 (N_2229,N_1549,N_1660);
nand U2230 (N_2230,N_1522,N_1971);
and U2231 (N_2231,N_1887,N_1845);
and U2232 (N_2232,N_1876,N_1572);
or U2233 (N_2233,N_1590,N_1786);
or U2234 (N_2234,N_1895,N_1983);
and U2235 (N_2235,N_1916,N_1774);
or U2236 (N_2236,N_1836,N_1973);
or U2237 (N_2237,N_1659,N_1541);
xor U2238 (N_2238,N_1735,N_1932);
nand U2239 (N_2239,N_1634,N_1750);
nor U2240 (N_2240,N_1638,N_1929);
nor U2241 (N_2241,N_1755,N_1926);
and U2242 (N_2242,N_1909,N_1570);
nor U2243 (N_2243,N_1819,N_1840);
nand U2244 (N_2244,N_1987,N_1800);
or U2245 (N_2245,N_1744,N_1509);
nor U2246 (N_2246,N_1608,N_1535);
nor U2247 (N_2247,N_1981,N_1989);
nand U2248 (N_2248,N_1795,N_1777);
nor U2249 (N_2249,N_1764,N_1902);
xor U2250 (N_2250,N_1602,N_1978);
nor U2251 (N_2251,N_1542,N_1694);
nor U2252 (N_2252,N_1693,N_1796);
and U2253 (N_2253,N_1717,N_1968);
or U2254 (N_2254,N_1569,N_1875);
nor U2255 (N_2255,N_1922,N_1595);
xnor U2256 (N_2256,N_1522,N_1721);
nor U2257 (N_2257,N_1807,N_1680);
nand U2258 (N_2258,N_1668,N_1925);
xnor U2259 (N_2259,N_1849,N_1958);
xor U2260 (N_2260,N_1606,N_1675);
nor U2261 (N_2261,N_1747,N_1779);
xor U2262 (N_2262,N_1506,N_1918);
and U2263 (N_2263,N_1540,N_1671);
xnor U2264 (N_2264,N_1507,N_1900);
xnor U2265 (N_2265,N_1746,N_1778);
nor U2266 (N_2266,N_1607,N_1980);
nand U2267 (N_2267,N_1949,N_1952);
nand U2268 (N_2268,N_1765,N_1502);
nor U2269 (N_2269,N_1501,N_1544);
nand U2270 (N_2270,N_1932,N_1616);
nand U2271 (N_2271,N_1552,N_1550);
xnor U2272 (N_2272,N_1837,N_1935);
xnor U2273 (N_2273,N_1612,N_1566);
xnor U2274 (N_2274,N_1688,N_1697);
nor U2275 (N_2275,N_1609,N_1666);
nand U2276 (N_2276,N_1792,N_1541);
nand U2277 (N_2277,N_1506,N_1985);
nand U2278 (N_2278,N_1552,N_1603);
nor U2279 (N_2279,N_1833,N_1865);
xor U2280 (N_2280,N_1972,N_1962);
or U2281 (N_2281,N_1816,N_1959);
and U2282 (N_2282,N_1861,N_1646);
nor U2283 (N_2283,N_1879,N_1612);
nand U2284 (N_2284,N_1999,N_1670);
or U2285 (N_2285,N_1628,N_1609);
nor U2286 (N_2286,N_1731,N_1796);
or U2287 (N_2287,N_1598,N_1924);
nand U2288 (N_2288,N_1791,N_1678);
xor U2289 (N_2289,N_1551,N_1805);
or U2290 (N_2290,N_1514,N_1801);
and U2291 (N_2291,N_1947,N_1680);
nand U2292 (N_2292,N_1997,N_1728);
or U2293 (N_2293,N_1995,N_1513);
and U2294 (N_2294,N_1950,N_1889);
and U2295 (N_2295,N_1554,N_1521);
or U2296 (N_2296,N_1915,N_1845);
or U2297 (N_2297,N_1539,N_1719);
nor U2298 (N_2298,N_1925,N_1985);
xor U2299 (N_2299,N_1581,N_1567);
xor U2300 (N_2300,N_1593,N_1923);
or U2301 (N_2301,N_1538,N_1664);
nor U2302 (N_2302,N_1577,N_1667);
or U2303 (N_2303,N_1667,N_1767);
or U2304 (N_2304,N_1835,N_1519);
nor U2305 (N_2305,N_1700,N_1758);
nor U2306 (N_2306,N_1763,N_1924);
nand U2307 (N_2307,N_1558,N_1690);
nor U2308 (N_2308,N_1787,N_1896);
or U2309 (N_2309,N_1906,N_1922);
or U2310 (N_2310,N_1595,N_1879);
nand U2311 (N_2311,N_1620,N_1792);
and U2312 (N_2312,N_1605,N_1759);
xnor U2313 (N_2313,N_1871,N_1506);
and U2314 (N_2314,N_1613,N_1769);
and U2315 (N_2315,N_1769,N_1520);
xnor U2316 (N_2316,N_1866,N_1894);
xor U2317 (N_2317,N_1683,N_1947);
nor U2318 (N_2318,N_1684,N_1803);
xnor U2319 (N_2319,N_1811,N_1859);
nor U2320 (N_2320,N_1934,N_1702);
xnor U2321 (N_2321,N_1703,N_1591);
nor U2322 (N_2322,N_1567,N_1578);
xnor U2323 (N_2323,N_1872,N_1596);
and U2324 (N_2324,N_1834,N_1898);
nand U2325 (N_2325,N_1836,N_1785);
xor U2326 (N_2326,N_1732,N_1992);
nor U2327 (N_2327,N_1810,N_1649);
nor U2328 (N_2328,N_1948,N_1550);
xnor U2329 (N_2329,N_1882,N_1965);
nand U2330 (N_2330,N_1941,N_1866);
nor U2331 (N_2331,N_1869,N_1990);
xnor U2332 (N_2332,N_1535,N_1914);
nor U2333 (N_2333,N_1517,N_1822);
nor U2334 (N_2334,N_1896,N_1575);
xnor U2335 (N_2335,N_1665,N_1808);
xnor U2336 (N_2336,N_1514,N_1998);
or U2337 (N_2337,N_1538,N_1591);
xor U2338 (N_2338,N_1653,N_1743);
and U2339 (N_2339,N_1827,N_1512);
xnor U2340 (N_2340,N_1981,N_1990);
xnor U2341 (N_2341,N_1915,N_1863);
and U2342 (N_2342,N_1868,N_1905);
nand U2343 (N_2343,N_1769,N_1700);
and U2344 (N_2344,N_1874,N_1979);
and U2345 (N_2345,N_1658,N_1706);
xnor U2346 (N_2346,N_1578,N_1557);
nand U2347 (N_2347,N_1647,N_1506);
or U2348 (N_2348,N_1591,N_1878);
xnor U2349 (N_2349,N_1536,N_1799);
and U2350 (N_2350,N_1636,N_1595);
nand U2351 (N_2351,N_1978,N_1664);
or U2352 (N_2352,N_1908,N_1551);
and U2353 (N_2353,N_1687,N_1736);
nor U2354 (N_2354,N_1532,N_1850);
nor U2355 (N_2355,N_1832,N_1650);
nor U2356 (N_2356,N_1916,N_1957);
and U2357 (N_2357,N_1949,N_1975);
nor U2358 (N_2358,N_1742,N_1625);
and U2359 (N_2359,N_1573,N_1651);
nor U2360 (N_2360,N_1857,N_1751);
xnor U2361 (N_2361,N_1858,N_1502);
xnor U2362 (N_2362,N_1788,N_1601);
and U2363 (N_2363,N_1615,N_1596);
nand U2364 (N_2364,N_1516,N_1800);
nor U2365 (N_2365,N_1886,N_1678);
xor U2366 (N_2366,N_1729,N_1758);
nor U2367 (N_2367,N_1707,N_1641);
and U2368 (N_2368,N_1909,N_1919);
or U2369 (N_2369,N_1885,N_1938);
nand U2370 (N_2370,N_1966,N_1594);
nand U2371 (N_2371,N_1845,N_1543);
or U2372 (N_2372,N_1744,N_1817);
xor U2373 (N_2373,N_1633,N_1606);
nand U2374 (N_2374,N_1960,N_1634);
nand U2375 (N_2375,N_1858,N_1727);
and U2376 (N_2376,N_1839,N_1703);
xnor U2377 (N_2377,N_1985,N_1710);
nor U2378 (N_2378,N_1665,N_1845);
xor U2379 (N_2379,N_1610,N_1681);
or U2380 (N_2380,N_1548,N_1854);
or U2381 (N_2381,N_1747,N_1922);
nor U2382 (N_2382,N_1820,N_1518);
and U2383 (N_2383,N_1829,N_1670);
or U2384 (N_2384,N_1559,N_1650);
nor U2385 (N_2385,N_1989,N_1917);
or U2386 (N_2386,N_1654,N_1675);
nor U2387 (N_2387,N_1933,N_1614);
xor U2388 (N_2388,N_1831,N_1733);
nor U2389 (N_2389,N_1774,N_1523);
xnor U2390 (N_2390,N_1712,N_1756);
xor U2391 (N_2391,N_1543,N_1713);
nand U2392 (N_2392,N_1883,N_1897);
nand U2393 (N_2393,N_1924,N_1556);
xnor U2394 (N_2394,N_1578,N_1659);
or U2395 (N_2395,N_1520,N_1522);
nand U2396 (N_2396,N_1568,N_1604);
nand U2397 (N_2397,N_1788,N_1774);
xnor U2398 (N_2398,N_1939,N_1838);
nor U2399 (N_2399,N_1998,N_1879);
xor U2400 (N_2400,N_1678,N_1692);
xnor U2401 (N_2401,N_1683,N_1504);
or U2402 (N_2402,N_1535,N_1840);
nand U2403 (N_2403,N_1668,N_1550);
nor U2404 (N_2404,N_1649,N_1954);
xnor U2405 (N_2405,N_1557,N_1971);
nand U2406 (N_2406,N_1761,N_1656);
xor U2407 (N_2407,N_1711,N_1859);
nor U2408 (N_2408,N_1513,N_1865);
xnor U2409 (N_2409,N_1872,N_1751);
nand U2410 (N_2410,N_1940,N_1864);
nor U2411 (N_2411,N_1871,N_1677);
and U2412 (N_2412,N_1653,N_1776);
or U2413 (N_2413,N_1500,N_1611);
xnor U2414 (N_2414,N_1890,N_1900);
xnor U2415 (N_2415,N_1943,N_1990);
or U2416 (N_2416,N_1880,N_1695);
and U2417 (N_2417,N_1883,N_1970);
and U2418 (N_2418,N_1839,N_1917);
and U2419 (N_2419,N_1561,N_1954);
nor U2420 (N_2420,N_1604,N_1767);
and U2421 (N_2421,N_1952,N_1753);
nor U2422 (N_2422,N_1803,N_1997);
or U2423 (N_2423,N_1860,N_1844);
or U2424 (N_2424,N_1686,N_1939);
or U2425 (N_2425,N_1776,N_1632);
nand U2426 (N_2426,N_1944,N_1543);
or U2427 (N_2427,N_1857,N_1752);
and U2428 (N_2428,N_1988,N_1744);
nand U2429 (N_2429,N_1625,N_1937);
xnor U2430 (N_2430,N_1639,N_1920);
or U2431 (N_2431,N_1844,N_1641);
and U2432 (N_2432,N_1615,N_1887);
or U2433 (N_2433,N_1646,N_1524);
and U2434 (N_2434,N_1532,N_1920);
nand U2435 (N_2435,N_1725,N_1895);
xor U2436 (N_2436,N_1880,N_1900);
nand U2437 (N_2437,N_1748,N_1759);
and U2438 (N_2438,N_1882,N_1659);
and U2439 (N_2439,N_1990,N_1635);
or U2440 (N_2440,N_1864,N_1838);
or U2441 (N_2441,N_1507,N_1957);
xor U2442 (N_2442,N_1964,N_1670);
and U2443 (N_2443,N_1977,N_1932);
xnor U2444 (N_2444,N_1933,N_1717);
and U2445 (N_2445,N_1554,N_1913);
nand U2446 (N_2446,N_1967,N_1524);
nand U2447 (N_2447,N_1947,N_1961);
nand U2448 (N_2448,N_1809,N_1530);
nor U2449 (N_2449,N_1592,N_1938);
xor U2450 (N_2450,N_1848,N_1845);
nand U2451 (N_2451,N_1723,N_1501);
or U2452 (N_2452,N_1652,N_1991);
nor U2453 (N_2453,N_1536,N_1951);
nand U2454 (N_2454,N_1661,N_1961);
nand U2455 (N_2455,N_1938,N_1791);
or U2456 (N_2456,N_1806,N_1997);
and U2457 (N_2457,N_1899,N_1751);
nand U2458 (N_2458,N_1921,N_1558);
xor U2459 (N_2459,N_1660,N_1576);
xor U2460 (N_2460,N_1896,N_1730);
nor U2461 (N_2461,N_1745,N_1898);
xor U2462 (N_2462,N_1654,N_1512);
nor U2463 (N_2463,N_1564,N_1974);
xnor U2464 (N_2464,N_1719,N_1614);
and U2465 (N_2465,N_1809,N_1580);
nor U2466 (N_2466,N_1769,N_1548);
nand U2467 (N_2467,N_1606,N_1656);
or U2468 (N_2468,N_1790,N_1766);
nor U2469 (N_2469,N_1821,N_1513);
or U2470 (N_2470,N_1661,N_1845);
nor U2471 (N_2471,N_1548,N_1663);
xnor U2472 (N_2472,N_1771,N_1561);
and U2473 (N_2473,N_1927,N_1529);
nor U2474 (N_2474,N_1522,N_1503);
nand U2475 (N_2475,N_1506,N_1609);
or U2476 (N_2476,N_1860,N_1653);
or U2477 (N_2477,N_1703,N_1687);
and U2478 (N_2478,N_1811,N_1936);
xnor U2479 (N_2479,N_1792,N_1505);
xor U2480 (N_2480,N_1611,N_1875);
and U2481 (N_2481,N_1574,N_1875);
xnor U2482 (N_2482,N_1945,N_1948);
nor U2483 (N_2483,N_1564,N_1609);
xor U2484 (N_2484,N_1773,N_1563);
xor U2485 (N_2485,N_1757,N_1544);
nor U2486 (N_2486,N_1554,N_1610);
nand U2487 (N_2487,N_1980,N_1920);
or U2488 (N_2488,N_1510,N_1721);
or U2489 (N_2489,N_1589,N_1558);
nor U2490 (N_2490,N_1669,N_1562);
nor U2491 (N_2491,N_1902,N_1940);
and U2492 (N_2492,N_1808,N_1666);
or U2493 (N_2493,N_1991,N_1567);
xnor U2494 (N_2494,N_1670,N_1841);
nand U2495 (N_2495,N_1775,N_1789);
nand U2496 (N_2496,N_1950,N_1552);
xor U2497 (N_2497,N_1697,N_1830);
or U2498 (N_2498,N_1644,N_1547);
or U2499 (N_2499,N_1750,N_1879);
and U2500 (N_2500,N_2368,N_2115);
and U2501 (N_2501,N_2113,N_2092);
and U2502 (N_2502,N_2342,N_2212);
or U2503 (N_2503,N_2074,N_2458);
xor U2504 (N_2504,N_2063,N_2420);
xnor U2505 (N_2505,N_2265,N_2130);
nand U2506 (N_2506,N_2390,N_2499);
or U2507 (N_2507,N_2371,N_2125);
or U2508 (N_2508,N_2207,N_2337);
nand U2509 (N_2509,N_2355,N_2197);
nor U2510 (N_2510,N_2041,N_2440);
nand U2511 (N_2511,N_2132,N_2021);
or U2512 (N_2512,N_2443,N_2338);
xnor U2513 (N_2513,N_2373,N_2426);
nand U2514 (N_2514,N_2104,N_2099);
nand U2515 (N_2515,N_2190,N_2419);
or U2516 (N_2516,N_2131,N_2225);
xor U2517 (N_2517,N_2112,N_2375);
nor U2518 (N_2518,N_2097,N_2055);
nor U2519 (N_2519,N_2129,N_2234);
nor U2520 (N_2520,N_2155,N_2363);
xnor U2521 (N_2521,N_2464,N_2404);
and U2522 (N_2522,N_2444,N_2106);
or U2523 (N_2523,N_2157,N_2459);
and U2524 (N_2524,N_2107,N_2076);
or U2525 (N_2525,N_2481,N_2300);
and U2526 (N_2526,N_2291,N_2033);
nand U2527 (N_2527,N_2386,N_2474);
nor U2528 (N_2528,N_2172,N_2066);
nand U2529 (N_2529,N_2057,N_2069);
or U2530 (N_2530,N_2196,N_2116);
nor U2531 (N_2531,N_2446,N_2396);
xnor U2532 (N_2532,N_2143,N_2242);
xor U2533 (N_2533,N_2455,N_2009);
nor U2534 (N_2534,N_2409,N_2203);
and U2535 (N_2535,N_2087,N_2414);
and U2536 (N_2536,N_2036,N_2179);
nor U2537 (N_2537,N_2269,N_2405);
nand U2538 (N_2538,N_2495,N_2306);
and U2539 (N_2539,N_2392,N_2438);
or U2540 (N_2540,N_2199,N_2216);
nand U2541 (N_2541,N_2456,N_2461);
and U2542 (N_2542,N_2428,N_2209);
and U2543 (N_2543,N_2309,N_2108);
xnor U2544 (N_2544,N_2410,N_2407);
and U2545 (N_2545,N_2360,N_2078);
nor U2546 (N_2546,N_2437,N_2353);
or U2547 (N_2547,N_2256,N_2003);
and U2548 (N_2548,N_2367,N_2093);
or U2549 (N_2549,N_2408,N_2475);
and U2550 (N_2550,N_2297,N_2156);
nor U2551 (N_2551,N_2303,N_2241);
or U2552 (N_2552,N_2255,N_2124);
and U2553 (N_2553,N_2029,N_2259);
or U2554 (N_2554,N_2311,N_2073);
nand U2555 (N_2555,N_2401,N_2151);
and U2556 (N_2556,N_2230,N_2096);
nor U2557 (N_2557,N_2340,N_2295);
or U2558 (N_2558,N_2202,N_2434);
or U2559 (N_2559,N_2079,N_2201);
nor U2560 (N_2560,N_2313,N_2416);
nor U2561 (N_2561,N_2288,N_2145);
nor U2562 (N_2562,N_2227,N_2307);
and U2563 (N_2563,N_2492,N_2469);
or U2564 (N_2564,N_2118,N_2090);
xor U2565 (N_2565,N_2171,N_2089);
or U2566 (N_2566,N_2482,N_2277);
and U2567 (N_2567,N_2028,N_2217);
xnor U2568 (N_2568,N_2232,N_2000);
and U2569 (N_2569,N_2284,N_2460);
nand U2570 (N_2570,N_2447,N_2394);
nor U2571 (N_2571,N_2483,N_2005);
and U2572 (N_2572,N_2356,N_2324);
xnor U2573 (N_2573,N_2065,N_2442);
or U2574 (N_2574,N_2173,N_2215);
nor U2575 (N_2575,N_2228,N_2180);
and U2576 (N_2576,N_2233,N_2214);
or U2577 (N_2577,N_2127,N_2039);
nand U2578 (N_2578,N_2035,N_2183);
nand U2579 (N_2579,N_2466,N_2161);
nand U2580 (N_2580,N_2347,N_2208);
nor U2581 (N_2581,N_2421,N_2372);
nor U2582 (N_2582,N_2048,N_2378);
nor U2583 (N_2583,N_2285,N_2123);
and U2584 (N_2584,N_2126,N_2266);
and U2585 (N_2585,N_2218,N_2162);
xnor U2586 (N_2586,N_2471,N_2080);
or U2587 (N_2587,N_2054,N_2182);
or U2588 (N_2588,N_2397,N_2398);
and U2589 (N_2589,N_2491,N_2168);
xnor U2590 (N_2590,N_2185,N_2484);
nor U2591 (N_2591,N_2240,N_2268);
xor U2592 (N_2592,N_2374,N_2067);
and U2593 (N_2593,N_2120,N_2321);
and U2594 (N_2594,N_2280,N_2463);
nor U2595 (N_2595,N_2134,N_2023);
xor U2596 (N_2596,N_2271,N_2279);
xnor U2597 (N_2597,N_2441,N_2453);
and U2598 (N_2598,N_2423,N_2015);
nand U2599 (N_2599,N_2301,N_2133);
and U2600 (N_2600,N_2263,N_2012);
xnor U2601 (N_2601,N_2071,N_2387);
or U2602 (N_2602,N_2333,N_2062);
and U2603 (N_2603,N_2494,N_2072);
and U2604 (N_2604,N_2247,N_2302);
or U2605 (N_2605,N_2184,N_2273);
and U2606 (N_2606,N_2343,N_2310);
xnor U2607 (N_2607,N_2429,N_2200);
nor U2608 (N_2608,N_2351,N_2457);
nand U2609 (N_2609,N_2010,N_2357);
and U2610 (N_2610,N_2478,N_2358);
nor U2611 (N_2611,N_2329,N_2350);
or U2612 (N_2612,N_2320,N_2019);
nor U2613 (N_2613,N_2485,N_2159);
nor U2614 (N_2614,N_2046,N_2293);
nor U2615 (N_2615,N_2117,N_2431);
and U2616 (N_2616,N_2417,N_2270);
nor U2617 (N_2617,N_2014,N_2045);
and U2618 (N_2618,N_2229,N_2348);
xor U2619 (N_2619,N_2341,N_2094);
nor U2620 (N_2620,N_2486,N_2448);
and U2621 (N_2621,N_2305,N_2002);
or U2622 (N_2622,N_2136,N_2052);
and U2623 (N_2623,N_2177,N_2181);
nor U2624 (N_2624,N_2498,N_2406);
nor U2625 (N_2625,N_2322,N_2439);
xnor U2626 (N_2626,N_2210,N_2163);
nand U2627 (N_2627,N_2206,N_2140);
or U2628 (N_2628,N_2379,N_2354);
xor U2629 (N_2629,N_2236,N_2026);
xor U2630 (N_2630,N_2415,N_2088);
nor U2631 (N_2631,N_2292,N_2344);
xor U2632 (N_2632,N_2211,N_2352);
nor U2633 (N_2633,N_2186,N_2135);
xor U2634 (N_2634,N_2473,N_2105);
xor U2635 (N_2635,N_2468,N_2020);
or U2636 (N_2636,N_2056,N_2146);
nor U2637 (N_2637,N_2403,N_2017);
nor U2638 (N_2638,N_2391,N_2245);
nor U2639 (N_2639,N_2169,N_2058);
and U2640 (N_2640,N_2102,N_2122);
xor U2641 (N_2641,N_2274,N_2487);
and U2642 (N_2642,N_2477,N_2275);
nand U2643 (N_2643,N_2189,N_2287);
nor U2644 (N_2644,N_2361,N_2025);
nor U2645 (N_2645,N_2221,N_2298);
nor U2646 (N_2646,N_2148,N_2308);
xnor U2647 (N_2647,N_2219,N_2433);
nor U2648 (N_2648,N_2490,N_2011);
nor U2649 (N_2649,N_2064,N_2164);
nor U2650 (N_2650,N_2328,N_2304);
nand U2651 (N_2651,N_2038,N_2142);
or U2652 (N_2652,N_2004,N_2091);
or U2653 (N_2653,N_2224,N_2138);
and U2654 (N_2654,N_2030,N_2339);
or U2655 (N_2655,N_2411,N_2061);
nor U2656 (N_2656,N_2100,N_2318);
or U2657 (N_2657,N_2170,N_2059);
xnor U2658 (N_2658,N_2497,N_2006);
and U2659 (N_2659,N_2384,N_2383);
nor U2660 (N_2660,N_2031,N_2213);
xor U2661 (N_2661,N_2278,N_2174);
or U2662 (N_2662,N_2489,N_2252);
and U2663 (N_2663,N_2472,N_2149);
xor U2664 (N_2664,N_2086,N_2267);
or U2665 (N_2665,N_2018,N_2204);
xnor U2666 (N_2666,N_2470,N_2412);
and U2667 (N_2667,N_2098,N_2111);
xnor U2668 (N_2668,N_2317,N_2034);
or U2669 (N_2669,N_2075,N_2042);
nor U2670 (N_2670,N_2253,N_2244);
and U2671 (N_2671,N_2257,N_2314);
nor U2672 (N_2672,N_2121,N_2312);
or U2673 (N_2673,N_2488,N_2334);
nor U2674 (N_2674,N_2399,N_2037);
and U2675 (N_2675,N_2262,N_2144);
nor U2676 (N_2676,N_2068,N_2449);
nor U2677 (N_2677,N_2496,N_2137);
xor U2678 (N_2678,N_2032,N_2335);
xor U2679 (N_2679,N_2141,N_2395);
nand U2680 (N_2680,N_2243,N_2016);
and U2681 (N_2681,N_2049,N_2047);
nor U2682 (N_2682,N_2422,N_2480);
or U2683 (N_2683,N_2381,N_2198);
and U2684 (N_2684,N_2479,N_2007);
and U2685 (N_2685,N_2283,N_2476);
nor U2686 (N_2686,N_2188,N_2024);
xnor U2687 (N_2687,N_2336,N_2194);
and U2688 (N_2688,N_2349,N_2220);
nand U2689 (N_2689,N_2346,N_2050);
xnor U2690 (N_2690,N_2070,N_2154);
or U2691 (N_2691,N_2109,N_2082);
and U2692 (N_2692,N_2187,N_2178);
and U2693 (N_2693,N_2326,N_2299);
or U2694 (N_2694,N_2128,N_2081);
xnor U2695 (N_2695,N_2493,N_2424);
nor U2696 (N_2696,N_2235,N_2451);
or U2697 (N_2697,N_2425,N_2246);
and U2698 (N_2698,N_2452,N_2250);
xor U2699 (N_2699,N_2260,N_2281);
or U2700 (N_2700,N_2327,N_2316);
and U2701 (N_2701,N_2195,N_2147);
and U2702 (N_2702,N_2237,N_2053);
and U2703 (N_2703,N_2231,N_2315);
nor U2704 (N_2704,N_2223,N_2150);
or U2705 (N_2705,N_2380,N_2393);
xnor U2706 (N_2706,N_2289,N_2119);
nand U2707 (N_2707,N_2332,N_2249);
nor U2708 (N_2708,N_2191,N_2192);
nand U2709 (N_2709,N_2366,N_2286);
nor U2710 (N_2710,N_2158,N_2238);
and U2711 (N_2711,N_2103,N_2044);
and U2712 (N_2712,N_2051,N_2462);
nand U2713 (N_2713,N_2258,N_2402);
or U2714 (N_2714,N_2114,N_2264);
or U2715 (N_2715,N_2345,N_2369);
xor U2716 (N_2716,N_2465,N_2382);
nor U2717 (N_2717,N_2251,N_2254);
nor U2718 (N_2718,N_2290,N_2084);
xor U2719 (N_2719,N_2110,N_2272);
xnor U2720 (N_2720,N_2282,N_2400);
xor U2721 (N_2721,N_2060,N_2325);
nand U2722 (N_2722,N_2364,N_2435);
and U2723 (N_2723,N_2467,N_2239);
nor U2724 (N_2724,N_2362,N_2450);
nand U2725 (N_2725,N_2176,N_2013);
xnor U2726 (N_2726,N_2043,N_2331);
nand U2727 (N_2727,N_2040,N_2077);
nand U2728 (N_2728,N_2085,N_2294);
and U2729 (N_2729,N_2248,N_2413);
nor U2730 (N_2730,N_2323,N_2376);
and U2731 (N_2731,N_2167,N_2418);
xnor U2732 (N_2732,N_2296,N_2359);
or U2733 (N_2733,N_2153,N_2436);
nor U2734 (N_2734,N_2226,N_2261);
or U2735 (N_2735,N_2365,N_2101);
and U2736 (N_2736,N_2432,N_2445);
or U2737 (N_2737,N_2388,N_2370);
and U2738 (N_2738,N_2152,N_2377);
or U2739 (N_2739,N_2166,N_2022);
nor U2740 (N_2740,N_2385,N_2001);
or U2741 (N_2741,N_2193,N_2083);
or U2742 (N_2742,N_2095,N_2175);
nand U2743 (N_2743,N_2139,N_2454);
xor U2744 (N_2744,N_2008,N_2276);
nor U2745 (N_2745,N_2430,N_2027);
nor U2746 (N_2746,N_2160,N_2427);
or U2747 (N_2747,N_2222,N_2389);
or U2748 (N_2748,N_2330,N_2205);
or U2749 (N_2749,N_2165,N_2319);
xnor U2750 (N_2750,N_2368,N_2199);
or U2751 (N_2751,N_2049,N_2325);
or U2752 (N_2752,N_2006,N_2395);
or U2753 (N_2753,N_2133,N_2411);
xnor U2754 (N_2754,N_2217,N_2330);
and U2755 (N_2755,N_2385,N_2187);
and U2756 (N_2756,N_2207,N_2363);
nand U2757 (N_2757,N_2243,N_2361);
xor U2758 (N_2758,N_2293,N_2479);
nor U2759 (N_2759,N_2496,N_2185);
xor U2760 (N_2760,N_2471,N_2367);
or U2761 (N_2761,N_2237,N_2417);
nor U2762 (N_2762,N_2009,N_2274);
nor U2763 (N_2763,N_2319,N_2240);
and U2764 (N_2764,N_2377,N_2479);
nand U2765 (N_2765,N_2115,N_2283);
nor U2766 (N_2766,N_2216,N_2213);
and U2767 (N_2767,N_2326,N_2267);
and U2768 (N_2768,N_2305,N_2450);
nand U2769 (N_2769,N_2171,N_2125);
nand U2770 (N_2770,N_2462,N_2490);
xnor U2771 (N_2771,N_2038,N_2174);
or U2772 (N_2772,N_2495,N_2048);
nand U2773 (N_2773,N_2467,N_2108);
xnor U2774 (N_2774,N_2283,N_2024);
and U2775 (N_2775,N_2053,N_2421);
or U2776 (N_2776,N_2218,N_2417);
or U2777 (N_2777,N_2138,N_2232);
nand U2778 (N_2778,N_2184,N_2460);
nor U2779 (N_2779,N_2142,N_2051);
xor U2780 (N_2780,N_2062,N_2125);
nor U2781 (N_2781,N_2378,N_2348);
or U2782 (N_2782,N_2437,N_2485);
nor U2783 (N_2783,N_2402,N_2468);
nand U2784 (N_2784,N_2096,N_2080);
xnor U2785 (N_2785,N_2270,N_2165);
nand U2786 (N_2786,N_2269,N_2025);
nand U2787 (N_2787,N_2276,N_2347);
xor U2788 (N_2788,N_2058,N_2035);
nor U2789 (N_2789,N_2444,N_2023);
nand U2790 (N_2790,N_2428,N_2062);
xnor U2791 (N_2791,N_2351,N_2266);
and U2792 (N_2792,N_2352,N_2132);
nand U2793 (N_2793,N_2326,N_2110);
nor U2794 (N_2794,N_2448,N_2375);
and U2795 (N_2795,N_2069,N_2186);
nand U2796 (N_2796,N_2049,N_2075);
nand U2797 (N_2797,N_2191,N_2110);
nand U2798 (N_2798,N_2145,N_2367);
or U2799 (N_2799,N_2386,N_2363);
nand U2800 (N_2800,N_2048,N_2316);
or U2801 (N_2801,N_2463,N_2479);
or U2802 (N_2802,N_2219,N_2143);
xor U2803 (N_2803,N_2440,N_2359);
xor U2804 (N_2804,N_2419,N_2013);
nand U2805 (N_2805,N_2400,N_2024);
nor U2806 (N_2806,N_2414,N_2232);
nor U2807 (N_2807,N_2005,N_2211);
nand U2808 (N_2808,N_2469,N_2148);
nand U2809 (N_2809,N_2372,N_2103);
and U2810 (N_2810,N_2474,N_2336);
xnor U2811 (N_2811,N_2431,N_2136);
nor U2812 (N_2812,N_2012,N_2186);
or U2813 (N_2813,N_2100,N_2330);
xnor U2814 (N_2814,N_2265,N_2163);
xor U2815 (N_2815,N_2498,N_2091);
xnor U2816 (N_2816,N_2098,N_2469);
or U2817 (N_2817,N_2110,N_2231);
nand U2818 (N_2818,N_2126,N_2395);
nand U2819 (N_2819,N_2114,N_2084);
nor U2820 (N_2820,N_2200,N_2397);
xnor U2821 (N_2821,N_2128,N_2115);
xnor U2822 (N_2822,N_2267,N_2365);
or U2823 (N_2823,N_2206,N_2220);
xor U2824 (N_2824,N_2272,N_2137);
or U2825 (N_2825,N_2456,N_2355);
nand U2826 (N_2826,N_2130,N_2185);
xnor U2827 (N_2827,N_2016,N_2164);
nand U2828 (N_2828,N_2480,N_2338);
and U2829 (N_2829,N_2101,N_2210);
nor U2830 (N_2830,N_2062,N_2314);
nand U2831 (N_2831,N_2084,N_2444);
and U2832 (N_2832,N_2230,N_2123);
or U2833 (N_2833,N_2391,N_2012);
nand U2834 (N_2834,N_2264,N_2207);
nand U2835 (N_2835,N_2202,N_2190);
nor U2836 (N_2836,N_2125,N_2475);
xor U2837 (N_2837,N_2068,N_2410);
and U2838 (N_2838,N_2351,N_2255);
nor U2839 (N_2839,N_2396,N_2115);
xnor U2840 (N_2840,N_2450,N_2330);
xnor U2841 (N_2841,N_2486,N_2221);
xnor U2842 (N_2842,N_2094,N_2049);
nand U2843 (N_2843,N_2127,N_2050);
or U2844 (N_2844,N_2403,N_2146);
nor U2845 (N_2845,N_2137,N_2374);
or U2846 (N_2846,N_2359,N_2300);
and U2847 (N_2847,N_2134,N_2380);
nand U2848 (N_2848,N_2276,N_2239);
xnor U2849 (N_2849,N_2326,N_2197);
nand U2850 (N_2850,N_2215,N_2367);
xor U2851 (N_2851,N_2078,N_2289);
nor U2852 (N_2852,N_2291,N_2036);
nand U2853 (N_2853,N_2051,N_2203);
or U2854 (N_2854,N_2327,N_2308);
nor U2855 (N_2855,N_2186,N_2305);
or U2856 (N_2856,N_2144,N_2116);
nor U2857 (N_2857,N_2019,N_2028);
and U2858 (N_2858,N_2080,N_2070);
nor U2859 (N_2859,N_2463,N_2097);
and U2860 (N_2860,N_2439,N_2418);
or U2861 (N_2861,N_2191,N_2188);
or U2862 (N_2862,N_2475,N_2380);
nor U2863 (N_2863,N_2300,N_2026);
nor U2864 (N_2864,N_2435,N_2046);
nand U2865 (N_2865,N_2468,N_2250);
or U2866 (N_2866,N_2088,N_2021);
xnor U2867 (N_2867,N_2038,N_2305);
nand U2868 (N_2868,N_2475,N_2130);
nand U2869 (N_2869,N_2432,N_2113);
xnor U2870 (N_2870,N_2324,N_2230);
and U2871 (N_2871,N_2374,N_2095);
xnor U2872 (N_2872,N_2423,N_2038);
nor U2873 (N_2873,N_2190,N_2165);
xor U2874 (N_2874,N_2024,N_2041);
nand U2875 (N_2875,N_2266,N_2140);
or U2876 (N_2876,N_2183,N_2203);
nand U2877 (N_2877,N_2040,N_2478);
and U2878 (N_2878,N_2250,N_2011);
or U2879 (N_2879,N_2239,N_2168);
nor U2880 (N_2880,N_2215,N_2294);
nor U2881 (N_2881,N_2034,N_2423);
xor U2882 (N_2882,N_2170,N_2438);
or U2883 (N_2883,N_2210,N_2325);
and U2884 (N_2884,N_2211,N_2073);
xnor U2885 (N_2885,N_2112,N_2040);
and U2886 (N_2886,N_2490,N_2152);
and U2887 (N_2887,N_2291,N_2048);
and U2888 (N_2888,N_2324,N_2210);
xor U2889 (N_2889,N_2060,N_2382);
and U2890 (N_2890,N_2050,N_2261);
xor U2891 (N_2891,N_2422,N_2351);
nor U2892 (N_2892,N_2053,N_2474);
and U2893 (N_2893,N_2030,N_2278);
or U2894 (N_2894,N_2411,N_2413);
and U2895 (N_2895,N_2445,N_2431);
nand U2896 (N_2896,N_2067,N_2281);
nand U2897 (N_2897,N_2214,N_2495);
and U2898 (N_2898,N_2345,N_2488);
and U2899 (N_2899,N_2066,N_2045);
and U2900 (N_2900,N_2261,N_2406);
and U2901 (N_2901,N_2046,N_2101);
nand U2902 (N_2902,N_2059,N_2082);
and U2903 (N_2903,N_2172,N_2384);
nor U2904 (N_2904,N_2134,N_2048);
nor U2905 (N_2905,N_2344,N_2285);
xnor U2906 (N_2906,N_2031,N_2326);
and U2907 (N_2907,N_2328,N_2161);
and U2908 (N_2908,N_2056,N_2481);
and U2909 (N_2909,N_2277,N_2139);
or U2910 (N_2910,N_2061,N_2332);
nor U2911 (N_2911,N_2363,N_2433);
nand U2912 (N_2912,N_2172,N_2151);
nor U2913 (N_2913,N_2333,N_2204);
nand U2914 (N_2914,N_2339,N_2142);
nand U2915 (N_2915,N_2282,N_2476);
xnor U2916 (N_2916,N_2125,N_2217);
nand U2917 (N_2917,N_2082,N_2035);
xnor U2918 (N_2918,N_2438,N_2040);
or U2919 (N_2919,N_2049,N_2014);
nor U2920 (N_2920,N_2142,N_2455);
or U2921 (N_2921,N_2307,N_2290);
nor U2922 (N_2922,N_2412,N_2059);
xor U2923 (N_2923,N_2214,N_2089);
or U2924 (N_2924,N_2120,N_2240);
nor U2925 (N_2925,N_2483,N_2214);
and U2926 (N_2926,N_2260,N_2453);
or U2927 (N_2927,N_2120,N_2436);
nor U2928 (N_2928,N_2446,N_2292);
xor U2929 (N_2929,N_2305,N_2423);
or U2930 (N_2930,N_2436,N_2260);
nand U2931 (N_2931,N_2407,N_2434);
nor U2932 (N_2932,N_2121,N_2282);
nand U2933 (N_2933,N_2369,N_2404);
and U2934 (N_2934,N_2134,N_2149);
xnor U2935 (N_2935,N_2154,N_2129);
or U2936 (N_2936,N_2061,N_2408);
xnor U2937 (N_2937,N_2334,N_2082);
xnor U2938 (N_2938,N_2033,N_2165);
xor U2939 (N_2939,N_2403,N_2421);
or U2940 (N_2940,N_2281,N_2094);
nor U2941 (N_2941,N_2409,N_2105);
or U2942 (N_2942,N_2456,N_2261);
nand U2943 (N_2943,N_2156,N_2344);
or U2944 (N_2944,N_2473,N_2437);
xnor U2945 (N_2945,N_2418,N_2412);
nand U2946 (N_2946,N_2134,N_2345);
and U2947 (N_2947,N_2260,N_2474);
and U2948 (N_2948,N_2276,N_2329);
nor U2949 (N_2949,N_2379,N_2065);
or U2950 (N_2950,N_2226,N_2356);
xor U2951 (N_2951,N_2009,N_2475);
nand U2952 (N_2952,N_2266,N_2447);
xor U2953 (N_2953,N_2445,N_2055);
or U2954 (N_2954,N_2068,N_2095);
nor U2955 (N_2955,N_2242,N_2189);
xor U2956 (N_2956,N_2262,N_2320);
and U2957 (N_2957,N_2364,N_2267);
nand U2958 (N_2958,N_2322,N_2409);
xnor U2959 (N_2959,N_2195,N_2266);
or U2960 (N_2960,N_2480,N_2287);
nand U2961 (N_2961,N_2262,N_2196);
xor U2962 (N_2962,N_2146,N_2221);
nand U2963 (N_2963,N_2261,N_2113);
nor U2964 (N_2964,N_2160,N_2487);
nor U2965 (N_2965,N_2363,N_2330);
nand U2966 (N_2966,N_2329,N_2499);
or U2967 (N_2967,N_2257,N_2086);
or U2968 (N_2968,N_2249,N_2116);
and U2969 (N_2969,N_2026,N_2389);
nand U2970 (N_2970,N_2492,N_2122);
or U2971 (N_2971,N_2024,N_2237);
xnor U2972 (N_2972,N_2050,N_2341);
and U2973 (N_2973,N_2485,N_2433);
nand U2974 (N_2974,N_2239,N_2393);
nor U2975 (N_2975,N_2044,N_2413);
and U2976 (N_2976,N_2255,N_2484);
or U2977 (N_2977,N_2142,N_2218);
nand U2978 (N_2978,N_2371,N_2085);
xnor U2979 (N_2979,N_2258,N_2208);
or U2980 (N_2980,N_2492,N_2273);
nand U2981 (N_2981,N_2412,N_2433);
nor U2982 (N_2982,N_2029,N_2106);
and U2983 (N_2983,N_2040,N_2115);
or U2984 (N_2984,N_2190,N_2125);
and U2985 (N_2985,N_2244,N_2000);
nor U2986 (N_2986,N_2412,N_2004);
nor U2987 (N_2987,N_2034,N_2393);
xor U2988 (N_2988,N_2142,N_2262);
nor U2989 (N_2989,N_2363,N_2478);
nor U2990 (N_2990,N_2343,N_2435);
nor U2991 (N_2991,N_2110,N_2402);
xnor U2992 (N_2992,N_2069,N_2156);
nand U2993 (N_2993,N_2348,N_2407);
nor U2994 (N_2994,N_2229,N_2290);
or U2995 (N_2995,N_2160,N_2444);
or U2996 (N_2996,N_2340,N_2219);
xnor U2997 (N_2997,N_2321,N_2147);
and U2998 (N_2998,N_2279,N_2145);
nor U2999 (N_2999,N_2237,N_2289);
nor U3000 (N_3000,N_2900,N_2662);
nand U3001 (N_3001,N_2548,N_2695);
nor U3002 (N_3002,N_2868,N_2941);
xor U3003 (N_3003,N_2894,N_2613);
and U3004 (N_3004,N_2607,N_2996);
nand U3005 (N_3005,N_2698,N_2534);
xor U3006 (N_3006,N_2539,N_2925);
or U3007 (N_3007,N_2656,N_2988);
and U3008 (N_3008,N_2778,N_2835);
or U3009 (N_3009,N_2571,N_2943);
nand U3010 (N_3010,N_2696,N_2545);
and U3011 (N_3011,N_2816,N_2886);
xnor U3012 (N_3012,N_2509,N_2744);
xnor U3013 (N_3013,N_2679,N_2960);
nor U3014 (N_3014,N_2724,N_2635);
nand U3015 (N_3015,N_2851,N_2917);
nor U3016 (N_3016,N_2985,N_2689);
xor U3017 (N_3017,N_2750,N_2508);
xnor U3018 (N_3018,N_2947,N_2617);
nor U3019 (N_3019,N_2991,N_2549);
and U3020 (N_3020,N_2809,N_2659);
nand U3021 (N_3021,N_2898,N_2680);
xnor U3022 (N_3022,N_2570,N_2560);
and U3023 (N_3023,N_2653,N_2939);
or U3024 (N_3024,N_2970,N_2675);
xnor U3025 (N_3025,N_2623,N_2528);
nor U3026 (N_3026,N_2830,N_2780);
or U3027 (N_3027,N_2628,N_2682);
or U3028 (N_3028,N_2507,N_2741);
and U3029 (N_3029,N_2688,N_2606);
or U3030 (N_3030,N_2621,N_2903);
nand U3031 (N_3031,N_2657,N_2832);
and U3032 (N_3032,N_2614,N_2998);
nand U3033 (N_3033,N_2702,N_2500);
xor U3034 (N_3034,N_2919,N_2537);
and U3035 (N_3035,N_2586,N_2541);
xor U3036 (N_3036,N_2928,N_2801);
nand U3037 (N_3037,N_2740,N_2746);
xnor U3038 (N_3038,N_2683,N_2701);
nor U3039 (N_3039,N_2874,N_2933);
xnor U3040 (N_3040,N_2557,N_2823);
and U3041 (N_3041,N_2561,N_2986);
and U3042 (N_3042,N_2805,N_2692);
or U3043 (N_3043,N_2803,N_2978);
nor U3044 (N_3044,N_2544,N_2578);
and U3045 (N_3045,N_2754,N_2833);
nand U3046 (N_3046,N_2799,N_2736);
or U3047 (N_3047,N_2759,N_2784);
or U3048 (N_3048,N_2515,N_2580);
and U3049 (N_3049,N_2971,N_2820);
nand U3050 (N_3050,N_2829,N_2665);
xnor U3051 (N_3051,N_2625,N_2834);
or U3052 (N_3052,N_2983,N_2739);
or U3053 (N_3053,N_2718,N_2556);
or U3054 (N_3054,N_2536,N_2563);
nand U3055 (N_3055,N_2768,N_2576);
and U3056 (N_3056,N_2569,N_2655);
or U3057 (N_3057,N_2639,N_2938);
and U3058 (N_3058,N_2620,N_2647);
and U3059 (N_3059,N_2891,N_2566);
nor U3060 (N_3060,N_2912,N_2822);
or U3061 (N_3061,N_2796,N_2574);
or U3062 (N_3062,N_2645,N_2824);
nand U3063 (N_3063,N_2913,N_2538);
nand U3064 (N_3064,N_2650,N_2989);
nand U3065 (N_3065,N_2932,N_2685);
and U3066 (N_3066,N_2715,N_2846);
nand U3067 (N_3067,N_2866,N_2742);
xor U3068 (N_3068,N_2853,N_2520);
or U3069 (N_3069,N_2860,N_2731);
nor U3070 (N_3070,N_2981,N_2961);
and U3071 (N_3071,N_2764,N_2783);
xnor U3072 (N_3072,N_2624,N_2703);
or U3073 (N_3073,N_2711,N_2871);
xor U3074 (N_3074,N_2940,N_2974);
and U3075 (N_3075,N_2502,N_2747);
and U3076 (N_3076,N_2717,N_2864);
xnor U3077 (N_3077,N_2890,N_2707);
xnor U3078 (N_3078,N_2564,N_2812);
nand U3079 (N_3079,N_2806,N_2920);
nor U3080 (N_3080,N_2562,N_2770);
and U3081 (N_3081,N_2734,N_2963);
nor U3082 (N_3082,N_2510,N_2957);
nand U3083 (N_3083,N_2831,N_2777);
or U3084 (N_3084,N_2849,N_2543);
nor U3085 (N_3085,N_2579,N_2622);
xnor U3086 (N_3086,N_2771,N_2969);
and U3087 (N_3087,N_2687,N_2880);
xor U3088 (N_3088,N_2787,N_2524);
and U3089 (N_3089,N_2547,N_2686);
nand U3090 (N_3090,N_2842,N_2899);
nor U3091 (N_3091,N_2700,N_2902);
and U3092 (N_3092,N_2859,N_2632);
or U3093 (N_3093,N_2513,N_2504);
and U3094 (N_3094,N_2881,N_2959);
nor U3095 (N_3095,N_2888,N_2755);
or U3096 (N_3096,N_2792,N_2758);
or U3097 (N_3097,N_2611,N_2914);
and U3098 (N_3098,N_2918,N_2877);
and U3099 (N_3099,N_2522,N_2559);
nand U3100 (N_3100,N_2637,N_2942);
xor U3101 (N_3101,N_2808,N_2814);
or U3102 (N_3102,N_2760,N_2964);
xnor U3103 (N_3103,N_2530,N_2885);
nand U3104 (N_3104,N_2945,N_2668);
and U3105 (N_3105,N_2529,N_2767);
xor U3106 (N_3106,N_2503,N_2514);
xnor U3107 (N_3107,N_2554,N_2798);
and U3108 (N_3108,N_2827,N_2521);
xor U3109 (N_3109,N_2568,N_2631);
and U3110 (N_3110,N_2870,N_2525);
xor U3111 (N_3111,N_2616,N_2793);
and U3112 (N_3112,N_2732,N_2555);
or U3113 (N_3113,N_2729,N_2934);
or U3114 (N_3114,N_2879,N_2838);
or U3115 (N_3115,N_2592,N_2896);
nor U3116 (N_3116,N_2716,N_2511);
and U3117 (N_3117,N_2876,N_2714);
nor U3118 (N_3118,N_2723,N_2597);
and U3119 (N_3119,N_2818,N_2905);
or U3120 (N_3120,N_2994,N_2911);
nor U3121 (N_3121,N_2709,N_2922);
nor U3122 (N_3122,N_2762,N_2519);
nor U3123 (N_3123,N_2980,N_2646);
nand U3124 (N_3124,N_2882,N_2836);
nand U3125 (N_3125,N_2769,N_2800);
nand U3126 (N_3126,N_2674,N_2861);
xor U3127 (N_3127,N_2641,N_2855);
and U3128 (N_3128,N_2648,N_2550);
nand U3129 (N_3129,N_2946,N_2847);
and U3130 (N_3130,N_2588,N_2869);
and U3131 (N_3131,N_2710,N_2501);
nand U3132 (N_3132,N_2526,N_2889);
nor U3133 (N_3133,N_2585,N_2825);
nand U3134 (N_3134,N_2813,N_2952);
nor U3135 (N_3135,N_2766,N_2531);
nand U3136 (N_3136,N_2897,N_2591);
nor U3137 (N_3137,N_2671,N_2927);
and U3138 (N_3138,N_2841,N_2713);
and U3139 (N_3139,N_2745,N_2542);
nor U3140 (N_3140,N_2527,N_2708);
and U3141 (N_3141,N_2733,N_2582);
nand U3142 (N_3142,N_2773,N_2596);
and U3143 (N_3143,N_2977,N_2546);
or U3144 (N_3144,N_2552,N_2909);
and U3145 (N_3145,N_2765,N_2763);
or U3146 (N_3146,N_2979,N_2958);
xor U3147 (N_3147,N_2779,N_2738);
nor U3148 (N_3148,N_2601,N_2856);
and U3149 (N_3149,N_2517,N_2791);
and U3150 (N_3150,N_2693,N_2790);
xor U3151 (N_3151,N_2776,N_2644);
nor U3152 (N_3152,N_2603,N_2844);
xor U3153 (N_3153,N_2600,N_2667);
nor U3154 (N_3154,N_2752,N_2727);
or U3155 (N_3155,N_2862,N_2984);
and U3156 (N_3156,N_2577,N_2987);
and U3157 (N_3157,N_2982,N_2719);
nor U3158 (N_3158,N_2908,N_2930);
or U3159 (N_3159,N_2737,N_2664);
xnor U3160 (N_3160,N_2730,N_2815);
and U3161 (N_3161,N_2948,N_2951);
nor U3162 (N_3162,N_2962,N_2873);
xnor U3163 (N_3163,N_2904,N_2867);
or U3164 (N_3164,N_2751,N_2627);
xor U3165 (N_3165,N_2781,N_2619);
or U3166 (N_3166,N_2558,N_2772);
nand U3167 (N_3167,N_2807,N_2992);
or U3168 (N_3168,N_2895,N_2512);
nand U3169 (N_3169,N_2540,N_2610);
xnor U3170 (N_3170,N_2626,N_2567);
xnor U3171 (N_3171,N_2965,N_2720);
xnor U3172 (N_3172,N_2923,N_2663);
or U3173 (N_3173,N_2921,N_2581);
xor U3174 (N_3174,N_2972,N_2735);
nor U3175 (N_3175,N_2535,N_2699);
or U3176 (N_3176,N_2975,N_2804);
nand U3177 (N_3177,N_2936,N_2743);
nand U3178 (N_3178,N_2937,N_2795);
and U3179 (N_3179,N_2602,N_2997);
nand U3180 (N_3180,N_2875,N_2629);
or U3181 (N_3181,N_2761,N_2518);
nand U3182 (N_3182,N_2848,N_2872);
and U3183 (N_3183,N_2666,N_2660);
xor U3184 (N_3184,N_2915,N_2649);
nand U3185 (N_3185,N_2583,N_2797);
xnor U3186 (N_3186,N_2852,N_2609);
nand U3187 (N_3187,N_2676,N_2929);
nor U3188 (N_3188,N_2658,N_2651);
nor U3189 (N_3189,N_2533,N_2990);
and U3190 (N_3190,N_2669,N_2785);
and U3191 (N_3191,N_2594,N_2633);
and U3192 (N_3192,N_2906,N_2976);
nand U3193 (N_3193,N_2843,N_2817);
nand U3194 (N_3194,N_2995,N_2892);
xor U3195 (N_3195,N_2722,N_2893);
or U3196 (N_3196,N_2678,N_2523);
and U3197 (N_3197,N_2757,N_2608);
xor U3198 (N_3198,N_2910,N_2725);
nor U3199 (N_3199,N_2950,N_2863);
xor U3200 (N_3200,N_2599,N_2949);
xnor U3201 (N_3201,N_2704,N_2774);
xor U3202 (N_3202,N_2630,N_2684);
and U3203 (N_3203,N_2967,N_2821);
or U3204 (N_3204,N_2640,N_2907);
nor U3205 (N_3205,N_2954,N_2670);
nand U3206 (N_3206,N_2505,N_2595);
or U3207 (N_3207,N_2584,N_2677);
xor U3208 (N_3208,N_2901,N_2944);
xor U3209 (N_3209,N_2916,N_2794);
nor U3210 (N_3210,N_2782,N_2589);
xnor U3211 (N_3211,N_2721,N_2955);
and U3212 (N_3212,N_2672,N_2605);
or U3213 (N_3213,N_2748,N_2612);
nand U3214 (N_3214,N_2697,N_2999);
or U3215 (N_3215,N_2618,N_2705);
xor U3216 (N_3216,N_2615,N_2865);
xor U3217 (N_3217,N_2786,N_2673);
and U3218 (N_3218,N_2850,N_2837);
nor U3219 (N_3219,N_2706,N_2652);
xor U3220 (N_3220,N_2802,N_2638);
nor U3221 (N_3221,N_2572,N_2828);
and U3222 (N_3222,N_2532,N_2966);
nor U3223 (N_3223,N_2883,N_2642);
and U3224 (N_3224,N_2840,N_2553);
xnor U3225 (N_3225,N_2924,N_2884);
nand U3226 (N_3226,N_2775,N_2973);
xor U3227 (N_3227,N_2598,N_2956);
xor U3228 (N_3228,N_2636,N_2749);
nand U3229 (N_3229,N_2845,N_2935);
or U3230 (N_3230,N_2728,N_2931);
or U3231 (N_3231,N_2593,N_2604);
xnor U3232 (N_3232,N_2858,N_2691);
and U3233 (N_3233,N_2826,N_2839);
nor U3234 (N_3234,N_2565,N_2661);
and U3235 (N_3235,N_2506,N_2993);
nand U3236 (N_3236,N_2690,N_2590);
or U3237 (N_3237,N_2819,N_2634);
and U3238 (N_3238,N_2968,N_2878);
nand U3239 (N_3239,N_2681,N_2643);
or U3240 (N_3240,N_2516,N_2575);
or U3241 (N_3241,N_2926,N_2810);
or U3242 (N_3242,N_2788,N_2953);
nor U3243 (N_3243,N_2654,N_2587);
nor U3244 (N_3244,N_2789,N_2753);
and U3245 (N_3245,N_2811,N_2854);
or U3246 (N_3246,N_2756,N_2551);
xor U3247 (N_3247,N_2726,N_2712);
nand U3248 (N_3248,N_2694,N_2573);
and U3249 (N_3249,N_2857,N_2887);
and U3250 (N_3250,N_2962,N_2603);
and U3251 (N_3251,N_2672,N_2888);
xnor U3252 (N_3252,N_2523,N_2668);
or U3253 (N_3253,N_2511,N_2639);
and U3254 (N_3254,N_2745,N_2566);
and U3255 (N_3255,N_2582,N_2806);
and U3256 (N_3256,N_2651,N_2701);
nand U3257 (N_3257,N_2794,N_2791);
nand U3258 (N_3258,N_2775,N_2979);
nand U3259 (N_3259,N_2509,N_2536);
xor U3260 (N_3260,N_2788,N_2747);
nand U3261 (N_3261,N_2656,N_2973);
nor U3262 (N_3262,N_2548,N_2931);
nand U3263 (N_3263,N_2703,N_2700);
or U3264 (N_3264,N_2723,N_2501);
or U3265 (N_3265,N_2890,N_2744);
or U3266 (N_3266,N_2532,N_2733);
nor U3267 (N_3267,N_2881,N_2834);
xnor U3268 (N_3268,N_2883,N_2670);
nand U3269 (N_3269,N_2874,N_2626);
xnor U3270 (N_3270,N_2749,N_2751);
nand U3271 (N_3271,N_2739,N_2527);
nor U3272 (N_3272,N_2686,N_2502);
xnor U3273 (N_3273,N_2708,N_2951);
xnor U3274 (N_3274,N_2622,N_2959);
or U3275 (N_3275,N_2950,N_2677);
or U3276 (N_3276,N_2893,N_2589);
or U3277 (N_3277,N_2540,N_2647);
nor U3278 (N_3278,N_2723,N_2653);
and U3279 (N_3279,N_2812,N_2994);
nand U3280 (N_3280,N_2628,N_2723);
xor U3281 (N_3281,N_2976,N_2998);
and U3282 (N_3282,N_2720,N_2504);
nand U3283 (N_3283,N_2596,N_2569);
nor U3284 (N_3284,N_2675,N_2540);
xor U3285 (N_3285,N_2652,N_2584);
and U3286 (N_3286,N_2515,N_2714);
nor U3287 (N_3287,N_2921,N_2657);
or U3288 (N_3288,N_2988,N_2745);
xnor U3289 (N_3289,N_2944,N_2856);
and U3290 (N_3290,N_2675,N_2941);
nor U3291 (N_3291,N_2856,N_2946);
xnor U3292 (N_3292,N_2774,N_2768);
nand U3293 (N_3293,N_2593,N_2811);
or U3294 (N_3294,N_2543,N_2812);
and U3295 (N_3295,N_2974,N_2933);
nand U3296 (N_3296,N_2766,N_2585);
nor U3297 (N_3297,N_2755,N_2897);
nand U3298 (N_3298,N_2748,N_2598);
xnor U3299 (N_3299,N_2516,N_2931);
and U3300 (N_3300,N_2867,N_2737);
and U3301 (N_3301,N_2873,N_2720);
nand U3302 (N_3302,N_2540,N_2746);
xnor U3303 (N_3303,N_2941,N_2900);
and U3304 (N_3304,N_2626,N_2797);
nor U3305 (N_3305,N_2816,N_2574);
or U3306 (N_3306,N_2914,N_2840);
and U3307 (N_3307,N_2968,N_2719);
and U3308 (N_3308,N_2574,N_2649);
or U3309 (N_3309,N_2704,N_2663);
or U3310 (N_3310,N_2585,N_2680);
and U3311 (N_3311,N_2710,N_2724);
nor U3312 (N_3312,N_2541,N_2519);
nor U3313 (N_3313,N_2768,N_2779);
nor U3314 (N_3314,N_2522,N_2643);
and U3315 (N_3315,N_2605,N_2670);
nand U3316 (N_3316,N_2848,N_2855);
nor U3317 (N_3317,N_2823,N_2665);
xnor U3318 (N_3318,N_2737,N_2505);
nand U3319 (N_3319,N_2962,N_2789);
nand U3320 (N_3320,N_2571,N_2762);
nor U3321 (N_3321,N_2762,N_2582);
nor U3322 (N_3322,N_2869,N_2795);
xor U3323 (N_3323,N_2815,N_2855);
or U3324 (N_3324,N_2733,N_2641);
and U3325 (N_3325,N_2873,N_2691);
and U3326 (N_3326,N_2943,N_2925);
and U3327 (N_3327,N_2615,N_2695);
xnor U3328 (N_3328,N_2755,N_2709);
nor U3329 (N_3329,N_2659,N_2938);
or U3330 (N_3330,N_2564,N_2802);
nor U3331 (N_3331,N_2551,N_2781);
or U3332 (N_3332,N_2659,N_2793);
or U3333 (N_3333,N_2707,N_2613);
nor U3334 (N_3334,N_2537,N_2983);
and U3335 (N_3335,N_2828,N_2550);
nand U3336 (N_3336,N_2687,N_2539);
xnor U3337 (N_3337,N_2804,N_2865);
nor U3338 (N_3338,N_2859,N_2875);
nor U3339 (N_3339,N_2562,N_2797);
nor U3340 (N_3340,N_2894,N_2791);
xnor U3341 (N_3341,N_2609,N_2640);
or U3342 (N_3342,N_2623,N_2610);
nand U3343 (N_3343,N_2638,N_2670);
nor U3344 (N_3344,N_2823,N_2529);
nor U3345 (N_3345,N_2839,N_2699);
nor U3346 (N_3346,N_2538,N_2636);
xnor U3347 (N_3347,N_2672,N_2688);
nor U3348 (N_3348,N_2971,N_2933);
nor U3349 (N_3349,N_2973,N_2903);
nand U3350 (N_3350,N_2672,N_2990);
and U3351 (N_3351,N_2840,N_2859);
nand U3352 (N_3352,N_2669,N_2956);
nor U3353 (N_3353,N_2696,N_2778);
nand U3354 (N_3354,N_2700,N_2827);
and U3355 (N_3355,N_2736,N_2714);
xnor U3356 (N_3356,N_2924,N_2661);
and U3357 (N_3357,N_2638,N_2945);
or U3358 (N_3358,N_2783,N_2811);
nand U3359 (N_3359,N_2612,N_2594);
or U3360 (N_3360,N_2822,N_2727);
nand U3361 (N_3361,N_2600,N_2639);
nand U3362 (N_3362,N_2500,N_2561);
and U3363 (N_3363,N_2655,N_2579);
or U3364 (N_3364,N_2826,N_2938);
or U3365 (N_3365,N_2680,N_2505);
nand U3366 (N_3366,N_2642,N_2770);
or U3367 (N_3367,N_2989,N_2586);
nand U3368 (N_3368,N_2963,N_2517);
xnor U3369 (N_3369,N_2525,N_2841);
and U3370 (N_3370,N_2960,N_2943);
and U3371 (N_3371,N_2682,N_2644);
nor U3372 (N_3372,N_2555,N_2680);
nand U3373 (N_3373,N_2534,N_2919);
and U3374 (N_3374,N_2978,N_2930);
nand U3375 (N_3375,N_2552,N_2738);
nand U3376 (N_3376,N_2856,N_2656);
or U3377 (N_3377,N_2952,N_2739);
or U3378 (N_3378,N_2529,N_2703);
xor U3379 (N_3379,N_2976,N_2578);
nor U3380 (N_3380,N_2964,N_2927);
nor U3381 (N_3381,N_2877,N_2615);
and U3382 (N_3382,N_2773,N_2942);
nand U3383 (N_3383,N_2961,N_2831);
nor U3384 (N_3384,N_2865,N_2939);
nand U3385 (N_3385,N_2933,N_2695);
nand U3386 (N_3386,N_2735,N_2865);
nor U3387 (N_3387,N_2714,N_2579);
nand U3388 (N_3388,N_2557,N_2648);
or U3389 (N_3389,N_2506,N_2720);
nand U3390 (N_3390,N_2890,N_2814);
and U3391 (N_3391,N_2679,N_2835);
or U3392 (N_3392,N_2574,N_2576);
xor U3393 (N_3393,N_2851,N_2945);
nor U3394 (N_3394,N_2869,N_2754);
nand U3395 (N_3395,N_2512,N_2804);
and U3396 (N_3396,N_2882,N_2748);
or U3397 (N_3397,N_2853,N_2692);
nor U3398 (N_3398,N_2727,N_2940);
xnor U3399 (N_3399,N_2734,N_2754);
nor U3400 (N_3400,N_2551,N_2625);
or U3401 (N_3401,N_2568,N_2518);
and U3402 (N_3402,N_2597,N_2588);
or U3403 (N_3403,N_2584,N_2819);
nor U3404 (N_3404,N_2777,N_2911);
and U3405 (N_3405,N_2843,N_2758);
nand U3406 (N_3406,N_2842,N_2534);
nor U3407 (N_3407,N_2996,N_2815);
xnor U3408 (N_3408,N_2985,N_2619);
or U3409 (N_3409,N_2618,N_2787);
nor U3410 (N_3410,N_2525,N_2880);
nor U3411 (N_3411,N_2913,N_2943);
nand U3412 (N_3412,N_2778,N_2573);
nand U3413 (N_3413,N_2585,N_2580);
nand U3414 (N_3414,N_2798,N_2618);
nand U3415 (N_3415,N_2901,N_2631);
nand U3416 (N_3416,N_2851,N_2782);
xnor U3417 (N_3417,N_2808,N_2643);
and U3418 (N_3418,N_2809,N_2734);
xor U3419 (N_3419,N_2513,N_2713);
nand U3420 (N_3420,N_2770,N_2644);
nand U3421 (N_3421,N_2601,N_2884);
xnor U3422 (N_3422,N_2800,N_2814);
and U3423 (N_3423,N_2898,N_2619);
nand U3424 (N_3424,N_2771,N_2932);
xnor U3425 (N_3425,N_2752,N_2837);
nand U3426 (N_3426,N_2801,N_2854);
xor U3427 (N_3427,N_2959,N_2692);
and U3428 (N_3428,N_2501,N_2812);
or U3429 (N_3429,N_2714,N_2529);
nor U3430 (N_3430,N_2807,N_2664);
and U3431 (N_3431,N_2897,N_2982);
nor U3432 (N_3432,N_2784,N_2505);
xnor U3433 (N_3433,N_2814,N_2945);
xnor U3434 (N_3434,N_2775,N_2839);
or U3435 (N_3435,N_2809,N_2644);
or U3436 (N_3436,N_2625,N_2544);
nor U3437 (N_3437,N_2678,N_2553);
nand U3438 (N_3438,N_2534,N_2961);
nor U3439 (N_3439,N_2694,N_2636);
or U3440 (N_3440,N_2645,N_2777);
xnor U3441 (N_3441,N_2876,N_2604);
nand U3442 (N_3442,N_2697,N_2818);
xnor U3443 (N_3443,N_2754,N_2577);
or U3444 (N_3444,N_2640,N_2727);
xnor U3445 (N_3445,N_2760,N_2726);
or U3446 (N_3446,N_2906,N_2787);
nand U3447 (N_3447,N_2732,N_2592);
nand U3448 (N_3448,N_2658,N_2876);
and U3449 (N_3449,N_2752,N_2942);
xor U3450 (N_3450,N_2624,N_2515);
and U3451 (N_3451,N_2819,N_2594);
or U3452 (N_3452,N_2959,N_2921);
or U3453 (N_3453,N_2976,N_2982);
or U3454 (N_3454,N_2561,N_2562);
and U3455 (N_3455,N_2986,N_2743);
and U3456 (N_3456,N_2764,N_2578);
nand U3457 (N_3457,N_2659,N_2736);
nor U3458 (N_3458,N_2663,N_2913);
or U3459 (N_3459,N_2853,N_2869);
nand U3460 (N_3460,N_2869,N_2779);
xor U3461 (N_3461,N_2773,N_2885);
xor U3462 (N_3462,N_2803,N_2991);
xor U3463 (N_3463,N_2910,N_2559);
nand U3464 (N_3464,N_2657,N_2872);
and U3465 (N_3465,N_2536,N_2548);
and U3466 (N_3466,N_2930,N_2919);
xnor U3467 (N_3467,N_2805,N_2968);
xor U3468 (N_3468,N_2973,N_2501);
and U3469 (N_3469,N_2856,N_2928);
or U3470 (N_3470,N_2731,N_2726);
nor U3471 (N_3471,N_2865,N_2612);
xor U3472 (N_3472,N_2973,N_2598);
or U3473 (N_3473,N_2599,N_2604);
nor U3474 (N_3474,N_2813,N_2769);
xor U3475 (N_3475,N_2537,N_2610);
nor U3476 (N_3476,N_2626,N_2963);
or U3477 (N_3477,N_2707,N_2761);
nor U3478 (N_3478,N_2697,N_2715);
and U3479 (N_3479,N_2596,N_2792);
and U3480 (N_3480,N_2909,N_2771);
nand U3481 (N_3481,N_2943,N_2964);
or U3482 (N_3482,N_2717,N_2584);
nor U3483 (N_3483,N_2590,N_2748);
or U3484 (N_3484,N_2545,N_2774);
xnor U3485 (N_3485,N_2829,N_2983);
or U3486 (N_3486,N_2741,N_2661);
or U3487 (N_3487,N_2669,N_2623);
nand U3488 (N_3488,N_2754,N_2920);
nor U3489 (N_3489,N_2802,N_2819);
nand U3490 (N_3490,N_2924,N_2668);
nand U3491 (N_3491,N_2988,N_2814);
nor U3492 (N_3492,N_2548,N_2855);
nand U3493 (N_3493,N_2521,N_2552);
or U3494 (N_3494,N_2786,N_2808);
nand U3495 (N_3495,N_2541,N_2714);
xnor U3496 (N_3496,N_2808,N_2968);
nor U3497 (N_3497,N_2511,N_2584);
xnor U3498 (N_3498,N_2549,N_2882);
nor U3499 (N_3499,N_2509,N_2880);
nor U3500 (N_3500,N_3484,N_3494);
or U3501 (N_3501,N_3089,N_3443);
nor U3502 (N_3502,N_3096,N_3265);
nor U3503 (N_3503,N_3223,N_3319);
nor U3504 (N_3504,N_3025,N_3182);
nand U3505 (N_3505,N_3134,N_3106);
or U3506 (N_3506,N_3444,N_3253);
nor U3507 (N_3507,N_3216,N_3100);
or U3508 (N_3508,N_3272,N_3151);
xor U3509 (N_3509,N_3120,N_3206);
and U3510 (N_3510,N_3191,N_3353);
xor U3511 (N_3511,N_3233,N_3424);
and U3512 (N_3512,N_3304,N_3413);
nand U3513 (N_3513,N_3465,N_3244);
nor U3514 (N_3514,N_3167,N_3333);
xnor U3515 (N_3515,N_3455,N_3072);
xor U3516 (N_3516,N_3458,N_3242);
nand U3517 (N_3517,N_3094,N_3175);
or U3518 (N_3518,N_3129,N_3160);
nand U3519 (N_3519,N_3247,N_3358);
nand U3520 (N_3520,N_3491,N_3267);
and U3521 (N_3521,N_3020,N_3483);
nand U3522 (N_3522,N_3044,N_3186);
xnor U3523 (N_3523,N_3325,N_3318);
xor U3524 (N_3524,N_3012,N_3021);
xor U3525 (N_3525,N_3158,N_3260);
and U3526 (N_3526,N_3196,N_3497);
nand U3527 (N_3527,N_3124,N_3212);
xor U3528 (N_3528,N_3097,N_3102);
and U3529 (N_3529,N_3306,N_3155);
and U3530 (N_3530,N_3084,N_3150);
and U3531 (N_3531,N_3329,N_3429);
nor U3532 (N_3532,N_3022,N_3049);
xor U3533 (N_3533,N_3245,N_3467);
xnor U3534 (N_3534,N_3009,N_3268);
xor U3535 (N_3535,N_3093,N_3074);
xnor U3536 (N_3536,N_3101,N_3468);
and U3537 (N_3537,N_3349,N_3414);
nor U3538 (N_3538,N_3449,N_3019);
nand U3539 (N_3539,N_3108,N_3143);
xor U3540 (N_3540,N_3411,N_3248);
xor U3541 (N_3541,N_3230,N_3461);
and U3542 (N_3542,N_3313,N_3017);
xnor U3543 (N_3543,N_3382,N_3371);
nand U3544 (N_3544,N_3261,N_3237);
nor U3545 (N_3545,N_3092,N_3126);
nor U3546 (N_3546,N_3477,N_3390);
nand U3547 (N_3547,N_3345,N_3067);
nor U3548 (N_3548,N_3128,N_3117);
nand U3549 (N_3549,N_3396,N_3460);
and U3550 (N_3550,N_3194,N_3352);
nor U3551 (N_3551,N_3190,N_3193);
or U3552 (N_3552,N_3399,N_3082);
or U3553 (N_3553,N_3023,N_3278);
nor U3554 (N_3554,N_3170,N_3273);
nand U3555 (N_3555,N_3290,N_3401);
xnor U3556 (N_3556,N_3240,N_3213);
nand U3557 (N_3557,N_3116,N_3320);
or U3558 (N_3558,N_3373,N_3033);
or U3559 (N_3559,N_3346,N_3400);
nor U3560 (N_3560,N_3149,N_3381);
and U3561 (N_3561,N_3380,N_3115);
xor U3562 (N_3562,N_3447,N_3252);
xor U3563 (N_3563,N_3328,N_3109);
nand U3564 (N_3564,N_3215,N_3470);
xnor U3565 (N_3565,N_3301,N_3254);
or U3566 (N_3566,N_3251,N_3030);
xor U3567 (N_3567,N_3422,N_3466);
nand U3568 (N_3568,N_3255,N_3479);
nand U3569 (N_3569,N_3492,N_3003);
or U3570 (N_3570,N_3331,N_3065);
and U3571 (N_3571,N_3433,N_3457);
xnor U3572 (N_3572,N_3173,N_3428);
or U3573 (N_3573,N_3256,N_3369);
nand U3574 (N_3574,N_3407,N_3241);
xor U3575 (N_3575,N_3047,N_3452);
or U3576 (N_3576,N_3176,N_3309);
or U3577 (N_3577,N_3259,N_3419);
nor U3578 (N_3578,N_3060,N_3192);
xor U3579 (N_3579,N_3168,N_3282);
and U3580 (N_3580,N_3051,N_3359);
and U3581 (N_3581,N_3499,N_3264);
xor U3582 (N_3582,N_3350,N_3037);
xnor U3583 (N_3583,N_3222,N_3184);
xor U3584 (N_3584,N_3263,N_3078);
or U3585 (N_3585,N_3360,N_3229);
nor U3586 (N_3586,N_3425,N_3163);
or U3587 (N_3587,N_3316,N_3276);
nand U3588 (N_3588,N_3062,N_3362);
nand U3589 (N_3589,N_3388,N_3148);
xnor U3590 (N_3590,N_3364,N_3228);
nor U3591 (N_3591,N_3383,N_3099);
or U3592 (N_3592,N_3481,N_3081);
xor U3593 (N_3593,N_3180,N_3462);
and U3594 (N_3594,N_3187,N_3157);
nor U3595 (N_3595,N_3498,N_3001);
nand U3596 (N_3596,N_3493,N_3339);
xnor U3597 (N_3597,N_3410,N_3136);
nand U3598 (N_3598,N_3367,N_3057);
nor U3599 (N_3599,N_3321,N_3225);
and U3600 (N_3600,N_3415,N_3405);
or U3601 (N_3601,N_3010,N_3324);
nand U3602 (N_3602,N_3370,N_3139);
xnor U3603 (N_3603,N_3008,N_3006);
nor U3604 (N_3604,N_3298,N_3137);
nand U3605 (N_3605,N_3398,N_3342);
and U3606 (N_3606,N_3469,N_3035);
and U3607 (N_3607,N_3351,N_3127);
and U3608 (N_3608,N_3208,N_3050);
nand U3609 (N_3609,N_3039,N_3210);
nand U3610 (N_3610,N_3327,N_3275);
nand U3611 (N_3611,N_3473,N_3283);
xor U3612 (N_3612,N_3292,N_3404);
nand U3613 (N_3613,N_3437,N_3271);
nand U3614 (N_3614,N_3418,N_3357);
or U3615 (N_3615,N_3323,N_3201);
nand U3616 (N_3616,N_3392,N_3438);
and U3617 (N_3617,N_3376,N_3207);
or U3618 (N_3618,N_3317,N_3337);
and U3619 (N_3619,N_3071,N_3294);
and U3620 (N_3620,N_3152,N_3475);
nor U3621 (N_3621,N_3027,N_3036);
and U3622 (N_3622,N_3188,N_3123);
or U3623 (N_3623,N_3164,N_3490);
or U3624 (N_3624,N_3159,N_3053);
xor U3625 (N_3625,N_3083,N_3246);
and U3626 (N_3626,N_3463,N_3250);
nor U3627 (N_3627,N_3054,N_3204);
nand U3628 (N_3628,N_3355,N_3073);
xnor U3629 (N_3629,N_3007,N_3013);
nor U3630 (N_3630,N_3436,N_3077);
nor U3631 (N_3631,N_3041,N_3393);
and U3632 (N_3632,N_3420,N_3121);
nor U3633 (N_3633,N_3293,N_3385);
nor U3634 (N_3634,N_3430,N_3202);
nor U3635 (N_3635,N_3091,N_3387);
or U3636 (N_3636,N_3166,N_3028);
nand U3637 (N_3637,N_3487,N_3311);
and U3638 (N_3638,N_3029,N_3200);
or U3639 (N_3639,N_3421,N_3131);
nand U3640 (N_3640,N_3257,N_3431);
and U3641 (N_3641,N_3079,N_3052);
nand U3642 (N_3642,N_3114,N_3238);
nand U3643 (N_3643,N_3464,N_3478);
nand U3644 (N_3644,N_3334,N_3243);
and U3645 (N_3645,N_3090,N_3075);
and U3646 (N_3646,N_3231,N_3434);
or U3647 (N_3647,N_3177,N_3235);
nor U3648 (N_3648,N_3219,N_3482);
xnor U3649 (N_3649,N_3132,N_3289);
or U3650 (N_3650,N_3338,N_3226);
or U3651 (N_3651,N_3227,N_3441);
nand U3652 (N_3652,N_3295,N_3002);
and U3653 (N_3653,N_3277,N_3379);
or U3654 (N_3654,N_3336,N_3171);
nor U3655 (N_3655,N_3104,N_3066);
xor U3656 (N_3656,N_3386,N_3209);
and U3657 (N_3657,N_3474,N_3119);
or U3658 (N_3658,N_3377,N_3061);
xnor U3659 (N_3659,N_3394,N_3111);
nor U3660 (N_3660,N_3000,N_3332);
nor U3661 (N_3661,N_3144,N_3423);
or U3662 (N_3662,N_3140,N_3107);
nor U3663 (N_3663,N_3105,N_3284);
nand U3664 (N_3664,N_3146,N_3085);
and U3665 (N_3665,N_3195,N_3004);
and U3666 (N_3666,N_3281,N_3296);
or U3667 (N_3667,N_3486,N_3403);
xor U3668 (N_3668,N_3417,N_3312);
and U3669 (N_3669,N_3068,N_3450);
nand U3670 (N_3670,N_3055,N_3198);
xnor U3671 (N_3671,N_3305,N_3395);
nor U3672 (N_3672,N_3118,N_3011);
nor U3673 (N_3673,N_3234,N_3310);
nor U3674 (N_3674,N_3174,N_3203);
xnor U3675 (N_3675,N_3014,N_3300);
nand U3676 (N_3676,N_3286,N_3368);
or U3677 (N_3677,N_3453,N_3070);
xnor U3678 (N_3678,N_3489,N_3239);
and U3679 (N_3679,N_3031,N_3348);
or U3680 (N_3680,N_3125,N_3064);
xor U3681 (N_3681,N_3375,N_3232);
xnor U3682 (N_3682,N_3005,N_3183);
or U3683 (N_3683,N_3416,N_3406);
nand U3684 (N_3684,N_3297,N_3042);
nor U3685 (N_3685,N_3220,N_3427);
or U3686 (N_3686,N_3480,N_3291);
xnor U3687 (N_3687,N_3221,N_3162);
nor U3688 (N_3688,N_3145,N_3056);
nand U3689 (N_3689,N_3038,N_3446);
nand U3690 (N_3690,N_3409,N_3307);
xnor U3691 (N_3691,N_3326,N_3076);
xnor U3692 (N_3692,N_3361,N_3026);
or U3693 (N_3693,N_3363,N_3269);
xor U3694 (N_3694,N_3165,N_3389);
xor U3695 (N_3695,N_3347,N_3408);
nand U3696 (N_3696,N_3258,N_3315);
nand U3697 (N_3697,N_3156,N_3032);
and U3698 (N_3698,N_3189,N_3185);
nor U3699 (N_3699,N_3302,N_3043);
or U3700 (N_3700,N_3288,N_3374);
or U3701 (N_3701,N_3112,N_3397);
xnor U3702 (N_3702,N_3426,N_3384);
xor U3703 (N_3703,N_3322,N_3459);
and U3704 (N_3704,N_3154,N_3147);
xor U3705 (N_3705,N_3016,N_3135);
xnor U3706 (N_3706,N_3314,N_3451);
nand U3707 (N_3707,N_3341,N_3356);
nand U3708 (N_3708,N_3199,N_3365);
xor U3709 (N_3709,N_3113,N_3045);
nand U3710 (N_3710,N_3303,N_3080);
nand U3711 (N_3711,N_3495,N_3161);
xnor U3712 (N_3712,N_3412,N_3103);
nand U3713 (N_3713,N_3391,N_3448);
or U3714 (N_3714,N_3432,N_3340);
nor U3715 (N_3715,N_3088,N_3435);
nor U3716 (N_3716,N_3217,N_3285);
nand U3717 (N_3717,N_3059,N_3040);
nor U3718 (N_3718,N_3330,N_3205);
xnor U3719 (N_3719,N_3485,N_3471);
xnor U3720 (N_3720,N_3372,N_3476);
or U3721 (N_3721,N_3046,N_3344);
or U3722 (N_3722,N_3058,N_3274);
nor U3723 (N_3723,N_3454,N_3249);
nand U3724 (N_3724,N_3018,N_3308);
or U3725 (N_3725,N_3442,N_3110);
nand U3726 (N_3726,N_3141,N_3402);
nor U3727 (N_3727,N_3095,N_3335);
nor U3728 (N_3728,N_3197,N_3024);
xnor U3729 (N_3729,N_3133,N_3279);
and U3730 (N_3730,N_3280,N_3287);
nand U3731 (N_3731,N_3472,N_3378);
or U3732 (N_3732,N_3266,N_3138);
and U3733 (N_3733,N_3069,N_3178);
and U3734 (N_3734,N_3086,N_3343);
nand U3735 (N_3735,N_3181,N_3439);
nand U3736 (N_3736,N_3063,N_3236);
nor U3737 (N_3737,N_3122,N_3034);
nor U3738 (N_3738,N_3169,N_3048);
or U3739 (N_3739,N_3354,N_3440);
or U3740 (N_3740,N_3262,N_3179);
nor U3741 (N_3741,N_3299,N_3211);
nand U3742 (N_3742,N_3098,N_3456);
nor U3743 (N_3743,N_3214,N_3130);
nand U3744 (N_3744,N_3488,N_3218);
or U3745 (N_3745,N_3496,N_3172);
nor U3746 (N_3746,N_3270,N_3142);
or U3747 (N_3747,N_3366,N_3153);
nor U3748 (N_3748,N_3445,N_3087);
xnor U3749 (N_3749,N_3015,N_3224);
nor U3750 (N_3750,N_3251,N_3204);
or U3751 (N_3751,N_3242,N_3146);
nand U3752 (N_3752,N_3159,N_3419);
nor U3753 (N_3753,N_3102,N_3021);
xnor U3754 (N_3754,N_3314,N_3002);
and U3755 (N_3755,N_3264,N_3422);
nand U3756 (N_3756,N_3285,N_3202);
and U3757 (N_3757,N_3471,N_3131);
nand U3758 (N_3758,N_3356,N_3195);
and U3759 (N_3759,N_3425,N_3421);
xnor U3760 (N_3760,N_3461,N_3440);
nand U3761 (N_3761,N_3429,N_3002);
nand U3762 (N_3762,N_3411,N_3146);
nor U3763 (N_3763,N_3312,N_3170);
nand U3764 (N_3764,N_3220,N_3160);
nor U3765 (N_3765,N_3180,N_3382);
xor U3766 (N_3766,N_3413,N_3482);
xor U3767 (N_3767,N_3180,N_3224);
nor U3768 (N_3768,N_3415,N_3278);
nor U3769 (N_3769,N_3339,N_3341);
nor U3770 (N_3770,N_3305,N_3142);
nand U3771 (N_3771,N_3133,N_3201);
or U3772 (N_3772,N_3037,N_3155);
xor U3773 (N_3773,N_3489,N_3409);
nor U3774 (N_3774,N_3305,N_3343);
nand U3775 (N_3775,N_3170,N_3276);
and U3776 (N_3776,N_3042,N_3050);
or U3777 (N_3777,N_3297,N_3188);
xor U3778 (N_3778,N_3240,N_3081);
nand U3779 (N_3779,N_3272,N_3251);
nand U3780 (N_3780,N_3421,N_3141);
and U3781 (N_3781,N_3482,N_3325);
and U3782 (N_3782,N_3310,N_3403);
nand U3783 (N_3783,N_3066,N_3442);
nor U3784 (N_3784,N_3368,N_3216);
nand U3785 (N_3785,N_3140,N_3495);
nor U3786 (N_3786,N_3218,N_3410);
or U3787 (N_3787,N_3239,N_3414);
and U3788 (N_3788,N_3391,N_3117);
and U3789 (N_3789,N_3213,N_3449);
and U3790 (N_3790,N_3002,N_3241);
nor U3791 (N_3791,N_3116,N_3099);
or U3792 (N_3792,N_3209,N_3452);
nand U3793 (N_3793,N_3008,N_3301);
xor U3794 (N_3794,N_3489,N_3321);
or U3795 (N_3795,N_3235,N_3344);
nand U3796 (N_3796,N_3109,N_3378);
xnor U3797 (N_3797,N_3184,N_3239);
nand U3798 (N_3798,N_3261,N_3470);
nand U3799 (N_3799,N_3043,N_3059);
nor U3800 (N_3800,N_3217,N_3216);
nor U3801 (N_3801,N_3002,N_3367);
nand U3802 (N_3802,N_3292,N_3438);
xor U3803 (N_3803,N_3198,N_3361);
and U3804 (N_3804,N_3027,N_3220);
or U3805 (N_3805,N_3056,N_3074);
nand U3806 (N_3806,N_3084,N_3437);
xnor U3807 (N_3807,N_3158,N_3307);
or U3808 (N_3808,N_3276,N_3349);
and U3809 (N_3809,N_3176,N_3283);
and U3810 (N_3810,N_3103,N_3155);
nand U3811 (N_3811,N_3075,N_3298);
nand U3812 (N_3812,N_3092,N_3435);
nand U3813 (N_3813,N_3130,N_3297);
nor U3814 (N_3814,N_3355,N_3294);
xor U3815 (N_3815,N_3050,N_3442);
or U3816 (N_3816,N_3460,N_3254);
or U3817 (N_3817,N_3135,N_3418);
nand U3818 (N_3818,N_3190,N_3054);
nand U3819 (N_3819,N_3290,N_3066);
nor U3820 (N_3820,N_3182,N_3125);
xor U3821 (N_3821,N_3298,N_3414);
nor U3822 (N_3822,N_3448,N_3330);
nand U3823 (N_3823,N_3164,N_3124);
and U3824 (N_3824,N_3360,N_3107);
nand U3825 (N_3825,N_3211,N_3307);
nand U3826 (N_3826,N_3340,N_3138);
or U3827 (N_3827,N_3162,N_3403);
nor U3828 (N_3828,N_3201,N_3357);
nor U3829 (N_3829,N_3318,N_3071);
or U3830 (N_3830,N_3119,N_3251);
and U3831 (N_3831,N_3253,N_3293);
or U3832 (N_3832,N_3437,N_3008);
nand U3833 (N_3833,N_3411,N_3446);
nand U3834 (N_3834,N_3291,N_3070);
and U3835 (N_3835,N_3089,N_3257);
or U3836 (N_3836,N_3054,N_3241);
or U3837 (N_3837,N_3281,N_3101);
nor U3838 (N_3838,N_3433,N_3403);
and U3839 (N_3839,N_3430,N_3465);
nor U3840 (N_3840,N_3477,N_3451);
xnor U3841 (N_3841,N_3386,N_3260);
nand U3842 (N_3842,N_3375,N_3421);
nor U3843 (N_3843,N_3363,N_3302);
and U3844 (N_3844,N_3204,N_3324);
nand U3845 (N_3845,N_3087,N_3335);
nand U3846 (N_3846,N_3071,N_3093);
or U3847 (N_3847,N_3379,N_3287);
xor U3848 (N_3848,N_3398,N_3358);
xor U3849 (N_3849,N_3045,N_3311);
nand U3850 (N_3850,N_3415,N_3290);
nor U3851 (N_3851,N_3300,N_3064);
nand U3852 (N_3852,N_3430,N_3050);
or U3853 (N_3853,N_3227,N_3054);
nand U3854 (N_3854,N_3441,N_3224);
xnor U3855 (N_3855,N_3059,N_3409);
or U3856 (N_3856,N_3450,N_3437);
and U3857 (N_3857,N_3235,N_3033);
xnor U3858 (N_3858,N_3173,N_3297);
nor U3859 (N_3859,N_3091,N_3438);
xor U3860 (N_3860,N_3139,N_3207);
xnor U3861 (N_3861,N_3151,N_3409);
nand U3862 (N_3862,N_3332,N_3269);
nand U3863 (N_3863,N_3007,N_3433);
nand U3864 (N_3864,N_3260,N_3415);
nand U3865 (N_3865,N_3086,N_3232);
and U3866 (N_3866,N_3499,N_3252);
nand U3867 (N_3867,N_3316,N_3255);
and U3868 (N_3868,N_3114,N_3054);
nor U3869 (N_3869,N_3396,N_3443);
or U3870 (N_3870,N_3362,N_3292);
and U3871 (N_3871,N_3070,N_3006);
nor U3872 (N_3872,N_3350,N_3359);
nand U3873 (N_3873,N_3348,N_3251);
or U3874 (N_3874,N_3271,N_3289);
nand U3875 (N_3875,N_3088,N_3026);
and U3876 (N_3876,N_3468,N_3204);
or U3877 (N_3877,N_3233,N_3477);
nor U3878 (N_3878,N_3083,N_3079);
nand U3879 (N_3879,N_3404,N_3032);
and U3880 (N_3880,N_3286,N_3219);
or U3881 (N_3881,N_3189,N_3431);
nand U3882 (N_3882,N_3298,N_3456);
or U3883 (N_3883,N_3337,N_3114);
nand U3884 (N_3884,N_3473,N_3155);
xnor U3885 (N_3885,N_3342,N_3400);
nor U3886 (N_3886,N_3092,N_3059);
nor U3887 (N_3887,N_3047,N_3322);
xnor U3888 (N_3888,N_3038,N_3334);
nand U3889 (N_3889,N_3479,N_3422);
nor U3890 (N_3890,N_3356,N_3338);
nor U3891 (N_3891,N_3090,N_3270);
or U3892 (N_3892,N_3270,N_3438);
and U3893 (N_3893,N_3040,N_3015);
nand U3894 (N_3894,N_3135,N_3481);
and U3895 (N_3895,N_3247,N_3073);
nor U3896 (N_3896,N_3259,N_3444);
and U3897 (N_3897,N_3446,N_3286);
and U3898 (N_3898,N_3138,N_3268);
nand U3899 (N_3899,N_3444,N_3379);
nor U3900 (N_3900,N_3368,N_3127);
nor U3901 (N_3901,N_3440,N_3472);
nand U3902 (N_3902,N_3293,N_3398);
xnor U3903 (N_3903,N_3455,N_3368);
and U3904 (N_3904,N_3264,N_3034);
nand U3905 (N_3905,N_3140,N_3257);
and U3906 (N_3906,N_3205,N_3399);
or U3907 (N_3907,N_3313,N_3426);
and U3908 (N_3908,N_3174,N_3449);
or U3909 (N_3909,N_3146,N_3387);
or U3910 (N_3910,N_3475,N_3015);
and U3911 (N_3911,N_3419,N_3206);
xor U3912 (N_3912,N_3390,N_3033);
nor U3913 (N_3913,N_3064,N_3423);
or U3914 (N_3914,N_3324,N_3036);
nand U3915 (N_3915,N_3029,N_3437);
xor U3916 (N_3916,N_3488,N_3175);
or U3917 (N_3917,N_3294,N_3455);
nand U3918 (N_3918,N_3073,N_3221);
nor U3919 (N_3919,N_3356,N_3122);
nor U3920 (N_3920,N_3087,N_3387);
xor U3921 (N_3921,N_3219,N_3499);
nor U3922 (N_3922,N_3122,N_3310);
nor U3923 (N_3923,N_3366,N_3361);
and U3924 (N_3924,N_3104,N_3409);
and U3925 (N_3925,N_3390,N_3465);
xnor U3926 (N_3926,N_3059,N_3286);
and U3927 (N_3927,N_3025,N_3113);
nand U3928 (N_3928,N_3351,N_3151);
nand U3929 (N_3929,N_3352,N_3385);
nand U3930 (N_3930,N_3314,N_3340);
nand U3931 (N_3931,N_3139,N_3231);
xor U3932 (N_3932,N_3484,N_3248);
and U3933 (N_3933,N_3311,N_3272);
nor U3934 (N_3934,N_3183,N_3091);
xor U3935 (N_3935,N_3097,N_3369);
xor U3936 (N_3936,N_3162,N_3048);
nand U3937 (N_3937,N_3310,N_3356);
xnor U3938 (N_3938,N_3419,N_3022);
xnor U3939 (N_3939,N_3116,N_3307);
nand U3940 (N_3940,N_3101,N_3188);
xnor U3941 (N_3941,N_3043,N_3396);
xor U3942 (N_3942,N_3258,N_3081);
nand U3943 (N_3943,N_3495,N_3329);
nor U3944 (N_3944,N_3017,N_3130);
and U3945 (N_3945,N_3204,N_3228);
nand U3946 (N_3946,N_3051,N_3289);
or U3947 (N_3947,N_3314,N_3305);
and U3948 (N_3948,N_3462,N_3195);
and U3949 (N_3949,N_3117,N_3172);
or U3950 (N_3950,N_3355,N_3459);
xnor U3951 (N_3951,N_3287,N_3285);
nand U3952 (N_3952,N_3114,N_3011);
nand U3953 (N_3953,N_3138,N_3282);
nand U3954 (N_3954,N_3307,N_3221);
or U3955 (N_3955,N_3482,N_3155);
xor U3956 (N_3956,N_3293,N_3280);
nand U3957 (N_3957,N_3146,N_3490);
nand U3958 (N_3958,N_3265,N_3182);
xnor U3959 (N_3959,N_3334,N_3187);
xnor U3960 (N_3960,N_3162,N_3164);
or U3961 (N_3961,N_3087,N_3093);
xor U3962 (N_3962,N_3306,N_3452);
and U3963 (N_3963,N_3418,N_3205);
and U3964 (N_3964,N_3245,N_3414);
nand U3965 (N_3965,N_3488,N_3407);
and U3966 (N_3966,N_3052,N_3275);
and U3967 (N_3967,N_3194,N_3477);
nand U3968 (N_3968,N_3321,N_3499);
or U3969 (N_3969,N_3045,N_3124);
or U3970 (N_3970,N_3444,N_3220);
nand U3971 (N_3971,N_3180,N_3371);
nand U3972 (N_3972,N_3247,N_3268);
nor U3973 (N_3973,N_3420,N_3081);
and U3974 (N_3974,N_3323,N_3483);
and U3975 (N_3975,N_3479,N_3215);
or U3976 (N_3976,N_3063,N_3429);
and U3977 (N_3977,N_3286,N_3382);
nand U3978 (N_3978,N_3303,N_3496);
xor U3979 (N_3979,N_3141,N_3089);
nand U3980 (N_3980,N_3094,N_3122);
xnor U3981 (N_3981,N_3094,N_3019);
or U3982 (N_3982,N_3355,N_3198);
and U3983 (N_3983,N_3141,N_3058);
nand U3984 (N_3984,N_3173,N_3121);
and U3985 (N_3985,N_3208,N_3444);
or U3986 (N_3986,N_3173,N_3201);
and U3987 (N_3987,N_3420,N_3116);
and U3988 (N_3988,N_3158,N_3388);
nor U3989 (N_3989,N_3133,N_3194);
and U3990 (N_3990,N_3147,N_3152);
xor U3991 (N_3991,N_3200,N_3431);
nor U3992 (N_3992,N_3214,N_3410);
nand U3993 (N_3993,N_3486,N_3098);
nand U3994 (N_3994,N_3360,N_3009);
and U3995 (N_3995,N_3394,N_3436);
nand U3996 (N_3996,N_3449,N_3438);
or U3997 (N_3997,N_3226,N_3032);
and U3998 (N_3998,N_3206,N_3455);
or U3999 (N_3999,N_3262,N_3420);
nand U4000 (N_4000,N_3702,N_3868);
nor U4001 (N_4001,N_3812,N_3568);
xor U4002 (N_4002,N_3594,N_3737);
xor U4003 (N_4003,N_3605,N_3513);
and U4004 (N_4004,N_3623,N_3682);
xor U4005 (N_4005,N_3571,N_3960);
nor U4006 (N_4006,N_3723,N_3769);
or U4007 (N_4007,N_3813,N_3668);
xor U4008 (N_4008,N_3907,N_3549);
nor U4009 (N_4009,N_3649,N_3806);
and U4010 (N_4010,N_3712,N_3562);
nor U4011 (N_4011,N_3899,N_3932);
nand U4012 (N_4012,N_3820,N_3785);
and U4013 (N_4013,N_3540,N_3997);
nand U4014 (N_4014,N_3503,N_3546);
xnor U4015 (N_4015,N_3697,N_3939);
nand U4016 (N_4016,N_3828,N_3535);
or U4017 (N_4017,N_3687,N_3940);
or U4018 (N_4018,N_3539,N_3916);
nor U4019 (N_4019,N_3840,N_3937);
xor U4020 (N_4020,N_3779,N_3629);
nor U4021 (N_4021,N_3545,N_3793);
xnor U4022 (N_4022,N_3816,N_3578);
and U4023 (N_4023,N_3517,N_3800);
or U4024 (N_4024,N_3598,N_3876);
and U4025 (N_4025,N_3710,N_3867);
and U4026 (N_4026,N_3835,N_3957);
and U4027 (N_4027,N_3659,N_3639);
and U4028 (N_4028,N_3902,N_3525);
nand U4029 (N_4029,N_3759,N_3972);
or U4030 (N_4030,N_3642,N_3859);
xnor U4031 (N_4031,N_3755,N_3652);
xnor U4032 (N_4032,N_3852,N_3830);
nand U4033 (N_4033,N_3938,N_3711);
xnor U4034 (N_4034,N_3945,N_3760);
nor U4035 (N_4035,N_3610,N_3921);
xor U4036 (N_4036,N_3834,N_3538);
nor U4037 (N_4037,N_3703,N_3574);
xor U4038 (N_4038,N_3903,N_3974);
xnor U4039 (N_4039,N_3688,N_3836);
nor U4040 (N_4040,N_3604,N_3678);
and U4041 (N_4041,N_3927,N_3608);
nor U4042 (N_4042,N_3507,N_3519);
nand U4043 (N_4043,N_3615,N_3500);
nor U4044 (N_4044,N_3991,N_3817);
nor U4045 (N_4045,N_3625,N_3695);
and U4046 (N_4046,N_3635,N_3602);
or U4047 (N_4047,N_3738,N_3827);
xor U4048 (N_4048,N_3632,N_3954);
xor U4049 (N_4049,N_3797,N_3626);
or U4050 (N_4050,N_3566,N_3883);
and U4051 (N_4051,N_3951,N_3727);
and U4052 (N_4052,N_3681,N_3796);
and U4053 (N_4053,N_3736,N_3998);
nand U4054 (N_4054,N_3512,N_3650);
and U4055 (N_4055,N_3700,N_3518);
nor U4056 (N_4056,N_3822,N_3734);
or U4057 (N_4057,N_3897,N_3742);
or U4058 (N_4058,N_3805,N_3728);
and U4059 (N_4059,N_3775,N_3637);
or U4060 (N_4060,N_3772,N_3558);
or U4061 (N_4061,N_3744,N_3587);
and U4062 (N_4062,N_3743,N_3524);
nand U4063 (N_4063,N_3798,N_3537);
nand U4064 (N_4064,N_3630,N_3829);
nor U4065 (N_4065,N_3508,N_3963);
nor U4066 (N_4066,N_3694,N_3962);
and U4067 (N_4067,N_3837,N_3582);
nand U4068 (N_4068,N_3502,N_3993);
xor U4069 (N_4069,N_3715,N_3882);
nand U4070 (N_4070,N_3941,N_3799);
nor U4071 (N_4071,N_3595,N_3655);
nand U4072 (N_4072,N_3689,N_3654);
or U4073 (N_4073,N_3893,N_3748);
nor U4074 (N_4074,N_3590,N_3819);
nor U4075 (N_4075,N_3633,N_3887);
or U4076 (N_4076,N_3912,N_3789);
xor U4077 (N_4077,N_3795,N_3923);
xor U4078 (N_4078,N_3643,N_3889);
or U4079 (N_4079,N_3976,N_3908);
xor U4080 (N_4080,N_3956,N_3871);
xnor U4081 (N_4081,N_3802,N_3950);
xnor U4082 (N_4082,N_3968,N_3705);
xor U4083 (N_4083,N_3851,N_3999);
or U4084 (N_4084,N_3870,N_3543);
nand U4085 (N_4085,N_3922,N_3911);
xor U4086 (N_4086,N_3888,N_3520);
or U4087 (N_4087,N_3551,N_3706);
xnor U4088 (N_4088,N_3641,N_3725);
nand U4089 (N_4089,N_3638,N_3801);
or U4090 (N_4090,N_3761,N_3909);
nand U4091 (N_4091,N_3698,N_3529);
and U4092 (N_4092,N_3560,N_3844);
or U4093 (N_4093,N_3614,N_3881);
and U4094 (N_4094,N_3784,N_3661);
or U4095 (N_4095,N_3684,N_3603);
or U4096 (N_4096,N_3606,N_3949);
and U4097 (N_4097,N_3901,N_3692);
or U4098 (N_4098,N_3669,N_3860);
nor U4099 (N_4099,N_3847,N_3570);
xor U4100 (N_4100,N_3588,N_3778);
or U4101 (N_4101,N_3541,N_3573);
or U4102 (N_4102,N_3644,N_3515);
nand U4103 (N_4103,N_3704,N_3803);
or U4104 (N_4104,N_3589,N_3777);
nor U4105 (N_4105,N_3690,N_3708);
nand U4106 (N_4106,N_3825,N_3961);
and U4107 (N_4107,N_3620,N_3826);
or U4108 (N_4108,N_3933,N_3823);
nor U4109 (N_4109,N_3624,N_3677);
or U4110 (N_4110,N_3717,N_3965);
or U4111 (N_4111,N_3707,N_3721);
or U4112 (N_4112,N_3579,N_3634);
and U4113 (N_4113,N_3861,N_3985);
nor U4114 (N_4114,N_3699,N_3658);
and U4115 (N_4115,N_3930,N_3880);
xor U4116 (N_4116,N_3955,N_3900);
xnor U4117 (N_4117,N_3771,N_3757);
or U4118 (N_4118,N_3832,N_3647);
and U4119 (N_4119,N_3651,N_3670);
xor U4120 (N_4120,N_3514,N_3885);
nand U4121 (N_4121,N_3730,N_3758);
nand U4122 (N_4122,N_3875,N_3718);
or U4123 (N_4123,N_3714,N_3733);
nor U4124 (N_4124,N_3596,N_3746);
and U4125 (N_4125,N_3653,N_3747);
nor U4126 (N_4126,N_3722,N_3586);
or U4127 (N_4127,N_3934,N_3989);
xnor U4128 (N_4128,N_3848,N_3865);
and U4129 (N_4129,N_3931,N_3522);
or U4130 (N_4130,N_3762,N_3745);
nor U4131 (N_4131,N_3988,N_3774);
nor U4132 (N_4132,N_3843,N_3996);
nand U4133 (N_4133,N_3983,N_3874);
or U4134 (N_4134,N_3905,N_3857);
nand U4135 (N_4135,N_3534,N_3929);
or U4136 (N_4136,N_3731,N_3966);
nand U4137 (N_4137,N_3782,N_3918);
nand U4138 (N_4138,N_3726,N_3942);
xnor U4139 (N_4139,N_3863,N_3947);
xor U4140 (N_4140,N_3808,N_3601);
or U4141 (N_4141,N_3729,N_3713);
xor U4142 (N_4142,N_3913,N_3628);
xor U4143 (N_4143,N_3580,N_3952);
or U4144 (N_4144,N_3794,N_3925);
nor U4145 (N_4145,N_3631,N_3686);
xor U4146 (N_4146,N_3809,N_3679);
nand U4147 (N_4147,N_3609,N_3948);
and U4148 (N_4148,N_3563,N_3831);
nor U4149 (N_4149,N_3676,N_3862);
nor U4150 (N_4150,N_3553,N_3982);
nand U4151 (N_4151,N_3572,N_3756);
nor U4152 (N_4152,N_3550,N_3716);
and U4153 (N_4153,N_3971,N_3839);
nor U4154 (N_4154,N_3510,N_3926);
nand U4155 (N_4155,N_3592,N_3667);
xor U4156 (N_4156,N_3719,N_3646);
nor U4157 (N_4157,N_3878,N_3662);
nand U4158 (N_4158,N_3898,N_3856);
xor U4159 (N_4159,N_3788,N_3842);
nand U4160 (N_4160,N_3523,N_3763);
and U4161 (N_4161,N_3564,N_3919);
and U4162 (N_4162,N_3599,N_3556);
and U4163 (N_4163,N_3527,N_3986);
and U4164 (N_4164,N_3724,N_3866);
or U4165 (N_4165,N_3928,N_3768);
or U4166 (N_4166,N_3750,N_3845);
xnor U4167 (N_4167,N_3969,N_3663);
and U4168 (N_4168,N_3627,N_3924);
nor U4169 (N_4169,N_3531,N_3685);
nand U4170 (N_4170,N_3765,N_3906);
nand U4171 (N_4171,N_3896,N_3561);
and U4172 (N_4172,N_3533,N_3884);
xnor U4173 (N_4173,N_3980,N_3886);
xor U4174 (N_4174,N_3548,N_3532);
nand U4175 (N_4175,N_3766,N_3877);
nor U4176 (N_4176,N_3753,N_3672);
nand U4177 (N_4177,N_3872,N_3767);
xnor U4178 (N_4178,N_3611,N_3990);
xor U4179 (N_4179,N_3987,N_3559);
nor U4180 (N_4180,N_3879,N_3910);
nand U4181 (N_4181,N_3555,N_3814);
nand U4182 (N_4182,N_3776,N_3890);
nand U4183 (N_4183,N_3790,N_3853);
or U4184 (N_4184,N_3552,N_3645);
xor U4185 (N_4185,N_3554,N_3739);
xor U4186 (N_4186,N_3977,N_3864);
nor U4187 (N_4187,N_3693,N_3577);
and U4188 (N_4188,N_3978,N_3984);
nor U4189 (N_4189,N_3607,N_3591);
or U4190 (N_4190,N_3838,N_3849);
or U4191 (N_4191,N_3873,N_3617);
nor U4192 (N_4192,N_3660,N_3516);
nor U4193 (N_4193,N_3869,N_3576);
xor U4194 (N_4194,N_3944,N_3557);
and U4195 (N_4195,N_3585,N_3581);
nand U4196 (N_4196,N_3674,N_3975);
nor U4197 (N_4197,N_3501,N_3970);
nor U4198 (N_4198,N_3696,N_3741);
nand U4199 (N_4199,N_3992,N_3846);
nor U4200 (N_4200,N_3973,N_3764);
and U4201 (N_4201,N_3749,N_3858);
and U4202 (N_4202,N_3953,N_3709);
nand U4203 (N_4203,N_3701,N_3612);
and U4204 (N_4204,N_3786,N_3967);
nand U4205 (N_4205,N_3521,N_3673);
nor U4206 (N_4206,N_3657,N_3979);
nand U4207 (N_4207,N_3509,N_3664);
nor U4208 (N_4208,N_3671,N_3680);
nor U4209 (N_4209,N_3773,N_3787);
xnor U4210 (N_4210,N_3584,N_3735);
nor U4211 (N_4211,N_3754,N_3824);
xnor U4212 (N_4212,N_3740,N_3506);
nand U4213 (N_4213,N_3981,N_3565);
nor U4214 (N_4214,N_3994,N_3995);
and U4215 (N_4215,N_3621,N_3544);
nand U4216 (N_4216,N_3855,N_3936);
or U4217 (N_4217,N_3619,N_3807);
or U4218 (N_4218,N_3943,N_3528);
nand U4219 (N_4219,N_3600,N_3622);
or U4220 (N_4220,N_3616,N_3666);
or U4221 (N_4221,N_3583,N_3511);
and U4222 (N_4222,N_3648,N_3720);
xor U4223 (N_4223,N_3613,N_3542);
or U4224 (N_4224,N_3504,N_3547);
nand U4225 (N_4225,N_3752,N_3804);
nor U4226 (N_4226,N_3683,N_3618);
nor U4227 (N_4227,N_3791,N_3854);
or U4228 (N_4228,N_3959,N_3815);
nor U4229 (N_4229,N_3935,N_3640);
xnor U4230 (N_4230,N_3567,N_3904);
nor U4231 (N_4231,N_3895,N_3920);
and U4232 (N_4232,N_3811,N_3569);
nor U4233 (N_4233,N_3841,N_3792);
and U4234 (N_4234,N_3783,N_3850);
nor U4235 (N_4235,N_3691,N_3597);
nand U4236 (N_4236,N_3958,N_3770);
or U4237 (N_4237,N_3530,N_3526);
or U4238 (N_4238,N_3964,N_3915);
nand U4239 (N_4239,N_3917,N_3656);
nor U4240 (N_4240,N_3780,N_3894);
nand U4241 (N_4241,N_3821,N_3946);
nor U4242 (N_4242,N_3575,N_3833);
and U4243 (N_4243,N_3810,N_3914);
nor U4244 (N_4244,N_3891,N_3818);
or U4245 (N_4245,N_3675,N_3593);
or U4246 (N_4246,N_3665,N_3781);
nor U4247 (N_4247,N_3505,N_3536);
nand U4248 (N_4248,N_3636,N_3732);
nor U4249 (N_4249,N_3751,N_3892);
or U4250 (N_4250,N_3833,N_3944);
nor U4251 (N_4251,N_3585,N_3682);
nor U4252 (N_4252,N_3662,N_3673);
xnor U4253 (N_4253,N_3931,N_3820);
nand U4254 (N_4254,N_3754,N_3619);
nor U4255 (N_4255,N_3766,N_3519);
and U4256 (N_4256,N_3913,N_3598);
nor U4257 (N_4257,N_3867,N_3521);
nor U4258 (N_4258,N_3699,N_3594);
and U4259 (N_4259,N_3663,N_3920);
or U4260 (N_4260,N_3907,N_3994);
nand U4261 (N_4261,N_3502,N_3729);
nor U4262 (N_4262,N_3616,N_3692);
or U4263 (N_4263,N_3593,N_3989);
nor U4264 (N_4264,N_3900,N_3635);
nor U4265 (N_4265,N_3655,N_3905);
xor U4266 (N_4266,N_3651,N_3968);
or U4267 (N_4267,N_3762,N_3838);
or U4268 (N_4268,N_3807,N_3625);
nand U4269 (N_4269,N_3570,N_3920);
nor U4270 (N_4270,N_3669,N_3745);
nor U4271 (N_4271,N_3967,N_3548);
nand U4272 (N_4272,N_3752,N_3710);
nand U4273 (N_4273,N_3953,N_3931);
nand U4274 (N_4274,N_3838,N_3936);
or U4275 (N_4275,N_3515,N_3837);
and U4276 (N_4276,N_3932,N_3510);
xor U4277 (N_4277,N_3596,N_3925);
nand U4278 (N_4278,N_3638,N_3921);
xnor U4279 (N_4279,N_3634,N_3915);
or U4280 (N_4280,N_3840,N_3890);
and U4281 (N_4281,N_3899,N_3826);
and U4282 (N_4282,N_3953,N_3973);
nand U4283 (N_4283,N_3956,N_3570);
or U4284 (N_4284,N_3528,N_3905);
or U4285 (N_4285,N_3922,N_3588);
nand U4286 (N_4286,N_3868,N_3859);
and U4287 (N_4287,N_3688,N_3888);
nand U4288 (N_4288,N_3657,N_3989);
and U4289 (N_4289,N_3947,N_3814);
and U4290 (N_4290,N_3817,N_3613);
and U4291 (N_4291,N_3711,N_3901);
nand U4292 (N_4292,N_3813,N_3763);
and U4293 (N_4293,N_3673,N_3683);
nor U4294 (N_4294,N_3611,N_3732);
or U4295 (N_4295,N_3832,N_3511);
and U4296 (N_4296,N_3534,N_3965);
nand U4297 (N_4297,N_3733,N_3818);
nand U4298 (N_4298,N_3624,N_3928);
and U4299 (N_4299,N_3962,N_3626);
xnor U4300 (N_4300,N_3565,N_3573);
and U4301 (N_4301,N_3736,N_3663);
and U4302 (N_4302,N_3524,N_3905);
and U4303 (N_4303,N_3543,N_3714);
or U4304 (N_4304,N_3754,N_3978);
nor U4305 (N_4305,N_3507,N_3857);
nand U4306 (N_4306,N_3572,N_3863);
or U4307 (N_4307,N_3785,N_3766);
and U4308 (N_4308,N_3790,N_3711);
and U4309 (N_4309,N_3711,N_3854);
xor U4310 (N_4310,N_3813,N_3712);
and U4311 (N_4311,N_3985,N_3614);
xnor U4312 (N_4312,N_3527,N_3796);
nand U4313 (N_4313,N_3712,N_3955);
xor U4314 (N_4314,N_3923,N_3894);
nor U4315 (N_4315,N_3673,N_3913);
nand U4316 (N_4316,N_3776,N_3900);
nor U4317 (N_4317,N_3634,N_3941);
and U4318 (N_4318,N_3662,N_3604);
xnor U4319 (N_4319,N_3971,N_3820);
xor U4320 (N_4320,N_3789,N_3803);
and U4321 (N_4321,N_3544,N_3537);
xnor U4322 (N_4322,N_3996,N_3710);
and U4323 (N_4323,N_3519,N_3933);
or U4324 (N_4324,N_3596,N_3983);
xnor U4325 (N_4325,N_3897,N_3822);
xnor U4326 (N_4326,N_3642,N_3827);
xor U4327 (N_4327,N_3710,N_3985);
xor U4328 (N_4328,N_3866,N_3668);
and U4329 (N_4329,N_3933,N_3749);
and U4330 (N_4330,N_3766,N_3848);
or U4331 (N_4331,N_3797,N_3953);
or U4332 (N_4332,N_3986,N_3887);
and U4333 (N_4333,N_3828,N_3583);
nor U4334 (N_4334,N_3715,N_3805);
nor U4335 (N_4335,N_3508,N_3606);
nand U4336 (N_4336,N_3879,N_3633);
nand U4337 (N_4337,N_3615,N_3717);
xnor U4338 (N_4338,N_3844,N_3944);
nor U4339 (N_4339,N_3560,N_3524);
nor U4340 (N_4340,N_3973,N_3640);
nor U4341 (N_4341,N_3817,N_3795);
or U4342 (N_4342,N_3545,N_3726);
nor U4343 (N_4343,N_3961,N_3619);
or U4344 (N_4344,N_3661,N_3853);
and U4345 (N_4345,N_3607,N_3558);
or U4346 (N_4346,N_3859,N_3775);
or U4347 (N_4347,N_3853,N_3517);
and U4348 (N_4348,N_3874,N_3756);
or U4349 (N_4349,N_3774,N_3792);
nor U4350 (N_4350,N_3624,N_3971);
xor U4351 (N_4351,N_3829,N_3934);
and U4352 (N_4352,N_3676,N_3756);
xor U4353 (N_4353,N_3868,N_3897);
nand U4354 (N_4354,N_3668,N_3926);
or U4355 (N_4355,N_3916,N_3840);
xnor U4356 (N_4356,N_3766,N_3968);
or U4357 (N_4357,N_3507,N_3760);
nor U4358 (N_4358,N_3596,N_3624);
xnor U4359 (N_4359,N_3701,N_3806);
nand U4360 (N_4360,N_3605,N_3522);
nor U4361 (N_4361,N_3582,N_3705);
nand U4362 (N_4362,N_3640,N_3932);
and U4363 (N_4363,N_3971,N_3526);
or U4364 (N_4364,N_3714,N_3720);
nor U4365 (N_4365,N_3569,N_3605);
nor U4366 (N_4366,N_3891,N_3519);
nand U4367 (N_4367,N_3878,N_3552);
nor U4368 (N_4368,N_3845,N_3819);
xnor U4369 (N_4369,N_3869,N_3662);
xnor U4370 (N_4370,N_3571,N_3530);
and U4371 (N_4371,N_3505,N_3600);
and U4372 (N_4372,N_3834,N_3893);
nand U4373 (N_4373,N_3796,N_3579);
nor U4374 (N_4374,N_3713,N_3802);
nand U4375 (N_4375,N_3584,N_3884);
and U4376 (N_4376,N_3974,N_3739);
and U4377 (N_4377,N_3899,N_3959);
nand U4378 (N_4378,N_3793,N_3526);
xor U4379 (N_4379,N_3568,N_3631);
and U4380 (N_4380,N_3819,N_3884);
and U4381 (N_4381,N_3771,N_3754);
xor U4382 (N_4382,N_3944,N_3912);
nor U4383 (N_4383,N_3627,N_3948);
nand U4384 (N_4384,N_3928,N_3970);
nor U4385 (N_4385,N_3537,N_3715);
or U4386 (N_4386,N_3574,N_3517);
nor U4387 (N_4387,N_3590,N_3993);
nand U4388 (N_4388,N_3643,N_3835);
xor U4389 (N_4389,N_3852,N_3556);
and U4390 (N_4390,N_3712,N_3819);
xor U4391 (N_4391,N_3568,N_3673);
nor U4392 (N_4392,N_3865,N_3648);
nor U4393 (N_4393,N_3646,N_3534);
or U4394 (N_4394,N_3705,N_3696);
nand U4395 (N_4395,N_3921,N_3654);
nand U4396 (N_4396,N_3731,N_3669);
and U4397 (N_4397,N_3668,N_3899);
xnor U4398 (N_4398,N_3760,N_3673);
or U4399 (N_4399,N_3951,N_3939);
nor U4400 (N_4400,N_3705,N_3813);
xor U4401 (N_4401,N_3652,N_3639);
nor U4402 (N_4402,N_3761,N_3755);
and U4403 (N_4403,N_3635,N_3968);
or U4404 (N_4404,N_3838,N_3839);
nor U4405 (N_4405,N_3949,N_3996);
or U4406 (N_4406,N_3584,N_3889);
xnor U4407 (N_4407,N_3884,N_3521);
nand U4408 (N_4408,N_3960,N_3621);
xnor U4409 (N_4409,N_3750,N_3869);
nand U4410 (N_4410,N_3559,N_3772);
nand U4411 (N_4411,N_3950,N_3832);
nor U4412 (N_4412,N_3548,N_3554);
xor U4413 (N_4413,N_3773,N_3811);
xnor U4414 (N_4414,N_3812,N_3943);
nand U4415 (N_4415,N_3733,N_3698);
and U4416 (N_4416,N_3888,N_3930);
and U4417 (N_4417,N_3709,N_3633);
or U4418 (N_4418,N_3649,N_3864);
nand U4419 (N_4419,N_3860,N_3967);
nand U4420 (N_4420,N_3988,N_3859);
nand U4421 (N_4421,N_3876,N_3663);
and U4422 (N_4422,N_3876,N_3909);
and U4423 (N_4423,N_3833,N_3977);
nand U4424 (N_4424,N_3574,N_3794);
xor U4425 (N_4425,N_3658,N_3742);
nand U4426 (N_4426,N_3959,N_3945);
nor U4427 (N_4427,N_3947,N_3605);
nand U4428 (N_4428,N_3632,N_3831);
xnor U4429 (N_4429,N_3526,N_3966);
or U4430 (N_4430,N_3612,N_3850);
nand U4431 (N_4431,N_3686,N_3659);
xor U4432 (N_4432,N_3814,N_3587);
or U4433 (N_4433,N_3602,N_3877);
xor U4434 (N_4434,N_3972,N_3547);
or U4435 (N_4435,N_3627,N_3570);
nand U4436 (N_4436,N_3701,N_3728);
xor U4437 (N_4437,N_3848,N_3866);
xnor U4438 (N_4438,N_3927,N_3508);
nor U4439 (N_4439,N_3780,N_3862);
xnor U4440 (N_4440,N_3577,N_3930);
or U4441 (N_4441,N_3890,N_3595);
and U4442 (N_4442,N_3806,N_3630);
and U4443 (N_4443,N_3680,N_3830);
nand U4444 (N_4444,N_3898,N_3680);
nor U4445 (N_4445,N_3583,N_3643);
or U4446 (N_4446,N_3783,N_3935);
and U4447 (N_4447,N_3856,N_3529);
nand U4448 (N_4448,N_3627,N_3760);
xor U4449 (N_4449,N_3976,N_3522);
nand U4450 (N_4450,N_3649,N_3761);
or U4451 (N_4451,N_3967,N_3857);
and U4452 (N_4452,N_3758,N_3910);
nor U4453 (N_4453,N_3956,N_3747);
xnor U4454 (N_4454,N_3943,N_3794);
xnor U4455 (N_4455,N_3752,N_3797);
nor U4456 (N_4456,N_3523,N_3829);
xor U4457 (N_4457,N_3858,N_3682);
nand U4458 (N_4458,N_3549,N_3791);
xnor U4459 (N_4459,N_3647,N_3803);
nor U4460 (N_4460,N_3884,N_3698);
xor U4461 (N_4461,N_3936,N_3799);
nor U4462 (N_4462,N_3754,N_3751);
nor U4463 (N_4463,N_3741,N_3765);
xnor U4464 (N_4464,N_3575,N_3876);
xor U4465 (N_4465,N_3776,N_3833);
and U4466 (N_4466,N_3625,N_3973);
or U4467 (N_4467,N_3811,N_3517);
and U4468 (N_4468,N_3932,N_3524);
nand U4469 (N_4469,N_3955,N_3833);
and U4470 (N_4470,N_3767,N_3765);
nand U4471 (N_4471,N_3779,N_3933);
nor U4472 (N_4472,N_3963,N_3724);
and U4473 (N_4473,N_3715,N_3923);
nor U4474 (N_4474,N_3792,N_3642);
and U4475 (N_4475,N_3994,N_3951);
or U4476 (N_4476,N_3776,N_3881);
xnor U4477 (N_4477,N_3894,N_3618);
xor U4478 (N_4478,N_3958,N_3721);
xor U4479 (N_4479,N_3638,N_3568);
or U4480 (N_4480,N_3769,N_3526);
or U4481 (N_4481,N_3932,N_3949);
nand U4482 (N_4482,N_3820,N_3658);
or U4483 (N_4483,N_3602,N_3837);
xnor U4484 (N_4484,N_3570,N_3709);
or U4485 (N_4485,N_3730,N_3681);
and U4486 (N_4486,N_3715,N_3953);
nor U4487 (N_4487,N_3637,N_3798);
and U4488 (N_4488,N_3637,N_3655);
nor U4489 (N_4489,N_3607,N_3562);
or U4490 (N_4490,N_3846,N_3918);
xor U4491 (N_4491,N_3754,N_3852);
or U4492 (N_4492,N_3898,N_3679);
or U4493 (N_4493,N_3570,N_3631);
xor U4494 (N_4494,N_3945,N_3667);
nand U4495 (N_4495,N_3606,N_3629);
xor U4496 (N_4496,N_3834,N_3781);
nand U4497 (N_4497,N_3531,N_3829);
xor U4498 (N_4498,N_3799,N_3876);
and U4499 (N_4499,N_3885,N_3665);
nor U4500 (N_4500,N_4031,N_4224);
or U4501 (N_4501,N_4192,N_4148);
xnor U4502 (N_4502,N_4338,N_4344);
nor U4503 (N_4503,N_4069,N_4411);
or U4504 (N_4504,N_4391,N_4313);
xor U4505 (N_4505,N_4329,N_4264);
and U4506 (N_4506,N_4387,N_4015);
and U4507 (N_4507,N_4191,N_4169);
xnor U4508 (N_4508,N_4484,N_4258);
and U4509 (N_4509,N_4158,N_4410);
nor U4510 (N_4510,N_4199,N_4257);
nand U4511 (N_4511,N_4195,N_4016);
nand U4512 (N_4512,N_4077,N_4030);
and U4513 (N_4513,N_4168,N_4172);
xnor U4514 (N_4514,N_4390,N_4049);
and U4515 (N_4515,N_4092,N_4143);
nor U4516 (N_4516,N_4185,N_4413);
xnor U4517 (N_4517,N_4342,N_4333);
nand U4518 (N_4518,N_4446,N_4210);
nand U4519 (N_4519,N_4383,N_4164);
nand U4520 (N_4520,N_4109,N_4220);
and U4521 (N_4521,N_4020,N_4240);
nand U4522 (N_4522,N_4305,N_4459);
and U4523 (N_4523,N_4331,N_4415);
nand U4524 (N_4524,N_4443,N_4126);
nand U4525 (N_4525,N_4428,N_4440);
or U4526 (N_4526,N_4438,N_4426);
or U4527 (N_4527,N_4217,N_4091);
or U4528 (N_4528,N_4237,N_4263);
or U4529 (N_4529,N_4214,N_4256);
xor U4530 (N_4530,N_4182,N_4178);
and U4531 (N_4531,N_4088,N_4419);
and U4532 (N_4532,N_4017,N_4207);
and U4533 (N_4533,N_4054,N_4475);
xnor U4534 (N_4534,N_4011,N_4341);
and U4535 (N_4535,N_4485,N_4078);
nor U4536 (N_4536,N_4412,N_4119);
xor U4537 (N_4537,N_4299,N_4442);
xnor U4538 (N_4538,N_4370,N_4420);
xnor U4539 (N_4539,N_4469,N_4032);
and U4540 (N_4540,N_4395,N_4055);
and U4541 (N_4541,N_4368,N_4425);
xor U4542 (N_4542,N_4361,N_4375);
or U4543 (N_4543,N_4334,N_4246);
nand U4544 (N_4544,N_4067,N_4066);
and U4545 (N_4545,N_4297,N_4254);
nor U4546 (N_4546,N_4277,N_4394);
or U4547 (N_4547,N_4141,N_4293);
nor U4548 (N_4548,N_4371,N_4177);
or U4549 (N_4549,N_4006,N_4311);
or U4550 (N_4550,N_4111,N_4400);
or U4551 (N_4551,N_4019,N_4068);
xor U4552 (N_4552,N_4346,N_4212);
and U4553 (N_4553,N_4047,N_4275);
nor U4554 (N_4554,N_4445,N_4118);
or U4555 (N_4555,N_4093,N_4325);
or U4556 (N_4556,N_4022,N_4320);
and U4557 (N_4557,N_4384,N_4145);
nand U4558 (N_4558,N_4267,N_4405);
and U4559 (N_4559,N_4348,N_4244);
nand U4560 (N_4560,N_4125,N_4318);
xor U4561 (N_4561,N_4480,N_4095);
nand U4562 (N_4562,N_4472,N_4447);
xor U4563 (N_4563,N_4187,N_4037);
or U4564 (N_4564,N_4386,N_4324);
and U4565 (N_4565,N_4481,N_4228);
xnor U4566 (N_4566,N_4340,N_4154);
or U4567 (N_4567,N_4202,N_4276);
and U4568 (N_4568,N_4347,N_4427);
and U4569 (N_4569,N_4429,N_4079);
nor U4570 (N_4570,N_4269,N_4130);
xor U4571 (N_4571,N_4468,N_4087);
nor U4572 (N_4572,N_4121,N_4456);
xor U4573 (N_4573,N_4360,N_4153);
xor U4574 (N_4574,N_4490,N_4494);
nor U4575 (N_4575,N_4493,N_4038);
and U4576 (N_4576,N_4012,N_4014);
xor U4577 (N_4577,N_4096,N_4479);
or U4578 (N_4578,N_4174,N_4222);
and U4579 (N_4579,N_4262,N_4142);
nor U4580 (N_4580,N_4421,N_4180);
xor U4581 (N_4581,N_4251,N_4245);
nand U4582 (N_4582,N_4234,N_4165);
nand U4583 (N_4583,N_4110,N_4302);
or U4584 (N_4584,N_4482,N_4441);
nor U4585 (N_4585,N_4204,N_4287);
nor U4586 (N_4586,N_4013,N_4124);
and U4587 (N_4587,N_4487,N_4108);
nand U4588 (N_4588,N_4358,N_4356);
nor U4589 (N_4589,N_4451,N_4407);
nor U4590 (N_4590,N_4050,N_4290);
nand U4591 (N_4591,N_4406,N_4206);
nand U4592 (N_4592,N_4498,N_4089);
and U4593 (N_4593,N_4128,N_4063);
xor U4594 (N_4594,N_4422,N_4448);
or U4595 (N_4595,N_4488,N_4235);
xnor U4596 (N_4596,N_4053,N_4044);
and U4597 (N_4597,N_4464,N_4175);
and U4598 (N_4598,N_4266,N_4401);
or U4599 (N_4599,N_4437,N_4028);
nand U4600 (N_4600,N_4103,N_4355);
nor U4601 (N_4601,N_4363,N_4381);
nand U4602 (N_4602,N_4166,N_4179);
nor U4603 (N_4603,N_4416,N_4197);
and U4604 (N_4604,N_4167,N_4034);
nand U4605 (N_4605,N_4173,N_4357);
and U4606 (N_4606,N_4144,N_4260);
nand U4607 (N_4607,N_4403,N_4114);
nand U4608 (N_4608,N_4460,N_4393);
or U4609 (N_4609,N_4366,N_4193);
nand U4610 (N_4610,N_4156,N_4052);
or U4611 (N_4611,N_4376,N_4230);
nand U4612 (N_4612,N_4045,N_4289);
nand U4613 (N_4613,N_4473,N_4051);
nand U4614 (N_4614,N_4218,N_4307);
xnor U4615 (N_4615,N_4389,N_4261);
and U4616 (N_4616,N_4382,N_4072);
or U4617 (N_4617,N_4483,N_4379);
or U4618 (N_4618,N_4135,N_4236);
nand U4619 (N_4619,N_4303,N_4388);
nand U4620 (N_4620,N_4352,N_4221);
or U4621 (N_4621,N_4116,N_4057);
and U4622 (N_4622,N_4281,N_4436);
nand U4623 (N_4623,N_4080,N_4137);
xor U4624 (N_4624,N_4280,N_4326);
xor U4625 (N_4625,N_4385,N_4397);
xnor U4626 (N_4626,N_4198,N_4139);
nor U4627 (N_4627,N_4339,N_4084);
xnor U4628 (N_4628,N_4408,N_4252);
or U4629 (N_4629,N_4147,N_4184);
nand U4630 (N_4630,N_4150,N_4497);
nor U4631 (N_4631,N_4399,N_4211);
and U4632 (N_4632,N_4056,N_4157);
nor U4633 (N_4633,N_4486,N_4319);
nor U4634 (N_4634,N_4076,N_4033);
nor U4635 (N_4635,N_4181,N_4452);
xor U4636 (N_4636,N_4470,N_4009);
nand U4637 (N_4637,N_4186,N_4227);
nand U4638 (N_4638,N_4216,N_4102);
and U4639 (N_4639,N_4136,N_4278);
xor U4640 (N_4640,N_4369,N_4176);
xor U4641 (N_4641,N_4306,N_4499);
and U4642 (N_4642,N_4042,N_4300);
or U4643 (N_4643,N_4353,N_4304);
or U4644 (N_4644,N_4113,N_4496);
nor U4645 (N_4645,N_4398,N_4225);
nor U4646 (N_4646,N_4433,N_4284);
and U4647 (N_4647,N_4350,N_4373);
xnor U4648 (N_4648,N_4495,N_4010);
xnor U4649 (N_4649,N_4127,N_4285);
nor U4650 (N_4650,N_4248,N_4492);
and U4651 (N_4651,N_4163,N_4082);
nand U4652 (N_4652,N_4349,N_4120);
nor U4653 (N_4653,N_4336,N_4453);
and U4654 (N_4654,N_4461,N_4081);
and U4655 (N_4655,N_4435,N_4454);
xor U4656 (N_4656,N_4359,N_4070);
and U4657 (N_4657,N_4414,N_4086);
xnor U4658 (N_4658,N_4268,N_4471);
xor U4659 (N_4659,N_4238,N_4098);
or U4660 (N_4660,N_4465,N_4328);
xor U4661 (N_4661,N_4354,N_4007);
and U4662 (N_4662,N_4170,N_4040);
or U4663 (N_4663,N_4036,N_4226);
or U4664 (N_4664,N_4418,N_4335);
xor U4665 (N_4665,N_4314,N_4265);
nor U4666 (N_4666,N_4117,N_4374);
nand U4667 (N_4667,N_4308,N_4146);
or U4668 (N_4668,N_4477,N_4250);
and U4669 (N_4669,N_4378,N_4160);
nand U4670 (N_4670,N_4463,N_4190);
and U4671 (N_4671,N_4291,N_4083);
xor U4672 (N_4672,N_4122,N_4271);
nand U4673 (N_4673,N_4058,N_4457);
nand U4674 (N_4674,N_4123,N_4242);
nor U4675 (N_4675,N_4296,N_4330);
nand U4676 (N_4676,N_4364,N_4467);
or U4677 (N_4677,N_4085,N_4474);
and U4678 (N_4678,N_4159,N_4219);
or U4679 (N_4679,N_4273,N_4005);
nand U4680 (N_4680,N_4321,N_4097);
or U4681 (N_4681,N_4138,N_4112);
xnor U4682 (N_4682,N_4309,N_4115);
or U4683 (N_4683,N_4048,N_4104);
and U4684 (N_4684,N_4194,N_4233);
or U4685 (N_4685,N_4310,N_4362);
nor U4686 (N_4686,N_4337,N_4466);
nand U4687 (N_4687,N_4196,N_4298);
and U4688 (N_4688,N_4021,N_4423);
xnor U4689 (N_4689,N_4409,N_4476);
nand U4690 (N_4690,N_4001,N_4243);
nand U4691 (N_4691,N_4155,N_4343);
nand U4692 (N_4692,N_4312,N_4380);
nand U4693 (N_4693,N_4396,N_4215);
xor U4694 (N_4694,N_4027,N_4223);
nand U4695 (N_4695,N_4188,N_4023);
xnor U4696 (N_4696,N_4152,N_4171);
and U4697 (N_4697,N_4043,N_4024);
or U4698 (N_4698,N_4450,N_4231);
xor U4699 (N_4699,N_4327,N_4105);
nand U4700 (N_4700,N_4259,N_4404);
nand U4701 (N_4701,N_4149,N_4255);
nor U4702 (N_4702,N_4372,N_4444);
or U4703 (N_4703,N_4151,N_4377);
nor U4704 (N_4704,N_4288,N_4239);
nor U4705 (N_4705,N_4434,N_4029);
or U4706 (N_4706,N_4008,N_4041);
xor U4707 (N_4707,N_4491,N_4332);
nand U4708 (N_4708,N_4229,N_4424);
nand U4709 (N_4709,N_4365,N_4003);
nor U4710 (N_4710,N_4133,N_4201);
nand U4711 (N_4711,N_4489,N_4129);
nand U4712 (N_4712,N_4162,N_4200);
or U4713 (N_4713,N_4099,N_4455);
nand U4714 (N_4714,N_4417,N_4213);
nand U4715 (N_4715,N_4253,N_4430);
or U4716 (N_4716,N_4132,N_4059);
or U4717 (N_4717,N_4249,N_4134);
or U4718 (N_4718,N_4161,N_4062);
xnor U4719 (N_4719,N_4402,N_4322);
xor U4720 (N_4720,N_4351,N_4345);
xnor U4721 (N_4721,N_4283,N_4107);
xnor U4722 (N_4722,N_4094,N_4060);
nor U4723 (N_4723,N_4323,N_4478);
or U4724 (N_4724,N_4061,N_4203);
nand U4725 (N_4725,N_4458,N_4315);
nor U4726 (N_4726,N_4439,N_4292);
nor U4727 (N_4727,N_4462,N_4274);
nand U4728 (N_4728,N_4367,N_4449);
nor U4729 (N_4729,N_4241,N_4209);
xnor U4730 (N_4730,N_4025,N_4071);
or U4731 (N_4731,N_4431,N_4189);
xor U4732 (N_4732,N_4282,N_4073);
xor U4733 (N_4733,N_4272,N_4039);
xor U4734 (N_4734,N_4432,N_4035);
or U4735 (N_4735,N_4018,N_4208);
nor U4736 (N_4736,N_4301,N_4294);
and U4737 (N_4737,N_4002,N_4075);
xor U4738 (N_4738,N_4101,N_4286);
and U4739 (N_4739,N_4140,N_4247);
nand U4740 (N_4740,N_4106,N_4279);
or U4741 (N_4741,N_4090,N_4270);
xor U4742 (N_4742,N_4232,N_4316);
or U4743 (N_4743,N_4046,N_4026);
nor U4744 (N_4744,N_4074,N_4131);
or U4745 (N_4745,N_4392,N_4000);
xor U4746 (N_4746,N_4004,N_4100);
or U4747 (N_4747,N_4317,N_4205);
xnor U4748 (N_4748,N_4295,N_4065);
nand U4749 (N_4749,N_4064,N_4183);
or U4750 (N_4750,N_4451,N_4239);
nand U4751 (N_4751,N_4486,N_4204);
nand U4752 (N_4752,N_4302,N_4382);
and U4753 (N_4753,N_4262,N_4030);
or U4754 (N_4754,N_4235,N_4455);
or U4755 (N_4755,N_4152,N_4414);
and U4756 (N_4756,N_4048,N_4067);
nand U4757 (N_4757,N_4122,N_4406);
xor U4758 (N_4758,N_4435,N_4085);
xnor U4759 (N_4759,N_4135,N_4060);
nor U4760 (N_4760,N_4079,N_4040);
nand U4761 (N_4761,N_4129,N_4469);
nor U4762 (N_4762,N_4328,N_4314);
and U4763 (N_4763,N_4052,N_4194);
xor U4764 (N_4764,N_4095,N_4036);
or U4765 (N_4765,N_4461,N_4401);
or U4766 (N_4766,N_4203,N_4174);
nand U4767 (N_4767,N_4004,N_4045);
or U4768 (N_4768,N_4360,N_4434);
and U4769 (N_4769,N_4352,N_4158);
or U4770 (N_4770,N_4416,N_4079);
nor U4771 (N_4771,N_4488,N_4364);
or U4772 (N_4772,N_4250,N_4466);
xor U4773 (N_4773,N_4130,N_4354);
xnor U4774 (N_4774,N_4080,N_4349);
or U4775 (N_4775,N_4415,N_4368);
and U4776 (N_4776,N_4282,N_4489);
nor U4777 (N_4777,N_4137,N_4024);
nor U4778 (N_4778,N_4443,N_4107);
xnor U4779 (N_4779,N_4340,N_4217);
and U4780 (N_4780,N_4085,N_4473);
nand U4781 (N_4781,N_4029,N_4124);
and U4782 (N_4782,N_4027,N_4038);
xnor U4783 (N_4783,N_4249,N_4054);
nor U4784 (N_4784,N_4016,N_4441);
and U4785 (N_4785,N_4328,N_4079);
nand U4786 (N_4786,N_4275,N_4354);
or U4787 (N_4787,N_4365,N_4299);
nand U4788 (N_4788,N_4225,N_4165);
nand U4789 (N_4789,N_4250,N_4026);
and U4790 (N_4790,N_4369,N_4437);
nand U4791 (N_4791,N_4493,N_4154);
or U4792 (N_4792,N_4443,N_4300);
nand U4793 (N_4793,N_4422,N_4398);
nand U4794 (N_4794,N_4134,N_4397);
or U4795 (N_4795,N_4349,N_4046);
or U4796 (N_4796,N_4374,N_4368);
nand U4797 (N_4797,N_4045,N_4306);
nor U4798 (N_4798,N_4305,N_4077);
nor U4799 (N_4799,N_4151,N_4011);
nand U4800 (N_4800,N_4091,N_4448);
and U4801 (N_4801,N_4461,N_4271);
and U4802 (N_4802,N_4140,N_4281);
or U4803 (N_4803,N_4099,N_4393);
and U4804 (N_4804,N_4370,N_4279);
or U4805 (N_4805,N_4160,N_4180);
xor U4806 (N_4806,N_4341,N_4220);
and U4807 (N_4807,N_4470,N_4312);
xor U4808 (N_4808,N_4136,N_4004);
and U4809 (N_4809,N_4239,N_4009);
nand U4810 (N_4810,N_4451,N_4353);
or U4811 (N_4811,N_4481,N_4350);
nand U4812 (N_4812,N_4160,N_4426);
nor U4813 (N_4813,N_4170,N_4228);
nand U4814 (N_4814,N_4201,N_4441);
and U4815 (N_4815,N_4070,N_4466);
and U4816 (N_4816,N_4023,N_4398);
nor U4817 (N_4817,N_4148,N_4141);
or U4818 (N_4818,N_4252,N_4130);
nor U4819 (N_4819,N_4289,N_4430);
and U4820 (N_4820,N_4185,N_4304);
xnor U4821 (N_4821,N_4307,N_4357);
xnor U4822 (N_4822,N_4316,N_4263);
nand U4823 (N_4823,N_4364,N_4360);
nor U4824 (N_4824,N_4179,N_4252);
nand U4825 (N_4825,N_4497,N_4175);
xnor U4826 (N_4826,N_4055,N_4287);
xor U4827 (N_4827,N_4276,N_4181);
and U4828 (N_4828,N_4277,N_4284);
nor U4829 (N_4829,N_4316,N_4438);
nor U4830 (N_4830,N_4197,N_4232);
and U4831 (N_4831,N_4257,N_4080);
nor U4832 (N_4832,N_4357,N_4251);
xor U4833 (N_4833,N_4409,N_4314);
or U4834 (N_4834,N_4045,N_4450);
or U4835 (N_4835,N_4282,N_4387);
nand U4836 (N_4836,N_4055,N_4265);
nor U4837 (N_4837,N_4177,N_4155);
or U4838 (N_4838,N_4464,N_4333);
xor U4839 (N_4839,N_4047,N_4132);
nand U4840 (N_4840,N_4108,N_4029);
xor U4841 (N_4841,N_4337,N_4381);
nor U4842 (N_4842,N_4038,N_4100);
xor U4843 (N_4843,N_4322,N_4035);
and U4844 (N_4844,N_4071,N_4323);
nand U4845 (N_4845,N_4205,N_4237);
nor U4846 (N_4846,N_4343,N_4172);
and U4847 (N_4847,N_4473,N_4062);
and U4848 (N_4848,N_4015,N_4293);
nand U4849 (N_4849,N_4471,N_4371);
nor U4850 (N_4850,N_4187,N_4076);
and U4851 (N_4851,N_4423,N_4156);
nand U4852 (N_4852,N_4262,N_4029);
or U4853 (N_4853,N_4047,N_4100);
or U4854 (N_4854,N_4161,N_4397);
xor U4855 (N_4855,N_4070,N_4243);
or U4856 (N_4856,N_4235,N_4377);
nor U4857 (N_4857,N_4121,N_4192);
and U4858 (N_4858,N_4324,N_4471);
nand U4859 (N_4859,N_4000,N_4020);
nor U4860 (N_4860,N_4102,N_4012);
xnor U4861 (N_4861,N_4285,N_4428);
xnor U4862 (N_4862,N_4054,N_4285);
and U4863 (N_4863,N_4071,N_4299);
or U4864 (N_4864,N_4480,N_4137);
xnor U4865 (N_4865,N_4111,N_4047);
xor U4866 (N_4866,N_4479,N_4333);
xnor U4867 (N_4867,N_4304,N_4366);
xor U4868 (N_4868,N_4452,N_4402);
and U4869 (N_4869,N_4440,N_4345);
xor U4870 (N_4870,N_4032,N_4117);
or U4871 (N_4871,N_4119,N_4409);
and U4872 (N_4872,N_4109,N_4021);
nand U4873 (N_4873,N_4279,N_4467);
or U4874 (N_4874,N_4048,N_4154);
xor U4875 (N_4875,N_4366,N_4423);
nor U4876 (N_4876,N_4115,N_4441);
nor U4877 (N_4877,N_4324,N_4131);
nand U4878 (N_4878,N_4435,N_4138);
and U4879 (N_4879,N_4497,N_4294);
nor U4880 (N_4880,N_4019,N_4222);
or U4881 (N_4881,N_4303,N_4391);
nand U4882 (N_4882,N_4378,N_4037);
nand U4883 (N_4883,N_4019,N_4161);
nand U4884 (N_4884,N_4019,N_4169);
and U4885 (N_4885,N_4420,N_4221);
xor U4886 (N_4886,N_4094,N_4173);
or U4887 (N_4887,N_4283,N_4148);
and U4888 (N_4888,N_4431,N_4068);
nor U4889 (N_4889,N_4349,N_4126);
nand U4890 (N_4890,N_4417,N_4204);
or U4891 (N_4891,N_4406,N_4237);
nand U4892 (N_4892,N_4495,N_4038);
nand U4893 (N_4893,N_4461,N_4177);
xor U4894 (N_4894,N_4022,N_4381);
nor U4895 (N_4895,N_4442,N_4023);
and U4896 (N_4896,N_4439,N_4276);
and U4897 (N_4897,N_4331,N_4458);
or U4898 (N_4898,N_4182,N_4196);
nor U4899 (N_4899,N_4438,N_4379);
or U4900 (N_4900,N_4356,N_4219);
or U4901 (N_4901,N_4037,N_4252);
and U4902 (N_4902,N_4372,N_4413);
and U4903 (N_4903,N_4283,N_4455);
nor U4904 (N_4904,N_4004,N_4263);
xor U4905 (N_4905,N_4200,N_4425);
and U4906 (N_4906,N_4315,N_4379);
xor U4907 (N_4907,N_4388,N_4382);
nor U4908 (N_4908,N_4102,N_4406);
xor U4909 (N_4909,N_4434,N_4305);
and U4910 (N_4910,N_4404,N_4421);
nand U4911 (N_4911,N_4074,N_4178);
nor U4912 (N_4912,N_4245,N_4003);
and U4913 (N_4913,N_4089,N_4201);
nand U4914 (N_4914,N_4034,N_4063);
nand U4915 (N_4915,N_4417,N_4158);
and U4916 (N_4916,N_4085,N_4098);
and U4917 (N_4917,N_4455,N_4232);
nor U4918 (N_4918,N_4499,N_4070);
and U4919 (N_4919,N_4162,N_4134);
nor U4920 (N_4920,N_4241,N_4168);
xnor U4921 (N_4921,N_4423,N_4462);
or U4922 (N_4922,N_4468,N_4474);
or U4923 (N_4923,N_4154,N_4434);
or U4924 (N_4924,N_4094,N_4385);
or U4925 (N_4925,N_4386,N_4364);
nor U4926 (N_4926,N_4186,N_4487);
or U4927 (N_4927,N_4336,N_4192);
or U4928 (N_4928,N_4349,N_4437);
nand U4929 (N_4929,N_4478,N_4348);
nor U4930 (N_4930,N_4115,N_4493);
nand U4931 (N_4931,N_4074,N_4291);
nor U4932 (N_4932,N_4351,N_4479);
and U4933 (N_4933,N_4124,N_4490);
xnor U4934 (N_4934,N_4205,N_4004);
and U4935 (N_4935,N_4035,N_4431);
and U4936 (N_4936,N_4367,N_4162);
xor U4937 (N_4937,N_4117,N_4075);
nand U4938 (N_4938,N_4479,N_4129);
and U4939 (N_4939,N_4232,N_4007);
or U4940 (N_4940,N_4035,N_4159);
and U4941 (N_4941,N_4459,N_4209);
or U4942 (N_4942,N_4439,N_4121);
and U4943 (N_4943,N_4492,N_4442);
nor U4944 (N_4944,N_4453,N_4330);
and U4945 (N_4945,N_4006,N_4226);
or U4946 (N_4946,N_4432,N_4493);
and U4947 (N_4947,N_4186,N_4076);
xnor U4948 (N_4948,N_4340,N_4126);
xnor U4949 (N_4949,N_4361,N_4421);
nor U4950 (N_4950,N_4102,N_4015);
nor U4951 (N_4951,N_4399,N_4108);
nor U4952 (N_4952,N_4486,N_4209);
nor U4953 (N_4953,N_4332,N_4468);
nand U4954 (N_4954,N_4199,N_4093);
or U4955 (N_4955,N_4211,N_4418);
nor U4956 (N_4956,N_4212,N_4366);
nand U4957 (N_4957,N_4261,N_4450);
nand U4958 (N_4958,N_4323,N_4435);
nor U4959 (N_4959,N_4400,N_4249);
xor U4960 (N_4960,N_4475,N_4471);
and U4961 (N_4961,N_4289,N_4039);
nand U4962 (N_4962,N_4387,N_4026);
nand U4963 (N_4963,N_4242,N_4285);
nand U4964 (N_4964,N_4155,N_4036);
nand U4965 (N_4965,N_4400,N_4402);
or U4966 (N_4966,N_4487,N_4486);
or U4967 (N_4967,N_4356,N_4394);
nand U4968 (N_4968,N_4109,N_4032);
xnor U4969 (N_4969,N_4375,N_4089);
xnor U4970 (N_4970,N_4302,N_4175);
nand U4971 (N_4971,N_4339,N_4133);
xor U4972 (N_4972,N_4149,N_4391);
xnor U4973 (N_4973,N_4295,N_4104);
or U4974 (N_4974,N_4028,N_4467);
or U4975 (N_4975,N_4041,N_4450);
xnor U4976 (N_4976,N_4004,N_4124);
nand U4977 (N_4977,N_4119,N_4214);
nand U4978 (N_4978,N_4441,N_4143);
nor U4979 (N_4979,N_4093,N_4407);
nor U4980 (N_4980,N_4009,N_4015);
or U4981 (N_4981,N_4057,N_4020);
and U4982 (N_4982,N_4323,N_4335);
nand U4983 (N_4983,N_4021,N_4367);
or U4984 (N_4984,N_4140,N_4165);
or U4985 (N_4985,N_4310,N_4165);
nand U4986 (N_4986,N_4323,N_4090);
nor U4987 (N_4987,N_4315,N_4330);
nand U4988 (N_4988,N_4259,N_4494);
or U4989 (N_4989,N_4199,N_4098);
xnor U4990 (N_4990,N_4131,N_4096);
or U4991 (N_4991,N_4273,N_4120);
xnor U4992 (N_4992,N_4218,N_4208);
and U4993 (N_4993,N_4238,N_4327);
nor U4994 (N_4994,N_4161,N_4096);
nor U4995 (N_4995,N_4054,N_4007);
or U4996 (N_4996,N_4317,N_4491);
xnor U4997 (N_4997,N_4397,N_4370);
xnor U4998 (N_4998,N_4414,N_4035);
nor U4999 (N_4999,N_4263,N_4245);
or U5000 (N_5000,N_4883,N_4876);
nor U5001 (N_5001,N_4763,N_4648);
nand U5002 (N_5002,N_4692,N_4867);
and U5003 (N_5003,N_4875,N_4540);
and U5004 (N_5004,N_4842,N_4793);
or U5005 (N_5005,N_4994,N_4739);
xnor U5006 (N_5006,N_4884,N_4526);
and U5007 (N_5007,N_4962,N_4957);
or U5008 (N_5008,N_4581,N_4528);
nor U5009 (N_5009,N_4986,N_4514);
nor U5010 (N_5010,N_4683,N_4885);
nor U5011 (N_5011,N_4729,N_4605);
nor U5012 (N_5012,N_4714,N_4592);
nand U5013 (N_5013,N_4837,N_4970);
nor U5014 (N_5014,N_4780,N_4652);
or U5015 (N_5015,N_4636,N_4621);
xnor U5016 (N_5016,N_4985,N_4787);
or U5017 (N_5017,N_4690,N_4678);
and U5018 (N_5018,N_4852,N_4749);
nor U5019 (N_5019,N_4944,N_4667);
nor U5020 (N_5020,N_4956,N_4688);
or U5021 (N_5021,N_4757,N_4608);
or U5022 (N_5022,N_4845,N_4762);
xor U5023 (N_5023,N_4542,N_4795);
and U5024 (N_5024,N_4719,N_4822);
or U5025 (N_5025,N_4811,N_4788);
or U5026 (N_5026,N_4784,N_4538);
nand U5027 (N_5027,N_4742,N_4825);
or U5028 (N_5028,N_4868,N_4503);
xor U5029 (N_5029,N_4653,N_4949);
nor U5030 (N_5030,N_4611,N_4619);
nor U5031 (N_5031,N_4930,N_4596);
xor U5032 (N_5032,N_4789,N_4534);
or U5033 (N_5033,N_4858,N_4992);
and U5034 (N_5034,N_4857,N_4946);
and U5035 (N_5035,N_4551,N_4800);
nand U5036 (N_5036,N_4576,N_4643);
or U5037 (N_5037,N_4897,N_4715);
or U5038 (N_5038,N_4703,N_4532);
xnor U5039 (N_5039,N_4604,N_4718);
nor U5040 (N_5040,N_4748,N_4755);
nand U5041 (N_5041,N_4623,N_4910);
xor U5042 (N_5042,N_4568,N_4732);
and U5043 (N_5043,N_4921,N_4695);
or U5044 (N_5044,N_4569,N_4754);
xor U5045 (N_5045,N_4824,N_4924);
or U5046 (N_5046,N_4785,N_4600);
nand U5047 (N_5047,N_4524,N_4812);
xor U5048 (N_5048,N_4878,N_4737);
nor U5049 (N_5049,N_4774,N_4996);
or U5050 (N_5050,N_4848,N_4861);
and U5051 (N_5051,N_4819,N_4575);
nand U5052 (N_5052,N_4846,N_4507);
xor U5053 (N_5053,N_4877,N_4658);
nand U5054 (N_5054,N_4676,N_4829);
nand U5055 (N_5055,N_4593,N_4726);
and U5056 (N_5056,N_4839,N_4738);
or U5057 (N_5057,N_4873,N_4736);
nor U5058 (N_5058,N_4505,N_4973);
nor U5059 (N_5059,N_4660,N_4555);
or U5060 (N_5060,N_4508,N_4993);
and U5061 (N_5061,N_4566,N_4934);
or U5062 (N_5062,N_4646,N_4642);
nand U5063 (N_5063,N_4898,N_4571);
or U5064 (N_5064,N_4834,N_4937);
xnor U5065 (N_5065,N_4630,N_4533);
nor U5066 (N_5066,N_4632,N_4606);
xor U5067 (N_5067,N_4797,N_4974);
or U5068 (N_5068,N_4908,N_4655);
and U5069 (N_5069,N_4887,N_4585);
nor U5070 (N_5070,N_4947,N_4645);
or U5071 (N_5071,N_4833,N_4556);
nand U5072 (N_5072,N_4727,N_4798);
nor U5073 (N_5073,N_4756,N_4603);
xnor U5074 (N_5074,N_4955,N_4782);
and U5075 (N_5075,N_4548,N_4693);
nand U5076 (N_5076,N_4740,N_4933);
and U5077 (N_5077,N_4620,N_4892);
or U5078 (N_5078,N_4982,N_4664);
nor U5079 (N_5079,N_4983,N_4677);
xor U5080 (N_5080,N_4851,N_4708);
nand U5081 (N_5081,N_4654,N_4778);
and U5082 (N_5082,N_4720,N_4586);
or U5083 (N_5083,N_4938,N_4779);
and U5084 (N_5084,N_4886,N_4731);
or U5085 (N_5085,N_4511,N_4768);
and U5086 (N_5086,N_4953,N_4689);
nor U5087 (N_5087,N_4578,N_4869);
and U5088 (N_5088,N_4670,N_4549);
nand U5089 (N_5089,N_4672,N_4554);
nor U5090 (N_5090,N_4753,N_4691);
nor U5091 (N_5091,N_4510,N_4988);
nor U5092 (N_5092,N_4502,N_4767);
nand U5093 (N_5093,N_4951,N_4669);
or U5094 (N_5094,N_4635,N_4577);
or U5095 (N_5095,N_4684,N_4710);
and U5096 (N_5096,N_4866,N_4790);
and U5097 (N_5097,N_4843,N_4971);
xnor U5098 (N_5098,N_4765,N_4500);
nand U5099 (N_5099,N_4871,N_4948);
and U5100 (N_5100,N_4929,N_4960);
nand U5101 (N_5101,N_4995,N_4709);
xnor U5102 (N_5102,N_4583,N_4560);
xor U5103 (N_5103,N_4922,N_4650);
nor U5104 (N_5104,N_4850,N_4711);
xnor U5105 (N_5105,N_4896,N_4844);
nor U5106 (N_5106,N_4639,N_4706);
and U5107 (N_5107,N_4752,N_4518);
nor U5108 (N_5108,N_4570,N_4882);
or U5109 (N_5109,N_4598,N_4751);
xnor U5110 (N_5110,N_4859,N_4814);
nand U5111 (N_5111,N_4890,N_4856);
xnor U5112 (N_5112,N_4794,N_4580);
and U5113 (N_5113,N_4567,N_4716);
nand U5114 (N_5114,N_4546,N_4745);
xor U5115 (N_5115,N_4997,N_4972);
or U5116 (N_5116,N_4894,N_4904);
nor U5117 (N_5117,N_4806,N_4616);
nand U5118 (N_5118,N_4909,N_4516);
nor U5119 (N_5119,N_4615,N_4622);
nand U5120 (N_5120,N_4584,N_4612);
and U5121 (N_5121,N_4853,N_4981);
or U5122 (N_5122,N_4820,N_4963);
nor U5123 (N_5123,N_4722,N_4668);
or U5124 (N_5124,N_4625,N_4631);
or U5125 (N_5125,N_4573,N_4936);
nand U5126 (N_5126,N_4657,N_4928);
nor U5127 (N_5127,N_4865,N_4893);
xor U5128 (N_5128,N_4557,N_4969);
xor U5129 (N_5129,N_4519,N_4772);
nor U5130 (N_5130,N_4582,N_4815);
nand U5131 (N_5131,N_4966,N_4527);
nor U5132 (N_5132,N_4881,N_4671);
nand U5133 (N_5133,N_4792,N_4515);
nor U5134 (N_5134,N_4541,N_4563);
and U5135 (N_5135,N_4545,N_4680);
xnor U5136 (N_5136,N_4818,N_4607);
xnor U5137 (N_5137,N_4553,N_4590);
nor U5138 (N_5138,N_4942,N_4939);
or U5139 (N_5139,N_4597,N_4879);
nor U5140 (N_5140,N_4624,N_4906);
or U5141 (N_5141,N_4991,N_4707);
nand U5142 (N_5142,N_4649,N_4665);
xor U5143 (N_5143,N_4945,N_4950);
and U5144 (N_5144,N_4591,N_4771);
nand U5145 (N_5145,N_4805,N_4796);
or U5146 (N_5146,N_4705,N_4803);
or U5147 (N_5147,N_4529,N_4558);
xor U5148 (N_5148,N_4899,N_4888);
nor U5149 (N_5149,N_4698,N_4987);
xor U5150 (N_5150,N_4759,N_4728);
nand U5151 (N_5151,N_4629,N_4874);
nand U5152 (N_5152,N_4562,N_4651);
or U5153 (N_5153,N_4958,N_4823);
or U5154 (N_5154,N_4730,N_4661);
or U5155 (N_5155,N_4506,N_4564);
or U5156 (N_5156,N_4535,N_4531);
xnor U5157 (N_5157,N_4517,N_4697);
nand U5158 (N_5158,N_4854,N_4901);
nand U5159 (N_5159,N_4968,N_4828);
or U5160 (N_5160,N_4952,N_4675);
and U5161 (N_5161,N_4862,N_4513);
nand U5162 (N_5162,N_4830,N_4918);
nor U5163 (N_5163,N_4595,N_4640);
and U5164 (N_5164,N_4864,N_4810);
nor U5165 (N_5165,N_4685,N_4610);
nor U5166 (N_5166,N_4773,N_4523);
nand U5167 (N_5167,N_4943,N_4932);
nand U5168 (N_5168,N_4589,N_4594);
and U5169 (N_5169,N_4602,N_4501);
or U5170 (N_5170,N_4537,N_4704);
or U5171 (N_5171,N_4965,N_4679);
nor U5172 (N_5172,N_4601,N_4723);
nor U5173 (N_5173,N_4978,N_4641);
nor U5174 (N_5174,N_4786,N_4725);
xor U5175 (N_5175,N_4666,N_4746);
or U5176 (N_5176,N_4832,N_4916);
nand U5177 (N_5177,N_4860,N_4976);
nor U5178 (N_5178,N_4741,N_4760);
xnor U5179 (N_5179,N_4801,N_4809);
and U5180 (N_5180,N_4764,N_4637);
nor U5181 (N_5181,N_4574,N_4552);
and U5182 (N_5182,N_4903,N_4917);
and U5183 (N_5183,N_4758,N_4686);
nor U5184 (N_5184,N_4539,N_4587);
nand U5185 (N_5185,N_4872,N_4980);
xor U5186 (N_5186,N_4599,N_4849);
nand U5187 (N_5187,N_4925,N_4847);
nor U5188 (N_5188,N_4659,N_4628);
or U5189 (N_5189,N_4813,N_4913);
nand U5190 (N_5190,N_4544,N_4975);
and U5191 (N_5191,N_4799,N_4776);
and U5192 (N_5192,N_4699,N_4734);
xnor U5193 (N_5193,N_4712,N_4579);
nor U5194 (N_5194,N_4735,N_4550);
nand U5195 (N_5195,N_4713,N_4536);
or U5196 (N_5196,N_4961,N_4990);
and U5197 (N_5197,N_4935,N_4681);
or U5198 (N_5198,N_4900,N_4804);
nand U5199 (N_5199,N_4831,N_4701);
nor U5200 (N_5200,N_4733,N_4572);
and U5201 (N_5201,N_4941,N_4902);
and U5202 (N_5202,N_4919,N_4998);
xnor U5203 (N_5203,N_4907,N_4769);
or U5204 (N_5204,N_4721,N_4816);
or U5205 (N_5205,N_4617,N_4520);
nand U5206 (N_5206,N_4559,N_4770);
or U5207 (N_5207,N_4870,N_4694);
xor U5208 (N_5208,N_4821,N_4880);
nand U5209 (N_5209,N_4863,N_4840);
nor U5210 (N_5210,N_4530,N_4895);
xnor U5211 (N_5211,N_4626,N_4743);
nand U5212 (N_5212,N_4977,N_4808);
nor U5213 (N_5213,N_4512,N_4940);
or U5214 (N_5214,N_4791,N_4912);
nand U5215 (N_5215,N_4855,N_4525);
or U5216 (N_5216,N_4989,N_4979);
nor U5217 (N_5217,N_4724,N_4702);
nand U5218 (N_5218,N_4644,N_4588);
or U5219 (N_5219,N_4999,N_4634);
nor U5220 (N_5220,N_4747,N_4783);
nand U5221 (N_5221,N_4905,N_4744);
nand U5222 (N_5222,N_4781,N_4633);
nand U5223 (N_5223,N_4777,N_4638);
and U5224 (N_5224,N_4802,N_4817);
or U5225 (N_5225,N_4682,N_4521);
and U5226 (N_5226,N_4522,N_4662);
nor U5227 (N_5227,N_4964,N_4609);
nor U5228 (N_5228,N_4614,N_4766);
or U5229 (N_5229,N_4967,N_4838);
nand U5230 (N_5230,N_4761,N_4889);
nand U5231 (N_5231,N_4841,N_4959);
or U5232 (N_5232,N_4547,N_4835);
and U5233 (N_5233,N_4915,N_4509);
or U5234 (N_5234,N_4647,N_4656);
or U5235 (N_5235,N_4807,N_4914);
nand U5236 (N_5236,N_4920,N_4613);
or U5237 (N_5237,N_4927,N_4504);
nor U5238 (N_5238,N_4673,N_4926);
or U5239 (N_5239,N_4561,N_4627);
nand U5240 (N_5240,N_4931,N_4827);
nand U5241 (N_5241,N_4923,N_4618);
nand U5242 (N_5242,N_4891,N_4696);
or U5243 (N_5243,N_4954,N_4565);
nand U5244 (N_5244,N_4543,N_4663);
nand U5245 (N_5245,N_4911,N_4826);
xor U5246 (N_5246,N_4984,N_4700);
xnor U5247 (N_5247,N_4750,N_4836);
or U5248 (N_5248,N_4775,N_4687);
or U5249 (N_5249,N_4674,N_4717);
and U5250 (N_5250,N_4863,N_4608);
and U5251 (N_5251,N_4521,N_4717);
xnor U5252 (N_5252,N_4594,N_4579);
xnor U5253 (N_5253,N_4700,N_4685);
or U5254 (N_5254,N_4772,N_4506);
nand U5255 (N_5255,N_4907,N_4860);
xor U5256 (N_5256,N_4716,N_4591);
and U5257 (N_5257,N_4523,N_4684);
or U5258 (N_5258,N_4965,N_4664);
nor U5259 (N_5259,N_4747,N_4952);
or U5260 (N_5260,N_4898,N_4824);
xor U5261 (N_5261,N_4658,N_4651);
nand U5262 (N_5262,N_4778,N_4810);
nand U5263 (N_5263,N_4791,N_4895);
xor U5264 (N_5264,N_4924,N_4821);
or U5265 (N_5265,N_4596,N_4844);
nor U5266 (N_5266,N_4800,N_4920);
or U5267 (N_5267,N_4850,N_4930);
or U5268 (N_5268,N_4648,N_4971);
nand U5269 (N_5269,N_4973,N_4942);
nor U5270 (N_5270,N_4527,N_4723);
nor U5271 (N_5271,N_4700,N_4550);
or U5272 (N_5272,N_4674,N_4536);
nor U5273 (N_5273,N_4642,N_4634);
nor U5274 (N_5274,N_4648,N_4568);
nor U5275 (N_5275,N_4716,N_4803);
nor U5276 (N_5276,N_4972,N_4638);
nor U5277 (N_5277,N_4830,N_4712);
nor U5278 (N_5278,N_4639,N_4801);
nand U5279 (N_5279,N_4645,N_4887);
nor U5280 (N_5280,N_4660,N_4597);
nand U5281 (N_5281,N_4779,N_4613);
and U5282 (N_5282,N_4823,N_4570);
or U5283 (N_5283,N_4881,N_4754);
nand U5284 (N_5284,N_4727,N_4543);
or U5285 (N_5285,N_4817,N_4962);
xor U5286 (N_5286,N_4529,N_4957);
and U5287 (N_5287,N_4709,N_4948);
nor U5288 (N_5288,N_4924,N_4555);
or U5289 (N_5289,N_4788,N_4748);
nand U5290 (N_5290,N_4931,N_4895);
nor U5291 (N_5291,N_4949,N_4980);
and U5292 (N_5292,N_4681,N_4937);
and U5293 (N_5293,N_4793,N_4976);
nor U5294 (N_5294,N_4551,N_4987);
or U5295 (N_5295,N_4705,N_4814);
and U5296 (N_5296,N_4672,N_4546);
and U5297 (N_5297,N_4916,N_4814);
nand U5298 (N_5298,N_4511,N_4991);
or U5299 (N_5299,N_4837,N_4869);
and U5300 (N_5300,N_4934,N_4940);
and U5301 (N_5301,N_4782,N_4666);
or U5302 (N_5302,N_4658,N_4931);
nor U5303 (N_5303,N_4928,N_4540);
xnor U5304 (N_5304,N_4758,N_4894);
and U5305 (N_5305,N_4655,N_4853);
nor U5306 (N_5306,N_4951,N_4847);
nand U5307 (N_5307,N_4987,N_4639);
and U5308 (N_5308,N_4871,N_4839);
nor U5309 (N_5309,N_4816,N_4688);
xnor U5310 (N_5310,N_4767,N_4844);
and U5311 (N_5311,N_4767,N_4709);
nand U5312 (N_5312,N_4707,N_4605);
and U5313 (N_5313,N_4753,N_4647);
or U5314 (N_5314,N_4691,N_4832);
nor U5315 (N_5315,N_4822,N_4958);
xnor U5316 (N_5316,N_4822,N_4905);
and U5317 (N_5317,N_4898,N_4836);
nand U5318 (N_5318,N_4705,N_4513);
nand U5319 (N_5319,N_4968,N_4762);
xor U5320 (N_5320,N_4808,N_4965);
and U5321 (N_5321,N_4867,N_4670);
or U5322 (N_5322,N_4910,N_4757);
xnor U5323 (N_5323,N_4925,N_4705);
and U5324 (N_5324,N_4644,N_4670);
nand U5325 (N_5325,N_4918,N_4834);
or U5326 (N_5326,N_4552,N_4819);
or U5327 (N_5327,N_4666,N_4949);
nand U5328 (N_5328,N_4687,N_4505);
nand U5329 (N_5329,N_4724,N_4582);
and U5330 (N_5330,N_4918,N_4827);
xor U5331 (N_5331,N_4899,N_4935);
xor U5332 (N_5332,N_4896,N_4868);
nor U5333 (N_5333,N_4992,N_4556);
nand U5334 (N_5334,N_4544,N_4814);
nor U5335 (N_5335,N_4580,N_4608);
nand U5336 (N_5336,N_4792,N_4584);
nor U5337 (N_5337,N_4748,N_4884);
nor U5338 (N_5338,N_4804,N_4690);
xnor U5339 (N_5339,N_4979,N_4820);
or U5340 (N_5340,N_4779,N_4814);
xor U5341 (N_5341,N_4636,N_4661);
or U5342 (N_5342,N_4508,N_4985);
and U5343 (N_5343,N_4793,N_4881);
xnor U5344 (N_5344,N_4687,N_4568);
nand U5345 (N_5345,N_4612,N_4720);
xor U5346 (N_5346,N_4715,N_4509);
or U5347 (N_5347,N_4758,N_4949);
and U5348 (N_5348,N_4662,N_4900);
nor U5349 (N_5349,N_4861,N_4921);
xnor U5350 (N_5350,N_4821,N_4575);
and U5351 (N_5351,N_4704,N_4605);
nand U5352 (N_5352,N_4842,N_4586);
nor U5353 (N_5353,N_4682,N_4677);
or U5354 (N_5354,N_4844,N_4989);
xnor U5355 (N_5355,N_4526,N_4647);
xnor U5356 (N_5356,N_4909,N_4618);
nor U5357 (N_5357,N_4591,N_4588);
xnor U5358 (N_5358,N_4813,N_4950);
xor U5359 (N_5359,N_4755,N_4876);
or U5360 (N_5360,N_4510,N_4846);
xnor U5361 (N_5361,N_4910,N_4974);
nor U5362 (N_5362,N_4907,N_4637);
or U5363 (N_5363,N_4613,N_4685);
or U5364 (N_5364,N_4908,N_4702);
or U5365 (N_5365,N_4945,N_4673);
and U5366 (N_5366,N_4721,N_4891);
xnor U5367 (N_5367,N_4500,N_4597);
nand U5368 (N_5368,N_4676,N_4681);
or U5369 (N_5369,N_4637,N_4576);
and U5370 (N_5370,N_4992,N_4692);
nand U5371 (N_5371,N_4928,N_4643);
nand U5372 (N_5372,N_4902,N_4998);
nor U5373 (N_5373,N_4607,N_4991);
nand U5374 (N_5374,N_4929,N_4603);
nand U5375 (N_5375,N_4594,N_4718);
or U5376 (N_5376,N_4587,N_4852);
or U5377 (N_5377,N_4645,N_4680);
and U5378 (N_5378,N_4607,N_4963);
nand U5379 (N_5379,N_4741,N_4528);
nand U5380 (N_5380,N_4953,N_4936);
or U5381 (N_5381,N_4802,N_4713);
and U5382 (N_5382,N_4558,N_4722);
nor U5383 (N_5383,N_4886,N_4565);
nor U5384 (N_5384,N_4734,N_4971);
nor U5385 (N_5385,N_4852,N_4824);
xnor U5386 (N_5386,N_4663,N_4959);
or U5387 (N_5387,N_4685,N_4806);
xor U5388 (N_5388,N_4978,N_4758);
or U5389 (N_5389,N_4505,N_4605);
and U5390 (N_5390,N_4946,N_4663);
xnor U5391 (N_5391,N_4634,N_4648);
nor U5392 (N_5392,N_4663,N_4671);
nand U5393 (N_5393,N_4768,N_4931);
xnor U5394 (N_5394,N_4856,N_4754);
nand U5395 (N_5395,N_4864,N_4668);
nand U5396 (N_5396,N_4884,N_4988);
nand U5397 (N_5397,N_4648,N_4729);
xnor U5398 (N_5398,N_4850,N_4517);
or U5399 (N_5399,N_4915,N_4795);
xor U5400 (N_5400,N_4694,N_4620);
nand U5401 (N_5401,N_4970,N_4728);
xor U5402 (N_5402,N_4993,N_4767);
xor U5403 (N_5403,N_4688,N_4930);
nand U5404 (N_5404,N_4849,N_4810);
nand U5405 (N_5405,N_4765,N_4563);
or U5406 (N_5406,N_4683,N_4953);
xor U5407 (N_5407,N_4788,N_4614);
or U5408 (N_5408,N_4714,N_4627);
and U5409 (N_5409,N_4779,N_4922);
or U5410 (N_5410,N_4997,N_4955);
nand U5411 (N_5411,N_4535,N_4552);
or U5412 (N_5412,N_4530,N_4893);
xnor U5413 (N_5413,N_4754,N_4532);
or U5414 (N_5414,N_4566,N_4914);
or U5415 (N_5415,N_4991,N_4546);
nand U5416 (N_5416,N_4948,N_4965);
and U5417 (N_5417,N_4990,N_4561);
nor U5418 (N_5418,N_4601,N_4680);
or U5419 (N_5419,N_4958,N_4876);
nor U5420 (N_5420,N_4918,N_4941);
or U5421 (N_5421,N_4599,N_4805);
xor U5422 (N_5422,N_4900,N_4536);
or U5423 (N_5423,N_4906,N_4852);
and U5424 (N_5424,N_4623,N_4866);
or U5425 (N_5425,N_4774,N_4596);
nor U5426 (N_5426,N_4732,N_4759);
and U5427 (N_5427,N_4750,N_4515);
or U5428 (N_5428,N_4790,N_4725);
nand U5429 (N_5429,N_4522,N_4943);
nand U5430 (N_5430,N_4780,N_4528);
nand U5431 (N_5431,N_4605,N_4920);
nand U5432 (N_5432,N_4871,N_4968);
nor U5433 (N_5433,N_4782,N_4523);
xor U5434 (N_5434,N_4904,N_4864);
nor U5435 (N_5435,N_4550,N_4629);
nor U5436 (N_5436,N_4859,N_4561);
xnor U5437 (N_5437,N_4854,N_4646);
and U5438 (N_5438,N_4565,N_4572);
xnor U5439 (N_5439,N_4545,N_4556);
nand U5440 (N_5440,N_4595,N_4884);
and U5441 (N_5441,N_4987,N_4730);
nor U5442 (N_5442,N_4930,N_4629);
nor U5443 (N_5443,N_4915,N_4995);
and U5444 (N_5444,N_4739,N_4998);
or U5445 (N_5445,N_4754,N_4577);
and U5446 (N_5446,N_4715,N_4522);
nor U5447 (N_5447,N_4951,N_4718);
nor U5448 (N_5448,N_4507,N_4708);
nand U5449 (N_5449,N_4583,N_4982);
and U5450 (N_5450,N_4819,N_4712);
or U5451 (N_5451,N_4512,N_4664);
nand U5452 (N_5452,N_4927,N_4814);
nor U5453 (N_5453,N_4608,N_4958);
nand U5454 (N_5454,N_4736,N_4829);
nor U5455 (N_5455,N_4795,N_4973);
or U5456 (N_5456,N_4980,N_4773);
and U5457 (N_5457,N_4707,N_4868);
or U5458 (N_5458,N_4925,N_4762);
and U5459 (N_5459,N_4914,N_4671);
or U5460 (N_5460,N_4598,N_4926);
xor U5461 (N_5461,N_4701,N_4844);
and U5462 (N_5462,N_4941,N_4516);
xor U5463 (N_5463,N_4943,N_4998);
nor U5464 (N_5464,N_4807,N_4773);
xor U5465 (N_5465,N_4767,N_4606);
and U5466 (N_5466,N_4688,N_4616);
and U5467 (N_5467,N_4706,N_4925);
or U5468 (N_5468,N_4708,N_4920);
nand U5469 (N_5469,N_4973,N_4815);
nand U5470 (N_5470,N_4944,N_4664);
nand U5471 (N_5471,N_4977,N_4704);
nand U5472 (N_5472,N_4824,N_4953);
and U5473 (N_5473,N_4607,N_4662);
nor U5474 (N_5474,N_4738,N_4930);
nand U5475 (N_5475,N_4611,N_4870);
xor U5476 (N_5476,N_4821,N_4930);
nand U5477 (N_5477,N_4522,N_4728);
nand U5478 (N_5478,N_4898,N_4621);
nand U5479 (N_5479,N_4742,N_4542);
xor U5480 (N_5480,N_4992,N_4781);
and U5481 (N_5481,N_4635,N_4506);
or U5482 (N_5482,N_4564,N_4584);
nor U5483 (N_5483,N_4906,N_4937);
nor U5484 (N_5484,N_4972,N_4607);
or U5485 (N_5485,N_4614,N_4696);
or U5486 (N_5486,N_4888,N_4607);
xor U5487 (N_5487,N_4639,N_4894);
or U5488 (N_5488,N_4945,N_4962);
nand U5489 (N_5489,N_4669,N_4522);
nor U5490 (N_5490,N_4604,N_4875);
or U5491 (N_5491,N_4916,N_4761);
nor U5492 (N_5492,N_4593,N_4623);
and U5493 (N_5493,N_4870,N_4645);
xor U5494 (N_5494,N_4694,N_4800);
xor U5495 (N_5495,N_4658,N_4600);
or U5496 (N_5496,N_4840,N_4563);
and U5497 (N_5497,N_4837,N_4729);
or U5498 (N_5498,N_4958,N_4762);
or U5499 (N_5499,N_4844,N_4588);
or U5500 (N_5500,N_5316,N_5418);
or U5501 (N_5501,N_5449,N_5045);
nor U5502 (N_5502,N_5168,N_5098);
nor U5503 (N_5503,N_5074,N_5201);
and U5504 (N_5504,N_5132,N_5269);
nand U5505 (N_5505,N_5477,N_5120);
xor U5506 (N_5506,N_5297,N_5333);
or U5507 (N_5507,N_5411,N_5178);
nand U5508 (N_5508,N_5003,N_5052);
nor U5509 (N_5509,N_5210,N_5208);
nand U5510 (N_5510,N_5092,N_5001);
nand U5511 (N_5511,N_5066,N_5007);
xnor U5512 (N_5512,N_5390,N_5101);
xnor U5513 (N_5513,N_5313,N_5249);
xor U5514 (N_5514,N_5474,N_5348);
xor U5515 (N_5515,N_5166,N_5028);
or U5516 (N_5516,N_5401,N_5457);
or U5517 (N_5517,N_5350,N_5085);
xnor U5518 (N_5518,N_5406,N_5072);
xor U5519 (N_5519,N_5374,N_5375);
or U5520 (N_5520,N_5135,N_5194);
xor U5521 (N_5521,N_5460,N_5343);
and U5522 (N_5522,N_5290,N_5469);
nand U5523 (N_5523,N_5090,N_5109);
nand U5524 (N_5524,N_5219,N_5421);
nor U5525 (N_5525,N_5499,N_5405);
nand U5526 (N_5526,N_5018,N_5145);
nor U5527 (N_5527,N_5429,N_5339);
or U5528 (N_5528,N_5044,N_5288);
and U5529 (N_5529,N_5464,N_5450);
and U5530 (N_5530,N_5142,N_5407);
or U5531 (N_5531,N_5461,N_5383);
and U5532 (N_5532,N_5041,N_5032);
nor U5533 (N_5533,N_5364,N_5211);
xnor U5534 (N_5534,N_5139,N_5177);
xnor U5535 (N_5535,N_5004,N_5221);
nor U5536 (N_5536,N_5199,N_5054);
nand U5537 (N_5537,N_5227,N_5015);
xor U5538 (N_5538,N_5012,N_5481);
or U5539 (N_5539,N_5257,N_5384);
nor U5540 (N_5540,N_5209,N_5344);
or U5541 (N_5541,N_5062,N_5472);
or U5542 (N_5542,N_5002,N_5238);
xor U5543 (N_5543,N_5053,N_5233);
nand U5544 (N_5544,N_5282,N_5129);
xnor U5545 (N_5545,N_5340,N_5315);
and U5546 (N_5546,N_5200,N_5428);
and U5547 (N_5547,N_5019,N_5058);
xor U5548 (N_5548,N_5439,N_5059);
xnor U5549 (N_5549,N_5274,N_5448);
nor U5550 (N_5550,N_5356,N_5320);
nor U5551 (N_5551,N_5043,N_5244);
nand U5552 (N_5552,N_5268,N_5106);
and U5553 (N_5553,N_5079,N_5223);
and U5554 (N_5554,N_5498,N_5115);
xor U5555 (N_5555,N_5281,N_5488);
xnor U5556 (N_5556,N_5061,N_5033);
and U5557 (N_5557,N_5330,N_5251);
nor U5558 (N_5558,N_5084,N_5089);
nand U5559 (N_5559,N_5110,N_5189);
or U5560 (N_5560,N_5172,N_5413);
and U5561 (N_5561,N_5185,N_5373);
nor U5562 (N_5562,N_5380,N_5453);
and U5563 (N_5563,N_5430,N_5321);
xnor U5564 (N_5564,N_5496,N_5262);
and U5565 (N_5565,N_5463,N_5051);
xnor U5566 (N_5566,N_5250,N_5036);
xnor U5567 (N_5567,N_5377,N_5347);
nor U5568 (N_5568,N_5403,N_5049);
nor U5569 (N_5569,N_5076,N_5196);
or U5570 (N_5570,N_5048,N_5021);
nor U5571 (N_5571,N_5363,N_5337);
nand U5572 (N_5572,N_5395,N_5497);
or U5573 (N_5573,N_5265,N_5157);
xnor U5574 (N_5574,N_5217,N_5197);
and U5575 (N_5575,N_5216,N_5327);
nand U5576 (N_5576,N_5434,N_5010);
xor U5577 (N_5577,N_5186,N_5482);
nor U5578 (N_5578,N_5080,N_5171);
nand U5579 (N_5579,N_5292,N_5191);
and U5580 (N_5580,N_5070,N_5494);
nor U5581 (N_5581,N_5286,N_5338);
nor U5582 (N_5582,N_5277,N_5241);
nor U5583 (N_5583,N_5298,N_5133);
xor U5584 (N_5584,N_5471,N_5314);
and U5585 (N_5585,N_5273,N_5475);
nor U5586 (N_5586,N_5423,N_5385);
nor U5587 (N_5587,N_5311,N_5440);
nor U5588 (N_5588,N_5393,N_5355);
and U5589 (N_5589,N_5151,N_5276);
and U5590 (N_5590,N_5170,N_5358);
or U5591 (N_5591,N_5240,N_5322);
nor U5592 (N_5592,N_5014,N_5468);
xnor U5593 (N_5593,N_5005,N_5218);
nor U5594 (N_5594,N_5400,N_5409);
nand U5595 (N_5595,N_5317,N_5144);
and U5596 (N_5596,N_5285,N_5427);
xnor U5597 (N_5597,N_5202,N_5328);
and U5598 (N_5598,N_5131,N_5404);
and U5599 (N_5599,N_5324,N_5220);
and U5600 (N_5600,N_5180,N_5035);
xor U5601 (N_5601,N_5183,N_5352);
nor U5602 (N_5602,N_5027,N_5181);
or U5603 (N_5603,N_5122,N_5303);
xor U5604 (N_5604,N_5226,N_5212);
or U5605 (N_5605,N_5483,N_5091);
or U5606 (N_5606,N_5071,N_5039);
or U5607 (N_5607,N_5153,N_5462);
nand U5608 (N_5608,N_5077,N_5150);
and U5609 (N_5609,N_5239,N_5064);
nor U5610 (N_5610,N_5459,N_5253);
xnor U5611 (N_5611,N_5466,N_5243);
or U5612 (N_5612,N_5230,N_5067);
or U5613 (N_5613,N_5480,N_5417);
nor U5614 (N_5614,N_5068,N_5422);
and U5615 (N_5615,N_5376,N_5437);
and U5616 (N_5616,N_5308,N_5394);
nor U5617 (N_5617,N_5368,N_5305);
nand U5618 (N_5618,N_5055,N_5029);
nand U5619 (N_5619,N_5312,N_5367);
and U5620 (N_5620,N_5278,N_5159);
xnor U5621 (N_5621,N_5161,N_5294);
nand U5622 (N_5622,N_5379,N_5047);
and U5623 (N_5623,N_5088,N_5037);
xnor U5624 (N_5624,N_5451,N_5438);
nand U5625 (N_5625,N_5456,N_5100);
or U5626 (N_5626,N_5366,N_5030);
and U5627 (N_5627,N_5458,N_5432);
nand U5628 (N_5628,N_5095,N_5491);
nand U5629 (N_5629,N_5040,N_5280);
or U5630 (N_5630,N_5152,N_5114);
nor U5631 (N_5631,N_5302,N_5046);
nor U5632 (N_5632,N_5446,N_5065);
and U5633 (N_5633,N_5369,N_5073);
nand U5634 (N_5634,N_5431,N_5473);
or U5635 (N_5635,N_5093,N_5156);
and U5636 (N_5636,N_5031,N_5354);
or U5637 (N_5637,N_5025,N_5104);
or U5638 (N_5638,N_5341,N_5165);
nand U5639 (N_5639,N_5126,N_5108);
or U5640 (N_5640,N_5301,N_5082);
or U5641 (N_5641,N_5214,N_5195);
nor U5642 (N_5642,N_5174,N_5184);
nor U5643 (N_5643,N_5487,N_5078);
nand U5644 (N_5644,N_5228,N_5293);
nand U5645 (N_5645,N_5397,N_5179);
nand U5646 (N_5646,N_5017,N_5130);
nand U5647 (N_5647,N_5489,N_5198);
nand U5648 (N_5648,N_5266,N_5231);
nor U5649 (N_5649,N_5204,N_5336);
xnor U5650 (N_5650,N_5163,N_5300);
xnor U5651 (N_5651,N_5329,N_5479);
nand U5652 (N_5652,N_5111,N_5096);
nand U5653 (N_5653,N_5207,N_5291);
xor U5654 (N_5654,N_5094,N_5123);
nand U5655 (N_5655,N_5441,N_5478);
and U5656 (N_5656,N_5206,N_5024);
or U5657 (N_5657,N_5299,N_5193);
or U5658 (N_5658,N_5325,N_5470);
xor U5659 (N_5659,N_5103,N_5175);
and U5660 (N_5660,N_5020,N_5391);
nor U5661 (N_5661,N_5442,N_5307);
and U5662 (N_5662,N_5008,N_5245);
nor U5663 (N_5663,N_5099,N_5234);
and U5664 (N_5664,N_5236,N_5396);
nand U5665 (N_5665,N_5215,N_5097);
nor U5666 (N_5666,N_5270,N_5086);
and U5667 (N_5667,N_5476,N_5435);
and U5668 (N_5668,N_5075,N_5455);
xnor U5669 (N_5669,N_5287,N_5452);
xor U5670 (N_5670,N_5237,N_5335);
xor U5671 (N_5671,N_5107,N_5190);
nand U5672 (N_5672,N_5203,N_5128);
xor U5673 (N_5673,N_5485,N_5022);
or U5674 (N_5674,N_5433,N_5247);
nand U5675 (N_5675,N_5116,N_5034);
nor U5676 (N_5676,N_5414,N_5495);
nor U5677 (N_5677,N_5187,N_5387);
xor U5678 (N_5678,N_5013,N_5147);
or U5679 (N_5679,N_5016,N_5143);
nand U5680 (N_5680,N_5304,N_5399);
nand U5681 (N_5681,N_5454,N_5360);
and U5682 (N_5682,N_5081,N_5362);
and U5683 (N_5683,N_5162,N_5138);
xnor U5684 (N_5684,N_5148,N_5087);
nand U5685 (N_5685,N_5484,N_5056);
and U5686 (N_5686,N_5388,N_5112);
nor U5687 (N_5687,N_5412,N_5365);
or U5688 (N_5688,N_5331,N_5445);
or U5689 (N_5689,N_5349,N_5486);
xnor U5690 (N_5690,N_5121,N_5176);
or U5691 (N_5691,N_5141,N_5370);
or U5692 (N_5692,N_5260,N_5117);
and U5693 (N_5693,N_5000,N_5359);
and U5694 (N_5694,N_5160,N_5158);
nand U5695 (N_5695,N_5275,N_5113);
and U5696 (N_5696,N_5493,N_5125);
nand U5697 (N_5697,N_5261,N_5426);
or U5698 (N_5698,N_5050,N_5083);
nor U5699 (N_5699,N_5222,N_5296);
nand U5700 (N_5700,N_5398,N_5124);
nand U5701 (N_5701,N_5492,N_5134);
nor U5702 (N_5702,N_5416,N_5408);
xnor U5703 (N_5703,N_5255,N_5271);
and U5704 (N_5704,N_5334,N_5382);
nor U5705 (N_5705,N_5490,N_5361);
and U5706 (N_5706,N_5182,N_5279);
and U5707 (N_5707,N_5155,N_5289);
nor U5708 (N_5708,N_5167,N_5467);
nand U5709 (N_5709,N_5272,N_5188);
xor U5710 (N_5710,N_5146,N_5105);
nor U5711 (N_5711,N_5410,N_5425);
xnor U5712 (N_5712,N_5057,N_5154);
or U5713 (N_5713,N_5137,N_5038);
nand U5714 (N_5714,N_5069,N_5323);
nand U5715 (N_5715,N_5192,N_5319);
nand U5716 (N_5716,N_5213,N_5267);
or U5717 (N_5717,N_5140,N_5127);
nor U5718 (N_5718,N_5443,N_5419);
and U5719 (N_5719,N_5436,N_5009);
or U5720 (N_5720,N_5386,N_5415);
nor U5721 (N_5721,N_5042,N_5254);
and U5722 (N_5722,N_5345,N_5295);
or U5723 (N_5723,N_5465,N_5444);
and U5724 (N_5724,N_5205,N_5011);
xnor U5725 (N_5725,N_5246,N_5353);
nor U5726 (N_5726,N_5309,N_5173);
nand U5727 (N_5727,N_5402,N_5371);
and U5728 (N_5728,N_5229,N_5332);
nand U5729 (N_5729,N_5424,N_5284);
or U5730 (N_5730,N_5119,N_5318);
or U5731 (N_5731,N_5420,N_5252);
nand U5732 (N_5732,N_5235,N_5232);
nand U5733 (N_5733,N_5102,N_5006);
or U5734 (N_5734,N_5224,N_5357);
nor U5735 (N_5735,N_5381,N_5326);
or U5736 (N_5736,N_5310,N_5263);
nand U5737 (N_5737,N_5169,N_5063);
nor U5738 (N_5738,N_5225,N_5389);
or U5739 (N_5739,N_5283,N_5259);
nand U5740 (N_5740,N_5023,N_5346);
or U5741 (N_5741,N_5372,N_5342);
and U5742 (N_5742,N_5264,N_5060);
nand U5743 (N_5743,N_5256,N_5136);
nand U5744 (N_5744,N_5378,N_5258);
xor U5745 (N_5745,N_5306,N_5164);
nand U5746 (N_5746,N_5149,N_5447);
or U5747 (N_5747,N_5118,N_5351);
or U5748 (N_5748,N_5026,N_5242);
or U5749 (N_5749,N_5248,N_5392);
nor U5750 (N_5750,N_5159,N_5126);
nand U5751 (N_5751,N_5016,N_5383);
or U5752 (N_5752,N_5381,N_5200);
nand U5753 (N_5753,N_5176,N_5295);
nand U5754 (N_5754,N_5001,N_5238);
nor U5755 (N_5755,N_5397,N_5494);
and U5756 (N_5756,N_5186,N_5051);
nand U5757 (N_5757,N_5289,N_5438);
or U5758 (N_5758,N_5032,N_5117);
nor U5759 (N_5759,N_5416,N_5141);
xor U5760 (N_5760,N_5111,N_5224);
xnor U5761 (N_5761,N_5494,N_5431);
or U5762 (N_5762,N_5253,N_5380);
nand U5763 (N_5763,N_5421,N_5175);
nor U5764 (N_5764,N_5157,N_5070);
and U5765 (N_5765,N_5192,N_5193);
and U5766 (N_5766,N_5203,N_5333);
nor U5767 (N_5767,N_5292,N_5023);
xor U5768 (N_5768,N_5176,N_5422);
nor U5769 (N_5769,N_5147,N_5189);
nand U5770 (N_5770,N_5064,N_5122);
xor U5771 (N_5771,N_5243,N_5120);
nor U5772 (N_5772,N_5468,N_5489);
nor U5773 (N_5773,N_5242,N_5228);
or U5774 (N_5774,N_5487,N_5341);
nand U5775 (N_5775,N_5474,N_5460);
nor U5776 (N_5776,N_5175,N_5311);
xor U5777 (N_5777,N_5416,N_5149);
xnor U5778 (N_5778,N_5376,N_5211);
nor U5779 (N_5779,N_5075,N_5404);
nor U5780 (N_5780,N_5254,N_5344);
and U5781 (N_5781,N_5035,N_5344);
xor U5782 (N_5782,N_5264,N_5364);
xor U5783 (N_5783,N_5430,N_5373);
nor U5784 (N_5784,N_5396,N_5413);
nor U5785 (N_5785,N_5175,N_5301);
or U5786 (N_5786,N_5147,N_5461);
nand U5787 (N_5787,N_5492,N_5189);
nand U5788 (N_5788,N_5418,N_5066);
nand U5789 (N_5789,N_5343,N_5487);
and U5790 (N_5790,N_5426,N_5064);
nor U5791 (N_5791,N_5266,N_5204);
or U5792 (N_5792,N_5188,N_5366);
xnor U5793 (N_5793,N_5365,N_5211);
xnor U5794 (N_5794,N_5067,N_5059);
nor U5795 (N_5795,N_5153,N_5284);
xnor U5796 (N_5796,N_5322,N_5168);
nor U5797 (N_5797,N_5395,N_5455);
and U5798 (N_5798,N_5092,N_5265);
nand U5799 (N_5799,N_5274,N_5497);
xnor U5800 (N_5800,N_5083,N_5435);
xnor U5801 (N_5801,N_5065,N_5032);
xnor U5802 (N_5802,N_5065,N_5059);
xor U5803 (N_5803,N_5446,N_5390);
xnor U5804 (N_5804,N_5483,N_5246);
nand U5805 (N_5805,N_5410,N_5236);
and U5806 (N_5806,N_5128,N_5066);
nor U5807 (N_5807,N_5336,N_5429);
nand U5808 (N_5808,N_5097,N_5420);
or U5809 (N_5809,N_5218,N_5022);
nand U5810 (N_5810,N_5374,N_5068);
xor U5811 (N_5811,N_5180,N_5124);
nand U5812 (N_5812,N_5181,N_5428);
xor U5813 (N_5813,N_5111,N_5392);
and U5814 (N_5814,N_5206,N_5322);
or U5815 (N_5815,N_5034,N_5449);
nor U5816 (N_5816,N_5147,N_5428);
or U5817 (N_5817,N_5252,N_5303);
nand U5818 (N_5818,N_5298,N_5307);
xor U5819 (N_5819,N_5005,N_5012);
nor U5820 (N_5820,N_5050,N_5211);
xor U5821 (N_5821,N_5228,N_5461);
xnor U5822 (N_5822,N_5002,N_5281);
or U5823 (N_5823,N_5477,N_5435);
or U5824 (N_5824,N_5217,N_5457);
nor U5825 (N_5825,N_5027,N_5237);
and U5826 (N_5826,N_5006,N_5352);
nand U5827 (N_5827,N_5423,N_5224);
xor U5828 (N_5828,N_5421,N_5280);
nand U5829 (N_5829,N_5069,N_5257);
nand U5830 (N_5830,N_5365,N_5329);
and U5831 (N_5831,N_5130,N_5346);
nand U5832 (N_5832,N_5127,N_5471);
or U5833 (N_5833,N_5163,N_5308);
or U5834 (N_5834,N_5476,N_5012);
nand U5835 (N_5835,N_5009,N_5216);
and U5836 (N_5836,N_5411,N_5153);
or U5837 (N_5837,N_5393,N_5359);
nor U5838 (N_5838,N_5360,N_5280);
nand U5839 (N_5839,N_5305,N_5014);
nor U5840 (N_5840,N_5136,N_5456);
nand U5841 (N_5841,N_5381,N_5154);
xor U5842 (N_5842,N_5140,N_5185);
and U5843 (N_5843,N_5080,N_5008);
and U5844 (N_5844,N_5346,N_5025);
and U5845 (N_5845,N_5401,N_5102);
or U5846 (N_5846,N_5434,N_5217);
or U5847 (N_5847,N_5029,N_5426);
or U5848 (N_5848,N_5026,N_5436);
xnor U5849 (N_5849,N_5289,N_5359);
nand U5850 (N_5850,N_5072,N_5386);
nor U5851 (N_5851,N_5231,N_5353);
and U5852 (N_5852,N_5273,N_5011);
nand U5853 (N_5853,N_5329,N_5411);
nor U5854 (N_5854,N_5371,N_5215);
and U5855 (N_5855,N_5229,N_5085);
xnor U5856 (N_5856,N_5319,N_5458);
or U5857 (N_5857,N_5005,N_5403);
xnor U5858 (N_5858,N_5435,N_5306);
nand U5859 (N_5859,N_5368,N_5350);
nor U5860 (N_5860,N_5370,N_5313);
or U5861 (N_5861,N_5469,N_5107);
or U5862 (N_5862,N_5161,N_5315);
nor U5863 (N_5863,N_5080,N_5380);
or U5864 (N_5864,N_5247,N_5195);
and U5865 (N_5865,N_5010,N_5330);
and U5866 (N_5866,N_5303,N_5249);
xor U5867 (N_5867,N_5439,N_5258);
nand U5868 (N_5868,N_5419,N_5214);
xnor U5869 (N_5869,N_5433,N_5351);
or U5870 (N_5870,N_5297,N_5229);
and U5871 (N_5871,N_5274,N_5256);
nand U5872 (N_5872,N_5476,N_5234);
nor U5873 (N_5873,N_5288,N_5215);
and U5874 (N_5874,N_5093,N_5198);
or U5875 (N_5875,N_5357,N_5133);
and U5876 (N_5876,N_5401,N_5002);
xor U5877 (N_5877,N_5214,N_5003);
nor U5878 (N_5878,N_5050,N_5060);
nand U5879 (N_5879,N_5160,N_5442);
nand U5880 (N_5880,N_5323,N_5457);
or U5881 (N_5881,N_5474,N_5066);
nand U5882 (N_5882,N_5217,N_5084);
xnor U5883 (N_5883,N_5140,N_5264);
xnor U5884 (N_5884,N_5334,N_5424);
and U5885 (N_5885,N_5001,N_5495);
or U5886 (N_5886,N_5001,N_5421);
xnor U5887 (N_5887,N_5263,N_5328);
nand U5888 (N_5888,N_5139,N_5443);
nand U5889 (N_5889,N_5138,N_5308);
or U5890 (N_5890,N_5076,N_5176);
xor U5891 (N_5891,N_5217,N_5058);
and U5892 (N_5892,N_5197,N_5410);
and U5893 (N_5893,N_5301,N_5445);
or U5894 (N_5894,N_5412,N_5481);
nand U5895 (N_5895,N_5168,N_5060);
nand U5896 (N_5896,N_5214,N_5237);
xor U5897 (N_5897,N_5282,N_5279);
and U5898 (N_5898,N_5484,N_5121);
nor U5899 (N_5899,N_5074,N_5007);
nand U5900 (N_5900,N_5447,N_5363);
nand U5901 (N_5901,N_5302,N_5266);
or U5902 (N_5902,N_5432,N_5393);
xnor U5903 (N_5903,N_5116,N_5232);
and U5904 (N_5904,N_5441,N_5130);
or U5905 (N_5905,N_5105,N_5303);
xnor U5906 (N_5906,N_5372,N_5410);
nor U5907 (N_5907,N_5406,N_5376);
and U5908 (N_5908,N_5010,N_5017);
or U5909 (N_5909,N_5163,N_5098);
nand U5910 (N_5910,N_5410,N_5166);
xnor U5911 (N_5911,N_5380,N_5165);
xnor U5912 (N_5912,N_5298,N_5004);
xor U5913 (N_5913,N_5018,N_5229);
or U5914 (N_5914,N_5136,N_5444);
or U5915 (N_5915,N_5432,N_5115);
or U5916 (N_5916,N_5466,N_5190);
nor U5917 (N_5917,N_5320,N_5213);
nand U5918 (N_5918,N_5255,N_5070);
nor U5919 (N_5919,N_5467,N_5269);
or U5920 (N_5920,N_5363,N_5423);
xnor U5921 (N_5921,N_5434,N_5343);
or U5922 (N_5922,N_5184,N_5227);
nand U5923 (N_5923,N_5078,N_5274);
or U5924 (N_5924,N_5296,N_5120);
or U5925 (N_5925,N_5131,N_5212);
xor U5926 (N_5926,N_5284,N_5493);
and U5927 (N_5927,N_5426,N_5175);
or U5928 (N_5928,N_5198,N_5256);
and U5929 (N_5929,N_5281,N_5022);
nand U5930 (N_5930,N_5105,N_5123);
or U5931 (N_5931,N_5273,N_5064);
or U5932 (N_5932,N_5167,N_5363);
or U5933 (N_5933,N_5171,N_5339);
and U5934 (N_5934,N_5172,N_5085);
and U5935 (N_5935,N_5441,N_5258);
or U5936 (N_5936,N_5063,N_5436);
or U5937 (N_5937,N_5068,N_5166);
xor U5938 (N_5938,N_5439,N_5083);
xnor U5939 (N_5939,N_5059,N_5153);
nor U5940 (N_5940,N_5079,N_5083);
xor U5941 (N_5941,N_5454,N_5311);
nand U5942 (N_5942,N_5386,N_5226);
xor U5943 (N_5943,N_5059,N_5297);
nand U5944 (N_5944,N_5192,N_5112);
or U5945 (N_5945,N_5430,N_5190);
nor U5946 (N_5946,N_5036,N_5030);
xor U5947 (N_5947,N_5023,N_5279);
nand U5948 (N_5948,N_5334,N_5110);
xnor U5949 (N_5949,N_5025,N_5141);
and U5950 (N_5950,N_5239,N_5451);
and U5951 (N_5951,N_5284,N_5288);
or U5952 (N_5952,N_5372,N_5082);
or U5953 (N_5953,N_5246,N_5354);
nor U5954 (N_5954,N_5029,N_5339);
and U5955 (N_5955,N_5044,N_5340);
or U5956 (N_5956,N_5027,N_5245);
nor U5957 (N_5957,N_5062,N_5192);
nor U5958 (N_5958,N_5032,N_5068);
xnor U5959 (N_5959,N_5217,N_5159);
xnor U5960 (N_5960,N_5094,N_5167);
xnor U5961 (N_5961,N_5424,N_5088);
and U5962 (N_5962,N_5261,N_5206);
nor U5963 (N_5963,N_5434,N_5368);
nand U5964 (N_5964,N_5043,N_5325);
xor U5965 (N_5965,N_5333,N_5189);
xor U5966 (N_5966,N_5391,N_5272);
and U5967 (N_5967,N_5076,N_5111);
nor U5968 (N_5968,N_5474,N_5162);
and U5969 (N_5969,N_5128,N_5231);
and U5970 (N_5970,N_5285,N_5458);
or U5971 (N_5971,N_5226,N_5467);
xor U5972 (N_5972,N_5277,N_5053);
xor U5973 (N_5973,N_5086,N_5050);
nor U5974 (N_5974,N_5456,N_5453);
nand U5975 (N_5975,N_5285,N_5372);
nand U5976 (N_5976,N_5084,N_5155);
and U5977 (N_5977,N_5047,N_5486);
or U5978 (N_5978,N_5263,N_5178);
nand U5979 (N_5979,N_5018,N_5240);
xor U5980 (N_5980,N_5055,N_5030);
xnor U5981 (N_5981,N_5277,N_5182);
and U5982 (N_5982,N_5177,N_5488);
xnor U5983 (N_5983,N_5106,N_5331);
nor U5984 (N_5984,N_5253,N_5309);
xnor U5985 (N_5985,N_5056,N_5231);
xnor U5986 (N_5986,N_5096,N_5211);
xor U5987 (N_5987,N_5363,N_5370);
xnor U5988 (N_5988,N_5296,N_5126);
xor U5989 (N_5989,N_5054,N_5021);
or U5990 (N_5990,N_5464,N_5423);
or U5991 (N_5991,N_5373,N_5472);
nand U5992 (N_5992,N_5039,N_5416);
and U5993 (N_5993,N_5143,N_5264);
and U5994 (N_5994,N_5167,N_5354);
nor U5995 (N_5995,N_5372,N_5390);
nand U5996 (N_5996,N_5371,N_5235);
nor U5997 (N_5997,N_5317,N_5292);
and U5998 (N_5998,N_5024,N_5276);
xnor U5999 (N_5999,N_5328,N_5327);
and U6000 (N_6000,N_5611,N_5849);
xnor U6001 (N_6001,N_5600,N_5883);
or U6002 (N_6002,N_5579,N_5652);
nor U6003 (N_6003,N_5898,N_5506);
xnor U6004 (N_6004,N_5881,N_5953);
xnor U6005 (N_6005,N_5892,N_5871);
and U6006 (N_6006,N_5662,N_5752);
nand U6007 (N_6007,N_5640,N_5590);
nor U6008 (N_6008,N_5516,N_5601);
nor U6009 (N_6009,N_5531,N_5974);
or U6010 (N_6010,N_5749,N_5700);
xnor U6011 (N_6011,N_5818,N_5938);
and U6012 (N_6012,N_5677,N_5573);
xnor U6013 (N_6013,N_5803,N_5594);
or U6014 (N_6014,N_5889,N_5696);
xor U6015 (N_6015,N_5934,N_5688);
xnor U6016 (N_6016,N_5575,N_5914);
and U6017 (N_6017,N_5857,N_5988);
and U6018 (N_6018,N_5853,N_5915);
xnor U6019 (N_6019,N_5679,N_5557);
nor U6020 (N_6020,N_5970,N_5599);
nor U6021 (N_6021,N_5949,N_5880);
nor U6022 (N_6022,N_5561,N_5709);
nor U6023 (N_6023,N_5870,N_5607);
or U6024 (N_6024,N_5543,N_5900);
or U6025 (N_6025,N_5577,N_5882);
and U6026 (N_6026,N_5859,N_5981);
and U6027 (N_6027,N_5998,N_5759);
nand U6028 (N_6028,N_5789,N_5913);
nor U6029 (N_6029,N_5642,N_5636);
nor U6030 (N_6030,N_5546,N_5643);
or U6031 (N_6031,N_5769,N_5608);
nor U6032 (N_6032,N_5549,N_5862);
xnor U6033 (N_6033,N_5893,N_5620);
xor U6034 (N_6034,N_5872,N_5899);
nand U6035 (N_6035,N_5514,N_5568);
nand U6036 (N_6036,N_5727,N_5523);
xnor U6037 (N_6037,N_5824,N_5508);
nand U6038 (N_6038,N_5537,N_5861);
xnor U6039 (N_6039,N_5796,N_5804);
nand U6040 (N_6040,N_5694,N_5723);
and U6041 (N_6041,N_5515,N_5618);
or U6042 (N_6042,N_5919,N_5774);
xnor U6043 (N_6043,N_5983,N_5864);
nor U6044 (N_6044,N_5526,N_5858);
xnor U6045 (N_6045,N_5683,N_5605);
and U6046 (N_6046,N_5702,N_5512);
nand U6047 (N_6047,N_5627,N_5631);
or U6048 (N_6048,N_5954,N_5732);
and U6049 (N_6049,N_5786,N_5558);
and U6050 (N_6050,N_5659,N_5879);
xor U6051 (N_6051,N_5588,N_5750);
xnor U6052 (N_6052,N_5517,N_5544);
xor U6053 (N_6053,N_5868,N_5814);
nand U6054 (N_6054,N_5639,N_5664);
xor U6055 (N_6055,N_5707,N_5958);
nor U6056 (N_6056,N_5741,N_5572);
and U6057 (N_6057,N_5907,N_5584);
and U6058 (N_6058,N_5684,N_5687);
and U6059 (N_6059,N_5667,N_5541);
nand U6060 (N_6060,N_5668,N_5658);
nor U6061 (N_6061,N_5978,N_5610);
xnor U6062 (N_6062,N_5591,N_5821);
nand U6063 (N_6063,N_5901,N_5597);
xnor U6064 (N_6064,N_5629,N_5613);
or U6065 (N_6065,N_5780,N_5830);
or U6066 (N_6066,N_5634,N_5772);
or U6067 (N_6067,N_5909,N_5563);
nor U6068 (N_6068,N_5875,N_5979);
nand U6069 (N_6069,N_5962,N_5873);
xor U6070 (N_6070,N_5690,N_5929);
xor U6071 (N_6071,N_5765,N_5648);
or U6072 (N_6072,N_5673,N_5784);
nor U6073 (N_6073,N_5950,N_5565);
nor U6074 (N_6074,N_5733,N_5856);
xor U6075 (N_6075,N_5994,N_5518);
or U6076 (N_6076,N_5767,N_5834);
or U6077 (N_6077,N_5805,N_5795);
or U6078 (N_6078,N_5947,N_5832);
nand U6079 (N_6079,N_5647,N_5746);
nor U6080 (N_6080,N_5972,N_5850);
nand U6081 (N_6081,N_5806,N_5595);
nor U6082 (N_6082,N_5867,N_5912);
and U6083 (N_6083,N_5852,N_5781);
nor U6084 (N_6084,N_5559,N_5501);
xnor U6085 (N_6085,N_5722,N_5606);
or U6086 (N_6086,N_5828,N_5720);
and U6087 (N_6087,N_5910,N_5930);
or U6088 (N_6088,N_5682,N_5848);
nand U6089 (N_6089,N_5725,N_5744);
or U6090 (N_6090,N_5843,N_5614);
nor U6091 (N_6091,N_5829,N_5997);
nor U6092 (N_6092,N_5977,N_5616);
or U6093 (N_6093,N_5718,N_5985);
nor U6094 (N_6094,N_5555,N_5582);
xnor U6095 (N_6095,N_5739,N_5793);
nand U6096 (N_6096,N_5822,N_5507);
and U6097 (N_6097,N_5908,N_5646);
and U6098 (N_6098,N_5788,N_5635);
xnor U6099 (N_6099,N_5760,N_5987);
nand U6100 (N_6100,N_5996,N_5952);
and U6101 (N_6101,N_5633,N_5538);
xnor U6102 (N_6102,N_5532,N_5866);
and U6103 (N_6103,N_5704,N_5812);
or U6104 (N_6104,N_5891,N_5603);
xor U6105 (N_6105,N_5976,N_5534);
nand U6106 (N_6106,N_5992,N_5956);
nor U6107 (N_6107,N_5705,N_5895);
nor U6108 (N_6108,N_5671,N_5835);
nor U6109 (N_6109,N_5808,N_5757);
or U6110 (N_6110,N_5982,N_5612);
nand U6111 (N_6111,N_5773,N_5714);
nor U6112 (N_6112,N_5622,N_5721);
nand U6113 (N_6113,N_5753,N_5927);
xnor U6114 (N_6114,N_5528,N_5693);
xnor U6115 (N_6115,N_5586,N_5995);
and U6116 (N_6116,N_5547,N_5840);
nor U6117 (N_6117,N_5548,N_5504);
and U6118 (N_6118,N_5916,N_5877);
xnor U6119 (N_6119,N_5969,N_5530);
or U6120 (N_6120,N_5713,N_5511);
nand U6121 (N_6121,N_5576,N_5837);
xnor U6122 (N_6122,N_5869,N_5681);
xor U6123 (N_6123,N_5503,N_5894);
and U6124 (N_6124,N_5560,N_5729);
and U6125 (N_6125,N_5585,N_5617);
nor U6126 (N_6126,N_5924,N_5776);
xor U6127 (N_6127,N_5500,N_5800);
nand U6128 (N_6128,N_5959,N_5931);
and U6129 (N_6129,N_5593,N_5797);
xnor U6130 (N_6130,N_5819,N_5698);
or U6131 (N_6131,N_5738,N_5663);
and U6132 (N_6132,N_5779,N_5933);
xor U6133 (N_6133,N_5918,N_5556);
and U6134 (N_6134,N_5654,N_5535);
or U6135 (N_6135,N_5728,N_5717);
or U6136 (N_6136,N_5851,N_5615);
nor U6137 (N_6137,N_5502,N_5903);
xnor U6138 (N_6138,N_5937,N_5825);
or U6139 (N_6139,N_5656,N_5533);
nand U6140 (N_6140,N_5975,N_5758);
or U6141 (N_6141,N_5621,N_5905);
nand U6142 (N_6142,N_5580,N_5798);
nor U6143 (N_6143,N_5708,N_5574);
nand U6144 (N_6144,N_5651,N_5672);
or U6145 (N_6145,N_5945,N_5742);
nand U6146 (N_6146,N_5645,N_5860);
and U6147 (N_6147,N_5520,N_5630);
or U6148 (N_6148,N_5971,N_5598);
nand U6149 (N_6149,N_5686,N_5942);
or U6150 (N_6150,N_5680,N_5666);
xor U6151 (N_6151,N_5587,N_5802);
nor U6152 (N_6152,N_5801,N_5878);
or U6153 (N_6153,N_5581,N_5820);
nor U6154 (N_6154,N_5941,N_5920);
nor U6155 (N_6155,N_5973,N_5695);
xor U6156 (N_6156,N_5715,N_5966);
xor U6157 (N_6157,N_5712,N_5562);
xnor U6158 (N_6158,N_5963,N_5886);
xor U6159 (N_6159,N_5521,N_5884);
nand U6160 (N_6160,N_5887,N_5510);
xnor U6161 (N_6161,N_5925,N_5566);
nand U6162 (N_6162,N_5785,N_5810);
or U6163 (N_6163,N_5578,N_5763);
or U6164 (N_6164,N_5644,N_5756);
nand U6165 (N_6165,N_5754,N_5792);
nor U6166 (N_6166,N_5813,N_5787);
or U6167 (N_6167,N_5554,N_5771);
nand U6168 (N_6168,N_5782,N_5811);
xnor U6169 (N_6169,N_5967,N_5626);
nor U6170 (N_6170,N_5940,N_5906);
and U6171 (N_6171,N_5838,N_5833);
nor U6172 (N_6172,N_5650,N_5553);
xnor U6173 (N_6173,N_5638,N_5527);
nand U6174 (N_6174,N_5604,N_5839);
xnor U6175 (N_6175,N_5653,N_5748);
nand U6176 (N_6176,N_5678,N_5689);
or U6177 (N_6177,N_5740,N_5734);
nand U6178 (N_6178,N_5799,N_5550);
nand U6179 (N_6179,N_5766,N_5670);
xnor U6180 (N_6180,N_5961,N_5619);
xor U6181 (N_6181,N_5632,N_5542);
xor U6182 (N_6182,N_5509,N_5790);
and U6183 (N_6183,N_5571,N_5536);
and U6184 (N_6184,N_5965,N_5567);
nand U6185 (N_6185,N_5637,N_5675);
and U6186 (N_6186,N_5710,N_5552);
and U6187 (N_6187,N_5697,N_5984);
nor U6188 (N_6188,N_5676,N_5836);
xor U6189 (N_6189,N_5762,N_5596);
and U6190 (N_6190,N_5991,N_5743);
xnor U6191 (N_6191,N_5964,N_5570);
nand U6192 (N_6192,N_5874,N_5778);
or U6193 (N_6193,N_5706,N_5816);
and U6194 (N_6194,N_5624,N_5524);
and U6195 (N_6195,N_5939,N_5569);
or U6196 (N_6196,N_5794,N_5854);
and U6197 (N_6197,N_5589,N_5649);
nand U6198 (N_6198,N_5817,N_5711);
nand U6199 (N_6199,N_5735,N_5846);
or U6200 (N_6200,N_5768,N_5863);
nand U6201 (N_6201,N_5522,N_5948);
or U6202 (N_6202,N_5660,N_5911);
nand U6203 (N_6203,N_5827,N_5525);
and U6204 (N_6204,N_5989,N_5809);
nand U6205 (N_6205,N_5885,N_5922);
nand U6206 (N_6206,N_5655,N_5691);
and U6207 (N_6207,N_5807,N_5703);
or U6208 (N_6208,N_5923,N_5826);
or U6209 (N_6209,N_5986,N_5674);
nor U6210 (N_6210,N_5731,N_5896);
nor U6211 (N_6211,N_5564,N_5770);
nand U6212 (N_6212,N_5505,N_5665);
nand U6213 (N_6213,N_5890,N_5946);
nand U6214 (N_6214,N_5539,N_5628);
or U6215 (N_6215,N_5951,N_5730);
nor U6216 (N_6216,N_5990,N_5726);
nand U6217 (N_6217,N_5791,N_5609);
or U6218 (N_6218,N_5699,N_5719);
xor U6219 (N_6219,N_5751,N_5980);
xnor U6220 (N_6220,N_5831,N_5716);
and U6221 (N_6221,N_5926,N_5623);
nand U6222 (N_6222,N_5692,N_5955);
or U6223 (N_6223,N_5935,N_5844);
xor U6224 (N_6224,N_5888,N_5815);
nand U6225 (N_6225,N_5845,N_5764);
or U6226 (N_6226,N_5902,N_5755);
nor U6227 (N_6227,N_5960,N_5936);
and U6228 (N_6228,N_5747,N_5545);
or U6229 (N_6229,N_5841,N_5999);
nor U6230 (N_6230,N_5724,N_5529);
nor U6231 (N_6231,N_5661,N_5540);
and U6232 (N_6232,N_5775,N_5761);
nand U6233 (N_6233,N_5783,N_5876);
nand U6234 (N_6234,N_5897,N_5625);
or U6235 (N_6235,N_5669,N_5745);
or U6236 (N_6236,N_5736,N_5917);
nor U6237 (N_6237,N_5685,N_5921);
or U6238 (N_6238,N_5602,N_5993);
and U6239 (N_6239,N_5737,N_5865);
nand U6240 (N_6240,N_5842,N_5583);
nand U6241 (N_6241,N_5928,N_5551);
xnor U6242 (N_6242,N_5519,N_5904);
nand U6243 (N_6243,N_5641,N_5657);
and U6244 (N_6244,N_5957,N_5701);
nand U6245 (N_6245,N_5855,N_5823);
or U6246 (N_6246,N_5932,N_5847);
nand U6247 (N_6247,N_5513,N_5943);
xnor U6248 (N_6248,N_5944,N_5968);
and U6249 (N_6249,N_5592,N_5777);
or U6250 (N_6250,N_5745,N_5822);
nand U6251 (N_6251,N_5748,N_5686);
or U6252 (N_6252,N_5837,N_5651);
xor U6253 (N_6253,N_5584,N_5755);
or U6254 (N_6254,N_5721,N_5895);
nand U6255 (N_6255,N_5975,N_5897);
and U6256 (N_6256,N_5923,N_5858);
nand U6257 (N_6257,N_5963,N_5859);
or U6258 (N_6258,N_5903,N_5928);
or U6259 (N_6259,N_5643,N_5825);
xnor U6260 (N_6260,N_5796,N_5961);
nor U6261 (N_6261,N_5925,N_5678);
xor U6262 (N_6262,N_5705,N_5860);
or U6263 (N_6263,N_5826,N_5740);
and U6264 (N_6264,N_5598,N_5682);
nor U6265 (N_6265,N_5647,N_5834);
or U6266 (N_6266,N_5972,N_5539);
and U6267 (N_6267,N_5772,N_5673);
and U6268 (N_6268,N_5779,N_5586);
and U6269 (N_6269,N_5632,N_5785);
or U6270 (N_6270,N_5527,N_5891);
nor U6271 (N_6271,N_5812,N_5593);
and U6272 (N_6272,N_5677,N_5885);
and U6273 (N_6273,N_5951,N_5676);
or U6274 (N_6274,N_5768,N_5742);
or U6275 (N_6275,N_5803,N_5853);
and U6276 (N_6276,N_5663,N_5980);
and U6277 (N_6277,N_5890,N_5500);
xor U6278 (N_6278,N_5927,N_5972);
nor U6279 (N_6279,N_5711,N_5825);
or U6280 (N_6280,N_5550,N_5556);
nand U6281 (N_6281,N_5782,N_5732);
xor U6282 (N_6282,N_5722,N_5892);
or U6283 (N_6283,N_5972,N_5512);
and U6284 (N_6284,N_5647,N_5580);
nand U6285 (N_6285,N_5551,N_5797);
or U6286 (N_6286,N_5659,N_5538);
nand U6287 (N_6287,N_5771,N_5930);
nand U6288 (N_6288,N_5955,N_5647);
xor U6289 (N_6289,N_5755,N_5834);
and U6290 (N_6290,N_5617,N_5982);
or U6291 (N_6291,N_5870,N_5627);
nand U6292 (N_6292,N_5501,N_5578);
and U6293 (N_6293,N_5799,N_5757);
or U6294 (N_6294,N_5764,N_5554);
or U6295 (N_6295,N_5672,N_5590);
or U6296 (N_6296,N_5599,N_5614);
and U6297 (N_6297,N_5896,N_5534);
xor U6298 (N_6298,N_5892,N_5675);
nor U6299 (N_6299,N_5713,N_5599);
xnor U6300 (N_6300,N_5529,N_5709);
nand U6301 (N_6301,N_5533,N_5558);
xnor U6302 (N_6302,N_5653,N_5710);
nand U6303 (N_6303,N_5596,N_5758);
or U6304 (N_6304,N_5533,N_5508);
nor U6305 (N_6305,N_5846,N_5740);
xor U6306 (N_6306,N_5551,N_5982);
and U6307 (N_6307,N_5784,N_5573);
xor U6308 (N_6308,N_5665,N_5761);
and U6309 (N_6309,N_5634,N_5985);
and U6310 (N_6310,N_5963,N_5779);
nor U6311 (N_6311,N_5960,N_5540);
and U6312 (N_6312,N_5879,N_5988);
and U6313 (N_6313,N_5981,N_5741);
or U6314 (N_6314,N_5533,N_5565);
xnor U6315 (N_6315,N_5860,N_5842);
or U6316 (N_6316,N_5885,N_5963);
nor U6317 (N_6317,N_5980,N_5822);
xnor U6318 (N_6318,N_5815,N_5640);
or U6319 (N_6319,N_5735,N_5796);
xnor U6320 (N_6320,N_5665,N_5570);
and U6321 (N_6321,N_5661,N_5984);
and U6322 (N_6322,N_5751,N_5715);
nand U6323 (N_6323,N_5996,N_5857);
and U6324 (N_6324,N_5985,N_5990);
nor U6325 (N_6325,N_5553,N_5651);
nor U6326 (N_6326,N_5807,N_5578);
nor U6327 (N_6327,N_5546,N_5670);
nor U6328 (N_6328,N_5953,N_5575);
xor U6329 (N_6329,N_5858,N_5956);
or U6330 (N_6330,N_5639,N_5755);
and U6331 (N_6331,N_5534,N_5970);
or U6332 (N_6332,N_5966,N_5768);
and U6333 (N_6333,N_5562,N_5663);
nor U6334 (N_6334,N_5722,N_5750);
or U6335 (N_6335,N_5581,N_5885);
or U6336 (N_6336,N_5636,N_5565);
or U6337 (N_6337,N_5530,N_5558);
and U6338 (N_6338,N_5962,N_5572);
nor U6339 (N_6339,N_5801,N_5847);
or U6340 (N_6340,N_5643,N_5563);
nor U6341 (N_6341,N_5966,N_5825);
or U6342 (N_6342,N_5823,N_5511);
or U6343 (N_6343,N_5877,N_5613);
and U6344 (N_6344,N_5500,N_5834);
nand U6345 (N_6345,N_5950,N_5632);
nor U6346 (N_6346,N_5584,N_5883);
nor U6347 (N_6347,N_5804,N_5594);
nor U6348 (N_6348,N_5606,N_5789);
xor U6349 (N_6349,N_5813,N_5532);
nor U6350 (N_6350,N_5514,N_5706);
xor U6351 (N_6351,N_5979,N_5909);
nand U6352 (N_6352,N_5656,N_5983);
xnor U6353 (N_6353,N_5909,N_5605);
nand U6354 (N_6354,N_5717,N_5570);
nor U6355 (N_6355,N_5673,N_5904);
nor U6356 (N_6356,N_5631,N_5781);
nor U6357 (N_6357,N_5592,N_5712);
nor U6358 (N_6358,N_5592,N_5804);
xnor U6359 (N_6359,N_5998,N_5549);
or U6360 (N_6360,N_5731,N_5592);
and U6361 (N_6361,N_5550,N_5690);
nand U6362 (N_6362,N_5900,N_5628);
xnor U6363 (N_6363,N_5529,N_5755);
nor U6364 (N_6364,N_5727,N_5903);
xor U6365 (N_6365,N_5510,N_5582);
or U6366 (N_6366,N_5742,N_5532);
and U6367 (N_6367,N_5664,N_5732);
and U6368 (N_6368,N_5833,N_5579);
xor U6369 (N_6369,N_5949,N_5987);
nor U6370 (N_6370,N_5514,N_5814);
nor U6371 (N_6371,N_5929,N_5815);
nand U6372 (N_6372,N_5774,N_5618);
nand U6373 (N_6373,N_5621,N_5973);
nand U6374 (N_6374,N_5786,N_5546);
and U6375 (N_6375,N_5614,N_5716);
nand U6376 (N_6376,N_5962,N_5570);
xor U6377 (N_6377,N_5682,N_5697);
nand U6378 (N_6378,N_5537,N_5638);
nand U6379 (N_6379,N_5816,N_5835);
and U6380 (N_6380,N_5688,N_5632);
and U6381 (N_6381,N_5777,N_5773);
nand U6382 (N_6382,N_5590,N_5921);
xor U6383 (N_6383,N_5636,N_5999);
xnor U6384 (N_6384,N_5967,N_5534);
nand U6385 (N_6385,N_5801,N_5852);
xor U6386 (N_6386,N_5989,N_5630);
nor U6387 (N_6387,N_5774,N_5544);
nand U6388 (N_6388,N_5800,N_5738);
xnor U6389 (N_6389,N_5755,N_5730);
xor U6390 (N_6390,N_5990,N_5997);
and U6391 (N_6391,N_5752,N_5980);
and U6392 (N_6392,N_5580,N_5848);
nand U6393 (N_6393,N_5673,N_5575);
xor U6394 (N_6394,N_5795,N_5910);
xor U6395 (N_6395,N_5714,N_5513);
and U6396 (N_6396,N_5670,N_5760);
and U6397 (N_6397,N_5774,N_5610);
nand U6398 (N_6398,N_5604,N_5631);
and U6399 (N_6399,N_5691,N_5635);
and U6400 (N_6400,N_5809,N_5583);
xor U6401 (N_6401,N_5663,N_5525);
nand U6402 (N_6402,N_5829,N_5931);
and U6403 (N_6403,N_5946,N_5652);
nand U6404 (N_6404,N_5950,N_5845);
and U6405 (N_6405,N_5954,N_5887);
nand U6406 (N_6406,N_5966,N_5604);
xor U6407 (N_6407,N_5763,N_5963);
and U6408 (N_6408,N_5733,N_5832);
nor U6409 (N_6409,N_5650,N_5584);
nor U6410 (N_6410,N_5563,N_5522);
nand U6411 (N_6411,N_5595,N_5723);
and U6412 (N_6412,N_5548,N_5590);
and U6413 (N_6413,N_5703,N_5677);
nand U6414 (N_6414,N_5697,N_5861);
nand U6415 (N_6415,N_5934,N_5747);
xor U6416 (N_6416,N_5651,N_5986);
nand U6417 (N_6417,N_5784,N_5729);
and U6418 (N_6418,N_5858,N_5579);
or U6419 (N_6419,N_5744,N_5643);
or U6420 (N_6420,N_5518,N_5512);
nand U6421 (N_6421,N_5741,N_5556);
nand U6422 (N_6422,N_5511,N_5694);
xor U6423 (N_6423,N_5770,N_5962);
nand U6424 (N_6424,N_5642,N_5518);
xor U6425 (N_6425,N_5808,N_5622);
nor U6426 (N_6426,N_5962,N_5622);
nor U6427 (N_6427,N_5914,N_5681);
nand U6428 (N_6428,N_5932,N_5999);
or U6429 (N_6429,N_5963,N_5797);
or U6430 (N_6430,N_5615,N_5708);
xnor U6431 (N_6431,N_5772,N_5794);
nand U6432 (N_6432,N_5629,N_5636);
nor U6433 (N_6433,N_5673,N_5705);
xor U6434 (N_6434,N_5962,N_5601);
and U6435 (N_6435,N_5909,N_5805);
xnor U6436 (N_6436,N_5561,N_5808);
nand U6437 (N_6437,N_5892,N_5947);
xor U6438 (N_6438,N_5928,N_5968);
or U6439 (N_6439,N_5664,N_5803);
and U6440 (N_6440,N_5688,N_5925);
nor U6441 (N_6441,N_5971,N_5562);
xor U6442 (N_6442,N_5556,N_5750);
nand U6443 (N_6443,N_5869,N_5883);
nand U6444 (N_6444,N_5684,N_5665);
or U6445 (N_6445,N_5951,N_5564);
nand U6446 (N_6446,N_5744,N_5973);
and U6447 (N_6447,N_5972,N_5953);
and U6448 (N_6448,N_5806,N_5530);
xnor U6449 (N_6449,N_5827,N_5869);
nand U6450 (N_6450,N_5925,N_5706);
or U6451 (N_6451,N_5923,N_5715);
xor U6452 (N_6452,N_5786,N_5870);
and U6453 (N_6453,N_5857,N_5571);
or U6454 (N_6454,N_5604,N_5987);
or U6455 (N_6455,N_5887,N_5894);
and U6456 (N_6456,N_5717,N_5580);
or U6457 (N_6457,N_5867,N_5900);
nor U6458 (N_6458,N_5734,N_5773);
nor U6459 (N_6459,N_5553,N_5958);
nand U6460 (N_6460,N_5548,N_5597);
and U6461 (N_6461,N_5719,N_5857);
xnor U6462 (N_6462,N_5743,N_5973);
and U6463 (N_6463,N_5912,N_5839);
nand U6464 (N_6464,N_5529,N_5741);
nor U6465 (N_6465,N_5587,N_5869);
nor U6466 (N_6466,N_5661,N_5709);
nor U6467 (N_6467,N_5575,N_5569);
or U6468 (N_6468,N_5607,N_5587);
or U6469 (N_6469,N_5643,N_5730);
xor U6470 (N_6470,N_5836,N_5812);
nor U6471 (N_6471,N_5815,N_5561);
nand U6472 (N_6472,N_5564,N_5833);
and U6473 (N_6473,N_5531,N_5652);
nor U6474 (N_6474,N_5737,N_5507);
and U6475 (N_6475,N_5529,N_5892);
or U6476 (N_6476,N_5789,N_5636);
or U6477 (N_6477,N_5791,N_5849);
nand U6478 (N_6478,N_5890,N_5610);
and U6479 (N_6479,N_5582,N_5953);
and U6480 (N_6480,N_5957,N_5719);
nor U6481 (N_6481,N_5732,N_5770);
nand U6482 (N_6482,N_5611,N_5801);
or U6483 (N_6483,N_5667,N_5615);
nor U6484 (N_6484,N_5907,N_5905);
nor U6485 (N_6485,N_5540,N_5814);
nand U6486 (N_6486,N_5831,N_5718);
nand U6487 (N_6487,N_5607,N_5977);
nor U6488 (N_6488,N_5943,N_5538);
or U6489 (N_6489,N_5815,N_5634);
nand U6490 (N_6490,N_5689,N_5644);
or U6491 (N_6491,N_5812,N_5822);
and U6492 (N_6492,N_5573,N_5791);
xnor U6493 (N_6493,N_5813,N_5911);
or U6494 (N_6494,N_5755,N_5516);
xnor U6495 (N_6495,N_5922,N_5527);
or U6496 (N_6496,N_5797,N_5751);
nor U6497 (N_6497,N_5722,N_5529);
or U6498 (N_6498,N_5795,N_5632);
or U6499 (N_6499,N_5911,N_5805);
nor U6500 (N_6500,N_6240,N_6292);
nand U6501 (N_6501,N_6259,N_6496);
and U6502 (N_6502,N_6333,N_6485);
nor U6503 (N_6503,N_6379,N_6410);
nand U6504 (N_6504,N_6144,N_6372);
xor U6505 (N_6505,N_6457,N_6251);
and U6506 (N_6506,N_6417,N_6010);
nand U6507 (N_6507,N_6081,N_6281);
xor U6508 (N_6508,N_6291,N_6235);
and U6509 (N_6509,N_6203,N_6201);
nor U6510 (N_6510,N_6392,N_6091);
and U6511 (N_6511,N_6335,N_6444);
xor U6512 (N_6512,N_6268,N_6214);
or U6513 (N_6513,N_6207,N_6229);
nor U6514 (N_6514,N_6471,N_6123);
or U6515 (N_6515,N_6362,N_6196);
and U6516 (N_6516,N_6257,N_6127);
nor U6517 (N_6517,N_6355,N_6059);
or U6518 (N_6518,N_6013,N_6323);
or U6519 (N_6519,N_6473,N_6418);
nor U6520 (N_6520,N_6193,N_6051);
nor U6521 (N_6521,N_6409,N_6087);
or U6522 (N_6522,N_6187,N_6337);
nand U6523 (N_6523,N_6408,N_6384);
and U6524 (N_6524,N_6395,N_6086);
and U6525 (N_6525,N_6137,N_6097);
or U6526 (N_6526,N_6480,N_6038);
nor U6527 (N_6527,N_6426,N_6027);
nor U6528 (N_6528,N_6244,N_6232);
or U6529 (N_6529,N_6407,N_6312);
and U6530 (N_6530,N_6233,N_6237);
xor U6531 (N_6531,N_6338,N_6146);
and U6532 (N_6532,N_6172,N_6357);
and U6533 (N_6533,N_6219,N_6239);
nand U6534 (N_6534,N_6495,N_6269);
nand U6535 (N_6535,N_6136,N_6446);
nor U6536 (N_6536,N_6393,N_6497);
xor U6537 (N_6537,N_6045,N_6103);
nor U6538 (N_6538,N_6162,N_6238);
nor U6539 (N_6539,N_6411,N_6065);
nor U6540 (N_6540,N_6467,N_6126);
and U6541 (N_6541,N_6298,N_6472);
nor U6542 (N_6542,N_6309,N_6275);
nand U6543 (N_6543,N_6068,N_6332);
and U6544 (N_6544,N_6370,N_6024);
or U6545 (N_6545,N_6018,N_6115);
or U6546 (N_6546,N_6433,N_6063);
and U6547 (N_6547,N_6425,N_6113);
nand U6548 (N_6548,N_6491,N_6208);
nand U6549 (N_6549,N_6255,N_6040);
nand U6550 (N_6550,N_6330,N_6397);
or U6551 (N_6551,N_6154,N_6061);
xnor U6552 (N_6552,N_6297,N_6276);
or U6553 (N_6553,N_6007,N_6004);
nor U6554 (N_6554,N_6353,N_6328);
xor U6555 (N_6555,N_6438,N_6270);
nor U6556 (N_6556,N_6058,N_6174);
nor U6557 (N_6557,N_6468,N_6035);
nand U6558 (N_6558,N_6033,N_6373);
nor U6559 (N_6559,N_6404,N_6195);
nand U6560 (N_6560,N_6169,N_6374);
nor U6561 (N_6561,N_6401,N_6340);
nand U6562 (N_6562,N_6181,N_6345);
nand U6563 (N_6563,N_6339,N_6290);
nand U6564 (N_6564,N_6124,N_6441);
nand U6565 (N_6565,N_6188,N_6028);
or U6566 (N_6566,N_6265,N_6145);
nor U6567 (N_6567,N_6118,N_6354);
and U6568 (N_6568,N_6047,N_6288);
nor U6569 (N_6569,N_6325,N_6246);
and U6570 (N_6570,N_6304,N_6073);
xnor U6571 (N_6571,N_6151,N_6221);
or U6572 (N_6572,N_6066,N_6498);
or U6573 (N_6573,N_6415,N_6076);
nand U6574 (N_6574,N_6250,N_6217);
or U6575 (N_6575,N_6069,N_6343);
and U6576 (N_6576,N_6450,N_6184);
xnor U6577 (N_6577,N_6488,N_6200);
or U6578 (N_6578,N_6106,N_6100);
and U6579 (N_6579,N_6133,N_6416);
xnor U6580 (N_6580,N_6029,N_6053);
or U6581 (N_6581,N_6331,N_6280);
nor U6582 (N_6582,N_6400,N_6216);
nand U6583 (N_6583,N_6037,N_6166);
xnor U6584 (N_6584,N_6279,N_6399);
nor U6585 (N_6585,N_6022,N_6483);
and U6586 (N_6586,N_6001,N_6088);
nor U6587 (N_6587,N_6342,N_6459);
nand U6588 (N_6588,N_6435,N_6191);
xnor U6589 (N_6589,N_6313,N_6341);
or U6590 (N_6590,N_6116,N_6322);
and U6591 (N_6591,N_6434,N_6025);
and U6592 (N_6592,N_6306,N_6356);
nand U6593 (N_6593,N_6095,N_6159);
or U6594 (N_6594,N_6228,N_6283);
nand U6595 (N_6595,N_6347,N_6023);
and U6596 (N_6596,N_6183,N_6352);
and U6597 (N_6597,N_6026,N_6102);
and U6598 (N_6598,N_6132,N_6083);
nor U6599 (N_6599,N_6148,N_6175);
nand U6600 (N_6600,N_6487,N_6294);
xnor U6601 (N_6601,N_6107,N_6256);
and U6602 (N_6602,N_6179,N_6054);
nand U6603 (N_6603,N_6267,N_6271);
xnor U6604 (N_6604,N_6463,N_6430);
or U6605 (N_6605,N_6226,N_6344);
nand U6606 (N_6606,N_6316,N_6336);
nand U6607 (N_6607,N_6163,N_6277);
or U6608 (N_6608,N_6346,N_6402);
and U6609 (N_6609,N_6419,N_6462);
and U6610 (N_6610,N_6261,N_6015);
nor U6611 (N_6611,N_6371,N_6079);
nand U6612 (N_6612,N_6460,N_6011);
or U6613 (N_6613,N_6249,N_6470);
nand U6614 (N_6614,N_6348,N_6224);
or U6615 (N_6615,N_6469,N_6248);
nor U6616 (N_6616,N_6398,N_6465);
and U6617 (N_6617,N_6489,N_6376);
or U6618 (N_6618,N_6412,N_6153);
xnor U6619 (N_6619,N_6300,N_6085);
and U6620 (N_6620,N_6139,N_6197);
nand U6621 (N_6621,N_6484,N_6456);
or U6622 (N_6622,N_6305,N_6016);
and U6623 (N_6623,N_6315,N_6262);
xnor U6624 (N_6624,N_6284,N_6366);
and U6625 (N_6625,N_6098,N_6388);
nand U6626 (N_6626,N_6032,N_6464);
and U6627 (N_6627,N_6167,N_6055);
nand U6628 (N_6628,N_6420,N_6178);
nand U6629 (N_6629,N_6381,N_6064);
nor U6630 (N_6630,N_6090,N_6108);
and U6631 (N_6631,N_6390,N_6486);
and U6632 (N_6632,N_6365,N_6252);
nor U6633 (N_6633,N_6014,N_6020);
or U6634 (N_6634,N_6245,N_6436);
nor U6635 (N_6635,N_6364,N_6260);
nor U6636 (N_6636,N_6084,N_6258);
nor U6637 (N_6637,N_6049,N_6317);
or U6638 (N_6638,N_6242,N_6272);
nand U6639 (N_6639,N_6114,N_6128);
nand U6640 (N_6640,N_6363,N_6129);
or U6641 (N_6641,N_6101,N_6044);
nor U6642 (N_6642,N_6445,N_6158);
xnor U6643 (N_6643,N_6006,N_6386);
xor U6644 (N_6644,N_6152,N_6302);
nand U6645 (N_6645,N_6093,N_6194);
nand U6646 (N_6646,N_6130,N_6171);
nand U6647 (N_6647,N_6067,N_6458);
or U6648 (N_6648,N_6396,N_6442);
nand U6649 (N_6649,N_6319,N_6424);
nor U6650 (N_6650,N_6150,N_6367);
or U6651 (N_6651,N_6094,N_6358);
nor U6652 (N_6652,N_6359,N_6432);
nand U6653 (N_6653,N_6293,N_6180);
and U6654 (N_6654,N_6156,N_6451);
nand U6655 (N_6655,N_6176,N_6494);
and U6656 (N_6656,N_6287,N_6039);
nand U6657 (N_6657,N_6147,N_6324);
nor U6658 (N_6658,N_6211,N_6314);
or U6659 (N_6659,N_6429,N_6492);
nand U6660 (N_6660,N_6198,N_6320);
xor U6661 (N_6661,N_6382,N_6383);
and U6662 (N_6662,N_6213,N_6282);
nor U6663 (N_6663,N_6227,N_6142);
and U6664 (N_6664,N_6140,N_6482);
nor U6665 (N_6665,N_6380,N_6052);
nor U6666 (N_6666,N_6448,N_6121);
xor U6667 (N_6667,N_6307,N_6177);
nor U6668 (N_6668,N_6406,N_6056);
xor U6669 (N_6669,N_6263,N_6421);
or U6670 (N_6670,N_6273,N_6134);
xnor U6671 (N_6671,N_6161,N_6215);
nand U6672 (N_6672,N_6241,N_6182);
nor U6673 (N_6673,N_6440,N_6385);
nor U6674 (N_6674,N_6135,N_6391);
nor U6675 (N_6675,N_6225,N_6349);
or U6676 (N_6676,N_6499,N_6110);
or U6677 (N_6677,N_6449,N_6375);
nor U6678 (N_6678,N_6206,N_6034);
and U6679 (N_6679,N_6173,N_6286);
or U6680 (N_6680,N_6264,N_6138);
nand U6681 (N_6681,N_6096,N_6368);
nand U6682 (N_6682,N_6003,N_6143);
or U6683 (N_6683,N_6243,N_6443);
or U6684 (N_6684,N_6046,N_6082);
xnor U6685 (N_6685,N_6199,N_6413);
and U6686 (N_6686,N_6050,N_6476);
and U6687 (N_6687,N_6168,N_6311);
and U6688 (N_6688,N_6042,N_6080);
nand U6689 (N_6689,N_6490,N_6301);
nor U6690 (N_6690,N_6389,N_6204);
nand U6691 (N_6691,N_6310,N_6048);
nor U6692 (N_6692,N_6454,N_6155);
nand U6693 (N_6693,N_6165,N_6428);
xnor U6694 (N_6694,N_6189,N_6062);
nor U6695 (N_6695,N_6036,N_6474);
xor U6696 (N_6696,N_6361,N_6478);
or U6697 (N_6697,N_6414,N_6117);
or U6698 (N_6698,N_6439,N_6296);
xnor U6699 (N_6699,N_6218,N_6477);
and U6700 (N_6700,N_6236,N_6031);
or U6701 (N_6701,N_6461,N_6021);
nand U6702 (N_6702,N_6008,N_6074);
or U6703 (N_6703,N_6403,N_6274);
xor U6704 (N_6704,N_6017,N_6289);
xnor U6705 (N_6705,N_6351,N_6120);
and U6706 (N_6706,N_6423,N_6231);
nor U6707 (N_6707,N_6479,N_6223);
nor U6708 (N_6708,N_6019,N_6030);
or U6709 (N_6709,N_6157,N_6190);
xnor U6710 (N_6710,N_6170,N_6104);
nand U6711 (N_6711,N_6431,N_6009);
nor U6712 (N_6712,N_6334,N_6405);
xnor U6713 (N_6713,N_6422,N_6447);
xor U6714 (N_6714,N_6481,N_6078);
and U6715 (N_6715,N_6105,N_6125);
nor U6716 (N_6716,N_6075,N_6192);
or U6717 (N_6717,N_6360,N_6387);
and U6718 (N_6718,N_6253,N_6475);
nor U6719 (N_6719,N_6285,N_6210);
nand U6720 (N_6720,N_6077,N_6185);
and U6721 (N_6721,N_6466,N_6149);
xnor U6722 (N_6722,N_6160,N_6378);
xor U6723 (N_6723,N_6266,N_6205);
nor U6724 (N_6724,N_6072,N_6164);
nor U6725 (N_6725,N_6254,N_6099);
or U6726 (N_6726,N_6278,N_6112);
nand U6727 (N_6727,N_6186,N_6222);
xor U6728 (N_6728,N_6202,N_6122);
and U6729 (N_6729,N_6141,N_6303);
or U6730 (N_6730,N_6109,N_6212);
and U6731 (N_6731,N_6220,N_6057);
and U6732 (N_6732,N_6308,N_6394);
and U6733 (N_6733,N_6234,N_6005);
xor U6734 (N_6734,N_6012,N_6318);
nor U6735 (N_6735,N_6329,N_6452);
nand U6736 (N_6736,N_6350,N_6326);
and U6737 (N_6737,N_6230,N_6299);
or U6738 (N_6738,N_6493,N_6453);
xnor U6739 (N_6739,N_6002,N_6369);
xnor U6740 (N_6740,N_6377,N_6247);
nor U6741 (N_6741,N_6427,N_6209);
and U6742 (N_6742,N_6089,N_6071);
and U6743 (N_6743,N_6437,N_6000);
xnor U6744 (N_6744,N_6111,N_6070);
and U6745 (N_6745,N_6131,N_6041);
nor U6746 (N_6746,N_6295,N_6043);
nand U6747 (N_6747,N_6092,N_6119);
nand U6748 (N_6748,N_6321,N_6455);
nor U6749 (N_6749,N_6060,N_6327);
nand U6750 (N_6750,N_6217,N_6210);
nor U6751 (N_6751,N_6447,N_6365);
nand U6752 (N_6752,N_6160,N_6235);
xor U6753 (N_6753,N_6161,N_6276);
nor U6754 (N_6754,N_6332,N_6356);
and U6755 (N_6755,N_6089,N_6405);
or U6756 (N_6756,N_6338,N_6228);
xor U6757 (N_6757,N_6055,N_6262);
and U6758 (N_6758,N_6141,N_6129);
xnor U6759 (N_6759,N_6494,N_6126);
or U6760 (N_6760,N_6106,N_6090);
nor U6761 (N_6761,N_6101,N_6310);
nand U6762 (N_6762,N_6497,N_6082);
xor U6763 (N_6763,N_6035,N_6146);
xor U6764 (N_6764,N_6146,N_6173);
or U6765 (N_6765,N_6194,N_6429);
or U6766 (N_6766,N_6330,N_6365);
or U6767 (N_6767,N_6226,N_6127);
nand U6768 (N_6768,N_6492,N_6443);
nor U6769 (N_6769,N_6260,N_6330);
and U6770 (N_6770,N_6377,N_6065);
and U6771 (N_6771,N_6286,N_6029);
or U6772 (N_6772,N_6175,N_6312);
nor U6773 (N_6773,N_6066,N_6294);
nor U6774 (N_6774,N_6340,N_6474);
or U6775 (N_6775,N_6322,N_6292);
xnor U6776 (N_6776,N_6329,N_6080);
and U6777 (N_6777,N_6191,N_6160);
nor U6778 (N_6778,N_6237,N_6039);
xor U6779 (N_6779,N_6355,N_6367);
and U6780 (N_6780,N_6189,N_6095);
and U6781 (N_6781,N_6322,N_6165);
nand U6782 (N_6782,N_6240,N_6431);
xor U6783 (N_6783,N_6307,N_6404);
xor U6784 (N_6784,N_6138,N_6313);
and U6785 (N_6785,N_6041,N_6234);
nand U6786 (N_6786,N_6203,N_6199);
nor U6787 (N_6787,N_6327,N_6232);
nand U6788 (N_6788,N_6458,N_6010);
nor U6789 (N_6789,N_6161,N_6358);
and U6790 (N_6790,N_6389,N_6394);
and U6791 (N_6791,N_6093,N_6438);
or U6792 (N_6792,N_6290,N_6143);
and U6793 (N_6793,N_6319,N_6044);
nor U6794 (N_6794,N_6023,N_6253);
or U6795 (N_6795,N_6057,N_6054);
or U6796 (N_6796,N_6463,N_6274);
or U6797 (N_6797,N_6419,N_6285);
and U6798 (N_6798,N_6421,N_6446);
and U6799 (N_6799,N_6431,N_6437);
nand U6800 (N_6800,N_6496,N_6044);
or U6801 (N_6801,N_6190,N_6162);
and U6802 (N_6802,N_6165,N_6471);
xor U6803 (N_6803,N_6348,N_6288);
xnor U6804 (N_6804,N_6385,N_6098);
nand U6805 (N_6805,N_6185,N_6269);
nor U6806 (N_6806,N_6404,N_6076);
nand U6807 (N_6807,N_6056,N_6405);
nand U6808 (N_6808,N_6406,N_6434);
xor U6809 (N_6809,N_6361,N_6146);
nor U6810 (N_6810,N_6310,N_6423);
and U6811 (N_6811,N_6149,N_6177);
nor U6812 (N_6812,N_6156,N_6195);
xor U6813 (N_6813,N_6118,N_6458);
nor U6814 (N_6814,N_6423,N_6307);
nor U6815 (N_6815,N_6223,N_6498);
xnor U6816 (N_6816,N_6281,N_6044);
nand U6817 (N_6817,N_6453,N_6161);
and U6818 (N_6818,N_6203,N_6207);
nand U6819 (N_6819,N_6094,N_6192);
xor U6820 (N_6820,N_6345,N_6188);
nand U6821 (N_6821,N_6352,N_6325);
xnor U6822 (N_6822,N_6298,N_6478);
nor U6823 (N_6823,N_6459,N_6057);
or U6824 (N_6824,N_6167,N_6420);
and U6825 (N_6825,N_6386,N_6086);
nor U6826 (N_6826,N_6191,N_6100);
and U6827 (N_6827,N_6125,N_6375);
nand U6828 (N_6828,N_6071,N_6437);
xor U6829 (N_6829,N_6168,N_6492);
xor U6830 (N_6830,N_6399,N_6260);
nand U6831 (N_6831,N_6020,N_6064);
and U6832 (N_6832,N_6322,N_6117);
xor U6833 (N_6833,N_6010,N_6062);
nor U6834 (N_6834,N_6445,N_6432);
or U6835 (N_6835,N_6454,N_6005);
or U6836 (N_6836,N_6110,N_6274);
xor U6837 (N_6837,N_6176,N_6136);
or U6838 (N_6838,N_6014,N_6327);
or U6839 (N_6839,N_6245,N_6268);
nand U6840 (N_6840,N_6046,N_6380);
nand U6841 (N_6841,N_6188,N_6327);
and U6842 (N_6842,N_6379,N_6099);
nand U6843 (N_6843,N_6146,N_6296);
nand U6844 (N_6844,N_6499,N_6077);
and U6845 (N_6845,N_6440,N_6293);
nand U6846 (N_6846,N_6401,N_6170);
and U6847 (N_6847,N_6057,N_6477);
nor U6848 (N_6848,N_6491,N_6120);
xnor U6849 (N_6849,N_6468,N_6284);
nor U6850 (N_6850,N_6051,N_6054);
and U6851 (N_6851,N_6261,N_6416);
and U6852 (N_6852,N_6202,N_6454);
xor U6853 (N_6853,N_6094,N_6427);
and U6854 (N_6854,N_6198,N_6406);
and U6855 (N_6855,N_6470,N_6321);
nand U6856 (N_6856,N_6211,N_6400);
nor U6857 (N_6857,N_6297,N_6380);
nand U6858 (N_6858,N_6303,N_6389);
nor U6859 (N_6859,N_6226,N_6011);
or U6860 (N_6860,N_6154,N_6440);
or U6861 (N_6861,N_6239,N_6091);
and U6862 (N_6862,N_6431,N_6189);
or U6863 (N_6863,N_6346,N_6429);
nand U6864 (N_6864,N_6136,N_6259);
or U6865 (N_6865,N_6349,N_6045);
xor U6866 (N_6866,N_6034,N_6045);
nand U6867 (N_6867,N_6407,N_6452);
nand U6868 (N_6868,N_6109,N_6206);
and U6869 (N_6869,N_6047,N_6098);
nor U6870 (N_6870,N_6208,N_6404);
xnor U6871 (N_6871,N_6171,N_6134);
or U6872 (N_6872,N_6033,N_6116);
or U6873 (N_6873,N_6161,N_6184);
or U6874 (N_6874,N_6232,N_6345);
nor U6875 (N_6875,N_6106,N_6107);
xor U6876 (N_6876,N_6387,N_6105);
or U6877 (N_6877,N_6321,N_6090);
nand U6878 (N_6878,N_6097,N_6003);
and U6879 (N_6879,N_6152,N_6082);
nand U6880 (N_6880,N_6377,N_6481);
nor U6881 (N_6881,N_6195,N_6349);
and U6882 (N_6882,N_6038,N_6247);
or U6883 (N_6883,N_6095,N_6394);
and U6884 (N_6884,N_6323,N_6203);
xnor U6885 (N_6885,N_6353,N_6499);
or U6886 (N_6886,N_6069,N_6210);
and U6887 (N_6887,N_6193,N_6130);
xnor U6888 (N_6888,N_6294,N_6065);
xnor U6889 (N_6889,N_6004,N_6050);
or U6890 (N_6890,N_6430,N_6421);
xnor U6891 (N_6891,N_6261,N_6353);
xnor U6892 (N_6892,N_6084,N_6163);
xnor U6893 (N_6893,N_6466,N_6160);
and U6894 (N_6894,N_6393,N_6495);
xnor U6895 (N_6895,N_6306,N_6452);
nand U6896 (N_6896,N_6013,N_6341);
and U6897 (N_6897,N_6245,N_6221);
xor U6898 (N_6898,N_6467,N_6190);
xnor U6899 (N_6899,N_6098,N_6224);
nand U6900 (N_6900,N_6374,N_6491);
or U6901 (N_6901,N_6305,N_6015);
nor U6902 (N_6902,N_6374,N_6372);
nand U6903 (N_6903,N_6290,N_6124);
nand U6904 (N_6904,N_6037,N_6376);
nor U6905 (N_6905,N_6187,N_6413);
xnor U6906 (N_6906,N_6146,N_6142);
nor U6907 (N_6907,N_6377,N_6287);
xor U6908 (N_6908,N_6440,N_6142);
nand U6909 (N_6909,N_6390,N_6474);
xor U6910 (N_6910,N_6134,N_6489);
or U6911 (N_6911,N_6493,N_6168);
xor U6912 (N_6912,N_6263,N_6169);
nand U6913 (N_6913,N_6351,N_6102);
and U6914 (N_6914,N_6207,N_6225);
nand U6915 (N_6915,N_6013,N_6220);
nor U6916 (N_6916,N_6257,N_6424);
and U6917 (N_6917,N_6354,N_6428);
and U6918 (N_6918,N_6045,N_6413);
or U6919 (N_6919,N_6311,N_6388);
nor U6920 (N_6920,N_6351,N_6362);
or U6921 (N_6921,N_6351,N_6318);
or U6922 (N_6922,N_6305,N_6253);
or U6923 (N_6923,N_6237,N_6390);
xnor U6924 (N_6924,N_6452,N_6459);
or U6925 (N_6925,N_6369,N_6180);
or U6926 (N_6926,N_6443,N_6417);
nor U6927 (N_6927,N_6309,N_6206);
xor U6928 (N_6928,N_6484,N_6214);
or U6929 (N_6929,N_6190,N_6079);
or U6930 (N_6930,N_6391,N_6224);
xnor U6931 (N_6931,N_6363,N_6074);
nand U6932 (N_6932,N_6484,N_6490);
xnor U6933 (N_6933,N_6359,N_6260);
or U6934 (N_6934,N_6141,N_6166);
or U6935 (N_6935,N_6022,N_6419);
and U6936 (N_6936,N_6046,N_6410);
or U6937 (N_6937,N_6020,N_6075);
nand U6938 (N_6938,N_6216,N_6241);
nor U6939 (N_6939,N_6239,N_6311);
nand U6940 (N_6940,N_6046,N_6348);
and U6941 (N_6941,N_6128,N_6077);
and U6942 (N_6942,N_6347,N_6356);
or U6943 (N_6943,N_6189,N_6290);
nor U6944 (N_6944,N_6403,N_6468);
nand U6945 (N_6945,N_6244,N_6396);
xor U6946 (N_6946,N_6076,N_6297);
and U6947 (N_6947,N_6304,N_6297);
xor U6948 (N_6948,N_6380,N_6477);
or U6949 (N_6949,N_6121,N_6182);
or U6950 (N_6950,N_6125,N_6465);
or U6951 (N_6951,N_6398,N_6383);
xnor U6952 (N_6952,N_6098,N_6323);
and U6953 (N_6953,N_6460,N_6349);
and U6954 (N_6954,N_6406,N_6226);
and U6955 (N_6955,N_6372,N_6228);
xor U6956 (N_6956,N_6487,N_6124);
nand U6957 (N_6957,N_6376,N_6227);
nand U6958 (N_6958,N_6170,N_6080);
nor U6959 (N_6959,N_6076,N_6020);
or U6960 (N_6960,N_6317,N_6431);
and U6961 (N_6961,N_6152,N_6083);
nor U6962 (N_6962,N_6285,N_6189);
or U6963 (N_6963,N_6170,N_6376);
or U6964 (N_6964,N_6459,N_6244);
or U6965 (N_6965,N_6038,N_6073);
and U6966 (N_6966,N_6368,N_6140);
and U6967 (N_6967,N_6331,N_6085);
and U6968 (N_6968,N_6458,N_6216);
or U6969 (N_6969,N_6417,N_6134);
xor U6970 (N_6970,N_6298,N_6237);
or U6971 (N_6971,N_6264,N_6141);
or U6972 (N_6972,N_6480,N_6114);
nor U6973 (N_6973,N_6158,N_6283);
nor U6974 (N_6974,N_6368,N_6424);
nand U6975 (N_6975,N_6150,N_6440);
nor U6976 (N_6976,N_6347,N_6495);
nand U6977 (N_6977,N_6420,N_6252);
nor U6978 (N_6978,N_6187,N_6211);
nor U6979 (N_6979,N_6467,N_6138);
xnor U6980 (N_6980,N_6458,N_6018);
xor U6981 (N_6981,N_6163,N_6413);
or U6982 (N_6982,N_6292,N_6294);
and U6983 (N_6983,N_6355,N_6065);
xnor U6984 (N_6984,N_6492,N_6159);
xor U6985 (N_6985,N_6441,N_6347);
and U6986 (N_6986,N_6043,N_6242);
nand U6987 (N_6987,N_6135,N_6098);
nand U6988 (N_6988,N_6000,N_6197);
and U6989 (N_6989,N_6063,N_6460);
or U6990 (N_6990,N_6074,N_6427);
nand U6991 (N_6991,N_6452,N_6130);
nand U6992 (N_6992,N_6145,N_6101);
nor U6993 (N_6993,N_6181,N_6414);
or U6994 (N_6994,N_6386,N_6483);
nor U6995 (N_6995,N_6283,N_6299);
xnor U6996 (N_6996,N_6301,N_6156);
nor U6997 (N_6997,N_6413,N_6421);
or U6998 (N_6998,N_6368,N_6116);
and U6999 (N_6999,N_6021,N_6048);
or U7000 (N_7000,N_6612,N_6966);
or U7001 (N_7001,N_6946,N_6643);
nand U7002 (N_7002,N_6658,N_6860);
or U7003 (N_7003,N_6929,N_6594);
nand U7004 (N_7004,N_6707,N_6665);
nand U7005 (N_7005,N_6950,N_6920);
and U7006 (N_7006,N_6818,N_6911);
xnor U7007 (N_7007,N_6502,N_6786);
nor U7008 (N_7008,N_6849,N_6627);
nor U7009 (N_7009,N_6930,N_6791);
xnor U7010 (N_7010,N_6826,N_6799);
and U7011 (N_7011,N_6616,N_6656);
or U7012 (N_7012,N_6905,N_6994);
and U7013 (N_7013,N_6728,N_6614);
and U7014 (N_7014,N_6916,N_6872);
and U7015 (N_7015,N_6809,N_6664);
or U7016 (N_7016,N_6582,N_6843);
nand U7017 (N_7017,N_6825,N_6764);
or U7018 (N_7018,N_6793,N_6592);
and U7019 (N_7019,N_6647,N_6673);
or U7020 (N_7020,N_6935,N_6589);
or U7021 (N_7021,N_6778,N_6628);
xor U7022 (N_7022,N_6514,N_6981);
or U7023 (N_7023,N_6524,N_6671);
xor U7024 (N_7024,N_6678,N_6549);
nor U7025 (N_7025,N_6918,N_6781);
and U7026 (N_7026,N_6962,N_6898);
and U7027 (N_7027,N_6827,N_6856);
or U7028 (N_7028,N_6895,N_6650);
nand U7029 (N_7029,N_6545,N_6753);
nor U7030 (N_7030,N_6590,N_6813);
or U7031 (N_7031,N_6765,N_6631);
nand U7032 (N_7032,N_6880,N_6749);
and U7033 (N_7033,N_6544,N_6700);
or U7034 (N_7034,N_6836,N_6894);
nand U7035 (N_7035,N_6882,N_6539);
nor U7036 (N_7036,N_6639,N_6638);
nand U7037 (N_7037,N_6912,N_6711);
nor U7038 (N_7038,N_6719,N_6941);
xor U7039 (N_7039,N_6967,N_6597);
nor U7040 (N_7040,N_6889,N_6522);
and U7041 (N_7041,N_6774,N_6997);
nand U7042 (N_7042,N_6610,N_6810);
and U7043 (N_7043,N_6525,N_6561);
or U7044 (N_7044,N_6542,N_6595);
or U7045 (N_7045,N_6585,N_6931);
xnor U7046 (N_7046,N_6833,N_6623);
nor U7047 (N_7047,N_6835,N_6657);
and U7048 (N_7048,N_6646,N_6988);
nand U7049 (N_7049,N_6928,N_6709);
xnor U7050 (N_7050,N_6800,N_6990);
and U7051 (N_7051,N_6903,N_6679);
xnor U7052 (N_7052,N_6901,N_6807);
and U7053 (N_7053,N_6571,N_6513);
nor U7054 (N_7054,N_6789,N_6821);
xor U7055 (N_7055,N_6831,N_6649);
xor U7056 (N_7056,N_6980,N_6755);
xnor U7057 (N_7057,N_6653,N_6863);
and U7058 (N_7058,N_6529,N_6998);
nor U7059 (N_7059,N_6566,N_6570);
and U7060 (N_7060,N_6685,N_6976);
nand U7061 (N_7061,N_6769,N_6668);
xor U7062 (N_7062,N_6986,N_6943);
and U7063 (N_7063,N_6521,N_6977);
and U7064 (N_7064,N_6557,N_6838);
nor U7065 (N_7065,N_6734,N_6878);
and U7066 (N_7066,N_6691,N_6572);
nor U7067 (N_7067,N_6805,N_6982);
xnor U7068 (N_7068,N_6927,N_6761);
xor U7069 (N_7069,N_6985,N_6694);
nand U7070 (N_7070,N_6758,N_6532);
nand U7071 (N_7071,N_6523,N_6580);
xnor U7072 (N_7072,N_6842,N_6900);
or U7073 (N_7073,N_6968,N_6690);
or U7074 (N_7074,N_6538,N_6747);
xor U7075 (N_7075,N_6559,N_6558);
or U7076 (N_7076,N_6716,N_6899);
nor U7077 (N_7077,N_6869,N_6617);
and U7078 (N_7078,N_6698,N_6748);
nand U7079 (N_7079,N_6562,N_6785);
and U7080 (N_7080,N_6507,N_6615);
or U7081 (N_7081,N_6987,N_6890);
nand U7082 (N_7082,N_6555,N_6727);
xor U7083 (N_7083,N_6969,N_6938);
or U7084 (N_7084,N_6787,N_6721);
nand U7085 (N_7085,N_6605,N_6515);
and U7086 (N_7086,N_6923,N_6548);
nand U7087 (N_7087,N_6752,N_6763);
and U7088 (N_7088,N_6501,N_6921);
and U7089 (N_7089,N_6955,N_6588);
xnor U7090 (N_7090,N_6788,N_6873);
nand U7091 (N_7091,N_6822,N_6546);
nor U7092 (N_7092,N_6645,N_6725);
and U7093 (N_7093,N_6634,N_6622);
nor U7094 (N_7094,N_6676,N_6924);
nand U7095 (N_7095,N_6926,N_6803);
or U7096 (N_7096,N_6971,N_6892);
and U7097 (N_7097,N_6888,N_6919);
xnor U7098 (N_7098,N_6543,N_6508);
and U7099 (N_7099,N_6754,N_6773);
or U7100 (N_7100,N_6573,N_6680);
or U7101 (N_7101,N_6531,N_6840);
xnor U7102 (N_7102,N_6670,N_6798);
nor U7103 (N_7103,N_6701,N_6995);
or U7104 (N_7104,N_6886,N_6942);
and U7105 (N_7105,N_6669,N_6584);
nand U7106 (N_7106,N_6815,N_6801);
and U7107 (N_7107,N_6984,N_6660);
xor U7108 (N_7108,N_6864,N_6858);
or U7109 (N_7109,N_6552,N_6904);
and U7110 (N_7110,N_6767,N_6794);
xor U7111 (N_7111,N_6723,N_6510);
nor U7112 (N_7112,N_6704,N_6934);
or U7113 (N_7113,N_6739,N_6677);
nor U7114 (N_7114,N_6732,N_6782);
and U7115 (N_7115,N_6951,N_6556);
or U7116 (N_7116,N_6817,N_6714);
nand U7117 (N_7117,N_6699,N_6611);
nor U7118 (N_7118,N_6599,N_6845);
xnor U7119 (N_7119,N_6848,N_6500);
or U7120 (N_7120,N_6688,N_6632);
nand U7121 (N_7121,N_6760,N_6506);
nand U7122 (N_7122,N_6578,N_6850);
xor U7123 (N_7123,N_6541,N_6925);
nor U7124 (N_7124,N_6766,N_6745);
nor U7125 (N_7125,N_6750,N_6738);
and U7126 (N_7126,N_6783,N_6576);
nand U7127 (N_7127,N_6563,N_6965);
or U7128 (N_7128,N_6839,N_6915);
and U7129 (N_7129,N_6624,N_6636);
xor U7130 (N_7130,N_6870,N_6652);
nor U7131 (N_7131,N_6855,N_6812);
or U7132 (N_7132,N_6762,N_6944);
xor U7133 (N_7133,N_6682,N_6596);
or U7134 (N_7134,N_6724,N_6936);
nand U7135 (N_7135,N_6587,N_6973);
xnor U7136 (N_7136,N_6983,N_6593);
xor U7137 (N_7137,N_6512,N_6746);
xor U7138 (N_7138,N_6841,N_6641);
xnor U7139 (N_7139,N_6874,N_6644);
xor U7140 (N_7140,N_6737,N_6681);
and U7141 (N_7141,N_6564,N_6829);
nor U7142 (N_7142,N_6846,N_6569);
nor U7143 (N_7143,N_6744,N_6866);
or U7144 (N_7144,N_6948,N_6996);
or U7145 (N_7145,N_6586,N_6875);
nor U7146 (N_7146,N_6796,N_6560);
or U7147 (N_7147,N_6527,N_6991);
nand U7148 (N_7148,N_6876,N_6674);
xnor U7149 (N_7149,N_6705,N_6713);
nand U7150 (N_7150,N_6715,N_6742);
xnor U7151 (N_7151,N_6567,N_6910);
and U7152 (N_7152,N_6516,N_6712);
nand U7153 (N_7153,N_6683,N_6600);
xor U7154 (N_7154,N_6537,N_6811);
nor U7155 (N_7155,N_6528,N_6702);
nor U7156 (N_7156,N_6625,N_6979);
and U7157 (N_7157,N_6802,N_6933);
nor U7158 (N_7158,N_6853,N_6603);
nor U7159 (N_7159,N_6814,N_6772);
xor U7160 (N_7160,N_6503,N_6651);
nand U7161 (N_7161,N_6891,N_6629);
xor U7162 (N_7162,N_6779,N_6871);
xor U7163 (N_7163,N_6893,N_6867);
and U7164 (N_7164,N_6844,N_6518);
nand U7165 (N_7165,N_6897,N_6575);
and U7166 (N_7166,N_6684,N_6630);
or U7167 (N_7167,N_6511,N_6854);
nor U7168 (N_7168,N_6945,N_6581);
nand U7169 (N_7169,N_6759,N_6743);
nand U7170 (N_7170,N_6663,N_6536);
xor U7171 (N_7171,N_6740,N_6686);
nand U7172 (N_7172,N_6620,N_6547);
or U7173 (N_7173,N_6914,N_6808);
and U7174 (N_7174,N_6731,N_6659);
or U7175 (N_7175,N_6703,N_6553);
nand U7176 (N_7176,N_6540,N_6949);
nor U7177 (N_7177,N_6917,N_6952);
xnor U7178 (N_7178,N_6533,N_6852);
or U7179 (N_7179,N_6520,N_6780);
or U7180 (N_7180,N_6751,N_6913);
or U7181 (N_7181,N_6654,N_6720);
xnor U7182 (N_7182,N_6633,N_6879);
xnor U7183 (N_7183,N_6865,N_6607);
nor U7184 (N_7184,N_6637,N_6862);
xor U7185 (N_7185,N_6618,N_6608);
nor U7186 (N_7186,N_6828,N_6861);
or U7187 (N_7187,N_6550,N_6859);
xor U7188 (N_7188,N_6777,N_6598);
and U7189 (N_7189,N_6722,N_6957);
xnor U7190 (N_7190,N_6974,N_6830);
nand U7191 (N_7191,N_6847,N_6733);
nand U7192 (N_7192,N_6609,N_6790);
nor U7193 (N_7193,N_6517,N_6837);
and U7194 (N_7194,N_6613,N_6519);
nand U7195 (N_7195,N_6907,N_6735);
xnor U7196 (N_7196,N_6851,N_6554);
or U7197 (N_7197,N_6989,N_6961);
and U7198 (N_7198,N_6565,N_6675);
nand U7199 (N_7199,N_6574,N_6741);
xor U7200 (N_7200,N_6922,N_6756);
or U7201 (N_7201,N_6689,N_6726);
or U7202 (N_7202,N_6908,N_6823);
or U7203 (N_7203,N_6963,N_6885);
nor U7204 (N_7204,N_6906,N_6583);
nor U7205 (N_7205,N_6978,N_6692);
xor U7206 (N_7206,N_6626,N_6797);
xor U7207 (N_7207,N_6832,N_6784);
or U7208 (N_7208,N_6717,N_6940);
nand U7209 (N_7209,N_6954,N_6887);
and U7210 (N_7210,N_6551,N_6509);
nor U7211 (N_7211,N_6992,N_6619);
nor U7212 (N_7212,N_6526,N_6606);
and U7213 (N_7213,N_6857,N_6792);
nor U7214 (N_7214,N_6956,N_6775);
nand U7215 (N_7215,N_6655,N_6667);
or U7216 (N_7216,N_6770,N_6909);
nor U7217 (N_7217,N_6648,N_6868);
nor U7218 (N_7218,N_6687,N_6729);
or U7219 (N_7219,N_6993,N_6964);
and U7220 (N_7220,N_6602,N_6568);
nand U7221 (N_7221,N_6939,N_6534);
and U7222 (N_7222,N_6696,N_6672);
nor U7223 (N_7223,N_6881,N_6975);
or U7224 (N_7224,N_6601,N_6706);
and U7225 (N_7225,N_6824,N_6718);
nand U7226 (N_7226,N_6972,N_6970);
nand U7227 (N_7227,N_6730,N_6577);
nand U7228 (N_7228,N_6884,N_6591);
nor U7229 (N_7229,N_6504,N_6795);
nand U7230 (N_7230,N_6947,N_6932);
nand U7231 (N_7231,N_6960,N_6710);
or U7232 (N_7232,N_6806,N_6896);
nor U7233 (N_7233,N_6820,N_6768);
xor U7234 (N_7234,N_6877,N_6902);
nand U7235 (N_7235,N_6604,N_6959);
nand U7236 (N_7236,N_6736,N_6579);
xnor U7237 (N_7237,N_6958,N_6883);
or U7238 (N_7238,N_6666,N_6776);
nor U7239 (N_7239,N_6505,N_6535);
nor U7240 (N_7240,N_6640,N_6697);
or U7241 (N_7241,N_6819,N_6771);
nand U7242 (N_7242,N_6530,N_6999);
xor U7243 (N_7243,N_6693,N_6953);
and U7244 (N_7244,N_6757,N_6834);
xnor U7245 (N_7245,N_6937,N_6642);
nand U7246 (N_7246,N_6635,N_6662);
nand U7247 (N_7247,N_6695,N_6621);
nand U7248 (N_7248,N_6708,N_6804);
nand U7249 (N_7249,N_6816,N_6661);
or U7250 (N_7250,N_6597,N_6956);
xnor U7251 (N_7251,N_6941,N_6848);
or U7252 (N_7252,N_6945,N_6771);
or U7253 (N_7253,N_6665,N_6893);
or U7254 (N_7254,N_6528,N_6845);
and U7255 (N_7255,N_6655,N_6645);
xnor U7256 (N_7256,N_6823,N_6854);
or U7257 (N_7257,N_6636,N_6538);
nor U7258 (N_7258,N_6922,N_6749);
xnor U7259 (N_7259,N_6865,N_6977);
nor U7260 (N_7260,N_6537,N_6858);
nor U7261 (N_7261,N_6627,N_6576);
and U7262 (N_7262,N_6865,N_6648);
and U7263 (N_7263,N_6895,N_6514);
nand U7264 (N_7264,N_6843,N_6528);
nor U7265 (N_7265,N_6941,N_6688);
and U7266 (N_7266,N_6640,N_6664);
nand U7267 (N_7267,N_6517,N_6635);
nand U7268 (N_7268,N_6808,N_6990);
nand U7269 (N_7269,N_6867,N_6988);
and U7270 (N_7270,N_6833,N_6758);
nor U7271 (N_7271,N_6805,N_6635);
xor U7272 (N_7272,N_6719,N_6805);
or U7273 (N_7273,N_6774,N_6501);
and U7274 (N_7274,N_6571,N_6633);
or U7275 (N_7275,N_6535,N_6654);
nand U7276 (N_7276,N_6880,N_6990);
xnor U7277 (N_7277,N_6903,N_6865);
nor U7278 (N_7278,N_6534,N_6949);
nand U7279 (N_7279,N_6927,N_6830);
and U7280 (N_7280,N_6686,N_6595);
or U7281 (N_7281,N_6744,N_6563);
nor U7282 (N_7282,N_6787,N_6617);
nand U7283 (N_7283,N_6813,N_6831);
nor U7284 (N_7284,N_6531,N_6501);
nand U7285 (N_7285,N_6885,N_6668);
nand U7286 (N_7286,N_6563,N_6547);
nor U7287 (N_7287,N_6960,N_6821);
nand U7288 (N_7288,N_6763,N_6561);
nand U7289 (N_7289,N_6925,N_6955);
nand U7290 (N_7290,N_6504,N_6958);
and U7291 (N_7291,N_6567,N_6712);
nor U7292 (N_7292,N_6714,N_6797);
and U7293 (N_7293,N_6654,N_6626);
nor U7294 (N_7294,N_6982,N_6516);
or U7295 (N_7295,N_6929,N_6937);
nand U7296 (N_7296,N_6588,N_6944);
nand U7297 (N_7297,N_6764,N_6677);
nand U7298 (N_7298,N_6585,N_6968);
and U7299 (N_7299,N_6847,N_6566);
or U7300 (N_7300,N_6762,N_6860);
xnor U7301 (N_7301,N_6532,N_6928);
nand U7302 (N_7302,N_6938,N_6750);
xor U7303 (N_7303,N_6827,N_6931);
nor U7304 (N_7304,N_6906,N_6886);
nor U7305 (N_7305,N_6761,N_6533);
or U7306 (N_7306,N_6561,N_6573);
nand U7307 (N_7307,N_6914,N_6873);
nor U7308 (N_7308,N_6799,N_6539);
nand U7309 (N_7309,N_6843,N_6515);
or U7310 (N_7310,N_6652,N_6758);
or U7311 (N_7311,N_6682,N_6510);
nand U7312 (N_7312,N_6969,N_6669);
nand U7313 (N_7313,N_6710,N_6996);
and U7314 (N_7314,N_6791,N_6794);
nor U7315 (N_7315,N_6740,N_6849);
xor U7316 (N_7316,N_6871,N_6537);
xor U7317 (N_7317,N_6670,N_6857);
and U7318 (N_7318,N_6645,N_6876);
nor U7319 (N_7319,N_6722,N_6522);
or U7320 (N_7320,N_6780,N_6702);
xnor U7321 (N_7321,N_6695,N_6967);
and U7322 (N_7322,N_6725,N_6960);
or U7323 (N_7323,N_6932,N_6609);
nor U7324 (N_7324,N_6835,N_6531);
or U7325 (N_7325,N_6890,N_6901);
nor U7326 (N_7326,N_6578,N_6505);
and U7327 (N_7327,N_6801,N_6886);
nand U7328 (N_7328,N_6542,N_6592);
xnor U7329 (N_7329,N_6711,N_6626);
nor U7330 (N_7330,N_6543,N_6950);
and U7331 (N_7331,N_6593,N_6562);
and U7332 (N_7332,N_6531,N_6640);
xnor U7333 (N_7333,N_6584,N_6719);
and U7334 (N_7334,N_6926,N_6618);
and U7335 (N_7335,N_6896,N_6509);
or U7336 (N_7336,N_6864,N_6622);
nor U7337 (N_7337,N_6948,N_6748);
nand U7338 (N_7338,N_6870,N_6982);
and U7339 (N_7339,N_6890,N_6894);
nor U7340 (N_7340,N_6882,N_6916);
or U7341 (N_7341,N_6779,N_6662);
xor U7342 (N_7342,N_6507,N_6622);
nor U7343 (N_7343,N_6913,N_6842);
or U7344 (N_7344,N_6554,N_6541);
or U7345 (N_7345,N_6978,N_6625);
nand U7346 (N_7346,N_6648,N_6552);
nor U7347 (N_7347,N_6942,N_6798);
nand U7348 (N_7348,N_6599,N_6789);
and U7349 (N_7349,N_6870,N_6548);
nand U7350 (N_7350,N_6755,N_6660);
xor U7351 (N_7351,N_6973,N_6776);
xnor U7352 (N_7352,N_6794,N_6508);
xnor U7353 (N_7353,N_6581,N_6906);
nand U7354 (N_7354,N_6650,N_6893);
and U7355 (N_7355,N_6558,N_6976);
or U7356 (N_7356,N_6619,N_6673);
nor U7357 (N_7357,N_6806,N_6949);
nand U7358 (N_7358,N_6864,N_6761);
and U7359 (N_7359,N_6524,N_6803);
or U7360 (N_7360,N_6659,N_6765);
and U7361 (N_7361,N_6882,N_6687);
or U7362 (N_7362,N_6934,N_6532);
nand U7363 (N_7363,N_6959,N_6904);
and U7364 (N_7364,N_6989,N_6672);
xor U7365 (N_7365,N_6835,N_6537);
or U7366 (N_7366,N_6709,N_6715);
nand U7367 (N_7367,N_6634,N_6718);
and U7368 (N_7368,N_6643,N_6968);
xor U7369 (N_7369,N_6539,N_6982);
nand U7370 (N_7370,N_6584,N_6552);
nor U7371 (N_7371,N_6810,N_6644);
nand U7372 (N_7372,N_6859,N_6974);
and U7373 (N_7373,N_6687,N_6838);
nand U7374 (N_7374,N_6860,N_6937);
nand U7375 (N_7375,N_6564,N_6995);
and U7376 (N_7376,N_6661,N_6914);
nor U7377 (N_7377,N_6712,N_6643);
nor U7378 (N_7378,N_6824,N_6711);
xor U7379 (N_7379,N_6589,N_6655);
nand U7380 (N_7380,N_6865,N_6905);
xor U7381 (N_7381,N_6783,N_6503);
xnor U7382 (N_7382,N_6929,N_6676);
and U7383 (N_7383,N_6503,N_6743);
or U7384 (N_7384,N_6768,N_6833);
or U7385 (N_7385,N_6832,N_6935);
and U7386 (N_7386,N_6968,N_6799);
or U7387 (N_7387,N_6926,N_6965);
nand U7388 (N_7388,N_6829,N_6792);
nand U7389 (N_7389,N_6920,N_6744);
nand U7390 (N_7390,N_6631,N_6812);
or U7391 (N_7391,N_6754,N_6594);
nand U7392 (N_7392,N_6929,N_6841);
nor U7393 (N_7393,N_6687,N_6706);
xnor U7394 (N_7394,N_6867,N_6848);
xor U7395 (N_7395,N_6973,N_6610);
xnor U7396 (N_7396,N_6861,N_6933);
or U7397 (N_7397,N_6832,N_6585);
or U7398 (N_7398,N_6821,N_6526);
and U7399 (N_7399,N_6625,N_6653);
or U7400 (N_7400,N_6503,N_6853);
nand U7401 (N_7401,N_6612,N_6539);
nand U7402 (N_7402,N_6759,N_6877);
nand U7403 (N_7403,N_6547,N_6973);
xor U7404 (N_7404,N_6808,N_6754);
and U7405 (N_7405,N_6937,N_6756);
or U7406 (N_7406,N_6518,N_6884);
nand U7407 (N_7407,N_6652,N_6762);
or U7408 (N_7408,N_6614,N_6741);
nor U7409 (N_7409,N_6969,N_6521);
and U7410 (N_7410,N_6793,N_6741);
nor U7411 (N_7411,N_6892,N_6520);
nand U7412 (N_7412,N_6595,N_6533);
xor U7413 (N_7413,N_6729,N_6559);
or U7414 (N_7414,N_6521,N_6774);
and U7415 (N_7415,N_6775,N_6508);
nor U7416 (N_7416,N_6796,N_6775);
xor U7417 (N_7417,N_6855,N_6548);
nand U7418 (N_7418,N_6625,N_6614);
nand U7419 (N_7419,N_6590,N_6658);
xnor U7420 (N_7420,N_6583,N_6607);
or U7421 (N_7421,N_6566,N_6762);
or U7422 (N_7422,N_6986,N_6666);
and U7423 (N_7423,N_6646,N_6744);
nor U7424 (N_7424,N_6976,N_6874);
xnor U7425 (N_7425,N_6842,N_6942);
nor U7426 (N_7426,N_6924,N_6679);
or U7427 (N_7427,N_6574,N_6788);
or U7428 (N_7428,N_6603,N_6881);
nand U7429 (N_7429,N_6556,N_6994);
nand U7430 (N_7430,N_6817,N_6971);
nand U7431 (N_7431,N_6904,N_6584);
and U7432 (N_7432,N_6550,N_6875);
or U7433 (N_7433,N_6519,N_6950);
or U7434 (N_7434,N_6897,N_6540);
or U7435 (N_7435,N_6744,N_6720);
nand U7436 (N_7436,N_6930,N_6604);
xor U7437 (N_7437,N_6542,N_6598);
xnor U7438 (N_7438,N_6663,N_6683);
nand U7439 (N_7439,N_6804,N_6930);
and U7440 (N_7440,N_6909,N_6849);
nor U7441 (N_7441,N_6532,N_6653);
nor U7442 (N_7442,N_6758,N_6651);
nand U7443 (N_7443,N_6587,N_6857);
xnor U7444 (N_7444,N_6701,N_6569);
xnor U7445 (N_7445,N_6746,N_6898);
and U7446 (N_7446,N_6810,N_6818);
and U7447 (N_7447,N_6954,N_6883);
nor U7448 (N_7448,N_6733,N_6634);
or U7449 (N_7449,N_6540,N_6595);
nor U7450 (N_7450,N_6768,N_6713);
nand U7451 (N_7451,N_6932,N_6975);
nand U7452 (N_7452,N_6810,N_6786);
nand U7453 (N_7453,N_6698,N_6928);
and U7454 (N_7454,N_6762,N_6997);
or U7455 (N_7455,N_6958,N_6523);
nor U7456 (N_7456,N_6858,N_6685);
or U7457 (N_7457,N_6514,N_6865);
nand U7458 (N_7458,N_6694,N_6999);
xnor U7459 (N_7459,N_6763,N_6633);
nor U7460 (N_7460,N_6760,N_6911);
nand U7461 (N_7461,N_6813,N_6870);
xor U7462 (N_7462,N_6814,N_6763);
xor U7463 (N_7463,N_6847,N_6891);
nor U7464 (N_7464,N_6840,N_6991);
and U7465 (N_7465,N_6864,N_6870);
or U7466 (N_7466,N_6700,N_6554);
xor U7467 (N_7467,N_6615,N_6580);
or U7468 (N_7468,N_6963,N_6655);
or U7469 (N_7469,N_6853,N_6828);
or U7470 (N_7470,N_6973,N_6509);
nor U7471 (N_7471,N_6937,N_6957);
nand U7472 (N_7472,N_6667,N_6971);
nor U7473 (N_7473,N_6976,N_6597);
xnor U7474 (N_7474,N_6665,N_6895);
or U7475 (N_7475,N_6808,N_6565);
nor U7476 (N_7476,N_6879,N_6775);
nor U7477 (N_7477,N_6722,N_6684);
and U7478 (N_7478,N_6679,N_6833);
nand U7479 (N_7479,N_6777,N_6710);
or U7480 (N_7480,N_6856,N_6951);
nand U7481 (N_7481,N_6505,N_6757);
or U7482 (N_7482,N_6702,N_6738);
and U7483 (N_7483,N_6908,N_6742);
or U7484 (N_7484,N_6880,N_6628);
or U7485 (N_7485,N_6708,N_6686);
or U7486 (N_7486,N_6918,N_6745);
nand U7487 (N_7487,N_6673,N_6995);
xor U7488 (N_7488,N_6630,N_6811);
nor U7489 (N_7489,N_6558,N_6772);
nor U7490 (N_7490,N_6911,N_6798);
and U7491 (N_7491,N_6945,N_6529);
xnor U7492 (N_7492,N_6603,N_6902);
nand U7493 (N_7493,N_6538,N_6815);
nand U7494 (N_7494,N_6568,N_6607);
xnor U7495 (N_7495,N_6530,N_6511);
and U7496 (N_7496,N_6957,N_6653);
and U7497 (N_7497,N_6702,N_6973);
or U7498 (N_7498,N_6738,N_6784);
or U7499 (N_7499,N_6530,N_6626);
nor U7500 (N_7500,N_7147,N_7410);
nand U7501 (N_7501,N_7019,N_7104);
nand U7502 (N_7502,N_7471,N_7442);
xor U7503 (N_7503,N_7214,N_7455);
or U7504 (N_7504,N_7129,N_7420);
xor U7505 (N_7505,N_7320,N_7392);
nor U7506 (N_7506,N_7218,N_7027);
nand U7507 (N_7507,N_7252,N_7154);
nor U7508 (N_7508,N_7444,N_7482);
nor U7509 (N_7509,N_7241,N_7174);
nor U7510 (N_7510,N_7059,N_7116);
and U7511 (N_7511,N_7254,N_7283);
or U7512 (N_7512,N_7013,N_7199);
or U7513 (N_7513,N_7441,N_7084);
nor U7514 (N_7514,N_7135,N_7036);
and U7515 (N_7515,N_7494,N_7128);
or U7516 (N_7516,N_7180,N_7220);
or U7517 (N_7517,N_7448,N_7412);
nand U7518 (N_7518,N_7060,N_7038);
and U7519 (N_7519,N_7487,N_7284);
xnor U7520 (N_7520,N_7078,N_7068);
xor U7521 (N_7521,N_7052,N_7243);
nand U7522 (N_7522,N_7237,N_7421);
or U7523 (N_7523,N_7480,N_7163);
or U7524 (N_7524,N_7089,N_7043);
xor U7525 (N_7525,N_7458,N_7271);
xor U7526 (N_7526,N_7427,N_7103);
and U7527 (N_7527,N_7073,N_7428);
and U7528 (N_7528,N_7253,N_7459);
nor U7529 (N_7529,N_7343,N_7273);
nand U7530 (N_7530,N_7045,N_7450);
and U7531 (N_7531,N_7379,N_7493);
nand U7532 (N_7532,N_7106,N_7323);
nor U7533 (N_7533,N_7247,N_7159);
nand U7534 (N_7534,N_7336,N_7461);
nand U7535 (N_7535,N_7091,N_7328);
and U7536 (N_7536,N_7325,N_7235);
xor U7537 (N_7537,N_7173,N_7145);
nand U7538 (N_7538,N_7258,N_7322);
xor U7539 (N_7539,N_7183,N_7404);
nand U7540 (N_7540,N_7489,N_7294);
nor U7541 (N_7541,N_7138,N_7338);
xnor U7542 (N_7542,N_7158,N_7492);
xor U7543 (N_7543,N_7209,N_7100);
and U7544 (N_7544,N_7033,N_7335);
nand U7545 (N_7545,N_7276,N_7035);
nor U7546 (N_7546,N_7403,N_7380);
xnor U7547 (N_7547,N_7113,N_7034);
nand U7548 (N_7548,N_7040,N_7249);
and U7549 (N_7549,N_7202,N_7341);
xnor U7550 (N_7550,N_7472,N_7460);
nand U7551 (N_7551,N_7049,N_7364);
xnor U7552 (N_7552,N_7292,N_7107);
nor U7553 (N_7553,N_7152,N_7346);
nand U7554 (N_7554,N_7288,N_7151);
or U7555 (N_7555,N_7405,N_7082);
or U7556 (N_7556,N_7327,N_7462);
xor U7557 (N_7557,N_7222,N_7474);
nor U7558 (N_7558,N_7190,N_7466);
and U7559 (N_7559,N_7313,N_7132);
nand U7560 (N_7560,N_7014,N_7272);
or U7561 (N_7561,N_7261,N_7074);
nor U7562 (N_7562,N_7340,N_7197);
or U7563 (N_7563,N_7446,N_7375);
nand U7564 (N_7564,N_7318,N_7136);
or U7565 (N_7565,N_7224,N_7080);
and U7566 (N_7566,N_7497,N_7498);
xor U7567 (N_7567,N_7064,N_7130);
xor U7568 (N_7568,N_7115,N_7293);
nand U7569 (N_7569,N_7495,N_7233);
or U7570 (N_7570,N_7026,N_7295);
xnor U7571 (N_7571,N_7246,N_7269);
and U7572 (N_7572,N_7361,N_7211);
and U7573 (N_7573,N_7433,N_7484);
nor U7574 (N_7574,N_7302,N_7285);
xnor U7575 (N_7575,N_7453,N_7331);
and U7576 (N_7576,N_7098,N_7232);
or U7577 (N_7577,N_7030,N_7216);
or U7578 (N_7578,N_7402,N_7170);
and U7579 (N_7579,N_7016,N_7161);
or U7580 (N_7580,N_7081,N_7345);
nand U7581 (N_7581,N_7473,N_7061);
and U7582 (N_7582,N_7390,N_7134);
nand U7583 (N_7583,N_7483,N_7131);
nor U7584 (N_7584,N_7058,N_7382);
and U7585 (N_7585,N_7101,N_7050);
nor U7586 (N_7586,N_7363,N_7150);
or U7587 (N_7587,N_7112,N_7457);
or U7588 (N_7588,N_7437,N_7469);
and U7589 (N_7589,N_7334,N_7260);
xnor U7590 (N_7590,N_7238,N_7093);
nor U7591 (N_7591,N_7426,N_7192);
xnor U7592 (N_7592,N_7406,N_7383);
or U7593 (N_7593,N_7053,N_7447);
nor U7594 (N_7594,N_7413,N_7349);
nand U7595 (N_7595,N_7417,N_7287);
nand U7596 (N_7596,N_7378,N_7465);
and U7597 (N_7597,N_7025,N_7278);
nand U7598 (N_7598,N_7371,N_7386);
or U7599 (N_7599,N_7296,N_7456);
nand U7600 (N_7600,N_7226,N_7401);
xnor U7601 (N_7601,N_7266,N_7308);
or U7602 (N_7602,N_7256,N_7319);
nor U7603 (N_7603,N_7002,N_7251);
nand U7604 (N_7604,N_7374,N_7125);
nand U7605 (N_7605,N_7187,N_7486);
and U7606 (N_7606,N_7029,N_7430);
nand U7607 (N_7607,N_7297,N_7157);
nand U7608 (N_7608,N_7184,N_7291);
nor U7609 (N_7609,N_7124,N_7434);
xnor U7610 (N_7610,N_7339,N_7179);
and U7611 (N_7611,N_7485,N_7468);
and U7612 (N_7612,N_7464,N_7267);
or U7613 (N_7613,N_7423,N_7095);
nor U7614 (N_7614,N_7221,N_7351);
nor U7615 (N_7615,N_7203,N_7481);
nand U7616 (N_7616,N_7146,N_7044);
and U7617 (N_7617,N_7085,N_7149);
xnor U7618 (N_7618,N_7017,N_7072);
or U7619 (N_7619,N_7369,N_7162);
or U7620 (N_7620,N_7281,N_7263);
and U7621 (N_7621,N_7141,N_7181);
or U7622 (N_7622,N_7204,N_7191);
nor U7623 (N_7623,N_7155,N_7309);
xnor U7624 (N_7624,N_7037,N_7153);
xor U7625 (N_7625,N_7164,N_7054);
nor U7626 (N_7626,N_7408,N_7398);
and U7627 (N_7627,N_7219,N_7117);
and U7628 (N_7628,N_7353,N_7206);
nand U7629 (N_7629,N_7217,N_7255);
nor U7630 (N_7630,N_7225,N_7397);
nand U7631 (N_7631,N_7094,N_7182);
nand U7632 (N_7632,N_7165,N_7477);
xor U7633 (N_7633,N_7300,N_7177);
or U7634 (N_7634,N_7223,N_7109);
or U7635 (N_7635,N_7440,N_7324);
or U7636 (N_7636,N_7227,N_7110);
xnor U7637 (N_7637,N_7000,N_7289);
xor U7638 (N_7638,N_7381,N_7264);
and U7639 (N_7639,N_7090,N_7188);
nand U7640 (N_7640,N_7265,N_7051);
or U7641 (N_7641,N_7242,N_7407);
and U7642 (N_7642,N_7126,N_7329);
and U7643 (N_7643,N_7056,N_7001);
and U7644 (N_7644,N_7395,N_7231);
nand U7645 (N_7645,N_7301,N_7372);
or U7646 (N_7646,N_7479,N_7148);
nor U7647 (N_7647,N_7262,N_7449);
xor U7648 (N_7648,N_7032,N_7286);
nor U7649 (N_7649,N_7385,N_7409);
and U7650 (N_7650,N_7496,N_7429);
nor U7651 (N_7651,N_7122,N_7195);
and U7652 (N_7652,N_7311,N_7005);
or U7653 (N_7653,N_7160,N_7021);
nor U7654 (N_7654,N_7229,N_7009);
nand U7655 (N_7655,N_7127,N_7055);
or U7656 (N_7656,N_7451,N_7007);
nor U7657 (N_7657,N_7282,N_7039);
nand U7658 (N_7658,N_7201,N_7020);
nor U7659 (N_7659,N_7042,N_7008);
and U7660 (N_7660,N_7394,N_7057);
nor U7661 (N_7661,N_7389,N_7317);
nor U7662 (N_7662,N_7377,N_7347);
nor U7663 (N_7663,N_7063,N_7077);
nand U7664 (N_7664,N_7337,N_7111);
xnor U7665 (N_7665,N_7259,N_7062);
nand U7666 (N_7666,N_7212,N_7366);
or U7667 (N_7667,N_7169,N_7399);
nor U7668 (N_7668,N_7079,N_7028);
or U7669 (N_7669,N_7333,N_7066);
nand U7670 (N_7670,N_7416,N_7424);
or U7671 (N_7671,N_7321,N_7393);
or U7672 (N_7672,N_7478,N_7373);
or U7673 (N_7673,N_7362,N_7015);
xor U7674 (N_7674,N_7376,N_7245);
or U7675 (N_7675,N_7352,N_7022);
xor U7676 (N_7676,N_7244,N_7355);
nand U7677 (N_7677,N_7445,N_7354);
nor U7678 (N_7678,N_7118,N_7279);
or U7679 (N_7679,N_7290,N_7041);
xnor U7680 (N_7680,N_7023,N_7194);
nor U7681 (N_7681,N_7065,N_7476);
nand U7682 (N_7682,N_7105,N_7010);
xnor U7683 (N_7683,N_7099,N_7280);
nor U7684 (N_7684,N_7193,N_7463);
xnor U7685 (N_7685,N_7488,N_7467);
or U7686 (N_7686,N_7047,N_7275);
nand U7687 (N_7687,N_7137,N_7411);
nand U7688 (N_7688,N_7344,N_7307);
xor U7689 (N_7689,N_7069,N_7491);
nor U7690 (N_7690,N_7006,N_7230);
xor U7691 (N_7691,N_7172,N_7419);
nand U7692 (N_7692,N_7312,N_7144);
or U7693 (N_7693,N_7248,N_7490);
xnor U7694 (N_7694,N_7418,N_7391);
and U7695 (N_7695,N_7257,N_7205);
xnor U7696 (N_7696,N_7143,N_7139);
and U7697 (N_7697,N_7370,N_7358);
xor U7698 (N_7698,N_7070,N_7018);
nand U7699 (N_7699,N_7425,N_7475);
xor U7700 (N_7700,N_7384,N_7310);
xnor U7701 (N_7701,N_7387,N_7303);
xnor U7702 (N_7702,N_7239,N_7305);
xnor U7703 (N_7703,N_7316,N_7167);
nor U7704 (N_7704,N_7200,N_7092);
nand U7705 (N_7705,N_7499,N_7360);
nor U7706 (N_7706,N_7189,N_7208);
nor U7707 (N_7707,N_7114,N_7314);
and U7708 (N_7708,N_7436,N_7196);
and U7709 (N_7709,N_7123,N_7198);
nand U7710 (N_7710,N_7422,N_7274);
or U7711 (N_7711,N_7207,N_7236);
and U7712 (N_7712,N_7228,N_7443);
and U7713 (N_7713,N_7268,N_7270);
or U7714 (N_7714,N_7004,N_7332);
or U7715 (N_7715,N_7210,N_7431);
nand U7716 (N_7716,N_7277,N_7400);
xnor U7717 (N_7717,N_7299,N_7306);
xor U7718 (N_7718,N_7031,N_7454);
and U7719 (N_7719,N_7175,N_7048);
xor U7720 (N_7720,N_7304,N_7024);
and U7721 (N_7721,N_7097,N_7213);
nor U7722 (N_7722,N_7166,N_7367);
or U7723 (N_7723,N_7075,N_7357);
nand U7724 (N_7724,N_7171,N_7133);
xor U7725 (N_7725,N_7011,N_7076);
nand U7726 (N_7726,N_7083,N_7185);
nor U7727 (N_7727,N_7414,N_7234);
or U7728 (N_7728,N_7102,N_7176);
nand U7729 (N_7729,N_7388,N_7439);
or U7730 (N_7730,N_7046,N_7350);
and U7731 (N_7731,N_7003,N_7250);
nor U7732 (N_7732,N_7156,N_7330);
nand U7733 (N_7733,N_7140,N_7452);
or U7734 (N_7734,N_7432,N_7356);
nand U7735 (N_7735,N_7121,N_7359);
nor U7736 (N_7736,N_7142,N_7470);
and U7737 (N_7737,N_7348,N_7298);
nand U7738 (N_7738,N_7368,N_7108);
or U7739 (N_7739,N_7178,N_7435);
or U7740 (N_7740,N_7186,N_7067);
and U7741 (N_7741,N_7120,N_7119);
and U7742 (N_7742,N_7168,N_7396);
nand U7743 (N_7743,N_7087,N_7088);
and U7744 (N_7744,N_7315,N_7365);
or U7745 (N_7745,N_7240,N_7071);
nand U7746 (N_7746,N_7012,N_7438);
or U7747 (N_7747,N_7086,N_7096);
nor U7748 (N_7748,N_7342,N_7215);
nor U7749 (N_7749,N_7415,N_7326);
and U7750 (N_7750,N_7334,N_7089);
nand U7751 (N_7751,N_7060,N_7103);
nand U7752 (N_7752,N_7359,N_7434);
and U7753 (N_7753,N_7033,N_7332);
nor U7754 (N_7754,N_7323,N_7337);
xor U7755 (N_7755,N_7493,N_7444);
xnor U7756 (N_7756,N_7434,N_7288);
and U7757 (N_7757,N_7207,N_7228);
nand U7758 (N_7758,N_7352,N_7481);
or U7759 (N_7759,N_7046,N_7432);
xor U7760 (N_7760,N_7193,N_7041);
and U7761 (N_7761,N_7492,N_7188);
or U7762 (N_7762,N_7448,N_7065);
nor U7763 (N_7763,N_7449,N_7486);
or U7764 (N_7764,N_7048,N_7165);
or U7765 (N_7765,N_7069,N_7150);
nand U7766 (N_7766,N_7084,N_7409);
xor U7767 (N_7767,N_7447,N_7315);
nor U7768 (N_7768,N_7372,N_7351);
nand U7769 (N_7769,N_7068,N_7410);
or U7770 (N_7770,N_7157,N_7312);
nor U7771 (N_7771,N_7186,N_7465);
nand U7772 (N_7772,N_7275,N_7481);
nand U7773 (N_7773,N_7017,N_7497);
xnor U7774 (N_7774,N_7453,N_7143);
or U7775 (N_7775,N_7165,N_7196);
nor U7776 (N_7776,N_7328,N_7242);
xnor U7777 (N_7777,N_7092,N_7294);
and U7778 (N_7778,N_7153,N_7149);
and U7779 (N_7779,N_7343,N_7192);
or U7780 (N_7780,N_7193,N_7035);
nand U7781 (N_7781,N_7207,N_7441);
or U7782 (N_7782,N_7038,N_7073);
and U7783 (N_7783,N_7085,N_7191);
xnor U7784 (N_7784,N_7075,N_7332);
xnor U7785 (N_7785,N_7292,N_7060);
nor U7786 (N_7786,N_7333,N_7406);
and U7787 (N_7787,N_7355,N_7302);
and U7788 (N_7788,N_7133,N_7226);
xor U7789 (N_7789,N_7284,N_7427);
nand U7790 (N_7790,N_7330,N_7476);
or U7791 (N_7791,N_7343,N_7000);
xor U7792 (N_7792,N_7197,N_7441);
xnor U7793 (N_7793,N_7129,N_7433);
and U7794 (N_7794,N_7102,N_7205);
nand U7795 (N_7795,N_7421,N_7259);
xnor U7796 (N_7796,N_7438,N_7378);
nand U7797 (N_7797,N_7481,N_7412);
nand U7798 (N_7798,N_7102,N_7090);
xor U7799 (N_7799,N_7224,N_7360);
and U7800 (N_7800,N_7018,N_7081);
xor U7801 (N_7801,N_7137,N_7180);
xnor U7802 (N_7802,N_7356,N_7460);
or U7803 (N_7803,N_7038,N_7142);
or U7804 (N_7804,N_7371,N_7309);
or U7805 (N_7805,N_7383,N_7218);
and U7806 (N_7806,N_7028,N_7051);
nor U7807 (N_7807,N_7178,N_7471);
nor U7808 (N_7808,N_7195,N_7300);
nor U7809 (N_7809,N_7488,N_7133);
nor U7810 (N_7810,N_7283,N_7289);
and U7811 (N_7811,N_7131,N_7346);
and U7812 (N_7812,N_7360,N_7265);
xnor U7813 (N_7813,N_7403,N_7015);
xnor U7814 (N_7814,N_7203,N_7058);
nor U7815 (N_7815,N_7261,N_7194);
and U7816 (N_7816,N_7274,N_7127);
xor U7817 (N_7817,N_7099,N_7161);
nor U7818 (N_7818,N_7114,N_7091);
nand U7819 (N_7819,N_7489,N_7281);
nor U7820 (N_7820,N_7013,N_7025);
xnor U7821 (N_7821,N_7479,N_7265);
nand U7822 (N_7822,N_7388,N_7159);
xor U7823 (N_7823,N_7349,N_7087);
nor U7824 (N_7824,N_7178,N_7272);
nor U7825 (N_7825,N_7455,N_7288);
nor U7826 (N_7826,N_7493,N_7253);
xor U7827 (N_7827,N_7122,N_7395);
nor U7828 (N_7828,N_7031,N_7282);
nor U7829 (N_7829,N_7334,N_7121);
xor U7830 (N_7830,N_7256,N_7360);
xnor U7831 (N_7831,N_7231,N_7014);
and U7832 (N_7832,N_7298,N_7300);
nor U7833 (N_7833,N_7235,N_7432);
nor U7834 (N_7834,N_7323,N_7499);
and U7835 (N_7835,N_7234,N_7395);
or U7836 (N_7836,N_7145,N_7358);
or U7837 (N_7837,N_7108,N_7116);
nor U7838 (N_7838,N_7147,N_7425);
nand U7839 (N_7839,N_7238,N_7359);
nor U7840 (N_7840,N_7237,N_7050);
or U7841 (N_7841,N_7358,N_7395);
nor U7842 (N_7842,N_7195,N_7197);
nand U7843 (N_7843,N_7431,N_7258);
or U7844 (N_7844,N_7011,N_7460);
and U7845 (N_7845,N_7295,N_7126);
or U7846 (N_7846,N_7399,N_7303);
xnor U7847 (N_7847,N_7215,N_7107);
and U7848 (N_7848,N_7451,N_7321);
nor U7849 (N_7849,N_7361,N_7122);
nand U7850 (N_7850,N_7022,N_7174);
xor U7851 (N_7851,N_7370,N_7282);
nand U7852 (N_7852,N_7408,N_7114);
xor U7853 (N_7853,N_7112,N_7324);
and U7854 (N_7854,N_7034,N_7062);
nor U7855 (N_7855,N_7277,N_7293);
or U7856 (N_7856,N_7456,N_7197);
xnor U7857 (N_7857,N_7108,N_7138);
xnor U7858 (N_7858,N_7483,N_7063);
nor U7859 (N_7859,N_7099,N_7294);
and U7860 (N_7860,N_7430,N_7310);
nand U7861 (N_7861,N_7221,N_7277);
nor U7862 (N_7862,N_7208,N_7036);
or U7863 (N_7863,N_7220,N_7148);
or U7864 (N_7864,N_7433,N_7486);
or U7865 (N_7865,N_7478,N_7026);
xor U7866 (N_7866,N_7484,N_7384);
or U7867 (N_7867,N_7068,N_7194);
nor U7868 (N_7868,N_7024,N_7277);
nor U7869 (N_7869,N_7426,N_7478);
and U7870 (N_7870,N_7416,N_7297);
and U7871 (N_7871,N_7102,N_7295);
or U7872 (N_7872,N_7206,N_7194);
and U7873 (N_7873,N_7001,N_7262);
and U7874 (N_7874,N_7370,N_7290);
nand U7875 (N_7875,N_7241,N_7191);
or U7876 (N_7876,N_7260,N_7188);
nand U7877 (N_7877,N_7292,N_7057);
and U7878 (N_7878,N_7070,N_7013);
and U7879 (N_7879,N_7437,N_7393);
nor U7880 (N_7880,N_7333,N_7174);
nand U7881 (N_7881,N_7141,N_7102);
and U7882 (N_7882,N_7441,N_7388);
xnor U7883 (N_7883,N_7149,N_7424);
nor U7884 (N_7884,N_7000,N_7155);
nor U7885 (N_7885,N_7361,N_7087);
and U7886 (N_7886,N_7192,N_7160);
xnor U7887 (N_7887,N_7421,N_7233);
xnor U7888 (N_7888,N_7176,N_7492);
and U7889 (N_7889,N_7276,N_7362);
and U7890 (N_7890,N_7036,N_7124);
nand U7891 (N_7891,N_7119,N_7030);
or U7892 (N_7892,N_7219,N_7071);
nand U7893 (N_7893,N_7442,N_7119);
nand U7894 (N_7894,N_7067,N_7291);
nor U7895 (N_7895,N_7470,N_7123);
nor U7896 (N_7896,N_7077,N_7422);
and U7897 (N_7897,N_7265,N_7460);
nand U7898 (N_7898,N_7024,N_7395);
nor U7899 (N_7899,N_7226,N_7108);
nor U7900 (N_7900,N_7024,N_7467);
and U7901 (N_7901,N_7371,N_7216);
and U7902 (N_7902,N_7492,N_7311);
xor U7903 (N_7903,N_7197,N_7328);
xor U7904 (N_7904,N_7443,N_7456);
nand U7905 (N_7905,N_7172,N_7398);
nor U7906 (N_7906,N_7176,N_7126);
or U7907 (N_7907,N_7143,N_7002);
xor U7908 (N_7908,N_7391,N_7218);
nand U7909 (N_7909,N_7369,N_7199);
or U7910 (N_7910,N_7323,N_7157);
xnor U7911 (N_7911,N_7156,N_7241);
nand U7912 (N_7912,N_7499,N_7142);
or U7913 (N_7913,N_7346,N_7231);
xnor U7914 (N_7914,N_7378,N_7436);
xor U7915 (N_7915,N_7475,N_7222);
or U7916 (N_7916,N_7441,N_7093);
nand U7917 (N_7917,N_7403,N_7489);
nand U7918 (N_7918,N_7278,N_7470);
or U7919 (N_7919,N_7254,N_7238);
or U7920 (N_7920,N_7450,N_7098);
nor U7921 (N_7921,N_7146,N_7181);
nor U7922 (N_7922,N_7462,N_7080);
xnor U7923 (N_7923,N_7367,N_7103);
nor U7924 (N_7924,N_7022,N_7146);
xor U7925 (N_7925,N_7006,N_7133);
xnor U7926 (N_7926,N_7214,N_7379);
and U7927 (N_7927,N_7257,N_7361);
xor U7928 (N_7928,N_7223,N_7260);
nor U7929 (N_7929,N_7023,N_7019);
xor U7930 (N_7930,N_7075,N_7497);
nor U7931 (N_7931,N_7397,N_7273);
and U7932 (N_7932,N_7435,N_7337);
and U7933 (N_7933,N_7262,N_7075);
nand U7934 (N_7934,N_7193,N_7482);
xnor U7935 (N_7935,N_7481,N_7058);
nor U7936 (N_7936,N_7472,N_7019);
nor U7937 (N_7937,N_7069,N_7036);
xor U7938 (N_7938,N_7395,N_7321);
and U7939 (N_7939,N_7442,N_7253);
nand U7940 (N_7940,N_7104,N_7003);
or U7941 (N_7941,N_7336,N_7144);
xor U7942 (N_7942,N_7227,N_7446);
or U7943 (N_7943,N_7461,N_7231);
xnor U7944 (N_7944,N_7081,N_7374);
nand U7945 (N_7945,N_7375,N_7111);
or U7946 (N_7946,N_7170,N_7171);
or U7947 (N_7947,N_7421,N_7128);
xnor U7948 (N_7948,N_7234,N_7131);
nor U7949 (N_7949,N_7437,N_7313);
or U7950 (N_7950,N_7357,N_7233);
and U7951 (N_7951,N_7062,N_7312);
xor U7952 (N_7952,N_7098,N_7353);
nand U7953 (N_7953,N_7372,N_7402);
or U7954 (N_7954,N_7135,N_7247);
or U7955 (N_7955,N_7379,N_7171);
nand U7956 (N_7956,N_7001,N_7415);
nand U7957 (N_7957,N_7413,N_7078);
and U7958 (N_7958,N_7120,N_7226);
and U7959 (N_7959,N_7111,N_7155);
xor U7960 (N_7960,N_7474,N_7457);
and U7961 (N_7961,N_7154,N_7464);
or U7962 (N_7962,N_7352,N_7312);
nand U7963 (N_7963,N_7181,N_7092);
or U7964 (N_7964,N_7411,N_7234);
or U7965 (N_7965,N_7125,N_7163);
nor U7966 (N_7966,N_7066,N_7432);
and U7967 (N_7967,N_7279,N_7426);
xnor U7968 (N_7968,N_7172,N_7137);
nand U7969 (N_7969,N_7086,N_7053);
nor U7970 (N_7970,N_7085,N_7354);
xor U7971 (N_7971,N_7167,N_7157);
nor U7972 (N_7972,N_7401,N_7267);
or U7973 (N_7973,N_7133,N_7476);
and U7974 (N_7974,N_7110,N_7231);
xnor U7975 (N_7975,N_7160,N_7396);
nand U7976 (N_7976,N_7023,N_7085);
and U7977 (N_7977,N_7304,N_7103);
nand U7978 (N_7978,N_7322,N_7396);
nor U7979 (N_7979,N_7277,N_7363);
and U7980 (N_7980,N_7489,N_7029);
or U7981 (N_7981,N_7483,N_7461);
nand U7982 (N_7982,N_7024,N_7241);
or U7983 (N_7983,N_7482,N_7347);
xor U7984 (N_7984,N_7245,N_7003);
xnor U7985 (N_7985,N_7448,N_7263);
nor U7986 (N_7986,N_7305,N_7303);
nor U7987 (N_7987,N_7317,N_7109);
xor U7988 (N_7988,N_7472,N_7227);
xnor U7989 (N_7989,N_7292,N_7393);
nor U7990 (N_7990,N_7110,N_7414);
nor U7991 (N_7991,N_7187,N_7130);
nand U7992 (N_7992,N_7353,N_7486);
nand U7993 (N_7993,N_7419,N_7487);
and U7994 (N_7994,N_7446,N_7401);
and U7995 (N_7995,N_7423,N_7131);
or U7996 (N_7996,N_7161,N_7075);
and U7997 (N_7997,N_7008,N_7027);
xor U7998 (N_7998,N_7239,N_7479);
or U7999 (N_7999,N_7234,N_7032);
nor U8000 (N_8000,N_7868,N_7581);
and U8001 (N_8001,N_7820,N_7779);
nor U8002 (N_8002,N_7613,N_7508);
nor U8003 (N_8003,N_7662,N_7735);
nor U8004 (N_8004,N_7853,N_7684);
or U8005 (N_8005,N_7722,N_7993);
and U8006 (N_8006,N_7915,N_7783);
nand U8007 (N_8007,N_7583,N_7523);
nor U8008 (N_8008,N_7616,N_7884);
nor U8009 (N_8009,N_7949,N_7622);
xor U8010 (N_8010,N_7894,N_7510);
nor U8011 (N_8011,N_7888,N_7570);
and U8012 (N_8012,N_7543,N_7528);
nor U8013 (N_8013,N_7869,N_7708);
xnor U8014 (N_8014,N_7924,N_7585);
xor U8015 (N_8015,N_7716,N_7749);
xor U8016 (N_8016,N_7969,N_7787);
nand U8017 (N_8017,N_7878,N_7641);
nand U8018 (N_8018,N_7950,N_7589);
or U8019 (N_8019,N_7947,N_7805);
and U8020 (N_8020,N_7914,N_7707);
or U8021 (N_8021,N_7815,N_7940);
nor U8022 (N_8022,N_7745,N_7923);
or U8023 (N_8023,N_7865,N_7800);
and U8024 (N_8024,N_7590,N_7657);
or U8025 (N_8025,N_7951,N_7864);
and U8026 (N_8026,N_7833,N_7655);
and U8027 (N_8027,N_7956,N_7531);
and U8028 (N_8028,N_7834,N_7999);
nand U8029 (N_8029,N_7628,N_7670);
nand U8030 (N_8030,N_7534,N_7921);
nand U8031 (N_8031,N_7627,N_7652);
xor U8032 (N_8032,N_7984,N_7677);
xnor U8033 (N_8033,N_7596,N_7535);
nand U8034 (N_8034,N_7636,N_7825);
nand U8035 (N_8035,N_7811,N_7766);
nand U8036 (N_8036,N_7690,N_7858);
nand U8037 (N_8037,N_7780,N_7651);
nor U8038 (N_8038,N_7633,N_7674);
nor U8039 (N_8039,N_7901,N_7598);
nand U8040 (N_8040,N_7866,N_7946);
or U8041 (N_8041,N_7703,N_7850);
and U8042 (N_8042,N_7506,N_7697);
or U8043 (N_8043,N_7916,N_7611);
nor U8044 (N_8044,N_7908,N_7597);
nand U8045 (N_8045,N_7863,N_7660);
nand U8046 (N_8046,N_7848,N_7656);
and U8047 (N_8047,N_7985,N_7930);
nor U8048 (N_8048,N_7742,N_7675);
and U8049 (N_8049,N_7927,N_7764);
or U8050 (N_8050,N_7577,N_7812);
xor U8051 (N_8051,N_7673,N_7553);
xnor U8052 (N_8052,N_7977,N_7773);
nand U8053 (N_8053,N_7502,N_7718);
nand U8054 (N_8054,N_7905,N_7887);
xor U8055 (N_8055,N_7644,N_7859);
or U8056 (N_8056,N_7992,N_7883);
nand U8057 (N_8057,N_7810,N_7939);
xnor U8058 (N_8058,N_7560,N_7608);
or U8059 (N_8059,N_7897,N_7918);
nor U8060 (N_8060,N_7711,N_7807);
nand U8061 (N_8061,N_7668,N_7587);
nor U8062 (N_8062,N_7871,N_7595);
xnor U8063 (N_8063,N_7981,N_7913);
nand U8064 (N_8064,N_7898,N_7952);
nand U8065 (N_8065,N_7639,N_7503);
nand U8066 (N_8066,N_7614,N_7998);
nor U8067 (N_8067,N_7731,N_7775);
and U8068 (N_8068,N_7615,N_7704);
or U8069 (N_8069,N_7791,N_7530);
nand U8070 (N_8070,N_7556,N_7709);
xnor U8071 (N_8071,N_7693,N_7756);
nand U8072 (N_8072,N_7664,N_7857);
nand U8073 (N_8073,N_7837,N_7720);
and U8074 (N_8074,N_7944,N_7514);
or U8075 (N_8075,N_7903,N_7907);
or U8076 (N_8076,N_7607,N_7686);
nor U8077 (N_8077,N_7527,N_7753);
nand U8078 (N_8078,N_7774,N_7654);
and U8079 (N_8079,N_7743,N_7542);
nor U8080 (N_8080,N_7824,N_7919);
or U8081 (N_8081,N_7715,N_7612);
or U8082 (N_8082,N_7885,N_7519);
nand U8083 (N_8083,N_7769,N_7548);
or U8084 (N_8084,N_7804,N_7705);
and U8085 (N_8085,N_7537,N_7699);
or U8086 (N_8086,N_7814,N_7591);
or U8087 (N_8087,N_7550,N_7700);
xnor U8088 (N_8088,N_7602,N_7971);
xnor U8089 (N_8089,N_7911,N_7909);
or U8090 (N_8090,N_7593,N_7557);
nand U8091 (N_8091,N_7549,N_7555);
xor U8092 (N_8092,N_7562,N_7788);
or U8093 (N_8093,N_7594,N_7852);
or U8094 (N_8094,N_7520,N_7855);
xnor U8095 (N_8095,N_7563,N_7890);
nor U8096 (N_8096,N_7521,N_7782);
nand U8097 (N_8097,N_7565,N_7757);
nor U8098 (N_8098,N_7659,N_7667);
or U8099 (N_8099,N_7736,N_7566);
nand U8100 (N_8100,N_7806,N_7879);
nor U8101 (N_8101,N_7712,N_7649);
and U8102 (N_8102,N_7663,N_7640);
nor U8103 (N_8103,N_7685,N_7819);
xnor U8104 (N_8104,N_7672,N_7854);
xnor U8105 (N_8105,N_7632,N_7610);
or U8106 (N_8106,N_7547,N_7576);
xor U8107 (N_8107,N_7706,N_7873);
or U8108 (N_8108,N_7741,N_7948);
xnor U8109 (N_8109,N_7793,N_7678);
xnor U8110 (N_8110,N_7899,N_7943);
or U8111 (N_8111,N_7803,N_7676);
and U8112 (N_8112,N_7822,N_7790);
xnor U8113 (N_8113,N_7737,N_7872);
xor U8114 (N_8114,N_7891,N_7532);
and U8115 (N_8115,N_7974,N_7669);
and U8116 (N_8116,N_7986,N_7829);
nor U8117 (N_8117,N_7605,N_7701);
xor U8118 (N_8118,N_7637,N_7955);
nor U8119 (N_8119,N_7768,N_7840);
or U8120 (N_8120,N_7642,N_7511);
xnor U8121 (N_8121,N_7661,N_7798);
xor U8122 (N_8122,N_7895,N_7875);
xnor U8123 (N_8123,N_7926,N_7692);
and U8124 (N_8124,N_7893,N_7823);
and U8125 (N_8125,N_7759,N_7827);
xnor U8126 (N_8126,N_7934,N_7846);
nand U8127 (N_8127,N_7710,N_7630);
and U8128 (N_8128,N_7845,N_7931);
xnor U8129 (N_8129,N_7726,N_7889);
and U8130 (N_8130,N_7922,N_7896);
or U8131 (N_8131,N_7938,N_7746);
and U8132 (N_8132,N_7729,N_7925);
or U8133 (N_8133,N_7886,N_7658);
xor U8134 (N_8134,N_7601,N_7509);
or U8135 (N_8135,N_7634,N_7933);
or U8136 (N_8136,N_7569,N_7653);
nor U8137 (N_8137,N_7995,N_7683);
xnor U8138 (N_8138,N_7802,N_7817);
xnor U8139 (N_8139,N_7963,N_7540);
nand U8140 (N_8140,N_7648,N_7580);
and U8141 (N_8141,N_7781,N_7862);
nor U8142 (N_8142,N_7629,N_7968);
xnor U8143 (N_8143,N_7723,N_7545);
xnor U8144 (N_8144,N_7504,N_7973);
nand U8145 (N_8145,N_7599,N_7906);
xor U8146 (N_8146,N_7719,N_7754);
xnor U8147 (N_8147,N_7721,N_7785);
or U8148 (N_8148,N_7513,N_7572);
xor U8149 (N_8149,N_7734,N_7606);
or U8150 (N_8150,N_7750,N_7839);
nor U8151 (N_8151,N_7600,N_7573);
or U8152 (N_8152,N_7799,N_7989);
nand U8153 (N_8153,N_7784,N_7727);
or U8154 (N_8154,N_7529,N_7567);
nor U8155 (N_8155,N_7541,N_7500);
nand U8156 (N_8156,N_7979,N_7588);
xnor U8157 (N_8157,N_7836,N_7920);
nor U8158 (N_8158,N_7666,N_7941);
nor U8159 (N_8159,N_7844,N_7816);
or U8160 (N_8160,N_7501,N_7945);
nand U8161 (N_8161,N_7776,N_7713);
or U8162 (N_8162,N_7524,N_7828);
and U8163 (N_8163,N_7631,N_7794);
nand U8164 (N_8164,N_7620,N_7904);
or U8165 (N_8165,N_7942,N_7847);
or U8166 (N_8166,N_7702,N_7730);
and U8167 (N_8167,N_7809,N_7752);
or U8168 (N_8168,N_7582,N_7961);
nand U8169 (N_8169,N_7801,N_7980);
nor U8170 (N_8170,N_7767,N_7619);
xor U8171 (N_8171,N_7571,N_7770);
nor U8172 (N_8172,N_7957,N_7763);
nor U8173 (N_8173,N_7876,N_7518);
nor U8174 (N_8174,N_7808,N_7987);
and U8175 (N_8175,N_7551,N_7517);
xor U8176 (N_8176,N_7691,N_7990);
or U8177 (N_8177,N_7680,N_7882);
or U8178 (N_8178,N_7625,N_7533);
nand U8179 (N_8179,N_7579,N_7826);
nand U8180 (N_8180,N_7643,N_7843);
and U8181 (N_8181,N_7953,N_7965);
nor U8182 (N_8182,N_7835,N_7512);
and U8183 (N_8183,N_7813,N_7976);
or U8184 (N_8184,N_7967,N_7983);
and U8185 (N_8185,N_7525,N_7621);
and U8186 (N_8186,N_7856,N_7758);
nor U8187 (N_8187,N_7958,N_7574);
xnor U8188 (N_8188,N_7860,N_7842);
or U8189 (N_8189,N_7698,N_7789);
xnor U8190 (N_8190,N_7538,N_7851);
xnor U8191 (N_8191,N_7717,N_7917);
nand U8192 (N_8192,N_7740,N_7568);
nor U8193 (N_8193,N_7765,N_7892);
and U8194 (N_8194,N_7539,N_7994);
or U8195 (N_8195,N_7910,N_7978);
and U8196 (N_8196,N_7755,N_7818);
or U8197 (N_8197,N_7912,N_7877);
or U8198 (N_8198,N_7578,N_7624);
or U8199 (N_8199,N_7584,N_7623);
or U8200 (N_8200,N_7728,N_7617);
xor U8201 (N_8201,N_7515,N_7797);
nor U8202 (N_8202,N_7650,N_7902);
or U8203 (N_8203,N_7960,N_7559);
xor U8204 (N_8204,N_7645,N_7694);
nor U8205 (N_8205,N_7618,N_7744);
xor U8206 (N_8206,N_7867,N_7786);
and U8207 (N_8207,N_7575,N_7687);
and U8208 (N_8208,N_7936,N_7609);
nand U8209 (N_8209,N_7841,N_7696);
and U8210 (N_8210,N_7688,N_7558);
xor U8211 (N_8211,N_7733,N_7880);
nand U8212 (N_8212,N_7964,N_7962);
or U8213 (N_8213,N_7937,N_7870);
nand U8214 (N_8214,N_7772,N_7982);
xor U8215 (N_8215,N_7536,N_7725);
nand U8216 (N_8216,N_7954,N_7522);
or U8217 (N_8217,N_7997,N_7795);
xnor U8218 (N_8218,N_7586,N_7671);
nand U8219 (N_8219,N_7592,N_7505);
nand U8220 (N_8220,N_7679,N_7552);
xor U8221 (N_8221,N_7972,N_7830);
xnor U8222 (N_8222,N_7832,N_7747);
or U8223 (N_8223,N_7544,N_7991);
or U8224 (N_8224,N_7739,N_7681);
and U8225 (N_8225,N_7738,N_7821);
xnor U8226 (N_8226,N_7646,N_7626);
and U8227 (N_8227,N_7647,N_7604);
nand U8228 (N_8228,N_7665,N_7561);
and U8229 (N_8229,N_7777,N_7849);
nand U8230 (N_8230,N_7861,N_7516);
xnor U8231 (N_8231,N_7996,N_7732);
or U8232 (N_8232,N_7874,N_7751);
xor U8233 (N_8233,N_7792,N_7970);
nor U8234 (N_8234,N_7762,N_7831);
nand U8235 (N_8235,N_7959,N_7881);
xnor U8236 (N_8236,N_7682,N_7975);
or U8237 (N_8237,N_7603,N_7761);
or U8238 (N_8238,N_7724,N_7778);
and U8239 (N_8239,N_7935,N_7929);
nand U8240 (N_8240,N_7966,N_7760);
nand U8241 (N_8241,N_7564,N_7771);
nor U8242 (N_8242,N_7900,N_7638);
xnor U8243 (N_8243,N_7748,N_7507);
nor U8244 (N_8244,N_7988,N_7546);
and U8245 (N_8245,N_7554,N_7635);
nor U8246 (N_8246,N_7838,N_7714);
or U8247 (N_8247,N_7695,N_7796);
or U8248 (N_8248,N_7689,N_7928);
xnor U8249 (N_8249,N_7932,N_7526);
nor U8250 (N_8250,N_7817,N_7661);
nor U8251 (N_8251,N_7856,N_7650);
nand U8252 (N_8252,N_7899,N_7879);
nor U8253 (N_8253,N_7654,N_7867);
xnor U8254 (N_8254,N_7562,N_7620);
xor U8255 (N_8255,N_7928,N_7548);
and U8256 (N_8256,N_7636,N_7514);
or U8257 (N_8257,N_7734,N_7743);
nand U8258 (N_8258,N_7585,N_7564);
or U8259 (N_8259,N_7996,N_7520);
nand U8260 (N_8260,N_7768,N_7612);
nand U8261 (N_8261,N_7635,N_7686);
nor U8262 (N_8262,N_7673,N_7937);
nor U8263 (N_8263,N_7821,N_7829);
or U8264 (N_8264,N_7763,N_7797);
xnor U8265 (N_8265,N_7674,N_7612);
and U8266 (N_8266,N_7736,N_7607);
or U8267 (N_8267,N_7769,N_7970);
nand U8268 (N_8268,N_7739,N_7902);
and U8269 (N_8269,N_7987,N_7835);
xnor U8270 (N_8270,N_7531,N_7675);
or U8271 (N_8271,N_7797,N_7943);
nand U8272 (N_8272,N_7775,N_7924);
nor U8273 (N_8273,N_7659,N_7902);
or U8274 (N_8274,N_7810,N_7911);
and U8275 (N_8275,N_7773,N_7519);
and U8276 (N_8276,N_7832,N_7739);
xor U8277 (N_8277,N_7636,N_7854);
nor U8278 (N_8278,N_7842,N_7963);
nor U8279 (N_8279,N_7615,N_7788);
and U8280 (N_8280,N_7577,N_7842);
or U8281 (N_8281,N_7920,N_7714);
and U8282 (N_8282,N_7613,N_7734);
and U8283 (N_8283,N_7577,N_7748);
and U8284 (N_8284,N_7592,N_7772);
or U8285 (N_8285,N_7990,N_7736);
nand U8286 (N_8286,N_7773,N_7941);
and U8287 (N_8287,N_7542,N_7809);
nor U8288 (N_8288,N_7663,N_7800);
or U8289 (N_8289,N_7625,N_7500);
xnor U8290 (N_8290,N_7862,N_7954);
xnor U8291 (N_8291,N_7827,N_7547);
nand U8292 (N_8292,N_7679,N_7723);
nor U8293 (N_8293,N_7685,N_7641);
and U8294 (N_8294,N_7551,N_7950);
nand U8295 (N_8295,N_7564,N_7503);
and U8296 (N_8296,N_7902,N_7622);
xor U8297 (N_8297,N_7503,N_7657);
xor U8298 (N_8298,N_7978,N_7633);
and U8299 (N_8299,N_7941,N_7989);
or U8300 (N_8300,N_7565,N_7877);
nor U8301 (N_8301,N_7656,N_7728);
xnor U8302 (N_8302,N_7664,N_7601);
or U8303 (N_8303,N_7719,N_7758);
xnor U8304 (N_8304,N_7670,N_7608);
xor U8305 (N_8305,N_7788,N_7851);
nor U8306 (N_8306,N_7540,N_7659);
xnor U8307 (N_8307,N_7769,N_7977);
nand U8308 (N_8308,N_7590,N_7814);
nand U8309 (N_8309,N_7758,N_7756);
and U8310 (N_8310,N_7771,N_7632);
xnor U8311 (N_8311,N_7709,N_7531);
or U8312 (N_8312,N_7669,N_7910);
nor U8313 (N_8313,N_7961,N_7694);
and U8314 (N_8314,N_7788,N_7722);
nand U8315 (N_8315,N_7752,N_7625);
nand U8316 (N_8316,N_7886,N_7924);
or U8317 (N_8317,N_7719,N_7685);
and U8318 (N_8318,N_7735,N_7917);
or U8319 (N_8319,N_7715,N_7927);
nor U8320 (N_8320,N_7785,N_7833);
or U8321 (N_8321,N_7761,N_7891);
xor U8322 (N_8322,N_7945,N_7803);
or U8323 (N_8323,N_7630,N_7588);
nand U8324 (N_8324,N_7622,N_7704);
nand U8325 (N_8325,N_7737,N_7823);
nand U8326 (N_8326,N_7706,N_7626);
nor U8327 (N_8327,N_7972,N_7994);
nand U8328 (N_8328,N_7552,N_7882);
xor U8329 (N_8329,N_7992,N_7731);
xor U8330 (N_8330,N_7814,N_7662);
or U8331 (N_8331,N_7530,N_7660);
nand U8332 (N_8332,N_7680,N_7919);
or U8333 (N_8333,N_7946,N_7611);
xnor U8334 (N_8334,N_7607,N_7956);
and U8335 (N_8335,N_7896,N_7733);
or U8336 (N_8336,N_7793,N_7737);
or U8337 (N_8337,N_7881,N_7875);
nand U8338 (N_8338,N_7842,N_7665);
nor U8339 (N_8339,N_7837,N_7706);
or U8340 (N_8340,N_7628,N_7895);
nor U8341 (N_8341,N_7991,N_7951);
xnor U8342 (N_8342,N_7535,N_7522);
nor U8343 (N_8343,N_7843,N_7505);
nand U8344 (N_8344,N_7654,N_7558);
nand U8345 (N_8345,N_7888,N_7945);
xor U8346 (N_8346,N_7987,N_7798);
xor U8347 (N_8347,N_7935,N_7628);
nor U8348 (N_8348,N_7883,N_7781);
nor U8349 (N_8349,N_7530,N_7648);
or U8350 (N_8350,N_7704,N_7739);
nand U8351 (N_8351,N_7665,N_7752);
or U8352 (N_8352,N_7734,N_7989);
or U8353 (N_8353,N_7631,N_7900);
xor U8354 (N_8354,N_7987,N_7733);
nor U8355 (N_8355,N_7581,N_7690);
and U8356 (N_8356,N_7575,N_7617);
xor U8357 (N_8357,N_7877,N_7786);
nor U8358 (N_8358,N_7894,N_7648);
nor U8359 (N_8359,N_7762,N_7858);
xor U8360 (N_8360,N_7885,N_7740);
xor U8361 (N_8361,N_7857,N_7859);
and U8362 (N_8362,N_7782,N_7607);
nor U8363 (N_8363,N_7949,N_7690);
or U8364 (N_8364,N_7733,N_7990);
and U8365 (N_8365,N_7959,N_7617);
xor U8366 (N_8366,N_7687,N_7896);
and U8367 (N_8367,N_7742,N_7924);
xnor U8368 (N_8368,N_7948,N_7996);
nand U8369 (N_8369,N_7623,N_7522);
or U8370 (N_8370,N_7899,N_7693);
nand U8371 (N_8371,N_7573,N_7585);
or U8372 (N_8372,N_7665,N_7632);
nor U8373 (N_8373,N_7723,N_7765);
xor U8374 (N_8374,N_7708,N_7607);
nand U8375 (N_8375,N_7717,N_7733);
nand U8376 (N_8376,N_7758,N_7790);
and U8377 (N_8377,N_7743,N_7732);
or U8378 (N_8378,N_7622,N_7731);
nand U8379 (N_8379,N_7650,N_7857);
nand U8380 (N_8380,N_7564,N_7799);
or U8381 (N_8381,N_7871,N_7949);
xnor U8382 (N_8382,N_7722,N_7557);
or U8383 (N_8383,N_7512,N_7845);
and U8384 (N_8384,N_7742,N_7662);
nand U8385 (N_8385,N_7884,N_7691);
nor U8386 (N_8386,N_7614,N_7967);
nand U8387 (N_8387,N_7929,N_7908);
and U8388 (N_8388,N_7826,N_7633);
or U8389 (N_8389,N_7728,N_7624);
and U8390 (N_8390,N_7817,N_7515);
and U8391 (N_8391,N_7800,N_7501);
xor U8392 (N_8392,N_7801,N_7889);
nor U8393 (N_8393,N_7686,N_7563);
and U8394 (N_8394,N_7971,N_7937);
nand U8395 (N_8395,N_7987,N_7601);
or U8396 (N_8396,N_7757,N_7726);
or U8397 (N_8397,N_7650,N_7658);
or U8398 (N_8398,N_7550,N_7871);
or U8399 (N_8399,N_7867,N_7895);
or U8400 (N_8400,N_7723,N_7707);
or U8401 (N_8401,N_7675,N_7810);
and U8402 (N_8402,N_7902,N_7874);
nand U8403 (N_8403,N_7668,N_7601);
nand U8404 (N_8404,N_7929,N_7911);
and U8405 (N_8405,N_7816,N_7736);
or U8406 (N_8406,N_7829,N_7533);
or U8407 (N_8407,N_7746,N_7970);
and U8408 (N_8408,N_7720,N_7854);
or U8409 (N_8409,N_7979,N_7929);
and U8410 (N_8410,N_7961,N_7873);
and U8411 (N_8411,N_7992,N_7712);
or U8412 (N_8412,N_7939,N_7713);
nand U8413 (N_8413,N_7976,N_7511);
or U8414 (N_8414,N_7763,N_7905);
xnor U8415 (N_8415,N_7522,N_7984);
xor U8416 (N_8416,N_7619,N_7749);
or U8417 (N_8417,N_7978,N_7926);
or U8418 (N_8418,N_7858,N_7952);
and U8419 (N_8419,N_7638,N_7951);
and U8420 (N_8420,N_7749,N_7656);
or U8421 (N_8421,N_7584,N_7610);
nor U8422 (N_8422,N_7542,N_7849);
or U8423 (N_8423,N_7558,N_7766);
nand U8424 (N_8424,N_7969,N_7603);
xor U8425 (N_8425,N_7542,N_7825);
xnor U8426 (N_8426,N_7747,N_7876);
nor U8427 (N_8427,N_7770,N_7968);
or U8428 (N_8428,N_7764,N_7932);
xnor U8429 (N_8429,N_7847,N_7810);
or U8430 (N_8430,N_7639,N_7923);
and U8431 (N_8431,N_7969,N_7970);
nor U8432 (N_8432,N_7598,N_7640);
nor U8433 (N_8433,N_7627,N_7681);
nor U8434 (N_8434,N_7608,N_7760);
or U8435 (N_8435,N_7865,N_7756);
and U8436 (N_8436,N_7995,N_7938);
or U8437 (N_8437,N_7571,N_7745);
nand U8438 (N_8438,N_7864,N_7677);
or U8439 (N_8439,N_7671,N_7530);
and U8440 (N_8440,N_7660,N_7982);
or U8441 (N_8441,N_7898,N_7951);
or U8442 (N_8442,N_7670,N_7740);
or U8443 (N_8443,N_7631,N_7753);
nand U8444 (N_8444,N_7821,N_7783);
or U8445 (N_8445,N_7940,N_7894);
nor U8446 (N_8446,N_7786,N_7767);
nand U8447 (N_8447,N_7934,N_7502);
and U8448 (N_8448,N_7693,N_7906);
or U8449 (N_8449,N_7547,N_7645);
nor U8450 (N_8450,N_7663,N_7677);
nor U8451 (N_8451,N_7675,N_7636);
and U8452 (N_8452,N_7702,N_7778);
and U8453 (N_8453,N_7957,N_7809);
and U8454 (N_8454,N_7817,N_7650);
xor U8455 (N_8455,N_7978,N_7562);
or U8456 (N_8456,N_7903,N_7926);
nand U8457 (N_8457,N_7914,N_7553);
nor U8458 (N_8458,N_7704,N_7649);
and U8459 (N_8459,N_7856,N_7546);
nor U8460 (N_8460,N_7727,N_7944);
or U8461 (N_8461,N_7808,N_7726);
nor U8462 (N_8462,N_7517,N_7667);
or U8463 (N_8463,N_7639,N_7513);
nor U8464 (N_8464,N_7935,N_7549);
xor U8465 (N_8465,N_7540,N_7563);
nand U8466 (N_8466,N_7731,N_7515);
nor U8467 (N_8467,N_7703,N_7960);
nor U8468 (N_8468,N_7836,N_7752);
xor U8469 (N_8469,N_7597,N_7575);
nand U8470 (N_8470,N_7740,N_7891);
nor U8471 (N_8471,N_7640,N_7696);
xor U8472 (N_8472,N_7806,N_7781);
and U8473 (N_8473,N_7798,N_7597);
nor U8474 (N_8474,N_7975,N_7915);
nor U8475 (N_8475,N_7620,N_7969);
nor U8476 (N_8476,N_7955,N_7694);
nor U8477 (N_8477,N_7761,N_7692);
and U8478 (N_8478,N_7544,N_7524);
or U8479 (N_8479,N_7854,N_7773);
and U8480 (N_8480,N_7958,N_7770);
and U8481 (N_8481,N_7635,N_7789);
nand U8482 (N_8482,N_7516,N_7806);
nand U8483 (N_8483,N_7867,N_7595);
and U8484 (N_8484,N_7523,N_7872);
and U8485 (N_8485,N_7602,N_7613);
nor U8486 (N_8486,N_7659,N_7919);
nor U8487 (N_8487,N_7699,N_7645);
nand U8488 (N_8488,N_7724,N_7625);
or U8489 (N_8489,N_7846,N_7795);
or U8490 (N_8490,N_7862,N_7901);
and U8491 (N_8491,N_7729,N_7638);
and U8492 (N_8492,N_7922,N_7732);
nor U8493 (N_8493,N_7978,N_7572);
nor U8494 (N_8494,N_7901,N_7816);
xor U8495 (N_8495,N_7607,N_7556);
and U8496 (N_8496,N_7950,N_7768);
and U8497 (N_8497,N_7962,N_7895);
xor U8498 (N_8498,N_7909,N_7832);
or U8499 (N_8499,N_7580,N_7834);
nor U8500 (N_8500,N_8073,N_8063);
nor U8501 (N_8501,N_8112,N_8438);
and U8502 (N_8502,N_8052,N_8211);
nand U8503 (N_8503,N_8371,N_8119);
nor U8504 (N_8504,N_8009,N_8306);
xnor U8505 (N_8505,N_8396,N_8417);
nand U8506 (N_8506,N_8373,N_8414);
nor U8507 (N_8507,N_8334,N_8226);
nand U8508 (N_8508,N_8499,N_8083);
nor U8509 (N_8509,N_8198,N_8014);
nand U8510 (N_8510,N_8240,N_8419);
xnor U8511 (N_8511,N_8107,N_8383);
nand U8512 (N_8512,N_8129,N_8425);
and U8513 (N_8513,N_8208,N_8053);
or U8514 (N_8514,N_8397,N_8166);
xnor U8515 (N_8515,N_8159,N_8313);
and U8516 (N_8516,N_8303,N_8487);
xor U8517 (N_8517,N_8199,N_8249);
nor U8518 (N_8518,N_8061,N_8104);
and U8519 (N_8519,N_8393,N_8262);
nor U8520 (N_8520,N_8178,N_8343);
and U8521 (N_8521,N_8344,N_8265);
and U8522 (N_8522,N_8153,N_8094);
nand U8523 (N_8523,N_8224,N_8082);
nand U8524 (N_8524,N_8353,N_8422);
and U8525 (N_8525,N_8118,N_8215);
xor U8526 (N_8526,N_8269,N_8151);
nand U8527 (N_8527,N_8367,N_8426);
or U8528 (N_8528,N_8455,N_8449);
nand U8529 (N_8529,N_8429,N_8365);
and U8530 (N_8530,N_8287,N_8039);
or U8531 (N_8531,N_8250,N_8185);
nor U8532 (N_8532,N_8321,N_8044);
nor U8533 (N_8533,N_8395,N_8441);
xnor U8534 (N_8534,N_8236,N_8304);
xor U8535 (N_8535,N_8464,N_8123);
and U8536 (N_8536,N_8225,N_8368);
and U8537 (N_8537,N_8292,N_8331);
nand U8538 (N_8538,N_8244,N_8184);
xor U8539 (N_8539,N_8217,N_8146);
or U8540 (N_8540,N_8308,N_8381);
and U8541 (N_8541,N_8357,N_8366);
and U8542 (N_8542,N_8372,N_8227);
xor U8543 (N_8543,N_8204,N_8348);
or U8544 (N_8544,N_8088,N_8207);
nor U8545 (N_8545,N_8336,N_8272);
or U8546 (N_8546,N_8124,N_8318);
and U8547 (N_8547,N_8162,N_8320);
nor U8548 (N_8548,N_8132,N_8314);
and U8549 (N_8549,N_8447,N_8209);
nand U8550 (N_8550,N_8310,N_8275);
nand U8551 (N_8551,N_8143,N_8278);
nand U8552 (N_8552,N_8445,N_8004);
nand U8553 (N_8553,N_8350,N_8477);
xnor U8554 (N_8554,N_8280,N_8347);
nor U8555 (N_8555,N_8183,N_8223);
nor U8556 (N_8556,N_8399,N_8327);
xor U8557 (N_8557,N_8376,N_8408);
or U8558 (N_8558,N_8089,N_8205);
xor U8559 (N_8559,N_8027,N_8488);
or U8560 (N_8560,N_8048,N_8420);
or U8561 (N_8561,N_8403,N_8261);
xnor U8562 (N_8562,N_8322,N_8147);
or U8563 (N_8563,N_8005,N_8152);
nor U8564 (N_8564,N_8160,N_8058);
nor U8565 (N_8565,N_8260,N_8349);
xor U8566 (N_8566,N_8043,N_8405);
xnor U8567 (N_8567,N_8157,N_8354);
or U8568 (N_8568,N_8181,N_8358);
nand U8569 (N_8569,N_8079,N_8382);
nor U8570 (N_8570,N_8241,N_8302);
or U8571 (N_8571,N_8125,N_8268);
nor U8572 (N_8572,N_8050,N_8461);
and U8573 (N_8573,N_8046,N_8497);
nor U8574 (N_8574,N_8006,N_8406);
nor U8575 (N_8575,N_8099,N_8361);
or U8576 (N_8576,N_8378,N_8440);
and U8577 (N_8577,N_8072,N_8093);
and U8578 (N_8578,N_8410,N_8324);
or U8579 (N_8579,N_8047,N_8271);
and U8580 (N_8580,N_8214,N_8003);
nor U8581 (N_8581,N_8297,N_8456);
nor U8582 (N_8582,N_8284,N_8270);
or U8583 (N_8583,N_8114,N_8404);
nand U8584 (N_8584,N_8031,N_8484);
nor U8585 (N_8585,N_8154,N_8174);
and U8586 (N_8586,N_8051,N_8385);
nor U8587 (N_8587,N_8036,N_8128);
or U8588 (N_8588,N_8235,N_8098);
xor U8589 (N_8589,N_8078,N_8409);
nand U8590 (N_8590,N_8283,N_8307);
or U8591 (N_8591,N_8282,N_8387);
nor U8592 (N_8592,N_8010,N_8281);
nand U8593 (N_8593,N_8191,N_8359);
and U8594 (N_8594,N_8253,N_8309);
nand U8595 (N_8595,N_8126,N_8168);
or U8596 (N_8596,N_8312,N_8264);
or U8597 (N_8597,N_8013,N_8459);
xnor U8598 (N_8598,N_8109,N_8345);
xor U8599 (N_8599,N_8401,N_8092);
xnor U8600 (N_8600,N_8000,N_8033);
nand U8601 (N_8601,N_8479,N_8351);
or U8602 (N_8602,N_8362,N_8469);
and U8603 (N_8603,N_8494,N_8220);
nand U8604 (N_8604,N_8038,N_8242);
xor U8605 (N_8605,N_8352,N_8444);
and U8606 (N_8606,N_8175,N_8407);
nor U8607 (N_8607,N_8356,N_8196);
and U8608 (N_8608,N_8374,N_8020);
or U8609 (N_8609,N_8096,N_8090);
and U8610 (N_8610,N_8173,N_8001);
nor U8611 (N_8611,N_8413,N_8187);
and U8612 (N_8612,N_8086,N_8256);
xnor U8613 (N_8613,N_8077,N_8498);
xnor U8614 (N_8614,N_8130,N_8024);
and U8615 (N_8615,N_8193,N_8450);
nor U8616 (N_8616,N_8491,N_8221);
or U8617 (N_8617,N_8301,N_8218);
nor U8618 (N_8618,N_8156,N_8267);
and U8619 (N_8619,N_8337,N_8040);
and U8620 (N_8620,N_8433,N_8200);
nor U8621 (N_8621,N_8120,N_8172);
and U8622 (N_8622,N_8462,N_8330);
nor U8623 (N_8623,N_8482,N_8192);
xnor U8624 (N_8624,N_8285,N_8471);
nand U8625 (N_8625,N_8025,N_8219);
xor U8626 (N_8626,N_8239,N_8189);
nor U8627 (N_8627,N_8231,N_8016);
nor U8628 (N_8628,N_8180,N_8234);
xnor U8629 (N_8629,N_8169,N_8255);
and U8630 (N_8630,N_8338,N_8190);
nand U8631 (N_8631,N_8305,N_8364);
nand U8632 (N_8632,N_8070,N_8045);
nor U8633 (N_8633,N_8391,N_8300);
and U8634 (N_8634,N_8465,N_8206);
nor U8635 (N_8635,N_8369,N_8415);
xnor U8636 (N_8636,N_8424,N_8476);
nand U8637 (N_8637,N_8329,N_8377);
nand U8638 (N_8638,N_8472,N_8158);
nand U8639 (N_8639,N_8493,N_8186);
nand U8640 (N_8640,N_8167,N_8478);
nor U8641 (N_8641,N_8274,N_8229);
nor U8642 (N_8642,N_8467,N_8103);
nor U8643 (N_8643,N_8384,N_8064);
and U8644 (N_8644,N_8238,N_8097);
and U8645 (N_8645,N_8121,N_8485);
nand U8646 (N_8646,N_8028,N_8188);
or U8647 (N_8647,N_8150,N_8115);
or U8648 (N_8648,N_8427,N_8116);
xor U8649 (N_8649,N_8339,N_8490);
nand U8650 (N_8650,N_8195,N_8007);
nor U8651 (N_8651,N_8210,N_8473);
and U8652 (N_8652,N_8202,N_8454);
nor U8653 (N_8653,N_8248,N_8237);
and U8654 (N_8654,N_8435,N_8108);
xnor U8655 (N_8655,N_8288,N_8134);
or U8656 (N_8656,N_8428,N_8182);
or U8657 (N_8657,N_8138,N_8144);
and U8658 (N_8658,N_8436,N_8453);
nor U8659 (N_8659,N_8294,N_8468);
and U8660 (N_8660,N_8136,N_8439);
xnor U8661 (N_8661,N_8075,N_8122);
nor U8662 (N_8662,N_8149,N_8049);
and U8663 (N_8663,N_8342,N_8475);
nand U8664 (N_8664,N_8355,N_8480);
or U8665 (N_8665,N_8370,N_8483);
nor U8666 (N_8666,N_8141,N_8111);
and U8667 (N_8667,N_8233,N_8012);
nand U8668 (N_8668,N_8100,N_8034);
nor U8669 (N_8669,N_8243,N_8068);
or U8670 (N_8670,N_8247,N_8216);
xor U8671 (N_8671,N_8035,N_8379);
nand U8672 (N_8672,N_8084,N_8222);
nand U8673 (N_8673,N_8411,N_8375);
nor U8674 (N_8674,N_8059,N_8201);
or U8675 (N_8675,N_8442,N_8194);
and U8676 (N_8676,N_8333,N_8142);
or U8677 (N_8677,N_8316,N_8332);
nor U8678 (N_8678,N_8245,N_8037);
or U8679 (N_8679,N_8011,N_8018);
xnor U8680 (N_8680,N_8257,N_8458);
nand U8681 (N_8681,N_8071,N_8105);
and U8682 (N_8682,N_8131,N_8402);
or U8683 (N_8683,N_8055,N_8091);
or U8684 (N_8684,N_8177,N_8296);
or U8685 (N_8685,N_8423,N_8443);
or U8686 (N_8686,N_8148,N_8254);
nand U8687 (N_8687,N_8460,N_8286);
nand U8688 (N_8688,N_8165,N_8133);
or U8689 (N_8689,N_8326,N_8054);
or U8690 (N_8690,N_8101,N_8060);
xor U8691 (N_8691,N_8466,N_8171);
nor U8692 (N_8692,N_8495,N_8032);
or U8693 (N_8693,N_8203,N_8026);
or U8694 (N_8694,N_8022,N_8434);
and U8695 (N_8695,N_8023,N_8492);
nand U8696 (N_8696,N_8127,N_8481);
nor U8697 (N_8697,N_8017,N_8139);
nand U8698 (N_8698,N_8360,N_8056);
xnor U8699 (N_8699,N_8452,N_8232);
and U8700 (N_8700,N_8021,N_8085);
and U8701 (N_8701,N_8062,N_8110);
nand U8702 (N_8702,N_8421,N_8323);
nor U8703 (N_8703,N_8029,N_8066);
and U8704 (N_8704,N_8252,N_8474);
or U8705 (N_8705,N_8412,N_8437);
nor U8706 (N_8706,N_8081,N_8113);
and U8707 (N_8707,N_8067,N_8315);
or U8708 (N_8708,N_8106,N_8380);
or U8709 (N_8709,N_8069,N_8489);
nor U8710 (N_8710,N_8486,N_8080);
nor U8711 (N_8711,N_8431,N_8448);
and U8712 (N_8712,N_8228,N_8386);
xor U8713 (N_8713,N_8164,N_8470);
and U8714 (N_8714,N_8266,N_8416);
or U8715 (N_8715,N_8325,N_8230);
nor U8716 (N_8716,N_8163,N_8335);
xnor U8717 (N_8717,N_8451,N_8145);
and U8718 (N_8718,N_8463,N_8392);
or U8719 (N_8719,N_8263,N_8341);
or U8720 (N_8720,N_8258,N_8328);
and U8721 (N_8721,N_8317,N_8295);
nand U8722 (N_8722,N_8246,N_8019);
xor U8723 (N_8723,N_8276,N_8418);
or U8724 (N_8724,N_8298,N_8277);
nor U8725 (N_8725,N_8346,N_8095);
xor U8726 (N_8726,N_8394,N_8117);
nand U8727 (N_8727,N_8293,N_8057);
or U8728 (N_8728,N_8446,N_8065);
xnor U8729 (N_8729,N_8311,N_8179);
xnor U8730 (N_8730,N_8289,N_8074);
or U8731 (N_8731,N_8251,N_8008);
nand U8732 (N_8732,N_8176,N_8042);
or U8733 (N_8733,N_8161,N_8388);
xnor U8734 (N_8734,N_8432,N_8002);
or U8735 (N_8735,N_8140,N_8299);
and U8736 (N_8736,N_8041,N_8291);
nand U8737 (N_8737,N_8102,N_8430);
nand U8738 (N_8738,N_8279,N_8137);
xnor U8739 (N_8739,N_8400,N_8398);
and U8740 (N_8740,N_8212,N_8213);
nand U8741 (N_8741,N_8390,N_8496);
or U8742 (N_8742,N_8015,N_8197);
xor U8743 (N_8743,N_8155,N_8363);
nand U8744 (N_8744,N_8273,N_8135);
or U8745 (N_8745,N_8030,N_8259);
xnor U8746 (N_8746,N_8170,N_8340);
and U8747 (N_8747,N_8319,N_8389);
nor U8748 (N_8748,N_8290,N_8076);
nor U8749 (N_8749,N_8457,N_8087);
nand U8750 (N_8750,N_8091,N_8419);
xor U8751 (N_8751,N_8187,N_8122);
xnor U8752 (N_8752,N_8385,N_8166);
nand U8753 (N_8753,N_8130,N_8389);
xor U8754 (N_8754,N_8246,N_8422);
xor U8755 (N_8755,N_8335,N_8151);
xor U8756 (N_8756,N_8176,N_8066);
nand U8757 (N_8757,N_8101,N_8029);
and U8758 (N_8758,N_8025,N_8026);
nor U8759 (N_8759,N_8055,N_8438);
xor U8760 (N_8760,N_8063,N_8183);
and U8761 (N_8761,N_8401,N_8100);
xnor U8762 (N_8762,N_8115,N_8476);
xnor U8763 (N_8763,N_8028,N_8364);
nand U8764 (N_8764,N_8077,N_8387);
nand U8765 (N_8765,N_8322,N_8398);
or U8766 (N_8766,N_8371,N_8120);
xnor U8767 (N_8767,N_8236,N_8133);
xnor U8768 (N_8768,N_8244,N_8494);
xnor U8769 (N_8769,N_8053,N_8254);
or U8770 (N_8770,N_8346,N_8043);
or U8771 (N_8771,N_8069,N_8180);
xor U8772 (N_8772,N_8498,N_8226);
nand U8773 (N_8773,N_8042,N_8264);
nand U8774 (N_8774,N_8408,N_8079);
nor U8775 (N_8775,N_8059,N_8382);
xor U8776 (N_8776,N_8084,N_8015);
or U8777 (N_8777,N_8431,N_8029);
nor U8778 (N_8778,N_8030,N_8185);
or U8779 (N_8779,N_8382,N_8039);
nor U8780 (N_8780,N_8392,N_8130);
nand U8781 (N_8781,N_8006,N_8131);
xor U8782 (N_8782,N_8091,N_8318);
nand U8783 (N_8783,N_8322,N_8244);
nor U8784 (N_8784,N_8222,N_8073);
or U8785 (N_8785,N_8484,N_8310);
nor U8786 (N_8786,N_8137,N_8476);
nor U8787 (N_8787,N_8479,N_8427);
xnor U8788 (N_8788,N_8041,N_8495);
and U8789 (N_8789,N_8493,N_8364);
nor U8790 (N_8790,N_8384,N_8101);
and U8791 (N_8791,N_8093,N_8431);
nand U8792 (N_8792,N_8339,N_8005);
nand U8793 (N_8793,N_8215,N_8244);
and U8794 (N_8794,N_8267,N_8341);
nand U8795 (N_8795,N_8257,N_8057);
nand U8796 (N_8796,N_8020,N_8162);
nand U8797 (N_8797,N_8012,N_8374);
nand U8798 (N_8798,N_8018,N_8045);
nor U8799 (N_8799,N_8395,N_8266);
and U8800 (N_8800,N_8139,N_8085);
xnor U8801 (N_8801,N_8191,N_8196);
and U8802 (N_8802,N_8496,N_8430);
xor U8803 (N_8803,N_8078,N_8195);
or U8804 (N_8804,N_8196,N_8451);
xor U8805 (N_8805,N_8050,N_8039);
or U8806 (N_8806,N_8404,N_8371);
or U8807 (N_8807,N_8401,N_8134);
and U8808 (N_8808,N_8074,N_8117);
nor U8809 (N_8809,N_8357,N_8225);
xor U8810 (N_8810,N_8399,N_8115);
xnor U8811 (N_8811,N_8303,N_8328);
and U8812 (N_8812,N_8060,N_8416);
nand U8813 (N_8813,N_8270,N_8066);
nor U8814 (N_8814,N_8336,N_8459);
and U8815 (N_8815,N_8394,N_8321);
nand U8816 (N_8816,N_8170,N_8085);
xnor U8817 (N_8817,N_8316,N_8357);
xor U8818 (N_8818,N_8483,N_8352);
or U8819 (N_8819,N_8093,N_8201);
nand U8820 (N_8820,N_8024,N_8071);
xor U8821 (N_8821,N_8152,N_8159);
nor U8822 (N_8822,N_8249,N_8189);
and U8823 (N_8823,N_8161,N_8251);
nor U8824 (N_8824,N_8321,N_8022);
nand U8825 (N_8825,N_8062,N_8168);
xnor U8826 (N_8826,N_8472,N_8074);
nor U8827 (N_8827,N_8465,N_8343);
nor U8828 (N_8828,N_8407,N_8405);
nand U8829 (N_8829,N_8029,N_8282);
and U8830 (N_8830,N_8212,N_8360);
or U8831 (N_8831,N_8093,N_8172);
or U8832 (N_8832,N_8394,N_8189);
nand U8833 (N_8833,N_8106,N_8207);
or U8834 (N_8834,N_8224,N_8113);
nor U8835 (N_8835,N_8346,N_8388);
nor U8836 (N_8836,N_8250,N_8423);
nor U8837 (N_8837,N_8346,N_8476);
and U8838 (N_8838,N_8314,N_8412);
or U8839 (N_8839,N_8204,N_8027);
nor U8840 (N_8840,N_8324,N_8348);
nor U8841 (N_8841,N_8378,N_8166);
and U8842 (N_8842,N_8236,N_8367);
nand U8843 (N_8843,N_8295,N_8491);
xor U8844 (N_8844,N_8281,N_8498);
or U8845 (N_8845,N_8233,N_8485);
or U8846 (N_8846,N_8377,N_8224);
and U8847 (N_8847,N_8034,N_8212);
nor U8848 (N_8848,N_8326,N_8393);
nor U8849 (N_8849,N_8151,N_8210);
or U8850 (N_8850,N_8411,N_8396);
and U8851 (N_8851,N_8407,N_8152);
xnor U8852 (N_8852,N_8186,N_8085);
nor U8853 (N_8853,N_8275,N_8364);
xnor U8854 (N_8854,N_8453,N_8330);
nor U8855 (N_8855,N_8217,N_8252);
xnor U8856 (N_8856,N_8193,N_8389);
nor U8857 (N_8857,N_8291,N_8467);
nor U8858 (N_8858,N_8193,N_8106);
xor U8859 (N_8859,N_8495,N_8366);
xor U8860 (N_8860,N_8254,N_8482);
xnor U8861 (N_8861,N_8470,N_8247);
or U8862 (N_8862,N_8087,N_8266);
nor U8863 (N_8863,N_8179,N_8292);
xor U8864 (N_8864,N_8364,N_8035);
nand U8865 (N_8865,N_8076,N_8295);
and U8866 (N_8866,N_8009,N_8062);
nand U8867 (N_8867,N_8159,N_8035);
nand U8868 (N_8868,N_8390,N_8123);
nor U8869 (N_8869,N_8425,N_8280);
or U8870 (N_8870,N_8380,N_8218);
nor U8871 (N_8871,N_8048,N_8456);
or U8872 (N_8872,N_8437,N_8355);
and U8873 (N_8873,N_8152,N_8461);
nor U8874 (N_8874,N_8217,N_8118);
xor U8875 (N_8875,N_8439,N_8278);
nor U8876 (N_8876,N_8122,N_8382);
nor U8877 (N_8877,N_8072,N_8401);
or U8878 (N_8878,N_8086,N_8482);
nor U8879 (N_8879,N_8172,N_8392);
or U8880 (N_8880,N_8248,N_8394);
xnor U8881 (N_8881,N_8392,N_8431);
nand U8882 (N_8882,N_8236,N_8060);
nor U8883 (N_8883,N_8167,N_8465);
nand U8884 (N_8884,N_8402,N_8363);
xnor U8885 (N_8885,N_8136,N_8232);
and U8886 (N_8886,N_8034,N_8273);
and U8887 (N_8887,N_8004,N_8447);
nand U8888 (N_8888,N_8191,N_8375);
or U8889 (N_8889,N_8111,N_8147);
or U8890 (N_8890,N_8133,N_8290);
nand U8891 (N_8891,N_8303,N_8225);
xnor U8892 (N_8892,N_8447,N_8125);
nor U8893 (N_8893,N_8446,N_8152);
or U8894 (N_8894,N_8462,N_8168);
nor U8895 (N_8895,N_8086,N_8109);
or U8896 (N_8896,N_8471,N_8341);
xnor U8897 (N_8897,N_8069,N_8294);
nor U8898 (N_8898,N_8480,N_8425);
nand U8899 (N_8899,N_8034,N_8454);
or U8900 (N_8900,N_8293,N_8255);
xnor U8901 (N_8901,N_8347,N_8337);
nor U8902 (N_8902,N_8148,N_8437);
nor U8903 (N_8903,N_8079,N_8366);
and U8904 (N_8904,N_8409,N_8292);
nand U8905 (N_8905,N_8111,N_8374);
nand U8906 (N_8906,N_8054,N_8234);
and U8907 (N_8907,N_8223,N_8110);
nor U8908 (N_8908,N_8011,N_8209);
nand U8909 (N_8909,N_8004,N_8493);
nand U8910 (N_8910,N_8446,N_8450);
xor U8911 (N_8911,N_8306,N_8162);
xor U8912 (N_8912,N_8321,N_8447);
nor U8913 (N_8913,N_8366,N_8351);
nand U8914 (N_8914,N_8028,N_8010);
or U8915 (N_8915,N_8265,N_8315);
nor U8916 (N_8916,N_8496,N_8435);
xor U8917 (N_8917,N_8031,N_8339);
and U8918 (N_8918,N_8288,N_8155);
nor U8919 (N_8919,N_8227,N_8060);
or U8920 (N_8920,N_8493,N_8046);
nand U8921 (N_8921,N_8210,N_8471);
nor U8922 (N_8922,N_8435,N_8343);
nand U8923 (N_8923,N_8259,N_8296);
nor U8924 (N_8924,N_8227,N_8219);
nand U8925 (N_8925,N_8405,N_8411);
xor U8926 (N_8926,N_8259,N_8337);
nor U8927 (N_8927,N_8190,N_8283);
nand U8928 (N_8928,N_8009,N_8312);
or U8929 (N_8929,N_8312,N_8407);
or U8930 (N_8930,N_8361,N_8266);
or U8931 (N_8931,N_8071,N_8225);
or U8932 (N_8932,N_8162,N_8469);
xor U8933 (N_8933,N_8375,N_8388);
nand U8934 (N_8934,N_8119,N_8055);
and U8935 (N_8935,N_8023,N_8376);
or U8936 (N_8936,N_8372,N_8334);
or U8937 (N_8937,N_8208,N_8158);
nand U8938 (N_8938,N_8201,N_8352);
or U8939 (N_8939,N_8333,N_8358);
nor U8940 (N_8940,N_8236,N_8121);
xor U8941 (N_8941,N_8152,N_8210);
and U8942 (N_8942,N_8058,N_8447);
and U8943 (N_8943,N_8220,N_8165);
nor U8944 (N_8944,N_8222,N_8198);
or U8945 (N_8945,N_8069,N_8126);
or U8946 (N_8946,N_8110,N_8437);
xnor U8947 (N_8947,N_8158,N_8064);
xor U8948 (N_8948,N_8260,N_8070);
and U8949 (N_8949,N_8343,N_8107);
nand U8950 (N_8950,N_8138,N_8162);
xor U8951 (N_8951,N_8465,N_8375);
and U8952 (N_8952,N_8344,N_8233);
xnor U8953 (N_8953,N_8333,N_8388);
xor U8954 (N_8954,N_8374,N_8003);
and U8955 (N_8955,N_8163,N_8141);
and U8956 (N_8956,N_8455,N_8393);
xor U8957 (N_8957,N_8344,N_8499);
nor U8958 (N_8958,N_8352,N_8141);
or U8959 (N_8959,N_8150,N_8492);
nor U8960 (N_8960,N_8449,N_8429);
and U8961 (N_8961,N_8241,N_8314);
or U8962 (N_8962,N_8183,N_8333);
xnor U8963 (N_8963,N_8286,N_8426);
nand U8964 (N_8964,N_8228,N_8344);
nor U8965 (N_8965,N_8302,N_8158);
nand U8966 (N_8966,N_8105,N_8319);
and U8967 (N_8967,N_8345,N_8241);
nor U8968 (N_8968,N_8111,N_8490);
and U8969 (N_8969,N_8145,N_8457);
xor U8970 (N_8970,N_8031,N_8393);
nand U8971 (N_8971,N_8427,N_8383);
or U8972 (N_8972,N_8352,N_8476);
xor U8973 (N_8973,N_8002,N_8480);
and U8974 (N_8974,N_8202,N_8370);
or U8975 (N_8975,N_8063,N_8356);
or U8976 (N_8976,N_8258,N_8188);
nor U8977 (N_8977,N_8181,N_8136);
nor U8978 (N_8978,N_8376,N_8243);
nor U8979 (N_8979,N_8182,N_8277);
and U8980 (N_8980,N_8118,N_8253);
xor U8981 (N_8981,N_8027,N_8432);
nand U8982 (N_8982,N_8384,N_8071);
and U8983 (N_8983,N_8318,N_8335);
and U8984 (N_8984,N_8085,N_8297);
nor U8985 (N_8985,N_8417,N_8303);
or U8986 (N_8986,N_8196,N_8017);
and U8987 (N_8987,N_8289,N_8434);
nand U8988 (N_8988,N_8091,N_8312);
and U8989 (N_8989,N_8054,N_8492);
nor U8990 (N_8990,N_8252,N_8484);
nor U8991 (N_8991,N_8031,N_8221);
nand U8992 (N_8992,N_8091,N_8274);
or U8993 (N_8993,N_8173,N_8332);
or U8994 (N_8994,N_8018,N_8362);
xor U8995 (N_8995,N_8011,N_8419);
and U8996 (N_8996,N_8259,N_8286);
and U8997 (N_8997,N_8154,N_8381);
or U8998 (N_8998,N_8192,N_8492);
and U8999 (N_8999,N_8231,N_8253);
or U9000 (N_9000,N_8668,N_8886);
nor U9001 (N_9001,N_8665,N_8870);
nor U9002 (N_9002,N_8897,N_8734);
and U9003 (N_9003,N_8909,N_8514);
and U9004 (N_9004,N_8509,N_8993);
nor U9005 (N_9005,N_8874,N_8920);
nand U9006 (N_9006,N_8823,N_8703);
nand U9007 (N_9007,N_8721,N_8917);
or U9008 (N_9008,N_8905,N_8607);
xor U9009 (N_9009,N_8597,N_8613);
or U9010 (N_9010,N_8506,N_8535);
and U9011 (N_9011,N_8912,N_8564);
nor U9012 (N_9012,N_8657,N_8804);
xnor U9013 (N_9013,N_8619,N_8902);
or U9014 (N_9014,N_8572,N_8966);
nor U9015 (N_9015,N_8772,N_8798);
xor U9016 (N_9016,N_8876,N_8853);
xor U9017 (N_9017,N_8933,N_8750);
xor U9018 (N_9018,N_8774,N_8697);
nor U9019 (N_9019,N_8805,N_8988);
xor U9020 (N_9020,N_8743,N_8531);
or U9021 (N_9021,N_8522,N_8543);
xor U9022 (N_9022,N_8907,N_8682);
or U9023 (N_9023,N_8625,N_8930);
nand U9024 (N_9024,N_8677,N_8960);
or U9025 (N_9025,N_8860,N_8985);
or U9026 (N_9026,N_8515,N_8761);
xnor U9027 (N_9027,N_8797,N_8633);
nor U9028 (N_9028,N_8827,N_8866);
or U9029 (N_9029,N_8767,N_8675);
nand U9030 (N_9030,N_8789,N_8887);
xnor U9031 (N_9031,N_8501,N_8710);
xor U9032 (N_9032,N_8626,N_8526);
nand U9033 (N_9033,N_8698,N_8537);
nor U9034 (N_9034,N_8661,N_8970);
nor U9035 (N_9035,N_8769,N_8932);
nor U9036 (N_9036,N_8673,N_8900);
or U9037 (N_9037,N_8948,N_8742);
nor U9038 (N_9038,N_8590,N_8819);
xor U9039 (N_9039,N_8906,N_8878);
nor U9040 (N_9040,N_8812,N_8503);
nor U9041 (N_9041,N_8521,N_8771);
or U9042 (N_9042,N_8719,N_8951);
nor U9043 (N_9043,N_8723,N_8760);
nand U9044 (N_9044,N_8645,N_8541);
and U9045 (N_9045,N_8554,N_8781);
or U9046 (N_9046,N_8570,N_8835);
nor U9047 (N_9047,N_8931,N_8623);
nor U9048 (N_9048,N_8938,N_8893);
nand U9049 (N_9049,N_8705,N_8502);
and U9050 (N_9050,N_8943,N_8962);
and U9051 (N_9051,N_8518,N_8552);
xnor U9052 (N_9052,N_8764,N_8504);
nand U9053 (N_9053,N_8660,N_8969);
nand U9054 (N_9054,N_8785,N_8810);
nor U9055 (N_9055,N_8696,N_8953);
xor U9056 (N_9056,N_8844,N_8791);
and U9057 (N_9057,N_8593,N_8620);
nor U9058 (N_9058,N_8641,N_8701);
or U9059 (N_9059,N_8542,N_8891);
nand U9060 (N_9060,N_8671,N_8957);
and U9061 (N_9061,N_8861,N_8699);
and U9062 (N_9062,N_8702,N_8651);
xnor U9063 (N_9063,N_8792,N_8763);
nand U9064 (N_9064,N_8777,N_8825);
nand U9065 (N_9065,N_8984,N_8881);
nor U9066 (N_9066,N_8756,N_8987);
nand U9067 (N_9067,N_8606,N_8865);
xor U9068 (N_9068,N_8632,N_8601);
nand U9069 (N_9069,N_8654,N_8565);
nor U9070 (N_9070,N_8867,N_8562);
and U9071 (N_9071,N_8811,N_8991);
nor U9072 (N_9072,N_8582,N_8744);
or U9073 (N_9073,N_8815,N_8855);
nor U9074 (N_9074,N_8868,N_8611);
and U9075 (N_9075,N_8954,N_8707);
and U9076 (N_9076,N_8599,N_8600);
and U9077 (N_9077,N_8924,N_8944);
nor U9078 (N_9078,N_8910,N_8643);
and U9079 (N_9079,N_8624,N_8759);
nand U9080 (N_9080,N_8755,N_8691);
nor U9081 (N_9081,N_8783,N_8879);
or U9082 (N_9082,N_8642,N_8901);
or U9083 (N_9083,N_8809,N_8929);
or U9084 (N_9084,N_8903,N_8637);
or U9085 (N_9085,N_8851,N_8813);
xnor U9086 (N_9086,N_8990,N_8708);
xor U9087 (N_9087,N_8534,N_8549);
nand U9088 (N_9088,N_8629,N_8500);
and U9089 (N_9089,N_8739,N_8834);
xor U9090 (N_9090,N_8529,N_8605);
nor U9091 (N_9091,N_8919,N_8892);
or U9092 (N_9092,N_8639,N_8816);
or U9093 (N_9093,N_8681,N_8945);
xnor U9094 (N_9094,N_8971,N_8553);
xnor U9095 (N_9095,N_8532,N_8545);
xor U9096 (N_9096,N_8687,N_8609);
or U9097 (N_9097,N_8894,N_8975);
nor U9098 (N_9098,N_8658,N_8652);
and U9099 (N_9099,N_8852,N_8830);
nand U9100 (N_9100,N_8826,N_8575);
xnor U9101 (N_9101,N_8822,N_8524);
or U9102 (N_9102,N_8776,N_8968);
and U9103 (N_9103,N_8621,N_8539);
xor U9104 (N_9104,N_8693,N_8753);
and U9105 (N_9105,N_8567,N_8690);
nand U9106 (N_9106,N_8616,N_8536);
nand U9107 (N_9107,N_8603,N_8680);
nor U9108 (N_9108,N_8807,N_8561);
and U9109 (N_9109,N_8936,N_8731);
xnor U9110 (N_9110,N_8836,N_8821);
or U9111 (N_9111,N_8726,N_8550);
nand U9112 (N_9112,N_8634,N_8847);
xor U9113 (N_9113,N_8981,N_8854);
and U9114 (N_9114,N_8588,N_8577);
and U9115 (N_9115,N_8982,N_8568);
xor U9116 (N_9116,N_8995,N_8662);
or U9117 (N_9117,N_8942,N_8749);
or U9118 (N_9118,N_8841,N_8875);
or U9119 (N_9119,N_8544,N_8628);
nor U9120 (N_9120,N_8926,N_8795);
nor U9121 (N_9121,N_8725,N_8558);
or U9122 (N_9122,N_8525,N_8997);
xnor U9123 (N_9123,N_8832,N_8747);
nor U9124 (N_9124,N_8846,N_8559);
xnor U9125 (N_9125,N_8678,N_8928);
and U9126 (N_9126,N_8689,N_8820);
nand U9127 (N_9127,N_8516,N_8869);
xor U9128 (N_9128,N_8730,N_8923);
xor U9129 (N_9129,N_8676,N_8937);
and U9130 (N_9130,N_8818,N_8838);
nor U9131 (N_9131,N_8779,N_8967);
or U9132 (N_9132,N_8873,N_8646);
or U9133 (N_9133,N_8700,N_8848);
nand U9134 (N_9134,N_8576,N_8800);
nor U9135 (N_9135,N_8947,N_8788);
nand U9136 (N_9136,N_8638,N_8569);
xor U9137 (N_9137,N_8890,N_8683);
and U9138 (N_9138,N_8794,N_8704);
nor U9139 (N_9139,N_8663,N_8956);
xnor U9140 (N_9140,N_8610,N_8915);
xor U9141 (N_9141,N_8512,N_8738);
nor U9142 (N_9142,N_8728,N_8899);
and U9143 (N_9143,N_8584,N_8612);
nand U9144 (N_9144,N_8883,N_8941);
and U9145 (N_9145,N_8862,N_8762);
nor U9146 (N_9146,N_8790,N_8980);
nand U9147 (N_9147,N_8801,N_8591);
xnor U9148 (N_9148,N_8972,N_8713);
or U9149 (N_9149,N_8729,N_8959);
nor U9150 (N_9150,N_8799,N_8806);
xor U9151 (N_9151,N_8934,N_8914);
and U9152 (N_9152,N_8950,N_8670);
nand U9153 (N_9153,N_8732,N_8692);
or U9154 (N_9154,N_8908,N_8655);
and U9155 (N_9155,N_8566,N_8857);
or U9156 (N_9156,N_8557,N_8608);
xnor U9157 (N_9157,N_8840,N_8647);
and U9158 (N_9158,N_8589,N_8508);
and U9159 (N_9159,N_8979,N_8527);
nand U9160 (N_9160,N_8858,N_8961);
nand U9161 (N_9161,N_8709,N_8921);
xor U9162 (N_9162,N_8679,N_8793);
or U9163 (N_9163,N_8829,N_8674);
xnor U9164 (N_9164,N_8712,N_8648);
and U9165 (N_9165,N_8911,N_8998);
nor U9166 (N_9166,N_8556,N_8745);
xnor U9167 (N_9167,N_8940,N_8973);
xnor U9168 (N_9168,N_8735,N_8754);
or U9169 (N_9169,N_8752,N_8630);
xor U9170 (N_9170,N_8555,N_8877);
nand U9171 (N_9171,N_8685,N_8839);
nand U9172 (N_9172,N_8751,N_8916);
nand U9173 (N_9173,N_8837,N_8617);
nor U9174 (N_9174,N_8775,N_8579);
nand U9175 (N_9175,N_8653,N_8737);
nand U9176 (N_9176,N_8814,N_8644);
nor U9177 (N_9177,N_8574,N_8952);
and U9178 (N_9178,N_8585,N_8672);
and U9179 (N_9179,N_8727,N_8664);
nor U9180 (N_9180,N_8859,N_8864);
or U9181 (N_9181,N_8802,N_8578);
xor U9182 (N_9182,N_8746,N_8547);
nand U9183 (N_9183,N_8640,N_8996);
and U9184 (N_9184,N_8656,N_8786);
nor U9185 (N_9185,N_8964,N_8635);
nor U9186 (N_9186,N_8817,N_8833);
or U9187 (N_9187,N_8520,N_8627);
nand U9188 (N_9188,N_8949,N_8856);
or U9189 (N_9189,N_8718,N_8989);
and U9190 (N_9190,N_8782,N_8885);
xnor U9191 (N_9191,N_8770,N_8530);
or U9192 (N_9192,N_8695,N_8884);
or U9193 (N_9193,N_8551,N_8935);
or U9194 (N_9194,N_8958,N_8803);
or U9195 (N_9195,N_8778,N_8604);
and U9196 (N_9196,N_8872,N_8733);
or U9197 (N_9197,N_8974,N_8882);
xor U9198 (N_9198,N_8898,N_8850);
or U9199 (N_9199,N_8592,N_8888);
nor U9200 (N_9200,N_8711,N_8824);
xor U9201 (N_9201,N_8849,N_8740);
nor U9202 (N_9202,N_8618,N_8507);
xnor U9203 (N_9203,N_8517,N_8649);
xnor U9204 (N_9204,N_8598,N_8863);
or U9205 (N_9205,N_8758,N_8983);
nand U9206 (N_9206,N_8880,N_8581);
and U9207 (N_9207,N_8533,N_8736);
or U9208 (N_9208,N_8538,N_8965);
nor U9209 (N_9209,N_8595,N_8540);
nor U9210 (N_9210,N_8828,N_8913);
or U9211 (N_9211,N_8845,N_8741);
or U9212 (N_9212,N_8636,N_8918);
and U9213 (N_9213,N_8684,N_8724);
and U9214 (N_9214,N_8622,N_8748);
xor U9215 (N_9215,N_8780,N_8717);
xor U9216 (N_9216,N_8773,N_8784);
or U9217 (N_9217,N_8895,N_8602);
or U9218 (N_9218,N_8714,N_8955);
xnor U9219 (N_9219,N_8528,N_8992);
and U9220 (N_9220,N_8716,N_8571);
and U9221 (N_9221,N_8994,N_8548);
and U9222 (N_9222,N_8511,N_8586);
or U9223 (N_9223,N_8922,N_8896);
xnor U9224 (N_9224,N_8766,N_8583);
or U9225 (N_9225,N_8505,N_8889);
nor U9226 (N_9226,N_8688,N_8631);
xnor U9227 (N_9227,N_8523,N_8843);
nor U9228 (N_9228,N_8978,N_8615);
or U9229 (N_9229,N_8686,N_8715);
and U9230 (N_9230,N_8666,N_8720);
and U9231 (N_9231,N_8706,N_8667);
or U9232 (N_9232,N_8796,N_8986);
and U9233 (N_9233,N_8939,N_8513);
nand U9234 (N_9234,N_8831,N_8510);
nor U9235 (N_9235,N_8614,N_8946);
nor U9236 (N_9236,N_8808,N_8563);
nor U9237 (N_9237,N_8768,N_8659);
nor U9238 (N_9238,N_8925,N_8587);
and U9239 (N_9239,N_8787,N_8977);
xnor U9240 (N_9240,N_8519,N_8650);
nor U9241 (N_9241,N_8765,N_8963);
nor U9242 (N_9242,N_8580,N_8669);
and U9243 (N_9243,N_8871,N_8927);
nor U9244 (N_9244,N_8596,N_8976);
or U9245 (N_9245,N_8573,N_8722);
nor U9246 (N_9246,N_8904,N_8999);
nand U9247 (N_9247,N_8546,N_8560);
nor U9248 (N_9248,N_8694,N_8757);
or U9249 (N_9249,N_8842,N_8594);
and U9250 (N_9250,N_8762,N_8501);
nor U9251 (N_9251,N_8754,N_8526);
nor U9252 (N_9252,N_8909,N_8868);
and U9253 (N_9253,N_8598,N_8851);
and U9254 (N_9254,N_8843,N_8747);
xnor U9255 (N_9255,N_8669,N_8845);
nand U9256 (N_9256,N_8897,N_8700);
nand U9257 (N_9257,N_8901,N_8927);
nor U9258 (N_9258,N_8736,N_8568);
and U9259 (N_9259,N_8714,N_8822);
nor U9260 (N_9260,N_8670,N_8750);
nor U9261 (N_9261,N_8881,N_8742);
xnor U9262 (N_9262,N_8918,N_8807);
and U9263 (N_9263,N_8686,N_8701);
nor U9264 (N_9264,N_8641,N_8960);
nand U9265 (N_9265,N_8841,N_8772);
and U9266 (N_9266,N_8766,N_8588);
nand U9267 (N_9267,N_8747,N_8995);
and U9268 (N_9268,N_8905,N_8541);
nor U9269 (N_9269,N_8674,N_8907);
nor U9270 (N_9270,N_8524,N_8928);
or U9271 (N_9271,N_8876,N_8946);
nor U9272 (N_9272,N_8870,N_8694);
nand U9273 (N_9273,N_8884,N_8842);
xnor U9274 (N_9274,N_8832,N_8983);
nor U9275 (N_9275,N_8865,N_8803);
and U9276 (N_9276,N_8613,N_8960);
or U9277 (N_9277,N_8526,N_8845);
nand U9278 (N_9278,N_8575,N_8714);
or U9279 (N_9279,N_8680,N_8745);
nor U9280 (N_9280,N_8679,N_8645);
xor U9281 (N_9281,N_8519,N_8510);
xnor U9282 (N_9282,N_8592,N_8971);
and U9283 (N_9283,N_8656,N_8920);
nor U9284 (N_9284,N_8727,N_8745);
and U9285 (N_9285,N_8598,N_8822);
nor U9286 (N_9286,N_8941,N_8510);
and U9287 (N_9287,N_8792,N_8661);
xnor U9288 (N_9288,N_8862,N_8815);
or U9289 (N_9289,N_8740,N_8541);
nor U9290 (N_9290,N_8653,N_8764);
or U9291 (N_9291,N_8780,N_8867);
xor U9292 (N_9292,N_8619,N_8864);
or U9293 (N_9293,N_8561,N_8918);
or U9294 (N_9294,N_8895,N_8721);
nor U9295 (N_9295,N_8818,N_8951);
or U9296 (N_9296,N_8867,N_8930);
nand U9297 (N_9297,N_8644,N_8839);
and U9298 (N_9298,N_8551,N_8619);
and U9299 (N_9299,N_8877,N_8895);
nand U9300 (N_9300,N_8595,N_8534);
or U9301 (N_9301,N_8900,N_8823);
nor U9302 (N_9302,N_8762,N_8816);
xor U9303 (N_9303,N_8986,N_8574);
nor U9304 (N_9304,N_8942,N_8833);
nor U9305 (N_9305,N_8529,N_8571);
nor U9306 (N_9306,N_8758,N_8725);
nor U9307 (N_9307,N_8913,N_8517);
nand U9308 (N_9308,N_8990,N_8748);
and U9309 (N_9309,N_8584,N_8564);
and U9310 (N_9310,N_8632,N_8754);
nor U9311 (N_9311,N_8752,N_8898);
or U9312 (N_9312,N_8584,N_8561);
nand U9313 (N_9313,N_8989,N_8619);
nor U9314 (N_9314,N_8879,N_8903);
xnor U9315 (N_9315,N_8758,N_8529);
nand U9316 (N_9316,N_8877,N_8522);
nand U9317 (N_9317,N_8888,N_8981);
xnor U9318 (N_9318,N_8613,N_8565);
nor U9319 (N_9319,N_8837,N_8692);
and U9320 (N_9320,N_8552,N_8947);
xnor U9321 (N_9321,N_8517,N_8536);
or U9322 (N_9322,N_8693,N_8580);
nand U9323 (N_9323,N_8943,N_8537);
xnor U9324 (N_9324,N_8587,N_8806);
xor U9325 (N_9325,N_8742,N_8536);
xor U9326 (N_9326,N_8515,N_8800);
and U9327 (N_9327,N_8756,N_8889);
or U9328 (N_9328,N_8687,N_8676);
xnor U9329 (N_9329,N_8990,N_8905);
or U9330 (N_9330,N_8640,N_8771);
nor U9331 (N_9331,N_8795,N_8702);
nor U9332 (N_9332,N_8567,N_8827);
or U9333 (N_9333,N_8722,N_8926);
nand U9334 (N_9334,N_8616,N_8875);
xnor U9335 (N_9335,N_8727,N_8832);
and U9336 (N_9336,N_8543,N_8618);
nor U9337 (N_9337,N_8820,N_8991);
and U9338 (N_9338,N_8572,N_8781);
and U9339 (N_9339,N_8632,N_8646);
nand U9340 (N_9340,N_8911,N_8944);
nand U9341 (N_9341,N_8579,N_8877);
nor U9342 (N_9342,N_8686,N_8582);
and U9343 (N_9343,N_8874,N_8541);
and U9344 (N_9344,N_8884,N_8995);
and U9345 (N_9345,N_8810,N_8984);
nand U9346 (N_9346,N_8869,N_8539);
xnor U9347 (N_9347,N_8945,N_8558);
nand U9348 (N_9348,N_8703,N_8649);
nand U9349 (N_9349,N_8584,N_8940);
or U9350 (N_9350,N_8977,N_8617);
xor U9351 (N_9351,N_8967,N_8517);
and U9352 (N_9352,N_8958,N_8878);
and U9353 (N_9353,N_8981,N_8708);
nand U9354 (N_9354,N_8849,N_8579);
and U9355 (N_9355,N_8807,N_8932);
and U9356 (N_9356,N_8891,N_8611);
nand U9357 (N_9357,N_8698,N_8727);
nor U9358 (N_9358,N_8974,N_8563);
nand U9359 (N_9359,N_8828,N_8665);
xor U9360 (N_9360,N_8743,N_8791);
nand U9361 (N_9361,N_8881,N_8553);
and U9362 (N_9362,N_8652,N_8991);
nand U9363 (N_9363,N_8776,N_8834);
and U9364 (N_9364,N_8991,N_8893);
xnor U9365 (N_9365,N_8951,N_8613);
or U9366 (N_9366,N_8599,N_8640);
nand U9367 (N_9367,N_8879,N_8611);
nor U9368 (N_9368,N_8981,N_8847);
and U9369 (N_9369,N_8776,N_8631);
and U9370 (N_9370,N_8920,N_8872);
or U9371 (N_9371,N_8641,N_8716);
nor U9372 (N_9372,N_8920,N_8775);
nor U9373 (N_9373,N_8556,N_8897);
nand U9374 (N_9374,N_8800,N_8806);
nand U9375 (N_9375,N_8638,N_8556);
nor U9376 (N_9376,N_8882,N_8992);
nand U9377 (N_9377,N_8810,N_8978);
xor U9378 (N_9378,N_8617,N_8674);
xnor U9379 (N_9379,N_8510,N_8848);
nand U9380 (N_9380,N_8729,N_8580);
xnor U9381 (N_9381,N_8612,N_8595);
and U9382 (N_9382,N_8748,N_8571);
nor U9383 (N_9383,N_8548,N_8780);
nand U9384 (N_9384,N_8631,N_8778);
xor U9385 (N_9385,N_8535,N_8802);
nor U9386 (N_9386,N_8673,N_8731);
and U9387 (N_9387,N_8599,N_8524);
nor U9388 (N_9388,N_8669,N_8955);
xnor U9389 (N_9389,N_8634,N_8970);
nand U9390 (N_9390,N_8722,N_8510);
nand U9391 (N_9391,N_8559,N_8688);
nand U9392 (N_9392,N_8637,N_8814);
or U9393 (N_9393,N_8579,N_8903);
nand U9394 (N_9394,N_8505,N_8597);
and U9395 (N_9395,N_8663,N_8924);
or U9396 (N_9396,N_8748,N_8987);
and U9397 (N_9397,N_8869,N_8815);
nor U9398 (N_9398,N_8597,N_8952);
xor U9399 (N_9399,N_8978,N_8943);
nor U9400 (N_9400,N_8861,N_8512);
nand U9401 (N_9401,N_8563,N_8955);
xnor U9402 (N_9402,N_8841,N_8822);
nor U9403 (N_9403,N_8921,N_8831);
nor U9404 (N_9404,N_8526,N_8554);
nand U9405 (N_9405,N_8526,N_8552);
nand U9406 (N_9406,N_8564,N_8565);
and U9407 (N_9407,N_8688,N_8608);
nor U9408 (N_9408,N_8795,N_8554);
xor U9409 (N_9409,N_8707,N_8765);
and U9410 (N_9410,N_8958,N_8873);
or U9411 (N_9411,N_8691,N_8980);
and U9412 (N_9412,N_8780,N_8675);
or U9413 (N_9413,N_8911,N_8878);
nand U9414 (N_9414,N_8651,N_8896);
or U9415 (N_9415,N_8643,N_8878);
nand U9416 (N_9416,N_8766,N_8713);
or U9417 (N_9417,N_8668,N_8566);
xor U9418 (N_9418,N_8717,N_8841);
and U9419 (N_9419,N_8624,N_8842);
nand U9420 (N_9420,N_8746,N_8929);
xor U9421 (N_9421,N_8705,N_8615);
and U9422 (N_9422,N_8740,N_8550);
nor U9423 (N_9423,N_8721,N_8706);
or U9424 (N_9424,N_8769,N_8774);
and U9425 (N_9425,N_8552,N_8932);
nor U9426 (N_9426,N_8721,N_8622);
or U9427 (N_9427,N_8802,N_8553);
nor U9428 (N_9428,N_8522,N_8938);
nand U9429 (N_9429,N_8886,N_8755);
nand U9430 (N_9430,N_8542,N_8619);
xnor U9431 (N_9431,N_8616,N_8577);
nand U9432 (N_9432,N_8750,N_8838);
or U9433 (N_9433,N_8989,N_8677);
or U9434 (N_9434,N_8539,N_8825);
nand U9435 (N_9435,N_8614,N_8996);
xor U9436 (N_9436,N_8982,N_8814);
nor U9437 (N_9437,N_8876,N_8846);
nand U9438 (N_9438,N_8640,N_8716);
nand U9439 (N_9439,N_8997,N_8885);
nand U9440 (N_9440,N_8834,N_8705);
or U9441 (N_9441,N_8559,N_8960);
nor U9442 (N_9442,N_8718,N_8816);
xnor U9443 (N_9443,N_8950,N_8973);
and U9444 (N_9444,N_8898,N_8832);
nor U9445 (N_9445,N_8563,N_8533);
nand U9446 (N_9446,N_8730,N_8525);
xor U9447 (N_9447,N_8808,N_8825);
xor U9448 (N_9448,N_8563,N_8858);
and U9449 (N_9449,N_8503,N_8572);
xnor U9450 (N_9450,N_8757,N_8911);
nor U9451 (N_9451,N_8885,N_8901);
xor U9452 (N_9452,N_8546,N_8949);
or U9453 (N_9453,N_8949,N_8779);
nor U9454 (N_9454,N_8578,N_8884);
or U9455 (N_9455,N_8626,N_8788);
and U9456 (N_9456,N_8717,N_8734);
nand U9457 (N_9457,N_8653,N_8752);
xor U9458 (N_9458,N_8720,N_8813);
and U9459 (N_9459,N_8726,N_8527);
nor U9460 (N_9460,N_8983,N_8696);
nand U9461 (N_9461,N_8679,N_8571);
xnor U9462 (N_9462,N_8993,N_8826);
or U9463 (N_9463,N_8765,N_8664);
nand U9464 (N_9464,N_8729,N_8916);
nor U9465 (N_9465,N_8765,N_8647);
nor U9466 (N_9466,N_8987,N_8876);
xor U9467 (N_9467,N_8556,N_8839);
nand U9468 (N_9468,N_8698,N_8942);
xor U9469 (N_9469,N_8649,N_8824);
nor U9470 (N_9470,N_8659,N_8847);
nor U9471 (N_9471,N_8540,N_8749);
xor U9472 (N_9472,N_8869,N_8743);
xnor U9473 (N_9473,N_8566,N_8546);
nand U9474 (N_9474,N_8520,N_8809);
or U9475 (N_9475,N_8708,N_8643);
xor U9476 (N_9476,N_8525,N_8887);
nor U9477 (N_9477,N_8508,N_8863);
or U9478 (N_9478,N_8569,N_8922);
nor U9479 (N_9479,N_8634,N_8771);
and U9480 (N_9480,N_8714,N_8744);
nor U9481 (N_9481,N_8679,N_8954);
xor U9482 (N_9482,N_8802,N_8587);
nand U9483 (N_9483,N_8943,N_8819);
or U9484 (N_9484,N_8611,N_8656);
nand U9485 (N_9485,N_8701,N_8958);
and U9486 (N_9486,N_8853,N_8646);
xor U9487 (N_9487,N_8854,N_8600);
and U9488 (N_9488,N_8534,N_8872);
or U9489 (N_9489,N_8736,N_8619);
xnor U9490 (N_9490,N_8581,N_8979);
nor U9491 (N_9491,N_8715,N_8922);
nor U9492 (N_9492,N_8864,N_8706);
nor U9493 (N_9493,N_8865,N_8586);
and U9494 (N_9494,N_8509,N_8943);
and U9495 (N_9495,N_8964,N_8908);
xor U9496 (N_9496,N_8577,N_8942);
nand U9497 (N_9497,N_8526,N_8624);
nor U9498 (N_9498,N_8829,N_8553);
and U9499 (N_9499,N_8612,N_8724);
or U9500 (N_9500,N_9289,N_9422);
nand U9501 (N_9501,N_9140,N_9241);
or U9502 (N_9502,N_9233,N_9042);
nor U9503 (N_9503,N_9460,N_9213);
xnor U9504 (N_9504,N_9310,N_9069);
nor U9505 (N_9505,N_9330,N_9483);
or U9506 (N_9506,N_9268,N_9141);
nand U9507 (N_9507,N_9031,N_9305);
nor U9508 (N_9508,N_9371,N_9368);
xnor U9509 (N_9509,N_9254,N_9291);
and U9510 (N_9510,N_9477,N_9232);
or U9511 (N_9511,N_9391,N_9252);
and U9512 (N_9512,N_9028,N_9411);
or U9513 (N_9513,N_9463,N_9376);
xnor U9514 (N_9514,N_9004,N_9156);
xor U9515 (N_9515,N_9261,N_9111);
nand U9516 (N_9516,N_9114,N_9340);
nor U9517 (N_9517,N_9064,N_9244);
nor U9518 (N_9518,N_9488,N_9467);
nor U9519 (N_9519,N_9365,N_9487);
or U9520 (N_9520,N_9033,N_9096);
xnor U9521 (N_9521,N_9209,N_9017);
nor U9522 (N_9522,N_9032,N_9492);
xor U9523 (N_9523,N_9360,N_9200);
and U9524 (N_9524,N_9021,N_9165);
or U9525 (N_9525,N_9377,N_9351);
and U9526 (N_9526,N_9274,N_9001);
nor U9527 (N_9527,N_9388,N_9191);
or U9528 (N_9528,N_9227,N_9195);
or U9529 (N_9529,N_9112,N_9041);
and U9530 (N_9530,N_9440,N_9426);
xnor U9531 (N_9531,N_9250,N_9326);
and U9532 (N_9532,N_9445,N_9364);
or U9533 (N_9533,N_9392,N_9037);
xnor U9534 (N_9534,N_9303,N_9089);
and U9535 (N_9535,N_9016,N_9188);
or U9536 (N_9536,N_9309,N_9234);
and U9537 (N_9537,N_9394,N_9217);
xnor U9538 (N_9538,N_9466,N_9007);
xor U9539 (N_9539,N_9399,N_9204);
nand U9540 (N_9540,N_9318,N_9137);
nor U9541 (N_9541,N_9409,N_9384);
nand U9542 (N_9542,N_9489,N_9459);
or U9543 (N_9543,N_9443,N_9157);
or U9544 (N_9544,N_9336,N_9150);
or U9545 (N_9545,N_9103,N_9434);
nor U9546 (N_9546,N_9138,N_9229);
xor U9547 (N_9547,N_9495,N_9038);
xor U9548 (N_9548,N_9446,N_9171);
nor U9549 (N_9549,N_9148,N_9108);
or U9550 (N_9550,N_9343,N_9239);
xnor U9551 (N_9551,N_9494,N_9243);
nand U9552 (N_9552,N_9224,N_9248);
nor U9553 (N_9553,N_9086,N_9363);
nor U9554 (N_9554,N_9005,N_9258);
nor U9555 (N_9555,N_9453,N_9283);
and U9556 (N_9556,N_9183,N_9199);
and U9557 (N_9557,N_9078,N_9170);
nor U9558 (N_9558,N_9350,N_9272);
nand U9559 (N_9559,N_9127,N_9290);
and U9560 (N_9560,N_9058,N_9079);
and U9561 (N_9561,N_9092,N_9202);
nor U9562 (N_9562,N_9382,N_9359);
nor U9563 (N_9563,N_9378,N_9410);
xor U9564 (N_9564,N_9369,N_9294);
xor U9565 (N_9565,N_9119,N_9120);
nand U9566 (N_9566,N_9315,N_9374);
nand U9567 (N_9567,N_9436,N_9237);
and U9568 (N_9568,N_9299,N_9347);
xor U9569 (N_9569,N_9295,N_9400);
nand U9570 (N_9570,N_9088,N_9383);
and U9571 (N_9571,N_9113,N_9065);
nor U9572 (N_9572,N_9471,N_9184);
and U9573 (N_9573,N_9068,N_9320);
nor U9574 (N_9574,N_9216,N_9415);
xor U9575 (N_9575,N_9266,N_9214);
and U9576 (N_9576,N_9050,N_9473);
nand U9577 (N_9577,N_9029,N_9370);
and U9578 (N_9578,N_9276,N_9063);
nor U9579 (N_9579,N_9334,N_9010);
and U9580 (N_9580,N_9132,N_9251);
xnor U9581 (N_9581,N_9339,N_9265);
or U9582 (N_9582,N_9052,N_9212);
nand U9583 (N_9583,N_9208,N_9301);
and U9584 (N_9584,N_9269,N_9462);
or U9585 (N_9585,N_9264,N_9332);
nand U9586 (N_9586,N_9327,N_9403);
xor U9587 (N_9587,N_9277,N_9284);
or U9588 (N_9588,N_9121,N_9297);
or U9589 (N_9589,N_9329,N_9313);
or U9590 (N_9590,N_9051,N_9448);
and U9591 (N_9591,N_9349,N_9348);
or U9592 (N_9592,N_9135,N_9231);
xnor U9593 (N_9593,N_9030,N_9099);
nand U9594 (N_9594,N_9133,N_9493);
xnor U9595 (N_9595,N_9172,N_9040);
xnor U9596 (N_9596,N_9091,N_9452);
or U9597 (N_9597,N_9389,N_9161);
nor U9598 (N_9598,N_9198,N_9366);
and U9599 (N_9599,N_9177,N_9149);
nor U9600 (N_9600,N_9090,N_9036);
and U9601 (N_9601,N_9357,N_9262);
and U9602 (N_9602,N_9201,N_9084);
and U9603 (N_9603,N_9444,N_9255);
or U9604 (N_9604,N_9168,N_9110);
xor U9605 (N_9605,N_9358,N_9014);
nor U9606 (N_9606,N_9438,N_9454);
and U9607 (N_9607,N_9273,N_9481);
nor U9608 (N_9608,N_9421,N_9047);
xor U9609 (N_9609,N_9093,N_9203);
nor U9610 (N_9610,N_9257,N_9129);
nor U9611 (N_9611,N_9053,N_9468);
and U9612 (N_9612,N_9196,N_9020);
and U9613 (N_9613,N_9484,N_9083);
nand U9614 (N_9614,N_9354,N_9151);
nand U9615 (N_9615,N_9026,N_9056);
or U9616 (N_9616,N_9134,N_9457);
or U9617 (N_9617,N_9152,N_9353);
xnor U9618 (N_9618,N_9442,N_9101);
xnor U9619 (N_9619,N_9375,N_9405);
and U9620 (N_9620,N_9285,N_9419);
nor U9621 (N_9621,N_9298,N_9338);
nand U9622 (N_9622,N_9228,N_9300);
nand U9623 (N_9623,N_9039,N_9102);
nor U9624 (N_9624,N_9025,N_9406);
or U9625 (N_9625,N_9167,N_9479);
or U9626 (N_9626,N_9450,N_9087);
nor U9627 (N_9627,N_9395,N_9397);
or U9628 (N_9628,N_9319,N_9249);
nor U9629 (N_9629,N_9278,N_9333);
xnor U9630 (N_9630,N_9465,N_9247);
nor U9631 (N_9631,N_9306,N_9186);
xnor U9632 (N_9632,N_9142,N_9345);
nand U9633 (N_9633,N_9190,N_9355);
nand U9634 (N_9634,N_9401,N_9476);
nand U9635 (N_9635,N_9176,N_9162);
or U9636 (N_9636,N_9282,N_9497);
nand U9637 (N_9637,N_9236,N_9420);
nand U9638 (N_9638,N_9433,N_9407);
or U9639 (N_9639,N_9180,N_9158);
nand U9640 (N_9640,N_9344,N_9304);
and U9641 (N_9641,N_9346,N_9116);
or U9642 (N_9642,N_9322,N_9166);
nand U9643 (N_9643,N_9179,N_9226);
nand U9644 (N_9644,N_9185,N_9131);
xnor U9645 (N_9645,N_9361,N_9230);
or U9646 (N_9646,N_9314,N_9387);
xnor U9647 (N_9647,N_9060,N_9024);
and U9648 (N_9648,N_9124,N_9011);
nand U9649 (N_9649,N_9428,N_9082);
or U9650 (N_9650,N_9035,N_9109);
nand U9651 (N_9651,N_9267,N_9490);
or U9652 (N_9652,N_9194,N_9317);
and U9653 (N_9653,N_9164,N_9270);
xor U9654 (N_9654,N_9066,N_9006);
nand U9655 (N_9655,N_9431,N_9342);
xnor U9656 (N_9656,N_9474,N_9246);
and U9657 (N_9657,N_9098,N_9074);
nor U9658 (N_9658,N_9192,N_9414);
or U9659 (N_9659,N_9023,N_9293);
and U9660 (N_9660,N_9015,N_9061);
nand U9661 (N_9661,N_9292,N_9173);
and U9662 (N_9662,N_9221,N_9043);
and U9663 (N_9663,N_9008,N_9193);
nand U9664 (N_9664,N_9432,N_9094);
or U9665 (N_9665,N_9367,N_9117);
or U9666 (N_9666,N_9097,N_9469);
or U9667 (N_9667,N_9381,N_9071);
and U9668 (N_9668,N_9491,N_9235);
or U9669 (N_9669,N_9012,N_9416);
and U9670 (N_9670,N_9070,N_9328);
and U9671 (N_9671,N_9104,N_9000);
nand U9672 (N_9672,N_9049,N_9316);
and U9673 (N_9673,N_9286,N_9210);
nand U9674 (N_9674,N_9181,N_9449);
nor U9675 (N_9675,N_9385,N_9335);
nand U9676 (N_9676,N_9478,N_9275);
nand U9677 (N_9677,N_9423,N_9280);
nand U9678 (N_9678,N_9393,N_9323);
xor U9679 (N_9679,N_9095,N_9380);
or U9680 (N_9680,N_9044,N_9027);
nor U9681 (N_9681,N_9076,N_9441);
and U9682 (N_9682,N_9219,N_9435);
nor U9683 (N_9683,N_9373,N_9175);
nor U9684 (N_9684,N_9379,N_9081);
nor U9685 (N_9685,N_9240,N_9022);
and U9686 (N_9686,N_9412,N_9372);
and U9687 (N_9687,N_9302,N_9238);
xnor U9688 (N_9688,N_9461,N_9034);
xor U9689 (N_9689,N_9223,N_9325);
xnor U9690 (N_9690,N_9386,N_9205);
xnor U9691 (N_9691,N_9263,N_9418);
and U9692 (N_9692,N_9144,N_9075);
nor U9693 (N_9693,N_9470,N_9062);
nor U9694 (N_9694,N_9055,N_9260);
xor U9695 (N_9695,N_9054,N_9281);
nor U9696 (N_9696,N_9077,N_9107);
and U9697 (N_9697,N_9404,N_9187);
nand U9698 (N_9698,N_9009,N_9106);
nor U9699 (N_9699,N_9126,N_9147);
nand U9700 (N_9700,N_9154,N_9143);
nor U9701 (N_9701,N_9207,N_9259);
and U9702 (N_9702,N_9245,N_9130);
nor U9703 (N_9703,N_9439,N_9324);
or U9704 (N_9704,N_9169,N_9159);
nor U9705 (N_9705,N_9136,N_9118);
and U9706 (N_9706,N_9287,N_9160);
or U9707 (N_9707,N_9072,N_9307);
nand U9708 (N_9708,N_9417,N_9045);
or U9709 (N_9709,N_9115,N_9390);
xnor U9710 (N_9710,N_9222,N_9425);
xor U9711 (N_9711,N_9480,N_9211);
nor U9712 (N_9712,N_9455,N_9123);
nand U9713 (N_9713,N_9413,N_9430);
nand U9714 (N_9714,N_9437,N_9472);
nand U9715 (N_9715,N_9174,N_9125);
and U9716 (N_9716,N_9182,N_9396);
and U9717 (N_9717,N_9163,N_9331);
nor U9718 (N_9718,N_9498,N_9456);
xor U9719 (N_9719,N_9486,N_9019);
nor U9720 (N_9720,N_9215,N_9145);
and U9721 (N_9721,N_9178,N_9128);
nand U9722 (N_9722,N_9408,N_9100);
and U9723 (N_9723,N_9067,N_9308);
and U9724 (N_9724,N_9312,N_9048);
or U9725 (N_9725,N_9458,N_9447);
nand U9726 (N_9726,N_9225,N_9499);
xor U9727 (N_9727,N_9218,N_9451);
nand U9728 (N_9728,N_9002,N_9059);
or U9729 (N_9729,N_9197,N_9402);
nor U9730 (N_9730,N_9122,N_9311);
xnor U9731 (N_9731,N_9362,N_9242);
nor U9732 (N_9732,N_9475,N_9206);
nand U9733 (N_9733,N_9296,N_9073);
and U9734 (N_9734,N_9105,N_9153);
and U9735 (N_9735,N_9018,N_9146);
xor U9736 (N_9736,N_9085,N_9253);
xnor U9737 (N_9737,N_9003,N_9279);
or U9738 (N_9738,N_9352,N_9337);
nor U9739 (N_9739,N_9139,N_9321);
xnor U9740 (N_9740,N_9271,N_9496);
xor U9741 (N_9741,N_9080,N_9427);
xnor U9742 (N_9742,N_9341,N_9189);
nand U9743 (N_9743,N_9220,N_9485);
nor U9744 (N_9744,N_9155,N_9256);
xor U9745 (N_9745,N_9424,N_9046);
nor U9746 (N_9746,N_9013,N_9356);
nor U9747 (N_9747,N_9288,N_9482);
nand U9748 (N_9748,N_9429,N_9464);
xnor U9749 (N_9749,N_9398,N_9057);
and U9750 (N_9750,N_9128,N_9472);
or U9751 (N_9751,N_9150,N_9305);
nor U9752 (N_9752,N_9234,N_9061);
nand U9753 (N_9753,N_9302,N_9005);
and U9754 (N_9754,N_9363,N_9390);
nor U9755 (N_9755,N_9139,N_9387);
nor U9756 (N_9756,N_9298,N_9281);
nand U9757 (N_9757,N_9459,N_9407);
or U9758 (N_9758,N_9393,N_9225);
nand U9759 (N_9759,N_9285,N_9117);
or U9760 (N_9760,N_9340,N_9144);
nor U9761 (N_9761,N_9211,N_9338);
or U9762 (N_9762,N_9025,N_9447);
xor U9763 (N_9763,N_9188,N_9045);
nor U9764 (N_9764,N_9029,N_9222);
xnor U9765 (N_9765,N_9414,N_9165);
xor U9766 (N_9766,N_9043,N_9454);
or U9767 (N_9767,N_9172,N_9125);
and U9768 (N_9768,N_9316,N_9484);
xor U9769 (N_9769,N_9070,N_9148);
or U9770 (N_9770,N_9183,N_9042);
nand U9771 (N_9771,N_9221,N_9037);
xor U9772 (N_9772,N_9472,N_9416);
or U9773 (N_9773,N_9450,N_9339);
or U9774 (N_9774,N_9055,N_9128);
nor U9775 (N_9775,N_9018,N_9427);
xnor U9776 (N_9776,N_9156,N_9466);
or U9777 (N_9777,N_9132,N_9103);
nand U9778 (N_9778,N_9171,N_9390);
and U9779 (N_9779,N_9135,N_9486);
xnor U9780 (N_9780,N_9255,N_9466);
nor U9781 (N_9781,N_9252,N_9353);
and U9782 (N_9782,N_9458,N_9360);
nor U9783 (N_9783,N_9445,N_9223);
xnor U9784 (N_9784,N_9182,N_9194);
nor U9785 (N_9785,N_9246,N_9338);
nor U9786 (N_9786,N_9174,N_9117);
or U9787 (N_9787,N_9391,N_9396);
nor U9788 (N_9788,N_9038,N_9306);
nor U9789 (N_9789,N_9190,N_9375);
or U9790 (N_9790,N_9426,N_9412);
xnor U9791 (N_9791,N_9466,N_9021);
nor U9792 (N_9792,N_9420,N_9250);
nor U9793 (N_9793,N_9014,N_9340);
xnor U9794 (N_9794,N_9011,N_9342);
or U9795 (N_9795,N_9441,N_9379);
nor U9796 (N_9796,N_9355,N_9150);
xnor U9797 (N_9797,N_9417,N_9351);
or U9798 (N_9798,N_9218,N_9118);
and U9799 (N_9799,N_9186,N_9104);
and U9800 (N_9800,N_9299,N_9366);
nor U9801 (N_9801,N_9451,N_9309);
xor U9802 (N_9802,N_9368,N_9319);
nor U9803 (N_9803,N_9249,N_9449);
and U9804 (N_9804,N_9296,N_9093);
and U9805 (N_9805,N_9015,N_9183);
xor U9806 (N_9806,N_9158,N_9021);
and U9807 (N_9807,N_9317,N_9413);
xor U9808 (N_9808,N_9190,N_9171);
and U9809 (N_9809,N_9005,N_9131);
and U9810 (N_9810,N_9145,N_9375);
nor U9811 (N_9811,N_9469,N_9451);
and U9812 (N_9812,N_9455,N_9394);
and U9813 (N_9813,N_9046,N_9237);
or U9814 (N_9814,N_9102,N_9262);
nor U9815 (N_9815,N_9285,N_9443);
nor U9816 (N_9816,N_9333,N_9392);
nor U9817 (N_9817,N_9002,N_9021);
xor U9818 (N_9818,N_9236,N_9010);
and U9819 (N_9819,N_9436,N_9219);
nor U9820 (N_9820,N_9072,N_9026);
or U9821 (N_9821,N_9311,N_9279);
nor U9822 (N_9822,N_9188,N_9209);
xor U9823 (N_9823,N_9189,N_9117);
nand U9824 (N_9824,N_9037,N_9235);
nor U9825 (N_9825,N_9118,N_9074);
and U9826 (N_9826,N_9403,N_9200);
and U9827 (N_9827,N_9343,N_9127);
nand U9828 (N_9828,N_9356,N_9497);
and U9829 (N_9829,N_9275,N_9203);
nand U9830 (N_9830,N_9329,N_9182);
or U9831 (N_9831,N_9036,N_9372);
xor U9832 (N_9832,N_9260,N_9148);
and U9833 (N_9833,N_9415,N_9041);
and U9834 (N_9834,N_9253,N_9288);
and U9835 (N_9835,N_9386,N_9214);
xor U9836 (N_9836,N_9369,N_9497);
and U9837 (N_9837,N_9058,N_9443);
xnor U9838 (N_9838,N_9322,N_9027);
nand U9839 (N_9839,N_9072,N_9281);
xor U9840 (N_9840,N_9443,N_9212);
nor U9841 (N_9841,N_9301,N_9347);
and U9842 (N_9842,N_9067,N_9040);
nand U9843 (N_9843,N_9161,N_9344);
xnor U9844 (N_9844,N_9433,N_9074);
or U9845 (N_9845,N_9359,N_9179);
nor U9846 (N_9846,N_9365,N_9249);
nor U9847 (N_9847,N_9424,N_9237);
nor U9848 (N_9848,N_9145,N_9298);
and U9849 (N_9849,N_9299,N_9330);
or U9850 (N_9850,N_9465,N_9023);
and U9851 (N_9851,N_9431,N_9366);
xor U9852 (N_9852,N_9307,N_9230);
nand U9853 (N_9853,N_9389,N_9331);
or U9854 (N_9854,N_9342,N_9369);
xor U9855 (N_9855,N_9194,N_9325);
or U9856 (N_9856,N_9355,N_9103);
nand U9857 (N_9857,N_9432,N_9222);
nand U9858 (N_9858,N_9140,N_9327);
xnor U9859 (N_9859,N_9489,N_9210);
and U9860 (N_9860,N_9304,N_9254);
xnor U9861 (N_9861,N_9453,N_9363);
and U9862 (N_9862,N_9083,N_9010);
or U9863 (N_9863,N_9210,N_9202);
nor U9864 (N_9864,N_9056,N_9027);
nor U9865 (N_9865,N_9105,N_9420);
xnor U9866 (N_9866,N_9099,N_9261);
nand U9867 (N_9867,N_9376,N_9097);
nor U9868 (N_9868,N_9219,N_9261);
xor U9869 (N_9869,N_9425,N_9008);
nor U9870 (N_9870,N_9184,N_9315);
nand U9871 (N_9871,N_9387,N_9411);
and U9872 (N_9872,N_9318,N_9323);
nand U9873 (N_9873,N_9067,N_9005);
xor U9874 (N_9874,N_9321,N_9137);
nand U9875 (N_9875,N_9223,N_9294);
and U9876 (N_9876,N_9459,N_9153);
or U9877 (N_9877,N_9283,N_9479);
or U9878 (N_9878,N_9125,N_9045);
nor U9879 (N_9879,N_9356,N_9091);
nor U9880 (N_9880,N_9007,N_9025);
nand U9881 (N_9881,N_9473,N_9192);
nand U9882 (N_9882,N_9249,N_9068);
nand U9883 (N_9883,N_9226,N_9136);
xor U9884 (N_9884,N_9398,N_9328);
nand U9885 (N_9885,N_9488,N_9058);
or U9886 (N_9886,N_9283,N_9074);
nor U9887 (N_9887,N_9226,N_9324);
or U9888 (N_9888,N_9441,N_9480);
and U9889 (N_9889,N_9325,N_9061);
nand U9890 (N_9890,N_9479,N_9102);
nand U9891 (N_9891,N_9451,N_9086);
nor U9892 (N_9892,N_9089,N_9029);
nand U9893 (N_9893,N_9438,N_9383);
and U9894 (N_9894,N_9077,N_9491);
or U9895 (N_9895,N_9190,N_9391);
nand U9896 (N_9896,N_9182,N_9332);
and U9897 (N_9897,N_9455,N_9047);
and U9898 (N_9898,N_9198,N_9459);
or U9899 (N_9899,N_9316,N_9414);
and U9900 (N_9900,N_9359,N_9453);
and U9901 (N_9901,N_9331,N_9114);
or U9902 (N_9902,N_9295,N_9192);
nand U9903 (N_9903,N_9145,N_9437);
nand U9904 (N_9904,N_9141,N_9009);
xnor U9905 (N_9905,N_9417,N_9151);
and U9906 (N_9906,N_9175,N_9363);
and U9907 (N_9907,N_9184,N_9121);
xnor U9908 (N_9908,N_9093,N_9082);
and U9909 (N_9909,N_9128,N_9493);
and U9910 (N_9910,N_9011,N_9256);
nor U9911 (N_9911,N_9337,N_9267);
nand U9912 (N_9912,N_9132,N_9171);
or U9913 (N_9913,N_9479,N_9279);
or U9914 (N_9914,N_9105,N_9341);
or U9915 (N_9915,N_9397,N_9321);
or U9916 (N_9916,N_9322,N_9126);
nand U9917 (N_9917,N_9274,N_9499);
nand U9918 (N_9918,N_9478,N_9018);
or U9919 (N_9919,N_9013,N_9399);
xor U9920 (N_9920,N_9428,N_9169);
nor U9921 (N_9921,N_9059,N_9307);
or U9922 (N_9922,N_9273,N_9217);
or U9923 (N_9923,N_9481,N_9093);
or U9924 (N_9924,N_9415,N_9295);
or U9925 (N_9925,N_9382,N_9380);
nor U9926 (N_9926,N_9356,N_9180);
or U9927 (N_9927,N_9113,N_9309);
or U9928 (N_9928,N_9221,N_9250);
and U9929 (N_9929,N_9453,N_9388);
nand U9930 (N_9930,N_9019,N_9136);
nand U9931 (N_9931,N_9110,N_9307);
or U9932 (N_9932,N_9176,N_9051);
xnor U9933 (N_9933,N_9004,N_9297);
xnor U9934 (N_9934,N_9047,N_9428);
nor U9935 (N_9935,N_9060,N_9369);
nand U9936 (N_9936,N_9148,N_9394);
xor U9937 (N_9937,N_9054,N_9192);
nor U9938 (N_9938,N_9009,N_9202);
nor U9939 (N_9939,N_9371,N_9330);
nand U9940 (N_9940,N_9281,N_9238);
nor U9941 (N_9941,N_9383,N_9333);
or U9942 (N_9942,N_9360,N_9044);
nor U9943 (N_9943,N_9035,N_9166);
or U9944 (N_9944,N_9338,N_9072);
and U9945 (N_9945,N_9109,N_9413);
and U9946 (N_9946,N_9121,N_9307);
or U9947 (N_9947,N_9301,N_9242);
nand U9948 (N_9948,N_9486,N_9148);
nand U9949 (N_9949,N_9174,N_9047);
xnor U9950 (N_9950,N_9247,N_9402);
and U9951 (N_9951,N_9112,N_9468);
nand U9952 (N_9952,N_9128,N_9365);
and U9953 (N_9953,N_9415,N_9366);
xnor U9954 (N_9954,N_9095,N_9353);
nand U9955 (N_9955,N_9371,N_9286);
or U9956 (N_9956,N_9180,N_9288);
xor U9957 (N_9957,N_9126,N_9380);
xnor U9958 (N_9958,N_9483,N_9314);
nor U9959 (N_9959,N_9061,N_9226);
nor U9960 (N_9960,N_9270,N_9272);
or U9961 (N_9961,N_9271,N_9067);
nor U9962 (N_9962,N_9488,N_9178);
and U9963 (N_9963,N_9071,N_9485);
and U9964 (N_9964,N_9371,N_9353);
xnor U9965 (N_9965,N_9125,N_9348);
nor U9966 (N_9966,N_9178,N_9464);
nand U9967 (N_9967,N_9091,N_9113);
nand U9968 (N_9968,N_9253,N_9116);
xnor U9969 (N_9969,N_9406,N_9150);
nand U9970 (N_9970,N_9132,N_9142);
nor U9971 (N_9971,N_9092,N_9093);
or U9972 (N_9972,N_9116,N_9322);
xor U9973 (N_9973,N_9315,N_9293);
and U9974 (N_9974,N_9486,N_9370);
nor U9975 (N_9975,N_9020,N_9484);
nand U9976 (N_9976,N_9475,N_9254);
or U9977 (N_9977,N_9081,N_9288);
nand U9978 (N_9978,N_9496,N_9365);
nor U9979 (N_9979,N_9125,N_9211);
and U9980 (N_9980,N_9042,N_9029);
or U9981 (N_9981,N_9146,N_9304);
or U9982 (N_9982,N_9157,N_9195);
nand U9983 (N_9983,N_9462,N_9434);
or U9984 (N_9984,N_9422,N_9177);
and U9985 (N_9985,N_9494,N_9174);
nor U9986 (N_9986,N_9417,N_9222);
and U9987 (N_9987,N_9282,N_9307);
nand U9988 (N_9988,N_9025,N_9146);
nor U9989 (N_9989,N_9351,N_9451);
or U9990 (N_9990,N_9150,N_9374);
xnor U9991 (N_9991,N_9376,N_9113);
xnor U9992 (N_9992,N_9145,N_9399);
or U9993 (N_9993,N_9405,N_9295);
or U9994 (N_9994,N_9119,N_9287);
nor U9995 (N_9995,N_9374,N_9316);
and U9996 (N_9996,N_9215,N_9321);
xor U9997 (N_9997,N_9402,N_9397);
nand U9998 (N_9998,N_9463,N_9189);
nand U9999 (N_9999,N_9331,N_9253);
nand UO_0 (O_0,N_9876,N_9608);
nand UO_1 (O_1,N_9503,N_9640);
nand UO_2 (O_2,N_9552,N_9538);
nand UO_3 (O_3,N_9953,N_9964);
and UO_4 (O_4,N_9705,N_9978);
xor UO_5 (O_5,N_9906,N_9872);
or UO_6 (O_6,N_9923,N_9899);
and UO_7 (O_7,N_9821,N_9860);
and UO_8 (O_8,N_9534,N_9992);
and UO_9 (O_9,N_9908,N_9516);
and UO_10 (O_10,N_9549,N_9502);
nor UO_11 (O_11,N_9930,N_9863);
nor UO_12 (O_12,N_9514,N_9556);
nor UO_13 (O_13,N_9785,N_9706);
nor UO_14 (O_14,N_9691,N_9629);
and UO_15 (O_15,N_9825,N_9735);
nor UO_16 (O_16,N_9717,N_9671);
or UO_17 (O_17,N_9797,N_9852);
nor UO_18 (O_18,N_9985,N_9827);
nor UO_19 (O_19,N_9975,N_9854);
or UO_20 (O_20,N_9960,N_9998);
and UO_21 (O_21,N_9783,N_9886);
xnor UO_22 (O_22,N_9989,N_9972);
xor UO_23 (O_23,N_9774,N_9840);
xor UO_24 (O_24,N_9553,N_9926);
nor UO_25 (O_25,N_9532,N_9941);
or UO_26 (O_26,N_9823,N_9855);
or UO_27 (O_27,N_9733,N_9858);
xor UO_28 (O_28,N_9834,N_9955);
nand UO_29 (O_29,N_9787,N_9995);
xor UO_30 (O_30,N_9635,N_9766);
xor UO_31 (O_31,N_9660,N_9742);
xor UO_32 (O_32,N_9842,N_9835);
nand UO_33 (O_33,N_9965,N_9518);
and UO_34 (O_34,N_9830,N_9554);
nor UO_35 (O_35,N_9524,N_9589);
nand UO_36 (O_36,N_9611,N_9818);
nand UO_37 (O_37,N_9548,N_9946);
or UO_38 (O_38,N_9604,N_9632);
or UO_39 (O_39,N_9619,N_9509);
or UO_40 (O_40,N_9932,N_9974);
or UO_41 (O_41,N_9719,N_9716);
nor UO_42 (O_42,N_9557,N_9994);
nor UO_43 (O_43,N_9723,N_9663);
xnor UO_44 (O_44,N_9674,N_9727);
nor UO_45 (O_45,N_9833,N_9748);
nor UO_46 (O_46,N_9555,N_9734);
nand UO_47 (O_47,N_9544,N_9917);
xnor UO_48 (O_48,N_9836,N_9507);
or UO_49 (O_49,N_9884,N_9869);
xor UO_50 (O_50,N_9857,N_9798);
and UO_51 (O_51,N_9637,N_9696);
xnor UO_52 (O_52,N_9636,N_9607);
and UO_53 (O_53,N_9982,N_9689);
xor UO_54 (O_54,N_9758,N_9750);
nand UO_55 (O_55,N_9943,N_9971);
xor UO_56 (O_56,N_9988,N_9618);
or UO_57 (O_57,N_9990,N_9800);
and UO_58 (O_58,N_9897,N_9997);
xnor UO_59 (O_59,N_9596,N_9668);
nor UO_60 (O_60,N_9752,N_9692);
nor UO_61 (O_61,N_9657,N_9769);
nor UO_62 (O_62,N_9676,N_9909);
and UO_63 (O_63,N_9747,N_9599);
or UO_64 (O_64,N_9642,N_9968);
or UO_65 (O_65,N_9952,N_9796);
and UO_66 (O_66,N_9583,N_9927);
xnor UO_67 (O_67,N_9763,N_9710);
or UO_68 (O_68,N_9581,N_9738);
or UO_69 (O_69,N_9933,N_9715);
and UO_70 (O_70,N_9614,N_9900);
nor UO_71 (O_71,N_9849,N_9693);
xnor UO_72 (O_72,N_9594,N_9725);
nand UO_73 (O_73,N_9891,N_9510);
or UO_74 (O_74,N_9648,N_9513);
and UO_75 (O_75,N_9537,N_9741);
xor UO_76 (O_76,N_9838,N_9853);
nand UO_77 (O_77,N_9517,N_9799);
nand UO_78 (O_78,N_9812,N_9625);
nor UO_79 (O_79,N_9770,N_9981);
nand UO_80 (O_80,N_9907,N_9686);
nor UO_81 (O_81,N_9786,N_9760);
nor UO_82 (O_82,N_9714,N_9874);
xnor UO_83 (O_83,N_9695,N_9568);
or UO_84 (O_84,N_9675,N_9948);
or UO_85 (O_85,N_9720,N_9832);
xor UO_86 (O_86,N_9814,N_9862);
or UO_87 (O_87,N_9605,N_9877);
xor UO_88 (O_88,N_9947,N_9672);
nand UO_89 (O_89,N_9579,N_9788);
xnor UO_90 (O_90,N_9662,N_9993);
xnor UO_91 (O_91,N_9646,N_9570);
nand UO_92 (O_92,N_9564,N_9745);
and UO_93 (O_93,N_9757,N_9655);
or UO_94 (O_94,N_9687,N_9681);
nand UO_95 (O_95,N_9688,N_9973);
nor UO_96 (O_96,N_9651,N_9620);
or UO_97 (O_97,N_9664,N_9624);
xnor UO_98 (O_98,N_9970,N_9639);
or UO_99 (O_99,N_9937,N_9977);
nand UO_100 (O_100,N_9574,N_9569);
xnor UO_101 (O_101,N_9580,N_9837);
nor UO_102 (O_102,N_9918,N_9819);
and UO_103 (O_103,N_9638,N_9698);
nor UO_104 (O_104,N_9744,N_9813);
xor UO_105 (O_105,N_9844,N_9916);
and UO_106 (O_106,N_9784,N_9794);
xor UO_107 (O_107,N_9966,N_9703);
nor UO_108 (O_108,N_9694,N_9575);
or UO_109 (O_109,N_9729,N_9606);
and UO_110 (O_110,N_9567,N_9896);
or UO_111 (O_111,N_9913,N_9914);
nand UO_112 (O_112,N_9983,N_9885);
xnor UO_113 (O_113,N_9929,N_9540);
nor UO_114 (O_114,N_9811,N_9724);
xor UO_115 (O_115,N_9616,N_9631);
xnor UO_116 (O_116,N_9561,N_9820);
or UO_117 (O_117,N_9803,N_9846);
or UO_118 (O_118,N_9609,N_9805);
xnor UO_119 (O_119,N_9709,N_9936);
nand UO_120 (O_120,N_9793,N_9904);
nand UO_121 (O_121,N_9559,N_9573);
or UO_122 (O_122,N_9673,N_9515);
nand UO_123 (O_123,N_9626,N_9740);
nor UO_124 (O_124,N_9654,N_9707);
or UO_125 (O_125,N_9647,N_9791);
nand UO_126 (O_126,N_9759,N_9521);
xnor UO_127 (O_127,N_9508,N_9731);
nor UO_128 (O_128,N_9684,N_9963);
and UO_129 (O_129,N_9721,N_9590);
nand UO_130 (O_130,N_9895,N_9523);
nor UO_131 (O_131,N_9547,N_9817);
nand UO_132 (O_132,N_9644,N_9781);
nand UO_133 (O_133,N_9653,N_9905);
nand UO_134 (O_134,N_9597,N_9887);
or UO_135 (O_135,N_9584,N_9856);
nor UO_136 (O_136,N_9749,N_9519);
or UO_137 (O_137,N_9980,N_9789);
or UO_138 (O_138,N_9652,N_9746);
or UO_139 (O_139,N_9969,N_9630);
or UO_140 (O_140,N_9822,N_9951);
nor UO_141 (O_141,N_9870,N_9586);
and UO_142 (O_142,N_9627,N_9726);
or UO_143 (O_143,N_9677,N_9950);
nand UO_144 (O_144,N_9685,N_9882);
xor UO_145 (O_145,N_9615,N_9773);
nand UO_146 (O_146,N_9683,N_9595);
nor UO_147 (O_147,N_9839,N_9621);
nand UO_148 (O_148,N_9542,N_9713);
or UO_149 (O_149,N_9712,N_9530);
xnor UO_150 (O_150,N_9535,N_9984);
or UO_151 (O_151,N_9563,N_9865);
and UO_152 (O_152,N_9986,N_9945);
xnor UO_153 (O_153,N_9831,N_9949);
xnor UO_154 (O_154,N_9679,N_9602);
xor UO_155 (O_155,N_9778,N_9711);
or UO_156 (O_156,N_9610,N_9566);
or UO_157 (O_157,N_9591,N_9987);
xor UO_158 (O_158,N_9873,N_9767);
nor UO_159 (O_159,N_9967,N_9658);
xnor UO_160 (O_160,N_9804,N_9828);
or UO_161 (O_161,N_9560,N_9558);
and UO_162 (O_162,N_9529,N_9919);
nor UO_163 (O_163,N_9824,N_9961);
xor UO_164 (O_164,N_9957,N_9976);
or UO_165 (O_165,N_9940,N_9931);
xnor UO_166 (O_166,N_9866,N_9565);
nand UO_167 (O_167,N_9925,N_9622);
nand UO_168 (O_168,N_9780,N_9768);
nand UO_169 (O_169,N_9843,N_9600);
and UO_170 (O_170,N_9765,N_9643);
xnor UO_171 (O_171,N_9939,N_9847);
and UO_172 (O_172,N_9612,N_9576);
nor UO_173 (O_173,N_9779,N_9861);
nand UO_174 (O_174,N_9934,N_9718);
and UO_175 (O_175,N_9649,N_9875);
nor UO_176 (O_176,N_9991,N_9522);
and UO_177 (O_177,N_9903,N_9678);
nand UO_178 (O_178,N_9525,N_9942);
nand UO_179 (O_179,N_9572,N_9809);
xnor UO_180 (O_180,N_9901,N_9506);
xor UO_181 (O_181,N_9656,N_9603);
xnor UO_182 (O_182,N_9730,N_9808);
xor UO_183 (O_183,N_9880,N_9928);
xnor UO_184 (O_184,N_9736,N_9665);
and UO_185 (O_185,N_9708,N_9511);
xnor UO_186 (O_186,N_9815,N_9902);
and UO_187 (O_187,N_9645,N_9910);
xnor UO_188 (O_188,N_9772,N_9859);
nand UO_189 (O_189,N_9776,N_9743);
and UO_190 (O_190,N_9697,N_9500);
nor UO_191 (O_191,N_9699,N_9753);
and UO_192 (O_192,N_9898,N_9527);
nand UO_193 (O_193,N_9883,N_9935);
and UO_194 (O_194,N_9578,N_9889);
nor UO_195 (O_195,N_9871,N_9915);
and UO_196 (O_196,N_9571,N_9944);
nor UO_197 (O_197,N_9911,N_9617);
xnor UO_198 (O_198,N_9501,N_9546);
nand UO_199 (O_199,N_9520,N_9661);
nand UO_200 (O_200,N_9878,N_9690);
or UO_201 (O_201,N_9641,N_9867);
and UO_202 (O_202,N_9881,N_9539);
xnor UO_203 (O_203,N_9938,N_9585);
and UO_204 (O_204,N_9533,N_9806);
and UO_205 (O_205,N_9958,N_9890);
and UO_206 (O_206,N_9623,N_9762);
or UO_207 (O_207,N_9962,N_9782);
nand UO_208 (O_208,N_9894,N_9634);
and UO_209 (O_209,N_9528,N_9761);
or UO_210 (O_210,N_9737,N_9551);
nand UO_211 (O_211,N_9924,N_9667);
nor UO_212 (O_212,N_9826,N_9577);
and UO_213 (O_213,N_9956,N_9841);
xnor UO_214 (O_214,N_9739,N_9601);
nand UO_215 (O_215,N_9893,N_9979);
xor UO_216 (O_216,N_9864,N_9751);
or UO_217 (O_217,N_9764,N_9848);
nor UO_218 (O_218,N_9562,N_9816);
or UO_219 (O_219,N_9732,N_9587);
nand UO_220 (O_220,N_9543,N_9659);
nand UO_221 (O_221,N_9633,N_9996);
and UO_222 (O_222,N_9845,N_9670);
xor UO_223 (O_223,N_9504,N_9920);
and UO_224 (O_224,N_9531,N_9851);
or UO_225 (O_225,N_9505,N_9722);
nand UO_226 (O_226,N_9628,N_9650);
nand UO_227 (O_227,N_9755,N_9582);
and UO_228 (O_228,N_9702,N_9545);
and UO_229 (O_229,N_9512,N_9704);
xor UO_230 (O_230,N_9810,N_9954);
or UO_231 (O_231,N_9593,N_9892);
nand UO_232 (O_232,N_9728,N_9802);
and UO_233 (O_233,N_9888,N_9795);
nor UO_234 (O_234,N_9775,N_9868);
or UO_235 (O_235,N_9526,N_9613);
or UO_236 (O_236,N_9598,N_9680);
xor UO_237 (O_237,N_9700,N_9754);
xor UO_238 (O_238,N_9588,N_9912);
nor UO_239 (O_239,N_9536,N_9550);
or UO_240 (O_240,N_9959,N_9771);
and UO_241 (O_241,N_9592,N_9756);
nor UO_242 (O_242,N_9541,N_9701);
and UO_243 (O_243,N_9682,N_9850);
or UO_244 (O_244,N_9669,N_9807);
nand UO_245 (O_245,N_9829,N_9999);
and UO_246 (O_246,N_9777,N_9879);
nor UO_247 (O_247,N_9666,N_9792);
xor UO_248 (O_248,N_9922,N_9801);
nand UO_249 (O_249,N_9790,N_9921);
or UO_250 (O_250,N_9962,N_9606);
and UO_251 (O_251,N_9635,N_9717);
nand UO_252 (O_252,N_9757,N_9628);
nor UO_253 (O_253,N_9603,N_9997);
nand UO_254 (O_254,N_9978,N_9766);
and UO_255 (O_255,N_9610,N_9797);
or UO_256 (O_256,N_9793,N_9907);
nor UO_257 (O_257,N_9583,N_9519);
or UO_258 (O_258,N_9824,N_9745);
nor UO_259 (O_259,N_9647,N_9719);
or UO_260 (O_260,N_9804,N_9765);
and UO_261 (O_261,N_9565,N_9620);
nor UO_262 (O_262,N_9520,N_9896);
nand UO_263 (O_263,N_9862,N_9603);
or UO_264 (O_264,N_9640,N_9518);
xnor UO_265 (O_265,N_9717,N_9689);
nor UO_266 (O_266,N_9752,N_9926);
and UO_267 (O_267,N_9651,N_9608);
xor UO_268 (O_268,N_9722,N_9699);
or UO_269 (O_269,N_9616,N_9856);
xor UO_270 (O_270,N_9539,N_9601);
and UO_271 (O_271,N_9971,N_9816);
xnor UO_272 (O_272,N_9950,N_9923);
and UO_273 (O_273,N_9660,N_9913);
or UO_274 (O_274,N_9972,N_9638);
nor UO_275 (O_275,N_9684,N_9663);
nand UO_276 (O_276,N_9672,N_9525);
nand UO_277 (O_277,N_9602,N_9800);
xnor UO_278 (O_278,N_9874,N_9817);
nand UO_279 (O_279,N_9620,N_9882);
nand UO_280 (O_280,N_9537,N_9795);
nor UO_281 (O_281,N_9785,N_9868);
xnor UO_282 (O_282,N_9633,N_9577);
and UO_283 (O_283,N_9587,N_9749);
and UO_284 (O_284,N_9900,N_9564);
xor UO_285 (O_285,N_9976,N_9764);
nand UO_286 (O_286,N_9919,N_9521);
and UO_287 (O_287,N_9685,N_9638);
xnor UO_288 (O_288,N_9948,N_9970);
and UO_289 (O_289,N_9694,N_9730);
or UO_290 (O_290,N_9545,N_9975);
nor UO_291 (O_291,N_9769,N_9870);
or UO_292 (O_292,N_9549,N_9548);
and UO_293 (O_293,N_9917,N_9740);
or UO_294 (O_294,N_9961,N_9529);
and UO_295 (O_295,N_9970,N_9887);
nand UO_296 (O_296,N_9866,N_9574);
or UO_297 (O_297,N_9567,N_9645);
xor UO_298 (O_298,N_9841,N_9711);
and UO_299 (O_299,N_9760,N_9837);
nand UO_300 (O_300,N_9600,N_9896);
and UO_301 (O_301,N_9850,N_9695);
nand UO_302 (O_302,N_9764,N_9855);
and UO_303 (O_303,N_9590,N_9718);
xor UO_304 (O_304,N_9976,N_9863);
nand UO_305 (O_305,N_9889,N_9613);
nand UO_306 (O_306,N_9876,N_9801);
xor UO_307 (O_307,N_9653,N_9930);
or UO_308 (O_308,N_9876,N_9701);
or UO_309 (O_309,N_9541,N_9522);
nand UO_310 (O_310,N_9690,N_9756);
xor UO_311 (O_311,N_9875,N_9660);
xor UO_312 (O_312,N_9757,N_9588);
nor UO_313 (O_313,N_9687,N_9696);
nand UO_314 (O_314,N_9657,N_9876);
or UO_315 (O_315,N_9628,N_9752);
nand UO_316 (O_316,N_9967,N_9612);
xnor UO_317 (O_317,N_9741,N_9934);
xnor UO_318 (O_318,N_9723,N_9739);
nor UO_319 (O_319,N_9582,N_9828);
xor UO_320 (O_320,N_9628,N_9685);
and UO_321 (O_321,N_9863,N_9754);
xor UO_322 (O_322,N_9688,N_9676);
xor UO_323 (O_323,N_9837,N_9868);
or UO_324 (O_324,N_9698,N_9872);
or UO_325 (O_325,N_9500,N_9680);
xor UO_326 (O_326,N_9854,N_9545);
or UO_327 (O_327,N_9528,N_9987);
or UO_328 (O_328,N_9599,N_9798);
nand UO_329 (O_329,N_9698,N_9857);
nor UO_330 (O_330,N_9905,N_9890);
xnor UO_331 (O_331,N_9650,N_9883);
nand UO_332 (O_332,N_9651,N_9614);
nor UO_333 (O_333,N_9543,N_9711);
and UO_334 (O_334,N_9850,N_9556);
nor UO_335 (O_335,N_9663,N_9549);
or UO_336 (O_336,N_9981,N_9729);
nor UO_337 (O_337,N_9959,N_9762);
nor UO_338 (O_338,N_9855,N_9684);
xor UO_339 (O_339,N_9883,N_9965);
xnor UO_340 (O_340,N_9891,N_9888);
nor UO_341 (O_341,N_9701,N_9838);
nand UO_342 (O_342,N_9601,N_9782);
nand UO_343 (O_343,N_9888,N_9556);
nand UO_344 (O_344,N_9538,N_9800);
nor UO_345 (O_345,N_9839,N_9693);
nand UO_346 (O_346,N_9882,N_9674);
nand UO_347 (O_347,N_9708,N_9784);
nand UO_348 (O_348,N_9907,N_9512);
xnor UO_349 (O_349,N_9713,N_9902);
nand UO_350 (O_350,N_9914,N_9902);
nor UO_351 (O_351,N_9694,N_9563);
or UO_352 (O_352,N_9603,N_9598);
and UO_353 (O_353,N_9708,N_9599);
xnor UO_354 (O_354,N_9769,N_9512);
and UO_355 (O_355,N_9883,N_9904);
xor UO_356 (O_356,N_9648,N_9909);
and UO_357 (O_357,N_9533,N_9668);
and UO_358 (O_358,N_9603,N_9925);
and UO_359 (O_359,N_9796,N_9788);
xnor UO_360 (O_360,N_9800,N_9796);
xor UO_361 (O_361,N_9685,N_9719);
xor UO_362 (O_362,N_9703,N_9871);
nor UO_363 (O_363,N_9997,N_9983);
nand UO_364 (O_364,N_9995,N_9728);
nand UO_365 (O_365,N_9534,N_9649);
nor UO_366 (O_366,N_9562,N_9744);
nand UO_367 (O_367,N_9657,N_9641);
xnor UO_368 (O_368,N_9864,N_9789);
nor UO_369 (O_369,N_9758,N_9565);
and UO_370 (O_370,N_9661,N_9685);
nor UO_371 (O_371,N_9800,N_9572);
or UO_372 (O_372,N_9724,N_9658);
or UO_373 (O_373,N_9799,N_9975);
and UO_374 (O_374,N_9979,N_9831);
nand UO_375 (O_375,N_9830,N_9993);
xnor UO_376 (O_376,N_9841,N_9796);
xor UO_377 (O_377,N_9592,N_9704);
xor UO_378 (O_378,N_9787,N_9923);
nor UO_379 (O_379,N_9519,N_9719);
nand UO_380 (O_380,N_9657,N_9623);
nor UO_381 (O_381,N_9751,N_9579);
or UO_382 (O_382,N_9541,N_9864);
xor UO_383 (O_383,N_9948,N_9632);
or UO_384 (O_384,N_9605,N_9572);
nand UO_385 (O_385,N_9617,N_9629);
or UO_386 (O_386,N_9606,N_9827);
nand UO_387 (O_387,N_9601,N_9617);
and UO_388 (O_388,N_9512,N_9726);
and UO_389 (O_389,N_9892,N_9880);
or UO_390 (O_390,N_9922,N_9662);
xor UO_391 (O_391,N_9809,N_9984);
nor UO_392 (O_392,N_9627,N_9811);
and UO_393 (O_393,N_9619,N_9839);
or UO_394 (O_394,N_9980,N_9993);
nor UO_395 (O_395,N_9687,N_9593);
and UO_396 (O_396,N_9954,N_9908);
xor UO_397 (O_397,N_9814,N_9750);
nand UO_398 (O_398,N_9577,N_9902);
or UO_399 (O_399,N_9947,N_9520);
nor UO_400 (O_400,N_9962,N_9890);
or UO_401 (O_401,N_9857,N_9889);
or UO_402 (O_402,N_9882,N_9932);
and UO_403 (O_403,N_9981,N_9831);
xnor UO_404 (O_404,N_9518,N_9738);
or UO_405 (O_405,N_9603,N_9629);
and UO_406 (O_406,N_9824,N_9559);
and UO_407 (O_407,N_9850,N_9559);
and UO_408 (O_408,N_9541,N_9943);
and UO_409 (O_409,N_9573,N_9851);
and UO_410 (O_410,N_9825,N_9952);
nor UO_411 (O_411,N_9736,N_9530);
or UO_412 (O_412,N_9731,N_9885);
or UO_413 (O_413,N_9918,N_9925);
nand UO_414 (O_414,N_9580,N_9785);
nand UO_415 (O_415,N_9974,N_9625);
and UO_416 (O_416,N_9890,N_9861);
nand UO_417 (O_417,N_9721,N_9509);
xor UO_418 (O_418,N_9940,N_9848);
nand UO_419 (O_419,N_9724,N_9733);
and UO_420 (O_420,N_9817,N_9919);
nand UO_421 (O_421,N_9701,N_9763);
and UO_422 (O_422,N_9637,N_9742);
xnor UO_423 (O_423,N_9832,N_9674);
or UO_424 (O_424,N_9848,N_9504);
nand UO_425 (O_425,N_9556,N_9934);
xor UO_426 (O_426,N_9649,N_9972);
and UO_427 (O_427,N_9706,N_9725);
nor UO_428 (O_428,N_9716,N_9705);
nor UO_429 (O_429,N_9508,N_9648);
xor UO_430 (O_430,N_9789,N_9988);
and UO_431 (O_431,N_9728,N_9733);
or UO_432 (O_432,N_9806,N_9911);
or UO_433 (O_433,N_9776,N_9553);
and UO_434 (O_434,N_9595,N_9824);
nor UO_435 (O_435,N_9660,N_9600);
xnor UO_436 (O_436,N_9830,N_9680);
nor UO_437 (O_437,N_9733,N_9575);
and UO_438 (O_438,N_9780,N_9651);
nor UO_439 (O_439,N_9738,N_9517);
or UO_440 (O_440,N_9603,N_9538);
nor UO_441 (O_441,N_9620,N_9563);
nand UO_442 (O_442,N_9995,N_9556);
nor UO_443 (O_443,N_9561,N_9797);
nand UO_444 (O_444,N_9752,N_9718);
nand UO_445 (O_445,N_9711,N_9820);
nand UO_446 (O_446,N_9974,N_9857);
nor UO_447 (O_447,N_9701,N_9601);
or UO_448 (O_448,N_9749,N_9811);
nor UO_449 (O_449,N_9679,N_9645);
xor UO_450 (O_450,N_9643,N_9842);
nand UO_451 (O_451,N_9551,N_9560);
nor UO_452 (O_452,N_9689,N_9522);
nand UO_453 (O_453,N_9755,N_9694);
or UO_454 (O_454,N_9689,N_9651);
or UO_455 (O_455,N_9588,N_9994);
and UO_456 (O_456,N_9866,N_9579);
nor UO_457 (O_457,N_9751,N_9542);
and UO_458 (O_458,N_9774,N_9936);
or UO_459 (O_459,N_9527,N_9772);
and UO_460 (O_460,N_9820,N_9661);
xor UO_461 (O_461,N_9974,N_9767);
nor UO_462 (O_462,N_9980,N_9813);
nor UO_463 (O_463,N_9759,N_9679);
and UO_464 (O_464,N_9977,N_9637);
or UO_465 (O_465,N_9790,N_9957);
and UO_466 (O_466,N_9586,N_9670);
or UO_467 (O_467,N_9929,N_9839);
or UO_468 (O_468,N_9532,N_9590);
and UO_469 (O_469,N_9746,N_9700);
nand UO_470 (O_470,N_9654,N_9591);
or UO_471 (O_471,N_9676,N_9622);
nor UO_472 (O_472,N_9533,N_9509);
and UO_473 (O_473,N_9978,N_9558);
nor UO_474 (O_474,N_9890,N_9920);
or UO_475 (O_475,N_9549,N_9807);
nor UO_476 (O_476,N_9976,N_9806);
or UO_477 (O_477,N_9783,N_9847);
and UO_478 (O_478,N_9791,N_9752);
and UO_479 (O_479,N_9902,N_9777);
xnor UO_480 (O_480,N_9960,N_9500);
xor UO_481 (O_481,N_9609,N_9811);
nand UO_482 (O_482,N_9810,N_9875);
xnor UO_483 (O_483,N_9602,N_9902);
nand UO_484 (O_484,N_9962,N_9916);
or UO_485 (O_485,N_9930,N_9635);
nor UO_486 (O_486,N_9954,N_9500);
nand UO_487 (O_487,N_9975,N_9752);
or UO_488 (O_488,N_9722,N_9972);
or UO_489 (O_489,N_9891,N_9850);
and UO_490 (O_490,N_9844,N_9563);
xor UO_491 (O_491,N_9557,N_9824);
nor UO_492 (O_492,N_9711,N_9800);
nand UO_493 (O_493,N_9968,N_9702);
and UO_494 (O_494,N_9761,N_9783);
xor UO_495 (O_495,N_9784,N_9894);
and UO_496 (O_496,N_9574,N_9770);
and UO_497 (O_497,N_9816,N_9833);
xnor UO_498 (O_498,N_9955,N_9848);
and UO_499 (O_499,N_9510,N_9650);
nand UO_500 (O_500,N_9618,N_9887);
or UO_501 (O_501,N_9717,N_9757);
nand UO_502 (O_502,N_9823,N_9913);
nand UO_503 (O_503,N_9720,N_9993);
or UO_504 (O_504,N_9792,N_9734);
xor UO_505 (O_505,N_9810,N_9752);
nand UO_506 (O_506,N_9783,N_9564);
or UO_507 (O_507,N_9863,N_9740);
nor UO_508 (O_508,N_9953,N_9548);
or UO_509 (O_509,N_9506,N_9530);
nand UO_510 (O_510,N_9783,N_9546);
nand UO_511 (O_511,N_9929,N_9740);
or UO_512 (O_512,N_9897,N_9657);
and UO_513 (O_513,N_9517,N_9505);
nor UO_514 (O_514,N_9972,N_9724);
nand UO_515 (O_515,N_9986,N_9753);
and UO_516 (O_516,N_9956,N_9722);
xor UO_517 (O_517,N_9632,N_9564);
and UO_518 (O_518,N_9695,N_9936);
xnor UO_519 (O_519,N_9916,N_9932);
and UO_520 (O_520,N_9967,N_9762);
and UO_521 (O_521,N_9641,N_9905);
and UO_522 (O_522,N_9655,N_9921);
xor UO_523 (O_523,N_9648,N_9986);
or UO_524 (O_524,N_9627,N_9997);
xnor UO_525 (O_525,N_9718,N_9813);
or UO_526 (O_526,N_9790,N_9816);
xor UO_527 (O_527,N_9800,N_9540);
xnor UO_528 (O_528,N_9783,N_9690);
and UO_529 (O_529,N_9648,N_9891);
and UO_530 (O_530,N_9658,N_9979);
xnor UO_531 (O_531,N_9980,N_9927);
nand UO_532 (O_532,N_9529,N_9580);
nand UO_533 (O_533,N_9861,N_9620);
nand UO_534 (O_534,N_9710,N_9695);
xnor UO_535 (O_535,N_9620,N_9604);
or UO_536 (O_536,N_9732,N_9745);
or UO_537 (O_537,N_9992,N_9703);
or UO_538 (O_538,N_9776,N_9710);
and UO_539 (O_539,N_9571,N_9745);
nor UO_540 (O_540,N_9644,N_9559);
nor UO_541 (O_541,N_9814,N_9818);
nor UO_542 (O_542,N_9966,N_9579);
nor UO_543 (O_543,N_9613,N_9587);
or UO_544 (O_544,N_9823,N_9598);
xor UO_545 (O_545,N_9765,N_9843);
nor UO_546 (O_546,N_9883,N_9756);
or UO_547 (O_547,N_9742,N_9789);
xor UO_548 (O_548,N_9907,N_9877);
or UO_549 (O_549,N_9819,N_9922);
xnor UO_550 (O_550,N_9799,N_9934);
nor UO_551 (O_551,N_9841,N_9745);
and UO_552 (O_552,N_9735,N_9524);
nand UO_553 (O_553,N_9778,N_9662);
nand UO_554 (O_554,N_9890,N_9799);
nor UO_555 (O_555,N_9587,N_9620);
nor UO_556 (O_556,N_9646,N_9755);
or UO_557 (O_557,N_9960,N_9958);
nand UO_558 (O_558,N_9644,N_9948);
or UO_559 (O_559,N_9748,N_9577);
xor UO_560 (O_560,N_9661,N_9771);
nand UO_561 (O_561,N_9863,N_9771);
nor UO_562 (O_562,N_9856,N_9954);
nand UO_563 (O_563,N_9974,N_9965);
and UO_564 (O_564,N_9721,N_9782);
nor UO_565 (O_565,N_9802,N_9686);
or UO_566 (O_566,N_9534,N_9829);
nor UO_567 (O_567,N_9564,N_9691);
xnor UO_568 (O_568,N_9961,N_9773);
nand UO_569 (O_569,N_9785,N_9920);
xor UO_570 (O_570,N_9752,N_9910);
nand UO_571 (O_571,N_9765,N_9745);
and UO_572 (O_572,N_9828,N_9632);
nand UO_573 (O_573,N_9787,N_9606);
xor UO_574 (O_574,N_9973,N_9852);
nor UO_575 (O_575,N_9576,N_9662);
nor UO_576 (O_576,N_9885,N_9947);
nor UO_577 (O_577,N_9982,N_9955);
and UO_578 (O_578,N_9766,N_9592);
or UO_579 (O_579,N_9825,N_9877);
or UO_580 (O_580,N_9998,N_9858);
nor UO_581 (O_581,N_9566,N_9954);
nor UO_582 (O_582,N_9705,N_9562);
nor UO_583 (O_583,N_9984,N_9634);
or UO_584 (O_584,N_9848,N_9937);
xor UO_585 (O_585,N_9918,N_9743);
xnor UO_586 (O_586,N_9832,N_9772);
nand UO_587 (O_587,N_9916,N_9986);
and UO_588 (O_588,N_9745,N_9932);
and UO_589 (O_589,N_9557,N_9588);
nor UO_590 (O_590,N_9742,N_9676);
nor UO_591 (O_591,N_9735,N_9503);
nor UO_592 (O_592,N_9965,N_9504);
xnor UO_593 (O_593,N_9819,N_9636);
xor UO_594 (O_594,N_9915,N_9857);
xor UO_595 (O_595,N_9519,N_9541);
nand UO_596 (O_596,N_9971,N_9846);
xor UO_597 (O_597,N_9570,N_9750);
nand UO_598 (O_598,N_9579,N_9958);
nor UO_599 (O_599,N_9811,N_9622);
and UO_600 (O_600,N_9952,N_9722);
nor UO_601 (O_601,N_9947,N_9637);
xnor UO_602 (O_602,N_9882,N_9912);
nand UO_603 (O_603,N_9756,N_9586);
nand UO_604 (O_604,N_9759,N_9890);
and UO_605 (O_605,N_9755,N_9763);
and UO_606 (O_606,N_9917,N_9732);
xnor UO_607 (O_607,N_9786,N_9603);
xor UO_608 (O_608,N_9832,N_9737);
xor UO_609 (O_609,N_9968,N_9731);
nor UO_610 (O_610,N_9905,N_9952);
nand UO_611 (O_611,N_9521,N_9787);
xor UO_612 (O_612,N_9751,N_9672);
and UO_613 (O_613,N_9841,N_9756);
or UO_614 (O_614,N_9719,N_9544);
nand UO_615 (O_615,N_9963,N_9990);
and UO_616 (O_616,N_9580,N_9973);
nor UO_617 (O_617,N_9785,N_9702);
or UO_618 (O_618,N_9549,N_9724);
xor UO_619 (O_619,N_9790,N_9743);
nand UO_620 (O_620,N_9832,N_9970);
xnor UO_621 (O_621,N_9524,N_9786);
xnor UO_622 (O_622,N_9643,N_9880);
nand UO_623 (O_623,N_9923,N_9664);
nand UO_624 (O_624,N_9617,N_9973);
nor UO_625 (O_625,N_9557,N_9733);
nor UO_626 (O_626,N_9770,N_9769);
nand UO_627 (O_627,N_9907,N_9987);
and UO_628 (O_628,N_9994,N_9903);
xor UO_629 (O_629,N_9953,N_9695);
and UO_630 (O_630,N_9680,N_9782);
and UO_631 (O_631,N_9879,N_9715);
and UO_632 (O_632,N_9994,N_9789);
or UO_633 (O_633,N_9712,N_9899);
xor UO_634 (O_634,N_9532,N_9841);
or UO_635 (O_635,N_9547,N_9897);
or UO_636 (O_636,N_9751,N_9619);
and UO_637 (O_637,N_9666,N_9551);
or UO_638 (O_638,N_9802,N_9982);
nand UO_639 (O_639,N_9934,N_9979);
and UO_640 (O_640,N_9729,N_9897);
or UO_641 (O_641,N_9942,N_9517);
nand UO_642 (O_642,N_9830,N_9563);
xor UO_643 (O_643,N_9590,N_9781);
xor UO_644 (O_644,N_9819,N_9877);
xor UO_645 (O_645,N_9565,N_9618);
and UO_646 (O_646,N_9967,N_9583);
nand UO_647 (O_647,N_9888,N_9730);
and UO_648 (O_648,N_9808,N_9929);
and UO_649 (O_649,N_9690,N_9577);
and UO_650 (O_650,N_9977,N_9569);
nor UO_651 (O_651,N_9888,N_9976);
nor UO_652 (O_652,N_9895,N_9957);
or UO_653 (O_653,N_9718,N_9784);
and UO_654 (O_654,N_9580,N_9832);
or UO_655 (O_655,N_9792,N_9786);
nor UO_656 (O_656,N_9995,N_9894);
or UO_657 (O_657,N_9600,N_9987);
nand UO_658 (O_658,N_9538,N_9964);
or UO_659 (O_659,N_9807,N_9601);
nor UO_660 (O_660,N_9716,N_9514);
and UO_661 (O_661,N_9820,N_9514);
nor UO_662 (O_662,N_9608,N_9580);
nand UO_663 (O_663,N_9846,N_9994);
and UO_664 (O_664,N_9531,N_9794);
nor UO_665 (O_665,N_9897,N_9502);
xnor UO_666 (O_666,N_9866,N_9505);
or UO_667 (O_667,N_9781,N_9653);
and UO_668 (O_668,N_9664,N_9797);
nand UO_669 (O_669,N_9666,N_9516);
nand UO_670 (O_670,N_9618,N_9760);
or UO_671 (O_671,N_9924,N_9844);
nand UO_672 (O_672,N_9992,N_9637);
nand UO_673 (O_673,N_9733,N_9674);
and UO_674 (O_674,N_9506,N_9858);
and UO_675 (O_675,N_9566,N_9744);
and UO_676 (O_676,N_9886,N_9557);
and UO_677 (O_677,N_9696,N_9643);
nand UO_678 (O_678,N_9935,N_9867);
nand UO_679 (O_679,N_9539,N_9614);
nor UO_680 (O_680,N_9686,N_9827);
and UO_681 (O_681,N_9992,N_9513);
and UO_682 (O_682,N_9548,N_9656);
and UO_683 (O_683,N_9750,N_9597);
xnor UO_684 (O_684,N_9956,N_9585);
or UO_685 (O_685,N_9509,N_9668);
nor UO_686 (O_686,N_9684,N_9515);
xnor UO_687 (O_687,N_9527,N_9811);
xnor UO_688 (O_688,N_9812,N_9617);
nand UO_689 (O_689,N_9601,N_9655);
nor UO_690 (O_690,N_9903,N_9553);
xnor UO_691 (O_691,N_9939,N_9678);
and UO_692 (O_692,N_9697,N_9508);
nor UO_693 (O_693,N_9656,N_9661);
and UO_694 (O_694,N_9713,N_9690);
xor UO_695 (O_695,N_9653,N_9844);
and UO_696 (O_696,N_9584,N_9796);
nand UO_697 (O_697,N_9554,N_9623);
nor UO_698 (O_698,N_9575,N_9546);
nand UO_699 (O_699,N_9856,N_9804);
nor UO_700 (O_700,N_9841,N_9820);
and UO_701 (O_701,N_9901,N_9794);
xor UO_702 (O_702,N_9760,N_9951);
nand UO_703 (O_703,N_9650,N_9676);
or UO_704 (O_704,N_9745,N_9619);
xnor UO_705 (O_705,N_9729,N_9904);
and UO_706 (O_706,N_9849,N_9994);
or UO_707 (O_707,N_9679,N_9921);
xnor UO_708 (O_708,N_9791,N_9686);
and UO_709 (O_709,N_9520,N_9963);
nor UO_710 (O_710,N_9726,N_9592);
nor UO_711 (O_711,N_9746,N_9664);
xnor UO_712 (O_712,N_9667,N_9843);
nor UO_713 (O_713,N_9911,N_9653);
and UO_714 (O_714,N_9858,N_9793);
nor UO_715 (O_715,N_9805,N_9797);
or UO_716 (O_716,N_9888,N_9659);
and UO_717 (O_717,N_9934,N_9647);
xnor UO_718 (O_718,N_9736,N_9735);
nand UO_719 (O_719,N_9903,N_9595);
and UO_720 (O_720,N_9524,N_9756);
xnor UO_721 (O_721,N_9575,N_9513);
or UO_722 (O_722,N_9659,N_9787);
xor UO_723 (O_723,N_9672,N_9757);
or UO_724 (O_724,N_9829,N_9774);
nor UO_725 (O_725,N_9678,N_9894);
or UO_726 (O_726,N_9958,N_9948);
xor UO_727 (O_727,N_9851,N_9616);
xor UO_728 (O_728,N_9670,N_9551);
and UO_729 (O_729,N_9891,N_9701);
nand UO_730 (O_730,N_9570,N_9783);
and UO_731 (O_731,N_9954,N_9670);
nand UO_732 (O_732,N_9741,N_9516);
nand UO_733 (O_733,N_9766,N_9697);
or UO_734 (O_734,N_9590,N_9961);
nor UO_735 (O_735,N_9795,N_9707);
or UO_736 (O_736,N_9507,N_9978);
nor UO_737 (O_737,N_9744,N_9954);
nor UO_738 (O_738,N_9637,N_9931);
or UO_739 (O_739,N_9635,N_9542);
nand UO_740 (O_740,N_9554,N_9992);
nand UO_741 (O_741,N_9776,N_9870);
nor UO_742 (O_742,N_9978,N_9848);
and UO_743 (O_743,N_9849,N_9674);
and UO_744 (O_744,N_9627,N_9661);
nand UO_745 (O_745,N_9529,N_9886);
and UO_746 (O_746,N_9975,N_9875);
or UO_747 (O_747,N_9510,N_9691);
or UO_748 (O_748,N_9795,N_9969);
xor UO_749 (O_749,N_9833,N_9689);
nor UO_750 (O_750,N_9983,N_9957);
or UO_751 (O_751,N_9636,N_9797);
nor UO_752 (O_752,N_9622,N_9543);
and UO_753 (O_753,N_9803,N_9911);
and UO_754 (O_754,N_9839,N_9649);
nand UO_755 (O_755,N_9516,N_9805);
xnor UO_756 (O_756,N_9605,N_9523);
nor UO_757 (O_757,N_9520,N_9911);
and UO_758 (O_758,N_9890,N_9941);
and UO_759 (O_759,N_9930,N_9632);
and UO_760 (O_760,N_9822,N_9782);
and UO_761 (O_761,N_9986,N_9931);
nor UO_762 (O_762,N_9785,N_9787);
xnor UO_763 (O_763,N_9632,N_9830);
and UO_764 (O_764,N_9973,N_9592);
nor UO_765 (O_765,N_9963,N_9993);
nand UO_766 (O_766,N_9968,N_9915);
nor UO_767 (O_767,N_9561,N_9541);
xor UO_768 (O_768,N_9959,N_9819);
nor UO_769 (O_769,N_9610,N_9759);
xnor UO_770 (O_770,N_9793,N_9625);
xor UO_771 (O_771,N_9572,N_9696);
and UO_772 (O_772,N_9789,N_9738);
nor UO_773 (O_773,N_9718,N_9779);
nor UO_774 (O_774,N_9774,N_9596);
xor UO_775 (O_775,N_9520,N_9945);
xnor UO_776 (O_776,N_9830,N_9526);
or UO_777 (O_777,N_9974,N_9860);
nand UO_778 (O_778,N_9992,N_9958);
and UO_779 (O_779,N_9826,N_9657);
nand UO_780 (O_780,N_9564,N_9998);
nand UO_781 (O_781,N_9982,N_9617);
nand UO_782 (O_782,N_9747,N_9800);
nand UO_783 (O_783,N_9784,N_9616);
and UO_784 (O_784,N_9654,N_9986);
or UO_785 (O_785,N_9562,N_9964);
or UO_786 (O_786,N_9906,N_9540);
and UO_787 (O_787,N_9639,N_9726);
nand UO_788 (O_788,N_9681,N_9762);
nand UO_789 (O_789,N_9671,N_9969);
nand UO_790 (O_790,N_9648,N_9542);
xor UO_791 (O_791,N_9653,N_9650);
nor UO_792 (O_792,N_9673,N_9794);
or UO_793 (O_793,N_9681,N_9904);
nor UO_794 (O_794,N_9836,N_9703);
nor UO_795 (O_795,N_9557,N_9952);
nand UO_796 (O_796,N_9613,N_9873);
xor UO_797 (O_797,N_9935,N_9988);
nand UO_798 (O_798,N_9678,N_9743);
or UO_799 (O_799,N_9519,N_9827);
xnor UO_800 (O_800,N_9908,N_9953);
or UO_801 (O_801,N_9831,N_9583);
or UO_802 (O_802,N_9583,N_9848);
nor UO_803 (O_803,N_9789,N_9953);
xor UO_804 (O_804,N_9729,N_9609);
xor UO_805 (O_805,N_9906,N_9986);
nor UO_806 (O_806,N_9542,N_9748);
and UO_807 (O_807,N_9979,N_9721);
and UO_808 (O_808,N_9869,N_9687);
nor UO_809 (O_809,N_9680,N_9556);
xor UO_810 (O_810,N_9754,N_9858);
nor UO_811 (O_811,N_9504,N_9757);
xor UO_812 (O_812,N_9673,N_9679);
and UO_813 (O_813,N_9855,N_9611);
and UO_814 (O_814,N_9766,N_9787);
nor UO_815 (O_815,N_9520,N_9509);
or UO_816 (O_816,N_9591,N_9911);
and UO_817 (O_817,N_9929,N_9971);
nand UO_818 (O_818,N_9608,N_9504);
and UO_819 (O_819,N_9743,N_9999);
xnor UO_820 (O_820,N_9926,N_9537);
nand UO_821 (O_821,N_9843,N_9618);
and UO_822 (O_822,N_9798,N_9943);
xnor UO_823 (O_823,N_9542,N_9909);
or UO_824 (O_824,N_9879,N_9781);
and UO_825 (O_825,N_9925,N_9749);
nand UO_826 (O_826,N_9933,N_9666);
and UO_827 (O_827,N_9689,N_9558);
and UO_828 (O_828,N_9631,N_9745);
nand UO_829 (O_829,N_9939,N_9667);
and UO_830 (O_830,N_9808,N_9732);
nor UO_831 (O_831,N_9591,N_9758);
and UO_832 (O_832,N_9656,N_9887);
nor UO_833 (O_833,N_9907,N_9528);
or UO_834 (O_834,N_9500,N_9841);
nand UO_835 (O_835,N_9686,N_9800);
and UO_836 (O_836,N_9618,N_9714);
xor UO_837 (O_837,N_9777,N_9927);
nand UO_838 (O_838,N_9846,N_9646);
and UO_839 (O_839,N_9639,N_9637);
nand UO_840 (O_840,N_9737,N_9521);
nor UO_841 (O_841,N_9709,N_9826);
nor UO_842 (O_842,N_9655,N_9779);
and UO_843 (O_843,N_9615,N_9720);
or UO_844 (O_844,N_9516,N_9952);
xor UO_845 (O_845,N_9630,N_9561);
nand UO_846 (O_846,N_9557,N_9804);
or UO_847 (O_847,N_9502,N_9602);
xor UO_848 (O_848,N_9959,N_9702);
nand UO_849 (O_849,N_9811,N_9855);
xor UO_850 (O_850,N_9717,N_9700);
xnor UO_851 (O_851,N_9927,N_9550);
xor UO_852 (O_852,N_9581,N_9819);
xnor UO_853 (O_853,N_9743,N_9534);
and UO_854 (O_854,N_9802,N_9803);
and UO_855 (O_855,N_9603,N_9601);
nor UO_856 (O_856,N_9746,N_9759);
nor UO_857 (O_857,N_9789,N_9976);
or UO_858 (O_858,N_9849,N_9773);
nand UO_859 (O_859,N_9682,N_9865);
or UO_860 (O_860,N_9631,N_9663);
nand UO_861 (O_861,N_9904,N_9602);
and UO_862 (O_862,N_9773,N_9783);
xnor UO_863 (O_863,N_9938,N_9571);
nand UO_864 (O_864,N_9660,N_9930);
nor UO_865 (O_865,N_9507,N_9644);
xnor UO_866 (O_866,N_9892,N_9570);
or UO_867 (O_867,N_9636,N_9852);
nand UO_868 (O_868,N_9926,N_9536);
xnor UO_869 (O_869,N_9926,N_9696);
and UO_870 (O_870,N_9841,N_9775);
or UO_871 (O_871,N_9807,N_9858);
nor UO_872 (O_872,N_9976,N_9644);
xor UO_873 (O_873,N_9903,N_9573);
xnor UO_874 (O_874,N_9538,N_9847);
and UO_875 (O_875,N_9590,N_9626);
nor UO_876 (O_876,N_9741,N_9687);
xnor UO_877 (O_877,N_9697,N_9593);
or UO_878 (O_878,N_9824,N_9737);
and UO_879 (O_879,N_9811,N_9544);
xor UO_880 (O_880,N_9726,N_9640);
nand UO_881 (O_881,N_9890,N_9752);
or UO_882 (O_882,N_9620,N_9813);
or UO_883 (O_883,N_9884,N_9961);
or UO_884 (O_884,N_9508,N_9774);
nand UO_885 (O_885,N_9882,N_9928);
and UO_886 (O_886,N_9801,N_9524);
nor UO_887 (O_887,N_9758,N_9675);
nand UO_888 (O_888,N_9734,N_9686);
nand UO_889 (O_889,N_9694,N_9701);
xor UO_890 (O_890,N_9615,N_9806);
xor UO_891 (O_891,N_9631,N_9881);
and UO_892 (O_892,N_9866,N_9665);
nor UO_893 (O_893,N_9591,N_9763);
xnor UO_894 (O_894,N_9734,N_9701);
nand UO_895 (O_895,N_9843,N_9603);
nor UO_896 (O_896,N_9583,N_9766);
or UO_897 (O_897,N_9818,N_9881);
nor UO_898 (O_898,N_9584,N_9845);
or UO_899 (O_899,N_9753,N_9695);
or UO_900 (O_900,N_9861,N_9610);
nor UO_901 (O_901,N_9916,N_9838);
or UO_902 (O_902,N_9950,N_9702);
and UO_903 (O_903,N_9865,N_9545);
xor UO_904 (O_904,N_9993,N_9737);
xor UO_905 (O_905,N_9583,N_9896);
and UO_906 (O_906,N_9595,N_9614);
and UO_907 (O_907,N_9825,N_9797);
xor UO_908 (O_908,N_9790,N_9973);
nand UO_909 (O_909,N_9900,N_9516);
nor UO_910 (O_910,N_9505,N_9670);
nand UO_911 (O_911,N_9724,N_9890);
nor UO_912 (O_912,N_9824,N_9969);
xnor UO_913 (O_913,N_9958,N_9565);
nand UO_914 (O_914,N_9568,N_9794);
nand UO_915 (O_915,N_9788,N_9786);
or UO_916 (O_916,N_9985,N_9888);
nand UO_917 (O_917,N_9918,N_9638);
xnor UO_918 (O_918,N_9705,N_9703);
and UO_919 (O_919,N_9903,N_9803);
xnor UO_920 (O_920,N_9649,N_9989);
nand UO_921 (O_921,N_9877,N_9883);
or UO_922 (O_922,N_9650,N_9540);
nand UO_923 (O_923,N_9849,N_9841);
nand UO_924 (O_924,N_9938,N_9939);
nor UO_925 (O_925,N_9937,N_9620);
nor UO_926 (O_926,N_9652,N_9953);
and UO_927 (O_927,N_9571,N_9993);
xnor UO_928 (O_928,N_9815,N_9555);
nor UO_929 (O_929,N_9562,N_9578);
and UO_930 (O_930,N_9623,N_9855);
nand UO_931 (O_931,N_9766,N_9710);
or UO_932 (O_932,N_9533,N_9688);
nand UO_933 (O_933,N_9989,N_9870);
nor UO_934 (O_934,N_9532,N_9588);
and UO_935 (O_935,N_9638,N_9727);
nand UO_936 (O_936,N_9751,N_9533);
nor UO_937 (O_937,N_9532,N_9775);
or UO_938 (O_938,N_9817,N_9665);
or UO_939 (O_939,N_9564,N_9661);
nor UO_940 (O_940,N_9877,N_9984);
nor UO_941 (O_941,N_9821,N_9838);
and UO_942 (O_942,N_9571,N_9758);
xnor UO_943 (O_943,N_9922,N_9875);
xor UO_944 (O_944,N_9801,N_9884);
xor UO_945 (O_945,N_9685,N_9846);
and UO_946 (O_946,N_9819,N_9674);
nand UO_947 (O_947,N_9797,N_9776);
or UO_948 (O_948,N_9952,N_9970);
xnor UO_949 (O_949,N_9656,N_9833);
nor UO_950 (O_950,N_9560,N_9775);
and UO_951 (O_951,N_9568,N_9583);
and UO_952 (O_952,N_9818,N_9543);
xor UO_953 (O_953,N_9747,N_9750);
and UO_954 (O_954,N_9569,N_9720);
and UO_955 (O_955,N_9620,N_9680);
or UO_956 (O_956,N_9852,N_9601);
or UO_957 (O_957,N_9614,N_9958);
and UO_958 (O_958,N_9644,N_9799);
and UO_959 (O_959,N_9725,N_9822);
or UO_960 (O_960,N_9552,N_9544);
xor UO_961 (O_961,N_9598,N_9613);
and UO_962 (O_962,N_9526,N_9844);
xnor UO_963 (O_963,N_9564,N_9692);
xor UO_964 (O_964,N_9936,N_9882);
nand UO_965 (O_965,N_9652,N_9925);
nand UO_966 (O_966,N_9949,N_9882);
xor UO_967 (O_967,N_9894,N_9741);
xnor UO_968 (O_968,N_9946,N_9534);
nor UO_969 (O_969,N_9738,N_9718);
and UO_970 (O_970,N_9880,N_9509);
and UO_971 (O_971,N_9915,N_9726);
or UO_972 (O_972,N_9941,N_9959);
or UO_973 (O_973,N_9878,N_9762);
nor UO_974 (O_974,N_9725,N_9735);
nor UO_975 (O_975,N_9590,N_9894);
nand UO_976 (O_976,N_9941,N_9696);
nor UO_977 (O_977,N_9786,N_9558);
or UO_978 (O_978,N_9714,N_9799);
or UO_979 (O_979,N_9690,N_9529);
and UO_980 (O_980,N_9801,N_9874);
xnor UO_981 (O_981,N_9889,N_9994);
nand UO_982 (O_982,N_9618,N_9739);
nand UO_983 (O_983,N_9891,N_9549);
nand UO_984 (O_984,N_9622,N_9918);
nand UO_985 (O_985,N_9820,N_9569);
nand UO_986 (O_986,N_9594,N_9654);
xnor UO_987 (O_987,N_9586,N_9648);
nand UO_988 (O_988,N_9980,N_9790);
nand UO_989 (O_989,N_9922,N_9609);
nand UO_990 (O_990,N_9944,N_9687);
xor UO_991 (O_991,N_9508,N_9862);
nor UO_992 (O_992,N_9645,N_9658);
nand UO_993 (O_993,N_9560,N_9801);
nand UO_994 (O_994,N_9813,N_9882);
and UO_995 (O_995,N_9931,N_9849);
nor UO_996 (O_996,N_9560,N_9652);
and UO_997 (O_997,N_9846,N_9963);
xnor UO_998 (O_998,N_9713,N_9717);
or UO_999 (O_999,N_9755,N_9764);
and UO_1000 (O_1000,N_9510,N_9978);
or UO_1001 (O_1001,N_9892,N_9654);
or UO_1002 (O_1002,N_9630,N_9974);
and UO_1003 (O_1003,N_9750,N_9961);
nand UO_1004 (O_1004,N_9850,N_9753);
xor UO_1005 (O_1005,N_9823,N_9542);
or UO_1006 (O_1006,N_9709,N_9706);
xnor UO_1007 (O_1007,N_9912,N_9812);
nor UO_1008 (O_1008,N_9776,N_9562);
nand UO_1009 (O_1009,N_9865,N_9962);
nand UO_1010 (O_1010,N_9796,N_9592);
nand UO_1011 (O_1011,N_9806,N_9734);
xor UO_1012 (O_1012,N_9929,N_9518);
and UO_1013 (O_1013,N_9881,N_9536);
xor UO_1014 (O_1014,N_9641,N_9565);
or UO_1015 (O_1015,N_9686,N_9585);
or UO_1016 (O_1016,N_9704,N_9652);
and UO_1017 (O_1017,N_9567,N_9635);
and UO_1018 (O_1018,N_9972,N_9613);
nor UO_1019 (O_1019,N_9805,N_9874);
nand UO_1020 (O_1020,N_9650,N_9805);
xor UO_1021 (O_1021,N_9716,N_9840);
and UO_1022 (O_1022,N_9626,N_9698);
nand UO_1023 (O_1023,N_9627,N_9897);
xor UO_1024 (O_1024,N_9537,N_9572);
nor UO_1025 (O_1025,N_9599,N_9950);
nor UO_1026 (O_1026,N_9654,N_9911);
nor UO_1027 (O_1027,N_9710,N_9664);
nor UO_1028 (O_1028,N_9728,N_9769);
and UO_1029 (O_1029,N_9827,N_9516);
and UO_1030 (O_1030,N_9833,N_9581);
xor UO_1031 (O_1031,N_9655,N_9705);
or UO_1032 (O_1032,N_9826,N_9964);
or UO_1033 (O_1033,N_9854,N_9621);
xnor UO_1034 (O_1034,N_9868,N_9618);
and UO_1035 (O_1035,N_9630,N_9722);
and UO_1036 (O_1036,N_9577,N_9806);
and UO_1037 (O_1037,N_9774,N_9678);
nor UO_1038 (O_1038,N_9975,N_9615);
xor UO_1039 (O_1039,N_9686,N_9933);
xor UO_1040 (O_1040,N_9789,N_9621);
nor UO_1041 (O_1041,N_9886,N_9829);
nor UO_1042 (O_1042,N_9716,N_9948);
nor UO_1043 (O_1043,N_9776,N_9729);
nor UO_1044 (O_1044,N_9702,N_9969);
nand UO_1045 (O_1045,N_9514,N_9525);
nor UO_1046 (O_1046,N_9697,N_9709);
or UO_1047 (O_1047,N_9819,N_9556);
xor UO_1048 (O_1048,N_9527,N_9837);
or UO_1049 (O_1049,N_9880,N_9538);
xnor UO_1050 (O_1050,N_9667,N_9818);
nor UO_1051 (O_1051,N_9939,N_9956);
and UO_1052 (O_1052,N_9699,N_9598);
and UO_1053 (O_1053,N_9654,N_9909);
nor UO_1054 (O_1054,N_9854,N_9506);
nor UO_1055 (O_1055,N_9798,N_9808);
and UO_1056 (O_1056,N_9681,N_9610);
xnor UO_1057 (O_1057,N_9807,N_9639);
nand UO_1058 (O_1058,N_9928,N_9718);
nand UO_1059 (O_1059,N_9908,N_9910);
or UO_1060 (O_1060,N_9873,N_9994);
nand UO_1061 (O_1061,N_9888,N_9722);
and UO_1062 (O_1062,N_9902,N_9559);
xnor UO_1063 (O_1063,N_9886,N_9792);
nand UO_1064 (O_1064,N_9506,N_9608);
xor UO_1065 (O_1065,N_9731,N_9641);
nor UO_1066 (O_1066,N_9522,N_9628);
or UO_1067 (O_1067,N_9772,N_9549);
and UO_1068 (O_1068,N_9627,N_9570);
or UO_1069 (O_1069,N_9576,N_9718);
nand UO_1070 (O_1070,N_9551,N_9671);
nor UO_1071 (O_1071,N_9787,N_9865);
nand UO_1072 (O_1072,N_9735,N_9836);
xnor UO_1073 (O_1073,N_9646,N_9588);
and UO_1074 (O_1074,N_9805,N_9780);
and UO_1075 (O_1075,N_9614,N_9766);
nor UO_1076 (O_1076,N_9774,N_9870);
or UO_1077 (O_1077,N_9607,N_9794);
nand UO_1078 (O_1078,N_9561,N_9778);
nand UO_1079 (O_1079,N_9792,N_9997);
or UO_1080 (O_1080,N_9581,N_9584);
nand UO_1081 (O_1081,N_9973,N_9624);
nand UO_1082 (O_1082,N_9807,N_9824);
or UO_1083 (O_1083,N_9917,N_9701);
xnor UO_1084 (O_1084,N_9538,N_9736);
xnor UO_1085 (O_1085,N_9680,N_9788);
and UO_1086 (O_1086,N_9813,N_9987);
nand UO_1087 (O_1087,N_9809,N_9640);
nand UO_1088 (O_1088,N_9788,N_9961);
xor UO_1089 (O_1089,N_9724,N_9632);
nand UO_1090 (O_1090,N_9501,N_9593);
or UO_1091 (O_1091,N_9571,N_9588);
and UO_1092 (O_1092,N_9587,N_9934);
and UO_1093 (O_1093,N_9518,N_9859);
xor UO_1094 (O_1094,N_9739,N_9625);
xor UO_1095 (O_1095,N_9789,N_9848);
xnor UO_1096 (O_1096,N_9929,N_9908);
and UO_1097 (O_1097,N_9779,N_9918);
or UO_1098 (O_1098,N_9547,N_9860);
and UO_1099 (O_1099,N_9504,N_9801);
nand UO_1100 (O_1100,N_9732,N_9985);
nor UO_1101 (O_1101,N_9509,N_9872);
nor UO_1102 (O_1102,N_9793,N_9654);
nand UO_1103 (O_1103,N_9950,N_9930);
nand UO_1104 (O_1104,N_9578,N_9824);
nor UO_1105 (O_1105,N_9930,N_9589);
or UO_1106 (O_1106,N_9681,N_9716);
or UO_1107 (O_1107,N_9811,N_9556);
nor UO_1108 (O_1108,N_9680,N_9965);
xnor UO_1109 (O_1109,N_9923,N_9926);
nor UO_1110 (O_1110,N_9985,N_9560);
nor UO_1111 (O_1111,N_9698,N_9686);
nand UO_1112 (O_1112,N_9710,N_9741);
nor UO_1113 (O_1113,N_9905,N_9599);
or UO_1114 (O_1114,N_9851,N_9570);
and UO_1115 (O_1115,N_9674,N_9904);
and UO_1116 (O_1116,N_9886,N_9690);
nand UO_1117 (O_1117,N_9533,N_9898);
nor UO_1118 (O_1118,N_9565,N_9545);
xor UO_1119 (O_1119,N_9853,N_9803);
nand UO_1120 (O_1120,N_9853,N_9544);
or UO_1121 (O_1121,N_9726,N_9664);
xor UO_1122 (O_1122,N_9862,N_9619);
and UO_1123 (O_1123,N_9808,N_9874);
and UO_1124 (O_1124,N_9902,N_9573);
nand UO_1125 (O_1125,N_9782,N_9619);
nor UO_1126 (O_1126,N_9586,N_9775);
nand UO_1127 (O_1127,N_9580,N_9579);
and UO_1128 (O_1128,N_9677,N_9892);
and UO_1129 (O_1129,N_9705,N_9722);
and UO_1130 (O_1130,N_9950,N_9830);
nor UO_1131 (O_1131,N_9815,N_9874);
or UO_1132 (O_1132,N_9996,N_9702);
and UO_1133 (O_1133,N_9687,N_9636);
or UO_1134 (O_1134,N_9665,N_9814);
or UO_1135 (O_1135,N_9540,N_9719);
or UO_1136 (O_1136,N_9962,N_9626);
and UO_1137 (O_1137,N_9540,N_9601);
xor UO_1138 (O_1138,N_9694,N_9793);
nand UO_1139 (O_1139,N_9834,N_9930);
nand UO_1140 (O_1140,N_9533,N_9506);
nor UO_1141 (O_1141,N_9769,N_9923);
xnor UO_1142 (O_1142,N_9761,N_9838);
and UO_1143 (O_1143,N_9509,N_9782);
nor UO_1144 (O_1144,N_9544,N_9753);
nand UO_1145 (O_1145,N_9530,N_9773);
nand UO_1146 (O_1146,N_9691,N_9575);
nand UO_1147 (O_1147,N_9700,N_9964);
xnor UO_1148 (O_1148,N_9754,N_9804);
or UO_1149 (O_1149,N_9799,N_9806);
and UO_1150 (O_1150,N_9705,N_9601);
nand UO_1151 (O_1151,N_9778,N_9959);
or UO_1152 (O_1152,N_9536,N_9906);
and UO_1153 (O_1153,N_9723,N_9531);
and UO_1154 (O_1154,N_9675,N_9710);
nand UO_1155 (O_1155,N_9620,N_9686);
and UO_1156 (O_1156,N_9853,N_9859);
xor UO_1157 (O_1157,N_9775,N_9838);
or UO_1158 (O_1158,N_9955,N_9937);
or UO_1159 (O_1159,N_9914,N_9666);
and UO_1160 (O_1160,N_9583,N_9887);
and UO_1161 (O_1161,N_9716,N_9877);
xor UO_1162 (O_1162,N_9951,N_9800);
xor UO_1163 (O_1163,N_9516,N_9531);
or UO_1164 (O_1164,N_9843,N_9581);
xor UO_1165 (O_1165,N_9642,N_9988);
and UO_1166 (O_1166,N_9633,N_9612);
xnor UO_1167 (O_1167,N_9557,N_9676);
nand UO_1168 (O_1168,N_9959,N_9923);
and UO_1169 (O_1169,N_9892,N_9672);
and UO_1170 (O_1170,N_9916,N_9867);
and UO_1171 (O_1171,N_9850,N_9724);
xnor UO_1172 (O_1172,N_9873,N_9567);
xnor UO_1173 (O_1173,N_9558,N_9580);
and UO_1174 (O_1174,N_9607,N_9534);
or UO_1175 (O_1175,N_9962,N_9642);
nand UO_1176 (O_1176,N_9514,N_9647);
nand UO_1177 (O_1177,N_9607,N_9781);
xnor UO_1178 (O_1178,N_9732,N_9837);
and UO_1179 (O_1179,N_9925,N_9897);
and UO_1180 (O_1180,N_9522,N_9523);
or UO_1181 (O_1181,N_9803,N_9705);
nor UO_1182 (O_1182,N_9904,N_9782);
and UO_1183 (O_1183,N_9868,N_9968);
and UO_1184 (O_1184,N_9820,N_9597);
and UO_1185 (O_1185,N_9982,N_9533);
xor UO_1186 (O_1186,N_9509,N_9832);
nand UO_1187 (O_1187,N_9783,N_9920);
nor UO_1188 (O_1188,N_9542,N_9683);
or UO_1189 (O_1189,N_9746,N_9595);
xnor UO_1190 (O_1190,N_9517,N_9694);
xor UO_1191 (O_1191,N_9538,N_9778);
and UO_1192 (O_1192,N_9559,N_9617);
or UO_1193 (O_1193,N_9591,N_9737);
and UO_1194 (O_1194,N_9878,N_9502);
and UO_1195 (O_1195,N_9758,N_9772);
xor UO_1196 (O_1196,N_9982,N_9653);
or UO_1197 (O_1197,N_9847,N_9500);
xor UO_1198 (O_1198,N_9657,N_9891);
nor UO_1199 (O_1199,N_9618,N_9545);
xnor UO_1200 (O_1200,N_9885,N_9517);
or UO_1201 (O_1201,N_9764,N_9503);
xor UO_1202 (O_1202,N_9562,N_9876);
nor UO_1203 (O_1203,N_9955,N_9604);
nand UO_1204 (O_1204,N_9690,N_9930);
nand UO_1205 (O_1205,N_9720,N_9754);
nand UO_1206 (O_1206,N_9884,N_9538);
or UO_1207 (O_1207,N_9761,N_9759);
and UO_1208 (O_1208,N_9604,N_9533);
xnor UO_1209 (O_1209,N_9874,N_9661);
and UO_1210 (O_1210,N_9945,N_9591);
nor UO_1211 (O_1211,N_9654,N_9596);
xnor UO_1212 (O_1212,N_9992,N_9983);
nor UO_1213 (O_1213,N_9730,N_9970);
and UO_1214 (O_1214,N_9968,N_9775);
xnor UO_1215 (O_1215,N_9528,N_9782);
or UO_1216 (O_1216,N_9680,N_9876);
xnor UO_1217 (O_1217,N_9954,N_9964);
xor UO_1218 (O_1218,N_9814,N_9601);
xnor UO_1219 (O_1219,N_9741,N_9594);
nand UO_1220 (O_1220,N_9505,N_9713);
nand UO_1221 (O_1221,N_9767,N_9879);
or UO_1222 (O_1222,N_9832,N_9922);
or UO_1223 (O_1223,N_9592,N_9841);
nor UO_1224 (O_1224,N_9834,N_9845);
nand UO_1225 (O_1225,N_9657,N_9762);
nor UO_1226 (O_1226,N_9965,N_9701);
and UO_1227 (O_1227,N_9550,N_9782);
xnor UO_1228 (O_1228,N_9636,N_9715);
nand UO_1229 (O_1229,N_9516,N_9616);
nand UO_1230 (O_1230,N_9981,N_9820);
nand UO_1231 (O_1231,N_9534,N_9538);
and UO_1232 (O_1232,N_9959,N_9990);
and UO_1233 (O_1233,N_9539,N_9763);
xnor UO_1234 (O_1234,N_9836,N_9899);
or UO_1235 (O_1235,N_9540,N_9555);
nand UO_1236 (O_1236,N_9615,N_9550);
nor UO_1237 (O_1237,N_9915,N_9669);
nor UO_1238 (O_1238,N_9776,N_9514);
xnor UO_1239 (O_1239,N_9656,N_9796);
xnor UO_1240 (O_1240,N_9612,N_9872);
nor UO_1241 (O_1241,N_9968,N_9884);
nand UO_1242 (O_1242,N_9668,N_9676);
nand UO_1243 (O_1243,N_9646,N_9897);
nand UO_1244 (O_1244,N_9650,N_9620);
nor UO_1245 (O_1245,N_9820,N_9654);
or UO_1246 (O_1246,N_9832,N_9866);
and UO_1247 (O_1247,N_9898,N_9788);
nand UO_1248 (O_1248,N_9990,N_9809);
nand UO_1249 (O_1249,N_9909,N_9931);
and UO_1250 (O_1250,N_9901,N_9668);
and UO_1251 (O_1251,N_9779,N_9673);
nor UO_1252 (O_1252,N_9968,N_9850);
nand UO_1253 (O_1253,N_9572,N_9716);
or UO_1254 (O_1254,N_9846,N_9623);
xnor UO_1255 (O_1255,N_9910,N_9513);
xnor UO_1256 (O_1256,N_9846,N_9793);
or UO_1257 (O_1257,N_9898,N_9959);
and UO_1258 (O_1258,N_9845,N_9635);
nor UO_1259 (O_1259,N_9680,N_9908);
and UO_1260 (O_1260,N_9657,N_9648);
or UO_1261 (O_1261,N_9792,N_9857);
and UO_1262 (O_1262,N_9879,N_9669);
and UO_1263 (O_1263,N_9524,N_9892);
xor UO_1264 (O_1264,N_9586,N_9980);
nor UO_1265 (O_1265,N_9526,N_9930);
nor UO_1266 (O_1266,N_9741,N_9562);
xnor UO_1267 (O_1267,N_9982,N_9750);
nand UO_1268 (O_1268,N_9930,N_9655);
or UO_1269 (O_1269,N_9615,N_9966);
nand UO_1270 (O_1270,N_9870,N_9506);
or UO_1271 (O_1271,N_9873,N_9802);
or UO_1272 (O_1272,N_9962,N_9941);
and UO_1273 (O_1273,N_9695,N_9884);
nand UO_1274 (O_1274,N_9721,N_9862);
and UO_1275 (O_1275,N_9881,N_9912);
nor UO_1276 (O_1276,N_9826,N_9922);
or UO_1277 (O_1277,N_9995,N_9773);
nor UO_1278 (O_1278,N_9873,N_9894);
xnor UO_1279 (O_1279,N_9842,N_9806);
nand UO_1280 (O_1280,N_9565,N_9588);
or UO_1281 (O_1281,N_9650,N_9811);
xnor UO_1282 (O_1282,N_9547,N_9875);
nand UO_1283 (O_1283,N_9846,N_9613);
xnor UO_1284 (O_1284,N_9608,N_9667);
and UO_1285 (O_1285,N_9702,N_9918);
nand UO_1286 (O_1286,N_9668,N_9845);
or UO_1287 (O_1287,N_9584,N_9913);
or UO_1288 (O_1288,N_9633,N_9836);
xnor UO_1289 (O_1289,N_9559,N_9734);
nor UO_1290 (O_1290,N_9809,N_9737);
nand UO_1291 (O_1291,N_9716,N_9602);
nor UO_1292 (O_1292,N_9570,N_9912);
xor UO_1293 (O_1293,N_9947,N_9525);
nor UO_1294 (O_1294,N_9833,N_9992);
or UO_1295 (O_1295,N_9948,N_9872);
xor UO_1296 (O_1296,N_9723,N_9610);
and UO_1297 (O_1297,N_9912,N_9682);
or UO_1298 (O_1298,N_9729,N_9681);
nand UO_1299 (O_1299,N_9703,N_9561);
nand UO_1300 (O_1300,N_9558,N_9994);
and UO_1301 (O_1301,N_9769,N_9651);
xnor UO_1302 (O_1302,N_9500,N_9622);
xnor UO_1303 (O_1303,N_9632,N_9891);
nand UO_1304 (O_1304,N_9922,N_9705);
xnor UO_1305 (O_1305,N_9928,N_9915);
nor UO_1306 (O_1306,N_9954,N_9925);
or UO_1307 (O_1307,N_9576,N_9854);
xor UO_1308 (O_1308,N_9668,N_9537);
nand UO_1309 (O_1309,N_9877,N_9631);
nand UO_1310 (O_1310,N_9699,N_9887);
and UO_1311 (O_1311,N_9530,N_9715);
nor UO_1312 (O_1312,N_9652,N_9871);
and UO_1313 (O_1313,N_9775,N_9821);
nor UO_1314 (O_1314,N_9661,N_9625);
and UO_1315 (O_1315,N_9765,N_9666);
or UO_1316 (O_1316,N_9873,N_9549);
nor UO_1317 (O_1317,N_9787,N_9515);
or UO_1318 (O_1318,N_9688,N_9992);
or UO_1319 (O_1319,N_9708,N_9785);
or UO_1320 (O_1320,N_9770,N_9527);
or UO_1321 (O_1321,N_9977,N_9685);
nor UO_1322 (O_1322,N_9966,N_9625);
nand UO_1323 (O_1323,N_9711,N_9964);
nor UO_1324 (O_1324,N_9855,N_9617);
nor UO_1325 (O_1325,N_9723,N_9806);
nor UO_1326 (O_1326,N_9649,N_9891);
and UO_1327 (O_1327,N_9731,N_9757);
xor UO_1328 (O_1328,N_9941,N_9999);
and UO_1329 (O_1329,N_9633,N_9585);
or UO_1330 (O_1330,N_9971,N_9987);
nand UO_1331 (O_1331,N_9798,N_9924);
or UO_1332 (O_1332,N_9619,N_9531);
nor UO_1333 (O_1333,N_9972,N_9948);
nand UO_1334 (O_1334,N_9705,N_9800);
xnor UO_1335 (O_1335,N_9908,N_9775);
nand UO_1336 (O_1336,N_9580,N_9538);
xnor UO_1337 (O_1337,N_9820,N_9642);
nor UO_1338 (O_1338,N_9764,N_9766);
and UO_1339 (O_1339,N_9666,N_9573);
nor UO_1340 (O_1340,N_9984,N_9669);
or UO_1341 (O_1341,N_9831,N_9857);
xnor UO_1342 (O_1342,N_9690,N_9837);
xor UO_1343 (O_1343,N_9827,N_9597);
xnor UO_1344 (O_1344,N_9591,N_9950);
nor UO_1345 (O_1345,N_9625,N_9916);
nor UO_1346 (O_1346,N_9747,N_9818);
nor UO_1347 (O_1347,N_9694,N_9991);
nand UO_1348 (O_1348,N_9827,N_9616);
xor UO_1349 (O_1349,N_9832,N_9760);
and UO_1350 (O_1350,N_9655,N_9587);
or UO_1351 (O_1351,N_9569,N_9771);
xnor UO_1352 (O_1352,N_9650,N_9886);
nor UO_1353 (O_1353,N_9942,N_9571);
or UO_1354 (O_1354,N_9723,N_9958);
nor UO_1355 (O_1355,N_9778,N_9900);
or UO_1356 (O_1356,N_9800,N_9819);
nand UO_1357 (O_1357,N_9802,N_9950);
nand UO_1358 (O_1358,N_9874,N_9816);
xnor UO_1359 (O_1359,N_9875,N_9876);
nor UO_1360 (O_1360,N_9515,N_9880);
or UO_1361 (O_1361,N_9742,N_9996);
xnor UO_1362 (O_1362,N_9908,N_9838);
or UO_1363 (O_1363,N_9712,N_9958);
and UO_1364 (O_1364,N_9549,N_9565);
xor UO_1365 (O_1365,N_9564,N_9633);
or UO_1366 (O_1366,N_9744,N_9581);
and UO_1367 (O_1367,N_9654,N_9954);
nor UO_1368 (O_1368,N_9619,N_9585);
nor UO_1369 (O_1369,N_9738,N_9912);
or UO_1370 (O_1370,N_9505,N_9522);
xor UO_1371 (O_1371,N_9937,N_9893);
and UO_1372 (O_1372,N_9721,N_9615);
or UO_1373 (O_1373,N_9527,N_9876);
nand UO_1374 (O_1374,N_9618,N_9687);
or UO_1375 (O_1375,N_9760,N_9691);
nand UO_1376 (O_1376,N_9506,N_9727);
nand UO_1377 (O_1377,N_9755,N_9823);
and UO_1378 (O_1378,N_9880,N_9841);
or UO_1379 (O_1379,N_9851,N_9980);
nand UO_1380 (O_1380,N_9747,N_9929);
or UO_1381 (O_1381,N_9646,N_9603);
and UO_1382 (O_1382,N_9872,N_9625);
or UO_1383 (O_1383,N_9573,N_9663);
nor UO_1384 (O_1384,N_9792,N_9564);
nor UO_1385 (O_1385,N_9785,N_9662);
nand UO_1386 (O_1386,N_9669,N_9810);
or UO_1387 (O_1387,N_9891,N_9748);
and UO_1388 (O_1388,N_9550,N_9878);
or UO_1389 (O_1389,N_9968,N_9943);
or UO_1390 (O_1390,N_9537,N_9773);
nor UO_1391 (O_1391,N_9626,N_9555);
nand UO_1392 (O_1392,N_9834,N_9668);
xnor UO_1393 (O_1393,N_9736,N_9641);
nor UO_1394 (O_1394,N_9818,N_9969);
xor UO_1395 (O_1395,N_9704,N_9879);
nor UO_1396 (O_1396,N_9706,N_9616);
or UO_1397 (O_1397,N_9872,N_9503);
and UO_1398 (O_1398,N_9701,N_9523);
xnor UO_1399 (O_1399,N_9543,N_9594);
xor UO_1400 (O_1400,N_9917,N_9500);
and UO_1401 (O_1401,N_9544,N_9852);
and UO_1402 (O_1402,N_9603,N_9774);
and UO_1403 (O_1403,N_9744,N_9924);
nor UO_1404 (O_1404,N_9952,N_9573);
nand UO_1405 (O_1405,N_9751,N_9740);
xnor UO_1406 (O_1406,N_9669,N_9625);
nand UO_1407 (O_1407,N_9652,N_9672);
and UO_1408 (O_1408,N_9886,N_9683);
xnor UO_1409 (O_1409,N_9994,N_9712);
or UO_1410 (O_1410,N_9528,N_9520);
and UO_1411 (O_1411,N_9836,N_9849);
and UO_1412 (O_1412,N_9531,N_9993);
nand UO_1413 (O_1413,N_9547,N_9688);
nor UO_1414 (O_1414,N_9972,N_9907);
nand UO_1415 (O_1415,N_9996,N_9859);
nand UO_1416 (O_1416,N_9875,N_9822);
nand UO_1417 (O_1417,N_9651,N_9851);
nand UO_1418 (O_1418,N_9584,N_9664);
xnor UO_1419 (O_1419,N_9533,N_9965);
nor UO_1420 (O_1420,N_9714,N_9961);
or UO_1421 (O_1421,N_9770,N_9525);
or UO_1422 (O_1422,N_9536,N_9865);
or UO_1423 (O_1423,N_9508,N_9505);
and UO_1424 (O_1424,N_9995,N_9990);
nor UO_1425 (O_1425,N_9581,N_9826);
xnor UO_1426 (O_1426,N_9925,N_9875);
and UO_1427 (O_1427,N_9974,N_9716);
and UO_1428 (O_1428,N_9752,N_9980);
nand UO_1429 (O_1429,N_9723,N_9715);
nor UO_1430 (O_1430,N_9956,N_9793);
nand UO_1431 (O_1431,N_9702,N_9805);
nor UO_1432 (O_1432,N_9970,N_9809);
nor UO_1433 (O_1433,N_9567,N_9596);
or UO_1434 (O_1434,N_9675,N_9904);
nand UO_1435 (O_1435,N_9633,N_9703);
and UO_1436 (O_1436,N_9657,N_9756);
nor UO_1437 (O_1437,N_9839,N_9713);
nand UO_1438 (O_1438,N_9714,N_9843);
and UO_1439 (O_1439,N_9667,N_9943);
or UO_1440 (O_1440,N_9656,N_9936);
xnor UO_1441 (O_1441,N_9955,N_9923);
xor UO_1442 (O_1442,N_9703,N_9994);
nor UO_1443 (O_1443,N_9766,N_9513);
and UO_1444 (O_1444,N_9518,N_9814);
nor UO_1445 (O_1445,N_9611,N_9969);
and UO_1446 (O_1446,N_9623,N_9881);
xor UO_1447 (O_1447,N_9702,N_9524);
and UO_1448 (O_1448,N_9690,N_9554);
or UO_1449 (O_1449,N_9763,N_9835);
nor UO_1450 (O_1450,N_9790,N_9912);
nor UO_1451 (O_1451,N_9684,N_9693);
nand UO_1452 (O_1452,N_9783,N_9829);
and UO_1453 (O_1453,N_9552,N_9788);
xnor UO_1454 (O_1454,N_9545,N_9645);
xnor UO_1455 (O_1455,N_9780,N_9544);
nor UO_1456 (O_1456,N_9595,N_9977);
or UO_1457 (O_1457,N_9845,N_9835);
and UO_1458 (O_1458,N_9559,N_9931);
and UO_1459 (O_1459,N_9844,N_9975);
nor UO_1460 (O_1460,N_9803,N_9774);
or UO_1461 (O_1461,N_9513,N_9707);
and UO_1462 (O_1462,N_9975,N_9999);
and UO_1463 (O_1463,N_9988,N_9671);
and UO_1464 (O_1464,N_9668,N_9865);
nand UO_1465 (O_1465,N_9815,N_9584);
and UO_1466 (O_1466,N_9897,N_9747);
nand UO_1467 (O_1467,N_9867,N_9629);
or UO_1468 (O_1468,N_9855,N_9516);
xnor UO_1469 (O_1469,N_9770,N_9655);
and UO_1470 (O_1470,N_9603,N_9516);
nand UO_1471 (O_1471,N_9797,N_9710);
nand UO_1472 (O_1472,N_9817,N_9745);
nor UO_1473 (O_1473,N_9987,N_9963);
nor UO_1474 (O_1474,N_9686,N_9850);
and UO_1475 (O_1475,N_9685,N_9743);
nor UO_1476 (O_1476,N_9625,N_9566);
or UO_1477 (O_1477,N_9595,N_9774);
or UO_1478 (O_1478,N_9614,N_9858);
nor UO_1479 (O_1479,N_9867,N_9838);
nand UO_1480 (O_1480,N_9956,N_9714);
xnor UO_1481 (O_1481,N_9636,N_9526);
xnor UO_1482 (O_1482,N_9809,N_9812);
nand UO_1483 (O_1483,N_9779,N_9955);
nor UO_1484 (O_1484,N_9760,N_9926);
or UO_1485 (O_1485,N_9721,N_9897);
xor UO_1486 (O_1486,N_9823,N_9701);
or UO_1487 (O_1487,N_9595,N_9577);
and UO_1488 (O_1488,N_9939,N_9985);
nor UO_1489 (O_1489,N_9507,N_9850);
xor UO_1490 (O_1490,N_9803,N_9682);
nor UO_1491 (O_1491,N_9572,N_9820);
or UO_1492 (O_1492,N_9955,N_9712);
or UO_1493 (O_1493,N_9728,N_9583);
and UO_1494 (O_1494,N_9681,N_9513);
and UO_1495 (O_1495,N_9911,N_9752);
xor UO_1496 (O_1496,N_9738,N_9785);
xor UO_1497 (O_1497,N_9737,N_9810);
and UO_1498 (O_1498,N_9553,N_9965);
xnor UO_1499 (O_1499,N_9588,N_9879);
endmodule