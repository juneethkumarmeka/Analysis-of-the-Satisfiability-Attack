module basic_750_5000_1000_2_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2530,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2560,N_2562,N_2564,N_2565,N_2567,N_2569,N_2570,N_2572,N_2574,N_2576,N_2578,N_2579,N_2580,N_2581,N_2583,N_2584,N_2585,N_2586,N_2588,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2636,N_2640,N_2642,N_2643,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2659,N_2660,N_2662,N_2663,N_2664,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2694,N_2695,N_2696,N_2699,N_2700,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2710,N_2711,N_2713,N_2714,N_2716,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2727,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2748,N_2749,N_2750,N_2751,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2760,N_2762,N_2763,N_2764,N_2765,N_2766,N_2768,N_2769,N_2771,N_2773,N_2774,N_2775,N_2777,N_2778,N_2779,N_2782,N_2783,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2792,N_2793,N_2795,N_2796,N_2797,N_2798,N_2799,N_2801,N_2802,N_2803,N_2804,N_2805,N_2807,N_2809,N_2811,N_2812,N_2813,N_2814,N_2816,N_2817,N_2818,N_2820,N_2821,N_2822,N_2823,N_2824,N_2827,N_2828,N_2829,N_2831,N_2832,N_2833,N_2834,N_2835,N_2838,N_2839,N_2840,N_2841,N_2842,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2869,N_2870,N_2871,N_2872,N_2873,N_2875,N_2876,N_2877,N_2878,N_2880,N_2881,N_2884,N_2885,N_2886,N_2887,N_2888,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2933,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2943,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2955,N_2956,N_2957,N_2958,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2971,N_2972,N_2973,N_2974,N_2977,N_2979,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2990,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3034,N_3035,N_3036,N_3037,N_3038,N_3040,N_3041,N_3042,N_3043,N_3044,N_3046,N_3047,N_3048,N_3049,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3067,N_3068,N_3069,N_3070,N_3071,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3081,N_3082,N_3083,N_3084,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3095,N_3096,N_3097,N_3098,N_3099,N_3101,N_3103,N_3104,N_3105,N_3106,N_3107,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3117,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3131,N_3132,N_3133,N_3134,N_3135,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3172,N_3173,N_3174,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3184,N_3186,N_3187,N_3188,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3200,N_3201,N_3202,N_3203,N_3205,N_3206,N_3207,N_3208,N_3210,N_3211,N_3212,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3230,N_3231,N_3232,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3263,N_3264,N_3266,N_3267,N_3268,N_3269,N_3272,N_3273,N_3274,N_3275,N_3277,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3298,N_3299,N_3300,N_3301,N_3303,N_3304,N_3305,N_3306,N_3308,N_3309,N_3310,N_3311,N_3313,N_3314,N_3316,N_3317,N_3319,N_3321,N_3323,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3340,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3363,N_3364,N_3365,N_3367,N_3368,N_3369,N_3371,N_3372,N_3373,N_3374,N_3375,N_3377,N_3378,N_3380,N_3381,N_3382,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3414,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3429,N_3430,N_3431,N_3432,N_3434,N_3435,N_3437,N_3438,N_3440,N_3441,N_3442,N_3443,N_3444,N_3446,N_3448,N_3449,N_3450,N_3451,N_3452,N_3454,N_3455,N_3457,N_3458,N_3459,N_3461,N_3462,N_3463,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3472,N_3473,N_3474,N_3476,N_3477,N_3478,N_3479,N_3480,N_3482,N_3483,N_3484,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3494,N_3495,N_3496,N_3497,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3508,N_3509,N_3510,N_3512,N_3513,N_3514,N_3515,N_3517,N_3518,N_3519,N_3520,N_3521,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3533,N_3535,N_3538,N_3539,N_3541,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3554,N_3555,N_3557,N_3558,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3572,N_3573,N_3574,N_3575,N_3577,N_3578,N_3580,N_3582,N_3586,N_3587,N_3589,N_3590,N_3592,N_3593,N_3594,N_3595,N_3597,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3661,N_3662,N_3663,N_3664,N_3665,N_3667,N_3668,N_3671,N_3672,N_3674,N_3675,N_3676,N_3679,N_3680,N_3681,N_3682,N_3684,N_3685,N_3687,N_3691,N_3692,N_3697,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3707,N_3708,N_3709,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3730,N_3732,N_3734,N_3736,N_3737,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3747,N_3749,N_3750,N_3751,N_3752,N_3753,N_3755,N_3756,N_3757,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3769,N_3770,N_3771,N_3772,N_3773,N_3775,N_3776,N_3777,N_3779,N_3780,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3792,N_3793,N_3794,N_3795,N_3797,N_3798,N_3799,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3811,N_3813,N_3815,N_3816,N_3817,N_3820,N_3821,N_3822,N_3823,N_3825,N_3826,N_3828,N_3829,N_3831,N_3832,N_3835,N_3836,N_3837,N_3839,N_3842,N_3843,N_3844,N_3845,N_3846,N_3848,N_3849,N_3850,N_3851,N_3855,N_3858,N_3859,N_3861,N_3862,N_3863,N_3865,N_3866,N_3867,N_3868,N_3870,N_3872,N_3873,N_3874,N_3875,N_3876,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3896,N_3897,N_3898,N_3901,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3965,N_3966,N_3968,N_3969,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3979,N_3980,N_3981,N_3983,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_4000,N_4001,N_4002,N_4003,N_4007,N_4008,N_4009,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4019,N_4020,N_4021,N_4023,N_4025,N_4026,N_4027,N_4028,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4041,N_4042,N_4044,N_4046,N_4047,N_4048,N_4049,N_4050,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4073,N_4074,N_4075,N_4076,N_4079,N_4080,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4161,N_4164,N_4165,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4180,N_4181,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4200,N_4201,N_4202,N_4203,N_4205,N_4206,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4219,N_4220,N_4221,N_4222,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4239,N_4241,N_4242,N_4243,N_4244,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4257,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4294,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4320,N_4321,N_4322,N_4323,N_4324,N_4326,N_4327,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4353,N_4354,N_4356,N_4357,N_4358,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4370,N_4372,N_4373,N_4375,N_4377,N_4378,N_4379,N_4380,N_4381,N_4383,N_4385,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4396,N_4397,N_4398,N_4399,N_4400,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4410,N_4411,N_4412,N_4413,N_4415,N_4417,N_4418,N_4419,N_4420,N_4422,N_4423,N_4425,N_4427,N_4430,N_4431,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4454,N_4455,N_4456,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4475,N_4477,N_4478,N_4479,N_4480,N_4481,N_4483,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4525,N_4526,N_4528,N_4529,N_4531,N_4532,N_4535,N_4537,N_4538,N_4540,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4555,N_4556,N_4557,N_4560,N_4561,N_4562,N_4563,N_4566,N_4567,N_4568,N_4569,N_4570,N_4572,N_4573,N_4574,N_4576,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4601,N_4602,N_4603,N_4608,N_4610,N_4611,N_4612,N_4613,N_4614,N_4616,N_4617,N_4618,N_4620,N_4621,N_4622,N_4624,N_4626,N_4627,N_4628,N_4630,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4641,N_4642,N_4644,N_4645,N_4646,N_4650,N_4652,N_4653,N_4654,N_4655,N_4656,N_4658,N_4659,N_4660,N_4661,N_4662,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4675,N_4676,N_4677,N_4678,N_4679,N_4681,N_4682,N_4683,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4693,N_4695,N_4696,N_4697,N_4698,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4718,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4739,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4750,N_4753,N_4754,N_4756,N_4759,N_4760,N_4761,N_4763,N_4767,N_4768,N_4769,N_4770,N_4771,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4782,N_4783,N_4785,N_4786,N_4787,N_4789,N_4790,N_4791,N_4792,N_4794,N_4795,N_4796,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4807,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4823,N_4825,N_4826,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4836,N_4837,N_4838,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4853,N_4857,N_4859,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4870,N_4872,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4890,N_4891,N_4893,N_4894,N_4897,N_4898,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4907,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4917,N_4918,N_4919,N_4920,N_4921,N_4923,N_4924,N_4925,N_4927,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4941,N_4942,N_4944,N_4945,N_4946,N_4947,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4970,N_4974,N_4975,N_4976,N_4979,N_4980,N_4982,N_4983,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_551,In_332);
nand U1 (N_1,In_596,In_726);
nor U2 (N_2,In_627,In_443);
nor U3 (N_3,In_31,In_734);
or U4 (N_4,In_529,In_167);
and U5 (N_5,In_483,In_188);
or U6 (N_6,In_418,In_24);
nor U7 (N_7,In_697,In_170);
and U8 (N_8,In_121,In_306);
and U9 (N_9,In_222,In_336);
and U10 (N_10,In_146,In_374);
and U11 (N_11,In_407,In_380);
nor U12 (N_12,In_67,In_581);
nand U13 (N_13,In_703,In_609);
and U14 (N_14,In_244,In_197);
and U15 (N_15,In_605,In_722);
or U16 (N_16,In_702,In_710);
nor U17 (N_17,In_484,In_232);
or U18 (N_18,In_216,In_355);
nor U19 (N_19,In_591,In_59);
and U20 (N_20,In_562,In_308);
or U21 (N_21,In_60,In_607);
xor U22 (N_22,In_158,In_471);
and U23 (N_23,In_61,In_177);
nor U24 (N_24,In_310,In_419);
and U25 (N_25,In_79,In_587);
and U26 (N_26,In_674,In_364);
nand U27 (N_27,In_223,In_494);
nor U28 (N_28,In_331,In_185);
nor U29 (N_29,In_112,In_558);
or U30 (N_30,In_745,In_454);
xor U31 (N_31,In_486,In_150);
nand U32 (N_32,In_26,In_267);
or U33 (N_33,In_462,In_39);
nand U34 (N_34,In_709,In_394);
or U35 (N_35,In_523,In_516);
nand U36 (N_36,In_472,In_157);
or U37 (N_37,In_594,In_744);
nand U38 (N_38,In_598,In_725);
nand U39 (N_39,In_208,In_700);
and U40 (N_40,In_47,In_411);
nor U41 (N_41,In_625,In_429);
or U42 (N_42,In_708,In_283);
and U43 (N_43,In_451,In_230);
nand U44 (N_44,In_477,In_329);
nand U45 (N_45,In_300,In_143);
or U46 (N_46,In_320,In_425);
nand U47 (N_47,In_475,In_48);
nor U48 (N_48,In_437,In_186);
or U49 (N_49,In_438,In_126);
nor U50 (N_50,In_651,In_388);
and U51 (N_51,In_560,In_108);
or U52 (N_52,In_162,In_246);
or U53 (N_53,In_730,In_402);
nor U54 (N_54,In_637,In_314);
nand U55 (N_55,In_18,In_219);
and U56 (N_56,In_473,In_271);
nor U57 (N_57,In_145,In_553);
and U58 (N_58,In_455,In_171);
and U59 (N_59,In_288,In_272);
or U60 (N_60,In_19,In_420);
nand U61 (N_61,In_628,In_559);
nand U62 (N_62,In_317,In_716);
nor U63 (N_63,In_589,In_362);
nor U64 (N_64,In_220,In_623);
and U65 (N_65,In_55,In_128);
and U66 (N_66,In_650,In_514);
and U67 (N_67,In_225,In_673);
nor U68 (N_68,In_554,In_528);
or U69 (N_69,In_139,In_34);
and U70 (N_70,In_301,In_262);
nor U71 (N_71,In_508,In_17);
nand U72 (N_72,In_511,In_612);
xnor U73 (N_73,In_292,In_382);
and U74 (N_74,In_692,In_37);
nand U75 (N_75,In_298,In_487);
nand U76 (N_76,In_346,In_735);
and U77 (N_77,In_504,In_182);
nor U78 (N_78,In_480,In_82);
and U79 (N_79,In_743,In_668);
or U80 (N_80,In_287,In_657);
or U81 (N_81,In_226,In_415);
nand U82 (N_82,In_236,In_600);
or U83 (N_83,In_42,In_379);
and U84 (N_84,In_681,In_384);
xnor U85 (N_85,In_187,In_638);
or U86 (N_86,In_72,In_662);
and U87 (N_87,In_369,In_10);
or U88 (N_88,In_166,In_100);
nor U89 (N_89,In_421,In_712);
or U90 (N_90,In_196,In_720);
nand U91 (N_91,In_290,In_169);
nor U92 (N_92,In_238,In_180);
and U93 (N_93,In_80,In_248);
nor U94 (N_94,In_647,In_493);
xor U95 (N_95,In_205,In_165);
or U96 (N_96,In_5,In_105);
or U97 (N_97,In_123,In_655);
or U98 (N_98,In_547,In_740);
nand U99 (N_99,In_356,In_168);
nand U100 (N_100,In_583,In_8);
or U101 (N_101,In_111,In_87);
and U102 (N_102,In_159,In_84);
and U103 (N_103,In_328,In_684);
or U104 (N_104,In_466,In_36);
and U105 (N_105,In_95,In_531);
and U106 (N_106,In_184,In_535);
nand U107 (N_107,In_467,In_445);
xor U108 (N_108,In_601,In_335);
and U109 (N_109,In_218,In_40);
and U110 (N_110,In_505,In_77);
and U111 (N_111,In_566,In_91);
nor U112 (N_112,In_255,In_303);
and U113 (N_113,In_405,In_142);
or U114 (N_114,In_237,In_387);
or U115 (N_115,In_358,In_253);
and U116 (N_116,In_330,In_731);
and U117 (N_117,In_400,In_497);
or U118 (N_118,In_416,In_198);
or U119 (N_119,In_254,In_339);
or U120 (N_120,In_319,In_570);
nand U121 (N_121,In_27,In_231);
nor U122 (N_122,In_406,In_682);
and U123 (N_123,In_663,In_93);
and U124 (N_124,In_643,In_620);
nand U125 (N_125,In_422,In_389);
and U126 (N_126,In_491,In_214);
and U127 (N_127,In_639,In_541);
and U128 (N_128,In_259,In_488);
nor U129 (N_129,In_327,In_615);
nand U130 (N_130,In_440,In_353);
and U131 (N_131,In_349,In_545);
and U132 (N_132,In_586,In_434);
xnor U133 (N_133,In_579,In_447);
nor U134 (N_134,In_699,In_45);
nor U135 (N_135,In_565,In_83);
or U136 (N_136,In_536,In_64);
nand U137 (N_137,In_33,In_106);
nor U138 (N_138,In_574,In_593);
nand U139 (N_139,In_468,In_334);
and U140 (N_140,In_485,In_132);
nor U141 (N_141,In_144,In_360);
nor U142 (N_142,In_137,In_441);
nor U143 (N_143,In_469,In_608);
nor U144 (N_144,In_599,In_245);
nand U145 (N_145,In_456,In_713);
nor U146 (N_146,In_147,In_11);
or U147 (N_147,In_432,In_696);
nand U148 (N_148,In_277,In_107);
or U149 (N_149,In_66,In_474);
nor U150 (N_150,In_706,In_526);
or U151 (N_151,In_660,In_359);
nor U152 (N_152,In_133,In_191);
or U153 (N_153,In_739,In_211);
xor U154 (N_154,In_148,In_385);
nor U155 (N_155,In_20,In_705);
nand U156 (N_156,In_375,In_124);
nand U157 (N_157,In_575,In_74);
or U158 (N_158,In_172,In_351);
nand U159 (N_159,In_96,In_717);
nand U160 (N_160,In_741,In_311);
or U161 (N_161,In_324,In_120);
and U162 (N_162,In_52,In_3);
nor U163 (N_163,In_683,In_548);
and U164 (N_164,In_632,In_645);
nand U165 (N_165,In_229,In_458);
and U166 (N_166,In_410,In_85);
nor U167 (N_167,In_373,In_302);
and U168 (N_168,In_264,In_496);
and U169 (N_169,In_179,In_436);
nor U170 (N_170,In_664,In_156);
nand U171 (N_171,In_109,In_749);
nand U172 (N_172,In_53,In_478);
nand U173 (N_173,In_41,In_688);
and U174 (N_174,In_280,In_14);
and U175 (N_175,In_368,In_687);
and U176 (N_176,In_338,In_397);
nor U177 (N_177,In_669,In_430);
nand U178 (N_178,In_403,In_517);
or U179 (N_179,In_54,In_195);
and U180 (N_180,In_695,In_6);
and U181 (N_181,In_733,In_178);
or U182 (N_182,In_518,In_727);
or U183 (N_183,In_190,In_648);
or U184 (N_184,In_715,In_701);
and U185 (N_185,In_213,In_401);
or U186 (N_186,In_318,In_439);
and U187 (N_187,In_16,In_103);
or U188 (N_188,In_435,In_240);
or U189 (N_189,In_527,In_649);
nand U190 (N_190,In_585,In_341);
nand U191 (N_191,In_260,In_21);
nor U192 (N_192,In_44,In_426);
or U193 (N_193,In_653,In_544);
and U194 (N_194,In_312,In_32);
nor U195 (N_195,In_621,In_141);
nand U196 (N_196,In_130,In_427);
nand U197 (N_197,In_577,In_689);
and U198 (N_198,In_134,In_204);
or U199 (N_199,In_125,In_665);
nand U200 (N_200,In_69,In_537);
nand U201 (N_201,In_452,In_619);
and U202 (N_202,In_556,In_630);
nor U203 (N_203,In_611,In_610);
nor U204 (N_204,In_275,In_568);
or U205 (N_205,In_194,In_381);
and U206 (N_206,In_297,In_424);
nor U207 (N_207,In_580,In_719);
nor U208 (N_208,In_299,In_578);
nor U209 (N_209,In_352,In_136);
and U210 (N_210,In_393,In_73);
or U211 (N_211,In_366,In_263);
and U212 (N_212,In_686,In_258);
nor U213 (N_213,In_489,In_256);
nor U214 (N_214,In_667,In_470);
and U215 (N_215,In_294,In_707);
nor U216 (N_216,In_652,In_476);
nor U217 (N_217,In_378,In_398);
nand U218 (N_218,In_1,In_461);
or U219 (N_219,In_433,In_671);
nand U220 (N_220,In_636,In_646);
nand U221 (N_221,In_365,In_659);
nand U222 (N_222,In_233,In_606);
or U223 (N_223,In_293,In_588);
nor U224 (N_224,In_274,In_465);
and U225 (N_225,In_370,In_654);
nor U226 (N_226,In_68,In_78);
nand U227 (N_227,In_65,In_295);
nand U228 (N_228,In_386,In_573);
nor U229 (N_229,In_738,In_503);
nor U230 (N_230,In_325,In_183);
xor U231 (N_231,In_509,In_428);
and U232 (N_232,In_448,In_155);
and U233 (N_233,In_92,In_110);
nor U234 (N_234,In_285,In_383);
or U235 (N_235,In_313,In_296);
or U236 (N_236,In_323,In_576);
or U237 (N_237,In_404,In_506);
or U238 (N_238,In_367,In_521);
nand U239 (N_239,In_391,In_519);
nand U240 (N_240,In_261,In_75);
and U241 (N_241,In_71,In_135);
or U242 (N_242,In_289,In_498);
nor U243 (N_243,In_101,In_492);
or U244 (N_244,In_515,In_685);
or U245 (N_245,In_337,In_315);
nor U246 (N_246,In_412,In_193);
or U247 (N_247,In_676,In_98);
and U248 (N_248,In_115,In_546);
or U249 (N_249,In_634,In_502);
nand U250 (N_250,In_266,In_217);
nor U251 (N_251,In_460,In_13);
or U252 (N_252,In_538,In_203);
nand U253 (N_253,In_631,In_43);
nand U254 (N_254,In_242,In_464);
or U255 (N_255,In_520,In_282);
and U256 (N_256,In_113,In_736);
nand U257 (N_257,In_181,In_495);
nor U258 (N_258,In_616,In_131);
nand U259 (N_259,In_626,In_446);
nor U260 (N_260,In_513,In_28);
nor U261 (N_261,In_279,In_678);
or U262 (N_262,In_542,In_206);
and U263 (N_263,In_201,In_62);
nor U264 (N_264,In_119,In_698);
or U265 (N_265,In_58,In_343);
nor U266 (N_266,In_189,In_561);
nor U267 (N_267,In_149,In_500);
nand U268 (N_268,In_291,In_25);
nand U269 (N_269,In_450,In_199);
nand U270 (N_270,In_152,In_215);
nor U271 (N_271,In_510,In_633);
or U272 (N_272,In_724,In_340);
nand U273 (N_273,In_89,In_56);
and U274 (N_274,In_549,In_9);
nor U275 (N_275,In_613,In_164);
and U276 (N_276,In_463,In_661);
nor U277 (N_277,In_552,In_129);
nand U278 (N_278,In_539,In_658);
or U279 (N_279,In_209,In_249);
nand U280 (N_280,In_677,In_200);
and U281 (N_281,In_563,In_224);
or U282 (N_282,In_390,In_540);
and U283 (N_283,In_276,In_442);
or U284 (N_284,In_22,In_250);
and U285 (N_285,In_675,In_748);
and U286 (N_286,In_592,In_278);
nand U287 (N_287,In_481,In_742);
nor U288 (N_288,In_641,In_63);
and U289 (N_289,In_102,In_522);
nand U290 (N_290,In_507,In_624);
nand U291 (N_291,In_371,In_670);
and U292 (N_292,In_714,In_163);
and U293 (N_293,In_499,In_414);
and U294 (N_294,In_679,In_88);
or U295 (N_295,In_543,In_114);
nor U296 (N_296,In_691,In_690);
or U297 (N_297,In_732,In_345);
and U298 (N_298,In_363,In_617);
or U299 (N_299,In_76,In_618);
xnor U300 (N_300,In_417,In_431);
nand U301 (N_301,In_457,In_550);
nand U302 (N_302,In_304,In_81);
and U303 (N_303,In_23,In_333);
and U304 (N_304,In_729,In_269);
nor U305 (N_305,In_192,In_251);
nor U306 (N_306,In_118,In_555);
or U307 (N_307,In_265,In_525);
or U308 (N_308,In_326,In_392);
nand U309 (N_309,In_30,In_512);
nor U310 (N_310,In_396,In_252);
xnor U311 (N_311,In_127,In_449);
nand U312 (N_312,In_409,In_604);
and U313 (N_313,In_117,In_737);
or U314 (N_314,In_357,In_322);
and U315 (N_315,In_728,In_140);
xor U316 (N_316,In_622,In_413);
and U317 (N_317,In_372,In_656);
nor U318 (N_318,In_51,In_453);
nand U319 (N_319,In_247,In_597);
or U320 (N_320,In_35,In_70);
and U321 (N_321,In_174,In_0);
nand U322 (N_322,In_482,In_490);
nor U323 (N_323,In_97,In_395);
nor U324 (N_324,In_138,In_361);
or U325 (N_325,In_635,In_582);
nand U326 (N_326,In_234,In_344);
and U327 (N_327,In_342,In_533);
or U328 (N_328,In_569,In_29);
nand U329 (N_329,In_273,In_99);
or U330 (N_330,In_694,In_644);
xnor U331 (N_331,In_321,In_747);
or U332 (N_332,In_672,In_104);
nor U333 (N_333,In_399,In_15);
nand U334 (N_334,In_12,In_239);
and U335 (N_335,In_268,In_316);
nor U336 (N_336,In_86,In_564);
nand U337 (N_337,In_210,In_348);
and U338 (N_338,In_584,In_602);
xor U339 (N_339,In_284,In_746);
nand U340 (N_340,In_642,In_680);
nor U341 (N_341,In_595,In_666);
or U342 (N_342,In_305,In_235);
nand U343 (N_343,In_444,In_202);
or U344 (N_344,In_286,In_241);
and U345 (N_345,In_173,In_501);
or U346 (N_346,In_49,In_459);
nand U347 (N_347,In_94,In_603);
nand U348 (N_348,In_270,In_376);
nand U349 (N_349,In_161,In_7);
nand U350 (N_350,In_704,In_154);
or U351 (N_351,In_524,In_567);
or U352 (N_352,In_307,In_711);
nor U353 (N_353,In_423,In_350);
or U354 (N_354,In_571,In_723);
nand U355 (N_355,In_175,In_377);
or U356 (N_356,In_281,In_153);
nand U357 (N_357,In_354,In_629);
xnor U358 (N_358,In_176,In_160);
nor U359 (N_359,In_572,In_212);
nand U360 (N_360,In_122,In_530);
nor U361 (N_361,In_557,In_693);
nand U362 (N_362,In_4,In_532);
or U363 (N_363,In_309,In_640);
or U364 (N_364,In_347,In_614);
and U365 (N_365,In_408,In_207);
nor U366 (N_366,In_151,In_57);
nand U367 (N_367,In_479,In_116);
nor U368 (N_368,In_50,In_228);
nand U369 (N_369,In_718,In_257);
nand U370 (N_370,In_2,In_46);
xor U371 (N_371,In_90,In_721);
and U372 (N_372,In_590,In_38);
or U373 (N_373,In_227,In_534);
nand U374 (N_374,In_243,In_221);
nor U375 (N_375,In_163,In_65);
nand U376 (N_376,In_536,In_200);
or U377 (N_377,In_133,In_729);
and U378 (N_378,In_507,In_163);
and U379 (N_379,In_53,In_179);
nand U380 (N_380,In_711,In_498);
nor U381 (N_381,In_669,In_595);
or U382 (N_382,In_114,In_257);
or U383 (N_383,In_83,In_496);
or U384 (N_384,In_305,In_316);
and U385 (N_385,In_675,In_471);
and U386 (N_386,In_651,In_708);
or U387 (N_387,In_602,In_512);
or U388 (N_388,In_619,In_719);
and U389 (N_389,In_686,In_208);
nor U390 (N_390,In_622,In_183);
and U391 (N_391,In_346,In_182);
xnor U392 (N_392,In_423,In_358);
nand U393 (N_393,In_23,In_577);
and U394 (N_394,In_380,In_124);
and U395 (N_395,In_569,In_261);
nor U396 (N_396,In_159,In_655);
or U397 (N_397,In_552,In_566);
and U398 (N_398,In_275,In_449);
and U399 (N_399,In_342,In_226);
or U400 (N_400,In_534,In_704);
and U401 (N_401,In_10,In_391);
and U402 (N_402,In_551,In_305);
and U403 (N_403,In_49,In_607);
nor U404 (N_404,In_285,In_641);
or U405 (N_405,In_499,In_205);
nor U406 (N_406,In_249,In_538);
nand U407 (N_407,In_9,In_256);
and U408 (N_408,In_182,In_299);
and U409 (N_409,In_647,In_7);
nand U410 (N_410,In_482,In_445);
nand U411 (N_411,In_155,In_457);
nand U412 (N_412,In_708,In_121);
and U413 (N_413,In_323,In_249);
nand U414 (N_414,In_205,In_54);
nor U415 (N_415,In_501,In_196);
nand U416 (N_416,In_215,In_524);
nand U417 (N_417,In_2,In_458);
nor U418 (N_418,In_205,In_713);
or U419 (N_419,In_547,In_643);
and U420 (N_420,In_545,In_265);
and U421 (N_421,In_43,In_11);
nand U422 (N_422,In_386,In_48);
nand U423 (N_423,In_598,In_488);
nand U424 (N_424,In_340,In_279);
nand U425 (N_425,In_10,In_683);
nor U426 (N_426,In_535,In_449);
and U427 (N_427,In_333,In_496);
nor U428 (N_428,In_648,In_131);
xor U429 (N_429,In_499,In_236);
or U430 (N_430,In_701,In_345);
and U431 (N_431,In_400,In_700);
nand U432 (N_432,In_67,In_428);
and U433 (N_433,In_705,In_189);
or U434 (N_434,In_93,In_95);
nor U435 (N_435,In_194,In_653);
nand U436 (N_436,In_679,In_321);
or U437 (N_437,In_170,In_554);
or U438 (N_438,In_448,In_239);
nand U439 (N_439,In_23,In_649);
nand U440 (N_440,In_274,In_471);
or U441 (N_441,In_569,In_353);
or U442 (N_442,In_289,In_269);
or U443 (N_443,In_66,In_528);
nand U444 (N_444,In_265,In_520);
nand U445 (N_445,In_207,In_653);
nand U446 (N_446,In_700,In_369);
nand U447 (N_447,In_95,In_194);
nand U448 (N_448,In_374,In_650);
and U449 (N_449,In_388,In_615);
and U450 (N_450,In_584,In_200);
nor U451 (N_451,In_537,In_125);
and U452 (N_452,In_544,In_575);
or U453 (N_453,In_180,In_195);
nor U454 (N_454,In_459,In_122);
nor U455 (N_455,In_413,In_134);
and U456 (N_456,In_245,In_615);
and U457 (N_457,In_526,In_412);
and U458 (N_458,In_639,In_733);
or U459 (N_459,In_736,In_138);
nand U460 (N_460,In_627,In_226);
nor U461 (N_461,In_27,In_540);
and U462 (N_462,In_183,In_383);
nor U463 (N_463,In_2,In_490);
or U464 (N_464,In_550,In_353);
nor U465 (N_465,In_148,In_205);
xnor U466 (N_466,In_332,In_1);
nand U467 (N_467,In_217,In_653);
or U468 (N_468,In_64,In_486);
or U469 (N_469,In_393,In_291);
nor U470 (N_470,In_20,In_451);
nor U471 (N_471,In_252,In_672);
and U472 (N_472,In_616,In_612);
or U473 (N_473,In_317,In_417);
and U474 (N_474,In_545,In_75);
and U475 (N_475,In_728,In_156);
or U476 (N_476,In_31,In_105);
nand U477 (N_477,In_611,In_469);
or U478 (N_478,In_164,In_172);
nor U479 (N_479,In_483,In_424);
or U480 (N_480,In_356,In_602);
and U481 (N_481,In_439,In_420);
nand U482 (N_482,In_170,In_487);
nor U483 (N_483,In_135,In_639);
nand U484 (N_484,In_669,In_32);
and U485 (N_485,In_45,In_539);
nand U486 (N_486,In_566,In_212);
nor U487 (N_487,In_740,In_719);
nand U488 (N_488,In_564,In_39);
nand U489 (N_489,In_431,In_146);
xnor U490 (N_490,In_529,In_729);
and U491 (N_491,In_474,In_48);
nor U492 (N_492,In_56,In_309);
nor U493 (N_493,In_672,In_500);
and U494 (N_494,In_82,In_460);
nand U495 (N_495,In_277,In_298);
or U496 (N_496,In_730,In_557);
and U497 (N_497,In_309,In_79);
and U498 (N_498,In_625,In_445);
and U499 (N_499,In_4,In_196);
nand U500 (N_500,In_475,In_148);
nand U501 (N_501,In_88,In_547);
or U502 (N_502,In_670,In_555);
and U503 (N_503,In_369,In_246);
and U504 (N_504,In_445,In_648);
nand U505 (N_505,In_707,In_138);
nand U506 (N_506,In_544,In_342);
nand U507 (N_507,In_621,In_317);
nand U508 (N_508,In_558,In_525);
and U509 (N_509,In_485,In_622);
nor U510 (N_510,In_382,In_646);
or U511 (N_511,In_529,In_393);
nor U512 (N_512,In_183,In_163);
nor U513 (N_513,In_382,In_99);
or U514 (N_514,In_621,In_279);
and U515 (N_515,In_263,In_68);
and U516 (N_516,In_141,In_473);
nand U517 (N_517,In_419,In_377);
and U518 (N_518,In_695,In_423);
and U519 (N_519,In_42,In_138);
nor U520 (N_520,In_154,In_621);
or U521 (N_521,In_629,In_687);
nor U522 (N_522,In_24,In_390);
or U523 (N_523,In_467,In_425);
nand U524 (N_524,In_447,In_264);
or U525 (N_525,In_321,In_368);
nor U526 (N_526,In_552,In_677);
or U527 (N_527,In_68,In_229);
and U528 (N_528,In_59,In_110);
nand U529 (N_529,In_404,In_143);
and U530 (N_530,In_459,In_33);
or U531 (N_531,In_455,In_633);
and U532 (N_532,In_133,In_639);
or U533 (N_533,In_117,In_481);
and U534 (N_534,In_749,In_524);
and U535 (N_535,In_83,In_36);
nand U536 (N_536,In_80,In_451);
nand U537 (N_537,In_43,In_552);
or U538 (N_538,In_340,In_100);
nor U539 (N_539,In_699,In_495);
nand U540 (N_540,In_398,In_424);
nand U541 (N_541,In_327,In_60);
and U542 (N_542,In_424,In_568);
or U543 (N_543,In_223,In_616);
nand U544 (N_544,In_60,In_102);
nand U545 (N_545,In_709,In_608);
or U546 (N_546,In_669,In_241);
nor U547 (N_547,In_550,In_195);
nand U548 (N_548,In_149,In_620);
nand U549 (N_549,In_33,In_305);
nand U550 (N_550,In_6,In_644);
or U551 (N_551,In_499,In_707);
or U552 (N_552,In_574,In_739);
nand U553 (N_553,In_57,In_140);
nor U554 (N_554,In_443,In_563);
xnor U555 (N_555,In_584,In_680);
nand U556 (N_556,In_45,In_40);
nor U557 (N_557,In_112,In_400);
and U558 (N_558,In_250,In_391);
and U559 (N_559,In_729,In_107);
and U560 (N_560,In_697,In_280);
nor U561 (N_561,In_261,In_318);
or U562 (N_562,In_247,In_256);
and U563 (N_563,In_182,In_102);
nand U564 (N_564,In_238,In_417);
and U565 (N_565,In_678,In_326);
nand U566 (N_566,In_219,In_210);
nor U567 (N_567,In_747,In_600);
nand U568 (N_568,In_436,In_572);
and U569 (N_569,In_60,In_454);
or U570 (N_570,In_136,In_272);
nor U571 (N_571,In_26,In_33);
nor U572 (N_572,In_524,In_460);
and U573 (N_573,In_226,In_96);
nor U574 (N_574,In_235,In_733);
nand U575 (N_575,In_261,In_731);
or U576 (N_576,In_381,In_345);
and U577 (N_577,In_540,In_535);
nand U578 (N_578,In_41,In_80);
nor U579 (N_579,In_484,In_59);
nand U580 (N_580,In_240,In_665);
nor U581 (N_581,In_582,In_414);
nand U582 (N_582,In_631,In_21);
and U583 (N_583,In_90,In_61);
nand U584 (N_584,In_331,In_70);
nand U585 (N_585,In_156,In_95);
and U586 (N_586,In_403,In_21);
nor U587 (N_587,In_61,In_660);
or U588 (N_588,In_708,In_392);
xnor U589 (N_589,In_161,In_250);
and U590 (N_590,In_622,In_411);
or U591 (N_591,In_65,In_139);
nand U592 (N_592,In_117,In_87);
and U593 (N_593,In_53,In_163);
nor U594 (N_594,In_602,In_159);
and U595 (N_595,In_615,In_461);
nand U596 (N_596,In_356,In_241);
nor U597 (N_597,In_401,In_124);
nor U598 (N_598,In_406,In_531);
or U599 (N_599,In_218,In_575);
nand U600 (N_600,In_125,In_463);
nor U601 (N_601,In_410,In_705);
or U602 (N_602,In_20,In_144);
and U603 (N_603,In_690,In_189);
nand U604 (N_604,In_542,In_697);
nand U605 (N_605,In_217,In_205);
and U606 (N_606,In_97,In_616);
or U607 (N_607,In_10,In_344);
and U608 (N_608,In_44,In_29);
nor U609 (N_609,In_510,In_135);
and U610 (N_610,In_579,In_615);
or U611 (N_611,In_545,In_512);
nand U612 (N_612,In_588,In_125);
xor U613 (N_613,In_606,In_526);
and U614 (N_614,In_740,In_612);
and U615 (N_615,In_387,In_456);
or U616 (N_616,In_574,In_493);
nand U617 (N_617,In_60,In_441);
and U618 (N_618,In_231,In_620);
xnor U619 (N_619,In_577,In_713);
and U620 (N_620,In_191,In_86);
or U621 (N_621,In_619,In_520);
nand U622 (N_622,In_403,In_730);
and U623 (N_623,In_238,In_517);
and U624 (N_624,In_396,In_659);
xor U625 (N_625,In_2,In_131);
xor U626 (N_626,In_564,In_584);
nor U627 (N_627,In_237,In_32);
nand U628 (N_628,In_236,In_419);
nand U629 (N_629,In_165,In_355);
nand U630 (N_630,In_69,In_196);
and U631 (N_631,In_492,In_410);
nand U632 (N_632,In_8,In_94);
and U633 (N_633,In_265,In_595);
nand U634 (N_634,In_83,In_149);
nand U635 (N_635,In_648,In_275);
or U636 (N_636,In_9,In_509);
nor U637 (N_637,In_714,In_105);
or U638 (N_638,In_109,In_565);
nor U639 (N_639,In_13,In_230);
or U640 (N_640,In_676,In_385);
nor U641 (N_641,In_727,In_223);
or U642 (N_642,In_404,In_341);
or U643 (N_643,In_59,In_415);
nor U644 (N_644,In_197,In_208);
or U645 (N_645,In_563,In_57);
and U646 (N_646,In_42,In_674);
and U647 (N_647,In_353,In_517);
and U648 (N_648,In_67,In_164);
and U649 (N_649,In_529,In_576);
nor U650 (N_650,In_57,In_533);
and U651 (N_651,In_326,In_229);
or U652 (N_652,In_730,In_89);
nand U653 (N_653,In_264,In_723);
and U654 (N_654,In_304,In_409);
nor U655 (N_655,In_266,In_355);
xor U656 (N_656,In_14,In_64);
nor U657 (N_657,In_102,In_482);
or U658 (N_658,In_397,In_662);
or U659 (N_659,In_445,In_350);
or U660 (N_660,In_370,In_103);
nor U661 (N_661,In_401,In_376);
nor U662 (N_662,In_63,In_718);
nor U663 (N_663,In_412,In_335);
or U664 (N_664,In_407,In_144);
nand U665 (N_665,In_535,In_442);
nor U666 (N_666,In_450,In_60);
nor U667 (N_667,In_290,In_479);
nand U668 (N_668,In_407,In_161);
or U669 (N_669,In_588,In_624);
and U670 (N_670,In_457,In_628);
nor U671 (N_671,In_420,In_193);
and U672 (N_672,In_82,In_27);
nor U673 (N_673,In_512,In_253);
nand U674 (N_674,In_219,In_215);
or U675 (N_675,In_520,In_505);
xor U676 (N_676,In_67,In_711);
nor U677 (N_677,In_735,In_217);
or U678 (N_678,In_485,In_729);
and U679 (N_679,In_429,In_496);
nand U680 (N_680,In_324,In_128);
nor U681 (N_681,In_686,In_698);
nor U682 (N_682,In_656,In_482);
nor U683 (N_683,In_229,In_435);
nor U684 (N_684,In_39,In_423);
nand U685 (N_685,In_506,In_712);
nor U686 (N_686,In_636,In_13);
and U687 (N_687,In_60,In_37);
nand U688 (N_688,In_248,In_197);
or U689 (N_689,In_285,In_122);
and U690 (N_690,In_421,In_683);
nand U691 (N_691,In_469,In_302);
nand U692 (N_692,In_379,In_407);
and U693 (N_693,In_740,In_618);
nand U694 (N_694,In_63,In_501);
and U695 (N_695,In_198,In_341);
nor U696 (N_696,In_77,In_728);
or U697 (N_697,In_8,In_226);
nand U698 (N_698,In_358,In_123);
nand U699 (N_699,In_709,In_275);
nor U700 (N_700,In_559,In_328);
nor U701 (N_701,In_181,In_550);
or U702 (N_702,In_741,In_295);
nor U703 (N_703,In_337,In_708);
or U704 (N_704,In_479,In_80);
nand U705 (N_705,In_527,In_565);
nor U706 (N_706,In_660,In_15);
nor U707 (N_707,In_584,In_175);
and U708 (N_708,In_496,In_519);
or U709 (N_709,In_497,In_347);
and U710 (N_710,In_167,In_124);
and U711 (N_711,In_562,In_238);
nor U712 (N_712,In_334,In_51);
nor U713 (N_713,In_183,In_643);
nand U714 (N_714,In_55,In_142);
nand U715 (N_715,In_87,In_157);
or U716 (N_716,In_326,In_716);
or U717 (N_717,In_401,In_226);
nor U718 (N_718,In_664,In_350);
nor U719 (N_719,In_535,In_537);
nor U720 (N_720,In_378,In_97);
or U721 (N_721,In_719,In_738);
nor U722 (N_722,In_258,In_311);
nand U723 (N_723,In_160,In_335);
and U724 (N_724,In_642,In_560);
nor U725 (N_725,In_726,In_107);
nand U726 (N_726,In_703,In_144);
or U727 (N_727,In_420,In_356);
nor U728 (N_728,In_146,In_32);
and U729 (N_729,In_273,In_620);
nor U730 (N_730,In_559,In_55);
and U731 (N_731,In_194,In_641);
nor U732 (N_732,In_198,In_542);
nand U733 (N_733,In_436,In_237);
or U734 (N_734,In_412,In_39);
and U735 (N_735,In_700,In_576);
nor U736 (N_736,In_195,In_547);
nand U737 (N_737,In_221,In_438);
or U738 (N_738,In_63,In_42);
and U739 (N_739,In_272,In_519);
nand U740 (N_740,In_666,In_557);
nand U741 (N_741,In_278,In_508);
nor U742 (N_742,In_165,In_354);
nor U743 (N_743,In_438,In_135);
nor U744 (N_744,In_362,In_407);
nand U745 (N_745,In_49,In_548);
nor U746 (N_746,In_135,In_468);
and U747 (N_747,In_202,In_44);
nor U748 (N_748,In_566,In_461);
or U749 (N_749,In_640,In_421);
or U750 (N_750,In_675,In_490);
or U751 (N_751,In_408,In_122);
and U752 (N_752,In_726,In_169);
or U753 (N_753,In_541,In_411);
and U754 (N_754,In_63,In_18);
nor U755 (N_755,In_366,In_269);
or U756 (N_756,In_367,In_514);
and U757 (N_757,In_452,In_510);
nand U758 (N_758,In_540,In_638);
nand U759 (N_759,In_418,In_355);
and U760 (N_760,In_144,In_489);
or U761 (N_761,In_346,In_539);
nor U762 (N_762,In_139,In_91);
and U763 (N_763,In_663,In_405);
and U764 (N_764,In_680,In_602);
nor U765 (N_765,In_733,In_420);
or U766 (N_766,In_20,In_112);
or U767 (N_767,In_605,In_571);
and U768 (N_768,In_699,In_485);
or U769 (N_769,In_380,In_338);
xor U770 (N_770,In_570,In_269);
and U771 (N_771,In_5,In_127);
and U772 (N_772,In_412,In_109);
or U773 (N_773,In_538,In_141);
or U774 (N_774,In_716,In_435);
nor U775 (N_775,In_346,In_265);
nor U776 (N_776,In_112,In_5);
nand U777 (N_777,In_200,In_133);
and U778 (N_778,In_540,In_138);
nor U779 (N_779,In_700,In_607);
or U780 (N_780,In_660,In_379);
nand U781 (N_781,In_648,In_281);
or U782 (N_782,In_89,In_682);
or U783 (N_783,In_477,In_136);
nor U784 (N_784,In_84,In_639);
or U785 (N_785,In_312,In_749);
or U786 (N_786,In_450,In_373);
nand U787 (N_787,In_88,In_530);
nand U788 (N_788,In_724,In_693);
nand U789 (N_789,In_102,In_703);
and U790 (N_790,In_478,In_222);
or U791 (N_791,In_442,In_427);
and U792 (N_792,In_261,In_395);
nand U793 (N_793,In_673,In_684);
nor U794 (N_794,In_370,In_547);
nor U795 (N_795,In_221,In_621);
and U796 (N_796,In_109,In_527);
and U797 (N_797,In_160,In_103);
nand U798 (N_798,In_648,In_725);
or U799 (N_799,In_93,In_733);
or U800 (N_800,In_338,In_625);
or U801 (N_801,In_611,In_304);
nor U802 (N_802,In_185,In_724);
nand U803 (N_803,In_259,In_633);
nor U804 (N_804,In_429,In_68);
nand U805 (N_805,In_671,In_491);
nor U806 (N_806,In_167,In_718);
nor U807 (N_807,In_287,In_335);
or U808 (N_808,In_497,In_191);
or U809 (N_809,In_108,In_166);
nand U810 (N_810,In_560,In_156);
nand U811 (N_811,In_390,In_355);
and U812 (N_812,In_269,In_185);
nor U813 (N_813,In_281,In_743);
or U814 (N_814,In_382,In_399);
nor U815 (N_815,In_222,In_6);
nor U816 (N_816,In_26,In_634);
nor U817 (N_817,In_154,In_200);
xor U818 (N_818,In_553,In_211);
nor U819 (N_819,In_451,In_37);
or U820 (N_820,In_603,In_585);
or U821 (N_821,In_162,In_369);
and U822 (N_822,In_533,In_29);
nand U823 (N_823,In_126,In_517);
xor U824 (N_824,In_255,In_428);
and U825 (N_825,In_166,In_170);
nand U826 (N_826,In_520,In_647);
or U827 (N_827,In_682,In_551);
nor U828 (N_828,In_41,In_575);
nor U829 (N_829,In_112,In_34);
and U830 (N_830,In_582,In_111);
and U831 (N_831,In_588,In_493);
or U832 (N_832,In_188,In_542);
nor U833 (N_833,In_394,In_420);
nor U834 (N_834,In_543,In_50);
nor U835 (N_835,In_390,In_240);
nand U836 (N_836,In_176,In_135);
nor U837 (N_837,In_613,In_34);
nor U838 (N_838,In_389,In_281);
and U839 (N_839,In_263,In_648);
nor U840 (N_840,In_459,In_151);
or U841 (N_841,In_294,In_228);
or U842 (N_842,In_238,In_133);
and U843 (N_843,In_629,In_220);
nand U844 (N_844,In_475,In_550);
or U845 (N_845,In_383,In_18);
nand U846 (N_846,In_152,In_91);
xor U847 (N_847,In_308,In_286);
or U848 (N_848,In_432,In_632);
and U849 (N_849,In_355,In_386);
nor U850 (N_850,In_299,In_72);
nand U851 (N_851,In_400,In_450);
or U852 (N_852,In_232,In_247);
and U853 (N_853,In_701,In_629);
nor U854 (N_854,In_78,In_538);
nor U855 (N_855,In_256,In_407);
nand U856 (N_856,In_525,In_434);
and U857 (N_857,In_397,In_9);
nand U858 (N_858,In_9,In_355);
nand U859 (N_859,In_479,In_349);
nor U860 (N_860,In_420,In_376);
and U861 (N_861,In_551,In_29);
or U862 (N_862,In_193,In_24);
nand U863 (N_863,In_275,In_337);
or U864 (N_864,In_645,In_144);
nor U865 (N_865,In_219,In_123);
or U866 (N_866,In_729,In_571);
and U867 (N_867,In_256,In_588);
nand U868 (N_868,In_288,In_509);
xor U869 (N_869,In_133,In_727);
nand U870 (N_870,In_493,In_351);
nor U871 (N_871,In_260,In_525);
nor U872 (N_872,In_673,In_348);
and U873 (N_873,In_214,In_606);
nand U874 (N_874,In_250,In_343);
nand U875 (N_875,In_275,In_176);
and U876 (N_876,In_245,In_34);
and U877 (N_877,In_354,In_491);
or U878 (N_878,In_409,In_309);
and U879 (N_879,In_74,In_220);
and U880 (N_880,In_45,In_117);
nand U881 (N_881,In_555,In_290);
nor U882 (N_882,In_149,In_176);
or U883 (N_883,In_746,In_316);
and U884 (N_884,In_164,In_710);
nand U885 (N_885,In_640,In_690);
or U886 (N_886,In_619,In_438);
nand U887 (N_887,In_525,In_696);
nand U888 (N_888,In_522,In_153);
nand U889 (N_889,In_448,In_250);
or U890 (N_890,In_56,In_558);
and U891 (N_891,In_47,In_414);
or U892 (N_892,In_123,In_223);
and U893 (N_893,In_545,In_357);
and U894 (N_894,In_8,In_592);
nand U895 (N_895,In_401,In_586);
or U896 (N_896,In_104,In_663);
nand U897 (N_897,In_226,In_253);
nor U898 (N_898,In_213,In_11);
or U899 (N_899,In_601,In_457);
and U900 (N_900,In_322,In_403);
nand U901 (N_901,In_119,In_184);
nor U902 (N_902,In_547,In_82);
nand U903 (N_903,In_133,In_129);
or U904 (N_904,In_659,In_366);
xor U905 (N_905,In_465,In_490);
and U906 (N_906,In_480,In_33);
xnor U907 (N_907,In_68,In_2);
nand U908 (N_908,In_557,In_156);
and U909 (N_909,In_118,In_471);
nand U910 (N_910,In_588,In_146);
and U911 (N_911,In_616,In_123);
or U912 (N_912,In_713,In_641);
nand U913 (N_913,In_585,In_402);
xor U914 (N_914,In_46,In_260);
or U915 (N_915,In_384,In_572);
xnor U916 (N_916,In_435,In_349);
or U917 (N_917,In_234,In_342);
and U918 (N_918,In_222,In_616);
nand U919 (N_919,In_282,In_642);
nor U920 (N_920,In_308,In_176);
xnor U921 (N_921,In_572,In_338);
nand U922 (N_922,In_81,In_421);
nand U923 (N_923,In_224,In_188);
or U924 (N_924,In_284,In_166);
and U925 (N_925,In_708,In_250);
xor U926 (N_926,In_668,In_463);
or U927 (N_927,In_583,In_634);
or U928 (N_928,In_28,In_196);
nand U929 (N_929,In_401,In_659);
nand U930 (N_930,In_153,In_345);
or U931 (N_931,In_331,In_52);
nand U932 (N_932,In_442,In_474);
or U933 (N_933,In_439,In_213);
and U934 (N_934,In_560,In_378);
nand U935 (N_935,In_241,In_193);
and U936 (N_936,In_100,In_111);
and U937 (N_937,In_598,In_703);
or U938 (N_938,In_560,In_537);
and U939 (N_939,In_19,In_377);
nand U940 (N_940,In_736,In_699);
nor U941 (N_941,In_343,In_148);
nand U942 (N_942,In_326,In_711);
nand U943 (N_943,In_367,In_455);
or U944 (N_944,In_587,In_203);
and U945 (N_945,In_438,In_720);
and U946 (N_946,In_81,In_392);
or U947 (N_947,In_588,In_434);
and U948 (N_948,In_308,In_191);
nor U949 (N_949,In_375,In_262);
nand U950 (N_950,In_472,In_388);
or U951 (N_951,In_510,In_676);
nor U952 (N_952,In_587,In_622);
nor U953 (N_953,In_38,In_359);
or U954 (N_954,In_702,In_431);
nand U955 (N_955,In_45,In_229);
and U956 (N_956,In_231,In_481);
nor U957 (N_957,In_401,In_696);
nand U958 (N_958,In_732,In_614);
and U959 (N_959,In_479,In_382);
or U960 (N_960,In_347,In_572);
nor U961 (N_961,In_142,In_743);
or U962 (N_962,In_673,In_310);
or U963 (N_963,In_339,In_315);
nor U964 (N_964,In_463,In_48);
nand U965 (N_965,In_15,In_702);
and U966 (N_966,In_611,In_513);
nor U967 (N_967,In_266,In_124);
or U968 (N_968,In_631,In_371);
or U969 (N_969,In_455,In_238);
and U970 (N_970,In_316,In_138);
xor U971 (N_971,In_441,In_578);
nor U972 (N_972,In_695,In_334);
and U973 (N_973,In_31,In_258);
nand U974 (N_974,In_690,In_61);
and U975 (N_975,In_621,In_186);
nand U976 (N_976,In_52,In_603);
and U977 (N_977,In_676,In_246);
nand U978 (N_978,In_30,In_25);
xor U979 (N_979,In_718,In_738);
or U980 (N_980,In_10,In_378);
or U981 (N_981,In_532,In_58);
and U982 (N_982,In_601,In_416);
or U983 (N_983,In_62,In_476);
xor U984 (N_984,In_61,In_367);
and U985 (N_985,In_100,In_427);
or U986 (N_986,In_545,In_252);
and U987 (N_987,In_377,In_187);
or U988 (N_988,In_337,In_87);
nand U989 (N_989,In_398,In_625);
nand U990 (N_990,In_538,In_601);
or U991 (N_991,In_408,In_536);
nand U992 (N_992,In_141,In_714);
nand U993 (N_993,In_509,In_423);
nor U994 (N_994,In_674,In_298);
nor U995 (N_995,In_228,In_100);
and U996 (N_996,In_557,In_486);
nor U997 (N_997,In_139,In_297);
and U998 (N_998,In_587,In_344);
nor U999 (N_999,In_693,In_199);
nand U1000 (N_1000,In_6,In_312);
or U1001 (N_1001,In_506,In_438);
and U1002 (N_1002,In_525,In_517);
nand U1003 (N_1003,In_82,In_318);
and U1004 (N_1004,In_420,In_141);
or U1005 (N_1005,In_9,In_514);
nor U1006 (N_1006,In_15,In_85);
and U1007 (N_1007,In_93,In_399);
or U1008 (N_1008,In_366,In_705);
and U1009 (N_1009,In_260,In_654);
nand U1010 (N_1010,In_7,In_453);
or U1011 (N_1011,In_500,In_301);
nand U1012 (N_1012,In_336,In_342);
nor U1013 (N_1013,In_554,In_54);
or U1014 (N_1014,In_207,In_636);
nand U1015 (N_1015,In_532,In_641);
and U1016 (N_1016,In_743,In_299);
xor U1017 (N_1017,In_692,In_139);
or U1018 (N_1018,In_159,In_119);
nand U1019 (N_1019,In_426,In_465);
or U1020 (N_1020,In_211,In_508);
and U1021 (N_1021,In_198,In_409);
nand U1022 (N_1022,In_390,In_40);
nand U1023 (N_1023,In_261,In_388);
nor U1024 (N_1024,In_173,In_275);
and U1025 (N_1025,In_142,In_548);
or U1026 (N_1026,In_23,In_688);
nand U1027 (N_1027,In_498,In_84);
nor U1028 (N_1028,In_648,In_103);
nor U1029 (N_1029,In_492,In_173);
and U1030 (N_1030,In_193,In_190);
nor U1031 (N_1031,In_500,In_306);
and U1032 (N_1032,In_349,In_555);
and U1033 (N_1033,In_666,In_400);
nand U1034 (N_1034,In_657,In_705);
or U1035 (N_1035,In_432,In_643);
xnor U1036 (N_1036,In_96,In_721);
or U1037 (N_1037,In_464,In_100);
nand U1038 (N_1038,In_201,In_748);
and U1039 (N_1039,In_479,In_159);
nand U1040 (N_1040,In_426,In_573);
and U1041 (N_1041,In_112,In_557);
nand U1042 (N_1042,In_636,In_410);
and U1043 (N_1043,In_345,In_291);
nor U1044 (N_1044,In_472,In_463);
or U1045 (N_1045,In_711,In_701);
nor U1046 (N_1046,In_45,In_527);
and U1047 (N_1047,In_272,In_95);
nor U1048 (N_1048,In_1,In_476);
nand U1049 (N_1049,In_447,In_496);
nor U1050 (N_1050,In_646,In_512);
and U1051 (N_1051,In_168,In_63);
or U1052 (N_1052,In_231,In_330);
nand U1053 (N_1053,In_402,In_9);
or U1054 (N_1054,In_306,In_26);
nand U1055 (N_1055,In_9,In_699);
nand U1056 (N_1056,In_624,In_332);
nor U1057 (N_1057,In_221,In_193);
and U1058 (N_1058,In_61,In_616);
and U1059 (N_1059,In_520,In_221);
nor U1060 (N_1060,In_499,In_590);
or U1061 (N_1061,In_501,In_338);
nor U1062 (N_1062,In_19,In_401);
nor U1063 (N_1063,In_527,In_68);
or U1064 (N_1064,In_446,In_411);
nand U1065 (N_1065,In_424,In_645);
nand U1066 (N_1066,In_50,In_388);
nor U1067 (N_1067,In_441,In_296);
and U1068 (N_1068,In_301,In_677);
nand U1069 (N_1069,In_59,In_735);
nand U1070 (N_1070,In_535,In_431);
or U1071 (N_1071,In_495,In_511);
nor U1072 (N_1072,In_375,In_286);
nand U1073 (N_1073,In_108,In_691);
and U1074 (N_1074,In_188,In_92);
nand U1075 (N_1075,In_81,In_466);
nor U1076 (N_1076,In_142,In_295);
nand U1077 (N_1077,In_621,In_23);
xor U1078 (N_1078,In_353,In_406);
nor U1079 (N_1079,In_648,In_118);
and U1080 (N_1080,In_147,In_266);
nor U1081 (N_1081,In_124,In_313);
and U1082 (N_1082,In_704,In_207);
nand U1083 (N_1083,In_339,In_327);
or U1084 (N_1084,In_114,In_574);
and U1085 (N_1085,In_382,In_279);
nand U1086 (N_1086,In_472,In_196);
nand U1087 (N_1087,In_211,In_144);
nand U1088 (N_1088,In_298,In_447);
or U1089 (N_1089,In_71,In_220);
nor U1090 (N_1090,In_237,In_541);
nor U1091 (N_1091,In_624,In_67);
nand U1092 (N_1092,In_683,In_95);
nor U1093 (N_1093,In_656,In_133);
and U1094 (N_1094,In_91,In_433);
nand U1095 (N_1095,In_518,In_451);
nor U1096 (N_1096,In_195,In_404);
nor U1097 (N_1097,In_48,In_669);
and U1098 (N_1098,In_702,In_185);
and U1099 (N_1099,In_32,In_651);
nand U1100 (N_1100,In_589,In_0);
or U1101 (N_1101,In_573,In_581);
nand U1102 (N_1102,In_188,In_250);
nor U1103 (N_1103,In_328,In_545);
nand U1104 (N_1104,In_113,In_185);
and U1105 (N_1105,In_501,In_142);
nor U1106 (N_1106,In_89,In_235);
and U1107 (N_1107,In_244,In_265);
nand U1108 (N_1108,In_209,In_431);
and U1109 (N_1109,In_221,In_466);
or U1110 (N_1110,In_59,In_124);
nand U1111 (N_1111,In_305,In_497);
nand U1112 (N_1112,In_325,In_311);
and U1113 (N_1113,In_110,In_97);
nor U1114 (N_1114,In_87,In_487);
and U1115 (N_1115,In_708,In_132);
xor U1116 (N_1116,In_364,In_262);
nand U1117 (N_1117,In_347,In_65);
nand U1118 (N_1118,In_649,In_600);
and U1119 (N_1119,In_129,In_539);
nand U1120 (N_1120,In_159,In_664);
or U1121 (N_1121,In_68,In_504);
and U1122 (N_1122,In_292,In_10);
nor U1123 (N_1123,In_644,In_620);
nor U1124 (N_1124,In_94,In_218);
and U1125 (N_1125,In_312,In_338);
xnor U1126 (N_1126,In_130,In_377);
and U1127 (N_1127,In_91,In_30);
and U1128 (N_1128,In_669,In_692);
or U1129 (N_1129,In_177,In_655);
nand U1130 (N_1130,In_715,In_125);
and U1131 (N_1131,In_56,In_147);
or U1132 (N_1132,In_143,In_110);
and U1133 (N_1133,In_417,In_55);
and U1134 (N_1134,In_567,In_59);
or U1135 (N_1135,In_303,In_252);
nand U1136 (N_1136,In_163,In_76);
nor U1137 (N_1137,In_433,In_669);
and U1138 (N_1138,In_696,In_701);
and U1139 (N_1139,In_416,In_106);
and U1140 (N_1140,In_236,In_695);
or U1141 (N_1141,In_460,In_552);
or U1142 (N_1142,In_91,In_221);
nor U1143 (N_1143,In_233,In_238);
nand U1144 (N_1144,In_476,In_360);
nand U1145 (N_1145,In_53,In_120);
nand U1146 (N_1146,In_444,In_536);
or U1147 (N_1147,In_163,In_466);
and U1148 (N_1148,In_365,In_673);
nor U1149 (N_1149,In_596,In_275);
nor U1150 (N_1150,In_555,In_130);
or U1151 (N_1151,In_393,In_747);
or U1152 (N_1152,In_494,In_498);
or U1153 (N_1153,In_566,In_450);
nand U1154 (N_1154,In_500,In_699);
and U1155 (N_1155,In_220,In_474);
or U1156 (N_1156,In_667,In_574);
or U1157 (N_1157,In_679,In_314);
nand U1158 (N_1158,In_470,In_702);
nor U1159 (N_1159,In_336,In_474);
nand U1160 (N_1160,In_587,In_268);
or U1161 (N_1161,In_262,In_326);
or U1162 (N_1162,In_545,In_355);
or U1163 (N_1163,In_643,In_443);
and U1164 (N_1164,In_142,In_728);
or U1165 (N_1165,In_79,In_538);
nor U1166 (N_1166,In_262,In_321);
nand U1167 (N_1167,In_379,In_214);
or U1168 (N_1168,In_738,In_632);
and U1169 (N_1169,In_715,In_237);
and U1170 (N_1170,In_44,In_437);
nor U1171 (N_1171,In_382,In_260);
or U1172 (N_1172,In_536,In_277);
nand U1173 (N_1173,In_170,In_77);
nor U1174 (N_1174,In_379,In_397);
and U1175 (N_1175,In_201,In_337);
or U1176 (N_1176,In_6,In_424);
nand U1177 (N_1177,In_259,In_679);
nor U1178 (N_1178,In_679,In_691);
nor U1179 (N_1179,In_345,In_8);
or U1180 (N_1180,In_348,In_392);
nor U1181 (N_1181,In_292,In_168);
nand U1182 (N_1182,In_652,In_19);
and U1183 (N_1183,In_543,In_456);
and U1184 (N_1184,In_713,In_227);
and U1185 (N_1185,In_67,In_176);
nand U1186 (N_1186,In_197,In_393);
xnor U1187 (N_1187,In_595,In_421);
nor U1188 (N_1188,In_483,In_127);
nand U1189 (N_1189,In_31,In_622);
nand U1190 (N_1190,In_629,In_228);
nor U1191 (N_1191,In_171,In_347);
nor U1192 (N_1192,In_701,In_594);
or U1193 (N_1193,In_314,In_254);
nand U1194 (N_1194,In_148,In_272);
nor U1195 (N_1195,In_528,In_183);
nand U1196 (N_1196,In_463,In_693);
and U1197 (N_1197,In_337,In_493);
nand U1198 (N_1198,In_567,In_161);
nor U1199 (N_1199,In_575,In_579);
or U1200 (N_1200,In_26,In_171);
nand U1201 (N_1201,In_275,In_126);
nor U1202 (N_1202,In_170,In_50);
or U1203 (N_1203,In_614,In_689);
xor U1204 (N_1204,In_211,In_493);
nor U1205 (N_1205,In_102,In_286);
or U1206 (N_1206,In_82,In_300);
nor U1207 (N_1207,In_256,In_742);
nor U1208 (N_1208,In_176,In_559);
nor U1209 (N_1209,In_565,In_163);
or U1210 (N_1210,In_387,In_537);
nand U1211 (N_1211,In_507,In_361);
and U1212 (N_1212,In_438,In_397);
and U1213 (N_1213,In_46,In_254);
or U1214 (N_1214,In_746,In_687);
or U1215 (N_1215,In_509,In_167);
nor U1216 (N_1216,In_557,In_565);
nor U1217 (N_1217,In_740,In_714);
nor U1218 (N_1218,In_125,In_652);
nand U1219 (N_1219,In_94,In_451);
and U1220 (N_1220,In_461,In_399);
or U1221 (N_1221,In_654,In_495);
nor U1222 (N_1222,In_540,In_46);
nor U1223 (N_1223,In_521,In_686);
or U1224 (N_1224,In_210,In_643);
or U1225 (N_1225,In_498,In_61);
or U1226 (N_1226,In_373,In_437);
and U1227 (N_1227,In_518,In_612);
nand U1228 (N_1228,In_732,In_339);
nand U1229 (N_1229,In_225,In_254);
and U1230 (N_1230,In_226,In_436);
nor U1231 (N_1231,In_527,In_657);
nand U1232 (N_1232,In_90,In_200);
nor U1233 (N_1233,In_461,In_361);
nor U1234 (N_1234,In_497,In_491);
nand U1235 (N_1235,In_127,In_681);
nand U1236 (N_1236,In_42,In_201);
nand U1237 (N_1237,In_132,In_312);
nor U1238 (N_1238,In_482,In_446);
or U1239 (N_1239,In_393,In_89);
nor U1240 (N_1240,In_604,In_699);
nand U1241 (N_1241,In_445,In_134);
or U1242 (N_1242,In_633,In_160);
nand U1243 (N_1243,In_7,In_276);
nand U1244 (N_1244,In_743,In_675);
and U1245 (N_1245,In_19,In_116);
nand U1246 (N_1246,In_480,In_225);
xnor U1247 (N_1247,In_554,In_686);
nor U1248 (N_1248,In_744,In_232);
nor U1249 (N_1249,In_79,In_641);
or U1250 (N_1250,In_212,In_134);
or U1251 (N_1251,In_14,In_53);
and U1252 (N_1252,In_197,In_134);
and U1253 (N_1253,In_171,In_41);
or U1254 (N_1254,In_388,In_330);
or U1255 (N_1255,In_381,In_88);
or U1256 (N_1256,In_376,In_460);
and U1257 (N_1257,In_310,In_98);
nor U1258 (N_1258,In_594,In_50);
nand U1259 (N_1259,In_12,In_199);
nand U1260 (N_1260,In_603,In_11);
nor U1261 (N_1261,In_379,In_648);
and U1262 (N_1262,In_557,In_131);
and U1263 (N_1263,In_651,In_50);
nor U1264 (N_1264,In_694,In_89);
and U1265 (N_1265,In_104,In_5);
and U1266 (N_1266,In_17,In_122);
nor U1267 (N_1267,In_641,In_592);
and U1268 (N_1268,In_289,In_569);
nor U1269 (N_1269,In_730,In_718);
xnor U1270 (N_1270,In_75,In_516);
or U1271 (N_1271,In_122,In_535);
nand U1272 (N_1272,In_368,In_375);
or U1273 (N_1273,In_679,In_121);
and U1274 (N_1274,In_654,In_345);
nor U1275 (N_1275,In_620,In_696);
nand U1276 (N_1276,In_598,In_655);
nand U1277 (N_1277,In_645,In_17);
nand U1278 (N_1278,In_350,In_735);
nand U1279 (N_1279,In_364,In_491);
and U1280 (N_1280,In_391,In_492);
xor U1281 (N_1281,In_458,In_326);
and U1282 (N_1282,In_34,In_188);
and U1283 (N_1283,In_243,In_135);
nor U1284 (N_1284,In_442,In_131);
nand U1285 (N_1285,In_474,In_322);
nand U1286 (N_1286,In_448,In_74);
and U1287 (N_1287,In_150,In_447);
nor U1288 (N_1288,In_633,In_184);
or U1289 (N_1289,In_104,In_375);
nor U1290 (N_1290,In_728,In_712);
nand U1291 (N_1291,In_21,In_67);
nor U1292 (N_1292,In_12,In_709);
or U1293 (N_1293,In_148,In_13);
or U1294 (N_1294,In_711,In_278);
nor U1295 (N_1295,In_639,In_309);
nor U1296 (N_1296,In_706,In_432);
and U1297 (N_1297,In_572,In_178);
and U1298 (N_1298,In_353,In_139);
nand U1299 (N_1299,In_50,In_4);
and U1300 (N_1300,In_745,In_99);
xor U1301 (N_1301,In_559,In_253);
xnor U1302 (N_1302,In_66,In_99);
nor U1303 (N_1303,In_474,In_617);
and U1304 (N_1304,In_553,In_189);
and U1305 (N_1305,In_710,In_518);
nor U1306 (N_1306,In_639,In_303);
or U1307 (N_1307,In_586,In_185);
or U1308 (N_1308,In_259,In_422);
nor U1309 (N_1309,In_519,In_526);
nor U1310 (N_1310,In_585,In_184);
or U1311 (N_1311,In_226,In_473);
and U1312 (N_1312,In_418,In_687);
nor U1313 (N_1313,In_295,In_215);
and U1314 (N_1314,In_186,In_748);
nor U1315 (N_1315,In_89,In_161);
nand U1316 (N_1316,In_167,In_75);
or U1317 (N_1317,In_705,In_21);
nand U1318 (N_1318,In_90,In_530);
and U1319 (N_1319,In_668,In_680);
and U1320 (N_1320,In_200,In_408);
nor U1321 (N_1321,In_725,In_89);
nand U1322 (N_1322,In_195,In_109);
nor U1323 (N_1323,In_528,In_220);
or U1324 (N_1324,In_703,In_94);
nand U1325 (N_1325,In_386,In_298);
xor U1326 (N_1326,In_342,In_389);
nor U1327 (N_1327,In_485,In_602);
nand U1328 (N_1328,In_704,In_330);
nand U1329 (N_1329,In_405,In_409);
nand U1330 (N_1330,In_634,In_202);
nand U1331 (N_1331,In_298,In_515);
or U1332 (N_1332,In_24,In_486);
nor U1333 (N_1333,In_112,In_78);
and U1334 (N_1334,In_505,In_283);
nand U1335 (N_1335,In_395,In_162);
nor U1336 (N_1336,In_308,In_67);
nor U1337 (N_1337,In_298,In_432);
and U1338 (N_1338,In_294,In_732);
nor U1339 (N_1339,In_386,In_540);
or U1340 (N_1340,In_745,In_388);
or U1341 (N_1341,In_413,In_387);
nand U1342 (N_1342,In_589,In_67);
or U1343 (N_1343,In_450,In_573);
nand U1344 (N_1344,In_565,In_269);
nor U1345 (N_1345,In_128,In_28);
and U1346 (N_1346,In_696,In_527);
or U1347 (N_1347,In_500,In_734);
nand U1348 (N_1348,In_459,In_510);
nand U1349 (N_1349,In_153,In_717);
nor U1350 (N_1350,In_702,In_531);
or U1351 (N_1351,In_603,In_101);
and U1352 (N_1352,In_21,In_596);
nor U1353 (N_1353,In_142,In_694);
nor U1354 (N_1354,In_404,In_446);
nand U1355 (N_1355,In_470,In_289);
nor U1356 (N_1356,In_164,In_511);
and U1357 (N_1357,In_179,In_122);
nor U1358 (N_1358,In_79,In_586);
nand U1359 (N_1359,In_33,In_282);
and U1360 (N_1360,In_181,In_228);
nand U1361 (N_1361,In_364,In_121);
or U1362 (N_1362,In_512,In_403);
or U1363 (N_1363,In_456,In_192);
and U1364 (N_1364,In_450,In_44);
nand U1365 (N_1365,In_662,In_281);
or U1366 (N_1366,In_212,In_75);
nand U1367 (N_1367,In_478,In_537);
and U1368 (N_1368,In_166,In_412);
nand U1369 (N_1369,In_695,In_272);
nand U1370 (N_1370,In_403,In_548);
or U1371 (N_1371,In_296,In_644);
and U1372 (N_1372,In_507,In_411);
xnor U1373 (N_1373,In_240,In_145);
and U1374 (N_1374,In_633,In_426);
and U1375 (N_1375,In_368,In_308);
nor U1376 (N_1376,In_479,In_174);
nor U1377 (N_1377,In_137,In_448);
nor U1378 (N_1378,In_614,In_307);
nor U1379 (N_1379,In_318,In_398);
nor U1380 (N_1380,In_711,In_279);
nand U1381 (N_1381,In_415,In_371);
nand U1382 (N_1382,In_375,In_546);
nor U1383 (N_1383,In_193,In_643);
nor U1384 (N_1384,In_156,In_101);
xnor U1385 (N_1385,In_208,In_622);
nor U1386 (N_1386,In_453,In_656);
nand U1387 (N_1387,In_327,In_90);
or U1388 (N_1388,In_671,In_538);
nor U1389 (N_1389,In_596,In_455);
or U1390 (N_1390,In_91,In_179);
or U1391 (N_1391,In_233,In_122);
or U1392 (N_1392,In_141,In_187);
nor U1393 (N_1393,In_170,In_642);
nand U1394 (N_1394,In_139,In_564);
nand U1395 (N_1395,In_544,In_637);
and U1396 (N_1396,In_94,In_450);
nor U1397 (N_1397,In_391,In_123);
or U1398 (N_1398,In_274,In_689);
or U1399 (N_1399,In_514,In_545);
nand U1400 (N_1400,In_604,In_58);
nor U1401 (N_1401,In_174,In_182);
or U1402 (N_1402,In_335,In_268);
and U1403 (N_1403,In_581,In_34);
or U1404 (N_1404,In_681,In_747);
or U1405 (N_1405,In_268,In_392);
or U1406 (N_1406,In_135,In_440);
nor U1407 (N_1407,In_207,In_566);
nand U1408 (N_1408,In_389,In_72);
or U1409 (N_1409,In_678,In_13);
nand U1410 (N_1410,In_408,In_242);
or U1411 (N_1411,In_478,In_235);
nor U1412 (N_1412,In_83,In_444);
nand U1413 (N_1413,In_61,In_213);
nand U1414 (N_1414,In_100,In_355);
and U1415 (N_1415,In_389,In_74);
nor U1416 (N_1416,In_494,In_468);
and U1417 (N_1417,In_672,In_639);
nor U1418 (N_1418,In_444,In_657);
and U1419 (N_1419,In_133,In_343);
nand U1420 (N_1420,In_308,In_374);
nand U1421 (N_1421,In_281,In_474);
nor U1422 (N_1422,In_13,In_461);
and U1423 (N_1423,In_310,In_127);
or U1424 (N_1424,In_600,In_223);
and U1425 (N_1425,In_486,In_600);
nor U1426 (N_1426,In_706,In_519);
nand U1427 (N_1427,In_729,In_543);
nor U1428 (N_1428,In_583,In_373);
or U1429 (N_1429,In_690,In_94);
nand U1430 (N_1430,In_172,In_400);
and U1431 (N_1431,In_195,In_467);
xor U1432 (N_1432,In_553,In_286);
nand U1433 (N_1433,In_445,In_460);
nand U1434 (N_1434,In_153,In_740);
and U1435 (N_1435,In_443,In_141);
nand U1436 (N_1436,In_614,In_668);
or U1437 (N_1437,In_210,In_720);
nor U1438 (N_1438,In_310,In_509);
nor U1439 (N_1439,In_326,In_28);
nor U1440 (N_1440,In_333,In_547);
or U1441 (N_1441,In_739,In_47);
nor U1442 (N_1442,In_46,In_353);
or U1443 (N_1443,In_358,In_15);
nor U1444 (N_1444,In_515,In_447);
nor U1445 (N_1445,In_200,In_46);
nand U1446 (N_1446,In_30,In_422);
or U1447 (N_1447,In_729,In_68);
nand U1448 (N_1448,In_691,In_541);
or U1449 (N_1449,In_604,In_123);
and U1450 (N_1450,In_35,In_530);
and U1451 (N_1451,In_352,In_641);
nor U1452 (N_1452,In_440,In_394);
and U1453 (N_1453,In_441,In_678);
and U1454 (N_1454,In_703,In_452);
or U1455 (N_1455,In_304,In_55);
or U1456 (N_1456,In_665,In_462);
nor U1457 (N_1457,In_397,In_214);
nor U1458 (N_1458,In_60,In_316);
nand U1459 (N_1459,In_709,In_551);
nand U1460 (N_1460,In_557,In_470);
nand U1461 (N_1461,In_676,In_234);
nand U1462 (N_1462,In_605,In_283);
and U1463 (N_1463,In_137,In_74);
and U1464 (N_1464,In_612,In_152);
or U1465 (N_1465,In_31,In_26);
nand U1466 (N_1466,In_470,In_648);
nor U1467 (N_1467,In_188,In_290);
nor U1468 (N_1468,In_511,In_110);
or U1469 (N_1469,In_302,In_522);
nand U1470 (N_1470,In_346,In_5);
and U1471 (N_1471,In_507,In_331);
or U1472 (N_1472,In_49,In_485);
and U1473 (N_1473,In_24,In_30);
nor U1474 (N_1474,In_15,In_297);
and U1475 (N_1475,In_187,In_537);
nor U1476 (N_1476,In_267,In_718);
or U1477 (N_1477,In_499,In_22);
or U1478 (N_1478,In_197,In_204);
and U1479 (N_1479,In_687,In_382);
or U1480 (N_1480,In_518,In_233);
and U1481 (N_1481,In_642,In_53);
xor U1482 (N_1482,In_511,In_302);
and U1483 (N_1483,In_361,In_372);
nor U1484 (N_1484,In_57,In_463);
and U1485 (N_1485,In_70,In_182);
nand U1486 (N_1486,In_102,In_517);
nor U1487 (N_1487,In_32,In_86);
nor U1488 (N_1488,In_623,In_443);
nand U1489 (N_1489,In_742,In_75);
nand U1490 (N_1490,In_622,In_194);
nand U1491 (N_1491,In_30,In_573);
or U1492 (N_1492,In_283,In_433);
and U1493 (N_1493,In_195,In_690);
nor U1494 (N_1494,In_693,In_469);
and U1495 (N_1495,In_475,In_250);
nor U1496 (N_1496,In_234,In_662);
nand U1497 (N_1497,In_529,In_116);
and U1498 (N_1498,In_515,In_318);
nor U1499 (N_1499,In_341,In_130);
and U1500 (N_1500,In_545,In_221);
nor U1501 (N_1501,In_607,In_114);
nor U1502 (N_1502,In_267,In_477);
or U1503 (N_1503,In_87,In_645);
and U1504 (N_1504,In_316,In_245);
or U1505 (N_1505,In_283,In_490);
xnor U1506 (N_1506,In_98,In_674);
nand U1507 (N_1507,In_33,In_260);
nor U1508 (N_1508,In_141,In_744);
nand U1509 (N_1509,In_370,In_121);
nand U1510 (N_1510,In_714,In_0);
nand U1511 (N_1511,In_473,In_570);
or U1512 (N_1512,In_695,In_155);
nor U1513 (N_1513,In_22,In_75);
nor U1514 (N_1514,In_382,In_40);
and U1515 (N_1515,In_168,In_448);
or U1516 (N_1516,In_665,In_495);
nand U1517 (N_1517,In_603,In_66);
and U1518 (N_1518,In_199,In_49);
nand U1519 (N_1519,In_586,In_292);
nand U1520 (N_1520,In_126,In_131);
nand U1521 (N_1521,In_117,In_671);
nor U1522 (N_1522,In_88,In_716);
nor U1523 (N_1523,In_104,In_678);
or U1524 (N_1524,In_383,In_3);
nand U1525 (N_1525,In_357,In_81);
nor U1526 (N_1526,In_663,In_520);
and U1527 (N_1527,In_574,In_680);
or U1528 (N_1528,In_8,In_92);
nand U1529 (N_1529,In_403,In_358);
xnor U1530 (N_1530,In_6,In_337);
nor U1531 (N_1531,In_686,In_341);
or U1532 (N_1532,In_674,In_84);
nor U1533 (N_1533,In_218,In_212);
or U1534 (N_1534,In_321,In_237);
and U1535 (N_1535,In_301,In_233);
nand U1536 (N_1536,In_75,In_112);
and U1537 (N_1537,In_662,In_426);
and U1538 (N_1538,In_391,In_672);
nand U1539 (N_1539,In_540,In_395);
and U1540 (N_1540,In_588,In_423);
nor U1541 (N_1541,In_536,In_540);
nand U1542 (N_1542,In_383,In_234);
and U1543 (N_1543,In_707,In_734);
and U1544 (N_1544,In_680,In_246);
nor U1545 (N_1545,In_719,In_749);
nor U1546 (N_1546,In_680,In_73);
or U1547 (N_1547,In_93,In_468);
and U1548 (N_1548,In_629,In_735);
nor U1549 (N_1549,In_466,In_437);
nor U1550 (N_1550,In_119,In_137);
xnor U1551 (N_1551,In_641,In_30);
and U1552 (N_1552,In_226,In_332);
or U1553 (N_1553,In_371,In_248);
nor U1554 (N_1554,In_165,In_366);
nand U1555 (N_1555,In_106,In_601);
and U1556 (N_1556,In_100,In_115);
or U1557 (N_1557,In_296,In_45);
or U1558 (N_1558,In_383,In_538);
and U1559 (N_1559,In_616,In_504);
nor U1560 (N_1560,In_252,In_523);
and U1561 (N_1561,In_637,In_31);
nand U1562 (N_1562,In_270,In_51);
nor U1563 (N_1563,In_360,In_443);
and U1564 (N_1564,In_514,In_576);
or U1565 (N_1565,In_298,In_683);
and U1566 (N_1566,In_114,In_208);
or U1567 (N_1567,In_704,In_386);
and U1568 (N_1568,In_733,In_46);
or U1569 (N_1569,In_70,In_305);
nor U1570 (N_1570,In_486,In_506);
or U1571 (N_1571,In_581,In_475);
nor U1572 (N_1572,In_51,In_570);
and U1573 (N_1573,In_463,In_409);
or U1574 (N_1574,In_340,In_456);
and U1575 (N_1575,In_225,In_132);
and U1576 (N_1576,In_583,In_666);
nand U1577 (N_1577,In_214,In_148);
or U1578 (N_1578,In_549,In_667);
or U1579 (N_1579,In_112,In_478);
nor U1580 (N_1580,In_710,In_570);
nand U1581 (N_1581,In_272,In_210);
or U1582 (N_1582,In_379,In_221);
or U1583 (N_1583,In_278,In_536);
or U1584 (N_1584,In_612,In_81);
or U1585 (N_1585,In_253,In_155);
or U1586 (N_1586,In_143,In_700);
nor U1587 (N_1587,In_13,In_390);
and U1588 (N_1588,In_245,In_692);
and U1589 (N_1589,In_312,In_232);
nand U1590 (N_1590,In_267,In_429);
nor U1591 (N_1591,In_362,In_0);
nor U1592 (N_1592,In_633,In_648);
nor U1593 (N_1593,In_703,In_165);
nor U1594 (N_1594,In_415,In_262);
nand U1595 (N_1595,In_576,In_558);
and U1596 (N_1596,In_385,In_331);
or U1597 (N_1597,In_458,In_118);
and U1598 (N_1598,In_308,In_679);
nand U1599 (N_1599,In_7,In_160);
nor U1600 (N_1600,In_377,In_392);
nor U1601 (N_1601,In_0,In_68);
or U1602 (N_1602,In_476,In_57);
nor U1603 (N_1603,In_556,In_321);
and U1604 (N_1604,In_540,In_714);
nor U1605 (N_1605,In_709,In_336);
or U1606 (N_1606,In_592,In_535);
nand U1607 (N_1607,In_624,In_636);
and U1608 (N_1608,In_586,In_174);
nand U1609 (N_1609,In_161,In_649);
or U1610 (N_1610,In_12,In_214);
and U1611 (N_1611,In_619,In_740);
nor U1612 (N_1612,In_347,In_608);
and U1613 (N_1613,In_736,In_422);
or U1614 (N_1614,In_578,In_18);
nand U1615 (N_1615,In_299,In_618);
and U1616 (N_1616,In_657,In_246);
or U1617 (N_1617,In_98,In_568);
and U1618 (N_1618,In_559,In_454);
or U1619 (N_1619,In_114,In_634);
and U1620 (N_1620,In_536,In_493);
nor U1621 (N_1621,In_677,In_454);
or U1622 (N_1622,In_564,In_521);
nor U1623 (N_1623,In_210,In_705);
or U1624 (N_1624,In_430,In_132);
nand U1625 (N_1625,In_417,In_450);
nand U1626 (N_1626,In_414,In_625);
and U1627 (N_1627,In_301,In_715);
nand U1628 (N_1628,In_213,In_188);
nor U1629 (N_1629,In_309,In_748);
nor U1630 (N_1630,In_294,In_265);
nand U1631 (N_1631,In_467,In_406);
or U1632 (N_1632,In_144,In_576);
nor U1633 (N_1633,In_84,In_474);
and U1634 (N_1634,In_134,In_202);
nand U1635 (N_1635,In_305,In_474);
and U1636 (N_1636,In_247,In_310);
and U1637 (N_1637,In_675,In_102);
nand U1638 (N_1638,In_557,In_715);
and U1639 (N_1639,In_471,In_268);
nand U1640 (N_1640,In_559,In_71);
and U1641 (N_1641,In_329,In_655);
and U1642 (N_1642,In_98,In_420);
nand U1643 (N_1643,In_42,In_313);
or U1644 (N_1644,In_317,In_151);
and U1645 (N_1645,In_107,In_297);
or U1646 (N_1646,In_198,In_279);
nor U1647 (N_1647,In_368,In_53);
nand U1648 (N_1648,In_611,In_454);
nand U1649 (N_1649,In_529,In_206);
and U1650 (N_1650,In_72,In_393);
nor U1651 (N_1651,In_222,In_339);
nand U1652 (N_1652,In_577,In_522);
nor U1653 (N_1653,In_747,In_264);
nor U1654 (N_1654,In_736,In_297);
nand U1655 (N_1655,In_471,In_180);
and U1656 (N_1656,In_453,In_337);
and U1657 (N_1657,In_492,In_302);
nor U1658 (N_1658,In_486,In_669);
nand U1659 (N_1659,In_524,In_462);
and U1660 (N_1660,In_337,In_544);
or U1661 (N_1661,In_25,In_366);
nand U1662 (N_1662,In_310,In_448);
nor U1663 (N_1663,In_38,In_718);
and U1664 (N_1664,In_44,In_273);
nor U1665 (N_1665,In_83,In_475);
nand U1666 (N_1666,In_732,In_241);
or U1667 (N_1667,In_98,In_540);
or U1668 (N_1668,In_616,In_139);
and U1669 (N_1669,In_600,In_437);
nor U1670 (N_1670,In_493,In_617);
nor U1671 (N_1671,In_619,In_744);
nand U1672 (N_1672,In_167,In_651);
nor U1673 (N_1673,In_304,In_602);
or U1674 (N_1674,In_115,In_327);
and U1675 (N_1675,In_238,In_134);
nor U1676 (N_1676,In_564,In_329);
nor U1677 (N_1677,In_465,In_1);
and U1678 (N_1678,In_21,In_220);
nor U1679 (N_1679,In_208,In_680);
xor U1680 (N_1680,In_238,In_182);
and U1681 (N_1681,In_74,In_704);
nor U1682 (N_1682,In_507,In_199);
nand U1683 (N_1683,In_449,In_437);
and U1684 (N_1684,In_286,In_507);
nor U1685 (N_1685,In_667,In_236);
nand U1686 (N_1686,In_266,In_391);
nor U1687 (N_1687,In_430,In_257);
or U1688 (N_1688,In_17,In_695);
and U1689 (N_1689,In_748,In_25);
or U1690 (N_1690,In_336,In_518);
or U1691 (N_1691,In_251,In_146);
and U1692 (N_1692,In_236,In_250);
nand U1693 (N_1693,In_629,In_517);
nand U1694 (N_1694,In_688,In_94);
nand U1695 (N_1695,In_165,In_10);
nor U1696 (N_1696,In_290,In_472);
or U1697 (N_1697,In_473,In_480);
and U1698 (N_1698,In_237,In_542);
nor U1699 (N_1699,In_2,In_125);
nor U1700 (N_1700,In_327,In_215);
and U1701 (N_1701,In_298,In_462);
or U1702 (N_1702,In_650,In_371);
nand U1703 (N_1703,In_529,In_666);
nor U1704 (N_1704,In_543,In_276);
nor U1705 (N_1705,In_52,In_231);
nand U1706 (N_1706,In_621,In_80);
and U1707 (N_1707,In_378,In_4);
or U1708 (N_1708,In_274,In_177);
and U1709 (N_1709,In_708,In_50);
and U1710 (N_1710,In_145,In_373);
nand U1711 (N_1711,In_566,In_512);
nand U1712 (N_1712,In_464,In_64);
nor U1713 (N_1713,In_73,In_134);
and U1714 (N_1714,In_316,In_298);
nor U1715 (N_1715,In_163,In_302);
or U1716 (N_1716,In_516,In_120);
nand U1717 (N_1717,In_271,In_684);
or U1718 (N_1718,In_293,In_47);
xor U1719 (N_1719,In_76,In_465);
or U1720 (N_1720,In_233,In_528);
xor U1721 (N_1721,In_678,In_1);
and U1722 (N_1722,In_73,In_43);
nor U1723 (N_1723,In_125,In_67);
nand U1724 (N_1724,In_467,In_28);
nor U1725 (N_1725,In_451,In_519);
nand U1726 (N_1726,In_72,In_480);
or U1727 (N_1727,In_627,In_220);
nand U1728 (N_1728,In_504,In_216);
nand U1729 (N_1729,In_640,In_212);
nand U1730 (N_1730,In_19,In_26);
nand U1731 (N_1731,In_160,In_376);
nor U1732 (N_1732,In_259,In_438);
nand U1733 (N_1733,In_596,In_185);
nor U1734 (N_1734,In_107,In_607);
and U1735 (N_1735,In_39,In_171);
nand U1736 (N_1736,In_565,In_657);
xor U1737 (N_1737,In_452,In_117);
nor U1738 (N_1738,In_556,In_4);
xor U1739 (N_1739,In_561,In_676);
nand U1740 (N_1740,In_188,In_247);
nand U1741 (N_1741,In_338,In_434);
nand U1742 (N_1742,In_189,In_618);
nor U1743 (N_1743,In_563,In_112);
nor U1744 (N_1744,In_628,In_722);
nor U1745 (N_1745,In_3,In_572);
xnor U1746 (N_1746,In_349,In_185);
xor U1747 (N_1747,In_256,In_292);
nor U1748 (N_1748,In_327,In_685);
nor U1749 (N_1749,In_161,In_437);
nor U1750 (N_1750,In_708,In_456);
nand U1751 (N_1751,In_72,In_49);
xnor U1752 (N_1752,In_80,In_708);
nand U1753 (N_1753,In_701,In_191);
and U1754 (N_1754,In_80,In_564);
and U1755 (N_1755,In_243,In_364);
and U1756 (N_1756,In_558,In_38);
nor U1757 (N_1757,In_32,In_575);
nand U1758 (N_1758,In_102,In_193);
nand U1759 (N_1759,In_612,In_270);
or U1760 (N_1760,In_46,In_681);
nand U1761 (N_1761,In_384,In_314);
nand U1762 (N_1762,In_97,In_657);
nor U1763 (N_1763,In_673,In_383);
or U1764 (N_1764,In_501,In_122);
or U1765 (N_1765,In_557,In_454);
or U1766 (N_1766,In_501,In_97);
nor U1767 (N_1767,In_468,In_178);
nand U1768 (N_1768,In_539,In_749);
nand U1769 (N_1769,In_47,In_234);
and U1770 (N_1770,In_57,In_411);
nand U1771 (N_1771,In_426,In_742);
and U1772 (N_1772,In_746,In_213);
nand U1773 (N_1773,In_177,In_490);
nor U1774 (N_1774,In_45,In_164);
nor U1775 (N_1775,In_680,In_600);
and U1776 (N_1776,In_320,In_268);
nor U1777 (N_1777,In_229,In_84);
and U1778 (N_1778,In_345,In_237);
or U1779 (N_1779,In_676,In_199);
nand U1780 (N_1780,In_187,In_191);
nor U1781 (N_1781,In_630,In_573);
nor U1782 (N_1782,In_305,In_74);
or U1783 (N_1783,In_211,In_641);
and U1784 (N_1784,In_288,In_120);
nor U1785 (N_1785,In_521,In_725);
nand U1786 (N_1786,In_472,In_95);
or U1787 (N_1787,In_491,In_553);
nand U1788 (N_1788,In_354,In_51);
or U1789 (N_1789,In_683,In_57);
xnor U1790 (N_1790,In_355,In_28);
or U1791 (N_1791,In_294,In_23);
nand U1792 (N_1792,In_148,In_729);
or U1793 (N_1793,In_105,In_561);
nor U1794 (N_1794,In_470,In_37);
or U1795 (N_1795,In_642,In_80);
and U1796 (N_1796,In_602,In_185);
and U1797 (N_1797,In_197,In_647);
and U1798 (N_1798,In_642,In_69);
or U1799 (N_1799,In_635,In_456);
and U1800 (N_1800,In_245,In_578);
and U1801 (N_1801,In_726,In_522);
nand U1802 (N_1802,In_87,In_293);
and U1803 (N_1803,In_59,In_447);
nand U1804 (N_1804,In_465,In_503);
nor U1805 (N_1805,In_164,In_18);
and U1806 (N_1806,In_315,In_136);
nor U1807 (N_1807,In_711,In_340);
or U1808 (N_1808,In_79,In_280);
nand U1809 (N_1809,In_159,In_483);
nor U1810 (N_1810,In_303,In_131);
and U1811 (N_1811,In_20,In_577);
nand U1812 (N_1812,In_436,In_181);
nor U1813 (N_1813,In_325,In_399);
xnor U1814 (N_1814,In_197,In_165);
nand U1815 (N_1815,In_303,In_317);
nor U1816 (N_1816,In_715,In_167);
nor U1817 (N_1817,In_386,In_593);
nor U1818 (N_1818,In_267,In_699);
and U1819 (N_1819,In_744,In_356);
and U1820 (N_1820,In_245,In_358);
and U1821 (N_1821,In_454,In_493);
or U1822 (N_1822,In_281,In_199);
nor U1823 (N_1823,In_43,In_224);
and U1824 (N_1824,In_67,In_656);
and U1825 (N_1825,In_413,In_115);
or U1826 (N_1826,In_36,In_341);
or U1827 (N_1827,In_595,In_694);
or U1828 (N_1828,In_745,In_665);
and U1829 (N_1829,In_702,In_724);
and U1830 (N_1830,In_336,In_48);
nor U1831 (N_1831,In_193,In_118);
nor U1832 (N_1832,In_205,In_514);
nand U1833 (N_1833,In_198,In_361);
nor U1834 (N_1834,In_405,In_352);
or U1835 (N_1835,In_97,In_47);
and U1836 (N_1836,In_543,In_411);
or U1837 (N_1837,In_119,In_42);
or U1838 (N_1838,In_71,In_645);
nand U1839 (N_1839,In_716,In_358);
or U1840 (N_1840,In_728,In_388);
or U1841 (N_1841,In_29,In_495);
or U1842 (N_1842,In_563,In_574);
or U1843 (N_1843,In_27,In_47);
nand U1844 (N_1844,In_550,In_180);
nand U1845 (N_1845,In_404,In_673);
and U1846 (N_1846,In_743,In_291);
nand U1847 (N_1847,In_143,In_229);
xor U1848 (N_1848,In_613,In_684);
nand U1849 (N_1849,In_233,In_42);
nor U1850 (N_1850,In_620,In_726);
and U1851 (N_1851,In_329,In_478);
or U1852 (N_1852,In_633,In_157);
nor U1853 (N_1853,In_429,In_350);
nand U1854 (N_1854,In_496,In_192);
xnor U1855 (N_1855,In_215,In_662);
or U1856 (N_1856,In_138,In_195);
or U1857 (N_1857,In_441,In_356);
and U1858 (N_1858,In_458,In_465);
nand U1859 (N_1859,In_494,In_438);
or U1860 (N_1860,In_333,In_521);
nand U1861 (N_1861,In_545,In_670);
and U1862 (N_1862,In_372,In_288);
or U1863 (N_1863,In_324,In_243);
and U1864 (N_1864,In_740,In_432);
or U1865 (N_1865,In_669,In_34);
nand U1866 (N_1866,In_438,In_415);
or U1867 (N_1867,In_610,In_20);
nor U1868 (N_1868,In_91,In_102);
nor U1869 (N_1869,In_674,In_565);
and U1870 (N_1870,In_124,In_356);
or U1871 (N_1871,In_651,In_691);
nor U1872 (N_1872,In_98,In_55);
and U1873 (N_1873,In_351,In_301);
and U1874 (N_1874,In_167,In_26);
nand U1875 (N_1875,In_625,In_598);
or U1876 (N_1876,In_364,In_18);
nor U1877 (N_1877,In_73,In_325);
nor U1878 (N_1878,In_539,In_698);
nor U1879 (N_1879,In_295,In_314);
nand U1880 (N_1880,In_365,In_454);
nand U1881 (N_1881,In_378,In_557);
and U1882 (N_1882,In_423,In_421);
and U1883 (N_1883,In_109,In_682);
and U1884 (N_1884,In_688,In_721);
nor U1885 (N_1885,In_83,In_629);
or U1886 (N_1886,In_496,In_380);
nor U1887 (N_1887,In_128,In_699);
nand U1888 (N_1888,In_221,In_380);
nor U1889 (N_1889,In_723,In_538);
and U1890 (N_1890,In_19,In_135);
xnor U1891 (N_1891,In_374,In_577);
and U1892 (N_1892,In_515,In_671);
nor U1893 (N_1893,In_530,In_272);
nor U1894 (N_1894,In_39,In_215);
nor U1895 (N_1895,In_486,In_460);
or U1896 (N_1896,In_384,In_18);
and U1897 (N_1897,In_660,In_601);
and U1898 (N_1898,In_550,In_461);
nor U1899 (N_1899,In_223,In_304);
and U1900 (N_1900,In_356,In_718);
nor U1901 (N_1901,In_222,In_371);
nand U1902 (N_1902,In_502,In_477);
or U1903 (N_1903,In_34,In_530);
nor U1904 (N_1904,In_212,In_589);
nor U1905 (N_1905,In_290,In_333);
nor U1906 (N_1906,In_338,In_74);
nand U1907 (N_1907,In_121,In_211);
nor U1908 (N_1908,In_668,In_189);
nor U1909 (N_1909,In_227,In_203);
nor U1910 (N_1910,In_612,In_509);
and U1911 (N_1911,In_212,In_96);
or U1912 (N_1912,In_354,In_313);
and U1913 (N_1913,In_614,In_110);
xor U1914 (N_1914,In_468,In_498);
xor U1915 (N_1915,In_428,In_88);
or U1916 (N_1916,In_430,In_335);
nand U1917 (N_1917,In_662,In_449);
and U1918 (N_1918,In_107,In_188);
or U1919 (N_1919,In_202,In_178);
and U1920 (N_1920,In_56,In_354);
or U1921 (N_1921,In_107,In_15);
nor U1922 (N_1922,In_411,In_651);
and U1923 (N_1923,In_345,In_537);
or U1924 (N_1924,In_339,In_459);
nor U1925 (N_1925,In_497,In_605);
and U1926 (N_1926,In_293,In_208);
nor U1927 (N_1927,In_128,In_435);
and U1928 (N_1928,In_206,In_466);
or U1929 (N_1929,In_295,In_605);
nor U1930 (N_1930,In_183,In_572);
and U1931 (N_1931,In_77,In_343);
nand U1932 (N_1932,In_594,In_643);
nor U1933 (N_1933,In_718,In_351);
and U1934 (N_1934,In_22,In_44);
nand U1935 (N_1935,In_116,In_683);
or U1936 (N_1936,In_299,In_366);
or U1937 (N_1937,In_9,In_438);
or U1938 (N_1938,In_238,In_669);
or U1939 (N_1939,In_217,In_695);
nor U1940 (N_1940,In_466,In_554);
or U1941 (N_1941,In_227,In_211);
and U1942 (N_1942,In_497,In_300);
or U1943 (N_1943,In_342,In_256);
nand U1944 (N_1944,In_56,In_153);
and U1945 (N_1945,In_299,In_94);
nand U1946 (N_1946,In_437,In_507);
and U1947 (N_1947,In_229,In_554);
nor U1948 (N_1948,In_347,In_678);
nand U1949 (N_1949,In_22,In_48);
nand U1950 (N_1950,In_121,In_38);
or U1951 (N_1951,In_532,In_711);
and U1952 (N_1952,In_340,In_363);
nor U1953 (N_1953,In_396,In_685);
nor U1954 (N_1954,In_360,In_287);
nor U1955 (N_1955,In_147,In_218);
and U1956 (N_1956,In_365,In_687);
or U1957 (N_1957,In_2,In_239);
or U1958 (N_1958,In_75,In_314);
or U1959 (N_1959,In_709,In_476);
or U1960 (N_1960,In_90,In_618);
nand U1961 (N_1961,In_663,In_572);
nor U1962 (N_1962,In_582,In_401);
and U1963 (N_1963,In_682,In_400);
and U1964 (N_1964,In_456,In_1);
nand U1965 (N_1965,In_422,In_157);
nand U1966 (N_1966,In_345,In_231);
nand U1967 (N_1967,In_265,In_254);
nand U1968 (N_1968,In_208,In_253);
or U1969 (N_1969,In_586,In_607);
xnor U1970 (N_1970,In_616,In_679);
nand U1971 (N_1971,In_671,In_360);
and U1972 (N_1972,In_696,In_408);
nand U1973 (N_1973,In_497,In_513);
nor U1974 (N_1974,In_53,In_690);
nand U1975 (N_1975,In_387,In_429);
nor U1976 (N_1976,In_303,In_348);
nor U1977 (N_1977,In_634,In_538);
and U1978 (N_1978,In_693,In_523);
nand U1979 (N_1979,In_422,In_40);
nor U1980 (N_1980,In_429,In_151);
and U1981 (N_1981,In_29,In_399);
nor U1982 (N_1982,In_547,In_68);
and U1983 (N_1983,In_287,In_589);
nand U1984 (N_1984,In_371,In_149);
nand U1985 (N_1985,In_78,In_212);
nand U1986 (N_1986,In_78,In_567);
nor U1987 (N_1987,In_399,In_126);
and U1988 (N_1988,In_453,In_336);
nand U1989 (N_1989,In_498,In_382);
nand U1990 (N_1990,In_157,In_744);
and U1991 (N_1991,In_357,In_689);
and U1992 (N_1992,In_678,In_184);
nor U1993 (N_1993,In_349,In_421);
and U1994 (N_1994,In_707,In_369);
nand U1995 (N_1995,In_686,In_46);
nand U1996 (N_1996,In_525,In_646);
nor U1997 (N_1997,In_337,In_504);
and U1998 (N_1998,In_294,In_748);
xnor U1999 (N_1999,In_119,In_354);
and U2000 (N_2000,In_77,In_531);
and U2001 (N_2001,In_350,In_273);
nor U2002 (N_2002,In_383,In_142);
nand U2003 (N_2003,In_5,In_236);
nor U2004 (N_2004,In_369,In_635);
and U2005 (N_2005,In_320,In_608);
and U2006 (N_2006,In_305,In_338);
and U2007 (N_2007,In_561,In_696);
and U2008 (N_2008,In_63,In_324);
nand U2009 (N_2009,In_501,In_141);
nor U2010 (N_2010,In_458,In_309);
nor U2011 (N_2011,In_621,In_562);
nor U2012 (N_2012,In_39,In_544);
nor U2013 (N_2013,In_670,In_376);
nand U2014 (N_2014,In_214,In_271);
and U2015 (N_2015,In_338,In_286);
nand U2016 (N_2016,In_35,In_704);
nand U2017 (N_2017,In_601,In_649);
nand U2018 (N_2018,In_233,In_52);
or U2019 (N_2019,In_625,In_722);
and U2020 (N_2020,In_263,In_741);
nor U2021 (N_2021,In_14,In_274);
and U2022 (N_2022,In_144,In_472);
or U2023 (N_2023,In_538,In_49);
nand U2024 (N_2024,In_739,In_245);
or U2025 (N_2025,In_466,In_325);
nor U2026 (N_2026,In_493,In_139);
or U2027 (N_2027,In_682,In_92);
nand U2028 (N_2028,In_41,In_142);
or U2029 (N_2029,In_545,In_418);
nor U2030 (N_2030,In_410,In_611);
or U2031 (N_2031,In_608,In_483);
nand U2032 (N_2032,In_145,In_503);
nor U2033 (N_2033,In_32,In_221);
nor U2034 (N_2034,In_605,In_98);
and U2035 (N_2035,In_718,In_101);
nand U2036 (N_2036,In_547,In_469);
nor U2037 (N_2037,In_26,In_652);
nor U2038 (N_2038,In_317,In_328);
or U2039 (N_2039,In_570,In_573);
nand U2040 (N_2040,In_578,In_114);
nor U2041 (N_2041,In_701,In_499);
and U2042 (N_2042,In_32,In_190);
and U2043 (N_2043,In_465,In_725);
nor U2044 (N_2044,In_440,In_174);
nor U2045 (N_2045,In_76,In_587);
or U2046 (N_2046,In_50,In_35);
or U2047 (N_2047,In_633,In_341);
nor U2048 (N_2048,In_342,In_287);
and U2049 (N_2049,In_627,In_579);
nor U2050 (N_2050,In_720,In_219);
nand U2051 (N_2051,In_654,In_4);
and U2052 (N_2052,In_454,In_200);
nand U2053 (N_2053,In_542,In_388);
nor U2054 (N_2054,In_250,In_503);
nor U2055 (N_2055,In_219,In_532);
nor U2056 (N_2056,In_151,In_399);
nand U2057 (N_2057,In_245,In_510);
or U2058 (N_2058,In_536,In_524);
xnor U2059 (N_2059,In_571,In_677);
nor U2060 (N_2060,In_188,In_216);
nand U2061 (N_2061,In_385,In_569);
nand U2062 (N_2062,In_641,In_736);
nor U2063 (N_2063,In_88,In_224);
or U2064 (N_2064,In_422,In_448);
and U2065 (N_2065,In_162,In_338);
xor U2066 (N_2066,In_578,In_279);
nand U2067 (N_2067,In_651,In_353);
or U2068 (N_2068,In_343,In_542);
nand U2069 (N_2069,In_397,In_143);
or U2070 (N_2070,In_36,In_27);
or U2071 (N_2071,In_48,In_196);
and U2072 (N_2072,In_219,In_30);
and U2073 (N_2073,In_394,In_452);
and U2074 (N_2074,In_709,In_307);
or U2075 (N_2075,In_542,In_722);
nand U2076 (N_2076,In_245,In_333);
and U2077 (N_2077,In_700,In_556);
or U2078 (N_2078,In_369,In_595);
nor U2079 (N_2079,In_330,In_452);
nor U2080 (N_2080,In_653,In_334);
nor U2081 (N_2081,In_117,In_584);
nor U2082 (N_2082,In_29,In_732);
nor U2083 (N_2083,In_311,In_241);
or U2084 (N_2084,In_386,In_430);
nand U2085 (N_2085,In_576,In_686);
nor U2086 (N_2086,In_266,In_573);
nand U2087 (N_2087,In_357,In_623);
or U2088 (N_2088,In_210,In_208);
nor U2089 (N_2089,In_216,In_175);
nand U2090 (N_2090,In_689,In_334);
nand U2091 (N_2091,In_412,In_237);
or U2092 (N_2092,In_685,In_664);
nand U2093 (N_2093,In_67,In_9);
or U2094 (N_2094,In_489,In_709);
and U2095 (N_2095,In_387,In_366);
nor U2096 (N_2096,In_556,In_648);
or U2097 (N_2097,In_154,In_603);
nor U2098 (N_2098,In_236,In_520);
and U2099 (N_2099,In_618,In_677);
and U2100 (N_2100,In_587,In_674);
nand U2101 (N_2101,In_58,In_729);
nand U2102 (N_2102,In_482,In_389);
nor U2103 (N_2103,In_206,In_602);
or U2104 (N_2104,In_246,In_312);
nor U2105 (N_2105,In_221,In_305);
or U2106 (N_2106,In_141,In_330);
nand U2107 (N_2107,In_339,In_442);
and U2108 (N_2108,In_498,In_288);
nor U2109 (N_2109,In_626,In_297);
nor U2110 (N_2110,In_207,In_84);
nand U2111 (N_2111,In_404,In_605);
and U2112 (N_2112,In_552,In_692);
nor U2113 (N_2113,In_511,In_187);
and U2114 (N_2114,In_531,In_247);
or U2115 (N_2115,In_308,In_730);
or U2116 (N_2116,In_663,In_418);
nor U2117 (N_2117,In_46,In_441);
and U2118 (N_2118,In_683,In_340);
and U2119 (N_2119,In_395,In_26);
nand U2120 (N_2120,In_77,In_434);
and U2121 (N_2121,In_646,In_620);
nor U2122 (N_2122,In_74,In_106);
or U2123 (N_2123,In_300,In_559);
and U2124 (N_2124,In_529,In_33);
and U2125 (N_2125,In_81,In_724);
nand U2126 (N_2126,In_543,In_432);
nor U2127 (N_2127,In_688,In_351);
nand U2128 (N_2128,In_339,In_101);
or U2129 (N_2129,In_491,In_208);
nand U2130 (N_2130,In_242,In_471);
xnor U2131 (N_2131,In_359,In_399);
and U2132 (N_2132,In_14,In_72);
nor U2133 (N_2133,In_349,In_345);
nor U2134 (N_2134,In_468,In_549);
or U2135 (N_2135,In_203,In_591);
or U2136 (N_2136,In_400,In_438);
and U2137 (N_2137,In_83,In_417);
nor U2138 (N_2138,In_20,In_605);
nand U2139 (N_2139,In_66,In_23);
or U2140 (N_2140,In_302,In_169);
or U2141 (N_2141,In_570,In_338);
or U2142 (N_2142,In_485,In_694);
nor U2143 (N_2143,In_557,In_66);
or U2144 (N_2144,In_90,In_326);
or U2145 (N_2145,In_317,In_440);
and U2146 (N_2146,In_245,In_61);
xnor U2147 (N_2147,In_484,In_716);
and U2148 (N_2148,In_536,In_262);
nor U2149 (N_2149,In_494,In_78);
nand U2150 (N_2150,In_330,In_536);
or U2151 (N_2151,In_363,In_46);
nor U2152 (N_2152,In_600,In_168);
or U2153 (N_2153,In_44,In_585);
nor U2154 (N_2154,In_369,In_275);
or U2155 (N_2155,In_89,In_269);
xnor U2156 (N_2156,In_607,In_141);
or U2157 (N_2157,In_323,In_26);
and U2158 (N_2158,In_715,In_321);
nand U2159 (N_2159,In_107,In_247);
or U2160 (N_2160,In_58,In_665);
or U2161 (N_2161,In_531,In_166);
nand U2162 (N_2162,In_659,In_477);
nand U2163 (N_2163,In_619,In_6);
nor U2164 (N_2164,In_360,In_436);
nand U2165 (N_2165,In_561,In_52);
and U2166 (N_2166,In_666,In_408);
and U2167 (N_2167,In_409,In_708);
nand U2168 (N_2168,In_652,In_13);
nor U2169 (N_2169,In_67,In_336);
nor U2170 (N_2170,In_511,In_532);
or U2171 (N_2171,In_32,In_106);
nor U2172 (N_2172,In_395,In_671);
nand U2173 (N_2173,In_338,In_623);
nand U2174 (N_2174,In_373,In_518);
or U2175 (N_2175,In_171,In_668);
nor U2176 (N_2176,In_217,In_283);
xor U2177 (N_2177,In_9,In_688);
or U2178 (N_2178,In_285,In_76);
and U2179 (N_2179,In_547,In_614);
nor U2180 (N_2180,In_177,In_22);
nand U2181 (N_2181,In_447,In_657);
nor U2182 (N_2182,In_92,In_503);
or U2183 (N_2183,In_650,In_539);
nand U2184 (N_2184,In_249,In_704);
and U2185 (N_2185,In_562,In_214);
nor U2186 (N_2186,In_570,In_238);
nand U2187 (N_2187,In_233,In_566);
nand U2188 (N_2188,In_24,In_564);
nor U2189 (N_2189,In_453,In_335);
or U2190 (N_2190,In_396,In_605);
and U2191 (N_2191,In_628,In_42);
nor U2192 (N_2192,In_171,In_590);
and U2193 (N_2193,In_439,In_145);
nor U2194 (N_2194,In_250,In_516);
nor U2195 (N_2195,In_740,In_286);
and U2196 (N_2196,In_530,In_93);
nor U2197 (N_2197,In_634,In_326);
and U2198 (N_2198,In_314,In_632);
nand U2199 (N_2199,In_220,In_414);
and U2200 (N_2200,In_128,In_32);
and U2201 (N_2201,In_42,In_396);
or U2202 (N_2202,In_459,In_284);
or U2203 (N_2203,In_363,In_613);
nor U2204 (N_2204,In_329,In_531);
nand U2205 (N_2205,In_204,In_576);
nor U2206 (N_2206,In_735,In_631);
nor U2207 (N_2207,In_144,In_182);
and U2208 (N_2208,In_129,In_82);
or U2209 (N_2209,In_382,In_639);
or U2210 (N_2210,In_279,In_248);
nand U2211 (N_2211,In_241,In_391);
nor U2212 (N_2212,In_123,In_442);
nor U2213 (N_2213,In_583,In_678);
nor U2214 (N_2214,In_137,In_688);
or U2215 (N_2215,In_234,In_111);
nand U2216 (N_2216,In_307,In_148);
nor U2217 (N_2217,In_343,In_56);
and U2218 (N_2218,In_348,In_527);
and U2219 (N_2219,In_496,In_157);
nor U2220 (N_2220,In_386,In_210);
and U2221 (N_2221,In_221,In_708);
or U2222 (N_2222,In_46,In_348);
or U2223 (N_2223,In_182,In_608);
and U2224 (N_2224,In_717,In_542);
or U2225 (N_2225,In_668,In_323);
nor U2226 (N_2226,In_46,In_326);
and U2227 (N_2227,In_596,In_218);
nor U2228 (N_2228,In_382,In_418);
or U2229 (N_2229,In_501,In_424);
or U2230 (N_2230,In_549,In_708);
nand U2231 (N_2231,In_444,In_502);
nor U2232 (N_2232,In_666,In_39);
and U2233 (N_2233,In_11,In_444);
nand U2234 (N_2234,In_144,In_678);
nand U2235 (N_2235,In_504,In_21);
nand U2236 (N_2236,In_100,In_536);
nand U2237 (N_2237,In_604,In_127);
nand U2238 (N_2238,In_74,In_97);
or U2239 (N_2239,In_647,In_193);
or U2240 (N_2240,In_489,In_280);
or U2241 (N_2241,In_195,In_645);
and U2242 (N_2242,In_305,In_593);
nand U2243 (N_2243,In_721,In_360);
nand U2244 (N_2244,In_604,In_454);
nand U2245 (N_2245,In_283,In_258);
or U2246 (N_2246,In_436,In_33);
and U2247 (N_2247,In_528,In_306);
nor U2248 (N_2248,In_330,In_622);
nor U2249 (N_2249,In_535,In_62);
and U2250 (N_2250,In_87,In_113);
nor U2251 (N_2251,In_243,In_249);
or U2252 (N_2252,In_59,In_287);
and U2253 (N_2253,In_498,In_299);
nor U2254 (N_2254,In_107,In_108);
xor U2255 (N_2255,In_443,In_679);
and U2256 (N_2256,In_38,In_490);
and U2257 (N_2257,In_35,In_526);
nor U2258 (N_2258,In_348,In_533);
nor U2259 (N_2259,In_637,In_130);
or U2260 (N_2260,In_508,In_644);
nand U2261 (N_2261,In_42,In_363);
and U2262 (N_2262,In_379,In_586);
nor U2263 (N_2263,In_683,In_321);
and U2264 (N_2264,In_492,In_382);
nor U2265 (N_2265,In_473,In_584);
nand U2266 (N_2266,In_587,In_605);
nand U2267 (N_2267,In_511,In_3);
nand U2268 (N_2268,In_466,In_428);
nor U2269 (N_2269,In_437,In_199);
and U2270 (N_2270,In_305,In_95);
nor U2271 (N_2271,In_586,In_588);
nand U2272 (N_2272,In_481,In_252);
nand U2273 (N_2273,In_1,In_618);
nor U2274 (N_2274,In_10,In_718);
nand U2275 (N_2275,In_34,In_75);
and U2276 (N_2276,In_394,In_622);
nor U2277 (N_2277,In_666,In_530);
nor U2278 (N_2278,In_468,In_541);
nand U2279 (N_2279,In_605,In_656);
nor U2280 (N_2280,In_598,In_649);
nor U2281 (N_2281,In_124,In_305);
or U2282 (N_2282,In_85,In_129);
xnor U2283 (N_2283,In_627,In_190);
nand U2284 (N_2284,In_739,In_153);
nor U2285 (N_2285,In_607,In_157);
and U2286 (N_2286,In_540,In_32);
and U2287 (N_2287,In_432,In_93);
nor U2288 (N_2288,In_378,In_718);
or U2289 (N_2289,In_2,In_353);
and U2290 (N_2290,In_655,In_74);
nand U2291 (N_2291,In_623,In_452);
nand U2292 (N_2292,In_704,In_301);
and U2293 (N_2293,In_571,In_379);
or U2294 (N_2294,In_298,In_730);
nand U2295 (N_2295,In_284,In_396);
nor U2296 (N_2296,In_160,In_162);
nand U2297 (N_2297,In_44,In_708);
and U2298 (N_2298,In_388,In_300);
and U2299 (N_2299,In_196,In_216);
or U2300 (N_2300,In_153,In_259);
nand U2301 (N_2301,In_728,In_614);
nor U2302 (N_2302,In_8,In_581);
nand U2303 (N_2303,In_129,In_191);
nand U2304 (N_2304,In_509,In_340);
and U2305 (N_2305,In_362,In_130);
nand U2306 (N_2306,In_1,In_144);
nand U2307 (N_2307,In_164,In_322);
nor U2308 (N_2308,In_748,In_407);
nand U2309 (N_2309,In_172,In_64);
nor U2310 (N_2310,In_289,In_221);
or U2311 (N_2311,In_209,In_73);
nand U2312 (N_2312,In_720,In_533);
and U2313 (N_2313,In_645,In_355);
and U2314 (N_2314,In_593,In_425);
nor U2315 (N_2315,In_551,In_63);
nand U2316 (N_2316,In_9,In_235);
or U2317 (N_2317,In_9,In_103);
and U2318 (N_2318,In_699,In_563);
or U2319 (N_2319,In_301,In_279);
nand U2320 (N_2320,In_739,In_39);
nand U2321 (N_2321,In_300,In_212);
or U2322 (N_2322,In_669,In_3);
and U2323 (N_2323,In_236,In_314);
nor U2324 (N_2324,In_494,In_346);
nand U2325 (N_2325,In_367,In_653);
nor U2326 (N_2326,In_152,In_284);
and U2327 (N_2327,In_487,In_283);
or U2328 (N_2328,In_78,In_711);
and U2329 (N_2329,In_493,In_698);
xnor U2330 (N_2330,In_121,In_63);
nor U2331 (N_2331,In_643,In_244);
or U2332 (N_2332,In_242,In_562);
nand U2333 (N_2333,In_290,In_639);
nand U2334 (N_2334,In_220,In_714);
nor U2335 (N_2335,In_192,In_138);
or U2336 (N_2336,In_93,In_187);
nand U2337 (N_2337,In_601,In_28);
and U2338 (N_2338,In_232,In_364);
nand U2339 (N_2339,In_719,In_664);
nor U2340 (N_2340,In_37,In_508);
nand U2341 (N_2341,In_203,In_471);
or U2342 (N_2342,In_746,In_456);
and U2343 (N_2343,In_350,In_411);
and U2344 (N_2344,In_142,In_273);
and U2345 (N_2345,In_439,In_444);
nor U2346 (N_2346,In_681,In_565);
and U2347 (N_2347,In_145,In_47);
and U2348 (N_2348,In_182,In_69);
nor U2349 (N_2349,In_724,In_657);
and U2350 (N_2350,In_658,In_476);
nand U2351 (N_2351,In_712,In_689);
nor U2352 (N_2352,In_489,In_135);
nor U2353 (N_2353,In_659,In_440);
and U2354 (N_2354,In_199,In_68);
nand U2355 (N_2355,In_631,In_692);
or U2356 (N_2356,In_440,In_505);
and U2357 (N_2357,In_169,In_550);
and U2358 (N_2358,In_506,In_575);
and U2359 (N_2359,In_523,In_691);
nand U2360 (N_2360,In_722,In_69);
nand U2361 (N_2361,In_517,In_9);
nand U2362 (N_2362,In_335,In_44);
and U2363 (N_2363,In_398,In_475);
or U2364 (N_2364,In_153,In_276);
nand U2365 (N_2365,In_130,In_354);
or U2366 (N_2366,In_4,In_409);
or U2367 (N_2367,In_131,In_233);
or U2368 (N_2368,In_637,In_351);
or U2369 (N_2369,In_85,In_154);
and U2370 (N_2370,In_440,In_337);
nand U2371 (N_2371,In_258,In_70);
or U2372 (N_2372,In_232,In_329);
nand U2373 (N_2373,In_529,In_40);
nand U2374 (N_2374,In_306,In_401);
nor U2375 (N_2375,In_748,In_258);
or U2376 (N_2376,In_249,In_350);
nor U2377 (N_2377,In_537,In_394);
nand U2378 (N_2378,In_350,In_666);
nor U2379 (N_2379,In_76,In_369);
and U2380 (N_2380,In_743,In_127);
or U2381 (N_2381,In_207,In_9);
and U2382 (N_2382,In_12,In_312);
xnor U2383 (N_2383,In_308,In_742);
or U2384 (N_2384,In_223,In_126);
nor U2385 (N_2385,In_386,In_380);
nand U2386 (N_2386,In_338,In_65);
and U2387 (N_2387,In_214,In_698);
nand U2388 (N_2388,In_120,In_126);
or U2389 (N_2389,In_60,In_139);
or U2390 (N_2390,In_270,In_414);
and U2391 (N_2391,In_150,In_579);
xnor U2392 (N_2392,In_504,In_229);
xnor U2393 (N_2393,In_413,In_116);
nor U2394 (N_2394,In_95,In_190);
nor U2395 (N_2395,In_455,In_210);
nand U2396 (N_2396,In_660,In_399);
nand U2397 (N_2397,In_250,In_715);
or U2398 (N_2398,In_143,In_114);
nor U2399 (N_2399,In_121,In_487);
or U2400 (N_2400,In_107,In_42);
and U2401 (N_2401,In_537,In_677);
and U2402 (N_2402,In_340,In_222);
nand U2403 (N_2403,In_133,In_310);
nor U2404 (N_2404,In_319,In_464);
nor U2405 (N_2405,In_264,In_469);
and U2406 (N_2406,In_293,In_229);
nor U2407 (N_2407,In_309,In_268);
nor U2408 (N_2408,In_725,In_702);
nor U2409 (N_2409,In_530,In_637);
and U2410 (N_2410,In_479,In_514);
nor U2411 (N_2411,In_97,In_709);
nor U2412 (N_2412,In_44,In_208);
and U2413 (N_2413,In_724,In_649);
and U2414 (N_2414,In_298,In_473);
or U2415 (N_2415,In_632,In_468);
or U2416 (N_2416,In_161,In_524);
xor U2417 (N_2417,In_620,In_731);
nor U2418 (N_2418,In_632,In_224);
nand U2419 (N_2419,In_747,In_349);
nand U2420 (N_2420,In_137,In_370);
nor U2421 (N_2421,In_249,In_104);
and U2422 (N_2422,In_483,In_44);
and U2423 (N_2423,In_66,In_154);
nand U2424 (N_2424,In_254,In_306);
and U2425 (N_2425,In_364,In_643);
nand U2426 (N_2426,In_312,In_676);
or U2427 (N_2427,In_346,In_57);
or U2428 (N_2428,In_472,In_164);
and U2429 (N_2429,In_559,In_645);
or U2430 (N_2430,In_559,In_650);
nor U2431 (N_2431,In_314,In_549);
and U2432 (N_2432,In_725,In_679);
nand U2433 (N_2433,In_571,In_28);
nand U2434 (N_2434,In_466,In_732);
and U2435 (N_2435,In_741,In_380);
or U2436 (N_2436,In_481,In_298);
nand U2437 (N_2437,In_58,In_747);
or U2438 (N_2438,In_121,In_352);
nand U2439 (N_2439,In_327,In_293);
or U2440 (N_2440,In_48,In_237);
and U2441 (N_2441,In_349,In_389);
or U2442 (N_2442,In_65,In_453);
nor U2443 (N_2443,In_398,In_729);
nand U2444 (N_2444,In_635,In_282);
or U2445 (N_2445,In_421,In_420);
and U2446 (N_2446,In_566,In_429);
and U2447 (N_2447,In_120,In_457);
nor U2448 (N_2448,In_275,In_201);
and U2449 (N_2449,In_672,In_637);
nor U2450 (N_2450,In_641,In_455);
xor U2451 (N_2451,In_181,In_462);
xor U2452 (N_2452,In_603,In_682);
nor U2453 (N_2453,In_616,In_569);
xor U2454 (N_2454,In_392,In_123);
nand U2455 (N_2455,In_205,In_128);
and U2456 (N_2456,In_288,In_104);
and U2457 (N_2457,In_332,In_378);
nor U2458 (N_2458,In_731,In_55);
or U2459 (N_2459,In_360,In_716);
nand U2460 (N_2460,In_414,In_314);
xor U2461 (N_2461,In_298,In_491);
and U2462 (N_2462,In_89,In_632);
or U2463 (N_2463,In_673,In_536);
and U2464 (N_2464,In_516,In_289);
nand U2465 (N_2465,In_504,In_74);
and U2466 (N_2466,In_385,In_153);
nand U2467 (N_2467,In_340,In_332);
nor U2468 (N_2468,In_564,In_374);
and U2469 (N_2469,In_735,In_70);
or U2470 (N_2470,In_35,In_296);
or U2471 (N_2471,In_11,In_666);
and U2472 (N_2472,In_697,In_408);
nand U2473 (N_2473,In_711,In_516);
xor U2474 (N_2474,In_78,In_113);
nand U2475 (N_2475,In_160,In_650);
nand U2476 (N_2476,In_157,In_733);
nor U2477 (N_2477,In_302,In_563);
or U2478 (N_2478,In_65,In_410);
and U2479 (N_2479,In_64,In_217);
nand U2480 (N_2480,In_560,In_298);
nand U2481 (N_2481,In_70,In_136);
nor U2482 (N_2482,In_516,In_116);
or U2483 (N_2483,In_705,In_82);
nand U2484 (N_2484,In_664,In_743);
and U2485 (N_2485,In_353,In_660);
nand U2486 (N_2486,In_607,In_153);
nor U2487 (N_2487,In_336,In_204);
nor U2488 (N_2488,In_339,In_279);
nand U2489 (N_2489,In_228,In_552);
nor U2490 (N_2490,In_494,In_76);
nor U2491 (N_2491,In_142,In_520);
nand U2492 (N_2492,In_338,In_662);
nor U2493 (N_2493,In_189,In_237);
nor U2494 (N_2494,In_219,In_642);
nor U2495 (N_2495,In_278,In_65);
and U2496 (N_2496,In_69,In_650);
xor U2497 (N_2497,In_104,In_131);
nor U2498 (N_2498,In_533,In_330);
nor U2499 (N_2499,In_273,In_476);
nand U2500 (N_2500,N_833,N_432);
and U2501 (N_2501,N_1918,N_577);
or U2502 (N_2502,N_1031,N_441);
nand U2503 (N_2503,N_1949,N_2226);
and U2504 (N_2504,N_2110,N_1715);
and U2505 (N_2505,N_425,N_2142);
nor U2506 (N_2506,N_2041,N_1576);
nor U2507 (N_2507,N_2449,N_2338);
nor U2508 (N_2508,N_1143,N_1919);
nand U2509 (N_2509,N_1177,N_1438);
and U2510 (N_2510,N_2088,N_300);
xor U2511 (N_2511,N_24,N_1421);
nor U2512 (N_2512,N_2114,N_354);
nand U2513 (N_2513,N_662,N_1633);
or U2514 (N_2514,N_1102,N_1185);
or U2515 (N_2515,N_240,N_1056);
nor U2516 (N_2516,N_696,N_1359);
nand U2517 (N_2517,N_1904,N_244);
and U2518 (N_2518,N_1701,N_418);
or U2519 (N_2519,N_1532,N_1261);
nor U2520 (N_2520,N_508,N_1330);
nand U2521 (N_2521,N_41,N_387);
nor U2522 (N_2522,N_2308,N_1216);
nand U2523 (N_2523,N_180,N_1740);
and U2524 (N_2524,N_586,N_1725);
or U2525 (N_2525,N_827,N_1231);
or U2526 (N_2526,N_1941,N_1235);
nand U2527 (N_2527,N_414,N_1246);
nor U2528 (N_2528,N_608,N_2363);
and U2529 (N_2529,N_603,N_1938);
and U2530 (N_2530,N_841,N_73);
and U2531 (N_2531,N_1119,N_1723);
and U2532 (N_2532,N_1150,N_5);
nor U2533 (N_2533,N_1360,N_897);
nor U2534 (N_2534,N_433,N_1053);
nand U2535 (N_2535,N_1166,N_849);
nor U2536 (N_2536,N_1478,N_2062);
and U2537 (N_2537,N_1923,N_1027);
nor U2538 (N_2538,N_2214,N_1545);
and U2539 (N_2539,N_457,N_2344);
or U2540 (N_2540,N_889,N_2440);
or U2541 (N_2541,N_1688,N_338);
nand U2542 (N_2542,N_1475,N_480);
and U2543 (N_2543,N_580,N_1064);
nor U2544 (N_2544,N_237,N_2419);
nand U2545 (N_2545,N_1889,N_1305);
or U2546 (N_2546,N_26,N_1319);
nand U2547 (N_2547,N_324,N_1113);
or U2548 (N_2548,N_1340,N_2270);
nor U2549 (N_2549,N_1005,N_1417);
nand U2550 (N_2550,N_1075,N_1326);
nor U2551 (N_2551,N_1123,N_1592);
and U2552 (N_2552,N_807,N_1623);
nand U2553 (N_2553,N_2345,N_436);
and U2554 (N_2554,N_2433,N_2324);
nand U2555 (N_2555,N_1186,N_1618);
or U2556 (N_2556,N_472,N_1074);
nor U2557 (N_2557,N_405,N_1347);
nor U2558 (N_2558,N_2165,N_2339);
nor U2559 (N_2559,N_2259,N_417);
nand U2560 (N_2560,N_1101,N_628);
or U2561 (N_2561,N_953,N_1401);
nand U2562 (N_2562,N_605,N_126);
or U2563 (N_2563,N_552,N_2286);
nand U2564 (N_2564,N_1415,N_200);
xor U2565 (N_2565,N_1893,N_380);
or U2566 (N_2566,N_2395,N_14);
or U2567 (N_2567,N_1010,N_398);
and U2568 (N_2568,N_231,N_2143);
nor U2569 (N_2569,N_815,N_1995);
or U2570 (N_2570,N_1139,N_1253);
and U2571 (N_2571,N_2359,N_495);
nor U2572 (N_2572,N_805,N_2375);
xnor U2573 (N_2573,N_774,N_2067);
nand U2574 (N_2574,N_1202,N_35);
nand U2575 (N_2575,N_341,N_1787);
nand U2576 (N_2576,N_455,N_1395);
or U2577 (N_2577,N_1982,N_2163);
or U2578 (N_2578,N_664,N_1868);
or U2579 (N_2579,N_370,N_1384);
nand U2580 (N_2580,N_393,N_207);
nor U2581 (N_2581,N_1881,N_77);
or U2582 (N_2582,N_263,N_1145);
nand U2583 (N_2583,N_1513,N_199);
or U2584 (N_2584,N_1501,N_1006);
and U2585 (N_2585,N_1214,N_994);
nor U2586 (N_2586,N_1552,N_383);
or U2587 (N_2587,N_1710,N_33);
nand U2588 (N_2588,N_2046,N_1989);
nand U2589 (N_2589,N_428,N_154);
or U2590 (N_2590,N_1888,N_624);
or U2591 (N_2591,N_799,N_957);
or U2592 (N_2592,N_554,N_968);
and U2593 (N_2593,N_1537,N_363);
nor U2594 (N_2594,N_1734,N_1443);
and U2595 (N_2595,N_189,N_1639);
or U2596 (N_2596,N_1174,N_771);
and U2597 (N_2597,N_2245,N_1577);
or U2598 (N_2598,N_2306,N_101);
nor U2599 (N_2599,N_1622,N_1392);
nand U2600 (N_2600,N_828,N_738);
and U2601 (N_2601,N_185,N_2034);
nand U2602 (N_2602,N_404,N_2118);
xnor U2603 (N_2603,N_1366,N_1568);
xnor U2604 (N_2604,N_214,N_1782);
nor U2605 (N_2605,N_1199,N_1014);
nor U2606 (N_2606,N_762,N_57);
and U2607 (N_2607,N_1328,N_167);
or U2608 (N_2608,N_1329,N_699);
nand U2609 (N_2609,N_162,N_672);
nand U2610 (N_2610,N_2304,N_1135);
or U2611 (N_2611,N_923,N_2006);
nor U2612 (N_2612,N_229,N_1505);
nor U2613 (N_2613,N_1737,N_1901);
and U2614 (N_2614,N_1019,N_1018);
nor U2615 (N_2615,N_2172,N_1280);
and U2616 (N_2616,N_937,N_1062);
nor U2617 (N_2617,N_626,N_1445);
and U2618 (N_2618,N_2277,N_1132);
and U2619 (N_2619,N_1915,N_1248);
xor U2620 (N_2620,N_491,N_962);
nor U2621 (N_2621,N_2438,N_2478);
and U2622 (N_2622,N_2129,N_1706);
nand U2623 (N_2623,N_137,N_854);
and U2624 (N_2624,N_2073,N_540);
and U2625 (N_2625,N_2009,N_2146);
nor U2626 (N_2626,N_1704,N_1374);
nor U2627 (N_2627,N_122,N_1653);
nand U2628 (N_2628,N_337,N_1114);
or U2629 (N_2629,N_325,N_1283);
and U2630 (N_2630,N_881,N_2406);
nand U2631 (N_2631,N_793,N_1509);
nand U2632 (N_2632,N_2014,N_1023);
and U2633 (N_2633,N_1301,N_1449);
or U2634 (N_2634,N_1015,N_2008);
nand U2635 (N_2635,N_1255,N_1615);
or U2636 (N_2636,N_913,N_1581);
and U2637 (N_2637,N_1678,N_4);
nand U2638 (N_2638,N_1112,N_1626);
and U2639 (N_2639,N_1378,N_560);
nand U2640 (N_2640,N_1167,N_582);
nor U2641 (N_2641,N_2373,N_682);
nand U2642 (N_2642,N_70,N_1130);
nor U2643 (N_2643,N_248,N_1614);
nand U2644 (N_2644,N_2414,N_847);
nand U2645 (N_2645,N_1908,N_2038);
or U2646 (N_2646,N_637,N_2250);
nor U2647 (N_2647,N_918,N_326);
or U2648 (N_2648,N_435,N_2398);
nor U2649 (N_2649,N_242,N_1827);
and U2650 (N_2650,N_1004,N_2313);
nand U2651 (N_2651,N_2276,N_802);
nor U2652 (N_2652,N_804,N_723);
and U2653 (N_2653,N_1816,N_1555);
nor U2654 (N_2654,N_298,N_329);
nand U2655 (N_2655,N_1036,N_2403);
and U2656 (N_2656,N_0,N_1407);
or U2657 (N_2657,N_2178,N_488);
or U2658 (N_2658,N_1495,N_612);
and U2659 (N_2659,N_195,N_673);
nor U2660 (N_2660,N_2232,N_1866);
nor U2661 (N_2661,N_1299,N_212);
or U2662 (N_2662,N_744,N_43);
nor U2663 (N_2663,N_76,N_1236);
nor U2664 (N_2664,N_933,N_2124);
and U2665 (N_2665,N_950,N_2271);
nand U2666 (N_2666,N_1353,N_1646);
and U2667 (N_2667,N_765,N_427);
nand U2668 (N_2668,N_1422,N_2240);
nand U2669 (N_2669,N_44,N_2474);
or U2670 (N_2670,N_1822,N_1815);
and U2671 (N_2671,N_446,N_2097);
nand U2672 (N_2672,N_442,N_1490);
nand U2673 (N_2673,N_1621,N_296);
and U2674 (N_2674,N_1778,N_259);
nor U2675 (N_2675,N_1203,N_1464);
nor U2676 (N_2676,N_2161,N_848);
nor U2677 (N_2677,N_518,N_1791);
nor U2678 (N_2678,N_2351,N_683);
and U2679 (N_2679,N_198,N_2379);
xor U2680 (N_2680,N_1922,N_1865);
and U2681 (N_2681,N_2461,N_676);
nor U2682 (N_2682,N_753,N_2136);
or U2683 (N_2683,N_1754,N_205);
or U2684 (N_2684,N_485,N_1875);
nand U2685 (N_2685,N_392,N_1218);
and U2686 (N_2686,N_1869,N_1189);
or U2687 (N_2687,N_1672,N_2452);
and U2688 (N_2688,N_1472,N_721);
nand U2689 (N_2689,N_257,N_32);
nand U2690 (N_2690,N_1811,N_2247);
nor U2691 (N_2691,N_1819,N_315);
nor U2692 (N_2692,N_2360,N_1763);
or U2693 (N_2693,N_688,N_1320);
nand U2694 (N_2694,N_1483,N_1970);
or U2695 (N_2695,N_1675,N_1388);
nand U2696 (N_2696,N_620,N_1821);
xor U2697 (N_2697,N_1382,N_1800);
and U2698 (N_2698,N_587,N_591);
or U2699 (N_2699,N_1440,N_168);
or U2700 (N_2700,N_410,N_12);
nor U2701 (N_2701,N_1450,N_1753);
and U2702 (N_2702,N_262,N_1659);
nand U2703 (N_2703,N_264,N_1536);
and U2704 (N_2704,N_1416,N_732);
nor U2705 (N_2705,N_1589,N_117);
or U2706 (N_2706,N_1194,N_1826);
or U2707 (N_2707,N_681,N_592);
or U2708 (N_2708,N_784,N_1500);
and U2709 (N_2709,N_2399,N_1482);
and U2710 (N_2710,N_941,N_1765);
nand U2711 (N_2711,N_665,N_914);
nand U2712 (N_2712,N_1461,N_1088);
nor U2713 (N_2713,N_289,N_1147);
nand U2714 (N_2714,N_1045,N_539);
nor U2715 (N_2715,N_1958,N_1683);
and U2716 (N_2716,N_1736,N_261);
nor U2717 (N_2717,N_45,N_917);
and U2718 (N_2718,N_1029,N_1488);
nor U2719 (N_2719,N_80,N_2007);
xnor U2720 (N_2720,N_2371,N_2358);
and U2721 (N_2721,N_415,N_1894);
nor U2722 (N_2722,N_2295,N_1220);
nor U2723 (N_2723,N_423,N_707);
nor U2724 (N_2724,N_992,N_2042);
xnor U2725 (N_2725,N_2203,N_479);
nor U2726 (N_2726,N_147,N_1562);
nand U2727 (N_2727,N_1095,N_187);
nand U2728 (N_2728,N_1582,N_1724);
nor U2729 (N_2729,N_2389,N_642);
and U2730 (N_2730,N_2310,N_1466);
nor U2731 (N_2731,N_743,N_2111);
nand U2732 (N_2732,N_1476,N_1493);
nor U2733 (N_2733,N_860,N_831);
or U2734 (N_2734,N_466,N_1183);
nand U2735 (N_2735,N_820,N_787);
and U2736 (N_2736,N_2076,N_622);
and U2737 (N_2737,N_1492,N_2170);
or U2738 (N_2738,N_986,N_2130);
or U2739 (N_2739,N_362,N_2294);
nor U2740 (N_2740,N_1376,N_2187);
and U2741 (N_2741,N_775,N_1979);
or U2742 (N_2742,N_829,N_1929);
and U2743 (N_2743,N_193,N_1900);
nand U2744 (N_2744,N_1733,N_1024);
nor U2745 (N_2745,N_385,N_669);
nor U2746 (N_2746,N_912,N_2191);
nand U2747 (N_2747,N_1162,N_600);
nand U2748 (N_2748,N_865,N_317);
and U2749 (N_2749,N_2156,N_2445);
nor U2750 (N_2750,N_555,N_54);
and U2751 (N_2751,N_2018,N_852);
nand U2752 (N_2752,N_1730,N_2181);
nor U2753 (N_2753,N_999,N_2095);
xor U2754 (N_2754,N_958,N_979);
nor U2755 (N_2755,N_1825,N_1148);
nand U2756 (N_2756,N_1520,N_1987);
nor U2757 (N_2757,N_1959,N_282);
nand U2758 (N_2758,N_2213,N_184);
or U2759 (N_2759,N_909,N_211);
or U2760 (N_2760,N_1354,N_733);
nor U2761 (N_2761,N_1161,N_1560);
or U2762 (N_2762,N_1664,N_2390);
nor U2763 (N_2763,N_638,N_2257);
and U2764 (N_2764,N_2031,N_2053);
nand U2765 (N_2765,N_1665,N_408);
nand U2766 (N_2766,N_2196,N_389);
and U2767 (N_2767,N_617,N_1057);
nor U2768 (N_2768,N_140,N_1504);
nor U2769 (N_2769,N_894,N_1686);
nor U2770 (N_2770,N_2349,N_120);
or U2771 (N_2771,N_2139,N_1097);
nor U2772 (N_2772,N_996,N_2422);
nor U2773 (N_2773,N_1533,N_1210);
or U2774 (N_2774,N_2140,N_1546);
nand U2775 (N_2775,N_1418,N_2356);
xnor U2776 (N_2776,N_78,N_112);
nand U2777 (N_2777,N_2497,N_1641);
nor U2778 (N_2778,N_2332,N_1300);
xnor U2779 (N_2779,N_520,N_110);
or U2780 (N_2780,N_987,N_928);
nor U2781 (N_2781,N_2446,N_704);
nor U2782 (N_2782,N_2437,N_1289);
xor U2783 (N_2783,N_2137,N_401);
or U2784 (N_2784,N_218,N_1327);
or U2785 (N_2785,N_1502,N_1403);
nand U2786 (N_2786,N_1506,N_481);
or U2787 (N_2787,N_834,N_2283);
or U2788 (N_2788,N_794,N_1510);
nand U2789 (N_2789,N_2377,N_977);
nor U2790 (N_2790,N_1830,N_2138);
nor U2791 (N_2791,N_1732,N_1975);
and U2792 (N_2792,N_1670,N_946);
or U2793 (N_2793,N_92,N_1850);
or U2794 (N_2794,N_50,N_100);
nand U2795 (N_2795,N_2391,N_2158);
nor U2796 (N_2796,N_2085,N_340);
or U2797 (N_2797,N_424,N_2296);
nand U2798 (N_2798,N_9,N_1717);
nor U2799 (N_2799,N_716,N_471);
nand U2800 (N_2800,N_1042,N_585);
nand U2801 (N_2801,N_2231,N_1292);
or U2802 (N_2802,N_1335,N_56);
nor U2803 (N_2803,N_208,N_692);
or U2804 (N_2804,N_421,N_376);
and U2805 (N_2805,N_1334,N_1441);
or U2806 (N_2806,N_1087,N_1566);
or U2807 (N_2807,N_1258,N_190);
nand U2808 (N_2808,N_1558,N_2325);
nand U2809 (N_2809,N_702,N_1981);
nor U2810 (N_2810,N_2092,N_619);
nor U2811 (N_2811,N_219,N_504);
nor U2812 (N_2812,N_1703,N_983);
nor U2813 (N_2813,N_2151,N_1991);
nor U2814 (N_2814,N_1976,N_1612);
nand U2815 (N_2815,N_2328,N_1195);
nand U2816 (N_2816,N_1585,N_407);
and U2817 (N_2817,N_443,N_1092);
nor U2818 (N_2818,N_97,N_23);
xnor U2819 (N_2819,N_356,N_2262);
and U2820 (N_2820,N_1914,N_49);
xor U2821 (N_2821,N_935,N_1063);
nand U2822 (N_2822,N_973,N_1078);
or U2823 (N_2823,N_1316,N_514);
nor U2824 (N_2824,N_227,N_2320);
nor U2825 (N_2825,N_995,N_1857);
and U2826 (N_2826,N_1898,N_2431);
and U2827 (N_2827,N_2427,N_1487);
nor U2828 (N_2828,N_1312,N_339);
or U2829 (N_2829,N_386,N_1314);
nor U2830 (N_2830,N_932,N_1902);
nand U2831 (N_2831,N_579,N_1992);
or U2832 (N_2832,N_419,N_192);
nor U2833 (N_2833,N_236,N_2468);
and U2834 (N_2834,N_675,N_292);
and U2835 (N_2835,N_754,N_879);
and U2836 (N_2836,N_647,N_291);
or U2837 (N_2837,N_29,N_867);
nand U2838 (N_2838,N_258,N_1735);
and U2839 (N_2839,N_2496,N_400);
and U2840 (N_2840,N_1645,N_234);
or U2841 (N_2841,N_1424,N_1636);
and U2842 (N_2842,N_2123,N_1133);
and U2843 (N_2843,N_569,N_141);
or U2844 (N_2844,N_1067,N_213);
or U2845 (N_2845,N_492,N_1597);
or U2846 (N_2846,N_1679,N_1554);
and U2847 (N_2847,N_630,N_1887);
and U2848 (N_2848,N_1109,N_715);
and U2849 (N_2849,N_1116,N_1932);
nand U2850 (N_2850,N_279,N_1468);
nand U2851 (N_2851,N_1808,N_1484);
and U2852 (N_2852,N_1267,N_143);
xnor U2853 (N_2853,N_2413,N_2162);
nor U2854 (N_2854,N_1640,N_2026);
or U2855 (N_2855,N_1001,N_2418);
or U2856 (N_2856,N_368,N_693);
nor U2857 (N_2857,N_1906,N_304);
or U2858 (N_2858,N_2204,N_2400);
or U2859 (N_2859,N_561,N_961);
or U2860 (N_2860,N_1948,N_186);
and U2861 (N_2861,N_1529,N_2166);
nor U2862 (N_2862,N_2303,N_1051);
xnor U2863 (N_2863,N_1567,N_985);
or U2864 (N_2864,N_748,N_2269);
and U2865 (N_2865,N_1911,N_1310);
nor U2866 (N_2866,N_1243,N_1954);
or U2867 (N_2867,N_2301,N_2116);
nand U2868 (N_2868,N_1530,N_1883);
nor U2869 (N_2869,N_1408,N_2244);
or U2870 (N_2870,N_808,N_2267);
nand U2871 (N_2871,N_371,N_604);
nor U2872 (N_2872,N_863,N_1459);
nor U2873 (N_2873,N_155,N_1322);
and U2874 (N_2874,N_366,N_1897);
nand U2875 (N_2875,N_2321,N_907);
or U2876 (N_2876,N_1870,N_249);
nor U2877 (N_2877,N_1100,N_374);
nand U2878 (N_2878,N_2049,N_836);
and U2879 (N_2879,N_66,N_1265);
or U2880 (N_2880,N_171,N_967);
xnor U2881 (N_2881,N_67,N_108);
nand U2882 (N_2882,N_293,N_1007);
or U2883 (N_2883,N_225,N_2155);
nor U2884 (N_2884,N_671,N_1939);
nand U2885 (N_2885,N_1663,N_1249);
nor U2886 (N_2886,N_247,N_360);
and U2887 (N_2887,N_1175,N_690);
and U2888 (N_2888,N_749,N_667);
nor U2889 (N_2889,N_874,N_2224);
nor U2890 (N_2890,N_2243,N_335);
and U2891 (N_2891,N_2274,N_1351);
nor U2892 (N_2892,N_1792,N_220);
and U2893 (N_2893,N_938,N_873);
and U2894 (N_2894,N_1598,N_1447);
or U2895 (N_2895,N_294,N_1543);
and U2896 (N_2896,N_997,N_825);
and U2897 (N_2897,N_1593,N_1785);
or U2898 (N_2898,N_1985,N_840);
nand U2899 (N_2899,N_886,N_1499);
or U2900 (N_2900,N_157,N_1234);
xor U2901 (N_2901,N_437,N_1867);
nor U2902 (N_2902,N_2479,N_87);
nand U2903 (N_2903,N_269,N_2424);
nor U2904 (N_2904,N_1059,N_188);
nor U2905 (N_2905,N_2218,N_1239);
and U2906 (N_2906,N_776,N_2189);
and U2907 (N_2907,N_2252,N_2086);
or U2908 (N_2908,N_1016,N_1874);
nor U2909 (N_2909,N_1245,N_550);
nor U2910 (N_2910,N_1783,N_1674);
or U2911 (N_2911,N_2012,N_618);
nor U2912 (N_2912,N_382,N_332);
nor U2913 (N_2913,N_1049,N_691);
nor U2914 (N_2914,N_884,N_125);
or U2915 (N_2915,N_698,N_929);
nand U2916 (N_2916,N_159,N_1169);
and U2917 (N_2917,N_1193,N_870);
or U2918 (N_2918,N_616,N_1070);
xor U2919 (N_2919,N_1437,N_355);
and U2920 (N_2920,N_1349,N_1226);
nor U2921 (N_2921,N_2337,N_1719);
and U2922 (N_2922,N_982,N_1012);
nor U2923 (N_2923,N_516,N_1047);
nor U2924 (N_2924,N_1190,N_1660);
nand U2925 (N_2925,N_150,N_1458);
and U2926 (N_2926,N_1494,N_1507);
or U2927 (N_2927,N_1017,N_486);
and U2928 (N_2928,N_2251,N_921);
or U2929 (N_2929,N_1629,N_562);
and U2930 (N_2930,N_1456,N_135);
or U2931 (N_2931,N_1756,N_2392);
and U2932 (N_2932,N_742,N_1750);
or U2933 (N_2933,N_2429,N_2037);
nand U2934 (N_2934,N_811,N_2182);
and U2935 (N_2935,N_1578,N_713);
and U2936 (N_2936,N_146,N_1396);
nor U2937 (N_2937,N_648,N_2347);
nor U2938 (N_2938,N_2011,N_763);
or U2939 (N_2939,N_1117,N_148);
xnor U2940 (N_2940,N_1933,N_1470);
nand U2941 (N_2941,N_902,N_2381);
and U2942 (N_2942,N_451,N_2176);
and U2943 (N_2943,N_2383,N_2368);
or U2944 (N_2944,N_2365,N_2005);
and U2945 (N_2945,N_328,N_53);
nor U2946 (N_2946,N_1721,N_464);
or U2947 (N_2947,N_278,N_2300);
nand U2948 (N_2948,N_2125,N_1096);
and U2949 (N_2949,N_1638,N_1572);
or U2950 (N_2950,N_2293,N_936);
and U2951 (N_2951,N_1515,N_658);
nor U2952 (N_2952,N_972,N_2463);
or U2953 (N_2953,N_2167,N_459);
nand U2954 (N_2954,N_351,N_955);
nand U2955 (N_2955,N_2070,N_1390);
nor U2956 (N_2956,N_1630,N_46);
nand U2957 (N_2957,N_1687,N_2415);
and U2958 (N_2958,N_1535,N_1068);
nand U2959 (N_2959,N_1768,N_1091);
nor U2960 (N_2960,N_2402,N_1757);
and U2961 (N_2961,N_581,N_2117);
and U2962 (N_2962,N_2367,N_718);
and U2963 (N_2963,N_2179,N_51);
nor U2964 (N_2964,N_226,N_1903);
nor U2965 (N_2965,N_2355,N_260);
nor U2966 (N_2966,N_571,N_1571);
nor U2967 (N_2967,N_1988,N_473);
nand U2968 (N_2968,N_989,N_779);
and U2969 (N_2969,N_2099,N_318);
and U2970 (N_2970,N_1164,N_1676);
nor U2971 (N_2971,N_1843,N_79);
and U2972 (N_2972,N_963,N_1159);
and U2973 (N_2973,N_359,N_89);
or U2974 (N_2974,N_2152,N_510);
or U2975 (N_2975,N_172,N_196);
and U2976 (N_2976,N_13,N_156);
nor U2977 (N_2977,N_2239,N_1285);
and U2978 (N_2978,N_270,N_1854);
nand U2979 (N_2979,N_2255,N_2412);
nor U2980 (N_2980,N_1368,N_589);
nand U2981 (N_2981,N_1350,N_2369);
nand U2982 (N_2982,N_1372,N_2104);
or U2983 (N_2983,N_1973,N_1943);
and U2984 (N_2984,N_1370,N_1471);
or U2985 (N_2985,N_641,N_1153);
nand U2986 (N_2986,N_1188,N_1624);
and U2987 (N_2987,N_1498,N_2004);
or U2988 (N_2988,N_310,N_1256);
nand U2989 (N_2989,N_489,N_1779);
nand U2990 (N_2990,N_1748,N_1853);
nand U2991 (N_2991,N_1474,N_1156);
nor U2992 (N_2992,N_2148,N_319);
or U2993 (N_2993,N_1178,N_151);
nor U2994 (N_2994,N_11,N_511);
xor U2995 (N_2995,N_2335,N_1357);
or U2996 (N_2996,N_243,N_1294);
and U2997 (N_2997,N_712,N_2173);
nor U2998 (N_2998,N_2183,N_1090);
nand U2999 (N_2999,N_643,N_2205);
and U3000 (N_3000,N_1616,N_1950);
nor U3001 (N_3001,N_2185,N_1890);
nor U3002 (N_3002,N_1878,N_202);
and U3003 (N_3003,N_1619,N_524);
or U3004 (N_3004,N_575,N_856);
nor U3005 (N_3005,N_36,N_1521);
or U3006 (N_3006,N_1601,N_557);
or U3007 (N_3007,N_719,N_644);
and U3008 (N_3008,N_131,N_1344);
and U3009 (N_3009,N_2043,N_649);
nand U3010 (N_3010,N_2253,N_559);
nor U3011 (N_3011,N_839,N_1647);
nor U3012 (N_3012,N_1298,N_2171);
nand U3013 (N_3013,N_2451,N_1877);
and U3014 (N_3014,N_1526,N_657);
nand U3015 (N_3015,N_88,N_574);
nand U3016 (N_3016,N_2459,N_568);
and U3017 (N_3017,N_2444,N_646);
nor U3018 (N_3018,N_611,N_1606);
nor U3019 (N_3019,N_872,N_2198);
and U3020 (N_3020,N_183,N_2471);
nor U3021 (N_3021,N_951,N_505);
and U3022 (N_3022,N_850,N_1760);
or U3023 (N_3023,N_517,N_594);
or U3024 (N_3024,N_1317,N_1104);
or U3025 (N_3025,N_1935,N_535);
and U3026 (N_3026,N_1293,N_851);
and U3027 (N_3027,N_2200,N_2264);
and U3028 (N_3028,N_1594,N_2397);
nand U3029 (N_3029,N_221,N_888);
nor U3030 (N_3030,N_1844,N_1885);
or U3031 (N_3031,N_880,N_727);
nor U3032 (N_3032,N_751,N_636);
or U3033 (N_3033,N_832,N_496);
and U3034 (N_3034,N_2287,N_1439);
nor U3035 (N_3035,N_1741,N_1040);
or U3036 (N_3036,N_966,N_869);
nor U3037 (N_3037,N_1654,N_2302);
nor U3038 (N_3038,N_2222,N_531);
xnor U3039 (N_3039,N_2485,N_2030);
nand U3040 (N_3040,N_2003,N_2473);
and U3041 (N_3041,N_1121,N_1182);
or U3042 (N_3042,N_891,N_119);
and U3043 (N_3043,N_1237,N_1946);
nor U3044 (N_3044,N_1849,N_1085);
nor U3045 (N_3045,N_2021,N_2020);
nor U3046 (N_3046,N_81,N_2455);
and U3047 (N_3047,N_770,N_1518);
nand U3048 (N_3048,N_730,N_1824);
and U3049 (N_3049,N_2372,N_121);
or U3050 (N_3050,N_527,N_1165);
nand U3051 (N_3051,N_1163,N_634);
and U3052 (N_3052,N_1544,N_2001);
or U3053 (N_3053,N_1512,N_2462);
nor U3054 (N_3054,N_1176,N_1747);
nor U3055 (N_3055,N_275,N_507);
nand U3056 (N_3056,N_2387,N_309);
and U3057 (N_3057,N_1355,N_281);
and U3058 (N_3058,N_1602,N_1207);
nor U3059 (N_3059,N_551,N_1684);
nand U3060 (N_3060,N_1556,N_1848);
or U3061 (N_3061,N_483,N_674);
or U3062 (N_3062,N_1196,N_1642);
and U3063 (N_3063,N_1009,N_1680);
and U3064 (N_3064,N_588,N_1297);
nand U3065 (N_3065,N_1081,N_1131);
and U3066 (N_3066,N_817,N_2280);
nand U3067 (N_3067,N_2442,N_175);
nor U3068 (N_3068,N_1477,N_1157);
xnor U3069 (N_3069,N_1043,N_1151);
and U3070 (N_3070,N_785,N_885);
nor U3071 (N_3071,N_327,N_714);
and U3072 (N_3072,N_548,N_526);
nand U3073 (N_3073,N_752,N_1467);
and U3074 (N_3074,N_164,N_1324);
nand U3075 (N_3075,N_2498,N_203);
xor U3076 (N_3076,N_2164,N_1599);
or U3077 (N_3077,N_892,N_1172);
nand U3078 (N_3078,N_2350,N_1393);
and U3079 (N_3079,N_871,N_2352);
nor U3080 (N_3080,N_656,N_1802);
nor U3081 (N_3081,N_903,N_1230);
nand U3082 (N_3082,N_2401,N_160);
nor U3083 (N_3083,N_474,N_843);
nand U3084 (N_3084,N_632,N_959);
or U3085 (N_3085,N_308,N_2260);
or U3086 (N_3086,N_1160,N_499);
or U3087 (N_3087,N_769,N_1356);
and U3088 (N_3088,N_449,N_1406);
and U3089 (N_3089,N_1035,N_1548);
nand U3090 (N_3090,N_1069,N_1726);
or U3091 (N_3091,N_1251,N_1561);
nor U3092 (N_3092,N_2202,N_942);
or U3093 (N_3093,N_980,N_118);
nand U3094 (N_3094,N_2386,N_1270);
xnor U3095 (N_3095,N_1540,N_1702);
nand U3096 (N_3096,N_246,N_1266);
or U3097 (N_3097,N_197,N_532);
or U3098 (N_3098,N_1124,N_924);
and U3099 (N_3099,N_2336,N_1118);
nor U3100 (N_3100,N_1046,N_1978);
and U3101 (N_3101,N_2194,N_1609);
and U3102 (N_3102,N_1457,N_1517);
and U3103 (N_3103,N_697,N_2329);
xnor U3104 (N_3104,N_2481,N_1997);
nor U3105 (N_3105,N_1588,N_2160);
nor U3106 (N_3106,N_1428,N_1662);
and U3107 (N_3107,N_467,N_2382);
and U3108 (N_3108,N_1241,N_663);
and U3109 (N_3109,N_2314,N_1940);
nor U3110 (N_3110,N_1586,N_823);
and U3111 (N_3111,N_750,N_361);
or U3112 (N_3112,N_679,N_1259);
nand U3113 (N_3113,N_2077,N_1228);
and U3114 (N_3114,N_2331,N_1971);
or U3115 (N_3115,N_576,N_469);
or U3116 (N_3116,N_1667,N_709);
nand U3117 (N_3117,N_1793,N_27);
nand U3118 (N_3118,N_1311,N_2047);
nand U3119 (N_3119,N_717,N_130);
or U3120 (N_3120,N_1436,N_678);
or U3121 (N_3121,N_1994,N_2483);
xor U3122 (N_3122,N_1569,N_1489);
and U3123 (N_3123,N_1631,N_494);
or U3124 (N_3124,N_2154,N_1491);
and U3125 (N_3125,N_822,N_2119);
xor U3126 (N_3126,N_1072,N_629);
nand U3127 (N_3127,N_21,N_1211);
nand U3128 (N_3128,N_63,N_174);
nand U3129 (N_3129,N_245,N_2268);
xor U3130 (N_3130,N_659,N_345);
and U3131 (N_3131,N_2206,N_1539);
nor U3132 (N_3132,N_1306,N_1998);
nor U3133 (N_3133,N_1739,N_990);
xnor U3134 (N_3134,N_344,N_689);
or U3135 (N_3135,N_558,N_1838);
or U3136 (N_3136,N_170,N_1879);
nand U3137 (N_3137,N_2195,N_2404);
nand U3138 (N_3138,N_635,N_91);
nand U3139 (N_3139,N_460,N_900);
nand U3140 (N_3140,N_145,N_2217);
nand U3141 (N_3141,N_687,N_757);
nand U3142 (N_3142,N_971,N_745);
and U3143 (N_3143,N_654,N_2258);
or U3144 (N_3144,N_2212,N_268);
nor U3145 (N_3145,N_1648,N_1872);
nor U3146 (N_3146,N_2450,N_1691);
nor U3147 (N_3147,N_487,N_1690);
nor U3148 (N_3148,N_2149,N_2177);
nor U3149 (N_3149,N_1103,N_2134);
or U3150 (N_3150,N_1925,N_1446);
and U3151 (N_3151,N_2054,N_1524);
or U3152 (N_3152,N_2109,N_2211);
and U3153 (N_3153,N_2475,N_911);
nor U3154 (N_3154,N_567,N_1144);
and U3155 (N_3155,N_1965,N_2333);
nand U3156 (N_3156,N_2279,N_391);
nor U3157 (N_3157,N_969,N_1570);
or U3158 (N_3158,N_1880,N_1275);
and U3159 (N_3159,N_2411,N_2228);
nand U3160 (N_3160,N_232,N_2343);
nand U3161 (N_3161,N_1080,N_1011);
nor U3162 (N_3162,N_1341,N_1731);
and U3163 (N_3163,N_395,N_149);
nand U3164 (N_3164,N_1434,N_1308);
nor U3165 (N_3165,N_974,N_926);
nand U3166 (N_3166,N_1079,N_1442);
xnor U3167 (N_3167,N_1700,N_1969);
and U3168 (N_3168,N_1181,N_798);
or U3169 (N_3169,N_173,N_365);
or U3170 (N_3170,N_47,N_1279);
and U3171 (N_3171,N_1528,N_2064);
nor U3172 (N_3172,N_1385,N_639);
and U3173 (N_3173,N_2288,N_1140);
and U3174 (N_3174,N_1632,N_529);
or U3175 (N_3175,N_297,N_916);
nor U3176 (N_3176,N_2416,N_2408);
nor U3177 (N_3177,N_2290,N_1806);
and U3178 (N_3178,N_2417,N_975);
and U3179 (N_3179,N_2108,N_2223);
or U3180 (N_3180,N_2495,N_2421);
nand U3181 (N_3181,N_93,N_1752);
nor U3182 (N_3182,N_2102,N_1373);
and U3183 (N_3183,N_803,N_311);
nor U3184 (N_3184,N_1432,N_375);
nand U3185 (N_3185,N_1227,N_1371);
or U3186 (N_3186,N_590,N_1224);
nand U3187 (N_3187,N_1751,N_768);
nor U3188 (N_3188,N_103,N_224);
and U3189 (N_3189,N_99,N_302);
or U3190 (N_3190,N_343,N_2311);
or U3191 (N_3191,N_2215,N_19);
and U3192 (N_3192,N_1876,N_2029);
or U3193 (N_3193,N_2454,N_1831);
nand U3194 (N_3194,N_1564,N_1673);
nand U3195 (N_3195,N_1420,N_1604);
nand U3196 (N_3196,N_465,N_2281);
nor U3197 (N_3197,N_1644,N_583);
nor U3198 (N_3198,N_816,N_1921);
nand U3199 (N_3199,N_2096,N_161);
and U3200 (N_3200,N_388,N_1770);
nor U3201 (N_3201,N_1907,N_336);
nand U3202 (N_3202,N_280,N_706);
and U3203 (N_3203,N_323,N_792);
or U3204 (N_3204,N_1774,N_1204);
or U3205 (N_3205,N_2299,N_1862);
and U3206 (N_3206,N_2000,N_1397);
or U3207 (N_3207,N_2225,N_700);
or U3208 (N_3208,N_837,N_2208);
or U3209 (N_3209,N_812,N_1771);
nand U3210 (N_3210,N_1219,N_2405);
xnor U3211 (N_3211,N_1899,N_255);
nor U3212 (N_3212,N_1711,N_1242);
and U3213 (N_3213,N_857,N_3);
nor U3214 (N_3214,N_1534,N_1262);
nor U3215 (N_3215,N_233,N_940);
xnor U3216 (N_3216,N_153,N_2131);
nor U3217 (N_3217,N_1232,N_1583);
nor U3218 (N_3218,N_2128,N_906);
nor U3219 (N_3219,N_1342,N_740);
nand U3220 (N_3220,N_2059,N_1346);
or U3221 (N_3221,N_1728,N_1990);
and U3222 (N_3222,N_1859,N_1620);
nor U3223 (N_3223,N_650,N_515);
nor U3224 (N_3224,N_728,N_927);
nor U3225 (N_3225,N_2219,N_684);
nand U3226 (N_3226,N_1677,N_572);
or U3227 (N_3227,N_1759,N_1722);
nor U3228 (N_3228,N_2127,N_411);
nor U3229 (N_3229,N_305,N_2089);
and U3230 (N_3230,N_1519,N_1086);
nor U3231 (N_3231,N_2052,N_2426);
or U3232 (N_3232,N_1149,N_1769);
and U3233 (N_3233,N_222,N_283);
and U3234 (N_3234,N_2227,N_152);
nand U3235 (N_3235,N_2458,N_444);
nand U3236 (N_3236,N_40,N_85);
or U3237 (N_3237,N_439,N_2248);
and U3238 (N_3238,N_796,N_2435);
and U3239 (N_3239,N_842,N_905);
nor U3240 (N_3240,N_1836,N_1026);
and U3241 (N_3241,N_1025,N_2348);
or U3242 (N_3242,N_2282,N_901);
or U3243 (N_3243,N_2361,N_2068);
or U3244 (N_3244,N_1864,N_1563);
nor U3245 (N_3245,N_1835,N_312);
or U3246 (N_3246,N_1637,N_342);
or U3247 (N_3247,N_1916,N_177);
and U3248 (N_3248,N_625,N_2436);
xnor U3249 (N_3249,N_875,N_685);
nand U3250 (N_3250,N_1276,N_2060);
nor U3251 (N_3251,N_855,N_179);
or U3252 (N_3252,N_286,N_2035);
or U3253 (N_3253,N_1054,N_2157);
and U3254 (N_3254,N_976,N_1720);
nand U3255 (N_3255,N_633,N_2056);
nor U3256 (N_3256,N_194,N_2315);
nand U3257 (N_3257,N_1331,N_2488);
and U3258 (N_3258,N_373,N_2341);
and U3259 (N_3259,N_1953,N_2023);
or U3260 (N_3260,N_1184,N_72);
nor U3261 (N_3261,N_1089,N_1380);
nand U3262 (N_3262,N_2153,N_978);
nand U3263 (N_3263,N_1309,N_2083);
or U3264 (N_3264,N_1465,N_537);
or U3265 (N_3265,N_737,N_655);
and U3266 (N_3266,N_1538,N_1961);
nand U3267 (N_3267,N_2316,N_2476);
or U3268 (N_3268,N_610,N_1000);
and U3269 (N_3269,N_578,N_1668);
nor U3270 (N_3270,N_523,N_2027);
or U3271 (N_3271,N_2045,N_1213);
or U3272 (N_3272,N_2234,N_69);
and U3273 (N_3273,N_1021,N_1200);
xor U3274 (N_3274,N_313,N_1398);
nor U3275 (N_3275,N_1650,N_447);
and U3276 (N_3276,N_991,N_725);
nor U3277 (N_3277,N_2327,N_1240);
nor U3278 (N_3278,N_2032,N_1749);
nor U3279 (N_3279,N_2121,N_1238);
and U3280 (N_3280,N_2482,N_1332);
or U3281 (N_3281,N_1960,N_1073);
nor U3282 (N_3282,N_1926,N_954);
and U3283 (N_3283,N_1972,N_1093);
or U3284 (N_3284,N_2309,N_124);
and U3285 (N_3285,N_8,N_898);
or U3286 (N_3286,N_1810,N_2180);
nand U3287 (N_3287,N_1410,N_238);
or U3288 (N_3288,N_627,N_169);
and U3289 (N_3289,N_939,N_1127);
nand U3290 (N_3290,N_2342,N_1847);
or U3291 (N_3291,N_1858,N_2122);
nor U3292 (N_3292,N_1128,N_204);
or U3293 (N_3293,N_1288,N_61);
and U3294 (N_3294,N_191,N_397);
xnor U3295 (N_3295,N_2216,N_652);
or U3296 (N_3296,N_1745,N_2469);
nor U3297 (N_3297,N_1233,N_1111);
xor U3298 (N_3298,N_1550,N_868);
nand U3299 (N_3299,N_756,N_1264);
and U3300 (N_3300,N_1574,N_2254);
or U3301 (N_3301,N_458,N_573);
nor U3302 (N_3302,N_107,N_1391);
and U3303 (N_3303,N_1812,N_1217);
nor U3304 (N_3304,N_949,N_2112);
nand U3305 (N_3305,N_1281,N_1799);
nand U3306 (N_3306,N_6,N_15);
and U3307 (N_3307,N_859,N_1379);
or U3308 (N_3308,N_2144,N_1861);
nand U3309 (N_3309,N_536,N_878);
and U3310 (N_3310,N_2192,N_2285);
and U3311 (N_3311,N_1685,N_862);
and U3312 (N_3312,N_1977,N_813);
and U3313 (N_3313,N_1784,N_493);
nor U3314 (N_3314,N_2420,N_142);
and U3315 (N_3315,N_31,N_1419);
nor U3316 (N_3316,N_1315,N_2428);
and U3317 (N_3317,N_2233,N_506);
nand U3318 (N_3318,N_1910,N_1986);
nor U3319 (N_3319,N_34,N_253);
and U3320 (N_3320,N_2188,N_1789);
or U3321 (N_3321,N_440,N_773);
and U3322 (N_3322,N_1453,N_1773);
nor U3323 (N_3323,N_394,N_2249);
nand U3324 (N_3324,N_2492,N_1579);
nand U3325 (N_3325,N_601,N_948);
nor U3326 (N_3326,N_448,N_1573);
and U3327 (N_3327,N_216,N_25);
nand U3328 (N_3328,N_1364,N_734);
or U3329 (N_3329,N_37,N_1833);
and U3330 (N_3330,N_1775,N_2175);
nor U3331 (N_3331,N_1587,N_104);
nor U3332 (N_3332,N_1302,N_1171);
nand U3333 (N_3333,N_2493,N_1338);
or U3334 (N_3334,N_1425,N_1129);
nor U3335 (N_3335,N_838,N_1947);
and U3336 (N_3336,N_115,N_1649);
xor U3337 (N_3337,N_500,N_1523);
and U3338 (N_3338,N_502,N_920);
or U3339 (N_3339,N_2298,N_2477);
or U3340 (N_3340,N_1274,N_82);
nand U3341 (N_3341,N_1605,N_853);
or U3342 (N_3342,N_307,N_90);
nor U3343 (N_3343,N_116,N_1206);
nor U3344 (N_3344,N_75,N_1048);
nand U3345 (N_3345,N_1738,N_686);
and U3346 (N_3346,N_970,N_1435);
and U3347 (N_3347,N_2241,N_429);
or U3348 (N_3348,N_1108,N_2312);
nand U3349 (N_3349,N_945,N_2448);
or U3350 (N_3350,N_522,N_1852);
and U3351 (N_3351,N_1634,N_1282);
nand U3352 (N_3352,N_252,N_454);
nand U3353 (N_3353,N_1595,N_1804);
and U3354 (N_3354,N_1361,N_1020);
nand U3355 (N_3355,N_2201,N_1596);
nand U3356 (N_3356,N_1823,N_521);
nand U3357 (N_3357,N_1936,N_2061);
nand U3358 (N_3358,N_1993,N_1856);
or U3359 (N_3359,N_138,N_651);
nand U3360 (N_3360,N_1607,N_136);
nor U3361 (N_3361,N_1244,N_1610);
or U3362 (N_3362,N_1818,N_1999);
and U3363 (N_3363,N_887,N_2013);
nand U3364 (N_3364,N_1625,N_1041);
and U3365 (N_3365,N_2305,N_2385);
nand U3366 (N_3366,N_206,N_1473);
and U3367 (N_3367,N_1661,N_127);
nand U3368 (N_3368,N_1912,N_1170);
or U3369 (N_3369,N_2396,N_95);
nor U3370 (N_3370,N_1790,N_1920);
nand U3371 (N_3371,N_2297,N_1400);
nand U3372 (N_3372,N_2484,N_1411);
nand U3373 (N_3373,N_2346,N_1404);
and U3374 (N_3374,N_530,N_2150);
or U3375 (N_3375,N_2058,N_528);
and U3376 (N_3376,N_2425,N_1152);
xnor U3377 (N_3377,N_1627,N_1713);
nand U3378 (N_3378,N_295,N_846);
or U3379 (N_3379,N_1796,N_68);
and U3380 (N_3380,N_767,N_759);
nor U3381 (N_3381,N_334,N_736);
or U3382 (N_3382,N_695,N_1952);
nand U3383 (N_3383,N_1817,N_789);
nand U3384 (N_3384,N_710,N_2120);
nor U3385 (N_3385,N_1065,N_181);
or U3386 (N_3386,N_1762,N_1996);
or U3387 (N_3387,N_1693,N_484);
nor U3388 (N_3388,N_1909,N_1692);
and U3389 (N_3389,N_1273,N_2322);
nor U3390 (N_3390,N_998,N_201);
and U3391 (N_3391,N_965,N_1221);
or U3392 (N_3392,N_1137,N_988);
or U3393 (N_3393,N_2221,N_809);
nand U3394 (N_3394,N_2050,N_549);
nor U3395 (N_3395,N_1758,N_1486);
or U3396 (N_3396,N_755,N_821);
and U3397 (N_3397,N_547,N_1032);
nor U3398 (N_3398,N_694,N_2048);
nand U3399 (N_3399,N_128,N_801);
and U3400 (N_3400,N_1788,N_1173);
nor U3401 (N_3401,N_726,N_1076);
nand U3402 (N_3402,N_1377,N_1252);
nand U3403 (N_3403,N_2407,N_1481);
nand U3404 (N_3404,N_1260,N_780);
or U3405 (N_3405,N_276,N_2106);
nor U3406 (N_3406,N_2272,N_1503);
or U3407 (N_3407,N_2364,N_1682);
or U3408 (N_3408,N_1828,N_2275);
or U3409 (N_3409,N_38,N_2499);
nor U3410 (N_3410,N_2487,N_2284);
nand U3411 (N_3411,N_1860,N_1776);
and U3412 (N_3412,N_330,N_1272);
nand U3413 (N_3413,N_254,N_2066);
nand U3414 (N_3414,N_1485,N_1613);
nor U3415 (N_3415,N_1575,N_1541);
or U3416 (N_3416,N_2237,N_288);
and U3417 (N_3417,N_956,N_1321);
or U3418 (N_3418,N_593,N_503);
nand U3419 (N_3419,N_2145,N_919);
nor U3420 (N_3420,N_1122,N_2340);
or U3421 (N_3421,N_1383,N_2098);
nand U3422 (N_3422,N_1115,N_2105);
nor U3423 (N_3423,N_2370,N_84);
and U3424 (N_3424,N_731,N_158);
nor U3425 (N_3425,N_2209,N_2236);
nand U3426 (N_3426,N_1944,N_2199);
or U3427 (N_3427,N_645,N_1761);
nand U3428 (N_3428,N_1451,N_2380);
nor U3429 (N_3429,N_764,N_384);
nor U3430 (N_3430,N_538,N_595);
or U3431 (N_3431,N_1657,N_1336);
nor U3432 (N_3432,N_2318,N_501);
or U3433 (N_3433,N_1358,N_452);
and U3434 (N_3434,N_861,N_1697);
or U3435 (N_3435,N_1786,N_797);
nand U3436 (N_3436,N_1497,N_563);
nor U3437 (N_3437,N_1277,N_277);
nand U3438 (N_3438,N_893,N_2135);
and U3439 (N_3439,N_735,N_71);
or U3440 (N_3440,N_2063,N_2242);
or U3441 (N_3441,N_2393,N_790);
xor U3442 (N_3442,N_456,N_470);
nor U3443 (N_3443,N_1873,N_1966);
and U3444 (N_3444,N_925,N_1448);
nand U3445 (N_3445,N_2081,N_981);
and U3446 (N_3446,N_1766,N_17);
or U3447 (N_3447,N_1142,N_1930);
nand U3448 (N_3448,N_2044,N_2366);
nor U3449 (N_3449,N_2423,N_703);
nand U3450 (N_3450,N_1527,N_1008);
or U3451 (N_3451,N_810,N_413);
nor U3452 (N_3452,N_1967,N_102);
nor U3453 (N_3453,N_65,N_299);
or U3454 (N_3454,N_1136,N_597);
nand U3455 (N_3455,N_320,N_422);
and U3456 (N_3456,N_2019,N_934);
or U3457 (N_3457,N_1842,N_348);
and U3458 (N_3458,N_2480,N_1839);
or U3459 (N_3459,N_2,N_2133);
xnor U3460 (N_3460,N_1807,N_30);
nor U3461 (N_3461,N_2017,N_1205);
nor U3462 (N_3462,N_1974,N_7);
and U3463 (N_3463,N_2388,N_896);
nand U3464 (N_3464,N_1855,N_1600);
or U3465 (N_3465,N_1522,N_1060);
nor U3466 (N_3466,N_1427,N_2080);
nand U3467 (N_3467,N_1962,N_2024);
or U3468 (N_3468,N_960,N_2291);
nor U3469 (N_3469,N_39,N_2036);
and U3470 (N_3470,N_2022,N_904);
nor U3471 (N_3471,N_1803,N_615);
nand U3472 (N_3472,N_1846,N_1744);
or U3473 (N_3473,N_1038,N_2263);
and U3474 (N_3474,N_1050,N_1643);
nand U3475 (N_3475,N_1603,N_228);
and U3476 (N_3476,N_2266,N_1022);
nand U3477 (N_3477,N_1125,N_826);
nor U3478 (N_3478,N_350,N_1287);
and U3479 (N_3479,N_2101,N_1841);
nand U3480 (N_3480,N_1709,N_818);
nand U3481 (N_3481,N_352,N_1983);
and U3482 (N_3482,N_1797,N_64);
nand U3483 (N_3483,N_58,N_1924);
nor U3484 (N_3484,N_758,N_1037);
and U3485 (N_3485,N_866,N_468);
nor U3486 (N_3486,N_1882,N_1367);
and U3487 (N_3487,N_1742,N_2289);
and U3488 (N_3488,N_83,N_1884);
and U3489 (N_3489,N_910,N_1937);
and U3490 (N_3490,N_2197,N_1559);
nand U3491 (N_3491,N_106,N_1917);
nand U3492 (N_3492,N_2040,N_22);
nor U3493 (N_3493,N_1146,N_134);
nand U3494 (N_3494,N_462,N_1455);
or U3495 (N_3495,N_86,N_1223);
nor U3496 (N_3496,N_303,N_1271);
or U3497 (N_3497,N_1871,N_1201);
or U3498 (N_3498,N_1452,N_1345);
nor U3499 (N_3499,N_1198,N_349);
and U3500 (N_3500,N_230,N_640);
or U3501 (N_3501,N_139,N_876);
or U3502 (N_3502,N_1044,N_1141);
nor U3503 (N_3503,N_1840,N_2466);
or U3504 (N_3504,N_209,N_565);
nor U3505 (N_3505,N_1409,N_1225);
nor U3506 (N_3506,N_599,N_2055);
xnor U3507 (N_3507,N_509,N_215);
nand U3508 (N_3508,N_705,N_399);
or U3509 (N_3509,N_2376,N_1413);
or U3510 (N_3510,N_2190,N_1608);
xnor U3511 (N_3511,N_182,N_1511);
and U3512 (N_3512,N_877,N_2051);
or U3513 (N_3513,N_52,N_1480);
nand U3514 (N_3514,N_1695,N_2467);
or U3515 (N_3515,N_1896,N_256);
and U3516 (N_3516,N_631,N_364);
or U3517 (N_3517,N_1635,N_1746);
and U3518 (N_3518,N_513,N_2010);
nand U3519 (N_3519,N_1549,N_241);
nor U3520 (N_3520,N_2489,N_1387);
and U3521 (N_3521,N_1155,N_2490);
nor U3522 (N_3522,N_541,N_720);
and U3523 (N_3523,N_2229,N_2278);
nand U3524 (N_3524,N_1286,N_915);
or U3525 (N_3525,N_1955,N_512);
and U3526 (N_3526,N_239,N_2207);
or U3527 (N_3527,N_1291,N_1651);
and U3528 (N_3528,N_2409,N_1814);
nand U3529 (N_3529,N_2025,N_2238);
nand U3530 (N_3530,N_372,N_2168);
nand U3531 (N_3531,N_1191,N_1777);
or U3532 (N_3532,N_761,N_1304);
and U3533 (N_3533,N_2235,N_2113);
nand U3534 (N_3534,N_321,N_1669);
xor U3535 (N_3535,N_1832,N_1479);
nor U3536 (N_3536,N_333,N_2147);
nor U3537 (N_3537,N_1671,N_1984);
nor U3538 (N_3538,N_781,N_1034);
or U3539 (N_3539,N_1399,N_1590);
or U3540 (N_3540,N_1343,N_772);
nand U3541 (N_3541,N_944,N_1698);
or U3542 (N_3542,N_1712,N_2230);
and U3543 (N_3543,N_1082,N_2057);
nor U3544 (N_3544,N_2210,N_1689);
or U3545 (N_3545,N_1652,N_346);
nand U3546 (N_3546,N_2292,N_1968);
or U3547 (N_3547,N_1851,N_1389);
or U3548 (N_3548,N_1120,N_777);
or U3549 (N_3549,N_1052,N_1845);
or U3550 (N_3550,N_1002,N_59);
nor U3551 (N_3551,N_10,N_1829);
and U3552 (N_3552,N_2374,N_2472);
nor U3553 (N_3553,N_1743,N_367);
nand U3554 (N_3554,N_1138,N_1764);
nand U3555 (N_3555,N_74,N_533);
or U3556 (N_3556,N_1496,N_2246);
nand U3557 (N_3557,N_412,N_1772);
or U3558 (N_3558,N_144,N_2186);
or U3559 (N_3559,N_2319,N_952);
or U3560 (N_3560,N_806,N_475);
nand U3561 (N_3561,N_2115,N_890);
xor U3562 (N_3562,N_1254,N_1290);
and U3563 (N_3563,N_883,N_274);
nand U3564 (N_3564,N_1107,N_1957);
and U3565 (N_3565,N_2439,N_1307);
nand U3566 (N_3566,N_1268,N_1180);
nand U3567 (N_3567,N_1433,N_741);
and U3568 (N_3568,N_1617,N_1013);
nor U3569 (N_3569,N_1580,N_2470);
nand U3570 (N_3570,N_1179,N_390);
nor U3571 (N_3571,N_1247,N_1071);
nor U3572 (N_3572,N_1269,N_1250);
nor U3573 (N_3573,N_2330,N_2362);
nor U3574 (N_3574,N_284,N_2087);
nand U3575 (N_3575,N_96,N_2457);
or U3576 (N_3576,N_94,N_596);
and U3577 (N_3577,N_396,N_1694);
nor U3578 (N_3578,N_114,N_1414);
nor U3579 (N_3579,N_1412,N_1681);
nor U3580 (N_3580,N_1956,N_2074);
nor U3581 (N_3581,N_498,N_722);
nand U3582 (N_3582,N_1565,N_609);
and U3583 (N_3583,N_1339,N_322);
nand U3584 (N_3584,N_830,N_570);
nor U3585 (N_3585,N_1696,N_2094);
or U3586 (N_3586,N_1192,N_2016);
nand U3587 (N_3587,N_1,N_1352);
and U3588 (N_3588,N_1516,N_545);
and U3589 (N_3589,N_379,N_584);
nand U3590 (N_3590,N_1708,N_378);
nor U3591 (N_3591,N_28,N_1658);
or U3592 (N_3592,N_316,N_1705);
nand U3593 (N_3593,N_1964,N_1365);
or U3594 (N_3594,N_406,N_314);
and U3595 (N_3595,N_598,N_1707);
nand U3596 (N_3596,N_2028,N_2082);
nor U3597 (N_3597,N_1942,N_1444);
and U3598 (N_3598,N_1813,N_2015);
nand U3599 (N_3599,N_2384,N_434);
nand U3600 (N_3600,N_882,N_1423);
and U3601 (N_3601,N_1303,N_1094);
nor U3602 (N_3602,N_111,N_964);
and U3603 (N_3603,N_477,N_2107);
and U3604 (N_3604,N_795,N_701);
nor U3605 (N_3605,N_176,N_2354);
nor U3606 (N_3606,N_2456,N_747);
nand U3607 (N_3607,N_607,N_2261);
nand U3608 (N_3608,N_2265,N_2410);
or U3609 (N_3609,N_2460,N_1084);
and U3610 (N_3610,N_1655,N_1098);
nand U3611 (N_3611,N_98,N_1426);
or U3612 (N_3612,N_2033,N_353);
nor U3613 (N_3613,N_2307,N_766);
nor U3614 (N_3614,N_123,N_606);
or U3615 (N_3615,N_1055,N_1729);
nor U3616 (N_3616,N_2084,N_273);
nand U3617 (N_3617,N_2443,N_2072);
and U3618 (N_3618,N_814,N_1208);
nor U3619 (N_3619,N_653,N_930);
nand U3620 (N_3620,N_1323,N_210);
and U3621 (N_3621,N_1551,N_819);
nand U3622 (N_3622,N_1077,N_430);
nand U3623 (N_3623,N_1656,N_2334);
and U3624 (N_3624,N_1980,N_786);
and U3625 (N_3625,N_482,N_2486);
or U3626 (N_3626,N_301,N_739);
nor U3627 (N_3627,N_377,N_1429);
or U3628 (N_3628,N_908,N_166);
and U3629 (N_3629,N_2141,N_450);
nor U3630 (N_3630,N_1837,N_613);
and U3631 (N_3631,N_165,N_1863);
xnor U3632 (N_3632,N_1931,N_2159);
or U3633 (N_3633,N_1110,N_1154);
or U3634 (N_3634,N_402,N_1460);
and U3635 (N_3635,N_357,N_113);
and U3636 (N_3636,N_1039,N_1197);
or U3637 (N_3637,N_544,N_1895);
or U3638 (N_3638,N_1105,N_564);
nand U3639 (N_3639,N_163,N_403);
or U3640 (N_3640,N_1945,N_1295);
xnor U3641 (N_3641,N_2039,N_2126);
and U3642 (N_3642,N_661,N_2220);
or U3643 (N_3643,N_1755,N_791);
nor U3644 (N_3644,N_1469,N_497);
xor U3645 (N_3645,N_931,N_1348);
or U3646 (N_3646,N_1795,N_1363);
nand U3647 (N_3647,N_800,N_2091);
nand U3648 (N_3648,N_1187,N_223);
or U3649 (N_3649,N_1716,N_2093);
nor U3650 (N_3650,N_1951,N_1381);
nor U3651 (N_3651,N_783,N_217);
nand U3652 (N_3652,N_490,N_553);
or U3653 (N_3653,N_1405,N_1369);
nand U3654 (N_3654,N_129,N_2326);
or U3655 (N_3655,N_1798,N_1557);
nor U3656 (N_3656,N_788,N_445);
nor U3657 (N_3657,N_711,N_1891);
and U3658 (N_3658,N_1628,N_1215);
or U3659 (N_3659,N_1584,N_1278);
or U3660 (N_3660,N_1333,N_461);
and U3661 (N_3661,N_1714,N_1375);
or U3662 (N_3662,N_331,N_1209);
and U3663 (N_3663,N_534,N_1313);
nand U3664 (N_3664,N_2193,N_2069);
nand U3665 (N_3665,N_381,N_677);
and U3666 (N_3666,N_1402,N_922);
xnor U3667 (N_3667,N_478,N_420);
or U3668 (N_3668,N_2465,N_566);
nand U3669 (N_3669,N_2378,N_666);
nand U3670 (N_3670,N_680,N_1809);
or U3671 (N_3671,N_1727,N_2184);
and U3672 (N_3672,N_1386,N_266);
nand U3673 (N_3673,N_2434,N_18);
nand U3674 (N_3674,N_895,N_943);
nand U3675 (N_3675,N_864,N_1591);
nor U3676 (N_3676,N_1263,N_519);
and U3677 (N_3677,N_178,N_1158);
or U3678 (N_3678,N_602,N_724);
and U3679 (N_3679,N_426,N_1003);
xnor U3680 (N_3680,N_1508,N_543);
nor U3681 (N_3681,N_1066,N_2464);
nor U3682 (N_3682,N_623,N_2256);
or U3683 (N_3683,N_2430,N_746);
nand U3684 (N_3684,N_1801,N_1892);
and U3685 (N_3685,N_1934,N_416);
nor U3686 (N_3686,N_984,N_1928);
and U3687 (N_3687,N_1296,N_290);
nand U3688 (N_3688,N_1033,N_1542);
nor U3689 (N_3689,N_2353,N_2357);
nand U3690 (N_3690,N_1525,N_670);
xnor U3691 (N_3691,N_358,N_2079);
or U3692 (N_3692,N_1780,N_1666);
nor U3693 (N_3693,N_1168,N_1030);
or U3694 (N_3694,N_2317,N_251);
and U3695 (N_3695,N_778,N_993);
and U3696 (N_3696,N_1257,N_235);
nand U3697 (N_3697,N_668,N_60);
nor U3698 (N_3698,N_453,N_1905);
and U3699 (N_3699,N_271,N_1106);
and U3700 (N_3700,N_2432,N_1553);
or U3701 (N_3701,N_1430,N_1126);
or U3702 (N_3702,N_542,N_1699);
xor U3703 (N_3703,N_409,N_2174);
and U3704 (N_3704,N_2453,N_20);
and U3705 (N_3705,N_1927,N_1284);
and U3706 (N_3706,N_899,N_2103);
or U3707 (N_3707,N_306,N_105);
and U3708 (N_3708,N_1805,N_2071);
or U3709 (N_3709,N_1212,N_1222);
or U3710 (N_3710,N_287,N_1462);
nand U3711 (N_3711,N_1083,N_1820);
nand U3712 (N_3712,N_1394,N_2065);
or U3713 (N_3713,N_1134,N_267);
or U3714 (N_3714,N_1325,N_347);
or U3715 (N_3715,N_265,N_1767);
nand U3716 (N_3716,N_2273,N_369);
or U3717 (N_3717,N_782,N_525);
nand U3718 (N_3718,N_272,N_614);
nand U3719 (N_3719,N_132,N_1514);
nor U3720 (N_3720,N_1794,N_556);
or U3721 (N_3721,N_2491,N_1337);
nand U3722 (N_3722,N_660,N_824);
and U3723 (N_3723,N_1834,N_431);
or U3724 (N_3724,N_1547,N_845);
and U3725 (N_3725,N_16,N_1781);
nand U3726 (N_3726,N_2441,N_1099);
xor U3727 (N_3727,N_729,N_2394);
nor U3728 (N_3728,N_476,N_1028);
or U3729 (N_3729,N_2078,N_48);
or U3730 (N_3730,N_2132,N_947);
and U3731 (N_3731,N_1886,N_708);
and U3732 (N_3732,N_55,N_2447);
nor U3733 (N_3733,N_62,N_2323);
or U3734 (N_3734,N_2075,N_1611);
or U3735 (N_3735,N_1913,N_1531);
nand U3736 (N_3736,N_546,N_1963);
nor U3737 (N_3737,N_285,N_2100);
and U3738 (N_3738,N_1718,N_463);
nand U3739 (N_3739,N_1431,N_2494);
and U3740 (N_3740,N_835,N_1058);
and U3741 (N_3741,N_438,N_2002);
nand U3742 (N_3742,N_621,N_858);
and U3743 (N_3743,N_109,N_1229);
and U3744 (N_3744,N_844,N_1318);
nor U3745 (N_3745,N_250,N_1061);
nor U3746 (N_3746,N_1454,N_2169);
nand U3747 (N_3747,N_42,N_1362);
nor U3748 (N_3748,N_133,N_1463);
or U3749 (N_3749,N_2090,N_760);
nand U3750 (N_3750,N_1275,N_393);
and U3751 (N_3751,N_1799,N_93);
nand U3752 (N_3752,N_1563,N_710);
or U3753 (N_3753,N_1132,N_1410);
xor U3754 (N_3754,N_2149,N_2127);
and U3755 (N_3755,N_1677,N_1239);
nor U3756 (N_3756,N_2283,N_94);
or U3757 (N_3757,N_788,N_900);
or U3758 (N_3758,N_616,N_1127);
and U3759 (N_3759,N_1700,N_2397);
and U3760 (N_3760,N_508,N_438);
and U3761 (N_3761,N_736,N_2415);
or U3762 (N_3762,N_2331,N_840);
nand U3763 (N_3763,N_1637,N_500);
or U3764 (N_3764,N_1796,N_2075);
and U3765 (N_3765,N_835,N_1989);
or U3766 (N_3766,N_68,N_1715);
and U3767 (N_3767,N_2081,N_542);
and U3768 (N_3768,N_698,N_76);
and U3769 (N_3769,N_1148,N_1565);
and U3770 (N_3770,N_2356,N_807);
or U3771 (N_3771,N_876,N_1874);
xnor U3772 (N_3772,N_1069,N_2343);
or U3773 (N_3773,N_1188,N_654);
nand U3774 (N_3774,N_310,N_1922);
and U3775 (N_3775,N_1428,N_1113);
nand U3776 (N_3776,N_117,N_910);
xor U3777 (N_3777,N_1121,N_946);
nand U3778 (N_3778,N_1111,N_1045);
and U3779 (N_3779,N_1351,N_1816);
nor U3780 (N_3780,N_2156,N_368);
or U3781 (N_3781,N_857,N_1044);
and U3782 (N_3782,N_1613,N_623);
or U3783 (N_3783,N_728,N_186);
nor U3784 (N_3784,N_1272,N_1443);
nor U3785 (N_3785,N_960,N_1550);
and U3786 (N_3786,N_2304,N_1823);
and U3787 (N_3787,N_564,N_39);
nand U3788 (N_3788,N_2344,N_1485);
and U3789 (N_3789,N_5,N_1439);
or U3790 (N_3790,N_2236,N_2364);
nand U3791 (N_3791,N_1485,N_214);
and U3792 (N_3792,N_433,N_1612);
or U3793 (N_3793,N_2282,N_760);
nor U3794 (N_3794,N_1862,N_292);
or U3795 (N_3795,N_1149,N_394);
or U3796 (N_3796,N_1288,N_1770);
nand U3797 (N_3797,N_2312,N_1628);
nand U3798 (N_3798,N_1169,N_267);
nor U3799 (N_3799,N_469,N_392);
or U3800 (N_3800,N_568,N_2052);
nand U3801 (N_3801,N_2080,N_692);
or U3802 (N_3802,N_512,N_1199);
or U3803 (N_3803,N_1006,N_1767);
or U3804 (N_3804,N_1019,N_1345);
nand U3805 (N_3805,N_2361,N_828);
and U3806 (N_3806,N_1512,N_1753);
and U3807 (N_3807,N_63,N_1976);
nor U3808 (N_3808,N_1692,N_976);
or U3809 (N_3809,N_2025,N_1924);
nand U3810 (N_3810,N_1504,N_85);
and U3811 (N_3811,N_90,N_2241);
and U3812 (N_3812,N_693,N_2153);
nand U3813 (N_3813,N_11,N_2160);
nand U3814 (N_3814,N_1177,N_2014);
nor U3815 (N_3815,N_262,N_511);
or U3816 (N_3816,N_588,N_1149);
nor U3817 (N_3817,N_956,N_2028);
and U3818 (N_3818,N_1732,N_2279);
nand U3819 (N_3819,N_1210,N_182);
nand U3820 (N_3820,N_920,N_1856);
nor U3821 (N_3821,N_233,N_984);
nand U3822 (N_3822,N_2224,N_349);
nand U3823 (N_3823,N_536,N_1488);
or U3824 (N_3824,N_179,N_975);
or U3825 (N_3825,N_1363,N_1176);
nor U3826 (N_3826,N_327,N_431);
or U3827 (N_3827,N_102,N_972);
xnor U3828 (N_3828,N_591,N_1585);
nor U3829 (N_3829,N_1157,N_260);
and U3830 (N_3830,N_189,N_16);
nor U3831 (N_3831,N_414,N_526);
nor U3832 (N_3832,N_584,N_876);
or U3833 (N_3833,N_1036,N_1881);
nor U3834 (N_3834,N_675,N_875);
nand U3835 (N_3835,N_2082,N_2189);
and U3836 (N_3836,N_2105,N_1096);
xnor U3837 (N_3837,N_72,N_1867);
and U3838 (N_3838,N_1121,N_814);
and U3839 (N_3839,N_1067,N_2423);
nor U3840 (N_3840,N_604,N_699);
nand U3841 (N_3841,N_293,N_1865);
and U3842 (N_3842,N_1879,N_2227);
and U3843 (N_3843,N_677,N_1523);
and U3844 (N_3844,N_1639,N_1708);
nor U3845 (N_3845,N_1261,N_1012);
and U3846 (N_3846,N_1348,N_291);
or U3847 (N_3847,N_1923,N_1065);
nand U3848 (N_3848,N_648,N_282);
or U3849 (N_3849,N_1279,N_169);
nand U3850 (N_3850,N_1610,N_299);
or U3851 (N_3851,N_551,N_1699);
nand U3852 (N_3852,N_138,N_34);
or U3853 (N_3853,N_2292,N_1921);
nand U3854 (N_3854,N_923,N_975);
nor U3855 (N_3855,N_2019,N_2178);
nor U3856 (N_3856,N_1963,N_26);
nand U3857 (N_3857,N_471,N_795);
nand U3858 (N_3858,N_2233,N_621);
nor U3859 (N_3859,N_2238,N_2475);
and U3860 (N_3860,N_2289,N_2436);
nand U3861 (N_3861,N_577,N_1017);
nor U3862 (N_3862,N_1653,N_1602);
nand U3863 (N_3863,N_1404,N_440);
nor U3864 (N_3864,N_2041,N_1326);
nor U3865 (N_3865,N_2358,N_1364);
and U3866 (N_3866,N_1776,N_752);
or U3867 (N_3867,N_256,N_1946);
or U3868 (N_3868,N_1393,N_276);
or U3869 (N_3869,N_2256,N_1591);
and U3870 (N_3870,N_2225,N_0);
and U3871 (N_3871,N_1746,N_1398);
or U3872 (N_3872,N_308,N_2358);
nor U3873 (N_3873,N_1614,N_1072);
nor U3874 (N_3874,N_2142,N_2314);
nor U3875 (N_3875,N_1673,N_711);
nand U3876 (N_3876,N_2447,N_1773);
and U3877 (N_3877,N_935,N_505);
nor U3878 (N_3878,N_1933,N_153);
nand U3879 (N_3879,N_543,N_2295);
nor U3880 (N_3880,N_308,N_1826);
nor U3881 (N_3881,N_1066,N_2321);
and U3882 (N_3882,N_2159,N_19);
nor U3883 (N_3883,N_1391,N_629);
or U3884 (N_3884,N_1669,N_1361);
nor U3885 (N_3885,N_1044,N_2153);
and U3886 (N_3886,N_520,N_2346);
or U3887 (N_3887,N_1290,N_170);
nor U3888 (N_3888,N_394,N_44);
or U3889 (N_3889,N_1851,N_5);
or U3890 (N_3890,N_437,N_1012);
nor U3891 (N_3891,N_2449,N_844);
nor U3892 (N_3892,N_2280,N_424);
nand U3893 (N_3893,N_1175,N_541);
nand U3894 (N_3894,N_2192,N_884);
and U3895 (N_3895,N_866,N_783);
nand U3896 (N_3896,N_1300,N_1510);
nor U3897 (N_3897,N_2169,N_1910);
nand U3898 (N_3898,N_44,N_312);
and U3899 (N_3899,N_1058,N_1066);
and U3900 (N_3900,N_1915,N_387);
and U3901 (N_3901,N_2292,N_1445);
nor U3902 (N_3902,N_1173,N_16);
and U3903 (N_3903,N_2305,N_1922);
and U3904 (N_3904,N_729,N_492);
nand U3905 (N_3905,N_1153,N_1604);
nor U3906 (N_3906,N_2193,N_1287);
and U3907 (N_3907,N_1611,N_101);
nand U3908 (N_3908,N_1577,N_1022);
or U3909 (N_3909,N_72,N_102);
xnor U3910 (N_3910,N_1592,N_472);
nor U3911 (N_3911,N_1119,N_1659);
or U3912 (N_3912,N_1353,N_482);
and U3913 (N_3913,N_1628,N_393);
or U3914 (N_3914,N_2442,N_1768);
nor U3915 (N_3915,N_177,N_983);
or U3916 (N_3916,N_120,N_644);
nand U3917 (N_3917,N_1468,N_2440);
and U3918 (N_3918,N_212,N_2242);
and U3919 (N_3919,N_1921,N_1811);
or U3920 (N_3920,N_1530,N_1335);
or U3921 (N_3921,N_2160,N_1939);
or U3922 (N_3922,N_925,N_5);
nand U3923 (N_3923,N_1178,N_2425);
nand U3924 (N_3924,N_11,N_385);
and U3925 (N_3925,N_928,N_452);
and U3926 (N_3926,N_2314,N_1591);
or U3927 (N_3927,N_1169,N_1840);
or U3928 (N_3928,N_1760,N_428);
nor U3929 (N_3929,N_381,N_1617);
nand U3930 (N_3930,N_1922,N_2055);
nand U3931 (N_3931,N_1523,N_462);
nor U3932 (N_3932,N_128,N_1943);
or U3933 (N_3933,N_1783,N_2397);
or U3934 (N_3934,N_2119,N_1669);
or U3935 (N_3935,N_524,N_12);
nand U3936 (N_3936,N_713,N_2230);
or U3937 (N_3937,N_2144,N_60);
and U3938 (N_3938,N_2071,N_1296);
nand U3939 (N_3939,N_307,N_868);
nor U3940 (N_3940,N_1927,N_2188);
and U3941 (N_3941,N_1303,N_796);
or U3942 (N_3942,N_1213,N_1924);
nor U3943 (N_3943,N_1067,N_169);
nand U3944 (N_3944,N_710,N_475);
and U3945 (N_3945,N_569,N_425);
nor U3946 (N_3946,N_1599,N_1347);
or U3947 (N_3947,N_1555,N_384);
or U3948 (N_3948,N_717,N_955);
and U3949 (N_3949,N_1874,N_2410);
nand U3950 (N_3950,N_604,N_1892);
or U3951 (N_3951,N_234,N_717);
nor U3952 (N_3952,N_1375,N_1864);
nand U3953 (N_3953,N_26,N_2085);
nor U3954 (N_3954,N_1949,N_2388);
nor U3955 (N_3955,N_2022,N_2364);
nand U3956 (N_3956,N_1442,N_2120);
nand U3957 (N_3957,N_2036,N_1495);
nor U3958 (N_3958,N_781,N_1267);
nand U3959 (N_3959,N_2056,N_346);
nand U3960 (N_3960,N_1368,N_730);
nor U3961 (N_3961,N_1217,N_322);
or U3962 (N_3962,N_1168,N_29);
nor U3963 (N_3963,N_499,N_123);
or U3964 (N_3964,N_2403,N_2202);
and U3965 (N_3965,N_1092,N_1218);
or U3966 (N_3966,N_1651,N_2031);
or U3967 (N_3967,N_83,N_1637);
nand U3968 (N_3968,N_1205,N_991);
nand U3969 (N_3969,N_1886,N_1944);
nor U3970 (N_3970,N_1347,N_1004);
and U3971 (N_3971,N_952,N_2085);
nor U3972 (N_3972,N_536,N_1000);
or U3973 (N_3973,N_1646,N_2424);
nor U3974 (N_3974,N_872,N_1952);
and U3975 (N_3975,N_1284,N_64);
nor U3976 (N_3976,N_1976,N_616);
or U3977 (N_3977,N_900,N_2354);
or U3978 (N_3978,N_221,N_1786);
nor U3979 (N_3979,N_257,N_875);
nor U3980 (N_3980,N_609,N_1352);
xnor U3981 (N_3981,N_2249,N_2069);
nand U3982 (N_3982,N_553,N_150);
and U3983 (N_3983,N_1668,N_1567);
nand U3984 (N_3984,N_2279,N_2047);
and U3985 (N_3985,N_2039,N_1816);
xor U3986 (N_3986,N_1018,N_1747);
nor U3987 (N_3987,N_290,N_311);
nor U3988 (N_3988,N_2303,N_2123);
or U3989 (N_3989,N_470,N_177);
nor U3990 (N_3990,N_1914,N_983);
and U3991 (N_3991,N_1840,N_2416);
or U3992 (N_3992,N_1768,N_2105);
and U3993 (N_3993,N_1697,N_1848);
or U3994 (N_3994,N_45,N_2283);
and U3995 (N_3995,N_131,N_521);
and U3996 (N_3996,N_2399,N_335);
nor U3997 (N_3997,N_2356,N_1979);
or U3998 (N_3998,N_2418,N_2001);
and U3999 (N_3999,N_1042,N_1706);
and U4000 (N_4000,N_544,N_1982);
or U4001 (N_4001,N_399,N_1267);
or U4002 (N_4002,N_1839,N_1302);
nand U4003 (N_4003,N_115,N_1120);
nand U4004 (N_4004,N_395,N_1110);
or U4005 (N_4005,N_729,N_1377);
xnor U4006 (N_4006,N_716,N_67);
nor U4007 (N_4007,N_917,N_1031);
nand U4008 (N_4008,N_1245,N_242);
and U4009 (N_4009,N_1049,N_1317);
nor U4010 (N_4010,N_1147,N_16);
and U4011 (N_4011,N_1490,N_1441);
and U4012 (N_4012,N_1571,N_2483);
or U4013 (N_4013,N_1809,N_150);
nor U4014 (N_4014,N_486,N_330);
or U4015 (N_4015,N_1493,N_272);
and U4016 (N_4016,N_2431,N_611);
xor U4017 (N_4017,N_2017,N_650);
nor U4018 (N_4018,N_1556,N_823);
nand U4019 (N_4019,N_787,N_1974);
nor U4020 (N_4020,N_1738,N_820);
nand U4021 (N_4021,N_1396,N_1603);
and U4022 (N_4022,N_642,N_549);
nor U4023 (N_4023,N_2077,N_1345);
nor U4024 (N_4024,N_1047,N_1956);
nor U4025 (N_4025,N_541,N_702);
nand U4026 (N_4026,N_1541,N_2481);
nand U4027 (N_4027,N_2184,N_701);
nand U4028 (N_4028,N_1677,N_1261);
or U4029 (N_4029,N_1696,N_1223);
or U4030 (N_4030,N_1716,N_1915);
or U4031 (N_4031,N_1415,N_2118);
nor U4032 (N_4032,N_981,N_1906);
or U4033 (N_4033,N_2001,N_833);
and U4034 (N_4034,N_2291,N_1632);
or U4035 (N_4035,N_168,N_1936);
and U4036 (N_4036,N_453,N_2147);
and U4037 (N_4037,N_60,N_2418);
nand U4038 (N_4038,N_1890,N_620);
or U4039 (N_4039,N_797,N_1488);
and U4040 (N_4040,N_956,N_1085);
and U4041 (N_4041,N_1411,N_2036);
and U4042 (N_4042,N_1830,N_2372);
and U4043 (N_4043,N_153,N_997);
nor U4044 (N_4044,N_1007,N_1310);
nand U4045 (N_4045,N_2254,N_1940);
nor U4046 (N_4046,N_259,N_1161);
nor U4047 (N_4047,N_2191,N_2105);
nor U4048 (N_4048,N_776,N_1380);
and U4049 (N_4049,N_1715,N_12);
and U4050 (N_4050,N_396,N_752);
nand U4051 (N_4051,N_2039,N_2157);
xor U4052 (N_4052,N_114,N_1991);
nor U4053 (N_4053,N_914,N_499);
nand U4054 (N_4054,N_376,N_103);
and U4055 (N_4055,N_280,N_2264);
and U4056 (N_4056,N_2110,N_460);
or U4057 (N_4057,N_91,N_17);
nand U4058 (N_4058,N_381,N_348);
nand U4059 (N_4059,N_1318,N_1369);
nor U4060 (N_4060,N_996,N_2313);
nor U4061 (N_4061,N_581,N_494);
nor U4062 (N_4062,N_1660,N_1401);
xnor U4063 (N_4063,N_1750,N_976);
nor U4064 (N_4064,N_123,N_753);
nand U4065 (N_4065,N_1914,N_1641);
or U4066 (N_4066,N_964,N_128);
nand U4067 (N_4067,N_2412,N_2090);
or U4068 (N_4068,N_1985,N_850);
and U4069 (N_4069,N_1233,N_340);
and U4070 (N_4070,N_842,N_1305);
nor U4071 (N_4071,N_1842,N_990);
nor U4072 (N_4072,N_1788,N_1371);
and U4073 (N_4073,N_237,N_1242);
and U4074 (N_4074,N_254,N_1633);
nor U4075 (N_4075,N_2014,N_2380);
nor U4076 (N_4076,N_2121,N_2129);
nand U4077 (N_4077,N_1657,N_2128);
and U4078 (N_4078,N_295,N_2267);
nand U4079 (N_4079,N_298,N_1333);
nor U4080 (N_4080,N_2292,N_1810);
and U4081 (N_4081,N_1523,N_1087);
nor U4082 (N_4082,N_1283,N_2321);
nand U4083 (N_4083,N_593,N_616);
nor U4084 (N_4084,N_917,N_300);
or U4085 (N_4085,N_535,N_1773);
xnor U4086 (N_4086,N_1947,N_1328);
or U4087 (N_4087,N_2184,N_2296);
nor U4088 (N_4088,N_2235,N_280);
and U4089 (N_4089,N_1315,N_1206);
and U4090 (N_4090,N_855,N_109);
and U4091 (N_4091,N_1853,N_1551);
and U4092 (N_4092,N_115,N_1990);
nor U4093 (N_4093,N_225,N_1279);
nor U4094 (N_4094,N_2303,N_59);
or U4095 (N_4095,N_67,N_927);
nor U4096 (N_4096,N_2151,N_194);
or U4097 (N_4097,N_1518,N_127);
nand U4098 (N_4098,N_917,N_1397);
nor U4099 (N_4099,N_1601,N_1123);
and U4100 (N_4100,N_989,N_2495);
nand U4101 (N_4101,N_2108,N_1021);
and U4102 (N_4102,N_1275,N_1812);
nor U4103 (N_4103,N_770,N_1804);
or U4104 (N_4104,N_605,N_2428);
or U4105 (N_4105,N_1600,N_2150);
nand U4106 (N_4106,N_1953,N_1204);
or U4107 (N_4107,N_2357,N_1558);
nand U4108 (N_4108,N_78,N_653);
nor U4109 (N_4109,N_1189,N_1483);
and U4110 (N_4110,N_1237,N_76);
or U4111 (N_4111,N_743,N_2238);
nor U4112 (N_4112,N_660,N_1451);
and U4113 (N_4113,N_321,N_1579);
and U4114 (N_4114,N_1053,N_587);
nand U4115 (N_4115,N_1932,N_2265);
nand U4116 (N_4116,N_2207,N_178);
nand U4117 (N_4117,N_1563,N_762);
and U4118 (N_4118,N_2204,N_492);
or U4119 (N_4119,N_1706,N_244);
or U4120 (N_4120,N_2101,N_188);
and U4121 (N_4121,N_1068,N_2327);
and U4122 (N_4122,N_1597,N_811);
and U4123 (N_4123,N_1561,N_1613);
or U4124 (N_4124,N_1538,N_1829);
nand U4125 (N_4125,N_1763,N_2383);
nor U4126 (N_4126,N_720,N_1989);
nand U4127 (N_4127,N_2227,N_1661);
or U4128 (N_4128,N_2418,N_2172);
nand U4129 (N_4129,N_2171,N_604);
nand U4130 (N_4130,N_504,N_1432);
xnor U4131 (N_4131,N_2234,N_1722);
and U4132 (N_4132,N_2,N_1184);
nor U4133 (N_4133,N_1904,N_2235);
and U4134 (N_4134,N_1802,N_1556);
nor U4135 (N_4135,N_2466,N_1860);
and U4136 (N_4136,N_1461,N_709);
or U4137 (N_4137,N_2422,N_1888);
nand U4138 (N_4138,N_1017,N_668);
and U4139 (N_4139,N_1214,N_1411);
or U4140 (N_4140,N_972,N_452);
xnor U4141 (N_4141,N_1549,N_1583);
nand U4142 (N_4142,N_1134,N_2065);
nor U4143 (N_4143,N_1511,N_1581);
nor U4144 (N_4144,N_795,N_1474);
and U4145 (N_4145,N_1876,N_1076);
nor U4146 (N_4146,N_2163,N_2057);
or U4147 (N_4147,N_1906,N_1498);
nor U4148 (N_4148,N_374,N_766);
nor U4149 (N_4149,N_1263,N_1130);
or U4150 (N_4150,N_1090,N_1593);
nand U4151 (N_4151,N_719,N_1603);
xor U4152 (N_4152,N_84,N_377);
or U4153 (N_4153,N_651,N_1792);
and U4154 (N_4154,N_1405,N_747);
or U4155 (N_4155,N_15,N_629);
and U4156 (N_4156,N_1650,N_1059);
and U4157 (N_4157,N_289,N_1389);
nand U4158 (N_4158,N_1131,N_1120);
nand U4159 (N_4159,N_344,N_647);
nor U4160 (N_4160,N_895,N_2238);
or U4161 (N_4161,N_1475,N_596);
nor U4162 (N_4162,N_2496,N_630);
nand U4163 (N_4163,N_654,N_1814);
nor U4164 (N_4164,N_1139,N_1394);
nor U4165 (N_4165,N_2035,N_2214);
nand U4166 (N_4166,N_1689,N_981);
and U4167 (N_4167,N_1883,N_1020);
nor U4168 (N_4168,N_2415,N_1396);
nand U4169 (N_4169,N_2061,N_1326);
nor U4170 (N_4170,N_204,N_1368);
nor U4171 (N_4171,N_1365,N_2267);
nor U4172 (N_4172,N_28,N_457);
or U4173 (N_4173,N_2147,N_106);
nand U4174 (N_4174,N_2319,N_2414);
and U4175 (N_4175,N_275,N_2241);
nor U4176 (N_4176,N_2081,N_656);
nor U4177 (N_4177,N_2153,N_1572);
and U4178 (N_4178,N_380,N_1024);
nor U4179 (N_4179,N_2052,N_918);
nor U4180 (N_4180,N_813,N_603);
nand U4181 (N_4181,N_1521,N_1622);
and U4182 (N_4182,N_754,N_448);
nand U4183 (N_4183,N_1651,N_543);
nor U4184 (N_4184,N_1761,N_1083);
or U4185 (N_4185,N_2329,N_257);
and U4186 (N_4186,N_493,N_959);
xnor U4187 (N_4187,N_1102,N_1515);
nor U4188 (N_4188,N_1742,N_1805);
and U4189 (N_4189,N_1208,N_1944);
nor U4190 (N_4190,N_456,N_1942);
nand U4191 (N_4191,N_865,N_1063);
or U4192 (N_4192,N_1449,N_2324);
and U4193 (N_4193,N_821,N_2272);
or U4194 (N_4194,N_613,N_1802);
or U4195 (N_4195,N_486,N_635);
or U4196 (N_4196,N_85,N_2130);
and U4197 (N_4197,N_1855,N_890);
or U4198 (N_4198,N_1771,N_2270);
or U4199 (N_4199,N_1915,N_1979);
nand U4200 (N_4200,N_717,N_658);
nand U4201 (N_4201,N_1539,N_758);
or U4202 (N_4202,N_1606,N_409);
and U4203 (N_4203,N_2078,N_1956);
or U4204 (N_4204,N_2184,N_1503);
nor U4205 (N_4205,N_2464,N_847);
and U4206 (N_4206,N_296,N_968);
and U4207 (N_4207,N_1337,N_261);
and U4208 (N_4208,N_309,N_590);
or U4209 (N_4209,N_2110,N_422);
nor U4210 (N_4210,N_1142,N_715);
or U4211 (N_4211,N_831,N_2360);
or U4212 (N_4212,N_163,N_1994);
nor U4213 (N_4213,N_740,N_1105);
nor U4214 (N_4214,N_1002,N_2099);
nor U4215 (N_4215,N_2452,N_74);
nand U4216 (N_4216,N_1784,N_2151);
or U4217 (N_4217,N_1408,N_1701);
xnor U4218 (N_4218,N_902,N_642);
or U4219 (N_4219,N_2084,N_1096);
nand U4220 (N_4220,N_2255,N_2206);
nand U4221 (N_4221,N_265,N_1929);
and U4222 (N_4222,N_1066,N_850);
and U4223 (N_4223,N_53,N_1467);
nor U4224 (N_4224,N_2194,N_1260);
xnor U4225 (N_4225,N_2146,N_1183);
nor U4226 (N_4226,N_437,N_1683);
nand U4227 (N_4227,N_1650,N_2456);
nand U4228 (N_4228,N_1096,N_1765);
nor U4229 (N_4229,N_309,N_482);
and U4230 (N_4230,N_1473,N_1262);
nand U4231 (N_4231,N_2456,N_954);
nor U4232 (N_4232,N_2490,N_377);
or U4233 (N_4233,N_2054,N_2217);
and U4234 (N_4234,N_2444,N_2311);
nand U4235 (N_4235,N_61,N_1865);
and U4236 (N_4236,N_608,N_233);
nand U4237 (N_4237,N_433,N_962);
or U4238 (N_4238,N_1432,N_2201);
and U4239 (N_4239,N_2224,N_1573);
or U4240 (N_4240,N_898,N_1589);
or U4241 (N_4241,N_2151,N_2388);
nand U4242 (N_4242,N_1193,N_608);
xnor U4243 (N_4243,N_671,N_1557);
nand U4244 (N_4244,N_2415,N_1588);
xor U4245 (N_4245,N_2206,N_1014);
or U4246 (N_4246,N_1487,N_2138);
nor U4247 (N_4247,N_1477,N_1012);
or U4248 (N_4248,N_1768,N_947);
nand U4249 (N_4249,N_574,N_275);
or U4250 (N_4250,N_681,N_826);
nand U4251 (N_4251,N_1667,N_396);
nor U4252 (N_4252,N_674,N_1439);
nand U4253 (N_4253,N_1580,N_2134);
or U4254 (N_4254,N_686,N_1863);
nor U4255 (N_4255,N_402,N_1431);
nand U4256 (N_4256,N_1450,N_2421);
or U4257 (N_4257,N_2355,N_507);
and U4258 (N_4258,N_2394,N_899);
nand U4259 (N_4259,N_964,N_1314);
and U4260 (N_4260,N_1765,N_827);
or U4261 (N_4261,N_2498,N_152);
nor U4262 (N_4262,N_2152,N_874);
and U4263 (N_4263,N_2086,N_2408);
and U4264 (N_4264,N_890,N_1079);
nor U4265 (N_4265,N_793,N_62);
or U4266 (N_4266,N_2480,N_840);
and U4267 (N_4267,N_1573,N_2035);
or U4268 (N_4268,N_1884,N_2378);
or U4269 (N_4269,N_628,N_1437);
or U4270 (N_4270,N_511,N_1636);
nand U4271 (N_4271,N_2119,N_22);
or U4272 (N_4272,N_898,N_69);
nor U4273 (N_4273,N_1549,N_1018);
nand U4274 (N_4274,N_2447,N_1751);
nor U4275 (N_4275,N_1587,N_1238);
nand U4276 (N_4276,N_2382,N_62);
or U4277 (N_4277,N_1055,N_1238);
nor U4278 (N_4278,N_1926,N_2115);
or U4279 (N_4279,N_478,N_494);
nand U4280 (N_4280,N_371,N_2424);
nor U4281 (N_4281,N_1159,N_1447);
nand U4282 (N_4282,N_1177,N_1616);
nand U4283 (N_4283,N_1396,N_2430);
nand U4284 (N_4284,N_107,N_607);
nor U4285 (N_4285,N_2325,N_1334);
or U4286 (N_4286,N_1312,N_1030);
or U4287 (N_4287,N_1202,N_438);
and U4288 (N_4288,N_927,N_702);
and U4289 (N_4289,N_393,N_125);
nor U4290 (N_4290,N_903,N_2088);
nand U4291 (N_4291,N_1098,N_2352);
and U4292 (N_4292,N_555,N_681);
nor U4293 (N_4293,N_2315,N_1182);
or U4294 (N_4294,N_2178,N_2230);
nand U4295 (N_4295,N_1056,N_963);
nor U4296 (N_4296,N_268,N_2436);
nor U4297 (N_4297,N_1406,N_353);
or U4298 (N_4298,N_1782,N_181);
or U4299 (N_4299,N_2486,N_1671);
or U4300 (N_4300,N_423,N_2075);
nor U4301 (N_4301,N_286,N_188);
and U4302 (N_4302,N_791,N_139);
or U4303 (N_4303,N_2289,N_584);
nand U4304 (N_4304,N_746,N_251);
nand U4305 (N_4305,N_2063,N_1101);
or U4306 (N_4306,N_1904,N_654);
nor U4307 (N_4307,N_2305,N_666);
or U4308 (N_4308,N_864,N_653);
nor U4309 (N_4309,N_1139,N_2267);
and U4310 (N_4310,N_2190,N_2375);
and U4311 (N_4311,N_1227,N_2374);
nor U4312 (N_4312,N_315,N_663);
and U4313 (N_4313,N_198,N_1617);
nand U4314 (N_4314,N_347,N_172);
or U4315 (N_4315,N_254,N_170);
and U4316 (N_4316,N_2271,N_414);
nor U4317 (N_4317,N_1326,N_620);
or U4318 (N_4318,N_1270,N_798);
nand U4319 (N_4319,N_279,N_174);
or U4320 (N_4320,N_1001,N_1082);
nor U4321 (N_4321,N_817,N_1655);
nor U4322 (N_4322,N_2110,N_1347);
or U4323 (N_4323,N_1501,N_792);
nand U4324 (N_4324,N_1014,N_1764);
nand U4325 (N_4325,N_608,N_1415);
or U4326 (N_4326,N_1063,N_2452);
nor U4327 (N_4327,N_254,N_1914);
or U4328 (N_4328,N_1027,N_1281);
nand U4329 (N_4329,N_1522,N_1570);
nand U4330 (N_4330,N_2316,N_1015);
xor U4331 (N_4331,N_276,N_2034);
nor U4332 (N_4332,N_2073,N_520);
nand U4333 (N_4333,N_619,N_934);
nor U4334 (N_4334,N_2235,N_843);
nor U4335 (N_4335,N_1428,N_1808);
and U4336 (N_4336,N_1868,N_2486);
and U4337 (N_4337,N_2215,N_1678);
nor U4338 (N_4338,N_1279,N_1511);
and U4339 (N_4339,N_1452,N_223);
nand U4340 (N_4340,N_594,N_1168);
nand U4341 (N_4341,N_522,N_960);
or U4342 (N_4342,N_1904,N_54);
nor U4343 (N_4343,N_1569,N_1527);
and U4344 (N_4344,N_448,N_938);
nor U4345 (N_4345,N_2252,N_45);
and U4346 (N_4346,N_1596,N_90);
and U4347 (N_4347,N_562,N_211);
and U4348 (N_4348,N_1492,N_833);
and U4349 (N_4349,N_812,N_1283);
nor U4350 (N_4350,N_483,N_1505);
nor U4351 (N_4351,N_1428,N_903);
or U4352 (N_4352,N_1558,N_1375);
nor U4353 (N_4353,N_2112,N_756);
nand U4354 (N_4354,N_913,N_1693);
xnor U4355 (N_4355,N_1373,N_1811);
nor U4356 (N_4356,N_2262,N_2053);
and U4357 (N_4357,N_1666,N_2348);
nand U4358 (N_4358,N_1345,N_1430);
nand U4359 (N_4359,N_1952,N_930);
or U4360 (N_4360,N_443,N_2054);
nor U4361 (N_4361,N_791,N_1737);
nand U4362 (N_4362,N_917,N_1845);
or U4363 (N_4363,N_158,N_412);
xnor U4364 (N_4364,N_94,N_1407);
nor U4365 (N_4365,N_302,N_1578);
nor U4366 (N_4366,N_1161,N_2453);
or U4367 (N_4367,N_791,N_293);
or U4368 (N_4368,N_491,N_894);
or U4369 (N_4369,N_1997,N_1019);
nor U4370 (N_4370,N_1881,N_2480);
nand U4371 (N_4371,N_762,N_1060);
and U4372 (N_4372,N_475,N_1769);
and U4373 (N_4373,N_1379,N_1864);
xnor U4374 (N_4374,N_1933,N_470);
nor U4375 (N_4375,N_2004,N_769);
and U4376 (N_4376,N_367,N_1029);
nand U4377 (N_4377,N_783,N_1047);
nor U4378 (N_4378,N_1247,N_150);
or U4379 (N_4379,N_756,N_2135);
and U4380 (N_4380,N_1044,N_2476);
or U4381 (N_4381,N_1605,N_151);
and U4382 (N_4382,N_1785,N_1683);
nand U4383 (N_4383,N_899,N_529);
nor U4384 (N_4384,N_1377,N_115);
nor U4385 (N_4385,N_78,N_1377);
nand U4386 (N_4386,N_1496,N_1964);
nor U4387 (N_4387,N_552,N_2130);
or U4388 (N_4388,N_780,N_1944);
nor U4389 (N_4389,N_1897,N_2498);
and U4390 (N_4390,N_649,N_2306);
and U4391 (N_4391,N_1352,N_2486);
nor U4392 (N_4392,N_200,N_2347);
and U4393 (N_4393,N_1675,N_1793);
or U4394 (N_4394,N_2302,N_260);
and U4395 (N_4395,N_1044,N_1414);
and U4396 (N_4396,N_845,N_2312);
or U4397 (N_4397,N_1334,N_1638);
nor U4398 (N_4398,N_1148,N_587);
nor U4399 (N_4399,N_1555,N_252);
xor U4400 (N_4400,N_2144,N_475);
nand U4401 (N_4401,N_1420,N_703);
and U4402 (N_4402,N_1355,N_1354);
xnor U4403 (N_4403,N_2349,N_763);
nor U4404 (N_4404,N_1697,N_1075);
and U4405 (N_4405,N_2228,N_729);
and U4406 (N_4406,N_853,N_1695);
nor U4407 (N_4407,N_1332,N_546);
or U4408 (N_4408,N_210,N_849);
nand U4409 (N_4409,N_2177,N_744);
or U4410 (N_4410,N_204,N_760);
and U4411 (N_4411,N_783,N_1491);
nand U4412 (N_4412,N_2412,N_686);
nand U4413 (N_4413,N_328,N_133);
nor U4414 (N_4414,N_1699,N_97);
nand U4415 (N_4415,N_1697,N_1812);
or U4416 (N_4416,N_643,N_1017);
nand U4417 (N_4417,N_432,N_1753);
and U4418 (N_4418,N_2126,N_255);
or U4419 (N_4419,N_1569,N_775);
or U4420 (N_4420,N_304,N_1632);
nor U4421 (N_4421,N_530,N_1999);
nor U4422 (N_4422,N_574,N_799);
nand U4423 (N_4423,N_2338,N_2206);
nor U4424 (N_4424,N_1722,N_1118);
or U4425 (N_4425,N_2238,N_1392);
nor U4426 (N_4426,N_492,N_821);
and U4427 (N_4427,N_481,N_1872);
and U4428 (N_4428,N_112,N_1627);
or U4429 (N_4429,N_518,N_147);
nand U4430 (N_4430,N_1981,N_28);
nand U4431 (N_4431,N_811,N_1889);
nor U4432 (N_4432,N_998,N_1419);
nor U4433 (N_4433,N_1114,N_430);
xor U4434 (N_4434,N_1894,N_941);
and U4435 (N_4435,N_101,N_1811);
nor U4436 (N_4436,N_1534,N_1487);
nand U4437 (N_4437,N_179,N_268);
or U4438 (N_4438,N_1408,N_2246);
and U4439 (N_4439,N_1704,N_1091);
nand U4440 (N_4440,N_955,N_339);
nand U4441 (N_4441,N_66,N_2303);
nand U4442 (N_4442,N_1390,N_103);
and U4443 (N_4443,N_1411,N_2382);
nor U4444 (N_4444,N_158,N_543);
and U4445 (N_4445,N_1568,N_679);
nand U4446 (N_4446,N_116,N_1673);
and U4447 (N_4447,N_2398,N_1043);
or U4448 (N_4448,N_2292,N_640);
nor U4449 (N_4449,N_408,N_1266);
and U4450 (N_4450,N_1083,N_2332);
nor U4451 (N_4451,N_2092,N_2498);
or U4452 (N_4452,N_1555,N_828);
or U4453 (N_4453,N_1814,N_1099);
or U4454 (N_4454,N_1389,N_551);
and U4455 (N_4455,N_2099,N_1136);
nor U4456 (N_4456,N_6,N_404);
or U4457 (N_4457,N_155,N_2463);
nor U4458 (N_4458,N_314,N_1575);
and U4459 (N_4459,N_1846,N_1537);
or U4460 (N_4460,N_2489,N_880);
nand U4461 (N_4461,N_1433,N_373);
nand U4462 (N_4462,N_2470,N_1324);
nor U4463 (N_4463,N_511,N_898);
nand U4464 (N_4464,N_1577,N_645);
and U4465 (N_4465,N_1984,N_8);
or U4466 (N_4466,N_2357,N_2459);
or U4467 (N_4467,N_1164,N_93);
nand U4468 (N_4468,N_1075,N_2166);
nor U4469 (N_4469,N_2139,N_479);
or U4470 (N_4470,N_1486,N_822);
and U4471 (N_4471,N_1246,N_2408);
nor U4472 (N_4472,N_1980,N_1045);
and U4473 (N_4473,N_1450,N_791);
nor U4474 (N_4474,N_2186,N_1600);
nand U4475 (N_4475,N_1333,N_1224);
and U4476 (N_4476,N_57,N_5);
xnor U4477 (N_4477,N_1356,N_1967);
nand U4478 (N_4478,N_1073,N_603);
nand U4479 (N_4479,N_8,N_2423);
nand U4480 (N_4480,N_1018,N_1020);
or U4481 (N_4481,N_121,N_322);
nand U4482 (N_4482,N_2139,N_490);
or U4483 (N_4483,N_1774,N_2218);
nand U4484 (N_4484,N_1039,N_1918);
nor U4485 (N_4485,N_50,N_1787);
nor U4486 (N_4486,N_183,N_1103);
nor U4487 (N_4487,N_928,N_1202);
or U4488 (N_4488,N_991,N_876);
and U4489 (N_4489,N_675,N_642);
nand U4490 (N_4490,N_85,N_1580);
or U4491 (N_4491,N_2278,N_1296);
nand U4492 (N_4492,N_809,N_191);
xnor U4493 (N_4493,N_574,N_2327);
and U4494 (N_4494,N_728,N_1501);
or U4495 (N_4495,N_195,N_263);
nor U4496 (N_4496,N_503,N_320);
nand U4497 (N_4497,N_2049,N_302);
and U4498 (N_4498,N_1922,N_1506);
nor U4499 (N_4499,N_2447,N_196);
nand U4500 (N_4500,N_362,N_1091);
and U4501 (N_4501,N_1840,N_346);
nor U4502 (N_4502,N_1121,N_1696);
nor U4503 (N_4503,N_2084,N_955);
and U4504 (N_4504,N_1845,N_1565);
nor U4505 (N_4505,N_571,N_1135);
and U4506 (N_4506,N_1055,N_2216);
or U4507 (N_4507,N_1531,N_850);
nor U4508 (N_4508,N_322,N_1794);
or U4509 (N_4509,N_197,N_421);
nor U4510 (N_4510,N_2335,N_2333);
nand U4511 (N_4511,N_1393,N_40);
and U4512 (N_4512,N_678,N_171);
or U4513 (N_4513,N_512,N_204);
nand U4514 (N_4514,N_359,N_789);
nand U4515 (N_4515,N_2048,N_631);
nand U4516 (N_4516,N_1169,N_1425);
or U4517 (N_4517,N_1025,N_153);
nor U4518 (N_4518,N_1748,N_1189);
or U4519 (N_4519,N_1827,N_896);
nand U4520 (N_4520,N_1744,N_826);
nor U4521 (N_4521,N_1544,N_2005);
nand U4522 (N_4522,N_1850,N_2497);
nand U4523 (N_4523,N_840,N_728);
nor U4524 (N_4524,N_1715,N_516);
nor U4525 (N_4525,N_1875,N_317);
nor U4526 (N_4526,N_948,N_1977);
or U4527 (N_4527,N_2324,N_886);
nand U4528 (N_4528,N_942,N_39);
nor U4529 (N_4529,N_480,N_2483);
nor U4530 (N_4530,N_1245,N_342);
nand U4531 (N_4531,N_241,N_1778);
nand U4532 (N_4532,N_886,N_1127);
or U4533 (N_4533,N_2112,N_830);
nand U4534 (N_4534,N_241,N_1651);
or U4535 (N_4535,N_1487,N_1709);
xor U4536 (N_4536,N_2154,N_276);
nor U4537 (N_4537,N_363,N_540);
and U4538 (N_4538,N_2032,N_86);
or U4539 (N_4539,N_253,N_423);
nand U4540 (N_4540,N_1399,N_566);
nor U4541 (N_4541,N_78,N_1889);
or U4542 (N_4542,N_1989,N_1252);
or U4543 (N_4543,N_1537,N_262);
nor U4544 (N_4544,N_1721,N_2000);
and U4545 (N_4545,N_427,N_1597);
and U4546 (N_4546,N_81,N_1497);
nor U4547 (N_4547,N_2432,N_1417);
and U4548 (N_4548,N_1481,N_849);
xor U4549 (N_4549,N_949,N_1969);
xor U4550 (N_4550,N_796,N_344);
nor U4551 (N_4551,N_1722,N_462);
nand U4552 (N_4552,N_606,N_2189);
or U4553 (N_4553,N_246,N_171);
nor U4554 (N_4554,N_668,N_548);
or U4555 (N_4555,N_69,N_1347);
nor U4556 (N_4556,N_2152,N_817);
and U4557 (N_4557,N_766,N_996);
and U4558 (N_4558,N_395,N_997);
and U4559 (N_4559,N_1026,N_1233);
and U4560 (N_4560,N_2175,N_1227);
and U4561 (N_4561,N_2404,N_1004);
nor U4562 (N_4562,N_2101,N_435);
nor U4563 (N_4563,N_437,N_1782);
nor U4564 (N_4564,N_868,N_532);
and U4565 (N_4565,N_1692,N_2335);
or U4566 (N_4566,N_439,N_1197);
nand U4567 (N_4567,N_242,N_29);
or U4568 (N_4568,N_1397,N_1313);
or U4569 (N_4569,N_983,N_210);
nand U4570 (N_4570,N_1208,N_757);
nand U4571 (N_4571,N_1067,N_469);
nor U4572 (N_4572,N_963,N_1376);
and U4573 (N_4573,N_464,N_1749);
nor U4574 (N_4574,N_1918,N_525);
nor U4575 (N_4575,N_1191,N_2418);
nor U4576 (N_4576,N_1481,N_1380);
and U4577 (N_4577,N_1633,N_1937);
nand U4578 (N_4578,N_1232,N_404);
and U4579 (N_4579,N_44,N_976);
nor U4580 (N_4580,N_404,N_528);
nor U4581 (N_4581,N_1973,N_2038);
nor U4582 (N_4582,N_733,N_916);
nor U4583 (N_4583,N_1645,N_382);
and U4584 (N_4584,N_1292,N_1116);
nand U4585 (N_4585,N_1897,N_1469);
and U4586 (N_4586,N_2356,N_756);
nand U4587 (N_4587,N_1237,N_2141);
or U4588 (N_4588,N_2101,N_2244);
or U4589 (N_4589,N_857,N_488);
and U4590 (N_4590,N_111,N_2452);
nand U4591 (N_4591,N_323,N_933);
nor U4592 (N_4592,N_629,N_2027);
and U4593 (N_4593,N_1932,N_1350);
nor U4594 (N_4594,N_37,N_1233);
or U4595 (N_4595,N_1221,N_2375);
and U4596 (N_4596,N_1701,N_906);
or U4597 (N_4597,N_987,N_1143);
and U4598 (N_4598,N_884,N_315);
nand U4599 (N_4599,N_1397,N_2);
nor U4600 (N_4600,N_755,N_496);
nor U4601 (N_4601,N_2111,N_1086);
or U4602 (N_4602,N_1960,N_2);
or U4603 (N_4603,N_651,N_1888);
nor U4604 (N_4604,N_2224,N_545);
nor U4605 (N_4605,N_982,N_79);
nand U4606 (N_4606,N_1591,N_1904);
nor U4607 (N_4607,N_1144,N_1969);
nor U4608 (N_4608,N_1473,N_314);
and U4609 (N_4609,N_1746,N_621);
or U4610 (N_4610,N_621,N_2203);
nand U4611 (N_4611,N_197,N_1281);
xor U4612 (N_4612,N_2261,N_1156);
nand U4613 (N_4613,N_280,N_2107);
and U4614 (N_4614,N_1917,N_1106);
nor U4615 (N_4615,N_1366,N_1035);
or U4616 (N_4616,N_120,N_1009);
nor U4617 (N_4617,N_1522,N_2183);
nor U4618 (N_4618,N_1949,N_1559);
nor U4619 (N_4619,N_2362,N_1076);
or U4620 (N_4620,N_504,N_111);
nand U4621 (N_4621,N_798,N_66);
and U4622 (N_4622,N_1706,N_453);
or U4623 (N_4623,N_1631,N_146);
xnor U4624 (N_4624,N_1465,N_2212);
and U4625 (N_4625,N_1973,N_1406);
nand U4626 (N_4626,N_2082,N_1179);
nor U4627 (N_4627,N_1479,N_506);
and U4628 (N_4628,N_84,N_258);
nor U4629 (N_4629,N_165,N_1621);
or U4630 (N_4630,N_65,N_2301);
and U4631 (N_4631,N_1514,N_431);
and U4632 (N_4632,N_533,N_2359);
nand U4633 (N_4633,N_1922,N_2014);
xnor U4634 (N_4634,N_1617,N_1908);
nand U4635 (N_4635,N_1907,N_11);
or U4636 (N_4636,N_2258,N_1426);
or U4637 (N_4637,N_1759,N_507);
or U4638 (N_4638,N_656,N_1801);
and U4639 (N_4639,N_539,N_2295);
nand U4640 (N_4640,N_2255,N_92);
nor U4641 (N_4641,N_2298,N_226);
or U4642 (N_4642,N_2424,N_1003);
and U4643 (N_4643,N_1417,N_1290);
nand U4644 (N_4644,N_517,N_2468);
nand U4645 (N_4645,N_980,N_2407);
and U4646 (N_4646,N_1120,N_267);
or U4647 (N_4647,N_1149,N_2206);
or U4648 (N_4648,N_2419,N_1498);
nand U4649 (N_4649,N_1178,N_1360);
nand U4650 (N_4650,N_699,N_591);
xor U4651 (N_4651,N_501,N_2083);
nand U4652 (N_4652,N_1819,N_646);
and U4653 (N_4653,N_1026,N_602);
or U4654 (N_4654,N_2081,N_88);
nand U4655 (N_4655,N_682,N_530);
nor U4656 (N_4656,N_1773,N_202);
nand U4657 (N_4657,N_2061,N_1827);
nand U4658 (N_4658,N_216,N_88);
or U4659 (N_4659,N_1826,N_1524);
and U4660 (N_4660,N_389,N_1168);
and U4661 (N_4661,N_1973,N_686);
nand U4662 (N_4662,N_520,N_2263);
nor U4663 (N_4663,N_2199,N_1711);
and U4664 (N_4664,N_506,N_496);
nor U4665 (N_4665,N_2223,N_884);
and U4666 (N_4666,N_158,N_763);
nand U4667 (N_4667,N_1111,N_211);
and U4668 (N_4668,N_1175,N_1332);
xnor U4669 (N_4669,N_1688,N_816);
nor U4670 (N_4670,N_2085,N_666);
nor U4671 (N_4671,N_1557,N_1014);
or U4672 (N_4672,N_2301,N_1243);
or U4673 (N_4673,N_326,N_1599);
or U4674 (N_4674,N_2184,N_2137);
or U4675 (N_4675,N_1027,N_1229);
and U4676 (N_4676,N_1661,N_2344);
and U4677 (N_4677,N_1212,N_353);
xnor U4678 (N_4678,N_810,N_1609);
or U4679 (N_4679,N_2477,N_1370);
nand U4680 (N_4680,N_1962,N_1244);
and U4681 (N_4681,N_2353,N_1849);
and U4682 (N_4682,N_311,N_1795);
nor U4683 (N_4683,N_1503,N_1343);
nand U4684 (N_4684,N_2324,N_1740);
nor U4685 (N_4685,N_1893,N_1066);
nand U4686 (N_4686,N_252,N_1250);
nand U4687 (N_4687,N_393,N_1090);
nor U4688 (N_4688,N_961,N_1252);
or U4689 (N_4689,N_2037,N_2093);
or U4690 (N_4690,N_2229,N_828);
nor U4691 (N_4691,N_707,N_212);
nand U4692 (N_4692,N_2128,N_744);
or U4693 (N_4693,N_562,N_1208);
or U4694 (N_4694,N_390,N_1629);
and U4695 (N_4695,N_2131,N_33);
or U4696 (N_4696,N_314,N_1137);
or U4697 (N_4697,N_1562,N_2392);
and U4698 (N_4698,N_2,N_1865);
or U4699 (N_4699,N_68,N_1407);
and U4700 (N_4700,N_734,N_989);
or U4701 (N_4701,N_1149,N_2268);
nand U4702 (N_4702,N_2435,N_2266);
or U4703 (N_4703,N_541,N_1141);
and U4704 (N_4704,N_466,N_1764);
nand U4705 (N_4705,N_2424,N_2012);
and U4706 (N_4706,N_1223,N_2419);
nor U4707 (N_4707,N_91,N_2357);
nand U4708 (N_4708,N_1296,N_2009);
nand U4709 (N_4709,N_863,N_542);
nor U4710 (N_4710,N_1118,N_554);
and U4711 (N_4711,N_804,N_1848);
and U4712 (N_4712,N_1595,N_1026);
or U4713 (N_4713,N_1542,N_601);
and U4714 (N_4714,N_1831,N_1941);
and U4715 (N_4715,N_781,N_1067);
xnor U4716 (N_4716,N_2290,N_2234);
or U4717 (N_4717,N_450,N_929);
nor U4718 (N_4718,N_2441,N_1505);
or U4719 (N_4719,N_2490,N_341);
or U4720 (N_4720,N_2433,N_566);
or U4721 (N_4721,N_14,N_775);
or U4722 (N_4722,N_857,N_88);
and U4723 (N_4723,N_696,N_820);
and U4724 (N_4724,N_67,N_2057);
nand U4725 (N_4725,N_853,N_963);
nor U4726 (N_4726,N_2014,N_911);
nand U4727 (N_4727,N_1114,N_1954);
nand U4728 (N_4728,N_132,N_1497);
nand U4729 (N_4729,N_556,N_162);
nand U4730 (N_4730,N_2311,N_1993);
and U4731 (N_4731,N_1308,N_2036);
and U4732 (N_4732,N_1925,N_2005);
nand U4733 (N_4733,N_892,N_252);
nand U4734 (N_4734,N_2182,N_248);
nor U4735 (N_4735,N_247,N_889);
nor U4736 (N_4736,N_1149,N_1406);
and U4737 (N_4737,N_1293,N_1729);
or U4738 (N_4738,N_20,N_2050);
nand U4739 (N_4739,N_1149,N_1008);
nor U4740 (N_4740,N_1951,N_764);
nor U4741 (N_4741,N_2052,N_780);
nand U4742 (N_4742,N_1139,N_20);
and U4743 (N_4743,N_1708,N_1680);
nor U4744 (N_4744,N_504,N_1753);
or U4745 (N_4745,N_617,N_537);
nor U4746 (N_4746,N_1091,N_1184);
or U4747 (N_4747,N_1103,N_1676);
and U4748 (N_4748,N_1424,N_2472);
nor U4749 (N_4749,N_1983,N_1445);
nand U4750 (N_4750,N_1907,N_511);
nor U4751 (N_4751,N_2430,N_441);
or U4752 (N_4752,N_1197,N_1782);
nor U4753 (N_4753,N_500,N_302);
nand U4754 (N_4754,N_741,N_251);
or U4755 (N_4755,N_666,N_314);
nand U4756 (N_4756,N_1659,N_935);
nand U4757 (N_4757,N_774,N_423);
nand U4758 (N_4758,N_1731,N_2323);
nor U4759 (N_4759,N_1637,N_746);
and U4760 (N_4760,N_7,N_1943);
and U4761 (N_4761,N_475,N_742);
nor U4762 (N_4762,N_148,N_149);
and U4763 (N_4763,N_694,N_734);
nand U4764 (N_4764,N_1935,N_59);
nand U4765 (N_4765,N_2323,N_1582);
and U4766 (N_4766,N_513,N_1150);
or U4767 (N_4767,N_1415,N_446);
xnor U4768 (N_4768,N_1189,N_2391);
nand U4769 (N_4769,N_2253,N_1129);
and U4770 (N_4770,N_322,N_417);
and U4771 (N_4771,N_1173,N_2165);
or U4772 (N_4772,N_627,N_2041);
nand U4773 (N_4773,N_813,N_2394);
or U4774 (N_4774,N_41,N_1004);
and U4775 (N_4775,N_1353,N_1829);
xnor U4776 (N_4776,N_1489,N_2162);
nand U4777 (N_4777,N_1170,N_1399);
nor U4778 (N_4778,N_2138,N_1902);
nand U4779 (N_4779,N_27,N_1108);
nor U4780 (N_4780,N_2158,N_214);
and U4781 (N_4781,N_1567,N_1833);
nand U4782 (N_4782,N_578,N_1553);
nand U4783 (N_4783,N_423,N_951);
and U4784 (N_4784,N_651,N_1800);
and U4785 (N_4785,N_696,N_631);
nor U4786 (N_4786,N_234,N_1871);
or U4787 (N_4787,N_2476,N_796);
and U4788 (N_4788,N_79,N_150);
nor U4789 (N_4789,N_123,N_207);
nor U4790 (N_4790,N_312,N_1012);
or U4791 (N_4791,N_1363,N_626);
nand U4792 (N_4792,N_1199,N_967);
or U4793 (N_4793,N_885,N_554);
or U4794 (N_4794,N_1783,N_1075);
nor U4795 (N_4795,N_401,N_52);
nand U4796 (N_4796,N_79,N_792);
nor U4797 (N_4797,N_536,N_2486);
xnor U4798 (N_4798,N_2429,N_420);
or U4799 (N_4799,N_2397,N_565);
or U4800 (N_4800,N_1367,N_71);
nand U4801 (N_4801,N_1551,N_1075);
nor U4802 (N_4802,N_1260,N_2002);
and U4803 (N_4803,N_2311,N_1553);
nor U4804 (N_4804,N_2040,N_1581);
and U4805 (N_4805,N_1160,N_1334);
nand U4806 (N_4806,N_1212,N_1624);
nor U4807 (N_4807,N_127,N_2228);
nor U4808 (N_4808,N_2163,N_785);
and U4809 (N_4809,N_1224,N_1182);
nand U4810 (N_4810,N_2323,N_1786);
and U4811 (N_4811,N_2423,N_2060);
and U4812 (N_4812,N_760,N_882);
or U4813 (N_4813,N_301,N_534);
nor U4814 (N_4814,N_1698,N_1238);
or U4815 (N_4815,N_468,N_718);
or U4816 (N_4816,N_1822,N_1444);
or U4817 (N_4817,N_854,N_670);
nor U4818 (N_4818,N_479,N_490);
and U4819 (N_4819,N_1235,N_1369);
and U4820 (N_4820,N_98,N_667);
nand U4821 (N_4821,N_1557,N_1950);
or U4822 (N_4822,N_2159,N_1734);
nor U4823 (N_4823,N_1366,N_1252);
nand U4824 (N_4824,N_621,N_794);
and U4825 (N_4825,N_885,N_475);
nand U4826 (N_4826,N_1709,N_1255);
nor U4827 (N_4827,N_397,N_1405);
nand U4828 (N_4828,N_471,N_969);
nor U4829 (N_4829,N_276,N_1578);
nor U4830 (N_4830,N_1257,N_440);
or U4831 (N_4831,N_1849,N_1825);
or U4832 (N_4832,N_685,N_1856);
or U4833 (N_4833,N_155,N_745);
nor U4834 (N_4834,N_170,N_6);
nor U4835 (N_4835,N_242,N_1429);
nor U4836 (N_4836,N_1327,N_604);
nor U4837 (N_4837,N_1918,N_1658);
nor U4838 (N_4838,N_2408,N_27);
or U4839 (N_4839,N_211,N_502);
and U4840 (N_4840,N_1337,N_562);
nand U4841 (N_4841,N_70,N_1879);
or U4842 (N_4842,N_1296,N_2006);
nand U4843 (N_4843,N_674,N_1364);
nor U4844 (N_4844,N_108,N_1084);
nor U4845 (N_4845,N_434,N_1086);
nand U4846 (N_4846,N_306,N_936);
nand U4847 (N_4847,N_1878,N_1791);
nand U4848 (N_4848,N_288,N_1680);
and U4849 (N_4849,N_1149,N_524);
nor U4850 (N_4850,N_651,N_2217);
nand U4851 (N_4851,N_2277,N_2371);
nand U4852 (N_4852,N_1933,N_1808);
and U4853 (N_4853,N_2065,N_93);
nor U4854 (N_4854,N_170,N_1276);
nor U4855 (N_4855,N_957,N_2299);
and U4856 (N_4856,N_949,N_1199);
xor U4857 (N_4857,N_2007,N_2465);
nand U4858 (N_4858,N_2256,N_2157);
nor U4859 (N_4859,N_2183,N_1459);
nand U4860 (N_4860,N_2393,N_220);
nor U4861 (N_4861,N_1746,N_1935);
and U4862 (N_4862,N_603,N_719);
nor U4863 (N_4863,N_1422,N_1230);
xor U4864 (N_4864,N_1709,N_1501);
nor U4865 (N_4865,N_1144,N_1470);
or U4866 (N_4866,N_1826,N_743);
and U4867 (N_4867,N_578,N_1965);
or U4868 (N_4868,N_2238,N_603);
and U4869 (N_4869,N_216,N_2220);
and U4870 (N_4870,N_1458,N_1526);
and U4871 (N_4871,N_942,N_704);
and U4872 (N_4872,N_1321,N_2367);
or U4873 (N_4873,N_2319,N_628);
nor U4874 (N_4874,N_1323,N_1997);
nand U4875 (N_4875,N_2138,N_2348);
or U4876 (N_4876,N_1737,N_1712);
or U4877 (N_4877,N_418,N_468);
nor U4878 (N_4878,N_2429,N_1242);
or U4879 (N_4879,N_1259,N_1657);
or U4880 (N_4880,N_257,N_1274);
nand U4881 (N_4881,N_1088,N_1401);
or U4882 (N_4882,N_1363,N_554);
and U4883 (N_4883,N_845,N_1383);
nand U4884 (N_4884,N_2481,N_1919);
and U4885 (N_4885,N_1096,N_2129);
nor U4886 (N_4886,N_1958,N_965);
nor U4887 (N_4887,N_1406,N_155);
or U4888 (N_4888,N_2262,N_697);
nor U4889 (N_4889,N_1562,N_482);
and U4890 (N_4890,N_49,N_1062);
nand U4891 (N_4891,N_1647,N_1383);
nor U4892 (N_4892,N_9,N_687);
and U4893 (N_4893,N_1125,N_1913);
or U4894 (N_4894,N_2293,N_545);
nand U4895 (N_4895,N_2457,N_594);
and U4896 (N_4896,N_55,N_387);
or U4897 (N_4897,N_1649,N_59);
or U4898 (N_4898,N_522,N_2385);
nor U4899 (N_4899,N_30,N_780);
and U4900 (N_4900,N_1719,N_1523);
nand U4901 (N_4901,N_1295,N_67);
or U4902 (N_4902,N_163,N_1320);
and U4903 (N_4903,N_2445,N_1744);
nand U4904 (N_4904,N_885,N_1000);
nor U4905 (N_4905,N_2317,N_161);
nand U4906 (N_4906,N_2485,N_1892);
nand U4907 (N_4907,N_743,N_2210);
xnor U4908 (N_4908,N_1360,N_956);
and U4909 (N_4909,N_1583,N_1379);
nand U4910 (N_4910,N_1345,N_1880);
and U4911 (N_4911,N_290,N_1207);
and U4912 (N_4912,N_440,N_1687);
nor U4913 (N_4913,N_23,N_2053);
nor U4914 (N_4914,N_1196,N_2464);
and U4915 (N_4915,N_605,N_2437);
or U4916 (N_4916,N_1191,N_246);
nor U4917 (N_4917,N_1428,N_2461);
or U4918 (N_4918,N_2396,N_1857);
nor U4919 (N_4919,N_1936,N_1914);
xor U4920 (N_4920,N_1860,N_2309);
and U4921 (N_4921,N_1772,N_370);
or U4922 (N_4922,N_789,N_1985);
nand U4923 (N_4923,N_1389,N_1331);
and U4924 (N_4924,N_679,N_233);
nor U4925 (N_4925,N_1135,N_384);
nand U4926 (N_4926,N_1327,N_820);
nand U4927 (N_4927,N_739,N_503);
nand U4928 (N_4928,N_1473,N_1698);
nor U4929 (N_4929,N_1951,N_1526);
and U4930 (N_4930,N_1915,N_1427);
nand U4931 (N_4931,N_1181,N_718);
and U4932 (N_4932,N_2453,N_1888);
and U4933 (N_4933,N_652,N_875);
nor U4934 (N_4934,N_2440,N_1147);
and U4935 (N_4935,N_684,N_1047);
or U4936 (N_4936,N_1737,N_617);
xnor U4937 (N_4937,N_2432,N_2458);
nand U4938 (N_4938,N_386,N_806);
and U4939 (N_4939,N_2425,N_153);
nor U4940 (N_4940,N_2275,N_919);
nand U4941 (N_4941,N_678,N_2068);
nand U4942 (N_4942,N_2038,N_2475);
or U4943 (N_4943,N_1959,N_1014);
nand U4944 (N_4944,N_49,N_1763);
nand U4945 (N_4945,N_1589,N_1924);
nor U4946 (N_4946,N_1564,N_1665);
or U4947 (N_4947,N_666,N_2302);
nor U4948 (N_4948,N_1924,N_892);
nor U4949 (N_4949,N_363,N_1870);
xnor U4950 (N_4950,N_2086,N_216);
nand U4951 (N_4951,N_2407,N_1063);
or U4952 (N_4952,N_316,N_1318);
and U4953 (N_4953,N_58,N_645);
nor U4954 (N_4954,N_216,N_1176);
nand U4955 (N_4955,N_1144,N_1750);
or U4956 (N_4956,N_1431,N_2237);
nor U4957 (N_4957,N_767,N_399);
or U4958 (N_4958,N_854,N_1765);
or U4959 (N_4959,N_1169,N_282);
or U4960 (N_4960,N_1187,N_2470);
and U4961 (N_4961,N_192,N_1699);
nor U4962 (N_4962,N_644,N_2180);
xnor U4963 (N_4963,N_1863,N_2454);
and U4964 (N_4964,N_518,N_909);
nand U4965 (N_4965,N_2169,N_566);
or U4966 (N_4966,N_963,N_2122);
nor U4967 (N_4967,N_1853,N_1916);
or U4968 (N_4968,N_182,N_1352);
or U4969 (N_4969,N_669,N_2103);
nor U4970 (N_4970,N_102,N_155);
nor U4971 (N_4971,N_340,N_1368);
or U4972 (N_4972,N_1152,N_1220);
nor U4973 (N_4973,N_1781,N_1859);
nand U4974 (N_4974,N_1329,N_2355);
nand U4975 (N_4975,N_1765,N_896);
nor U4976 (N_4976,N_1161,N_1884);
and U4977 (N_4977,N_1122,N_112);
xnor U4978 (N_4978,N_895,N_1965);
and U4979 (N_4979,N_771,N_2142);
nor U4980 (N_4980,N_921,N_2112);
or U4981 (N_4981,N_169,N_1641);
or U4982 (N_4982,N_1181,N_583);
and U4983 (N_4983,N_1175,N_1322);
or U4984 (N_4984,N_995,N_2261);
nand U4985 (N_4985,N_1746,N_824);
or U4986 (N_4986,N_1805,N_923);
or U4987 (N_4987,N_769,N_2414);
nand U4988 (N_4988,N_90,N_159);
and U4989 (N_4989,N_2341,N_2345);
nor U4990 (N_4990,N_1088,N_1302);
nor U4991 (N_4991,N_396,N_1507);
nor U4992 (N_4992,N_1300,N_1938);
and U4993 (N_4993,N_1893,N_1577);
nand U4994 (N_4994,N_2467,N_348);
or U4995 (N_4995,N_2057,N_1352);
or U4996 (N_4996,N_886,N_2415);
nand U4997 (N_4997,N_227,N_2432);
and U4998 (N_4998,N_1161,N_2329);
and U4999 (N_4999,N_247,N_48);
nor UO_0 (O_0,N_3974,N_4415);
and UO_1 (O_1,N_4966,N_3120);
nand UO_2 (O_2,N_2736,N_2691);
nor UO_3 (O_3,N_3505,N_4329);
or UO_4 (O_4,N_2939,N_2554);
nor UO_5 (O_5,N_2873,N_3725);
nor UO_6 (O_6,N_4811,N_4783);
nor UO_7 (O_7,N_4094,N_3957);
or UO_8 (O_8,N_3526,N_2847);
or UO_9 (O_9,N_4342,N_4921);
nor UO_10 (O_10,N_2611,N_2539);
or UO_11 (O_11,N_4799,N_2890);
nor UO_12 (O_12,N_2858,N_3027);
and UO_13 (O_13,N_4028,N_4324);
and UO_14 (O_14,N_4067,N_4795);
and UO_15 (O_15,N_4830,N_3155);
or UO_16 (O_16,N_4241,N_3828);
nor UO_17 (O_17,N_4167,N_4176);
and UO_18 (O_18,N_4612,N_4846);
and UO_19 (O_19,N_3646,N_4299);
xor UO_20 (O_20,N_4956,N_4598);
or UO_21 (O_21,N_4654,N_3482);
nor UO_22 (O_22,N_3296,N_2943);
nand UO_23 (O_23,N_4767,N_2948);
or UO_24 (O_24,N_4924,N_4222);
nor UO_25 (O_25,N_3060,N_2738);
nand UO_26 (O_26,N_4904,N_3950);
nand UO_27 (O_27,N_4080,N_3406);
and UO_28 (O_28,N_3879,N_3223);
and UO_29 (O_29,N_4820,N_3121);
nand UO_30 (O_30,N_4705,N_3412);
nand UO_31 (O_31,N_3608,N_2813);
nor UO_32 (O_32,N_3560,N_4488);
nor UO_33 (O_33,N_2696,N_2788);
nand UO_34 (O_34,N_2766,N_4644);
nand UO_35 (O_35,N_4351,N_3034);
nor UO_36 (O_36,N_4456,N_4447);
or UO_37 (O_37,N_4817,N_2532);
nor UO_38 (O_38,N_4962,N_3038);
nand UO_39 (O_39,N_4778,N_3249);
or UO_40 (O_40,N_4601,N_4064);
or UO_41 (O_41,N_4932,N_4847);
or UO_42 (O_42,N_4596,N_3492);
or UO_43 (O_43,N_4261,N_3645);
nor UO_44 (O_44,N_3726,N_3306);
nand UO_45 (O_45,N_4347,N_4215);
and UO_46 (O_46,N_3358,N_3594);
and UO_47 (O_47,N_4075,N_4511);
nor UO_48 (O_48,N_2885,N_3317);
or UO_49 (O_49,N_2763,N_4423);
and UO_50 (O_50,N_3260,N_3294);
nor UO_51 (O_51,N_3618,N_4066);
and UO_52 (O_52,N_3593,N_4667);
nand UO_53 (O_53,N_4520,N_4406);
nor UO_54 (O_54,N_3079,N_2872);
nor UO_55 (O_55,N_3510,N_4315);
and UO_56 (O_56,N_2869,N_4231);
and UO_57 (O_57,N_3805,N_4056);
nor UO_58 (O_58,N_4117,N_4508);
nor UO_59 (O_59,N_2855,N_3227);
or UO_60 (O_60,N_3046,N_3763);
or UO_61 (O_61,N_4336,N_4137);
or UO_62 (O_62,N_4002,N_3365);
nand UO_63 (O_63,N_4732,N_3384);
nand UO_64 (O_64,N_3813,N_4602);
and UO_65 (O_65,N_4513,N_4053);
and UO_66 (O_66,N_4760,N_4302);
nand UO_67 (O_67,N_4655,N_4380);
or UO_68 (O_68,N_3232,N_3414);
nor UO_69 (O_69,N_3032,N_3019);
nor UO_70 (O_70,N_3037,N_2723);
and UO_71 (O_71,N_3135,N_3164);
or UO_72 (O_72,N_4910,N_2961);
nor UO_73 (O_73,N_2588,N_3975);
or UO_74 (O_74,N_3273,N_4071);
nand UO_75 (O_75,N_3859,N_3627);
and UO_76 (O_76,N_4111,N_3539);
and UO_77 (O_77,N_2936,N_3044);
or UO_78 (O_78,N_2623,N_4410);
nor UO_79 (O_79,N_3811,N_2684);
nand UO_80 (O_80,N_4819,N_3866);
nor UO_81 (O_81,N_4686,N_3577);
nor UO_82 (O_82,N_2982,N_4776);
nand UO_83 (O_83,N_3587,N_3104);
or UO_84 (O_84,N_2553,N_4041);
nor UO_85 (O_85,N_4116,N_3968);
and UO_86 (O_86,N_2514,N_2903);
and UO_87 (O_87,N_2945,N_4313);
nor UO_88 (O_88,N_3520,N_3054);
nand UO_89 (O_89,N_3008,N_3491);
nand UO_90 (O_90,N_4568,N_3782);
nor UO_91 (O_91,N_3875,N_4985);
nand UO_92 (O_92,N_3422,N_3377);
xnor UO_93 (O_93,N_4519,N_4739);
nand UO_94 (O_94,N_2632,N_4195);
nor UO_95 (O_95,N_2547,N_2528);
nand UO_96 (O_96,N_4566,N_3711);
or UO_97 (O_97,N_3573,N_3623);
nor UO_98 (O_98,N_3238,N_3600);
xor UO_99 (O_99,N_3247,N_2821);
nand UO_100 (O_100,N_4281,N_2545);
or UO_101 (O_101,N_3115,N_3518);
nor UO_102 (O_102,N_4247,N_4707);
or UO_103 (O_103,N_4844,N_3258);
or UO_104 (O_104,N_2543,N_4092);
and UO_105 (O_105,N_3014,N_2867);
or UO_106 (O_106,N_4301,N_4079);
and UO_107 (O_107,N_4934,N_3500);
nor UO_108 (O_108,N_4688,N_4367);
nor UO_109 (O_109,N_4128,N_3373);
or UO_110 (O_110,N_4422,N_4227);
nor UO_111 (O_111,N_3001,N_3960);
nor UO_112 (O_112,N_4768,N_4164);
and UO_113 (O_113,N_2977,N_3277);
nor UO_114 (O_114,N_3648,N_3332);
nand UO_115 (O_115,N_3061,N_2621);
nor UO_116 (O_116,N_2914,N_4753);
and UO_117 (O_117,N_2831,N_2930);
nor UO_118 (O_118,N_2560,N_3980);
nand UO_119 (O_119,N_2871,N_4123);
and UO_120 (O_120,N_2768,N_3088);
or UO_121 (O_121,N_3166,N_4528);
nand UO_122 (O_122,N_2718,N_4316);
or UO_123 (O_123,N_3031,N_4493);
nor UO_124 (O_124,N_3567,N_3991);
and UO_125 (O_125,N_2591,N_4933);
or UO_126 (O_126,N_4983,N_3884);
xnor UO_127 (O_127,N_2619,N_3267);
or UO_128 (O_128,N_3657,N_4622);
or UO_129 (O_129,N_3056,N_3440);
nor UO_130 (O_130,N_3216,N_4177);
and UO_131 (O_131,N_3714,N_4288);
nor UO_132 (O_132,N_3281,N_3443);
nor UO_133 (O_133,N_2909,N_3681);
and UO_134 (O_134,N_2779,N_4480);
and UO_135 (O_135,N_4032,N_4818);
nand UO_136 (O_136,N_4014,N_3192);
and UO_137 (O_137,N_3552,N_2842);
or UO_138 (O_138,N_3301,N_4061);
or UO_139 (O_139,N_4475,N_3767);
and UO_140 (O_140,N_4201,N_3636);
nand UO_141 (O_141,N_3769,N_4341);
nor UO_142 (O_142,N_4702,N_2668);
nor UO_143 (O_143,N_2968,N_4802);
or UO_144 (O_144,N_3770,N_4798);
nand UO_145 (O_145,N_4597,N_2710);
or UO_146 (O_146,N_4431,N_4681);
or UO_147 (O_147,N_4614,N_3890);
and UO_148 (O_148,N_4698,N_2992);
nor UO_149 (O_149,N_2824,N_3671);
and UO_150 (O_150,N_3621,N_4990);
nor UO_151 (O_151,N_4455,N_4991);
nor UO_152 (O_152,N_3269,N_4547);
or UO_153 (O_153,N_3210,N_3125);
nand UO_154 (O_154,N_3291,N_2829);
and UO_155 (O_155,N_4893,N_2857);
nand UO_156 (O_156,N_4399,N_3638);
or UO_157 (O_157,N_3602,N_3868);
nand UO_158 (O_158,N_4146,N_4112);
nand UO_159 (O_159,N_4463,N_3918);
nand UO_160 (O_160,N_2570,N_3394);
xnor UO_161 (O_161,N_3119,N_4861);
nor UO_162 (O_162,N_4354,N_3603);
or UO_163 (O_163,N_3605,N_4348);
nor UO_164 (O_164,N_4282,N_4362);
or UO_165 (O_165,N_3945,N_4546);
nor UO_166 (O_166,N_2937,N_4570);
nor UO_167 (O_167,N_3521,N_3156);
nand UO_168 (O_168,N_3551,N_2530);
nand UO_169 (O_169,N_3760,N_4259);
and UO_170 (O_170,N_4544,N_2845);
nand UO_171 (O_171,N_3367,N_2986);
and UO_172 (O_172,N_4805,N_3795);
nand UO_173 (O_173,N_2783,N_4787);
nand UO_174 (O_174,N_3855,N_4314);
and UO_175 (O_175,N_4900,N_3504);
nand UO_176 (O_176,N_2908,N_3272);
or UO_177 (O_177,N_3972,N_2957);
nand UO_178 (O_178,N_3761,N_4938);
and UO_179 (O_179,N_4086,N_2878);
and UO_180 (O_180,N_3624,N_4665);
or UO_181 (O_181,N_2946,N_3882);
or UO_182 (O_182,N_2834,N_3207);
nand UO_183 (O_183,N_2714,N_3176);
nand UO_184 (O_184,N_4200,N_2955);
or UO_185 (O_185,N_3589,N_4063);
or UO_186 (O_186,N_4803,N_4782);
or UO_187 (O_187,N_4697,N_3397);
or UO_188 (O_188,N_3004,N_3344);
and UO_189 (O_189,N_2804,N_3766);
or UO_190 (O_190,N_2671,N_4572);
nor UO_191 (O_191,N_4838,N_3922);
nand UO_192 (O_192,N_2523,N_2994);
and UO_193 (O_193,N_2549,N_3508);
or UO_194 (O_194,N_2507,N_3123);
nor UO_195 (O_195,N_3029,N_4538);
and UO_196 (O_196,N_3640,N_4930);
or UO_197 (O_197,N_3303,N_3310);
nor UO_198 (O_198,N_3821,N_4621);
nor UO_199 (O_199,N_3529,N_3279);
nor UO_200 (O_200,N_2649,N_4349);
or UO_201 (O_201,N_2505,N_2854);
nor UO_202 (O_202,N_4865,N_4890);
nand UO_203 (O_203,N_3730,N_2984);
xor UO_204 (O_204,N_3152,N_4756);
nor UO_205 (O_205,N_4545,N_4451);
and UO_206 (O_206,N_4228,N_4434);
or UO_207 (O_207,N_2600,N_4175);
nor UO_208 (O_208,N_4543,N_2748);
nor UO_209 (O_209,N_3992,N_2525);
nor UO_210 (O_210,N_4393,N_4718);
or UO_211 (O_211,N_4187,N_2574);
nor UO_212 (O_212,N_2615,N_2983);
or UO_213 (O_213,N_3878,N_3998);
or UO_214 (O_214,N_3949,N_4155);
and UO_215 (O_215,N_3351,N_3467);
or UO_216 (O_216,N_3611,N_4611);
or UO_217 (O_217,N_4280,N_3804);
or UO_218 (O_218,N_2865,N_3647);
and UO_219 (O_219,N_2593,N_3665);
and UO_220 (O_220,N_2848,N_3011);
or UO_221 (O_221,N_4391,N_3886);
or UO_222 (O_222,N_3951,N_2771);
nor UO_223 (O_223,N_4486,N_4344);
or UO_224 (O_224,N_4026,N_4083);
nand UO_225 (O_225,N_3653,N_3101);
or UO_226 (O_226,N_3385,N_3025);
nand UO_227 (O_227,N_4427,N_3146);
nor UO_228 (O_228,N_2860,N_3224);
nor UO_229 (O_229,N_3134,N_4124);
xor UO_230 (O_230,N_4189,N_3336);
or UO_231 (O_231,N_3528,N_3843);
or UO_232 (O_232,N_2596,N_4859);
and UO_233 (O_233,N_4323,N_4340);
nand UO_234 (O_234,N_2966,N_4481);
nor UO_235 (O_235,N_4791,N_3196);
or UO_236 (O_236,N_4877,N_3092);
and UO_237 (O_237,N_4180,N_3969);
xnor UO_238 (O_238,N_3087,N_4318);
nor UO_239 (O_239,N_3654,N_4672);
nand UO_240 (O_240,N_3486,N_3757);
or UO_241 (O_241,N_4095,N_3783);
nand UO_242 (O_242,N_2603,N_4696);
and UO_243 (O_243,N_4551,N_4330);
nor UO_244 (O_244,N_4521,N_4120);
and UO_245 (O_245,N_4425,N_4633);
and UO_246 (O_246,N_4326,N_4430);
xor UO_247 (O_247,N_3892,N_4557);
or UO_248 (O_248,N_4653,N_4800);
nand UO_249 (O_249,N_4514,N_2733);
and UO_250 (O_250,N_3180,N_2729);
nand UO_251 (O_251,N_2500,N_2660);
or UO_252 (O_252,N_4131,N_4610);
nand UO_253 (O_253,N_3905,N_4274);
nand UO_254 (O_254,N_4375,N_2636);
nor UO_255 (O_255,N_4309,N_3077);
nand UO_256 (O_256,N_2790,N_2690);
nand UO_257 (O_257,N_4049,N_4635);
or UO_258 (O_258,N_4870,N_4722);
nor UO_259 (O_259,N_2713,N_3755);
nor UO_260 (O_260,N_3117,N_3075);
nor UO_261 (O_261,N_3245,N_4392);
and UO_262 (O_262,N_4219,N_4279);
nor UO_263 (O_263,N_2998,N_3449);
or UO_264 (O_264,N_4068,N_2546);
nor UO_265 (O_265,N_3873,N_3280);
nor UO_266 (O_266,N_4306,N_4003);
or UO_267 (O_267,N_2663,N_3062);
nor UO_268 (O_268,N_4715,N_4660);
nor UO_269 (O_269,N_4874,N_4343);
nand UO_270 (O_270,N_3168,N_4937);
nor UO_271 (O_271,N_4101,N_3354);
nor UO_272 (O_272,N_2695,N_3114);
or UO_273 (O_273,N_4136,N_4173);
or UO_274 (O_274,N_4770,N_4054);
and UO_275 (O_275,N_4065,N_4673);
nand UO_276 (O_276,N_3097,N_4959);
nor UO_277 (O_277,N_3253,N_3173);
nor UO_278 (O_278,N_4225,N_3561);
or UO_279 (O_279,N_3836,N_3124);
nand UO_280 (O_280,N_4439,N_2898);
nor UO_281 (O_281,N_3523,N_4213);
nor UO_282 (O_282,N_2562,N_2659);
or UO_283 (O_283,N_2996,N_3667);
nor UO_284 (O_284,N_4594,N_2652);
or UO_285 (O_285,N_3017,N_2888);
or UO_286 (O_286,N_4998,N_2664);
and UO_287 (O_287,N_3986,N_3582);
nand UO_288 (O_288,N_4823,N_3468);
nand UO_289 (O_289,N_2777,N_4211);
nand UO_290 (O_290,N_2760,N_4492);
and UO_291 (O_291,N_3463,N_2958);
nor UO_292 (O_292,N_4897,N_3675);
nor UO_293 (O_293,N_4505,N_4454);
and UO_294 (O_294,N_4992,N_2662);
nand UO_295 (O_295,N_4581,N_3359);
nor UO_296 (O_296,N_4471,N_3182);
and UO_297 (O_297,N_4942,N_4152);
and UO_298 (O_298,N_3243,N_4007);
nand UO_299 (O_299,N_3133,N_3501);
and UO_300 (O_300,N_3773,N_2877);
nand UO_301 (O_301,N_3137,N_3987);
or UO_302 (O_302,N_4742,N_3352);
nand UO_303 (O_303,N_4015,N_4230);
and UO_304 (O_304,N_3544,N_2745);
and UO_305 (O_305,N_2923,N_3093);
and UO_306 (O_306,N_4361,N_3787);
and UO_307 (O_307,N_3802,N_4853);
or UO_308 (O_308,N_3939,N_4084);
and UO_309 (O_309,N_2624,N_4449);
or UO_310 (O_310,N_4031,N_4987);
nor UO_311 (O_311,N_4262,N_3459);
and UO_312 (O_312,N_2558,N_3664);
and UO_313 (O_313,N_4950,N_4055);
or UO_314 (O_314,N_4412,N_4307);
or UO_315 (O_315,N_3314,N_4501);
and UO_316 (O_316,N_2902,N_3241);
nand UO_317 (O_317,N_2730,N_3053);
or UO_318 (O_318,N_4927,N_2602);
and UO_319 (O_319,N_4769,N_3254);
and UO_320 (O_320,N_4902,N_4019);
nand UO_321 (O_321,N_3448,N_4321);
and UO_322 (O_322,N_3865,N_3424);
nor UO_323 (O_323,N_3826,N_4181);
xor UO_324 (O_324,N_4011,N_3993);
nand UO_325 (O_325,N_4935,N_3512);
or UO_326 (O_326,N_3111,N_3396);
or UO_327 (O_327,N_4358,N_4695);
nand UO_328 (O_328,N_2702,N_3465);
nand UO_329 (O_329,N_3403,N_3211);
and UO_330 (O_330,N_3801,N_3700);
or UO_331 (O_331,N_4503,N_4303);
nand UO_332 (O_332,N_3215,N_3067);
and UO_333 (O_333,N_4468,N_3081);
nand UO_334 (O_334,N_2985,N_3432);
and UO_335 (O_335,N_3708,N_3010);
or UO_336 (O_336,N_2751,N_4266);
xor UO_337 (O_337,N_4196,N_4331);
or UO_338 (O_338,N_3806,N_4628);
nor UO_339 (O_339,N_3680,N_3609);
or UO_340 (O_340,N_3765,N_4372);
or UO_341 (O_341,N_4154,N_3113);
and UO_342 (O_342,N_3926,N_2816);
or UO_343 (O_343,N_3153,N_4394);
nor UO_344 (O_344,N_4277,N_4138);
and UO_345 (O_345,N_4774,N_3862);
nor UO_346 (O_346,N_4560,N_3419);
and UO_347 (O_347,N_3065,N_3474);
nor UO_348 (O_348,N_4483,N_2764);
or UO_349 (O_349,N_2917,N_4567);
and UO_350 (O_350,N_4467,N_4452);
or UO_351 (O_351,N_3817,N_4518);
and UO_352 (O_352,N_3920,N_3222);
nand UO_353 (O_353,N_3469,N_2541);
or UO_354 (O_354,N_4150,N_4580);
or UO_355 (O_355,N_2817,N_4246);
and UO_356 (O_356,N_2578,N_3533);
or UO_357 (O_357,N_2724,N_3874);
or UO_358 (O_358,N_3679,N_4831);
or UO_359 (O_359,N_4139,N_3786);
and UO_360 (O_360,N_3042,N_2604);
or UO_361 (O_361,N_2920,N_4460);
or UO_362 (O_362,N_3887,N_4143);
and UO_363 (O_363,N_2642,N_4104);
nand UO_364 (O_364,N_4147,N_3891);
nand UO_365 (O_365,N_4158,N_4165);
xnor UO_366 (O_366,N_4305,N_2884);
and UO_367 (O_367,N_4988,N_2526);
and UO_368 (O_368,N_2993,N_4417);
and UO_369 (O_369,N_3024,N_3558);
xor UO_370 (O_370,N_2653,N_2509);
and UO_371 (O_371,N_3083,N_3547);
or UO_372 (O_372,N_3590,N_4775);
nand UO_373 (O_373,N_4490,N_4419);
or UO_374 (O_374,N_2667,N_3845);
and UO_375 (O_375,N_3178,N_4121);
nor UO_376 (O_376,N_3018,N_4796);
nand UO_377 (O_377,N_4841,N_3230);
nor UO_378 (O_378,N_3712,N_3256);
and UO_379 (O_379,N_4656,N_4733);
and UO_380 (O_380,N_2823,N_3462);
or UO_381 (O_381,N_4583,N_4012);
nor UO_382 (O_382,N_3292,N_3692);
nand UO_383 (O_383,N_3952,N_3488);
and UO_384 (O_384,N_2896,N_2540);
and UO_385 (O_385,N_4886,N_4944);
nor UO_386 (O_386,N_2866,N_3194);
and UO_387 (O_387,N_2677,N_3933);
nor UO_388 (O_388,N_4171,N_4346);
and UO_389 (O_389,N_4085,N_2536);
and UO_390 (O_390,N_3059,N_4864);
nand UO_391 (O_391,N_3823,N_4388);
nor UO_392 (O_392,N_2537,N_3250);
nand UO_393 (O_393,N_4701,N_2670);
and UO_394 (O_394,N_3722,N_3154);
nor UO_395 (O_395,N_2681,N_3997);
nand UO_396 (O_396,N_4203,N_4887);
and UO_397 (O_397,N_3342,N_4446);
nand UO_398 (O_398,N_2907,N_2595);
nand UO_399 (O_399,N_4951,N_2682);
nor UO_400 (O_400,N_4076,N_3822);
nor UO_401 (O_401,N_2801,N_3005);
nor UO_402 (O_402,N_4917,N_4814);
nand UO_403 (O_403,N_4297,N_4214);
xor UO_404 (O_404,N_2956,N_4995);
or UO_405 (O_405,N_3350,N_4828);
nand UO_406 (O_406,N_3564,N_4478);
and UO_407 (O_407,N_3793,N_2592);
or UO_408 (O_408,N_3842,N_2886);
nand UO_409 (O_409,N_3048,N_3497);
nand UO_410 (O_410,N_4194,N_3290);
or UO_411 (O_411,N_3282,N_3321);
or UO_412 (O_412,N_4573,N_2527);
or UO_413 (O_413,N_3055,N_3747);
nor UO_414 (O_414,N_3699,N_3378);
nor UO_415 (O_415,N_3411,N_4191);
or UO_416 (O_416,N_2963,N_4706);
and UO_417 (O_417,N_3953,N_3549);
nor UO_418 (O_418,N_4727,N_4857);
nand UO_419 (O_419,N_4954,N_4920);
nor UO_420 (O_420,N_3548,N_2731);
and UO_421 (O_421,N_4709,N_2556);
nand UO_422 (O_422,N_4107,N_4249);
or UO_423 (O_423,N_3779,N_3399);
or UO_424 (O_424,N_4042,N_3913);
nand UO_425 (O_425,N_4023,N_3357);
or UO_426 (O_426,N_2940,N_3401);
xor UO_427 (O_427,N_4140,N_2775);
nand UO_428 (O_428,N_2597,N_2915);
nor UO_429 (O_429,N_3184,N_3928);
nor UO_430 (O_430,N_3930,N_3837);
nand UO_431 (O_431,N_3327,N_3644);
or UO_432 (O_432,N_4098,N_4289);
and UO_433 (O_433,N_4445,N_4794);
and UO_434 (O_434,N_4849,N_4502);
or UO_435 (O_435,N_3142,N_2876);
xor UO_436 (O_436,N_4789,N_4074);
nand UO_437 (O_437,N_2564,N_4848);
and UO_438 (O_438,N_3346,N_4365);
or UO_439 (O_439,N_4729,N_2705);
nand UO_440 (O_440,N_4025,N_3353);
nor UO_441 (O_441,N_4437,N_3479);
and UO_442 (O_442,N_4273,N_3737);
and UO_443 (O_443,N_3237,N_2538);
and UO_444 (O_444,N_3487,N_4464);
and UO_445 (O_445,N_2792,N_3880);
and UO_446 (O_446,N_4947,N_4276);
and UO_447 (O_447,N_4532,N_3455);
and UO_448 (O_448,N_2565,N_3546);
nand UO_449 (O_449,N_4980,N_3555);
or UO_450 (O_450,N_4397,N_2828);
nand UO_451 (O_451,N_4089,N_4713);
or UO_452 (O_452,N_3407,N_3226);
nand UO_453 (O_453,N_3139,N_2735);
or UO_454 (O_454,N_4837,N_4009);
nand UO_455 (O_455,N_4650,N_3617);
or UO_456 (O_456,N_3200,N_4691);
nand UO_457 (O_457,N_2795,N_2997);
or UO_458 (O_458,N_4197,N_2778);
nor UO_459 (O_459,N_4047,N_2544);
nand UO_460 (O_460,N_4843,N_3400);
and UO_461 (O_461,N_2913,N_2614);
or UO_462 (O_462,N_2762,N_2927);
nor UO_463 (O_463,N_3068,N_4979);
or UO_464 (O_464,N_4716,N_2933);
nor UO_465 (O_465,N_3601,N_3295);
nor UO_466 (O_466,N_3867,N_3752);
nor UO_467 (O_467,N_4370,N_3105);
nor UO_468 (O_468,N_4278,N_2513);
nand UO_469 (O_469,N_3535,N_3219);
nand UO_470 (O_470,N_3495,N_4148);
nand UO_471 (O_471,N_3450,N_4008);
nor UO_472 (O_472,N_4300,N_3808);
xor UO_473 (O_473,N_4271,N_3186);
nand UO_474 (O_474,N_2687,N_4448);
nor UO_475 (O_475,N_3484,N_3231);
or UO_476 (O_476,N_3002,N_2807);
nand UO_477 (O_477,N_3515,N_2517);
or UO_478 (O_478,N_4466,N_2949);
nand UO_479 (O_479,N_3356,N_3911);
nor UO_480 (O_480,N_3047,N_4443);
and UO_481 (O_481,N_4190,N_3089);
and UO_482 (O_482,N_3160,N_3333);
nand UO_483 (O_483,N_4804,N_4440);
or UO_484 (O_484,N_2765,N_4498);
nor UO_485 (O_485,N_3792,N_3530);
or UO_486 (O_486,N_3943,N_4287);
nand UO_487 (O_487,N_3509,N_3251);
or UO_488 (O_488,N_4122,N_4905);
and UO_489 (O_489,N_2754,N_4634);
nor UO_490 (O_490,N_2594,N_3218);
and UO_491 (O_491,N_4668,N_4687);
and UO_492 (O_492,N_3883,N_4582);
nor UO_493 (O_493,N_4052,N_3283);
and UO_494 (O_494,N_4949,N_2893);
nand UO_495 (O_495,N_3662,N_2605);
or UO_496 (O_496,N_3374,N_4678);
and UO_497 (O_497,N_2931,N_2572);
or UO_498 (O_498,N_3935,N_3850);
nor UO_499 (O_499,N_4510,N_2625);
or UO_500 (O_500,N_4723,N_2925);
nand UO_501 (O_501,N_3041,N_3299);
and UO_502 (O_502,N_4110,N_2542);
nor UO_503 (O_503,N_4345,N_4226);
nor UO_504 (O_504,N_2550,N_2964);
and UO_505 (O_505,N_3191,N_4377);
nand UO_506 (O_506,N_2969,N_3717);
or UO_507 (O_507,N_3217,N_4381);
or UO_508 (O_508,N_4777,N_2694);
nor UO_509 (O_509,N_2515,N_4353);
xor UO_510 (O_510,N_4491,N_3753);
and UO_511 (O_511,N_4958,N_4875);
and UO_512 (O_512,N_2656,N_4790);
and UO_513 (O_513,N_2628,N_3461);
or UO_514 (O_514,N_4710,N_4507);
and UO_515 (O_515,N_2512,N_2987);
or UO_516 (O_516,N_2567,N_4963);
nand UO_517 (O_517,N_3015,N_4442);
or UO_518 (O_518,N_3898,N_2938);
or UO_519 (O_519,N_2524,N_4252);
nand UO_520 (O_520,N_2599,N_3418);
and UO_521 (O_521,N_3996,N_3764);
and UO_522 (O_522,N_4239,N_3572);
nor UO_523 (O_523,N_2789,N_4641);
nor UO_524 (O_524,N_4379,N_4642);
or UO_525 (O_525,N_3684,N_3923);
nand UO_526 (O_526,N_2585,N_4224);
nand UO_527 (O_527,N_3472,N_4389);
nand UO_528 (O_528,N_3388,N_3470);
nor UO_529 (O_529,N_4587,N_4390);
nor UO_530 (O_530,N_2535,N_4363);
nor UO_531 (O_531,N_4311,N_4832);
nand UO_532 (O_532,N_2725,N_3661);
and UO_533 (O_533,N_4616,N_3563);
nand UO_534 (O_534,N_4773,N_2580);
and UO_535 (O_535,N_4270,N_3404);
nor UO_536 (O_536,N_4465,N_2839);
or UO_537 (O_537,N_3340,N_4118);
nand UO_538 (O_538,N_2786,N_4579);
nand UO_539 (O_539,N_3701,N_3261);
and UO_540 (O_540,N_4914,N_2846);
or UO_541 (O_541,N_3831,N_4036);
xor UO_542 (O_542,N_4936,N_2737);
or UO_543 (O_543,N_3174,N_4133);
or UO_544 (O_544,N_3566,N_2576);
nor UO_545 (O_545,N_2676,N_4470);
or UO_546 (O_546,N_4073,N_4901);
and UO_547 (O_547,N_3707,N_4512);
and UO_548 (O_548,N_4387,N_2887);
nor UO_549 (O_549,N_3538,N_2607);
nor UO_550 (O_550,N_3595,N_2981);
or UO_551 (O_551,N_2640,N_3426);
nand UO_552 (O_552,N_4048,N_3132);
nor UO_553 (O_553,N_3656,N_3480);
nand UO_554 (O_554,N_4113,N_2675);
or UO_555 (O_555,N_4613,N_2557);
and UO_556 (O_556,N_3846,N_4968);
nor UO_557 (O_557,N_3973,N_4267);
nand UO_558 (O_558,N_2655,N_2899);
nor UO_559 (O_559,N_3776,N_4125);
nand UO_560 (O_560,N_3622,N_4885);
nand UO_561 (O_561,N_4725,N_4754);
or UO_562 (O_562,N_3257,N_3395);
and UO_563 (O_563,N_3099,N_2785);
nor UO_564 (O_564,N_2750,N_4771);
or UO_565 (O_565,N_4542,N_3651);
nor UO_566 (O_566,N_4106,N_4529);
or UO_567 (O_567,N_2741,N_4720);
nand UO_568 (O_568,N_4728,N_3652);
or UO_569 (O_569,N_3541,N_3309);
and UO_570 (O_570,N_3734,N_4743);
or UO_571 (O_571,N_3057,N_3628);
or UO_572 (O_572,N_2551,N_3723);
and UO_573 (O_573,N_4097,N_4169);
nand UO_574 (O_574,N_3635,N_4420);
and UO_575 (O_575,N_3829,N_4620);
and UO_576 (O_576,N_2891,N_3167);
and UO_577 (O_577,N_3408,N_4556);
and UO_578 (O_578,N_3316,N_4473);
or UO_579 (O_579,N_4156,N_4711);
nand UO_580 (O_580,N_4590,N_3007);
and UO_581 (O_581,N_3863,N_4208);
or UO_582 (O_582,N_3127,N_2633);
or UO_583 (O_583,N_3931,N_2758);
nor UO_584 (O_584,N_3169,N_3550);
nand UO_585 (O_585,N_3876,N_4941);
and UO_586 (O_586,N_2721,N_4523);
nor UO_587 (O_587,N_2648,N_3921);
nand UO_588 (O_588,N_4731,N_4585);
or UO_589 (O_589,N_3586,N_3188);
nand UO_590 (O_590,N_4221,N_4919);
or UO_591 (O_591,N_3762,N_2833);
or UO_592 (O_592,N_4652,N_4404);
and UO_593 (O_593,N_3709,N_2797);
or UO_594 (O_594,N_3912,N_4599);
and UO_595 (O_595,N_3893,N_3064);
nor UO_596 (O_596,N_3434,N_2521);
nor UO_597 (O_597,N_2811,N_2861);
nand UO_598 (O_598,N_4779,N_3298);
nand UO_599 (O_599,N_3742,N_3300);
or UO_600 (O_600,N_4685,N_2503);
nor UO_601 (O_601,N_4976,N_4105);
nor UO_602 (O_602,N_3718,N_4090);
or UO_603 (O_603,N_4537,N_4703);
or UO_604 (O_604,N_2864,N_4734);
nand UO_605 (O_605,N_2919,N_4918);
and UO_606 (O_606,N_4748,N_4931);
and UO_607 (O_607,N_2688,N_4676);
nand UO_608 (O_608,N_4700,N_3958);
and UO_609 (O_609,N_3909,N_4099);
and UO_610 (O_610,N_3221,N_4157);
or UO_611 (O_611,N_2769,N_3275);
nor UO_612 (O_612,N_4825,N_4833);
or UO_613 (O_613,N_4100,N_3904);
nor UO_614 (O_614,N_3502,N_4842);
or UO_615 (O_615,N_4646,N_3570);
nand UO_616 (O_616,N_2838,N_4333);
nand UO_617 (O_617,N_4096,N_4626);
or UO_618 (O_618,N_3932,N_4884);
and UO_619 (O_619,N_3441,N_2643);
and UO_620 (O_620,N_4911,N_4264);
and UO_621 (O_621,N_4119,N_4269);
nand UO_622 (O_622,N_3691,N_3924);
or UO_623 (O_623,N_3305,N_4496);
and UO_624 (O_624,N_3239,N_3981);
or UO_625 (O_625,N_2941,N_2841);
nand UO_626 (O_626,N_4265,N_4970);
nand UO_627 (O_627,N_3743,N_4308);
and UO_628 (O_628,N_4174,N_4161);
nand UO_629 (O_629,N_2979,N_4232);
nand UO_630 (O_630,N_4967,N_4260);
and UO_631 (O_631,N_4216,N_2511);
nand UO_632 (O_632,N_3368,N_3990);
or UO_633 (O_633,N_3179,N_3849);
nand UO_634 (O_634,N_3234,N_4953);
nand UO_635 (O_635,N_2952,N_2835);
nor UO_636 (O_636,N_3071,N_4745);
or UO_637 (O_637,N_4737,N_2753);
or UO_638 (O_638,N_3051,N_4589);
nand UO_639 (O_639,N_3334,N_3816);
and UO_640 (O_640,N_4880,N_2679);
or UO_641 (O_641,N_3323,N_2965);
nor UO_642 (O_642,N_4070,N_3633);
or UO_643 (O_643,N_4724,N_4268);
and UO_644 (O_644,N_4746,N_2974);
nor UO_645 (O_645,N_3925,N_4516);
nand UO_646 (O_646,N_2851,N_2704);
and UO_647 (O_647,N_3897,N_3995);
nand UO_648 (O_648,N_3798,N_2683);
nand UO_649 (O_649,N_3319,N_4129);
or UO_650 (O_650,N_4891,N_3288);
nor UO_651 (O_651,N_3095,N_4898);
and UO_652 (O_652,N_4286,N_2720);
or UO_653 (O_653,N_3147,N_3255);
or UO_654 (O_654,N_3557,N_4531);
xnor UO_655 (O_655,N_3476,N_4982);
nand UO_656 (O_656,N_2999,N_2708);
nand UO_657 (O_657,N_3908,N_4021);
nor UO_658 (O_658,N_4233,N_2972);
nand UO_659 (O_659,N_4290,N_3989);
nor UO_660 (O_660,N_4712,N_4168);
xor UO_661 (O_661,N_2618,N_4955);
and UO_662 (O_662,N_3363,N_2579);
or UO_663 (O_663,N_3963,N_3190);
and UO_664 (O_664,N_3961,N_3165);
or UO_665 (O_665,N_3740,N_3023);
and UO_666 (O_666,N_4881,N_4744);
nor UO_667 (O_667,N_4645,N_2590);
nor UO_668 (O_668,N_3799,N_3181);
or UO_669 (O_669,N_3197,N_3466);
and UO_670 (O_670,N_3934,N_3626);
nand UO_671 (O_671,N_3382,N_4812);
or UO_672 (O_672,N_4945,N_4485);
and UO_673 (O_673,N_3750,N_2749);
or UO_674 (O_674,N_3129,N_2897);
nor UO_675 (O_675,N_3078,N_4396);
and UO_676 (O_676,N_4821,N_3732);
and UO_677 (O_677,N_3149,N_2650);
or UO_678 (O_678,N_3205,N_3438);
nand UO_679 (O_679,N_2853,N_3639);
and UO_680 (O_680,N_4206,N_3446);
or UO_681 (O_681,N_4664,N_3266);
or UO_682 (O_682,N_3437,N_4172);
and UO_683 (O_683,N_2988,N_2895);
or UO_684 (O_684,N_3794,N_3000);
and UO_685 (O_685,N_2814,N_2973);
nand UO_686 (O_686,N_3637,N_4552);
nand UO_687 (O_687,N_3335,N_3201);
xnor UO_688 (O_688,N_4912,N_4472);
or UO_689 (O_689,N_3430,N_4459);
nand UO_690 (O_690,N_4487,N_4996);
nand UO_691 (O_691,N_4735,N_4636);
and UO_692 (O_692,N_3927,N_4960);
and UO_693 (O_693,N_3150,N_2812);
nor UO_694 (O_694,N_4141,N_4671);
nand UO_695 (O_695,N_3503,N_3203);
nand UO_696 (O_696,N_2892,N_4093);
or UO_697 (O_697,N_3264,N_4127);
or UO_698 (O_698,N_4450,N_2569);
or UO_699 (O_699,N_3452,N_3971);
nor UO_700 (O_700,N_4526,N_3832);
xnor UO_701 (O_701,N_4704,N_3036);
nand UO_702 (O_702,N_2647,N_2971);
nand UO_703 (O_703,N_3676,N_4975);
or UO_704 (O_704,N_4786,N_2802);
and UO_705 (O_705,N_4913,N_3496);
nand UO_706 (O_706,N_4586,N_3263);
nor UO_707 (O_707,N_4403,N_3797);
and UO_708 (O_708,N_3527,N_4997);
and UO_709 (O_709,N_4198,N_3872);
nor UO_710 (O_710,N_3371,N_3917);
nand UO_711 (O_711,N_3364,N_3715);
and UO_712 (O_712,N_4682,N_2918);
nor UO_713 (O_713,N_4879,N_2799);
or UO_714 (O_714,N_4563,N_3881);
or UO_715 (O_715,N_3163,N_4750);
nand UO_716 (O_716,N_3612,N_3940);
or UO_717 (O_717,N_4909,N_2555);
and UO_718 (O_718,N_3630,N_3741);
nor UO_719 (O_719,N_4876,N_4438);
nand UO_720 (O_720,N_2706,N_4845);
or UO_721 (O_721,N_2630,N_4350);
and UO_722 (O_722,N_3944,N_2739);
nand UO_723 (O_723,N_2504,N_3728);
and UO_724 (O_724,N_2910,N_3574);
or UO_725 (O_725,N_3026,N_3244);
nand UO_726 (O_726,N_3293,N_3629);
and UO_727 (O_727,N_4250,N_4035);
nand UO_728 (O_728,N_4986,N_3965);
or UO_729 (O_729,N_4661,N_3756);
xor UO_730 (O_730,N_3442,N_4816);
nand UO_731 (O_731,N_4405,N_3851);
or UO_732 (O_732,N_2757,N_2862);
nor UO_733 (O_733,N_4525,N_4555);
nand UO_734 (O_734,N_3161,N_4327);
nor UO_735 (O_735,N_4535,N_4013);
nand UO_736 (O_736,N_2506,N_2743);
or UO_737 (O_737,N_4894,N_4638);
nor UO_738 (O_738,N_2502,N_3444);
nor UO_739 (O_739,N_4807,N_2755);
and UO_740 (O_740,N_3421,N_3458);
or UO_741 (O_741,N_3938,N_2672);
and UO_742 (O_742,N_4939,N_2586);
and UO_743 (O_743,N_4217,N_3387);
and UO_744 (O_744,N_4569,N_2522);
nor UO_745 (O_745,N_3206,N_4675);
nand UO_746 (O_746,N_4153,N_4145);
and UO_747 (O_747,N_4130,N_2612);
nor UO_748 (O_748,N_4030,N_3329);
or UO_749 (O_749,N_2870,N_4553);
and UO_750 (O_750,N_3607,N_4243);
and UO_751 (O_751,N_3807,N_2711);
nor UO_752 (O_752,N_2601,N_2674);
or UO_753 (O_753,N_2774,N_3956);
and UO_754 (O_754,N_3285,N_4373);
nand UO_755 (O_755,N_4595,N_2746);
and UO_756 (O_756,N_3604,N_4000);
and UO_757 (O_757,N_3331,N_4016);
and UO_758 (O_758,N_4436,N_3668);
nand UO_759 (O_759,N_4294,N_4761);
nor UO_760 (O_760,N_4193,N_4378);
or UO_761 (O_761,N_3641,N_4046);
nor UO_762 (O_762,N_4253,N_2796);
and UO_763 (O_763,N_2548,N_2803);
or UO_764 (O_764,N_4017,N_4801);
and UO_765 (O_765,N_4683,N_4809);
nand UO_766 (O_766,N_2707,N_4185);
or UO_767 (O_767,N_4044,N_3979);
nor UO_768 (O_768,N_4576,N_3268);
nor UO_769 (O_769,N_3785,N_3772);
nor UO_770 (O_770,N_3246,N_4310);
xor UO_771 (O_771,N_3361,N_4593);
nand UO_772 (O_772,N_3896,N_2552);
nand UO_773 (O_773,N_2699,N_3393);
nand UO_774 (O_774,N_3236,N_4630);
nor UO_775 (O_775,N_4540,N_4659);
nand UO_776 (O_776,N_2756,N_3524);
or UO_777 (O_777,N_4584,N_3126);
nand UO_778 (O_778,N_2881,N_4714);
nand UO_779 (O_779,N_4504,N_4335);
or UO_780 (O_780,N_4202,N_3016);
or UO_781 (O_781,N_3771,N_3252);
and UO_782 (O_782,N_3685,N_3514);
nand UO_783 (O_783,N_4670,N_3575);
nor UO_784 (O_784,N_4108,N_2742);
or UO_785 (O_785,N_3330,N_4522);
nand UO_786 (O_786,N_4517,N_3259);
or UO_787 (O_787,N_3284,N_4883);
nor UO_788 (O_788,N_3780,N_4248);
or UO_789 (O_789,N_4617,N_2905);
nand UO_790 (O_790,N_3349,N_2719);
nor UO_791 (O_791,N_3702,N_3228);
nor UO_792 (O_792,N_4283,N_3381);
nand UO_793 (O_793,N_3519,N_3947);
nand UO_794 (O_794,N_3220,N_3429);
xnor UO_795 (O_795,N_4400,N_4479);
and UO_796 (O_796,N_4666,N_3343);
or UO_797 (O_797,N_4441,N_3788);
nand UO_798 (O_798,N_4298,N_4548);
nand UO_799 (O_799,N_3848,N_4408);
nand UO_800 (O_800,N_3035,N_2990);
or UO_801 (O_801,N_3610,N_4304);
or UO_802 (O_802,N_3242,N_4296);
nor UO_803 (O_803,N_4050,N_3901);
or UO_804 (O_804,N_3326,N_3919);
and UO_805 (O_805,N_2722,N_4462);
nand UO_806 (O_806,N_3311,N_3490);
or UO_807 (O_807,N_2912,N_3634);
nor UO_808 (O_808,N_2646,N_4062);
nand UO_809 (O_809,N_2850,N_3907);
or UO_810 (O_810,N_2926,N_3672);
nand UO_811 (O_811,N_3337,N_3090);
nor UO_812 (O_812,N_2608,N_3148);
nand UO_813 (O_813,N_3106,N_3478);
nand UO_814 (O_814,N_4578,N_3839);
or UO_815 (O_815,N_3916,N_2916);
nand UO_816 (O_816,N_4603,N_4693);
or UO_817 (O_817,N_4730,N_3208);
and UO_818 (O_818,N_2716,N_4961);
nor UO_819 (O_819,N_3825,N_2822);
nand UO_820 (O_820,N_3143,N_4495);
nor UO_821 (O_821,N_3187,N_3858);
or UO_822 (O_822,N_2634,N_3043);
nor UO_823 (O_823,N_4813,N_3304);
nor UO_824 (O_824,N_3674,N_3122);
and UO_825 (O_825,N_4458,N_3988);
nor UO_826 (O_826,N_4418,N_3513);
nand UO_827 (O_827,N_4836,N_2950);
or UO_828 (O_828,N_4763,N_3431);
and UO_829 (O_829,N_3663,N_2928);
or UO_830 (O_830,N_3063,N_3483);
xor UO_831 (O_831,N_4364,N_3937);
nand UO_832 (O_832,N_4088,N_2673);
nor UO_833 (O_833,N_3983,N_4134);
and UO_834 (O_834,N_3435,N_2692);
nor UO_835 (O_835,N_4780,N_3499);
nand UO_836 (O_836,N_4662,N_2609);
nand UO_837 (O_837,N_3744,N_3009);
and UO_838 (O_838,N_3193,N_3006);
nor UO_839 (O_839,N_4592,N_4037);
nand UO_840 (O_840,N_3313,N_4132);
nor UO_841 (O_841,N_4020,N_3369);
xor UO_842 (O_842,N_3649,N_2840);
nor UO_843 (O_843,N_4322,N_3784);
nor UO_844 (O_844,N_2832,N_2734);
or UO_845 (O_845,N_2534,N_3375);
nor UO_846 (O_846,N_4368,N_4411);
nand UO_847 (O_847,N_3704,N_2631);
nor UO_848 (O_848,N_4317,N_3815);
nand UO_849 (O_849,N_3098,N_3141);
and UO_850 (O_850,N_3289,N_3597);
and UO_851 (O_851,N_4038,N_4109);
nor UO_852 (O_852,N_2680,N_2700);
or UO_853 (O_853,N_4989,N_3109);
or UO_854 (O_854,N_3451,N_4497);
nand UO_855 (O_855,N_3325,N_3844);
or UO_856 (O_856,N_3554,N_2651);
nor UO_857 (O_857,N_2820,N_2904);
and UO_858 (O_858,N_3235,N_3138);
nand UO_859 (O_859,N_4251,N_4205);
and UO_860 (O_860,N_3195,N_3977);
or UO_861 (O_861,N_4220,N_3835);
and UO_862 (O_862,N_3069,N_3172);
nor UO_863 (O_863,N_4810,N_4383);
and UO_864 (O_864,N_2805,N_3145);
nor UO_865 (O_865,N_2995,N_3360);
or UO_866 (O_866,N_4209,N_4469);
nor UO_867 (O_867,N_3716,N_4506);
nor UO_868 (O_868,N_3473,N_3003);
nand UO_869 (O_869,N_4059,N_2626);
or UO_870 (O_870,N_4792,N_3021);
nand UO_871 (O_871,N_2782,N_4385);
nand UO_872 (O_872,N_2951,N_3420);
nand UO_873 (O_873,N_3592,N_3903);
xnor UO_874 (O_874,N_3494,N_3144);
nor UO_875 (O_875,N_2901,N_4337);
and UO_876 (O_876,N_4669,N_2809);
and UO_877 (O_877,N_4229,N_2787);
nor UO_878 (O_878,N_2947,N_2583);
or UO_879 (O_879,N_3861,N_3489);
and UO_880 (O_880,N_3568,N_3889);
or UO_881 (O_881,N_3091,N_4965);
or UO_882 (O_882,N_2657,N_3959);
or UO_883 (O_883,N_3777,N_2967);
and UO_884 (O_884,N_2827,N_2613);
nand UO_885 (O_885,N_3380,N_3625);
or UO_886 (O_886,N_3820,N_2924);
or UO_887 (O_887,N_3103,N_4034);
or UO_888 (O_888,N_4332,N_3885);
nor UO_889 (O_889,N_4689,N_4272);
nor UO_890 (O_890,N_4444,N_4254);
nand UO_891 (O_891,N_3578,N_3894);
and UO_892 (O_892,N_2894,N_3070);
or UO_893 (O_893,N_3477,N_3240);
and UO_894 (O_894,N_3074,N_4946);
nand UO_895 (O_895,N_4407,N_3659);
or UO_896 (O_896,N_3454,N_2622);
and UO_897 (O_897,N_2727,N_4759);
nand UO_898 (O_898,N_4862,N_3941);
or UO_899 (O_899,N_3906,N_2844);
nor UO_900 (O_900,N_4291,N_2863);
and UO_901 (O_901,N_3151,N_4618);
or UO_902 (O_902,N_4574,N_2935);
nand UO_903 (O_903,N_4257,N_3372);
nand UO_904 (O_904,N_3398,N_4001);
and UO_905 (O_905,N_4639,N_4878);
and UO_906 (O_906,N_4210,N_4999);
and UO_907 (O_907,N_4677,N_3409);
nor UO_908 (O_908,N_4561,N_3703);
and UO_909 (O_909,N_3910,N_2929);
and UO_910 (O_910,N_3012,N_4087);
or UO_911 (O_911,N_3759,N_3410);
or UO_912 (O_912,N_3423,N_4741);
or UO_913 (O_913,N_3697,N_4562);
nor UO_914 (O_914,N_3198,N_3049);
nand UO_915 (O_915,N_4057,N_3225);
nand UO_916 (O_916,N_3613,N_4159);
nor UO_917 (O_917,N_3028,N_3976);
nor UO_918 (O_918,N_4923,N_3274);
and UO_919 (O_919,N_2669,N_4549);
or UO_920 (O_920,N_4785,N_4608);
nor UO_921 (O_921,N_3727,N_4840);
xnor UO_922 (O_922,N_4242,N_4974);
and UO_923 (O_923,N_4658,N_3402);
nor UO_924 (O_924,N_3569,N_3328);
and UO_925 (O_925,N_3158,N_3751);
and UO_926 (O_926,N_3076,N_3658);
and UO_927 (O_927,N_4624,N_3682);
or UO_928 (O_928,N_2516,N_2849);
nand UO_929 (O_929,N_2620,N_3545);
nand UO_930 (O_930,N_4461,N_3157);
nor UO_931 (O_931,N_3131,N_4747);
and UO_932 (O_932,N_3565,N_2856);
nor UO_933 (O_933,N_4915,N_2773);
and UO_934 (O_934,N_3112,N_3705);
or UO_935 (O_935,N_3745,N_2793);
nor UO_936 (O_936,N_4114,N_4721);
nand UO_937 (O_937,N_3599,N_3994);
and UO_938 (O_938,N_3942,N_4736);
and UO_939 (O_939,N_2911,N_4863);
nand UO_940 (O_940,N_3389,N_3775);
xnor UO_941 (O_941,N_4170,N_4888);
and UO_942 (O_942,N_4398,N_3096);
nor UO_943 (O_943,N_4952,N_3620);
or UO_944 (O_944,N_3082,N_4334);
nand UO_945 (O_945,N_4515,N_4489);
nand UO_946 (O_946,N_2875,N_3248);
nor UO_947 (O_947,N_3084,N_4929);
nand UO_948 (O_948,N_3655,N_4826);
nand UO_949 (O_949,N_2629,N_3212);
or UO_950 (O_950,N_3948,N_3128);
nand UO_951 (O_951,N_2962,N_3517);
and UO_952 (O_952,N_4925,N_3202);
nor UO_953 (O_953,N_3030,N_3140);
and UO_954 (O_954,N_4357,N_3347);
or UO_955 (O_955,N_2922,N_4188);
nand UO_956 (O_956,N_3308,N_3803);
and UO_957 (O_957,N_3736,N_4433);
or UO_958 (O_958,N_2654,N_3749);
and UO_959 (O_959,N_4027,N_2703);
and UO_960 (O_960,N_2818,N_4142);
xor UO_961 (O_961,N_2616,N_3580);
nand UO_962 (O_962,N_4069,N_3955);
nor UO_963 (O_963,N_3073,N_3052);
and UO_964 (O_964,N_3110,N_2666);
nand UO_965 (O_965,N_4366,N_4591);
or UO_966 (O_966,N_2880,N_3562);
or UO_967 (O_967,N_2533,N_4499);
nor UO_968 (O_968,N_3107,N_3386);
nand UO_969 (O_969,N_3457,N_4550);
or UO_970 (O_970,N_4244,N_3159);
nor UO_971 (O_971,N_3721,N_4356);
and UO_972 (O_972,N_2744,N_3020);
xnor UO_973 (O_973,N_3425,N_3338);
and UO_974 (O_974,N_3525,N_3687);
nand UO_975 (O_975,N_2510,N_4275);
and UO_976 (O_976,N_4186,N_2900);
and UO_977 (O_977,N_4872,N_4500);
nand UO_978 (O_978,N_3390,N_4149);
and UO_979 (O_979,N_3170,N_3966);
nor UO_980 (O_980,N_4477,N_2953);
and UO_981 (O_981,N_4292,N_4413);
and UO_982 (O_982,N_3040,N_4320);
nor UO_983 (O_983,N_4060,N_4039);
nand UO_984 (O_984,N_2584,N_4212);
and UO_985 (O_985,N_3914,N_4903);
nand UO_986 (O_986,N_3348,N_4964);
nor UO_987 (O_987,N_2581,N_3619);
nand UO_988 (O_988,N_3392,N_2798);
and UO_989 (O_989,N_4679,N_4829);
nand UO_990 (O_990,N_3177,N_3724);
and UO_991 (O_991,N_4627,N_4690);
and UO_992 (O_992,N_3870,N_3713);
nand UO_993 (O_993,N_4263,N_4435);
or UO_994 (O_994,N_4126,N_3962);
nor UO_995 (O_995,N_4866,N_3345);
nand UO_996 (O_996,N_2610,N_2689);
nand UO_997 (O_997,N_2732,N_3287);
and UO_998 (O_998,N_4637,N_3720);
or UO_999 (O_999,N_4033,N_4907);
endmodule