module basic_500_3000_500_6_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_475,In_69);
nand U1 (N_1,In_140,In_496);
and U2 (N_2,In_224,In_251);
xnor U3 (N_3,In_487,In_186);
xor U4 (N_4,In_486,In_248);
xor U5 (N_5,In_209,In_42);
nand U6 (N_6,In_219,In_371);
nor U7 (N_7,In_112,In_270);
or U8 (N_8,In_20,In_25);
or U9 (N_9,In_181,In_192);
nor U10 (N_10,In_234,In_163);
nor U11 (N_11,In_348,In_454);
and U12 (N_12,In_483,In_457);
nand U13 (N_13,In_471,In_214);
nand U14 (N_14,In_168,In_334);
nand U15 (N_15,In_262,In_32);
nand U16 (N_16,In_449,In_221);
or U17 (N_17,In_474,In_281);
nor U18 (N_18,In_161,In_398);
nor U19 (N_19,In_309,In_62);
and U20 (N_20,In_350,In_9);
or U21 (N_21,In_421,In_462);
and U22 (N_22,In_172,In_225);
nand U23 (N_23,In_19,In_440);
or U24 (N_24,In_66,In_28);
or U25 (N_25,In_217,In_109);
and U26 (N_26,In_282,In_443);
or U27 (N_27,In_170,In_324);
and U28 (N_28,In_263,In_469);
nand U29 (N_29,In_2,In_177);
nand U30 (N_30,In_293,In_272);
nand U31 (N_31,In_426,In_236);
or U32 (N_32,In_295,In_456);
nand U33 (N_33,In_299,In_461);
nor U34 (N_34,In_108,In_415);
and U35 (N_35,In_126,In_372);
or U36 (N_36,In_199,In_265);
or U37 (N_37,In_308,In_446);
or U38 (N_38,In_458,In_448);
nand U39 (N_39,In_169,In_97);
and U40 (N_40,In_329,In_478);
nor U41 (N_41,In_431,In_273);
nor U42 (N_42,In_476,In_365);
nor U43 (N_43,In_485,In_283);
nor U44 (N_44,In_325,In_271);
nor U45 (N_45,In_358,In_392);
and U46 (N_46,In_148,In_326);
nand U47 (N_47,In_274,In_4);
xor U48 (N_48,In_359,In_342);
and U49 (N_49,In_388,In_328);
and U50 (N_50,In_89,In_114);
or U51 (N_51,In_179,In_407);
nor U52 (N_52,In_226,In_497);
or U53 (N_53,In_285,In_304);
or U54 (N_54,In_400,In_178);
nor U55 (N_55,In_11,In_472);
nand U56 (N_56,In_246,In_164);
nor U57 (N_57,In_119,In_240);
and U58 (N_58,In_76,In_351);
xnor U59 (N_59,In_43,In_242);
and U60 (N_60,In_105,In_302);
or U61 (N_61,In_74,In_191);
or U62 (N_62,In_387,In_482);
nor U63 (N_63,In_215,In_316);
nand U64 (N_64,In_57,In_331);
xnor U65 (N_65,In_53,In_297);
nand U66 (N_66,In_85,In_205);
nor U67 (N_67,In_13,In_8);
or U68 (N_68,In_465,In_480);
or U69 (N_69,In_54,In_292);
nor U70 (N_70,In_238,In_174);
or U71 (N_71,In_55,In_175);
and U72 (N_72,In_202,In_127);
nor U73 (N_73,In_31,In_430);
nor U74 (N_74,In_152,In_40);
nand U75 (N_75,In_187,In_44);
nand U76 (N_76,In_210,In_362);
or U77 (N_77,In_154,In_7);
nand U78 (N_78,In_68,In_373);
nor U79 (N_79,In_58,In_417);
nand U80 (N_80,In_255,In_420);
nor U81 (N_81,In_452,In_190);
and U82 (N_82,In_307,In_88);
nor U83 (N_83,In_150,In_466);
xnor U84 (N_84,In_444,In_113);
or U85 (N_85,In_17,In_216);
nor U86 (N_86,In_142,In_418);
and U87 (N_87,In_137,In_123);
nor U88 (N_88,In_338,In_59);
nand U89 (N_89,In_312,In_185);
nor U90 (N_90,In_241,In_322);
nand U91 (N_91,In_39,In_481);
and U92 (N_92,In_367,In_197);
xor U93 (N_93,In_1,In_38);
xor U94 (N_94,In_343,In_162);
nand U95 (N_95,In_253,In_80);
nor U96 (N_96,In_499,In_239);
nor U97 (N_97,In_428,In_155);
and U98 (N_98,In_333,In_376);
and U99 (N_99,In_337,In_132);
nand U100 (N_100,In_353,In_451);
or U101 (N_101,In_135,In_455);
nor U102 (N_102,In_327,In_296);
or U103 (N_103,In_414,In_409);
or U104 (N_104,In_26,In_294);
and U105 (N_105,In_93,In_412);
nor U106 (N_106,In_442,In_259);
xnor U107 (N_107,In_361,In_346);
xnor U108 (N_108,In_211,In_498);
nand U109 (N_109,In_220,In_463);
and U110 (N_110,In_291,In_130);
nand U111 (N_111,In_491,In_196);
xor U112 (N_112,In_266,In_46);
nand U113 (N_113,In_336,In_35);
xor U114 (N_114,In_194,In_268);
or U115 (N_115,In_134,In_94);
nor U116 (N_116,In_22,In_52);
and U117 (N_117,In_419,In_206);
nand U118 (N_118,In_208,In_73);
and U119 (N_119,In_165,In_237);
and U120 (N_120,In_345,In_167);
or U121 (N_121,In_403,In_157);
and U122 (N_122,In_118,In_51);
or U123 (N_123,In_397,In_406);
or U124 (N_124,In_21,In_120);
nand U125 (N_125,In_101,In_385);
nor U126 (N_126,In_479,In_212);
and U127 (N_127,In_102,In_314);
and U128 (N_128,In_404,In_363);
nand U129 (N_129,In_231,In_258);
and U130 (N_130,In_171,In_50);
or U131 (N_131,In_233,In_413);
or U132 (N_132,In_48,In_61);
or U133 (N_133,In_67,In_98);
and U134 (N_134,In_184,In_131);
or U135 (N_135,In_193,In_484);
nor U136 (N_136,In_425,In_30);
nand U137 (N_137,In_432,In_111);
nand U138 (N_138,In_305,In_117);
nor U139 (N_139,In_427,In_422);
nand U140 (N_140,In_284,In_453);
and U141 (N_141,In_301,In_357);
nand U142 (N_142,In_235,In_144);
or U143 (N_143,In_34,In_278);
and U144 (N_144,In_122,In_12);
nand U145 (N_145,In_189,In_267);
or U146 (N_146,In_411,In_250);
or U147 (N_147,In_405,In_160);
or U148 (N_148,In_15,In_393);
and U149 (N_149,In_355,In_288);
nand U150 (N_150,In_96,In_276);
or U151 (N_151,In_201,In_408);
or U152 (N_152,In_203,In_64);
and U153 (N_153,In_396,In_245);
and U154 (N_154,In_222,In_213);
and U155 (N_155,In_423,In_341);
xnor U156 (N_156,In_390,In_92);
nor U157 (N_157,In_124,In_156);
or U158 (N_158,In_303,In_252);
xnor U159 (N_159,In_344,In_340);
nor U160 (N_160,In_493,In_286);
and U161 (N_161,In_0,In_149);
xor U162 (N_162,In_29,In_99);
nor U163 (N_163,In_488,In_10);
nor U164 (N_164,In_103,In_433);
xnor U165 (N_165,In_5,In_87);
or U166 (N_166,In_381,In_104);
xor U167 (N_167,In_438,In_72);
nor U168 (N_168,In_489,In_37);
nor U169 (N_169,In_468,In_159);
xnor U170 (N_170,In_3,In_230);
or U171 (N_171,In_287,In_82);
or U172 (N_172,In_429,In_339);
nor U173 (N_173,In_244,In_347);
nor U174 (N_174,In_24,In_391);
nand U175 (N_175,In_410,In_77);
nand U176 (N_176,In_153,In_352);
and U177 (N_177,In_386,In_145);
xor U178 (N_178,In_424,In_402);
xor U179 (N_179,In_477,In_204);
or U180 (N_180,In_289,In_116);
and U181 (N_181,In_133,In_147);
xnor U182 (N_182,In_495,In_378);
nor U183 (N_183,In_382,In_439);
nand U184 (N_184,In_264,In_173);
nor U185 (N_185,In_473,In_467);
or U186 (N_186,In_16,In_106);
or U187 (N_187,In_141,In_138);
nor U188 (N_188,In_257,In_47);
and U189 (N_189,In_182,In_136);
and U190 (N_190,In_490,In_260);
or U191 (N_191,In_279,In_261);
or U192 (N_192,In_311,In_23);
and U193 (N_193,In_354,In_166);
nor U194 (N_194,In_143,In_107);
nor U195 (N_195,In_366,In_115);
nor U196 (N_196,In_218,In_232);
and U197 (N_197,In_229,In_223);
nor U198 (N_198,In_280,In_277);
or U199 (N_199,In_56,In_86);
and U200 (N_200,In_375,In_14);
nand U201 (N_201,In_227,In_364);
nor U202 (N_202,In_349,In_450);
and U203 (N_203,In_33,In_436);
and U204 (N_204,In_18,In_79);
nor U205 (N_205,In_91,In_315);
and U206 (N_206,In_198,In_317);
nand U207 (N_207,In_395,In_41);
or U208 (N_208,In_319,In_243);
or U209 (N_209,In_60,In_383);
nand U210 (N_210,In_71,In_437);
nand U211 (N_211,In_183,In_389);
nor U212 (N_212,In_275,In_401);
nand U213 (N_213,In_464,In_313);
nand U214 (N_214,In_445,In_368);
nor U215 (N_215,In_176,In_256);
nor U216 (N_216,In_435,In_254);
and U217 (N_217,In_27,In_320);
or U218 (N_218,In_200,In_180);
or U219 (N_219,In_460,In_36);
nor U220 (N_220,In_441,In_49);
and U221 (N_221,In_300,In_310);
nand U222 (N_222,In_335,In_332);
nand U223 (N_223,In_434,In_63);
nand U224 (N_224,In_158,In_470);
or U225 (N_225,In_360,In_125);
nand U226 (N_226,In_269,In_83);
nor U227 (N_227,In_384,In_45);
nor U228 (N_228,In_380,In_65);
or U229 (N_229,In_139,In_399);
and U230 (N_230,In_306,In_330);
nand U231 (N_231,In_84,In_146);
nand U232 (N_232,In_6,In_494);
nand U233 (N_233,In_129,In_370);
and U234 (N_234,In_290,In_394);
nor U235 (N_235,In_369,In_416);
nand U236 (N_236,In_81,In_207);
or U237 (N_237,In_321,In_90);
nor U238 (N_238,In_379,In_195);
and U239 (N_239,In_356,In_249);
nand U240 (N_240,In_78,In_70);
nor U241 (N_241,In_121,In_188);
or U242 (N_242,In_377,In_323);
nor U243 (N_243,In_492,In_298);
and U244 (N_244,In_247,In_374);
nor U245 (N_245,In_459,In_447);
nand U246 (N_246,In_318,In_100);
or U247 (N_247,In_228,In_110);
and U248 (N_248,In_128,In_75);
or U249 (N_249,In_151,In_95);
nor U250 (N_250,In_494,In_169);
nor U251 (N_251,In_225,In_12);
and U252 (N_252,In_60,In_211);
nand U253 (N_253,In_73,In_299);
or U254 (N_254,In_271,In_159);
and U255 (N_255,In_462,In_296);
and U256 (N_256,In_78,In_389);
and U257 (N_257,In_371,In_260);
or U258 (N_258,In_87,In_177);
nand U259 (N_259,In_267,In_232);
xor U260 (N_260,In_490,In_252);
or U261 (N_261,In_79,In_459);
nor U262 (N_262,In_148,In_447);
nand U263 (N_263,In_445,In_481);
xor U264 (N_264,In_474,In_286);
nand U265 (N_265,In_296,In_463);
and U266 (N_266,In_360,In_494);
nand U267 (N_267,In_61,In_498);
nor U268 (N_268,In_257,In_464);
and U269 (N_269,In_153,In_401);
or U270 (N_270,In_222,In_460);
nand U271 (N_271,In_300,In_20);
nand U272 (N_272,In_3,In_167);
xnor U273 (N_273,In_94,In_341);
and U274 (N_274,In_154,In_341);
nand U275 (N_275,In_160,In_395);
and U276 (N_276,In_49,In_233);
or U277 (N_277,In_169,In_201);
and U278 (N_278,In_192,In_315);
and U279 (N_279,In_63,In_79);
nor U280 (N_280,In_215,In_438);
and U281 (N_281,In_205,In_297);
nand U282 (N_282,In_102,In_207);
nand U283 (N_283,In_461,In_79);
or U284 (N_284,In_293,In_352);
nand U285 (N_285,In_139,In_137);
nand U286 (N_286,In_174,In_391);
and U287 (N_287,In_297,In_89);
nor U288 (N_288,In_368,In_165);
or U289 (N_289,In_208,In_484);
nor U290 (N_290,In_336,In_379);
or U291 (N_291,In_86,In_483);
nand U292 (N_292,In_365,In_83);
nand U293 (N_293,In_261,In_217);
or U294 (N_294,In_349,In_430);
or U295 (N_295,In_75,In_125);
nor U296 (N_296,In_268,In_449);
and U297 (N_297,In_478,In_193);
or U298 (N_298,In_236,In_105);
or U299 (N_299,In_363,In_382);
or U300 (N_300,In_423,In_323);
nand U301 (N_301,In_417,In_222);
xnor U302 (N_302,In_284,In_411);
nand U303 (N_303,In_37,In_99);
and U304 (N_304,In_115,In_376);
and U305 (N_305,In_416,In_384);
and U306 (N_306,In_291,In_478);
nor U307 (N_307,In_432,In_28);
or U308 (N_308,In_193,In_153);
xnor U309 (N_309,In_148,In_298);
or U310 (N_310,In_0,In_480);
or U311 (N_311,In_174,In_261);
or U312 (N_312,In_473,In_272);
and U313 (N_313,In_82,In_21);
or U314 (N_314,In_116,In_154);
and U315 (N_315,In_77,In_457);
and U316 (N_316,In_410,In_147);
xor U317 (N_317,In_214,In_83);
nor U318 (N_318,In_134,In_408);
nand U319 (N_319,In_382,In_452);
nand U320 (N_320,In_27,In_348);
and U321 (N_321,In_419,In_293);
nand U322 (N_322,In_290,In_369);
and U323 (N_323,In_490,In_290);
and U324 (N_324,In_464,In_250);
or U325 (N_325,In_396,In_407);
nand U326 (N_326,In_253,In_52);
and U327 (N_327,In_92,In_353);
nand U328 (N_328,In_477,In_363);
or U329 (N_329,In_36,In_53);
xor U330 (N_330,In_320,In_385);
and U331 (N_331,In_294,In_20);
nor U332 (N_332,In_339,In_354);
xnor U333 (N_333,In_292,In_96);
or U334 (N_334,In_458,In_193);
nand U335 (N_335,In_113,In_189);
nor U336 (N_336,In_431,In_483);
nand U337 (N_337,In_375,In_267);
xor U338 (N_338,In_247,In_314);
and U339 (N_339,In_147,In_475);
or U340 (N_340,In_292,In_436);
and U341 (N_341,In_369,In_108);
and U342 (N_342,In_216,In_141);
and U343 (N_343,In_126,In_101);
nand U344 (N_344,In_415,In_113);
nand U345 (N_345,In_434,In_270);
or U346 (N_346,In_389,In_150);
nor U347 (N_347,In_307,In_191);
nand U348 (N_348,In_48,In_318);
or U349 (N_349,In_328,In_454);
and U350 (N_350,In_14,In_419);
and U351 (N_351,In_5,In_90);
nor U352 (N_352,In_103,In_169);
and U353 (N_353,In_322,In_154);
xnor U354 (N_354,In_474,In_431);
nor U355 (N_355,In_206,In_204);
and U356 (N_356,In_90,In_476);
and U357 (N_357,In_352,In_336);
or U358 (N_358,In_280,In_316);
nand U359 (N_359,In_410,In_48);
nor U360 (N_360,In_217,In_456);
nor U361 (N_361,In_275,In_372);
or U362 (N_362,In_407,In_206);
and U363 (N_363,In_155,In_219);
xnor U364 (N_364,In_276,In_170);
nand U365 (N_365,In_324,In_62);
and U366 (N_366,In_143,In_349);
or U367 (N_367,In_54,In_150);
nor U368 (N_368,In_58,In_127);
and U369 (N_369,In_452,In_116);
nand U370 (N_370,In_219,In_87);
nor U371 (N_371,In_3,In_11);
and U372 (N_372,In_127,In_418);
and U373 (N_373,In_486,In_97);
and U374 (N_374,In_255,In_188);
and U375 (N_375,In_345,In_288);
and U376 (N_376,In_93,In_142);
nor U377 (N_377,In_400,In_480);
or U378 (N_378,In_403,In_350);
nand U379 (N_379,In_86,In_333);
and U380 (N_380,In_120,In_13);
nand U381 (N_381,In_456,In_183);
nand U382 (N_382,In_218,In_299);
and U383 (N_383,In_97,In_87);
and U384 (N_384,In_196,In_3);
or U385 (N_385,In_239,In_299);
nor U386 (N_386,In_230,In_384);
and U387 (N_387,In_488,In_174);
nand U388 (N_388,In_35,In_338);
or U389 (N_389,In_162,In_131);
or U390 (N_390,In_117,In_460);
xor U391 (N_391,In_208,In_252);
nand U392 (N_392,In_418,In_101);
nor U393 (N_393,In_246,In_493);
or U394 (N_394,In_163,In_364);
nand U395 (N_395,In_165,In_441);
and U396 (N_396,In_202,In_493);
nor U397 (N_397,In_57,In_155);
or U398 (N_398,In_355,In_454);
nand U399 (N_399,In_63,In_98);
or U400 (N_400,In_97,In_273);
or U401 (N_401,In_268,In_219);
and U402 (N_402,In_109,In_472);
and U403 (N_403,In_292,In_187);
nor U404 (N_404,In_430,In_0);
and U405 (N_405,In_239,In_311);
nand U406 (N_406,In_114,In_216);
nor U407 (N_407,In_82,In_356);
nor U408 (N_408,In_441,In_111);
nand U409 (N_409,In_269,In_205);
or U410 (N_410,In_257,In_495);
nor U411 (N_411,In_116,In_276);
and U412 (N_412,In_496,In_423);
or U413 (N_413,In_391,In_158);
and U414 (N_414,In_455,In_269);
nand U415 (N_415,In_377,In_101);
nand U416 (N_416,In_28,In_97);
xnor U417 (N_417,In_36,In_230);
and U418 (N_418,In_145,In_140);
or U419 (N_419,In_452,In_403);
nand U420 (N_420,In_80,In_89);
and U421 (N_421,In_231,In_404);
nand U422 (N_422,In_470,In_326);
nor U423 (N_423,In_211,In_434);
or U424 (N_424,In_9,In_269);
nand U425 (N_425,In_220,In_147);
or U426 (N_426,In_213,In_466);
and U427 (N_427,In_101,In_330);
and U428 (N_428,In_281,In_407);
nor U429 (N_429,In_454,In_26);
nor U430 (N_430,In_394,In_435);
xnor U431 (N_431,In_360,In_166);
nand U432 (N_432,In_383,In_71);
nor U433 (N_433,In_399,In_282);
xor U434 (N_434,In_66,In_408);
or U435 (N_435,In_69,In_405);
nor U436 (N_436,In_88,In_140);
or U437 (N_437,In_18,In_389);
or U438 (N_438,In_249,In_474);
nand U439 (N_439,In_71,In_312);
or U440 (N_440,In_356,In_412);
and U441 (N_441,In_76,In_53);
and U442 (N_442,In_81,In_361);
nor U443 (N_443,In_209,In_67);
nor U444 (N_444,In_158,In_0);
or U445 (N_445,In_184,In_361);
and U446 (N_446,In_50,In_472);
and U447 (N_447,In_160,In_10);
nand U448 (N_448,In_367,In_24);
or U449 (N_449,In_218,In_345);
and U450 (N_450,In_134,In_65);
or U451 (N_451,In_70,In_176);
xor U452 (N_452,In_168,In_24);
or U453 (N_453,In_188,In_246);
nor U454 (N_454,In_99,In_72);
nand U455 (N_455,In_390,In_315);
nor U456 (N_456,In_315,In_189);
and U457 (N_457,In_60,In_475);
nor U458 (N_458,In_75,In_105);
nor U459 (N_459,In_253,In_130);
and U460 (N_460,In_498,In_371);
xnor U461 (N_461,In_231,In_399);
and U462 (N_462,In_476,In_344);
nand U463 (N_463,In_223,In_461);
xor U464 (N_464,In_379,In_443);
and U465 (N_465,In_124,In_111);
xnor U466 (N_466,In_495,In_362);
and U467 (N_467,In_42,In_18);
and U468 (N_468,In_58,In_395);
nand U469 (N_469,In_391,In_204);
nor U470 (N_470,In_6,In_278);
nor U471 (N_471,In_164,In_213);
xor U472 (N_472,In_208,In_419);
or U473 (N_473,In_136,In_48);
xor U474 (N_474,In_89,In_423);
nand U475 (N_475,In_255,In_268);
and U476 (N_476,In_469,In_158);
nand U477 (N_477,In_226,In_49);
and U478 (N_478,In_19,In_222);
and U479 (N_479,In_33,In_445);
and U480 (N_480,In_468,In_431);
nand U481 (N_481,In_179,In_204);
nor U482 (N_482,In_391,In_1);
or U483 (N_483,In_180,In_268);
nor U484 (N_484,In_461,In_138);
and U485 (N_485,In_122,In_133);
nand U486 (N_486,In_112,In_379);
and U487 (N_487,In_44,In_179);
nand U488 (N_488,In_280,In_4);
or U489 (N_489,In_375,In_360);
nand U490 (N_490,In_312,In_373);
xor U491 (N_491,In_440,In_244);
nor U492 (N_492,In_199,In_338);
nand U493 (N_493,In_313,In_312);
nand U494 (N_494,In_272,In_276);
or U495 (N_495,In_361,In_125);
nor U496 (N_496,In_85,In_194);
xor U497 (N_497,In_481,In_252);
and U498 (N_498,In_122,In_358);
nor U499 (N_499,In_236,In_419);
nor U500 (N_500,N_368,N_404);
nand U501 (N_501,N_48,N_253);
and U502 (N_502,N_2,N_29);
nand U503 (N_503,N_73,N_63);
nor U504 (N_504,N_160,N_250);
xnor U505 (N_505,N_42,N_262);
nor U506 (N_506,N_164,N_139);
or U507 (N_507,N_247,N_421);
or U508 (N_508,N_102,N_449);
or U509 (N_509,N_369,N_292);
nor U510 (N_510,N_85,N_349);
or U511 (N_511,N_269,N_242);
xnor U512 (N_512,N_482,N_177);
or U513 (N_513,N_162,N_335);
nand U514 (N_514,N_394,N_180);
nor U515 (N_515,N_26,N_153);
xnor U516 (N_516,N_83,N_255);
nand U517 (N_517,N_3,N_82);
nor U518 (N_518,N_18,N_283);
nand U519 (N_519,N_190,N_235);
nor U520 (N_520,N_375,N_193);
or U521 (N_521,N_141,N_259);
nand U522 (N_522,N_121,N_330);
nor U523 (N_523,N_216,N_422);
or U524 (N_524,N_445,N_59);
nor U525 (N_525,N_274,N_40);
or U526 (N_526,N_148,N_100);
nor U527 (N_527,N_474,N_336);
xnor U528 (N_528,N_24,N_293);
nor U529 (N_529,N_420,N_205);
or U530 (N_530,N_296,N_110);
or U531 (N_531,N_308,N_472);
or U532 (N_532,N_294,N_75);
and U533 (N_533,N_306,N_265);
or U534 (N_534,N_290,N_62);
nand U535 (N_535,N_328,N_33);
nand U536 (N_536,N_489,N_146);
nand U537 (N_537,N_185,N_476);
nor U538 (N_538,N_457,N_490);
nand U539 (N_539,N_96,N_58);
xor U540 (N_540,N_300,N_116);
nand U541 (N_541,N_480,N_66);
or U542 (N_542,N_383,N_60);
nor U543 (N_543,N_252,N_390);
nor U544 (N_544,N_166,N_355);
and U545 (N_545,N_80,N_178);
nor U546 (N_546,N_311,N_264);
or U547 (N_547,N_373,N_443);
xnor U548 (N_548,N_54,N_98);
nor U549 (N_549,N_270,N_416);
nor U550 (N_550,N_423,N_413);
and U551 (N_551,N_345,N_95);
nand U552 (N_552,N_138,N_402);
nand U553 (N_553,N_9,N_34);
xor U554 (N_554,N_133,N_387);
and U555 (N_555,N_84,N_465);
nand U556 (N_556,N_277,N_268);
or U557 (N_557,N_359,N_441);
and U558 (N_558,N_179,N_393);
or U559 (N_559,N_409,N_101);
nor U560 (N_560,N_266,N_124);
or U561 (N_561,N_494,N_329);
nor U562 (N_562,N_462,N_254);
nand U563 (N_563,N_52,N_151);
and U564 (N_564,N_475,N_49);
nand U565 (N_565,N_27,N_200);
nand U566 (N_566,N_8,N_378);
nor U567 (N_567,N_466,N_384);
nor U568 (N_568,N_318,N_140);
nor U569 (N_569,N_487,N_45);
or U570 (N_570,N_174,N_468);
xnor U571 (N_571,N_463,N_32);
nor U572 (N_572,N_256,N_439);
and U573 (N_573,N_309,N_154);
and U574 (N_574,N_458,N_240);
nor U575 (N_575,N_107,N_415);
and U576 (N_576,N_198,N_497);
xor U577 (N_577,N_284,N_407);
nor U578 (N_578,N_212,N_68);
and U579 (N_579,N_78,N_218);
nor U580 (N_580,N_71,N_232);
and U581 (N_581,N_324,N_15);
or U582 (N_582,N_271,N_94);
and U583 (N_583,N_131,N_209);
and U584 (N_584,N_55,N_234);
nand U585 (N_585,N_65,N_231);
nor U586 (N_586,N_279,N_453);
nand U587 (N_587,N_374,N_76);
and U588 (N_588,N_183,N_481);
nor U589 (N_589,N_321,N_50);
or U590 (N_590,N_347,N_187);
and U591 (N_591,N_286,N_419);
or U592 (N_592,N_167,N_282);
and U593 (N_593,N_471,N_245);
or U594 (N_594,N_291,N_228);
and U595 (N_595,N_137,N_244);
nor U596 (N_596,N_496,N_135);
and U597 (N_597,N_348,N_477);
and U598 (N_598,N_114,N_109);
xnor U599 (N_599,N_464,N_194);
nor U600 (N_600,N_74,N_399);
nor U601 (N_601,N_273,N_280);
and U602 (N_602,N_342,N_120);
nand U603 (N_603,N_352,N_484);
nand U604 (N_604,N_248,N_376);
nor U605 (N_605,N_365,N_455);
xor U606 (N_606,N_10,N_434);
nand U607 (N_607,N_479,N_128);
or U608 (N_608,N_176,N_323);
nor U609 (N_609,N_186,N_281);
and U610 (N_610,N_346,N_338);
or U611 (N_611,N_424,N_312);
nor U612 (N_612,N_181,N_201);
nor U613 (N_613,N_339,N_4);
nor U614 (N_614,N_470,N_20);
nor U615 (N_615,N_31,N_17);
and U616 (N_616,N_221,N_275);
nand U617 (N_617,N_459,N_112);
nand U618 (N_618,N_360,N_446);
nor U619 (N_619,N_103,N_326);
nand U620 (N_620,N_237,N_316);
nand U621 (N_621,N_21,N_440);
xor U622 (N_622,N_363,N_353);
nand U623 (N_623,N_426,N_57);
or U624 (N_624,N_410,N_217);
or U625 (N_625,N_191,N_56);
nor U626 (N_626,N_351,N_81);
or U627 (N_627,N_315,N_157);
nand U628 (N_628,N_173,N_39);
and U629 (N_629,N_276,N_391);
or U630 (N_630,N_343,N_456);
or U631 (N_631,N_230,N_331);
nand U632 (N_632,N_469,N_77);
or U633 (N_633,N_227,N_272);
or U634 (N_634,N_436,N_366);
or U635 (N_635,N_215,N_431);
nor U636 (N_636,N_88,N_207);
nor U637 (N_637,N_208,N_25);
xor U638 (N_638,N_192,N_493);
and U639 (N_639,N_367,N_89);
and U640 (N_640,N_35,N_298);
or U641 (N_641,N_142,N_222);
nor U642 (N_642,N_396,N_28);
nand U643 (N_643,N_263,N_447);
nor U644 (N_644,N_6,N_305);
nor U645 (N_645,N_92,N_22);
or U646 (N_646,N_46,N_129);
and U647 (N_647,N_392,N_182);
xnor U648 (N_648,N_287,N_302);
or U649 (N_649,N_119,N_203);
nand U650 (N_650,N_307,N_202);
xor U651 (N_651,N_196,N_188);
xor U652 (N_652,N_113,N_397);
or U653 (N_653,N_19,N_372);
or U654 (N_654,N_225,N_389);
nor U655 (N_655,N_249,N_319);
xor U656 (N_656,N_461,N_362);
nor U657 (N_657,N_223,N_132);
xnor U658 (N_658,N_213,N_467);
and U659 (N_659,N_219,N_354);
and U660 (N_660,N_149,N_144);
and U661 (N_661,N_233,N_350);
nor U662 (N_662,N_246,N_418);
nor U663 (N_663,N_488,N_23);
nand U664 (N_664,N_451,N_93);
nor U665 (N_665,N_382,N_432);
xor U666 (N_666,N_485,N_122);
and U667 (N_667,N_134,N_498);
nand U668 (N_668,N_386,N_406);
or U669 (N_669,N_184,N_425);
or U670 (N_670,N_161,N_67);
and U671 (N_671,N_195,N_152);
nor U672 (N_672,N_168,N_197);
or U673 (N_673,N_364,N_322);
xnor U674 (N_674,N_38,N_143);
nor U675 (N_675,N_379,N_91);
nand U676 (N_676,N_70,N_332);
nor U677 (N_677,N_108,N_243);
xnor U678 (N_678,N_229,N_314);
nor U679 (N_679,N_370,N_429);
nor U680 (N_680,N_159,N_1);
and U681 (N_681,N_320,N_437);
and U682 (N_682,N_87,N_171);
nor U683 (N_683,N_486,N_297);
nand U684 (N_684,N_51,N_267);
or U685 (N_685,N_452,N_5);
or U686 (N_686,N_204,N_403);
xnor U687 (N_687,N_442,N_64);
nand U688 (N_688,N_414,N_454);
nand U689 (N_689,N_156,N_199);
or U690 (N_690,N_43,N_30);
nand U691 (N_691,N_13,N_86);
or U692 (N_692,N_163,N_172);
nand U693 (N_693,N_427,N_211);
and U694 (N_694,N_123,N_170);
or U695 (N_695,N_126,N_117);
nor U696 (N_696,N_214,N_127);
nand U697 (N_697,N_16,N_450);
or U698 (N_698,N_395,N_206);
nor U699 (N_699,N_130,N_340);
nor U700 (N_700,N_289,N_155);
nor U701 (N_701,N_491,N_41);
nor U702 (N_702,N_261,N_433);
nand U703 (N_703,N_483,N_356);
or U704 (N_704,N_257,N_299);
xnor U705 (N_705,N_388,N_295);
and U706 (N_706,N_325,N_260);
and U707 (N_707,N_220,N_444);
and U708 (N_708,N_435,N_11);
and U709 (N_709,N_288,N_165);
and U710 (N_710,N_150,N_430);
xnor U711 (N_711,N_428,N_499);
nor U712 (N_712,N_236,N_460);
and U713 (N_713,N_344,N_106);
nand U714 (N_714,N_175,N_47);
nand U715 (N_715,N_478,N_412);
xor U716 (N_716,N_44,N_448);
and U717 (N_717,N_210,N_12);
nor U718 (N_718,N_304,N_337);
and U719 (N_719,N_72,N_145);
nor U720 (N_720,N_7,N_301);
xnor U721 (N_721,N_118,N_37);
and U722 (N_722,N_97,N_53);
nand U723 (N_723,N_405,N_371);
nand U724 (N_724,N_251,N_104);
nor U725 (N_725,N_358,N_327);
nor U726 (N_726,N_158,N_90);
or U727 (N_727,N_241,N_239);
and U728 (N_728,N_317,N_417);
nor U729 (N_729,N_278,N_69);
nor U730 (N_730,N_238,N_380);
nor U731 (N_731,N_333,N_14);
and U732 (N_732,N_495,N_226);
nand U733 (N_733,N_438,N_147);
xor U734 (N_734,N_361,N_0);
or U735 (N_735,N_115,N_125);
nand U736 (N_736,N_341,N_408);
or U737 (N_737,N_111,N_313);
nand U738 (N_738,N_224,N_492);
nand U739 (N_739,N_136,N_285);
nand U740 (N_740,N_36,N_357);
and U741 (N_741,N_99,N_401);
nand U742 (N_742,N_377,N_303);
or U743 (N_743,N_411,N_381);
xnor U744 (N_744,N_400,N_258);
and U745 (N_745,N_79,N_169);
nand U746 (N_746,N_398,N_385);
and U747 (N_747,N_310,N_334);
or U748 (N_748,N_105,N_473);
nand U749 (N_749,N_189,N_61);
or U750 (N_750,N_130,N_359);
or U751 (N_751,N_3,N_148);
or U752 (N_752,N_444,N_441);
nor U753 (N_753,N_316,N_151);
nor U754 (N_754,N_327,N_332);
or U755 (N_755,N_76,N_349);
nand U756 (N_756,N_355,N_55);
or U757 (N_757,N_124,N_132);
and U758 (N_758,N_391,N_408);
nand U759 (N_759,N_138,N_75);
nand U760 (N_760,N_237,N_277);
nand U761 (N_761,N_239,N_197);
and U762 (N_762,N_361,N_153);
and U763 (N_763,N_196,N_278);
nor U764 (N_764,N_339,N_207);
and U765 (N_765,N_39,N_451);
nor U766 (N_766,N_216,N_200);
and U767 (N_767,N_163,N_206);
xor U768 (N_768,N_469,N_12);
nand U769 (N_769,N_429,N_297);
and U770 (N_770,N_182,N_341);
and U771 (N_771,N_323,N_331);
nand U772 (N_772,N_282,N_46);
nor U773 (N_773,N_236,N_117);
and U774 (N_774,N_371,N_340);
nor U775 (N_775,N_279,N_31);
and U776 (N_776,N_67,N_328);
or U777 (N_777,N_111,N_418);
and U778 (N_778,N_355,N_84);
or U779 (N_779,N_249,N_321);
nand U780 (N_780,N_104,N_314);
or U781 (N_781,N_496,N_459);
nand U782 (N_782,N_235,N_418);
or U783 (N_783,N_428,N_41);
nand U784 (N_784,N_379,N_9);
and U785 (N_785,N_19,N_288);
xnor U786 (N_786,N_457,N_431);
or U787 (N_787,N_258,N_386);
nand U788 (N_788,N_181,N_371);
nor U789 (N_789,N_285,N_375);
nor U790 (N_790,N_328,N_267);
and U791 (N_791,N_253,N_265);
nor U792 (N_792,N_133,N_314);
or U793 (N_793,N_143,N_127);
nor U794 (N_794,N_351,N_124);
nor U795 (N_795,N_273,N_433);
nor U796 (N_796,N_179,N_352);
and U797 (N_797,N_313,N_486);
or U798 (N_798,N_428,N_110);
nor U799 (N_799,N_237,N_21);
xor U800 (N_800,N_221,N_317);
nand U801 (N_801,N_123,N_410);
or U802 (N_802,N_42,N_448);
and U803 (N_803,N_217,N_467);
nand U804 (N_804,N_289,N_10);
or U805 (N_805,N_214,N_16);
nor U806 (N_806,N_443,N_130);
nor U807 (N_807,N_452,N_245);
xor U808 (N_808,N_275,N_237);
nor U809 (N_809,N_337,N_302);
or U810 (N_810,N_386,N_468);
nor U811 (N_811,N_295,N_474);
nor U812 (N_812,N_144,N_314);
and U813 (N_813,N_395,N_292);
nand U814 (N_814,N_166,N_34);
nor U815 (N_815,N_265,N_249);
xor U816 (N_816,N_356,N_147);
nand U817 (N_817,N_190,N_494);
nor U818 (N_818,N_272,N_68);
nand U819 (N_819,N_310,N_370);
or U820 (N_820,N_226,N_437);
nor U821 (N_821,N_20,N_375);
nand U822 (N_822,N_109,N_163);
nor U823 (N_823,N_198,N_116);
and U824 (N_824,N_174,N_495);
and U825 (N_825,N_2,N_131);
nor U826 (N_826,N_303,N_235);
and U827 (N_827,N_219,N_4);
nor U828 (N_828,N_494,N_63);
nand U829 (N_829,N_388,N_211);
xnor U830 (N_830,N_149,N_162);
or U831 (N_831,N_154,N_0);
and U832 (N_832,N_267,N_115);
nand U833 (N_833,N_228,N_69);
or U834 (N_834,N_143,N_112);
nand U835 (N_835,N_256,N_404);
nor U836 (N_836,N_83,N_465);
nand U837 (N_837,N_135,N_181);
or U838 (N_838,N_193,N_392);
nor U839 (N_839,N_338,N_196);
nor U840 (N_840,N_162,N_494);
and U841 (N_841,N_485,N_465);
nand U842 (N_842,N_168,N_485);
nand U843 (N_843,N_117,N_43);
nand U844 (N_844,N_398,N_330);
or U845 (N_845,N_360,N_238);
or U846 (N_846,N_285,N_219);
and U847 (N_847,N_432,N_251);
or U848 (N_848,N_478,N_383);
or U849 (N_849,N_172,N_227);
nand U850 (N_850,N_25,N_399);
and U851 (N_851,N_130,N_205);
nor U852 (N_852,N_26,N_265);
nand U853 (N_853,N_103,N_351);
nor U854 (N_854,N_359,N_321);
and U855 (N_855,N_190,N_480);
nand U856 (N_856,N_381,N_28);
nand U857 (N_857,N_322,N_307);
and U858 (N_858,N_470,N_399);
nand U859 (N_859,N_21,N_361);
nand U860 (N_860,N_435,N_91);
or U861 (N_861,N_58,N_154);
and U862 (N_862,N_58,N_122);
nor U863 (N_863,N_138,N_453);
nand U864 (N_864,N_81,N_222);
and U865 (N_865,N_365,N_435);
xor U866 (N_866,N_159,N_465);
and U867 (N_867,N_370,N_317);
nor U868 (N_868,N_290,N_228);
nand U869 (N_869,N_64,N_475);
nand U870 (N_870,N_35,N_222);
nor U871 (N_871,N_220,N_463);
nor U872 (N_872,N_399,N_373);
or U873 (N_873,N_284,N_370);
nand U874 (N_874,N_440,N_375);
or U875 (N_875,N_184,N_233);
nand U876 (N_876,N_311,N_441);
nor U877 (N_877,N_433,N_300);
or U878 (N_878,N_39,N_487);
or U879 (N_879,N_49,N_42);
nand U880 (N_880,N_267,N_334);
nor U881 (N_881,N_435,N_58);
xnor U882 (N_882,N_287,N_190);
nor U883 (N_883,N_89,N_378);
and U884 (N_884,N_134,N_420);
xor U885 (N_885,N_147,N_274);
or U886 (N_886,N_369,N_390);
and U887 (N_887,N_234,N_337);
nor U888 (N_888,N_415,N_61);
or U889 (N_889,N_103,N_315);
and U890 (N_890,N_242,N_488);
and U891 (N_891,N_294,N_124);
nor U892 (N_892,N_369,N_331);
and U893 (N_893,N_33,N_263);
and U894 (N_894,N_482,N_310);
nor U895 (N_895,N_448,N_344);
nor U896 (N_896,N_382,N_160);
nor U897 (N_897,N_132,N_18);
nand U898 (N_898,N_328,N_93);
or U899 (N_899,N_227,N_368);
or U900 (N_900,N_405,N_275);
nor U901 (N_901,N_357,N_462);
nand U902 (N_902,N_131,N_197);
and U903 (N_903,N_243,N_74);
and U904 (N_904,N_397,N_312);
or U905 (N_905,N_334,N_364);
or U906 (N_906,N_334,N_330);
or U907 (N_907,N_294,N_240);
and U908 (N_908,N_151,N_57);
nand U909 (N_909,N_415,N_240);
nand U910 (N_910,N_208,N_498);
or U911 (N_911,N_405,N_13);
nor U912 (N_912,N_13,N_353);
or U913 (N_913,N_128,N_231);
or U914 (N_914,N_305,N_347);
xnor U915 (N_915,N_218,N_190);
and U916 (N_916,N_52,N_459);
xnor U917 (N_917,N_332,N_121);
nand U918 (N_918,N_156,N_39);
nand U919 (N_919,N_208,N_210);
nor U920 (N_920,N_444,N_334);
nor U921 (N_921,N_164,N_431);
nand U922 (N_922,N_176,N_230);
or U923 (N_923,N_64,N_306);
nor U924 (N_924,N_70,N_362);
or U925 (N_925,N_98,N_314);
nor U926 (N_926,N_181,N_489);
and U927 (N_927,N_376,N_366);
or U928 (N_928,N_168,N_377);
nor U929 (N_929,N_302,N_319);
or U930 (N_930,N_6,N_116);
xor U931 (N_931,N_385,N_436);
nor U932 (N_932,N_288,N_357);
and U933 (N_933,N_361,N_145);
xnor U934 (N_934,N_324,N_476);
nand U935 (N_935,N_124,N_276);
or U936 (N_936,N_470,N_122);
nor U937 (N_937,N_460,N_426);
nand U938 (N_938,N_244,N_320);
xnor U939 (N_939,N_272,N_323);
nor U940 (N_940,N_45,N_176);
and U941 (N_941,N_52,N_493);
nor U942 (N_942,N_396,N_498);
or U943 (N_943,N_85,N_469);
or U944 (N_944,N_444,N_94);
xor U945 (N_945,N_194,N_401);
nand U946 (N_946,N_316,N_451);
nor U947 (N_947,N_259,N_315);
nand U948 (N_948,N_242,N_132);
and U949 (N_949,N_493,N_102);
nor U950 (N_950,N_116,N_109);
or U951 (N_951,N_394,N_430);
xnor U952 (N_952,N_306,N_76);
and U953 (N_953,N_384,N_303);
or U954 (N_954,N_280,N_419);
nor U955 (N_955,N_429,N_185);
nand U956 (N_956,N_404,N_353);
xor U957 (N_957,N_15,N_359);
nor U958 (N_958,N_218,N_100);
or U959 (N_959,N_359,N_485);
and U960 (N_960,N_448,N_1);
nor U961 (N_961,N_19,N_69);
or U962 (N_962,N_450,N_246);
or U963 (N_963,N_212,N_241);
and U964 (N_964,N_496,N_266);
or U965 (N_965,N_98,N_482);
nor U966 (N_966,N_122,N_345);
nand U967 (N_967,N_491,N_19);
and U968 (N_968,N_287,N_12);
xor U969 (N_969,N_156,N_151);
nor U970 (N_970,N_290,N_307);
nand U971 (N_971,N_375,N_13);
and U972 (N_972,N_119,N_311);
nor U973 (N_973,N_250,N_193);
nand U974 (N_974,N_314,N_173);
nand U975 (N_975,N_499,N_338);
nor U976 (N_976,N_367,N_421);
and U977 (N_977,N_305,N_499);
or U978 (N_978,N_357,N_353);
or U979 (N_979,N_2,N_230);
nor U980 (N_980,N_165,N_327);
nor U981 (N_981,N_151,N_76);
or U982 (N_982,N_149,N_15);
and U983 (N_983,N_486,N_89);
and U984 (N_984,N_157,N_486);
and U985 (N_985,N_125,N_216);
nand U986 (N_986,N_214,N_344);
and U987 (N_987,N_383,N_395);
nand U988 (N_988,N_270,N_20);
nand U989 (N_989,N_2,N_326);
xor U990 (N_990,N_364,N_135);
or U991 (N_991,N_240,N_459);
nor U992 (N_992,N_167,N_53);
and U993 (N_993,N_202,N_401);
xnor U994 (N_994,N_77,N_398);
nand U995 (N_995,N_267,N_110);
nand U996 (N_996,N_102,N_279);
and U997 (N_997,N_165,N_169);
and U998 (N_998,N_154,N_428);
nor U999 (N_999,N_366,N_67);
or U1000 (N_1000,N_641,N_726);
nand U1001 (N_1001,N_604,N_605);
nand U1002 (N_1002,N_615,N_628);
nand U1003 (N_1003,N_926,N_553);
nand U1004 (N_1004,N_540,N_775);
nor U1005 (N_1005,N_886,N_613);
and U1006 (N_1006,N_913,N_829);
and U1007 (N_1007,N_784,N_690);
or U1008 (N_1008,N_729,N_734);
nand U1009 (N_1009,N_779,N_502);
and U1010 (N_1010,N_906,N_688);
nor U1011 (N_1011,N_698,N_697);
xnor U1012 (N_1012,N_921,N_706);
or U1013 (N_1013,N_918,N_981);
or U1014 (N_1014,N_822,N_953);
and U1015 (N_1015,N_670,N_889);
nand U1016 (N_1016,N_550,N_679);
nand U1017 (N_1017,N_555,N_671);
and U1018 (N_1018,N_972,N_601);
nor U1019 (N_1019,N_600,N_687);
nand U1020 (N_1020,N_838,N_957);
or U1021 (N_1021,N_620,N_885);
xnor U1022 (N_1022,N_507,N_716);
xnor U1023 (N_1023,N_989,N_609);
or U1024 (N_1024,N_539,N_730);
xor U1025 (N_1025,N_586,N_661);
xor U1026 (N_1026,N_614,N_871);
nand U1027 (N_1027,N_846,N_535);
and U1028 (N_1028,N_572,N_956);
xor U1029 (N_1029,N_854,N_669);
nor U1030 (N_1030,N_941,N_587);
nor U1031 (N_1031,N_895,N_533);
nand U1032 (N_1032,N_797,N_635);
or U1033 (N_1033,N_530,N_917);
nand U1034 (N_1034,N_722,N_606);
xnor U1035 (N_1035,N_993,N_839);
and U1036 (N_1036,N_691,N_610);
or U1037 (N_1037,N_929,N_982);
and U1038 (N_1038,N_924,N_789);
nor U1039 (N_1039,N_908,N_720);
or U1040 (N_1040,N_888,N_719);
nand U1041 (N_1041,N_975,N_799);
nor U1042 (N_1042,N_684,N_802);
or U1043 (N_1043,N_674,N_905);
nor U1044 (N_1044,N_893,N_509);
xor U1045 (N_1045,N_616,N_686);
nand U1046 (N_1046,N_780,N_579);
or U1047 (N_1047,N_623,N_599);
and U1048 (N_1048,N_894,N_649);
and U1049 (N_1049,N_814,N_642);
nand U1050 (N_1050,N_753,N_875);
nor U1051 (N_1051,N_629,N_723);
or U1052 (N_1052,N_618,N_996);
nor U1053 (N_1053,N_899,N_884);
nor U1054 (N_1054,N_531,N_503);
xnor U1055 (N_1055,N_834,N_717);
nand U1056 (N_1056,N_939,N_971);
nor U1057 (N_1057,N_765,N_934);
nand U1058 (N_1058,N_583,N_644);
xor U1059 (N_1059,N_995,N_808);
nor U1060 (N_1060,N_693,N_845);
xnor U1061 (N_1061,N_997,N_974);
nor U1062 (N_1062,N_580,N_980);
and U1063 (N_1063,N_840,N_912);
nand U1064 (N_1064,N_853,N_567);
or U1065 (N_1065,N_842,N_933);
nor U1066 (N_1066,N_872,N_949);
nand U1067 (N_1067,N_713,N_529);
and U1068 (N_1068,N_633,N_725);
and U1069 (N_1069,N_986,N_807);
and U1070 (N_1070,N_677,N_762);
nor U1071 (N_1071,N_947,N_560);
nand U1072 (N_1072,N_831,N_733);
nor U1073 (N_1073,N_936,N_754);
and U1074 (N_1074,N_803,N_904);
and U1075 (N_1075,N_955,N_685);
nor U1076 (N_1076,N_741,N_666);
and U1077 (N_1077,N_903,N_653);
nand U1078 (N_1078,N_788,N_901);
xor U1079 (N_1079,N_536,N_621);
and U1080 (N_1080,N_896,N_864);
and U1081 (N_1081,N_863,N_522);
and U1082 (N_1082,N_658,N_563);
and U1083 (N_1083,N_774,N_805);
xnor U1084 (N_1084,N_513,N_983);
nor U1085 (N_1085,N_678,N_590);
nand U1086 (N_1086,N_792,N_630);
nand U1087 (N_1087,N_962,N_874);
xnor U1088 (N_1088,N_546,N_935);
and U1089 (N_1089,N_701,N_800);
nand U1090 (N_1090,N_856,N_940);
nand U1091 (N_1091,N_988,N_865);
or U1092 (N_1092,N_636,N_923);
nor U1093 (N_1093,N_708,N_712);
or U1094 (N_1094,N_558,N_813);
nor U1095 (N_1095,N_785,N_773);
or U1096 (N_1096,N_862,N_817);
nand U1097 (N_1097,N_634,N_760);
nand U1098 (N_1098,N_809,N_736);
nor U1099 (N_1099,N_768,N_549);
and U1100 (N_1100,N_878,N_882);
nor U1101 (N_1101,N_891,N_920);
nand U1102 (N_1102,N_657,N_541);
nand U1103 (N_1103,N_819,N_591);
or U1104 (N_1104,N_782,N_897);
xnor U1105 (N_1105,N_619,N_909);
or U1106 (N_1106,N_596,N_617);
and U1107 (N_1107,N_692,N_750);
nand U1108 (N_1108,N_727,N_738);
xor U1109 (N_1109,N_945,N_647);
nor U1110 (N_1110,N_648,N_624);
nor U1111 (N_1111,N_577,N_952);
and U1112 (N_1112,N_561,N_919);
and U1113 (N_1113,N_787,N_739);
nor U1114 (N_1114,N_559,N_746);
or U1115 (N_1115,N_512,N_728);
nand U1116 (N_1116,N_810,N_999);
nor U1117 (N_1117,N_565,N_931);
and U1118 (N_1118,N_847,N_764);
nor U1119 (N_1119,N_597,N_639);
and U1120 (N_1120,N_704,N_824);
and U1121 (N_1121,N_883,N_689);
nand U1122 (N_1122,N_626,N_927);
nand U1123 (N_1123,N_611,N_681);
nand U1124 (N_1124,N_818,N_506);
nor U1125 (N_1125,N_710,N_622);
nand U1126 (N_1126,N_576,N_826);
nand U1127 (N_1127,N_735,N_976);
nand U1128 (N_1128,N_702,N_967);
nand U1129 (N_1129,N_767,N_724);
and U1130 (N_1130,N_742,N_528);
xor U1131 (N_1131,N_925,N_510);
or U1132 (N_1132,N_569,N_756);
or U1133 (N_1133,N_964,N_711);
nor U1134 (N_1134,N_763,N_538);
nand U1135 (N_1135,N_578,N_973);
xor U1136 (N_1136,N_830,N_602);
and U1137 (N_1137,N_961,N_870);
or U1138 (N_1138,N_770,N_815);
or U1139 (N_1139,N_631,N_823);
nand U1140 (N_1140,N_595,N_625);
or U1141 (N_1141,N_584,N_715);
and U1142 (N_1142,N_682,N_777);
and U1143 (N_1143,N_769,N_796);
and U1144 (N_1144,N_547,N_844);
xnor U1145 (N_1145,N_643,N_571);
or U1146 (N_1146,N_588,N_793);
xnor U1147 (N_1147,N_757,N_755);
nand U1148 (N_1148,N_992,N_835);
nand U1149 (N_1149,N_593,N_519);
nor U1150 (N_1150,N_852,N_752);
or U1151 (N_1151,N_585,N_958);
nand U1152 (N_1152,N_907,N_672);
or U1153 (N_1153,N_857,N_612);
or U1154 (N_1154,N_843,N_520);
or U1155 (N_1155,N_695,N_676);
nand U1156 (N_1156,N_749,N_632);
nand U1157 (N_1157,N_968,N_650);
and U1158 (N_1158,N_970,N_850);
xor U1159 (N_1159,N_627,N_915);
and U1160 (N_1160,N_979,N_879);
or U1161 (N_1161,N_603,N_552);
xnor U1162 (N_1162,N_922,N_902);
and U1163 (N_1163,N_751,N_806);
nor U1164 (N_1164,N_900,N_598);
nor U1165 (N_1165,N_887,N_990);
nor U1166 (N_1166,N_705,N_556);
nand U1167 (N_1167,N_532,N_573);
nor U1168 (N_1168,N_545,N_654);
and U1169 (N_1169,N_721,N_948);
nor U1170 (N_1170,N_744,N_662);
nand U1171 (N_1171,N_747,N_943);
nand U1172 (N_1172,N_523,N_855);
nand U1173 (N_1173,N_816,N_740);
and U1174 (N_1174,N_525,N_543);
nor U1175 (N_1175,N_527,N_637);
xnor U1176 (N_1176,N_709,N_828);
nand U1177 (N_1177,N_517,N_759);
nand U1178 (N_1178,N_570,N_521);
nand U1179 (N_1179,N_832,N_978);
nor U1180 (N_1180,N_833,N_638);
and U1181 (N_1181,N_858,N_798);
and U1182 (N_1182,N_700,N_987);
or U1183 (N_1183,N_514,N_673);
nor U1184 (N_1184,N_994,N_821);
nand U1185 (N_1185,N_914,N_737);
nand U1186 (N_1186,N_783,N_772);
or U1187 (N_1187,N_849,N_965);
nor U1188 (N_1188,N_869,N_663);
nand U1189 (N_1189,N_801,N_680);
nor U1190 (N_1190,N_969,N_640);
nor U1191 (N_1191,N_811,N_790);
xor U1192 (N_1192,N_694,N_544);
xnor U1193 (N_1193,N_675,N_836);
xor U1194 (N_1194,N_656,N_954);
and U1195 (N_1195,N_942,N_984);
nand U1196 (N_1196,N_505,N_518);
and U1197 (N_1197,N_537,N_582);
and U1198 (N_1198,N_592,N_574);
nand U1199 (N_1199,N_718,N_881);
nor U1200 (N_1200,N_557,N_861);
or U1201 (N_1201,N_551,N_778);
and U1202 (N_1202,N_991,N_745);
or U1203 (N_1203,N_877,N_960);
xor U1204 (N_1204,N_963,N_707);
and U1205 (N_1205,N_786,N_867);
or U1206 (N_1206,N_916,N_841);
or U1207 (N_1207,N_703,N_589);
nand U1208 (N_1208,N_659,N_515);
nand U1209 (N_1209,N_511,N_928);
nor U1210 (N_1210,N_731,N_938);
xnor U1211 (N_1211,N_959,N_664);
xor U1212 (N_1212,N_890,N_998);
nand U1213 (N_1213,N_714,N_564);
xnor U1214 (N_1214,N_554,N_743);
or U1215 (N_1215,N_851,N_761);
nand U1216 (N_1216,N_665,N_795);
and U1217 (N_1217,N_526,N_668);
nor U1218 (N_1218,N_868,N_848);
nand U1219 (N_1219,N_542,N_950);
nor U1220 (N_1220,N_937,N_946);
or U1221 (N_1221,N_966,N_607);
nand U1222 (N_1222,N_944,N_766);
nor U1223 (N_1223,N_859,N_898);
nand U1224 (N_1224,N_524,N_655);
nor U1225 (N_1225,N_500,N_696);
or U1226 (N_1226,N_667,N_504);
nand U1227 (N_1227,N_646,N_860);
or U1228 (N_1228,N_645,N_837);
or U1229 (N_1229,N_892,N_910);
and U1230 (N_1230,N_791,N_977);
or U1231 (N_1231,N_876,N_594);
nand U1232 (N_1232,N_985,N_683);
nor U1233 (N_1233,N_812,N_575);
and U1234 (N_1234,N_758,N_566);
nor U1235 (N_1235,N_825,N_776);
nand U1236 (N_1236,N_794,N_562);
or U1237 (N_1237,N_951,N_501);
or U1238 (N_1238,N_911,N_652);
nor U1239 (N_1239,N_534,N_651);
nor U1240 (N_1240,N_608,N_820);
and U1241 (N_1241,N_581,N_516);
nor U1242 (N_1242,N_771,N_873);
and U1243 (N_1243,N_568,N_732);
nor U1244 (N_1244,N_827,N_748);
nand U1245 (N_1245,N_932,N_660);
and U1246 (N_1246,N_804,N_508);
or U1247 (N_1247,N_699,N_781);
nand U1248 (N_1248,N_866,N_548);
nor U1249 (N_1249,N_880,N_930);
nand U1250 (N_1250,N_759,N_687);
nand U1251 (N_1251,N_899,N_834);
or U1252 (N_1252,N_892,N_786);
nor U1253 (N_1253,N_521,N_869);
nor U1254 (N_1254,N_945,N_614);
nor U1255 (N_1255,N_844,N_716);
or U1256 (N_1256,N_992,N_968);
nand U1257 (N_1257,N_727,N_649);
nor U1258 (N_1258,N_691,N_794);
or U1259 (N_1259,N_902,N_537);
nor U1260 (N_1260,N_842,N_880);
nand U1261 (N_1261,N_823,N_518);
and U1262 (N_1262,N_620,N_696);
xnor U1263 (N_1263,N_556,N_782);
nor U1264 (N_1264,N_702,N_732);
nand U1265 (N_1265,N_720,N_784);
or U1266 (N_1266,N_561,N_606);
and U1267 (N_1267,N_893,N_807);
and U1268 (N_1268,N_987,N_734);
and U1269 (N_1269,N_749,N_910);
nand U1270 (N_1270,N_674,N_937);
nor U1271 (N_1271,N_545,N_788);
nor U1272 (N_1272,N_562,N_813);
xor U1273 (N_1273,N_956,N_629);
or U1274 (N_1274,N_843,N_780);
xnor U1275 (N_1275,N_569,N_790);
or U1276 (N_1276,N_587,N_507);
or U1277 (N_1277,N_713,N_635);
or U1278 (N_1278,N_616,N_651);
and U1279 (N_1279,N_841,N_733);
or U1280 (N_1280,N_584,N_858);
and U1281 (N_1281,N_810,N_761);
or U1282 (N_1282,N_794,N_571);
nand U1283 (N_1283,N_859,N_870);
or U1284 (N_1284,N_683,N_731);
xor U1285 (N_1285,N_537,N_717);
nor U1286 (N_1286,N_803,N_651);
nor U1287 (N_1287,N_504,N_777);
nand U1288 (N_1288,N_542,N_654);
xnor U1289 (N_1289,N_539,N_763);
nor U1290 (N_1290,N_582,N_730);
xor U1291 (N_1291,N_550,N_926);
or U1292 (N_1292,N_895,N_548);
nand U1293 (N_1293,N_786,N_778);
or U1294 (N_1294,N_653,N_631);
and U1295 (N_1295,N_773,N_551);
nand U1296 (N_1296,N_990,N_938);
xnor U1297 (N_1297,N_750,N_892);
and U1298 (N_1298,N_573,N_773);
or U1299 (N_1299,N_830,N_911);
nand U1300 (N_1300,N_889,N_681);
nor U1301 (N_1301,N_524,N_936);
nand U1302 (N_1302,N_805,N_607);
nor U1303 (N_1303,N_953,N_696);
nor U1304 (N_1304,N_578,N_598);
and U1305 (N_1305,N_735,N_979);
nand U1306 (N_1306,N_862,N_565);
and U1307 (N_1307,N_964,N_598);
nand U1308 (N_1308,N_914,N_882);
nand U1309 (N_1309,N_974,N_670);
and U1310 (N_1310,N_563,N_822);
nor U1311 (N_1311,N_797,N_917);
or U1312 (N_1312,N_741,N_906);
or U1313 (N_1313,N_872,N_622);
xor U1314 (N_1314,N_842,N_962);
and U1315 (N_1315,N_676,N_872);
and U1316 (N_1316,N_617,N_523);
nor U1317 (N_1317,N_523,N_841);
and U1318 (N_1318,N_951,N_825);
nor U1319 (N_1319,N_820,N_719);
nand U1320 (N_1320,N_574,N_754);
nor U1321 (N_1321,N_595,N_618);
and U1322 (N_1322,N_783,N_761);
nor U1323 (N_1323,N_791,N_836);
and U1324 (N_1324,N_553,N_567);
or U1325 (N_1325,N_706,N_956);
and U1326 (N_1326,N_967,N_524);
xnor U1327 (N_1327,N_744,N_610);
nand U1328 (N_1328,N_788,N_962);
and U1329 (N_1329,N_559,N_790);
and U1330 (N_1330,N_939,N_808);
nor U1331 (N_1331,N_588,N_532);
xnor U1332 (N_1332,N_710,N_822);
or U1333 (N_1333,N_749,N_729);
nand U1334 (N_1334,N_876,N_941);
and U1335 (N_1335,N_781,N_991);
and U1336 (N_1336,N_694,N_782);
nand U1337 (N_1337,N_567,N_520);
or U1338 (N_1338,N_957,N_619);
and U1339 (N_1339,N_770,N_745);
xnor U1340 (N_1340,N_569,N_641);
and U1341 (N_1341,N_951,N_671);
nor U1342 (N_1342,N_733,N_627);
and U1343 (N_1343,N_786,N_676);
xnor U1344 (N_1344,N_743,N_525);
xnor U1345 (N_1345,N_679,N_601);
xnor U1346 (N_1346,N_654,N_873);
and U1347 (N_1347,N_642,N_831);
nor U1348 (N_1348,N_546,N_802);
nand U1349 (N_1349,N_938,N_758);
or U1350 (N_1350,N_614,N_565);
nand U1351 (N_1351,N_563,N_882);
nand U1352 (N_1352,N_890,N_956);
nand U1353 (N_1353,N_867,N_567);
xnor U1354 (N_1354,N_585,N_667);
or U1355 (N_1355,N_628,N_887);
xor U1356 (N_1356,N_799,N_761);
or U1357 (N_1357,N_591,N_767);
and U1358 (N_1358,N_845,N_596);
or U1359 (N_1359,N_610,N_732);
or U1360 (N_1360,N_586,N_761);
or U1361 (N_1361,N_771,N_518);
and U1362 (N_1362,N_811,N_590);
nand U1363 (N_1363,N_935,N_766);
or U1364 (N_1364,N_646,N_647);
nor U1365 (N_1365,N_719,N_751);
nand U1366 (N_1366,N_922,N_770);
nor U1367 (N_1367,N_540,N_883);
or U1368 (N_1368,N_881,N_581);
nand U1369 (N_1369,N_820,N_972);
or U1370 (N_1370,N_828,N_683);
nor U1371 (N_1371,N_944,N_616);
and U1372 (N_1372,N_642,N_625);
or U1373 (N_1373,N_951,N_674);
nand U1374 (N_1374,N_746,N_621);
nor U1375 (N_1375,N_873,N_890);
or U1376 (N_1376,N_595,N_997);
nand U1377 (N_1377,N_715,N_847);
or U1378 (N_1378,N_925,N_701);
and U1379 (N_1379,N_522,N_564);
nor U1380 (N_1380,N_998,N_582);
nand U1381 (N_1381,N_976,N_943);
and U1382 (N_1382,N_731,N_863);
or U1383 (N_1383,N_523,N_960);
nor U1384 (N_1384,N_648,N_691);
or U1385 (N_1385,N_954,N_789);
and U1386 (N_1386,N_981,N_546);
and U1387 (N_1387,N_596,N_676);
nor U1388 (N_1388,N_998,N_805);
or U1389 (N_1389,N_939,N_823);
xnor U1390 (N_1390,N_808,N_621);
nand U1391 (N_1391,N_890,N_771);
and U1392 (N_1392,N_519,N_791);
nor U1393 (N_1393,N_584,N_850);
and U1394 (N_1394,N_549,N_909);
nor U1395 (N_1395,N_629,N_937);
or U1396 (N_1396,N_826,N_693);
and U1397 (N_1397,N_558,N_664);
xnor U1398 (N_1398,N_548,N_586);
or U1399 (N_1399,N_921,N_593);
or U1400 (N_1400,N_808,N_942);
or U1401 (N_1401,N_699,N_546);
or U1402 (N_1402,N_903,N_698);
or U1403 (N_1403,N_934,N_956);
nand U1404 (N_1404,N_972,N_527);
nand U1405 (N_1405,N_883,N_692);
nor U1406 (N_1406,N_572,N_801);
or U1407 (N_1407,N_557,N_952);
xnor U1408 (N_1408,N_812,N_996);
or U1409 (N_1409,N_763,N_722);
or U1410 (N_1410,N_531,N_642);
and U1411 (N_1411,N_718,N_505);
nand U1412 (N_1412,N_859,N_709);
or U1413 (N_1413,N_973,N_807);
nor U1414 (N_1414,N_858,N_937);
or U1415 (N_1415,N_787,N_670);
and U1416 (N_1416,N_904,N_652);
or U1417 (N_1417,N_960,N_617);
and U1418 (N_1418,N_525,N_946);
xnor U1419 (N_1419,N_844,N_625);
and U1420 (N_1420,N_615,N_715);
nor U1421 (N_1421,N_779,N_918);
or U1422 (N_1422,N_726,N_667);
nor U1423 (N_1423,N_728,N_954);
and U1424 (N_1424,N_687,N_879);
or U1425 (N_1425,N_533,N_664);
nand U1426 (N_1426,N_753,N_869);
and U1427 (N_1427,N_687,N_659);
xor U1428 (N_1428,N_914,N_574);
nor U1429 (N_1429,N_808,N_816);
and U1430 (N_1430,N_698,N_615);
xnor U1431 (N_1431,N_936,N_631);
or U1432 (N_1432,N_512,N_884);
nand U1433 (N_1433,N_704,N_810);
nor U1434 (N_1434,N_929,N_807);
nand U1435 (N_1435,N_742,N_645);
or U1436 (N_1436,N_960,N_810);
and U1437 (N_1437,N_741,N_764);
nor U1438 (N_1438,N_598,N_624);
nand U1439 (N_1439,N_789,N_505);
and U1440 (N_1440,N_596,N_958);
or U1441 (N_1441,N_944,N_613);
nand U1442 (N_1442,N_922,N_567);
nor U1443 (N_1443,N_622,N_816);
or U1444 (N_1444,N_879,N_844);
xor U1445 (N_1445,N_736,N_735);
xor U1446 (N_1446,N_816,N_926);
nand U1447 (N_1447,N_728,N_818);
and U1448 (N_1448,N_632,N_621);
xor U1449 (N_1449,N_634,N_589);
nand U1450 (N_1450,N_673,N_663);
nor U1451 (N_1451,N_969,N_766);
nand U1452 (N_1452,N_774,N_897);
and U1453 (N_1453,N_642,N_584);
nand U1454 (N_1454,N_705,N_684);
nor U1455 (N_1455,N_994,N_757);
nor U1456 (N_1456,N_876,N_669);
and U1457 (N_1457,N_524,N_572);
or U1458 (N_1458,N_955,N_627);
or U1459 (N_1459,N_973,N_734);
nand U1460 (N_1460,N_813,N_939);
or U1461 (N_1461,N_614,N_543);
nor U1462 (N_1462,N_611,N_688);
and U1463 (N_1463,N_945,N_894);
nand U1464 (N_1464,N_795,N_544);
or U1465 (N_1465,N_735,N_555);
and U1466 (N_1466,N_811,N_671);
or U1467 (N_1467,N_618,N_809);
nand U1468 (N_1468,N_910,N_701);
nand U1469 (N_1469,N_523,N_800);
nand U1470 (N_1470,N_696,N_579);
xor U1471 (N_1471,N_523,N_731);
or U1472 (N_1472,N_629,N_979);
or U1473 (N_1473,N_628,N_906);
nand U1474 (N_1474,N_874,N_782);
nor U1475 (N_1475,N_885,N_715);
nor U1476 (N_1476,N_506,N_919);
and U1477 (N_1477,N_656,N_673);
nand U1478 (N_1478,N_812,N_813);
nor U1479 (N_1479,N_572,N_653);
nand U1480 (N_1480,N_584,N_680);
and U1481 (N_1481,N_777,N_695);
nand U1482 (N_1482,N_796,N_562);
and U1483 (N_1483,N_596,N_792);
nor U1484 (N_1484,N_750,N_501);
or U1485 (N_1485,N_600,N_516);
and U1486 (N_1486,N_783,N_827);
and U1487 (N_1487,N_882,N_804);
and U1488 (N_1488,N_959,N_556);
nor U1489 (N_1489,N_853,N_825);
xor U1490 (N_1490,N_923,N_746);
and U1491 (N_1491,N_809,N_794);
or U1492 (N_1492,N_861,N_529);
nor U1493 (N_1493,N_853,N_935);
xor U1494 (N_1494,N_775,N_985);
and U1495 (N_1495,N_951,N_978);
nor U1496 (N_1496,N_513,N_923);
and U1497 (N_1497,N_708,N_553);
and U1498 (N_1498,N_862,N_780);
nor U1499 (N_1499,N_942,N_631);
or U1500 (N_1500,N_1218,N_1080);
nor U1501 (N_1501,N_1306,N_1471);
and U1502 (N_1502,N_1204,N_1011);
and U1503 (N_1503,N_1372,N_1376);
nor U1504 (N_1504,N_1115,N_1320);
nor U1505 (N_1505,N_1422,N_1323);
or U1506 (N_1506,N_1481,N_1234);
and U1507 (N_1507,N_1223,N_1339);
and U1508 (N_1508,N_1280,N_1059);
nor U1509 (N_1509,N_1499,N_1336);
and U1510 (N_1510,N_1463,N_1007);
nor U1511 (N_1511,N_1495,N_1328);
nor U1512 (N_1512,N_1180,N_1464);
nor U1513 (N_1513,N_1267,N_1033);
or U1514 (N_1514,N_1497,N_1069);
or U1515 (N_1515,N_1181,N_1206);
nor U1516 (N_1516,N_1379,N_1082);
nand U1517 (N_1517,N_1288,N_1003);
xor U1518 (N_1518,N_1066,N_1341);
nor U1519 (N_1519,N_1386,N_1091);
and U1520 (N_1520,N_1403,N_1151);
or U1521 (N_1521,N_1261,N_1197);
xor U1522 (N_1522,N_1165,N_1441);
nor U1523 (N_1523,N_1237,N_1296);
and U1524 (N_1524,N_1483,N_1345);
or U1525 (N_1525,N_1251,N_1325);
and U1526 (N_1526,N_1006,N_1119);
nand U1527 (N_1527,N_1108,N_1294);
nor U1528 (N_1528,N_1032,N_1461);
nor U1529 (N_1529,N_1149,N_1125);
nand U1530 (N_1530,N_1021,N_1298);
nor U1531 (N_1531,N_1063,N_1430);
nor U1532 (N_1532,N_1466,N_1076);
and U1533 (N_1533,N_1214,N_1365);
nand U1534 (N_1534,N_1484,N_1240);
or U1535 (N_1535,N_1433,N_1233);
nand U1536 (N_1536,N_1492,N_1144);
xor U1537 (N_1537,N_1040,N_1213);
and U1538 (N_1538,N_1434,N_1459);
or U1539 (N_1539,N_1259,N_1161);
nand U1540 (N_1540,N_1418,N_1286);
xnor U1541 (N_1541,N_1049,N_1061);
nor U1542 (N_1542,N_1030,N_1447);
and U1543 (N_1543,N_1085,N_1107);
nand U1544 (N_1544,N_1392,N_1385);
xor U1545 (N_1545,N_1332,N_1494);
or U1546 (N_1546,N_1147,N_1239);
nand U1547 (N_1547,N_1046,N_1384);
nor U1548 (N_1548,N_1127,N_1402);
nor U1549 (N_1549,N_1230,N_1360);
or U1550 (N_1550,N_1162,N_1020);
or U1551 (N_1551,N_1216,N_1278);
and U1552 (N_1552,N_1176,N_1319);
nand U1553 (N_1553,N_1419,N_1112);
nor U1554 (N_1554,N_1035,N_1406);
nor U1555 (N_1555,N_1122,N_1302);
nand U1556 (N_1556,N_1014,N_1383);
or U1557 (N_1557,N_1052,N_1293);
nand U1558 (N_1558,N_1462,N_1196);
nand U1559 (N_1559,N_1452,N_1093);
or U1560 (N_1560,N_1106,N_1388);
and U1561 (N_1561,N_1169,N_1245);
or U1562 (N_1562,N_1166,N_1203);
nor U1563 (N_1563,N_1292,N_1362);
xor U1564 (N_1564,N_1351,N_1221);
and U1565 (N_1565,N_1142,N_1427);
and U1566 (N_1566,N_1205,N_1283);
and U1567 (N_1567,N_1238,N_1289);
or U1568 (N_1568,N_1359,N_1015);
nor U1569 (N_1569,N_1055,N_1044);
or U1570 (N_1570,N_1005,N_1295);
and U1571 (N_1571,N_1363,N_1358);
nor U1572 (N_1572,N_1153,N_1279);
and U1573 (N_1573,N_1490,N_1172);
nor U1574 (N_1574,N_1331,N_1075);
and U1575 (N_1575,N_1311,N_1160);
and U1576 (N_1576,N_1042,N_1235);
and U1577 (N_1577,N_1355,N_1211);
nor U1578 (N_1578,N_1310,N_1013);
nor U1579 (N_1579,N_1375,N_1329);
nor U1580 (N_1580,N_1201,N_1408);
nor U1581 (N_1581,N_1192,N_1225);
and U1582 (N_1582,N_1034,N_1140);
or U1583 (N_1583,N_1473,N_1154);
or U1584 (N_1584,N_1099,N_1232);
nor U1585 (N_1585,N_1002,N_1070);
nor U1586 (N_1586,N_1190,N_1171);
or U1587 (N_1587,N_1404,N_1307);
and U1588 (N_1588,N_1269,N_1493);
nor U1589 (N_1589,N_1326,N_1148);
xnor U1590 (N_1590,N_1198,N_1486);
nand U1591 (N_1591,N_1256,N_1215);
nand U1592 (N_1592,N_1395,N_1361);
nor U1593 (N_1593,N_1152,N_1079);
nand U1594 (N_1594,N_1023,N_1182);
and U1595 (N_1595,N_1167,N_1134);
or U1596 (N_1596,N_1027,N_1231);
and U1597 (N_1597,N_1110,N_1432);
nor U1598 (N_1598,N_1420,N_1087);
or U1599 (N_1599,N_1116,N_1094);
xnor U1600 (N_1600,N_1100,N_1103);
nor U1601 (N_1601,N_1048,N_1413);
nand U1602 (N_1602,N_1487,N_1390);
or U1603 (N_1603,N_1194,N_1448);
nand U1604 (N_1604,N_1443,N_1368);
nor U1605 (N_1605,N_1193,N_1444);
or U1606 (N_1606,N_1429,N_1356);
xnor U1607 (N_1607,N_1414,N_1405);
or U1608 (N_1608,N_1271,N_1482);
nor U1609 (N_1609,N_1120,N_1022);
or U1610 (N_1610,N_1253,N_1019);
nand U1611 (N_1611,N_1353,N_1062);
or U1612 (N_1612,N_1017,N_1210);
or U1613 (N_1613,N_1469,N_1423);
or U1614 (N_1614,N_1141,N_1474);
or U1615 (N_1615,N_1209,N_1489);
and U1616 (N_1616,N_1174,N_1284);
nor U1617 (N_1617,N_1199,N_1138);
and U1618 (N_1618,N_1123,N_1491);
nor U1619 (N_1619,N_1391,N_1380);
nor U1620 (N_1620,N_1426,N_1188);
or U1621 (N_1621,N_1092,N_1064);
xor U1622 (N_1622,N_1342,N_1073);
and U1623 (N_1623,N_1349,N_1184);
or U1624 (N_1624,N_1200,N_1291);
or U1625 (N_1625,N_1246,N_1428);
or U1626 (N_1626,N_1410,N_1453);
and U1627 (N_1627,N_1400,N_1129);
or U1628 (N_1628,N_1337,N_1409);
or U1629 (N_1629,N_1065,N_1377);
nor U1630 (N_1630,N_1281,N_1313);
and U1631 (N_1631,N_1244,N_1333);
or U1632 (N_1632,N_1071,N_1010);
nor U1633 (N_1633,N_1118,N_1089);
or U1634 (N_1634,N_1425,N_1304);
or U1635 (N_1635,N_1440,N_1460);
xnor U1636 (N_1636,N_1131,N_1163);
nand U1637 (N_1637,N_1137,N_1257);
and U1638 (N_1638,N_1258,N_1101);
and U1639 (N_1639,N_1476,N_1366);
nand U1640 (N_1640,N_1401,N_1277);
or U1641 (N_1641,N_1290,N_1096);
nor U1642 (N_1642,N_1369,N_1037);
nand U1643 (N_1643,N_1185,N_1393);
nor U1644 (N_1644,N_1450,N_1378);
nor U1645 (N_1645,N_1111,N_1114);
nand U1646 (N_1646,N_1327,N_1242);
or U1647 (N_1647,N_1109,N_1449);
or U1648 (N_1648,N_1478,N_1241);
nor U1649 (N_1649,N_1217,N_1164);
and U1650 (N_1650,N_1097,N_1054);
or U1651 (N_1651,N_1268,N_1431);
or U1652 (N_1652,N_1399,N_1407);
xor U1653 (N_1653,N_1025,N_1475);
nand U1654 (N_1654,N_1272,N_1456);
nor U1655 (N_1655,N_1439,N_1236);
and U1656 (N_1656,N_1155,N_1031);
xor U1657 (N_1657,N_1248,N_1126);
xnor U1658 (N_1658,N_1057,N_1050);
nand U1659 (N_1659,N_1227,N_1117);
or U1660 (N_1660,N_1041,N_1446);
nor U1661 (N_1661,N_1266,N_1145);
and U1662 (N_1662,N_1043,N_1202);
xor U1663 (N_1663,N_1330,N_1036);
nor U1664 (N_1664,N_1299,N_1053);
nand U1665 (N_1665,N_1477,N_1146);
or U1666 (N_1666,N_1128,N_1029);
or U1667 (N_1667,N_1287,N_1394);
nor U1668 (N_1668,N_1273,N_1472);
nor U1669 (N_1669,N_1098,N_1170);
nor U1670 (N_1670,N_1016,N_1157);
and U1671 (N_1671,N_1354,N_1156);
or U1672 (N_1672,N_1135,N_1343);
and U1673 (N_1673,N_1018,N_1308);
xor U1674 (N_1674,N_1189,N_1322);
nand U1675 (N_1675,N_1421,N_1265);
xor U1676 (N_1676,N_1183,N_1367);
nand U1677 (N_1677,N_1305,N_1415);
and U1678 (N_1678,N_1324,N_1077);
and U1679 (N_1679,N_1350,N_1270);
or U1680 (N_1680,N_1334,N_1488);
or U1681 (N_1681,N_1121,N_1297);
nand U1682 (N_1682,N_1274,N_1250);
or U1683 (N_1683,N_1132,N_1454);
and U1684 (N_1684,N_1067,N_1178);
nor U1685 (N_1685,N_1045,N_1276);
xnor U1686 (N_1686,N_1348,N_1424);
and U1687 (N_1687,N_1445,N_1102);
and U1688 (N_1688,N_1028,N_1451);
nand U1689 (N_1689,N_1060,N_1412);
and U1690 (N_1690,N_1309,N_1442);
nand U1691 (N_1691,N_1090,N_1047);
and U1692 (N_1692,N_1374,N_1321);
nor U1693 (N_1693,N_1397,N_1387);
or U1694 (N_1694,N_1143,N_1396);
or U1695 (N_1695,N_1026,N_1187);
or U1696 (N_1696,N_1254,N_1315);
and U1697 (N_1697,N_1136,N_1262);
xor U1698 (N_1698,N_1470,N_1072);
or U1699 (N_1699,N_1078,N_1219);
nand U1700 (N_1700,N_1357,N_1058);
or U1701 (N_1701,N_1458,N_1024);
or U1702 (N_1702,N_1243,N_1373);
nor U1703 (N_1703,N_1247,N_1104);
and U1704 (N_1704,N_1195,N_1220);
xnor U1705 (N_1705,N_1485,N_1004);
nor U1706 (N_1706,N_1222,N_1496);
and U1707 (N_1707,N_1318,N_1371);
and U1708 (N_1708,N_1340,N_1175);
or U1709 (N_1709,N_1457,N_1438);
and U1710 (N_1710,N_1000,N_1285);
nand U1711 (N_1711,N_1364,N_1467);
nand U1712 (N_1712,N_1084,N_1335);
or U1713 (N_1713,N_1051,N_1263);
and U1714 (N_1714,N_1411,N_1186);
xor U1715 (N_1715,N_1074,N_1249);
nor U1716 (N_1716,N_1382,N_1207);
nand U1717 (N_1717,N_1224,N_1133);
nor U1718 (N_1718,N_1039,N_1455);
nand U1719 (N_1719,N_1346,N_1177);
or U1720 (N_1720,N_1083,N_1300);
nand U1721 (N_1721,N_1381,N_1095);
nor U1722 (N_1722,N_1344,N_1226);
xor U1723 (N_1723,N_1158,N_1317);
or U1724 (N_1724,N_1316,N_1150);
nand U1725 (N_1725,N_1168,N_1437);
or U1726 (N_1726,N_1229,N_1130);
and U1727 (N_1727,N_1212,N_1314);
nand U1728 (N_1728,N_1338,N_1370);
or U1729 (N_1729,N_1105,N_1008);
or U1730 (N_1730,N_1252,N_1191);
or U1731 (N_1731,N_1312,N_1282);
xnor U1732 (N_1732,N_1113,N_1301);
nor U1733 (N_1733,N_1173,N_1435);
nand U1734 (N_1734,N_1139,N_1416);
nand U1735 (N_1735,N_1086,N_1465);
nor U1736 (N_1736,N_1124,N_1398);
and U1737 (N_1737,N_1159,N_1179);
xnor U1738 (N_1738,N_1009,N_1056);
or U1739 (N_1739,N_1001,N_1275);
or U1740 (N_1740,N_1264,N_1068);
and U1741 (N_1741,N_1468,N_1347);
xor U1742 (N_1742,N_1352,N_1255);
and U1743 (N_1743,N_1417,N_1303);
nand U1744 (N_1744,N_1208,N_1480);
nor U1745 (N_1745,N_1012,N_1081);
or U1746 (N_1746,N_1038,N_1479);
nand U1747 (N_1747,N_1228,N_1260);
nand U1748 (N_1748,N_1436,N_1389);
and U1749 (N_1749,N_1088,N_1498);
nor U1750 (N_1750,N_1094,N_1395);
nor U1751 (N_1751,N_1211,N_1310);
or U1752 (N_1752,N_1066,N_1005);
or U1753 (N_1753,N_1333,N_1087);
and U1754 (N_1754,N_1233,N_1148);
or U1755 (N_1755,N_1180,N_1468);
xnor U1756 (N_1756,N_1292,N_1331);
or U1757 (N_1757,N_1235,N_1018);
or U1758 (N_1758,N_1256,N_1106);
nor U1759 (N_1759,N_1303,N_1284);
nor U1760 (N_1760,N_1487,N_1476);
nand U1761 (N_1761,N_1280,N_1090);
nor U1762 (N_1762,N_1294,N_1216);
or U1763 (N_1763,N_1244,N_1094);
nand U1764 (N_1764,N_1375,N_1445);
nor U1765 (N_1765,N_1200,N_1396);
nand U1766 (N_1766,N_1489,N_1118);
xor U1767 (N_1767,N_1001,N_1402);
nor U1768 (N_1768,N_1092,N_1044);
nor U1769 (N_1769,N_1121,N_1102);
nand U1770 (N_1770,N_1261,N_1451);
or U1771 (N_1771,N_1294,N_1496);
xor U1772 (N_1772,N_1110,N_1207);
or U1773 (N_1773,N_1122,N_1466);
nor U1774 (N_1774,N_1148,N_1036);
and U1775 (N_1775,N_1164,N_1345);
and U1776 (N_1776,N_1268,N_1029);
and U1777 (N_1777,N_1076,N_1090);
nor U1778 (N_1778,N_1398,N_1014);
nor U1779 (N_1779,N_1270,N_1384);
nor U1780 (N_1780,N_1128,N_1406);
or U1781 (N_1781,N_1481,N_1360);
nand U1782 (N_1782,N_1022,N_1385);
nor U1783 (N_1783,N_1146,N_1287);
and U1784 (N_1784,N_1452,N_1345);
or U1785 (N_1785,N_1066,N_1244);
nor U1786 (N_1786,N_1454,N_1303);
nor U1787 (N_1787,N_1436,N_1365);
or U1788 (N_1788,N_1010,N_1073);
nor U1789 (N_1789,N_1167,N_1343);
and U1790 (N_1790,N_1280,N_1369);
and U1791 (N_1791,N_1247,N_1387);
nor U1792 (N_1792,N_1067,N_1200);
nand U1793 (N_1793,N_1210,N_1396);
or U1794 (N_1794,N_1421,N_1102);
nor U1795 (N_1795,N_1263,N_1274);
nor U1796 (N_1796,N_1156,N_1359);
and U1797 (N_1797,N_1185,N_1178);
nor U1798 (N_1798,N_1043,N_1462);
xnor U1799 (N_1799,N_1261,N_1230);
nand U1800 (N_1800,N_1394,N_1146);
nor U1801 (N_1801,N_1243,N_1435);
and U1802 (N_1802,N_1082,N_1356);
xor U1803 (N_1803,N_1103,N_1211);
and U1804 (N_1804,N_1465,N_1220);
and U1805 (N_1805,N_1337,N_1126);
nand U1806 (N_1806,N_1318,N_1078);
xor U1807 (N_1807,N_1061,N_1412);
and U1808 (N_1808,N_1222,N_1268);
nand U1809 (N_1809,N_1229,N_1399);
or U1810 (N_1810,N_1163,N_1107);
nand U1811 (N_1811,N_1001,N_1073);
or U1812 (N_1812,N_1416,N_1320);
nor U1813 (N_1813,N_1431,N_1222);
nand U1814 (N_1814,N_1247,N_1089);
nor U1815 (N_1815,N_1386,N_1171);
or U1816 (N_1816,N_1257,N_1291);
xnor U1817 (N_1817,N_1340,N_1384);
nor U1818 (N_1818,N_1178,N_1143);
nor U1819 (N_1819,N_1475,N_1447);
nor U1820 (N_1820,N_1345,N_1349);
and U1821 (N_1821,N_1366,N_1269);
and U1822 (N_1822,N_1399,N_1302);
nand U1823 (N_1823,N_1377,N_1071);
or U1824 (N_1824,N_1418,N_1211);
nand U1825 (N_1825,N_1296,N_1407);
nand U1826 (N_1826,N_1133,N_1272);
nor U1827 (N_1827,N_1259,N_1418);
nand U1828 (N_1828,N_1315,N_1173);
nor U1829 (N_1829,N_1036,N_1477);
or U1830 (N_1830,N_1164,N_1303);
or U1831 (N_1831,N_1080,N_1014);
or U1832 (N_1832,N_1293,N_1133);
nor U1833 (N_1833,N_1249,N_1362);
and U1834 (N_1834,N_1210,N_1049);
or U1835 (N_1835,N_1289,N_1189);
xor U1836 (N_1836,N_1123,N_1293);
nand U1837 (N_1837,N_1064,N_1072);
and U1838 (N_1838,N_1285,N_1498);
nand U1839 (N_1839,N_1332,N_1124);
nor U1840 (N_1840,N_1292,N_1282);
nand U1841 (N_1841,N_1187,N_1073);
and U1842 (N_1842,N_1399,N_1363);
and U1843 (N_1843,N_1193,N_1473);
and U1844 (N_1844,N_1004,N_1357);
and U1845 (N_1845,N_1357,N_1167);
nand U1846 (N_1846,N_1099,N_1438);
or U1847 (N_1847,N_1100,N_1212);
xor U1848 (N_1848,N_1306,N_1379);
or U1849 (N_1849,N_1262,N_1411);
nor U1850 (N_1850,N_1211,N_1155);
or U1851 (N_1851,N_1251,N_1337);
nor U1852 (N_1852,N_1036,N_1316);
nor U1853 (N_1853,N_1279,N_1223);
or U1854 (N_1854,N_1132,N_1487);
nand U1855 (N_1855,N_1067,N_1155);
nor U1856 (N_1856,N_1094,N_1025);
or U1857 (N_1857,N_1486,N_1138);
nor U1858 (N_1858,N_1092,N_1131);
xor U1859 (N_1859,N_1144,N_1219);
and U1860 (N_1860,N_1248,N_1183);
nand U1861 (N_1861,N_1336,N_1050);
nor U1862 (N_1862,N_1456,N_1258);
nand U1863 (N_1863,N_1120,N_1426);
or U1864 (N_1864,N_1104,N_1337);
or U1865 (N_1865,N_1009,N_1385);
nand U1866 (N_1866,N_1286,N_1001);
and U1867 (N_1867,N_1019,N_1134);
xor U1868 (N_1868,N_1327,N_1197);
nor U1869 (N_1869,N_1326,N_1383);
nand U1870 (N_1870,N_1323,N_1310);
or U1871 (N_1871,N_1432,N_1035);
and U1872 (N_1872,N_1274,N_1363);
and U1873 (N_1873,N_1066,N_1115);
nand U1874 (N_1874,N_1374,N_1380);
and U1875 (N_1875,N_1385,N_1230);
nor U1876 (N_1876,N_1415,N_1189);
xnor U1877 (N_1877,N_1087,N_1419);
nand U1878 (N_1878,N_1095,N_1216);
or U1879 (N_1879,N_1067,N_1286);
or U1880 (N_1880,N_1330,N_1112);
nor U1881 (N_1881,N_1135,N_1211);
nand U1882 (N_1882,N_1254,N_1068);
nand U1883 (N_1883,N_1257,N_1106);
nor U1884 (N_1884,N_1322,N_1051);
nand U1885 (N_1885,N_1210,N_1386);
nor U1886 (N_1886,N_1029,N_1088);
nor U1887 (N_1887,N_1254,N_1303);
and U1888 (N_1888,N_1448,N_1216);
and U1889 (N_1889,N_1003,N_1231);
nand U1890 (N_1890,N_1418,N_1109);
xnor U1891 (N_1891,N_1398,N_1386);
and U1892 (N_1892,N_1405,N_1011);
nor U1893 (N_1893,N_1293,N_1131);
nor U1894 (N_1894,N_1002,N_1143);
or U1895 (N_1895,N_1432,N_1238);
nor U1896 (N_1896,N_1357,N_1253);
nor U1897 (N_1897,N_1131,N_1248);
or U1898 (N_1898,N_1493,N_1051);
nor U1899 (N_1899,N_1016,N_1495);
and U1900 (N_1900,N_1273,N_1109);
nand U1901 (N_1901,N_1391,N_1198);
or U1902 (N_1902,N_1123,N_1187);
or U1903 (N_1903,N_1191,N_1345);
nand U1904 (N_1904,N_1441,N_1420);
and U1905 (N_1905,N_1008,N_1033);
and U1906 (N_1906,N_1333,N_1028);
nand U1907 (N_1907,N_1240,N_1261);
nand U1908 (N_1908,N_1210,N_1032);
nor U1909 (N_1909,N_1246,N_1466);
nor U1910 (N_1910,N_1183,N_1390);
nand U1911 (N_1911,N_1260,N_1376);
nor U1912 (N_1912,N_1414,N_1343);
and U1913 (N_1913,N_1011,N_1473);
xnor U1914 (N_1914,N_1129,N_1309);
nand U1915 (N_1915,N_1387,N_1245);
or U1916 (N_1916,N_1343,N_1449);
nand U1917 (N_1917,N_1132,N_1288);
nand U1918 (N_1918,N_1400,N_1075);
and U1919 (N_1919,N_1400,N_1475);
and U1920 (N_1920,N_1282,N_1382);
nand U1921 (N_1921,N_1459,N_1169);
and U1922 (N_1922,N_1111,N_1254);
nor U1923 (N_1923,N_1446,N_1002);
nor U1924 (N_1924,N_1055,N_1105);
and U1925 (N_1925,N_1246,N_1448);
or U1926 (N_1926,N_1065,N_1109);
nor U1927 (N_1927,N_1279,N_1426);
or U1928 (N_1928,N_1230,N_1387);
nand U1929 (N_1929,N_1211,N_1308);
or U1930 (N_1930,N_1485,N_1227);
nor U1931 (N_1931,N_1200,N_1244);
xnor U1932 (N_1932,N_1236,N_1352);
nand U1933 (N_1933,N_1467,N_1431);
and U1934 (N_1934,N_1148,N_1186);
or U1935 (N_1935,N_1118,N_1473);
nand U1936 (N_1936,N_1447,N_1040);
nand U1937 (N_1937,N_1144,N_1442);
xnor U1938 (N_1938,N_1228,N_1442);
or U1939 (N_1939,N_1368,N_1091);
or U1940 (N_1940,N_1235,N_1420);
nor U1941 (N_1941,N_1069,N_1373);
nor U1942 (N_1942,N_1464,N_1178);
nor U1943 (N_1943,N_1084,N_1126);
nor U1944 (N_1944,N_1452,N_1175);
or U1945 (N_1945,N_1119,N_1178);
nand U1946 (N_1946,N_1281,N_1309);
nand U1947 (N_1947,N_1444,N_1227);
and U1948 (N_1948,N_1012,N_1261);
nand U1949 (N_1949,N_1396,N_1033);
and U1950 (N_1950,N_1089,N_1085);
or U1951 (N_1951,N_1280,N_1106);
nor U1952 (N_1952,N_1211,N_1488);
and U1953 (N_1953,N_1209,N_1432);
and U1954 (N_1954,N_1496,N_1473);
nand U1955 (N_1955,N_1111,N_1235);
nor U1956 (N_1956,N_1274,N_1474);
or U1957 (N_1957,N_1418,N_1057);
nand U1958 (N_1958,N_1138,N_1380);
nor U1959 (N_1959,N_1039,N_1077);
nor U1960 (N_1960,N_1470,N_1250);
and U1961 (N_1961,N_1186,N_1236);
nor U1962 (N_1962,N_1311,N_1097);
nor U1963 (N_1963,N_1295,N_1432);
and U1964 (N_1964,N_1084,N_1433);
nand U1965 (N_1965,N_1466,N_1380);
nor U1966 (N_1966,N_1183,N_1232);
nand U1967 (N_1967,N_1190,N_1097);
nor U1968 (N_1968,N_1315,N_1348);
and U1969 (N_1969,N_1242,N_1186);
nand U1970 (N_1970,N_1169,N_1147);
nand U1971 (N_1971,N_1413,N_1068);
nand U1972 (N_1972,N_1462,N_1419);
and U1973 (N_1973,N_1446,N_1454);
or U1974 (N_1974,N_1150,N_1187);
nand U1975 (N_1975,N_1483,N_1488);
and U1976 (N_1976,N_1078,N_1089);
nor U1977 (N_1977,N_1396,N_1185);
and U1978 (N_1978,N_1347,N_1227);
or U1979 (N_1979,N_1372,N_1174);
and U1980 (N_1980,N_1412,N_1169);
nand U1981 (N_1981,N_1283,N_1019);
and U1982 (N_1982,N_1177,N_1423);
nand U1983 (N_1983,N_1167,N_1318);
nor U1984 (N_1984,N_1298,N_1103);
and U1985 (N_1985,N_1459,N_1403);
or U1986 (N_1986,N_1011,N_1480);
nand U1987 (N_1987,N_1231,N_1095);
nand U1988 (N_1988,N_1460,N_1380);
or U1989 (N_1989,N_1358,N_1467);
nor U1990 (N_1990,N_1321,N_1459);
nor U1991 (N_1991,N_1323,N_1088);
nor U1992 (N_1992,N_1054,N_1214);
or U1993 (N_1993,N_1006,N_1475);
xor U1994 (N_1994,N_1492,N_1395);
or U1995 (N_1995,N_1404,N_1475);
and U1996 (N_1996,N_1419,N_1147);
nand U1997 (N_1997,N_1290,N_1154);
nor U1998 (N_1998,N_1002,N_1327);
nor U1999 (N_1999,N_1053,N_1185);
and U2000 (N_2000,N_1707,N_1714);
nand U2001 (N_2001,N_1764,N_1863);
nand U2002 (N_2002,N_1900,N_1547);
nand U2003 (N_2003,N_1517,N_1561);
and U2004 (N_2004,N_1568,N_1655);
nand U2005 (N_2005,N_1526,N_1948);
and U2006 (N_2006,N_1838,N_1984);
nand U2007 (N_2007,N_1605,N_1706);
nor U2008 (N_2008,N_1708,N_1562);
nand U2009 (N_2009,N_1993,N_1869);
or U2010 (N_2010,N_1534,N_1814);
nor U2011 (N_2011,N_1783,N_1961);
nor U2012 (N_2012,N_1668,N_1638);
and U2013 (N_2013,N_1724,N_1693);
and U2014 (N_2014,N_1761,N_1701);
and U2015 (N_2015,N_1542,N_1712);
nand U2016 (N_2016,N_1659,N_1632);
nor U2017 (N_2017,N_1620,N_1933);
xnor U2018 (N_2018,N_1621,N_1716);
nor U2019 (N_2019,N_1841,N_1760);
and U2020 (N_2020,N_1540,N_1992);
or U2021 (N_2021,N_1776,N_1998);
nor U2022 (N_2022,N_1868,N_1514);
nor U2023 (N_2023,N_1766,N_1593);
and U2024 (N_2024,N_1923,N_1539);
and U2025 (N_2025,N_1821,N_1913);
nor U2026 (N_2026,N_1559,N_1894);
xnor U2027 (N_2027,N_1504,N_1815);
nor U2028 (N_2028,N_1934,N_1951);
and U2029 (N_2029,N_1690,N_1881);
nor U2030 (N_2030,N_1626,N_1942);
and U2031 (N_2031,N_1789,N_1813);
nand U2032 (N_2032,N_1850,N_1935);
xor U2033 (N_2033,N_1891,N_1730);
nand U2034 (N_2034,N_1557,N_1955);
and U2035 (N_2035,N_1695,N_1633);
and U2036 (N_2036,N_1975,N_1674);
nor U2037 (N_2037,N_1886,N_1737);
xnor U2038 (N_2038,N_1954,N_1558);
nor U2039 (N_2039,N_1572,N_1851);
nand U2040 (N_2040,N_1920,N_1973);
nand U2041 (N_2041,N_1936,N_1926);
or U2042 (N_2042,N_1883,N_1738);
xnor U2043 (N_2043,N_1782,N_1908);
nor U2044 (N_2044,N_1664,N_1711);
nor U2045 (N_2045,N_1796,N_1909);
xnor U2046 (N_2046,N_1616,N_1617);
nand U2047 (N_2047,N_1888,N_1986);
nor U2048 (N_2048,N_1609,N_1587);
nand U2049 (N_2049,N_1535,N_1571);
nor U2050 (N_2050,N_1677,N_1682);
or U2051 (N_2051,N_1567,N_1755);
xor U2052 (N_2052,N_1892,N_1748);
nand U2053 (N_2053,N_1550,N_1545);
and U2054 (N_2054,N_1667,N_1692);
or U2055 (N_2055,N_1594,N_1702);
and U2056 (N_2056,N_1924,N_1671);
and U2057 (N_2057,N_1739,N_1778);
nor U2058 (N_2058,N_1732,N_1689);
and U2059 (N_2059,N_1719,N_1928);
nand U2060 (N_2060,N_1591,N_1548);
and U2061 (N_2061,N_1600,N_1549);
or U2062 (N_2062,N_1808,N_1735);
or U2063 (N_2063,N_1864,N_1956);
or U2064 (N_2064,N_1861,N_1612);
xnor U2065 (N_2065,N_1925,N_1641);
nor U2066 (N_2066,N_1585,N_1752);
nand U2067 (N_2067,N_1902,N_1663);
nor U2068 (N_2068,N_1912,N_1699);
and U2069 (N_2069,N_1510,N_1790);
and U2070 (N_2070,N_1862,N_1709);
nand U2071 (N_2071,N_1503,N_1791);
and U2072 (N_2072,N_1827,N_1803);
or U2073 (N_2073,N_1983,N_1994);
xnor U2074 (N_2074,N_1939,N_1987);
xor U2075 (N_2075,N_1854,N_1871);
and U2076 (N_2076,N_1577,N_1524);
or U2077 (N_2077,N_1635,N_1823);
and U2078 (N_2078,N_1642,N_1687);
and U2079 (N_2079,N_1844,N_1670);
nand U2080 (N_2080,N_1625,N_1999);
xnor U2081 (N_2081,N_1775,N_1884);
or U2082 (N_2082,N_1905,N_1965);
nor U2083 (N_2083,N_1753,N_1688);
and U2084 (N_2084,N_1964,N_1847);
and U2085 (N_2085,N_1977,N_1798);
xnor U2086 (N_2086,N_1565,N_1606);
and U2087 (N_2087,N_1756,N_1929);
xor U2088 (N_2088,N_1763,N_1876);
xor U2089 (N_2089,N_1582,N_1650);
and U2090 (N_2090,N_1804,N_1713);
or U2091 (N_2091,N_1529,N_1959);
xor U2092 (N_2092,N_1976,N_1624);
or U2093 (N_2093,N_1904,N_1957);
and U2094 (N_2094,N_1696,N_1982);
and U2095 (N_2095,N_1793,N_1527);
and U2096 (N_2096,N_1556,N_1684);
xnor U2097 (N_2097,N_1710,N_1607);
and U2098 (N_2098,N_1774,N_1859);
and U2099 (N_2099,N_1786,N_1648);
nand U2100 (N_2100,N_1508,N_1686);
or U2101 (N_2101,N_1907,N_1873);
nand U2102 (N_2102,N_1817,N_1511);
or U2103 (N_2103,N_1849,N_1801);
and U2104 (N_2104,N_1980,N_1613);
or U2105 (N_2105,N_1656,N_1678);
or U2106 (N_2106,N_1564,N_1802);
nor U2107 (N_2107,N_1501,N_1903);
and U2108 (N_2108,N_1836,N_1744);
nand U2109 (N_2109,N_1509,N_1727);
or U2110 (N_2110,N_1967,N_1537);
or U2111 (N_2111,N_1889,N_1809);
and U2112 (N_2112,N_1552,N_1521);
or U2113 (N_2113,N_1516,N_1820);
nand U2114 (N_2114,N_1771,N_1971);
nor U2115 (N_2115,N_1754,N_1704);
or U2116 (N_2116,N_1953,N_1887);
nand U2117 (N_2117,N_1570,N_1874);
nor U2118 (N_2118,N_1728,N_1749);
nand U2119 (N_2119,N_1855,N_1691);
or U2120 (N_2120,N_1518,N_1734);
nand U2121 (N_2121,N_1882,N_1672);
nor U2122 (N_2122,N_1541,N_1870);
xnor U2123 (N_2123,N_1531,N_1584);
and U2124 (N_2124,N_1543,N_1831);
nand U2125 (N_2125,N_1566,N_1940);
xnor U2126 (N_2126,N_1603,N_1825);
or U2127 (N_2127,N_1588,N_1840);
or U2128 (N_2128,N_1742,N_1758);
nand U2129 (N_2129,N_1512,N_1828);
and U2130 (N_2130,N_1769,N_1937);
xnor U2131 (N_2131,N_1901,N_1602);
or U2132 (N_2132,N_1921,N_1919);
and U2133 (N_2133,N_1736,N_1833);
nand U2134 (N_2134,N_1917,N_1860);
and U2135 (N_2135,N_1898,N_1636);
or U2136 (N_2136,N_1914,N_1899);
nor U2137 (N_2137,N_1597,N_1997);
or U2138 (N_2138,N_1931,N_1880);
nor U2139 (N_2139,N_1797,N_1569);
xor U2140 (N_2140,N_1995,N_1822);
or U2141 (N_2141,N_1826,N_1877);
nor U2142 (N_2142,N_1694,N_1949);
or U2143 (N_2143,N_1507,N_1819);
nand U2144 (N_2144,N_1845,N_1596);
xor U2145 (N_2145,N_1563,N_1772);
nor U2146 (N_2146,N_1519,N_1513);
or U2147 (N_2147,N_1867,N_1974);
or U2148 (N_2148,N_1653,N_1779);
nand U2149 (N_2149,N_1500,N_1578);
nand U2150 (N_2150,N_1818,N_1731);
nand U2151 (N_2151,N_1573,N_1720);
xnor U2152 (N_2152,N_1614,N_1795);
nand U2153 (N_2153,N_1705,N_1794);
nor U2154 (N_2154,N_1673,N_1890);
or U2155 (N_2155,N_1792,N_1536);
nand U2156 (N_2156,N_1698,N_1969);
or U2157 (N_2157,N_1996,N_1832);
and U2158 (N_2158,N_1645,N_1978);
or U2159 (N_2159,N_1979,N_1824);
nand U2160 (N_2160,N_1858,N_1878);
nand U2161 (N_2161,N_1989,N_1628);
xor U2162 (N_2162,N_1576,N_1595);
and U2163 (N_2163,N_1598,N_1679);
nor U2164 (N_2164,N_1740,N_1788);
and U2165 (N_2165,N_1647,N_1812);
nor U2166 (N_2166,N_1623,N_1843);
or U2167 (N_2167,N_1560,N_1781);
nor U2168 (N_2168,N_1837,N_1733);
xor U2169 (N_2169,N_1586,N_1528);
or U2170 (N_2170,N_1872,N_1768);
xnor U2171 (N_2171,N_1634,N_1896);
nor U2172 (N_2172,N_1985,N_1780);
xor U2173 (N_2173,N_1746,N_1723);
nand U2174 (N_2174,N_1665,N_1717);
nor U2175 (N_2175,N_1660,N_1649);
and U2176 (N_2176,N_1601,N_1640);
nor U2177 (N_2177,N_1685,N_1750);
xor U2178 (N_2178,N_1885,N_1842);
nand U2179 (N_2179,N_1950,N_1522);
or U2180 (N_2180,N_1589,N_1922);
nand U2181 (N_2181,N_1972,N_1579);
nor U2182 (N_2182,N_1651,N_1968);
nand U2183 (N_2183,N_1800,N_1806);
nor U2184 (N_2184,N_1866,N_1773);
nor U2185 (N_2185,N_1963,N_1608);
nor U2186 (N_2186,N_1703,N_1910);
nand U2187 (N_2187,N_1676,N_1683);
or U2188 (N_2188,N_1960,N_1643);
and U2189 (N_2189,N_1532,N_1525);
xor U2190 (N_2190,N_1533,N_1941);
nor U2191 (N_2191,N_1852,N_1631);
or U2192 (N_2192,N_1875,N_1865);
or U2193 (N_2193,N_1810,N_1610);
and U2194 (N_2194,N_1622,N_1918);
or U2195 (N_2195,N_1745,N_1574);
nand U2196 (N_2196,N_1943,N_1627);
xnor U2197 (N_2197,N_1544,N_1799);
nand U2198 (N_2198,N_1988,N_1857);
nor U2199 (N_2199,N_1805,N_1654);
nand U2200 (N_2200,N_1834,N_1946);
xnor U2201 (N_2201,N_1930,N_1835);
xnor U2202 (N_2202,N_1743,N_1615);
or U2203 (N_2203,N_1657,N_1970);
and U2204 (N_2204,N_1583,N_1757);
and U2205 (N_2205,N_1555,N_1990);
or U2206 (N_2206,N_1697,N_1816);
nor U2207 (N_2207,N_1729,N_1915);
xnor U2208 (N_2208,N_1944,N_1515);
nand U2209 (N_2209,N_1680,N_1581);
and U2210 (N_2210,N_1893,N_1947);
nand U2211 (N_2211,N_1592,N_1658);
nand U2212 (N_2212,N_1741,N_1952);
nor U2213 (N_2213,N_1785,N_1726);
nor U2214 (N_2214,N_1945,N_1715);
nor U2215 (N_2215,N_1718,N_1681);
or U2216 (N_2216,N_1669,N_1652);
or U2217 (N_2217,N_1646,N_1722);
and U2218 (N_2218,N_1767,N_1932);
and U2219 (N_2219,N_1604,N_1853);
or U2220 (N_2220,N_1611,N_1762);
and U2221 (N_2221,N_1784,N_1506);
xnor U2222 (N_2222,N_1747,N_1759);
nand U2223 (N_2223,N_1639,N_1590);
nand U2224 (N_2224,N_1991,N_1554);
nand U2225 (N_2225,N_1551,N_1700);
nor U2226 (N_2226,N_1505,N_1829);
nand U2227 (N_2227,N_1751,N_1906);
nand U2228 (N_2228,N_1839,N_1830);
nor U2229 (N_2229,N_1927,N_1553);
or U2230 (N_2230,N_1846,N_1787);
nand U2231 (N_2231,N_1538,N_1962);
and U2232 (N_2232,N_1637,N_1580);
and U2233 (N_2233,N_1721,N_1895);
nor U2234 (N_2234,N_1644,N_1811);
nand U2235 (N_2235,N_1502,N_1765);
and U2236 (N_2236,N_1575,N_1897);
or U2237 (N_2237,N_1958,N_1848);
nand U2238 (N_2238,N_1530,N_1938);
or U2239 (N_2239,N_1966,N_1523);
and U2240 (N_2240,N_1666,N_1725);
or U2241 (N_2241,N_1618,N_1916);
and U2242 (N_2242,N_1770,N_1661);
nand U2243 (N_2243,N_1856,N_1807);
or U2244 (N_2244,N_1879,N_1599);
and U2245 (N_2245,N_1630,N_1911);
nor U2246 (N_2246,N_1629,N_1662);
nand U2247 (N_2247,N_1981,N_1777);
nor U2248 (N_2248,N_1619,N_1675);
and U2249 (N_2249,N_1520,N_1546);
xor U2250 (N_2250,N_1607,N_1796);
nor U2251 (N_2251,N_1993,N_1523);
and U2252 (N_2252,N_1998,N_1648);
and U2253 (N_2253,N_1548,N_1531);
nand U2254 (N_2254,N_1587,N_1781);
xnor U2255 (N_2255,N_1970,N_1528);
nor U2256 (N_2256,N_1659,N_1501);
and U2257 (N_2257,N_1564,N_1752);
or U2258 (N_2258,N_1659,N_1897);
nor U2259 (N_2259,N_1574,N_1655);
nor U2260 (N_2260,N_1900,N_1875);
and U2261 (N_2261,N_1830,N_1758);
or U2262 (N_2262,N_1640,N_1681);
nand U2263 (N_2263,N_1562,N_1722);
or U2264 (N_2264,N_1621,N_1869);
nor U2265 (N_2265,N_1890,N_1964);
xnor U2266 (N_2266,N_1511,N_1926);
nor U2267 (N_2267,N_1926,N_1554);
nand U2268 (N_2268,N_1844,N_1897);
xnor U2269 (N_2269,N_1911,N_1823);
nor U2270 (N_2270,N_1741,N_1837);
or U2271 (N_2271,N_1927,N_1694);
and U2272 (N_2272,N_1949,N_1839);
nand U2273 (N_2273,N_1702,N_1751);
nand U2274 (N_2274,N_1796,N_1676);
nor U2275 (N_2275,N_1580,N_1861);
nand U2276 (N_2276,N_1568,N_1961);
nor U2277 (N_2277,N_1886,N_1563);
and U2278 (N_2278,N_1562,N_1745);
xnor U2279 (N_2279,N_1883,N_1835);
xnor U2280 (N_2280,N_1961,N_1721);
nand U2281 (N_2281,N_1943,N_1967);
nand U2282 (N_2282,N_1687,N_1734);
and U2283 (N_2283,N_1854,N_1914);
or U2284 (N_2284,N_1724,N_1906);
or U2285 (N_2285,N_1769,N_1837);
or U2286 (N_2286,N_1776,N_1621);
and U2287 (N_2287,N_1720,N_1887);
nor U2288 (N_2288,N_1610,N_1631);
nand U2289 (N_2289,N_1959,N_1952);
and U2290 (N_2290,N_1631,N_1834);
or U2291 (N_2291,N_1977,N_1795);
or U2292 (N_2292,N_1823,N_1774);
nand U2293 (N_2293,N_1513,N_1582);
xor U2294 (N_2294,N_1629,N_1540);
and U2295 (N_2295,N_1674,N_1958);
xnor U2296 (N_2296,N_1553,N_1731);
and U2297 (N_2297,N_1797,N_1933);
or U2298 (N_2298,N_1947,N_1839);
and U2299 (N_2299,N_1671,N_1599);
nor U2300 (N_2300,N_1928,N_1950);
nor U2301 (N_2301,N_1608,N_1813);
and U2302 (N_2302,N_1501,N_1565);
nor U2303 (N_2303,N_1864,N_1850);
nor U2304 (N_2304,N_1980,N_1644);
nand U2305 (N_2305,N_1668,N_1734);
or U2306 (N_2306,N_1778,N_1587);
nor U2307 (N_2307,N_1694,N_1801);
nand U2308 (N_2308,N_1517,N_1985);
or U2309 (N_2309,N_1816,N_1807);
and U2310 (N_2310,N_1517,N_1639);
xor U2311 (N_2311,N_1893,N_1781);
or U2312 (N_2312,N_1695,N_1946);
xnor U2313 (N_2313,N_1920,N_1588);
nor U2314 (N_2314,N_1559,N_1789);
nand U2315 (N_2315,N_1936,N_1802);
nor U2316 (N_2316,N_1675,N_1609);
or U2317 (N_2317,N_1943,N_1925);
and U2318 (N_2318,N_1516,N_1550);
nor U2319 (N_2319,N_1852,N_1885);
nand U2320 (N_2320,N_1742,N_1525);
or U2321 (N_2321,N_1618,N_1712);
nor U2322 (N_2322,N_1870,N_1732);
nor U2323 (N_2323,N_1969,N_1528);
nand U2324 (N_2324,N_1921,N_1906);
and U2325 (N_2325,N_1573,N_1619);
nor U2326 (N_2326,N_1942,N_1904);
or U2327 (N_2327,N_1934,N_1513);
nor U2328 (N_2328,N_1616,N_1560);
nor U2329 (N_2329,N_1585,N_1587);
nand U2330 (N_2330,N_1678,N_1664);
xnor U2331 (N_2331,N_1841,N_1630);
nand U2332 (N_2332,N_1909,N_1532);
and U2333 (N_2333,N_1711,N_1602);
nor U2334 (N_2334,N_1622,N_1747);
and U2335 (N_2335,N_1531,N_1971);
nand U2336 (N_2336,N_1552,N_1882);
nand U2337 (N_2337,N_1677,N_1570);
nor U2338 (N_2338,N_1786,N_1882);
nor U2339 (N_2339,N_1757,N_1910);
nand U2340 (N_2340,N_1599,N_1757);
xor U2341 (N_2341,N_1833,N_1864);
or U2342 (N_2342,N_1537,N_1503);
nand U2343 (N_2343,N_1855,N_1804);
or U2344 (N_2344,N_1862,N_1810);
or U2345 (N_2345,N_1886,N_1622);
nand U2346 (N_2346,N_1625,N_1969);
nor U2347 (N_2347,N_1555,N_1580);
nand U2348 (N_2348,N_1563,N_1810);
nand U2349 (N_2349,N_1762,N_1706);
nor U2350 (N_2350,N_1919,N_1816);
nand U2351 (N_2351,N_1854,N_1654);
or U2352 (N_2352,N_1907,N_1502);
and U2353 (N_2353,N_1524,N_1941);
xnor U2354 (N_2354,N_1857,N_1837);
or U2355 (N_2355,N_1593,N_1725);
nand U2356 (N_2356,N_1858,N_1589);
nand U2357 (N_2357,N_1804,N_1872);
or U2358 (N_2358,N_1536,N_1627);
and U2359 (N_2359,N_1670,N_1750);
nor U2360 (N_2360,N_1591,N_1690);
nand U2361 (N_2361,N_1778,N_1940);
nand U2362 (N_2362,N_1552,N_1846);
xnor U2363 (N_2363,N_1663,N_1529);
nor U2364 (N_2364,N_1669,N_1808);
nand U2365 (N_2365,N_1668,N_1557);
nor U2366 (N_2366,N_1545,N_1554);
and U2367 (N_2367,N_1713,N_1781);
nand U2368 (N_2368,N_1584,N_1788);
and U2369 (N_2369,N_1995,N_1520);
or U2370 (N_2370,N_1898,N_1579);
or U2371 (N_2371,N_1945,N_1888);
or U2372 (N_2372,N_1734,N_1502);
xor U2373 (N_2373,N_1863,N_1574);
nand U2374 (N_2374,N_1934,N_1843);
nand U2375 (N_2375,N_1749,N_1994);
or U2376 (N_2376,N_1704,N_1516);
and U2377 (N_2377,N_1573,N_1811);
and U2378 (N_2378,N_1784,N_1981);
nand U2379 (N_2379,N_1727,N_1994);
and U2380 (N_2380,N_1522,N_1564);
nor U2381 (N_2381,N_1663,N_1759);
nor U2382 (N_2382,N_1872,N_1963);
or U2383 (N_2383,N_1627,N_1663);
nor U2384 (N_2384,N_1502,N_1926);
and U2385 (N_2385,N_1749,N_1561);
or U2386 (N_2386,N_1650,N_1555);
or U2387 (N_2387,N_1829,N_1640);
xor U2388 (N_2388,N_1815,N_1569);
nor U2389 (N_2389,N_1683,N_1822);
and U2390 (N_2390,N_1550,N_1508);
and U2391 (N_2391,N_1572,N_1999);
and U2392 (N_2392,N_1743,N_1955);
nor U2393 (N_2393,N_1943,N_1551);
nand U2394 (N_2394,N_1840,N_1632);
xnor U2395 (N_2395,N_1792,N_1946);
xnor U2396 (N_2396,N_1508,N_1514);
or U2397 (N_2397,N_1598,N_1803);
nand U2398 (N_2398,N_1800,N_1638);
or U2399 (N_2399,N_1911,N_1644);
and U2400 (N_2400,N_1784,N_1601);
nor U2401 (N_2401,N_1552,N_1873);
nand U2402 (N_2402,N_1674,N_1951);
nor U2403 (N_2403,N_1811,N_1769);
xor U2404 (N_2404,N_1551,N_1812);
or U2405 (N_2405,N_1656,N_1699);
or U2406 (N_2406,N_1660,N_1900);
or U2407 (N_2407,N_1864,N_1737);
or U2408 (N_2408,N_1889,N_1742);
and U2409 (N_2409,N_1947,N_1621);
and U2410 (N_2410,N_1995,N_1800);
and U2411 (N_2411,N_1999,N_1771);
nor U2412 (N_2412,N_1635,N_1632);
or U2413 (N_2413,N_1880,N_1530);
xor U2414 (N_2414,N_1619,N_1827);
and U2415 (N_2415,N_1747,N_1987);
xnor U2416 (N_2416,N_1515,N_1666);
nor U2417 (N_2417,N_1565,N_1720);
or U2418 (N_2418,N_1893,N_1875);
or U2419 (N_2419,N_1593,N_1590);
nor U2420 (N_2420,N_1810,N_1627);
nand U2421 (N_2421,N_1899,N_1848);
or U2422 (N_2422,N_1564,N_1989);
nor U2423 (N_2423,N_1943,N_1855);
nand U2424 (N_2424,N_1664,N_1730);
or U2425 (N_2425,N_1611,N_1966);
nor U2426 (N_2426,N_1871,N_1923);
and U2427 (N_2427,N_1885,N_1820);
nor U2428 (N_2428,N_1927,N_1906);
nand U2429 (N_2429,N_1836,N_1802);
nor U2430 (N_2430,N_1523,N_1810);
and U2431 (N_2431,N_1707,N_1734);
and U2432 (N_2432,N_1553,N_1804);
xnor U2433 (N_2433,N_1905,N_1858);
nand U2434 (N_2434,N_1715,N_1506);
nor U2435 (N_2435,N_1544,N_1641);
and U2436 (N_2436,N_1978,N_1739);
nand U2437 (N_2437,N_1563,N_1661);
and U2438 (N_2438,N_1913,N_1797);
nor U2439 (N_2439,N_1520,N_1715);
xnor U2440 (N_2440,N_1770,N_1645);
nor U2441 (N_2441,N_1538,N_1875);
and U2442 (N_2442,N_1684,N_1746);
or U2443 (N_2443,N_1873,N_1719);
or U2444 (N_2444,N_1853,N_1521);
xor U2445 (N_2445,N_1628,N_1650);
nor U2446 (N_2446,N_1693,N_1748);
nor U2447 (N_2447,N_1810,N_1541);
nand U2448 (N_2448,N_1829,N_1848);
nand U2449 (N_2449,N_1967,N_1876);
and U2450 (N_2450,N_1692,N_1722);
or U2451 (N_2451,N_1919,N_1650);
or U2452 (N_2452,N_1740,N_1608);
or U2453 (N_2453,N_1581,N_1750);
nor U2454 (N_2454,N_1726,N_1925);
nand U2455 (N_2455,N_1534,N_1516);
and U2456 (N_2456,N_1800,N_1879);
nor U2457 (N_2457,N_1791,N_1748);
xor U2458 (N_2458,N_1870,N_1798);
and U2459 (N_2459,N_1636,N_1751);
nand U2460 (N_2460,N_1527,N_1827);
nand U2461 (N_2461,N_1784,N_1812);
or U2462 (N_2462,N_1527,N_1736);
nor U2463 (N_2463,N_1842,N_1900);
nor U2464 (N_2464,N_1557,N_1700);
nand U2465 (N_2465,N_1989,N_1717);
nand U2466 (N_2466,N_1979,N_1923);
and U2467 (N_2467,N_1843,N_1738);
nand U2468 (N_2468,N_1829,N_1961);
nand U2469 (N_2469,N_1519,N_1885);
or U2470 (N_2470,N_1770,N_1653);
nand U2471 (N_2471,N_1933,N_1781);
or U2472 (N_2472,N_1915,N_1514);
or U2473 (N_2473,N_1822,N_1703);
and U2474 (N_2474,N_1944,N_1689);
xnor U2475 (N_2475,N_1728,N_1929);
or U2476 (N_2476,N_1958,N_1524);
and U2477 (N_2477,N_1575,N_1880);
or U2478 (N_2478,N_1902,N_1606);
xor U2479 (N_2479,N_1949,N_1989);
and U2480 (N_2480,N_1797,N_1522);
nor U2481 (N_2481,N_1666,N_1755);
or U2482 (N_2482,N_1944,N_1660);
and U2483 (N_2483,N_1882,N_1947);
or U2484 (N_2484,N_1926,N_1969);
or U2485 (N_2485,N_1669,N_1500);
xnor U2486 (N_2486,N_1918,N_1550);
xor U2487 (N_2487,N_1910,N_1587);
or U2488 (N_2488,N_1547,N_1854);
xor U2489 (N_2489,N_1831,N_1507);
nand U2490 (N_2490,N_1631,N_1988);
or U2491 (N_2491,N_1545,N_1566);
and U2492 (N_2492,N_1819,N_1845);
and U2493 (N_2493,N_1543,N_1732);
xnor U2494 (N_2494,N_1521,N_1956);
xnor U2495 (N_2495,N_1541,N_1844);
nor U2496 (N_2496,N_1888,N_1703);
xor U2497 (N_2497,N_1810,N_1811);
or U2498 (N_2498,N_1864,N_1545);
nor U2499 (N_2499,N_1814,N_1500);
nor U2500 (N_2500,N_2320,N_2352);
or U2501 (N_2501,N_2351,N_2417);
nand U2502 (N_2502,N_2424,N_2202);
and U2503 (N_2503,N_2107,N_2201);
nand U2504 (N_2504,N_2440,N_2458);
nor U2505 (N_2505,N_2270,N_2473);
or U2506 (N_2506,N_2355,N_2476);
nor U2507 (N_2507,N_2260,N_2442);
and U2508 (N_2508,N_2124,N_2447);
and U2509 (N_2509,N_2113,N_2378);
and U2510 (N_2510,N_2361,N_2380);
nand U2511 (N_2511,N_2388,N_2077);
nor U2512 (N_2512,N_2171,N_2407);
nand U2513 (N_2513,N_2478,N_2266);
nand U2514 (N_2514,N_2446,N_2136);
and U2515 (N_2515,N_2411,N_2108);
or U2516 (N_2516,N_2335,N_2105);
and U2517 (N_2517,N_2340,N_2034);
or U2518 (N_2518,N_2200,N_2032);
and U2519 (N_2519,N_2049,N_2131);
and U2520 (N_2520,N_2252,N_2382);
and U2521 (N_2521,N_2120,N_2204);
nor U2522 (N_2522,N_2371,N_2375);
nand U2523 (N_2523,N_2373,N_2233);
nor U2524 (N_2524,N_2067,N_2481);
nor U2525 (N_2525,N_2064,N_2017);
nor U2526 (N_2526,N_2474,N_2291);
nand U2527 (N_2527,N_2228,N_2236);
or U2528 (N_2528,N_2285,N_2438);
and U2529 (N_2529,N_2104,N_2413);
nor U2530 (N_2530,N_2102,N_2237);
xor U2531 (N_2531,N_2428,N_2086);
or U2532 (N_2532,N_2144,N_2357);
and U2533 (N_2533,N_2448,N_2353);
xor U2534 (N_2534,N_2044,N_2268);
nor U2535 (N_2535,N_2115,N_2039);
and U2536 (N_2536,N_2000,N_2287);
xor U2537 (N_2537,N_2362,N_2129);
nor U2538 (N_2538,N_2274,N_2301);
nor U2539 (N_2539,N_2379,N_2364);
and U2540 (N_2540,N_2385,N_2170);
and U2541 (N_2541,N_2167,N_2246);
nor U2542 (N_2542,N_2217,N_2394);
nand U2543 (N_2543,N_2145,N_2484);
or U2544 (N_2544,N_2042,N_2057);
nor U2545 (N_2545,N_2321,N_2384);
or U2546 (N_2546,N_2306,N_2265);
xor U2547 (N_2547,N_2273,N_2479);
nor U2548 (N_2548,N_2213,N_2269);
nor U2549 (N_2549,N_2035,N_2486);
or U2550 (N_2550,N_2023,N_2106);
or U2551 (N_2551,N_2467,N_2307);
and U2552 (N_2552,N_2232,N_2336);
nand U2553 (N_2553,N_2283,N_2020);
xor U2554 (N_2554,N_2047,N_2286);
nor U2555 (N_2555,N_2161,N_2162);
or U2556 (N_2556,N_2038,N_2419);
nand U2557 (N_2557,N_2189,N_2396);
and U2558 (N_2558,N_2368,N_2156);
nand U2559 (N_2559,N_2416,N_2096);
and U2560 (N_2560,N_2464,N_2303);
or U2561 (N_2561,N_2408,N_2322);
xor U2562 (N_2562,N_2358,N_2101);
nand U2563 (N_2563,N_2249,N_2247);
nor U2564 (N_2564,N_2346,N_2400);
nand U2565 (N_2565,N_2074,N_2463);
nand U2566 (N_2566,N_2429,N_2130);
or U2567 (N_2567,N_2480,N_2281);
and U2568 (N_2568,N_2278,N_2192);
and U2569 (N_2569,N_2312,N_2126);
and U2570 (N_2570,N_2215,N_2051);
nand U2571 (N_2571,N_2060,N_2127);
and U2572 (N_2572,N_2316,N_2152);
nor U2573 (N_2573,N_2001,N_2002);
or U2574 (N_2574,N_2433,N_2423);
or U2575 (N_2575,N_2079,N_2172);
or U2576 (N_2576,N_2100,N_2179);
nor U2577 (N_2577,N_2025,N_2040);
nor U2578 (N_2578,N_2142,N_2469);
and U2579 (N_2579,N_2177,N_2212);
xor U2580 (N_2580,N_2453,N_2289);
xor U2581 (N_2581,N_2435,N_2462);
xor U2582 (N_2582,N_2327,N_2333);
xor U2583 (N_2583,N_2391,N_2191);
or U2584 (N_2584,N_2461,N_2186);
nor U2585 (N_2585,N_2043,N_2495);
nor U2586 (N_2586,N_2185,N_2205);
or U2587 (N_2587,N_2445,N_2359);
nand U2588 (N_2588,N_2016,N_2045);
nor U2589 (N_2589,N_2477,N_2377);
nand U2590 (N_2590,N_2451,N_2354);
and U2591 (N_2591,N_2006,N_2147);
and U2592 (N_2592,N_2493,N_2311);
and U2593 (N_2593,N_2482,N_2343);
nand U2594 (N_2594,N_2157,N_2313);
nand U2595 (N_2595,N_2024,N_2367);
nand U2596 (N_2596,N_2135,N_2392);
nand U2597 (N_2597,N_2255,N_2374);
and U2598 (N_2598,N_2123,N_2398);
and U2599 (N_2599,N_2084,N_2360);
xnor U2600 (N_2600,N_2347,N_2138);
xnor U2601 (N_2601,N_2250,N_2342);
nand U2602 (N_2602,N_2279,N_2422);
or U2603 (N_2603,N_2095,N_2363);
and U2604 (N_2604,N_2436,N_2224);
or U2605 (N_2605,N_2365,N_2053);
xor U2606 (N_2606,N_2018,N_2409);
xnor U2607 (N_2607,N_2366,N_2248);
xor U2608 (N_2608,N_2028,N_2219);
or U2609 (N_2609,N_2206,N_2103);
xnor U2610 (N_2610,N_2421,N_2284);
or U2611 (N_2611,N_2091,N_2082);
xor U2612 (N_2612,N_2022,N_2395);
and U2613 (N_2613,N_2198,N_2176);
nand U2614 (N_2614,N_2425,N_2376);
and U2615 (N_2615,N_2491,N_2323);
and U2616 (N_2616,N_2386,N_2207);
xor U2617 (N_2617,N_2406,N_2116);
nand U2618 (N_2618,N_2263,N_2071);
nand U2619 (N_2619,N_2261,N_2004);
nor U2620 (N_2620,N_2262,N_2121);
nor U2621 (N_2621,N_2099,N_2166);
nor U2622 (N_2622,N_2339,N_2065);
nand U2623 (N_2623,N_2210,N_2036);
nor U2624 (N_2624,N_2292,N_2180);
nand U2625 (N_2625,N_2221,N_2143);
xnor U2626 (N_2626,N_2399,N_2117);
nand U2627 (N_2627,N_2208,N_2056);
nor U2628 (N_2628,N_2093,N_2090);
nor U2629 (N_2629,N_2146,N_2452);
and U2630 (N_2630,N_2370,N_2280);
nand U2631 (N_2631,N_2154,N_2488);
nor U2632 (N_2632,N_2401,N_2196);
nand U2633 (N_2633,N_2194,N_2439);
or U2634 (N_2634,N_2489,N_2070);
xor U2635 (N_2635,N_2405,N_2112);
or U2636 (N_2636,N_2173,N_2111);
and U2637 (N_2637,N_2348,N_2150);
nand U2638 (N_2638,N_2139,N_2133);
and U2639 (N_2639,N_2220,N_2432);
and U2640 (N_2640,N_2223,N_2345);
nor U2641 (N_2641,N_2149,N_2331);
or U2642 (N_2642,N_2037,N_2188);
and U2643 (N_2643,N_2054,N_2456);
or U2644 (N_2644,N_2328,N_2471);
and U2645 (N_2645,N_2193,N_2109);
nand U2646 (N_2646,N_2089,N_2454);
or U2647 (N_2647,N_2465,N_2141);
nor U2648 (N_2648,N_2197,N_2159);
and U2649 (N_2649,N_2072,N_2497);
xor U2650 (N_2650,N_2169,N_2470);
nand U2651 (N_2651,N_2329,N_2257);
or U2652 (N_2652,N_2402,N_2258);
and U2653 (N_2653,N_2238,N_2087);
xnor U2654 (N_2654,N_2277,N_2492);
or U2655 (N_2655,N_2183,N_2098);
or U2656 (N_2656,N_2350,N_2021);
or U2657 (N_2657,N_2325,N_2317);
nor U2658 (N_2658,N_2076,N_2330);
or U2659 (N_2659,N_2012,N_2326);
and U2660 (N_2660,N_2460,N_2231);
nor U2661 (N_2661,N_2472,N_2441);
and U2662 (N_2662,N_2068,N_2390);
xor U2663 (N_2663,N_2387,N_2005);
nor U2664 (N_2664,N_2319,N_2214);
and U2665 (N_2665,N_2181,N_2218);
or U2666 (N_2666,N_2305,N_2097);
or U2667 (N_2667,N_2052,N_2008);
or U2668 (N_2668,N_2494,N_2349);
xor U2669 (N_2669,N_2485,N_2299);
nand U2670 (N_2670,N_2443,N_2055);
and U2671 (N_2671,N_2059,N_2013);
nand U2672 (N_2672,N_2222,N_2455);
or U2673 (N_2673,N_2209,N_2468);
xor U2674 (N_2674,N_2226,N_2094);
nand U2675 (N_2675,N_2080,N_2088);
and U2676 (N_2676,N_2073,N_2341);
and U2677 (N_2677,N_2264,N_2225);
or U2678 (N_2678,N_2404,N_2069);
and U2679 (N_2679,N_2164,N_2254);
nand U2680 (N_2680,N_2487,N_2414);
nand U2681 (N_2681,N_2203,N_2412);
xor U2682 (N_2682,N_2431,N_2128);
or U2683 (N_2683,N_2244,N_2410);
and U2684 (N_2684,N_2083,N_2010);
nor U2685 (N_2685,N_2163,N_2048);
and U2686 (N_2686,N_2490,N_2014);
and U2687 (N_2687,N_2061,N_2256);
or U2688 (N_2688,N_2062,N_2383);
nor U2689 (N_2689,N_2403,N_2230);
nand U2690 (N_2690,N_2216,N_2075);
or U2691 (N_2691,N_2430,N_2160);
or U2692 (N_2692,N_2174,N_2397);
and U2693 (N_2693,N_2199,N_2243);
nand U2694 (N_2694,N_2011,N_2334);
nand U2695 (N_2695,N_2148,N_2239);
nor U2696 (N_2696,N_2125,N_2134);
nor U2697 (N_2697,N_2332,N_2033);
nor U2698 (N_2698,N_2081,N_2276);
and U2699 (N_2699,N_2066,N_2019);
nor U2700 (N_2700,N_2168,N_2466);
or U2701 (N_2701,N_2003,N_2031);
nor U2702 (N_2702,N_2415,N_2297);
nand U2703 (N_2703,N_2119,N_2229);
nand U2704 (N_2704,N_2434,N_2184);
nand U2705 (N_2705,N_2251,N_2498);
or U2706 (N_2706,N_2381,N_2240);
nand U2707 (N_2707,N_2063,N_2393);
nand U2708 (N_2708,N_2300,N_2241);
nand U2709 (N_2709,N_2450,N_2195);
or U2710 (N_2710,N_2227,N_2211);
or U2711 (N_2711,N_2437,N_2483);
nor U2712 (N_2712,N_2137,N_2151);
or U2713 (N_2713,N_2175,N_2182);
or U2714 (N_2714,N_2110,N_2058);
or U2715 (N_2715,N_2132,N_2308);
nor U2716 (N_2716,N_2318,N_2309);
nor U2717 (N_2717,N_2449,N_2294);
or U2718 (N_2718,N_2140,N_2027);
nand U2719 (N_2719,N_2389,N_2253);
or U2720 (N_2720,N_2041,N_2457);
or U2721 (N_2721,N_2118,N_2271);
nor U2722 (N_2722,N_2496,N_2372);
nand U2723 (N_2723,N_2030,N_2007);
nor U2724 (N_2724,N_2298,N_2272);
nand U2725 (N_2725,N_2085,N_2302);
nand U2726 (N_2726,N_2499,N_2078);
and U2727 (N_2727,N_2234,N_2245);
nor U2728 (N_2728,N_2344,N_2296);
and U2729 (N_2729,N_2282,N_2242);
and U2730 (N_2730,N_2259,N_2295);
or U2731 (N_2731,N_2337,N_2475);
xor U2732 (N_2732,N_2459,N_2288);
nor U2733 (N_2733,N_2293,N_2114);
and U2734 (N_2734,N_2275,N_2324);
nand U2735 (N_2735,N_2009,N_2235);
nand U2736 (N_2736,N_2290,N_2338);
or U2737 (N_2737,N_2369,N_2310);
xor U2738 (N_2738,N_2015,N_2122);
and U2739 (N_2739,N_2427,N_2165);
or U2740 (N_2740,N_2092,N_2026);
nor U2741 (N_2741,N_2153,N_2444);
xnor U2742 (N_2742,N_2314,N_2046);
or U2743 (N_2743,N_2356,N_2155);
and U2744 (N_2744,N_2158,N_2304);
xnor U2745 (N_2745,N_2315,N_2187);
and U2746 (N_2746,N_2190,N_2420);
xor U2747 (N_2747,N_2178,N_2418);
nand U2748 (N_2748,N_2267,N_2050);
nor U2749 (N_2749,N_2426,N_2029);
or U2750 (N_2750,N_2458,N_2445);
or U2751 (N_2751,N_2424,N_2015);
or U2752 (N_2752,N_2358,N_2469);
or U2753 (N_2753,N_2196,N_2456);
or U2754 (N_2754,N_2205,N_2232);
nand U2755 (N_2755,N_2054,N_2162);
nand U2756 (N_2756,N_2370,N_2136);
or U2757 (N_2757,N_2045,N_2174);
nand U2758 (N_2758,N_2232,N_2460);
nor U2759 (N_2759,N_2093,N_2292);
and U2760 (N_2760,N_2438,N_2462);
xnor U2761 (N_2761,N_2336,N_2087);
xnor U2762 (N_2762,N_2084,N_2152);
and U2763 (N_2763,N_2479,N_2357);
nand U2764 (N_2764,N_2391,N_2380);
and U2765 (N_2765,N_2225,N_2014);
and U2766 (N_2766,N_2242,N_2088);
or U2767 (N_2767,N_2085,N_2257);
nand U2768 (N_2768,N_2076,N_2302);
nand U2769 (N_2769,N_2360,N_2495);
or U2770 (N_2770,N_2008,N_2341);
nor U2771 (N_2771,N_2440,N_2149);
and U2772 (N_2772,N_2331,N_2085);
or U2773 (N_2773,N_2399,N_2192);
nand U2774 (N_2774,N_2119,N_2091);
or U2775 (N_2775,N_2195,N_2314);
nand U2776 (N_2776,N_2096,N_2260);
and U2777 (N_2777,N_2068,N_2032);
or U2778 (N_2778,N_2490,N_2107);
and U2779 (N_2779,N_2051,N_2227);
and U2780 (N_2780,N_2047,N_2441);
nor U2781 (N_2781,N_2024,N_2484);
and U2782 (N_2782,N_2345,N_2122);
or U2783 (N_2783,N_2212,N_2219);
or U2784 (N_2784,N_2230,N_2342);
nand U2785 (N_2785,N_2030,N_2360);
nand U2786 (N_2786,N_2338,N_2434);
xnor U2787 (N_2787,N_2087,N_2192);
and U2788 (N_2788,N_2344,N_2105);
or U2789 (N_2789,N_2099,N_2468);
nor U2790 (N_2790,N_2366,N_2106);
xor U2791 (N_2791,N_2103,N_2463);
and U2792 (N_2792,N_2433,N_2431);
xor U2793 (N_2793,N_2017,N_2435);
nor U2794 (N_2794,N_2260,N_2050);
or U2795 (N_2795,N_2075,N_2338);
nor U2796 (N_2796,N_2245,N_2193);
or U2797 (N_2797,N_2317,N_2292);
or U2798 (N_2798,N_2195,N_2413);
nor U2799 (N_2799,N_2374,N_2366);
nand U2800 (N_2800,N_2476,N_2026);
and U2801 (N_2801,N_2441,N_2167);
nand U2802 (N_2802,N_2269,N_2026);
or U2803 (N_2803,N_2169,N_2372);
nor U2804 (N_2804,N_2308,N_2429);
nor U2805 (N_2805,N_2377,N_2201);
xnor U2806 (N_2806,N_2295,N_2493);
or U2807 (N_2807,N_2151,N_2282);
nand U2808 (N_2808,N_2107,N_2293);
nand U2809 (N_2809,N_2132,N_2208);
and U2810 (N_2810,N_2082,N_2065);
nor U2811 (N_2811,N_2269,N_2445);
xor U2812 (N_2812,N_2144,N_2010);
or U2813 (N_2813,N_2137,N_2452);
or U2814 (N_2814,N_2293,N_2111);
nor U2815 (N_2815,N_2408,N_2162);
or U2816 (N_2816,N_2142,N_2441);
xnor U2817 (N_2817,N_2149,N_2105);
or U2818 (N_2818,N_2313,N_2319);
nand U2819 (N_2819,N_2290,N_2143);
and U2820 (N_2820,N_2407,N_2432);
xnor U2821 (N_2821,N_2049,N_2407);
xnor U2822 (N_2822,N_2390,N_2049);
or U2823 (N_2823,N_2062,N_2469);
xor U2824 (N_2824,N_2366,N_2019);
and U2825 (N_2825,N_2397,N_2386);
nand U2826 (N_2826,N_2112,N_2073);
and U2827 (N_2827,N_2335,N_2324);
or U2828 (N_2828,N_2186,N_2456);
nor U2829 (N_2829,N_2361,N_2076);
and U2830 (N_2830,N_2219,N_2262);
xnor U2831 (N_2831,N_2406,N_2010);
nand U2832 (N_2832,N_2272,N_2078);
nor U2833 (N_2833,N_2456,N_2361);
and U2834 (N_2834,N_2065,N_2049);
nor U2835 (N_2835,N_2009,N_2484);
nor U2836 (N_2836,N_2086,N_2054);
and U2837 (N_2837,N_2444,N_2151);
nor U2838 (N_2838,N_2355,N_2374);
xor U2839 (N_2839,N_2198,N_2069);
and U2840 (N_2840,N_2405,N_2388);
xor U2841 (N_2841,N_2293,N_2095);
nor U2842 (N_2842,N_2273,N_2373);
or U2843 (N_2843,N_2158,N_2256);
or U2844 (N_2844,N_2264,N_2224);
or U2845 (N_2845,N_2386,N_2454);
nor U2846 (N_2846,N_2108,N_2460);
and U2847 (N_2847,N_2346,N_2003);
and U2848 (N_2848,N_2351,N_2179);
nor U2849 (N_2849,N_2295,N_2260);
nor U2850 (N_2850,N_2005,N_2128);
or U2851 (N_2851,N_2487,N_2265);
nand U2852 (N_2852,N_2171,N_2448);
and U2853 (N_2853,N_2220,N_2266);
nand U2854 (N_2854,N_2206,N_2412);
or U2855 (N_2855,N_2078,N_2117);
and U2856 (N_2856,N_2344,N_2153);
or U2857 (N_2857,N_2162,N_2282);
nand U2858 (N_2858,N_2351,N_2493);
and U2859 (N_2859,N_2463,N_2201);
nor U2860 (N_2860,N_2215,N_2460);
or U2861 (N_2861,N_2224,N_2475);
or U2862 (N_2862,N_2254,N_2242);
and U2863 (N_2863,N_2451,N_2045);
nand U2864 (N_2864,N_2425,N_2444);
nor U2865 (N_2865,N_2351,N_2445);
or U2866 (N_2866,N_2262,N_2024);
nor U2867 (N_2867,N_2282,N_2120);
or U2868 (N_2868,N_2304,N_2094);
nand U2869 (N_2869,N_2262,N_2128);
nor U2870 (N_2870,N_2320,N_2481);
nor U2871 (N_2871,N_2333,N_2224);
nor U2872 (N_2872,N_2117,N_2256);
and U2873 (N_2873,N_2144,N_2374);
and U2874 (N_2874,N_2493,N_2314);
xnor U2875 (N_2875,N_2229,N_2286);
and U2876 (N_2876,N_2429,N_2215);
nand U2877 (N_2877,N_2267,N_2209);
and U2878 (N_2878,N_2183,N_2192);
and U2879 (N_2879,N_2015,N_2416);
nor U2880 (N_2880,N_2024,N_2315);
nor U2881 (N_2881,N_2004,N_2486);
nand U2882 (N_2882,N_2156,N_2191);
or U2883 (N_2883,N_2124,N_2057);
nand U2884 (N_2884,N_2479,N_2202);
nor U2885 (N_2885,N_2346,N_2259);
nor U2886 (N_2886,N_2376,N_2058);
or U2887 (N_2887,N_2462,N_2111);
nor U2888 (N_2888,N_2423,N_2047);
nand U2889 (N_2889,N_2005,N_2100);
nor U2890 (N_2890,N_2024,N_2346);
xor U2891 (N_2891,N_2497,N_2141);
and U2892 (N_2892,N_2215,N_2018);
nand U2893 (N_2893,N_2441,N_2402);
nand U2894 (N_2894,N_2142,N_2333);
xor U2895 (N_2895,N_2102,N_2381);
or U2896 (N_2896,N_2150,N_2412);
nand U2897 (N_2897,N_2348,N_2027);
and U2898 (N_2898,N_2086,N_2036);
xnor U2899 (N_2899,N_2100,N_2107);
or U2900 (N_2900,N_2184,N_2099);
xor U2901 (N_2901,N_2053,N_2359);
and U2902 (N_2902,N_2237,N_2287);
nand U2903 (N_2903,N_2070,N_2496);
and U2904 (N_2904,N_2142,N_2163);
or U2905 (N_2905,N_2408,N_2136);
nor U2906 (N_2906,N_2226,N_2451);
and U2907 (N_2907,N_2164,N_2220);
nand U2908 (N_2908,N_2412,N_2346);
or U2909 (N_2909,N_2332,N_2214);
nor U2910 (N_2910,N_2182,N_2061);
or U2911 (N_2911,N_2199,N_2414);
nand U2912 (N_2912,N_2315,N_2366);
nor U2913 (N_2913,N_2261,N_2361);
or U2914 (N_2914,N_2474,N_2164);
nor U2915 (N_2915,N_2282,N_2230);
or U2916 (N_2916,N_2044,N_2259);
and U2917 (N_2917,N_2369,N_2457);
or U2918 (N_2918,N_2117,N_2068);
nand U2919 (N_2919,N_2026,N_2489);
and U2920 (N_2920,N_2325,N_2322);
nand U2921 (N_2921,N_2450,N_2159);
nand U2922 (N_2922,N_2093,N_2065);
nor U2923 (N_2923,N_2220,N_2054);
and U2924 (N_2924,N_2281,N_2424);
or U2925 (N_2925,N_2235,N_2398);
and U2926 (N_2926,N_2010,N_2246);
or U2927 (N_2927,N_2254,N_2200);
nor U2928 (N_2928,N_2391,N_2140);
and U2929 (N_2929,N_2419,N_2480);
nor U2930 (N_2930,N_2299,N_2207);
xnor U2931 (N_2931,N_2194,N_2467);
or U2932 (N_2932,N_2277,N_2485);
nand U2933 (N_2933,N_2250,N_2025);
nand U2934 (N_2934,N_2262,N_2280);
xor U2935 (N_2935,N_2445,N_2175);
nor U2936 (N_2936,N_2320,N_2492);
or U2937 (N_2937,N_2486,N_2362);
or U2938 (N_2938,N_2058,N_2289);
nand U2939 (N_2939,N_2445,N_2171);
nand U2940 (N_2940,N_2198,N_2317);
nand U2941 (N_2941,N_2399,N_2163);
and U2942 (N_2942,N_2397,N_2322);
and U2943 (N_2943,N_2465,N_2331);
or U2944 (N_2944,N_2034,N_2239);
xnor U2945 (N_2945,N_2416,N_2135);
and U2946 (N_2946,N_2179,N_2334);
and U2947 (N_2947,N_2289,N_2020);
nand U2948 (N_2948,N_2231,N_2341);
nor U2949 (N_2949,N_2414,N_2480);
nor U2950 (N_2950,N_2444,N_2056);
or U2951 (N_2951,N_2077,N_2057);
and U2952 (N_2952,N_2282,N_2403);
nor U2953 (N_2953,N_2286,N_2275);
and U2954 (N_2954,N_2145,N_2259);
nor U2955 (N_2955,N_2107,N_2473);
nor U2956 (N_2956,N_2119,N_2024);
nor U2957 (N_2957,N_2056,N_2203);
or U2958 (N_2958,N_2324,N_2075);
nand U2959 (N_2959,N_2214,N_2386);
nand U2960 (N_2960,N_2039,N_2469);
or U2961 (N_2961,N_2112,N_2351);
xor U2962 (N_2962,N_2053,N_2456);
xor U2963 (N_2963,N_2122,N_2100);
nand U2964 (N_2964,N_2153,N_2450);
and U2965 (N_2965,N_2440,N_2391);
xnor U2966 (N_2966,N_2280,N_2064);
nand U2967 (N_2967,N_2233,N_2206);
nor U2968 (N_2968,N_2095,N_2276);
and U2969 (N_2969,N_2311,N_2327);
nand U2970 (N_2970,N_2492,N_2378);
nor U2971 (N_2971,N_2158,N_2037);
nor U2972 (N_2972,N_2496,N_2316);
nor U2973 (N_2973,N_2179,N_2094);
nor U2974 (N_2974,N_2471,N_2371);
nor U2975 (N_2975,N_2473,N_2165);
xnor U2976 (N_2976,N_2312,N_2002);
or U2977 (N_2977,N_2467,N_2419);
nor U2978 (N_2978,N_2033,N_2214);
nor U2979 (N_2979,N_2358,N_2422);
or U2980 (N_2980,N_2283,N_2253);
or U2981 (N_2981,N_2009,N_2329);
or U2982 (N_2982,N_2107,N_2182);
nor U2983 (N_2983,N_2117,N_2022);
xor U2984 (N_2984,N_2020,N_2431);
xnor U2985 (N_2985,N_2019,N_2275);
and U2986 (N_2986,N_2168,N_2399);
nand U2987 (N_2987,N_2430,N_2328);
nand U2988 (N_2988,N_2006,N_2211);
nor U2989 (N_2989,N_2220,N_2239);
or U2990 (N_2990,N_2245,N_2248);
or U2991 (N_2991,N_2228,N_2423);
or U2992 (N_2992,N_2430,N_2041);
nand U2993 (N_2993,N_2035,N_2218);
and U2994 (N_2994,N_2288,N_2259);
or U2995 (N_2995,N_2130,N_2188);
and U2996 (N_2996,N_2273,N_2202);
nor U2997 (N_2997,N_2033,N_2231);
or U2998 (N_2998,N_2464,N_2309);
or U2999 (N_2999,N_2488,N_2006);
and UO_0 (O_0,N_2961,N_2966);
nand UO_1 (O_1,N_2768,N_2586);
nor UO_2 (O_2,N_2678,N_2913);
nor UO_3 (O_3,N_2905,N_2700);
and UO_4 (O_4,N_2536,N_2967);
and UO_5 (O_5,N_2695,N_2657);
nand UO_6 (O_6,N_2790,N_2522);
or UO_7 (O_7,N_2526,N_2774);
nand UO_8 (O_8,N_2643,N_2892);
or UO_9 (O_9,N_2540,N_2562);
or UO_10 (O_10,N_2772,N_2754);
or UO_11 (O_11,N_2617,N_2706);
nand UO_12 (O_12,N_2635,N_2735);
nand UO_13 (O_13,N_2809,N_2982);
and UO_14 (O_14,N_2654,N_2650);
nand UO_15 (O_15,N_2680,N_2957);
nor UO_16 (O_16,N_2777,N_2642);
nor UO_17 (O_17,N_2721,N_2723);
nand UO_18 (O_18,N_2552,N_2510);
or UO_19 (O_19,N_2965,N_2683);
or UO_20 (O_20,N_2807,N_2704);
xor UO_21 (O_21,N_2501,N_2902);
nor UO_22 (O_22,N_2716,N_2715);
or UO_23 (O_23,N_2516,N_2749);
nor UO_24 (O_24,N_2925,N_2823);
and UO_25 (O_25,N_2887,N_2588);
xnor UO_26 (O_26,N_2949,N_2849);
and UO_27 (O_27,N_2585,N_2831);
or UO_28 (O_28,N_2856,N_2527);
or UO_29 (O_29,N_2659,N_2572);
nand UO_30 (O_30,N_2780,N_2545);
and UO_31 (O_31,N_2885,N_2820);
or UO_32 (O_32,N_2791,N_2514);
nor UO_33 (O_33,N_2784,N_2752);
nor UO_34 (O_34,N_2532,N_2983);
or UO_35 (O_35,N_2933,N_2800);
or UO_36 (O_36,N_2782,N_2857);
and UO_37 (O_37,N_2582,N_2688);
or UO_38 (O_38,N_2893,N_2558);
or UO_39 (O_39,N_2833,N_2661);
xnor UO_40 (O_40,N_2505,N_2684);
nand UO_41 (O_41,N_2665,N_2811);
or UO_42 (O_42,N_2616,N_2655);
or UO_43 (O_43,N_2679,N_2796);
nand UO_44 (O_44,N_2534,N_2845);
and UO_45 (O_45,N_2513,N_2675);
and UO_46 (O_46,N_2740,N_2955);
xor UO_47 (O_47,N_2681,N_2544);
and UO_48 (O_48,N_2568,N_2935);
nand UO_49 (O_49,N_2546,N_2810);
nor UO_50 (O_50,N_2741,N_2550);
or UO_51 (O_51,N_2578,N_2725);
or UO_52 (O_52,N_2995,N_2563);
or UO_53 (O_53,N_2824,N_2641);
nand UO_54 (O_54,N_2795,N_2753);
nor UO_55 (O_55,N_2794,N_2511);
nor UO_56 (O_56,N_2686,N_2828);
xnor UO_57 (O_57,N_2757,N_2970);
xor UO_58 (O_58,N_2822,N_2812);
nand UO_59 (O_59,N_2920,N_2668);
nor UO_60 (O_60,N_2669,N_2787);
nand UO_61 (O_61,N_2613,N_2537);
nor UO_62 (O_62,N_2636,N_2731);
nand UO_63 (O_63,N_2997,N_2980);
nor UO_64 (O_64,N_2692,N_2817);
and UO_65 (O_65,N_2660,N_2712);
and UO_66 (O_66,N_2512,N_2848);
or UO_67 (O_67,N_2797,N_2648);
or UO_68 (O_68,N_2687,N_2633);
or UO_69 (O_69,N_2717,N_2909);
or UO_70 (O_70,N_2879,N_2798);
nor UO_71 (O_71,N_2663,N_2576);
nor UO_72 (O_72,N_2917,N_2976);
and UO_73 (O_73,N_2506,N_2775);
and UO_74 (O_74,N_2803,N_2884);
or UO_75 (O_75,N_2509,N_2870);
nand UO_76 (O_76,N_2622,N_2555);
or UO_77 (O_77,N_2804,N_2869);
and UO_78 (O_78,N_2541,N_2951);
or UO_79 (O_79,N_2677,N_2921);
and UO_80 (O_80,N_2587,N_2747);
or UO_81 (O_81,N_2685,N_2785);
or UO_82 (O_82,N_2689,N_2763);
nor UO_83 (O_83,N_2714,N_2569);
xor UO_84 (O_84,N_2531,N_2947);
or UO_85 (O_85,N_2941,N_2639);
or UO_86 (O_86,N_2589,N_2606);
or UO_87 (O_87,N_2567,N_2600);
and UO_88 (O_88,N_2696,N_2652);
or UO_89 (O_89,N_2929,N_2878);
and UO_90 (O_90,N_2535,N_2829);
and UO_91 (O_91,N_2738,N_2500);
nor UO_92 (O_92,N_2503,N_2923);
and UO_93 (O_93,N_2533,N_2720);
and UO_94 (O_94,N_2530,N_2524);
and UO_95 (O_95,N_2838,N_2728);
and UO_96 (O_96,N_2894,N_2889);
xor UO_97 (O_97,N_2515,N_2814);
or UO_98 (O_98,N_2610,N_2727);
and UO_99 (O_99,N_2990,N_2998);
and UO_100 (O_100,N_2901,N_2750);
nor UO_101 (O_101,N_2904,N_2821);
and UO_102 (O_102,N_2919,N_2872);
nor UO_103 (O_103,N_2637,N_2960);
nand UO_104 (O_104,N_2840,N_2805);
or UO_105 (O_105,N_2888,N_2698);
nor UO_106 (O_106,N_2788,N_2786);
nor UO_107 (O_107,N_2553,N_2504);
and UO_108 (O_108,N_2881,N_2547);
and UO_109 (O_109,N_2602,N_2592);
and UO_110 (O_110,N_2579,N_2624);
nand UO_111 (O_111,N_2584,N_2525);
nand UO_112 (O_112,N_2575,N_2979);
or UO_113 (O_113,N_2882,N_2508);
or UO_114 (O_114,N_2528,N_2649);
nand UO_115 (O_115,N_2758,N_2710);
or UO_116 (O_116,N_2851,N_2626);
and UO_117 (O_117,N_2808,N_2937);
nand UO_118 (O_118,N_2959,N_2762);
xor UO_119 (O_119,N_2718,N_2865);
or UO_120 (O_120,N_2815,N_2631);
nor UO_121 (O_121,N_2672,N_2694);
and UO_122 (O_122,N_2673,N_2682);
nand UO_123 (O_123,N_2928,N_2945);
and UO_124 (O_124,N_2936,N_2978);
xor UO_125 (O_125,N_2908,N_2598);
nand UO_126 (O_126,N_2618,N_2597);
nor UO_127 (O_127,N_2953,N_2975);
nand UO_128 (O_128,N_2732,N_2644);
xor UO_129 (O_129,N_2972,N_2765);
and UO_130 (O_130,N_2591,N_2866);
nor UO_131 (O_131,N_2994,N_2981);
and UO_132 (O_132,N_2609,N_2926);
and UO_133 (O_133,N_2615,N_2867);
and UO_134 (O_134,N_2852,N_2806);
and UO_135 (O_135,N_2746,N_2903);
or UO_136 (O_136,N_2854,N_2583);
and UO_137 (O_137,N_2577,N_2939);
nand UO_138 (O_138,N_2934,N_2580);
or UO_139 (O_139,N_2880,N_2656);
or UO_140 (O_140,N_2628,N_2724);
or UO_141 (O_141,N_2897,N_2991);
and UO_142 (O_142,N_2907,N_2899);
or UO_143 (O_143,N_2662,N_2719);
or UO_144 (O_144,N_2799,N_2973);
nand UO_145 (O_145,N_2502,N_2566);
nor UO_146 (O_146,N_2858,N_2915);
and UO_147 (O_147,N_2962,N_2846);
or UO_148 (O_148,N_2911,N_2847);
nand UO_149 (O_149,N_2940,N_2733);
and UO_150 (O_150,N_2601,N_2938);
nor UO_151 (O_151,N_2574,N_2573);
nor UO_152 (O_152,N_2596,N_2590);
nor UO_153 (O_153,N_2507,N_2607);
and UO_154 (O_154,N_2664,N_2756);
nor UO_155 (O_155,N_2709,N_2956);
or UO_156 (O_156,N_2958,N_2581);
and UO_157 (O_157,N_2968,N_2638);
or UO_158 (O_158,N_2760,N_2729);
nor UO_159 (O_159,N_2627,N_2634);
nand UO_160 (O_160,N_2910,N_2674);
or UO_161 (O_161,N_2755,N_2873);
nor UO_162 (O_162,N_2860,N_2691);
nand UO_163 (O_163,N_2819,N_2924);
nor UO_164 (O_164,N_2651,N_2801);
and UO_165 (O_165,N_2942,N_2877);
nand UO_166 (O_166,N_2843,N_2842);
xor UO_167 (O_167,N_2766,N_2548);
and UO_168 (O_168,N_2789,N_2999);
or UO_169 (O_169,N_2918,N_2671);
nand UO_170 (O_170,N_2861,N_2538);
or UO_171 (O_171,N_2818,N_2561);
nor UO_172 (O_172,N_2625,N_2930);
or UO_173 (O_173,N_2977,N_2726);
or UO_174 (O_174,N_2542,N_2705);
nand UO_175 (O_175,N_2521,N_2783);
nor UO_176 (O_176,N_2543,N_2871);
nand UO_177 (O_177,N_2701,N_2987);
and UO_178 (O_178,N_2612,N_2946);
nand UO_179 (O_179,N_2868,N_2557);
nand UO_180 (O_180,N_2640,N_2539);
nand UO_181 (O_181,N_2771,N_2736);
nand UO_182 (O_182,N_2781,N_2974);
nand UO_183 (O_183,N_2839,N_2922);
and UO_184 (O_184,N_2813,N_2985);
and UO_185 (O_185,N_2841,N_2703);
or UO_186 (O_186,N_2739,N_2850);
nor UO_187 (O_187,N_2876,N_2912);
or UO_188 (O_188,N_2702,N_2520);
and UO_189 (O_189,N_2517,N_2699);
or UO_190 (O_190,N_2707,N_2943);
nor UO_191 (O_191,N_2556,N_2730);
nand UO_192 (O_192,N_2874,N_2834);
nand UO_193 (O_193,N_2611,N_2944);
or UO_194 (O_194,N_2864,N_2751);
and UO_195 (O_195,N_2855,N_2599);
or UO_196 (O_196,N_2594,N_2896);
or UO_197 (O_197,N_2963,N_2551);
and UO_198 (O_198,N_2554,N_2620);
nand UO_199 (O_199,N_2745,N_2996);
and UO_200 (O_200,N_2950,N_2883);
or UO_201 (O_201,N_2969,N_2708);
or UO_202 (O_202,N_2778,N_2621);
and UO_203 (O_203,N_2776,N_2875);
and UO_204 (O_204,N_2825,N_2886);
and UO_205 (O_205,N_2529,N_2632);
or UO_206 (O_206,N_2564,N_2916);
nand UO_207 (O_207,N_2802,N_2853);
and UO_208 (O_208,N_2742,N_2827);
or UO_209 (O_209,N_2769,N_2779);
or UO_210 (O_210,N_2630,N_2549);
nand UO_211 (O_211,N_2859,N_2666);
nor UO_212 (O_212,N_2619,N_2743);
and UO_213 (O_213,N_2900,N_2890);
and UO_214 (O_214,N_2898,N_2676);
and UO_215 (O_215,N_2773,N_2931);
xnor UO_216 (O_216,N_2914,N_2646);
or UO_217 (O_217,N_2988,N_2993);
or UO_218 (O_218,N_2984,N_2570);
nor UO_219 (O_219,N_2614,N_2986);
and UO_220 (O_220,N_2604,N_2830);
nor UO_221 (O_221,N_2734,N_2971);
or UO_222 (O_222,N_2748,N_2895);
nor UO_223 (O_223,N_2792,N_2759);
and UO_224 (O_224,N_2645,N_2711);
or UO_225 (O_225,N_2826,N_2793);
and UO_226 (O_226,N_2523,N_2658);
and UO_227 (O_227,N_2836,N_2737);
and UO_228 (O_228,N_2767,N_2608);
nor UO_229 (O_229,N_2605,N_2770);
and UO_230 (O_230,N_2837,N_2518);
xnor UO_231 (O_231,N_2690,N_2629);
nand UO_232 (O_232,N_2519,N_2565);
or UO_233 (O_233,N_2670,N_2948);
nor UO_234 (O_234,N_2693,N_2764);
nor UO_235 (O_235,N_2647,N_2571);
or UO_236 (O_236,N_2816,N_2832);
xor UO_237 (O_237,N_2992,N_2560);
xor UO_238 (O_238,N_2744,N_2623);
and UO_239 (O_239,N_2862,N_2593);
xnor UO_240 (O_240,N_2954,N_2595);
xnor UO_241 (O_241,N_2761,N_2989);
nand UO_242 (O_242,N_2863,N_2952);
nor UO_243 (O_243,N_2697,N_2653);
nand UO_244 (O_244,N_2667,N_2559);
nand UO_245 (O_245,N_2835,N_2932);
nor UO_246 (O_246,N_2603,N_2713);
nand UO_247 (O_247,N_2906,N_2844);
nand UO_248 (O_248,N_2927,N_2891);
and UO_249 (O_249,N_2964,N_2722);
and UO_250 (O_250,N_2721,N_2607);
nand UO_251 (O_251,N_2764,N_2949);
nor UO_252 (O_252,N_2525,N_2953);
nor UO_253 (O_253,N_2514,N_2806);
and UO_254 (O_254,N_2798,N_2704);
nand UO_255 (O_255,N_2833,N_2521);
and UO_256 (O_256,N_2589,N_2930);
nor UO_257 (O_257,N_2802,N_2765);
or UO_258 (O_258,N_2883,N_2901);
and UO_259 (O_259,N_2519,N_2683);
nand UO_260 (O_260,N_2888,N_2606);
or UO_261 (O_261,N_2507,N_2681);
nand UO_262 (O_262,N_2925,N_2855);
and UO_263 (O_263,N_2839,N_2729);
nand UO_264 (O_264,N_2669,N_2979);
or UO_265 (O_265,N_2555,N_2999);
nand UO_266 (O_266,N_2642,N_2846);
and UO_267 (O_267,N_2627,N_2767);
or UO_268 (O_268,N_2579,N_2963);
nand UO_269 (O_269,N_2865,N_2795);
or UO_270 (O_270,N_2819,N_2641);
nand UO_271 (O_271,N_2792,N_2725);
and UO_272 (O_272,N_2771,N_2764);
nand UO_273 (O_273,N_2888,N_2986);
nand UO_274 (O_274,N_2580,N_2877);
or UO_275 (O_275,N_2612,N_2636);
nand UO_276 (O_276,N_2674,N_2517);
or UO_277 (O_277,N_2887,N_2767);
nor UO_278 (O_278,N_2684,N_2988);
or UO_279 (O_279,N_2980,N_2831);
or UO_280 (O_280,N_2921,N_2538);
and UO_281 (O_281,N_2503,N_2792);
xnor UO_282 (O_282,N_2830,N_2665);
nor UO_283 (O_283,N_2935,N_2542);
nor UO_284 (O_284,N_2836,N_2544);
nand UO_285 (O_285,N_2748,N_2691);
nor UO_286 (O_286,N_2693,N_2901);
xnor UO_287 (O_287,N_2827,N_2937);
xnor UO_288 (O_288,N_2764,N_2740);
or UO_289 (O_289,N_2774,N_2612);
nand UO_290 (O_290,N_2683,N_2983);
and UO_291 (O_291,N_2704,N_2624);
and UO_292 (O_292,N_2586,N_2600);
and UO_293 (O_293,N_2912,N_2654);
or UO_294 (O_294,N_2833,N_2648);
or UO_295 (O_295,N_2929,N_2962);
nor UO_296 (O_296,N_2522,N_2963);
and UO_297 (O_297,N_2703,N_2688);
nor UO_298 (O_298,N_2626,N_2655);
and UO_299 (O_299,N_2751,N_2998);
nand UO_300 (O_300,N_2781,N_2654);
xnor UO_301 (O_301,N_2623,N_2697);
nor UO_302 (O_302,N_2532,N_2562);
nor UO_303 (O_303,N_2600,N_2565);
xnor UO_304 (O_304,N_2900,N_2822);
and UO_305 (O_305,N_2707,N_2800);
nand UO_306 (O_306,N_2730,N_2654);
nor UO_307 (O_307,N_2847,N_2549);
nor UO_308 (O_308,N_2913,N_2922);
and UO_309 (O_309,N_2658,N_2559);
or UO_310 (O_310,N_2701,N_2813);
nor UO_311 (O_311,N_2875,N_2541);
nand UO_312 (O_312,N_2777,N_2963);
or UO_313 (O_313,N_2760,N_2995);
or UO_314 (O_314,N_2538,N_2550);
or UO_315 (O_315,N_2724,N_2846);
and UO_316 (O_316,N_2810,N_2764);
nor UO_317 (O_317,N_2588,N_2869);
nand UO_318 (O_318,N_2912,N_2847);
nor UO_319 (O_319,N_2950,N_2715);
and UO_320 (O_320,N_2788,N_2853);
nor UO_321 (O_321,N_2854,N_2710);
nand UO_322 (O_322,N_2858,N_2965);
and UO_323 (O_323,N_2852,N_2543);
and UO_324 (O_324,N_2819,N_2642);
and UO_325 (O_325,N_2526,N_2763);
or UO_326 (O_326,N_2759,N_2748);
or UO_327 (O_327,N_2811,N_2956);
and UO_328 (O_328,N_2829,N_2640);
nand UO_329 (O_329,N_2556,N_2972);
xnor UO_330 (O_330,N_2577,N_2831);
and UO_331 (O_331,N_2652,N_2945);
nand UO_332 (O_332,N_2711,N_2791);
nand UO_333 (O_333,N_2770,N_2544);
nand UO_334 (O_334,N_2614,N_2679);
nor UO_335 (O_335,N_2940,N_2707);
nor UO_336 (O_336,N_2611,N_2756);
or UO_337 (O_337,N_2551,N_2678);
or UO_338 (O_338,N_2962,N_2692);
nor UO_339 (O_339,N_2940,N_2939);
or UO_340 (O_340,N_2597,N_2742);
and UO_341 (O_341,N_2940,N_2937);
or UO_342 (O_342,N_2619,N_2501);
nor UO_343 (O_343,N_2743,N_2508);
and UO_344 (O_344,N_2530,N_2982);
and UO_345 (O_345,N_2625,N_2786);
or UO_346 (O_346,N_2574,N_2834);
or UO_347 (O_347,N_2929,N_2576);
nand UO_348 (O_348,N_2866,N_2693);
xnor UO_349 (O_349,N_2905,N_2625);
xor UO_350 (O_350,N_2651,N_2697);
nand UO_351 (O_351,N_2512,N_2510);
and UO_352 (O_352,N_2691,N_2839);
or UO_353 (O_353,N_2823,N_2596);
nand UO_354 (O_354,N_2530,N_2784);
and UO_355 (O_355,N_2572,N_2749);
nor UO_356 (O_356,N_2535,N_2817);
or UO_357 (O_357,N_2846,N_2701);
nor UO_358 (O_358,N_2872,N_2505);
or UO_359 (O_359,N_2731,N_2807);
or UO_360 (O_360,N_2637,N_2626);
or UO_361 (O_361,N_2874,N_2501);
xnor UO_362 (O_362,N_2622,N_2867);
nand UO_363 (O_363,N_2752,N_2626);
or UO_364 (O_364,N_2947,N_2975);
nor UO_365 (O_365,N_2843,N_2536);
or UO_366 (O_366,N_2838,N_2659);
nand UO_367 (O_367,N_2598,N_2566);
nor UO_368 (O_368,N_2562,N_2684);
xnor UO_369 (O_369,N_2718,N_2517);
and UO_370 (O_370,N_2764,N_2842);
nand UO_371 (O_371,N_2790,N_2989);
nand UO_372 (O_372,N_2587,N_2636);
xnor UO_373 (O_373,N_2595,N_2809);
and UO_374 (O_374,N_2767,N_2749);
and UO_375 (O_375,N_2769,N_2721);
and UO_376 (O_376,N_2969,N_2938);
and UO_377 (O_377,N_2673,N_2557);
nand UO_378 (O_378,N_2746,N_2561);
nor UO_379 (O_379,N_2726,N_2734);
and UO_380 (O_380,N_2668,N_2809);
nand UO_381 (O_381,N_2966,N_2905);
nand UO_382 (O_382,N_2977,N_2576);
or UO_383 (O_383,N_2679,N_2800);
nand UO_384 (O_384,N_2746,N_2959);
nand UO_385 (O_385,N_2695,N_2830);
nor UO_386 (O_386,N_2597,N_2541);
or UO_387 (O_387,N_2941,N_2758);
nor UO_388 (O_388,N_2642,N_2813);
xor UO_389 (O_389,N_2926,N_2961);
xnor UO_390 (O_390,N_2556,N_2565);
and UO_391 (O_391,N_2860,N_2598);
nor UO_392 (O_392,N_2793,N_2524);
or UO_393 (O_393,N_2526,N_2585);
and UO_394 (O_394,N_2823,N_2637);
or UO_395 (O_395,N_2978,N_2513);
nand UO_396 (O_396,N_2942,N_2688);
nor UO_397 (O_397,N_2972,N_2878);
nand UO_398 (O_398,N_2504,N_2832);
and UO_399 (O_399,N_2699,N_2522);
or UO_400 (O_400,N_2746,N_2853);
or UO_401 (O_401,N_2800,N_2859);
nand UO_402 (O_402,N_2571,N_2645);
or UO_403 (O_403,N_2802,N_2916);
nor UO_404 (O_404,N_2577,N_2850);
nand UO_405 (O_405,N_2832,N_2935);
and UO_406 (O_406,N_2883,N_2843);
and UO_407 (O_407,N_2699,N_2846);
and UO_408 (O_408,N_2756,N_2678);
nand UO_409 (O_409,N_2753,N_2912);
xor UO_410 (O_410,N_2578,N_2842);
or UO_411 (O_411,N_2655,N_2959);
nor UO_412 (O_412,N_2509,N_2546);
nor UO_413 (O_413,N_2536,N_2834);
or UO_414 (O_414,N_2741,N_2952);
nand UO_415 (O_415,N_2732,N_2819);
and UO_416 (O_416,N_2803,N_2518);
or UO_417 (O_417,N_2676,N_2760);
and UO_418 (O_418,N_2757,N_2529);
or UO_419 (O_419,N_2571,N_2673);
nand UO_420 (O_420,N_2679,N_2764);
nor UO_421 (O_421,N_2805,N_2864);
xnor UO_422 (O_422,N_2739,N_2909);
and UO_423 (O_423,N_2707,N_2860);
or UO_424 (O_424,N_2809,N_2939);
nor UO_425 (O_425,N_2870,N_2600);
xnor UO_426 (O_426,N_2563,N_2702);
nor UO_427 (O_427,N_2548,N_2738);
nand UO_428 (O_428,N_2637,N_2604);
or UO_429 (O_429,N_2561,N_2581);
and UO_430 (O_430,N_2592,N_2557);
xnor UO_431 (O_431,N_2945,N_2562);
xnor UO_432 (O_432,N_2513,N_2896);
and UO_433 (O_433,N_2798,N_2977);
nor UO_434 (O_434,N_2579,N_2953);
nand UO_435 (O_435,N_2802,N_2933);
or UO_436 (O_436,N_2843,N_2811);
or UO_437 (O_437,N_2745,N_2598);
or UO_438 (O_438,N_2762,N_2792);
xnor UO_439 (O_439,N_2864,N_2741);
or UO_440 (O_440,N_2828,N_2953);
nand UO_441 (O_441,N_2831,N_2778);
or UO_442 (O_442,N_2961,N_2870);
or UO_443 (O_443,N_2544,N_2917);
nand UO_444 (O_444,N_2835,N_2839);
and UO_445 (O_445,N_2587,N_2921);
nand UO_446 (O_446,N_2717,N_2639);
nand UO_447 (O_447,N_2938,N_2581);
and UO_448 (O_448,N_2624,N_2611);
xnor UO_449 (O_449,N_2613,N_2881);
nor UO_450 (O_450,N_2866,N_2521);
xor UO_451 (O_451,N_2728,N_2848);
nor UO_452 (O_452,N_2858,N_2626);
xor UO_453 (O_453,N_2733,N_2894);
xor UO_454 (O_454,N_2574,N_2956);
nand UO_455 (O_455,N_2580,N_2762);
nand UO_456 (O_456,N_2905,N_2977);
and UO_457 (O_457,N_2654,N_2820);
or UO_458 (O_458,N_2811,N_2868);
and UO_459 (O_459,N_2686,N_2619);
nor UO_460 (O_460,N_2837,N_2911);
nand UO_461 (O_461,N_2788,N_2934);
or UO_462 (O_462,N_2500,N_2910);
and UO_463 (O_463,N_2601,N_2551);
nor UO_464 (O_464,N_2533,N_2785);
and UO_465 (O_465,N_2585,N_2798);
nor UO_466 (O_466,N_2995,N_2650);
xor UO_467 (O_467,N_2639,N_2945);
xnor UO_468 (O_468,N_2806,N_2951);
or UO_469 (O_469,N_2578,N_2968);
xnor UO_470 (O_470,N_2808,N_2972);
and UO_471 (O_471,N_2950,N_2994);
nor UO_472 (O_472,N_2650,N_2809);
or UO_473 (O_473,N_2995,N_2805);
nor UO_474 (O_474,N_2537,N_2784);
nand UO_475 (O_475,N_2649,N_2668);
and UO_476 (O_476,N_2897,N_2533);
nor UO_477 (O_477,N_2514,N_2601);
nand UO_478 (O_478,N_2949,N_2752);
and UO_479 (O_479,N_2911,N_2917);
nor UO_480 (O_480,N_2652,N_2769);
nand UO_481 (O_481,N_2558,N_2738);
nand UO_482 (O_482,N_2717,N_2967);
and UO_483 (O_483,N_2576,N_2603);
nor UO_484 (O_484,N_2568,N_2608);
or UO_485 (O_485,N_2826,N_2729);
nor UO_486 (O_486,N_2549,N_2898);
nand UO_487 (O_487,N_2513,N_2751);
nor UO_488 (O_488,N_2672,N_2624);
and UO_489 (O_489,N_2928,N_2645);
nand UO_490 (O_490,N_2668,N_2695);
or UO_491 (O_491,N_2608,N_2725);
or UO_492 (O_492,N_2941,N_2669);
or UO_493 (O_493,N_2636,N_2589);
or UO_494 (O_494,N_2554,N_2799);
nand UO_495 (O_495,N_2637,N_2994);
nor UO_496 (O_496,N_2538,N_2553);
and UO_497 (O_497,N_2655,N_2628);
xor UO_498 (O_498,N_2660,N_2918);
nand UO_499 (O_499,N_2506,N_2871);
endmodule