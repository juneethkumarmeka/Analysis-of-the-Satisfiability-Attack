module basic_500_3000_500_4_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_124,In_285);
or U1 (N_1,In_304,In_419);
nand U2 (N_2,In_230,In_108);
nor U3 (N_3,In_421,In_121);
nor U4 (N_4,In_312,In_307);
or U5 (N_5,In_449,In_387);
nand U6 (N_6,In_8,In_223);
and U7 (N_7,In_136,In_401);
nor U8 (N_8,In_212,In_250);
or U9 (N_9,In_26,In_226);
nor U10 (N_10,In_478,In_98);
nand U11 (N_11,In_468,In_93);
xnor U12 (N_12,In_350,In_262);
nor U13 (N_13,In_110,In_62);
or U14 (N_14,In_282,In_374);
nand U15 (N_15,In_201,In_426);
nor U16 (N_16,In_126,In_288);
and U17 (N_17,In_247,In_259);
nand U18 (N_18,In_5,In_398);
and U19 (N_19,In_209,In_111);
and U20 (N_20,In_393,In_443);
and U21 (N_21,In_415,In_327);
nand U22 (N_22,In_35,In_21);
nand U23 (N_23,In_138,In_188);
nand U24 (N_24,In_204,In_129);
and U25 (N_25,In_391,In_127);
and U26 (N_26,In_73,In_324);
xnor U27 (N_27,In_107,In_376);
nand U28 (N_28,In_182,In_9);
nor U29 (N_29,In_221,In_337);
nand U30 (N_30,In_116,In_220);
nor U31 (N_31,In_491,In_89);
or U32 (N_32,In_195,In_271);
or U33 (N_33,In_79,In_329);
and U34 (N_34,In_57,In_397);
and U35 (N_35,In_444,In_433);
nor U36 (N_36,In_144,In_119);
nor U37 (N_37,In_135,In_280);
or U38 (N_38,In_276,In_248);
nor U39 (N_39,In_395,In_261);
nor U40 (N_40,In_298,In_345);
or U41 (N_41,In_6,In_46);
nor U42 (N_42,In_94,In_355);
nand U43 (N_43,In_75,In_464);
and U44 (N_44,In_161,In_428);
or U45 (N_45,In_211,In_180);
and U46 (N_46,In_186,In_80);
and U47 (N_47,In_302,In_403);
or U48 (N_48,In_323,In_319);
and U49 (N_49,In_30,In_370);
nor U50 (N_50,In_495,In_326);
and U51 (N_51,In_18,In_382);
or U52 (N_52,In_103,In_364);
nand U53 (N_53,In_390,In_325);
or U54 (N_54,In_76,In_236);
or U55 (N_55,In_11,In_109);
and U56 (N_56,In_294,In_424);
or U57 (N_57,In_333,In_342);
and U58 (N_58,In_163,In_214);
nor U59 (N_59,In_493,In_205);
and U60 (N_60,In_192,In_358);
nor U61 (N_61,In_361,In_470);
and U62 (N_62,In_490,In_232);
or U63 (N_63,In_77,In_318);
and U64 (N_64,In_199,In_392);
nor U65 (N_65,In_438,In_412);
nor U66 (N_66,In_279,In_19);
and U67 (N_67,In_469,In_472);
or U68 (N_68,In_281,In_152);
or U69 (N_69,In_17,In_141);
and U70 (N_70,In_362,In_134);
and U71 (N_71,In_331,In_215);
nand U72 (N_72,In_191,In_287);
nand U73 (N_73,In_71,In_356);
nand U74 (N_74,In_12,In_32);
or U75 (N_75,In_239,In_434);
or U76 (N_76,In_123,In_224);
nor U77 (N_77,In_146,In_15);
and U78 (N_78,In_269,In_448);
or U79 (N_79,In_70,In_310);
nor U80 (N_80,In_100,In_359);
nor U81 (N_81,In_145,In_335);
or U82 (N_82,In_386,In_499);
nand U83 (N_83,In_4,In_187);
or U84 (N_84,In_227,In_260);
and U85 (N_85,In_128,In_407);
or U86 (N_86,In_456,In_427);
nand U87 (N_87,In_213,In_117);
and U88 (N_88,In_167,In_194);
or U89 (N_89,In_413,In_66);
nand U90 (N_90,In_441,In_10);
and U91 (N_91,In_408,In_241);
and U92 (N_92,In_475,In_455);
nand U93 (N_93,In_237,In_436);
and U94 (N_94,In_314,In_473);
and U95 (N_95,In_90,In_59);
nand U96 (N_96,In_341,In_176);
and U97 (N_97,In_466,In_137);
and U98 (N_98,In_91,In_133);
nor U99 (N_99,In_0,In_25);
or U100 (N_100,In_185,In_297);
or U101 (N_101,In_1,In_458);
and U102 (N_102,In_439,In_430);
nor U103 (N_103,In_340,In_104);
and U104 (N_104,In_131,In_388);
and U105 (N_105,In_33,In_38);
nand U106 (N_106,In_368,In_140);
nand U107 (N_107,In_229,In_166);
nand U108 (N_108,In_164,In_306);
or U109 (N_109,In_159,In_139);
nor U110 (N_110,In_252,In_384);
nand U111 (N_111,In_292,In_172);
or U112 (N_112,In_153,In_348);
nor U113 (N_113,In_251,In_485);
nor U114 (N_114,In_151,In_277);
nor U115 (N_115,In_385,In_206);
xor U116 (N_116,In_488,In_483);
nor U117 (N_117,In_184,In_267);
and U118 (N_118,In_474,In_243);
nor U119 (N_119,In_50,In_183);
nor U120 (N_120,In_411,In_169);
nor U121 (N_121,In_437,In_346);
nand U122 (N_122,In_190,In_425);
and U123 (N_123,In_132,In_486);
and U124 (N_124,In_492,In_344);
or U125 (N_125,In_270,In_489);
and U126 (N_126,In_465,In_263);
nor U127 (N_127,In_414,In_200);
or U128 (N_128,In_45,In_467);
nand U129 (N_129,In_208,In_7);
or U130 (N_130,In_290,In_300);
nor U131 (N_131,In_375,In_189);
and U132 (N_132,In_41,In_404);
or U133 (N_133,In_431,In_60);
or U134 (N_134,In_115,In_257);
or U135 (N_135,In_351,In_394);
nand U136 (N_136,In_160,In_148);
nor U137 (N_137,In_278,In_339);
and U138 (N_138,In_330,In_150);
and U139 (N_139,In_245,In_13);
or U140 (N_140,In_23,In_367);
and U141 (N_141,In_258,In_410);
nor U142 (N_142,In_156,In_101);
nor U143 (N_143,In_378,In_497);
or U144 (N_144,In_55,In_445);
or U145 (N_145,In_99,In_380);
and U146 (N_146,In_36,In_389);
nand U147 (N_147,In_225,In_354);
nand U148 (N_148,In_246,In_87);
nand U149 (N_149,In_78,In_154);
or U150 (N_150,In_363,In_82);
nor U151 (N_151,In_228,In_296);
nand U152 (N_152,In_171,In_496);
nor U153 (N_153,In_112,In_357);
or U154 (N_154,In_202,In_429);
nor U155 (N_155,In_400,In_471);
nand U156 (N_156,In_175,In_63);
or U157 (N_157,In_396,In_446);
or U158 (N_158,In_453,In_210);
nand U159 (N_159,In_315,In_238);
or U160 (N_160,In_106,In_22);
and U161 (N_161,In_84,In_72);
nand U162 (N_162,In_417,In_24);
nor U163 (N_163,In_274,In_264);
or U164 (N_164,In_487,In_273);
and U165 (N_165,In_40,In_416);
nand U166 (N_166,In_321,In_39);
nor U167 (N_167,In_313,In_147);
nor U168 (N_168,In_83,In_61);
nand U169 (N_169,In_463,In_371);
nand U170 (N_170,In_435,In_69);
nand U171 (N_171,In_197,In_97);
and U172 (N_172,In_405,In_420);
nand U173 (N_173,In_20,In_343);
or U174 (N_174,In_402,In_462);
or U175 (N_175,In_219,In_74);
nor U176 (N_176,In_56,In_34);
or U177 (N_177,In_142,In_143);
nor U178 (N_178,In_299,In_253);
and U179 (N_179,In_31,In_322);
or U180 (N_180,In_193,In_303);
nor U181 (N_181,In_440,In_311);
and U182 (N_182,In_48,In_162);
nor U183 (N_183,In_480,In_203);
or U184 (N_184,In_432,In_461);
or U185 (N_185,In_242,In_320);
nor U186 (N_186,In_452,In_317);
or U187 (N_187,In_482,In_338);
or U188 (N_188,In_157,In_173);
and U189 (N_189,In_353,In_29);
nand U190 (N_190,In_265,In_293);
nand U191 (N_191,In_377,In_118);
and U192 (N_192,In_178,In_81);
or U193 (N_193,In_181,In_308);
and U194 (N_194,In_179,In_301);
nand U195 (N_195,In_328,In_222);
nor U196 (N_196,In_409,In_96);
and U197 (N_197,In_177,In_305);
or U198 (N_198,In_256,In_360);
nand U199 (N_199,In_28,In_447);
and U200 (N_200,In_334,In_379);
or U201 (N_201,In_347,In_43);
nand U202 (N_202,In_120,In_494);
nand U203 (N_203,In_381,In_442);
nand U204 (N_204,In_336,In_130);
or U205 (N_205,In_174,In_459);
and U206 (N_206,In_406,In_2);
and U207 (N_207,In_383,In_240);
and U208 (N_208,In_102,In_309);
or U209 (N_209,In_479,In_451);
or U210 (N_210,In_234,In_113);
nand U211 (N_211,In_255,In_3);
nor U212 (N_212,In_86,In_231);
nand U213 (N_213,In_168,In_457);
or U214 (N_214,In_332,In_54);
and U215 (N_215,In_122,In_399);
nor U216 (N_216,In_460,In_42);
and U217 (N_217,In_47,In_27);
nor U218 (N_218,In_58,In_316);
nand U219 (N_219,In_423,In_372);
nor U220 (N_220,In_295,In_95);
nand U221 (N_221,In_198,In_291);
or U222 (N_222,In_286,In_272);
and U223 (N_223,In_149,In_125);
or U224 (N_224,In_289,In_484);
nor U225 (N_225,In_477,In_268);
nor U226 (N_226,In_67,In_266);
or U227 (N_227,In_373,In_352);
nor U228 (N_228,In_450,In_283);
or U229 (N_229,In_52,In_158);
or U230 (N_230,In_14,In_498);
nor U231 (N_231,In_65,In_114);
or U232 (N_232,In_218,In_476);
or U233 (N_233,In_349,In_244);
and U234 (N_234,In_249,In_64);
and U235 (N_235,In_254,In_37);
nor U236 (N_236,In_235,In_454);
and U237 (N_237,In_68,In_49);
nor U238 (N_238,In_207,In_105);
nand U239 (N_239,In_16,In_92);
nand U240 (N_240,In_233,In_366);
nand U241 (N_241,In_422,In_217);
and U242 (N_242,In_216,In_165);
and U243 (N_243,In_155,In_85);
or U244 (N_244,In_369,In_88);
or U245 (N_245,In_284,In_44);
nor U246 (N_246,In_365,In_418);
or U247 (N_247,In_196,In_481);
nand U248 (N_248,In_170,In_53);
or U249 (N_249,In_275,In_51);
nand U250 (N_250,In_155,In_189);
nor U251 (N_251,In_304,In_167);
nand U252 (N_252,In_134,In_324);
nor U253 (N_253,In_16,In_290);
and U254 (N_254,In_323,In_97);
and U255 (N_255,In_444,In_313);
and U256 (N_256,In_43,In_209);
nand U257 (N_257,In_144,In_45);
nor U258 (N_258,In_312,In_443);
and U259 (N_259,In_118,In_158);
nand U260 (N_260,In_127,In_197);
nor U261 (N_261,In_348,In_439);
nand U262 (N_262,In_428,In_396);
nand U263 (N_263,In_209,In_131);
or U264 (N_264,In_380,In_486);
nand U265 (N_265,In_99,In_214);
and U266 (N_266,In_105,In_190);
and U267 (N_267,In_73,In_171);
nand U268 (N_268,In_11,In_8);
nand U269 (N_269,In_77,In_414);
and U270 (N_270,In_10,In_54);
or U271 (N_271,In_98,In_433);
nand U272 (N_272,In_72,In_198);
or U273 (N_273,In_487,In_457);
nor U274 (N_274,In_14,In_267);
and U275 (N_275,In_236,In_158);
and U276 (N_276,In_265,In_372);
or U277 (N_277,In_243,In_156);
and U278 (N_278,In_323,In_166);
nor U279 (N_279,In_38,In_470);
nand U280 (N_280,In_237,In_7);
or U281 (N_281,In_277,In_446);
nand U282 (N_282,In_359,In_115);
or U283 (N_283,In_440,In_461);
or U284 (N_284,In_385,In_454);
nor U285 (N_285,In_405,In_72);
nand U286 (N_286,In_304,In_456);
nand U287 (N_287,In_84,In_365);
and U288 (N_288,In_289,In_320);
nand U289 (N_289,In_153,In_220);
nand U290 (N_290,In_91,In_495);
and U291 (N_291,In_254,In_393);
nor U292 (N_292,In_106,In_91);
or U293 (N_293,In_311,In_468);
nand U294 (N_294,In_346,In_66);
nor U295 (N_295,In_295,In_330);
and U296 (N_296,In_218,In_489);
and U297 (N_297,In_420,In_491);
nor U298 (N_298,In_354,In_431);
or U299 (N_299,In_103,In_396);
or U300 (N_300,In_41,In_303);
or U301 (N_301,In_115,In_268);
nand U302 (N_302,In_190,In_483);
and U303 (N_303,In_376,In_280);
and U304 (N_304,In_29,In_99);
and U305 (N_305,In_172,In_140);
and U306 (N_306,In_66,In_386);
nor U307 (N_307,In_145,In_125);
and U308 (N_308,In_53,In_39);
or U309 (N_309,In_162,In_23);
and U310 (N_310,In_350,In_178);
or U311 (N_311,In_88,In_95);
nor U312 (N_312,In_394,In_363);
and U313 (N_313,In_158,In_325);
and U314 (N_314,In_419,In_369);
nor U315 (N_315,In_236,In_254);
nand U316 (N_316,In_365,In_280);
nor U317 (N_317,In_314,In_85);
and U318 (N_318,In_33,In_200);
and U319 (N_319,In_106,In_221);
and U320 (N_320,In_210,In_255);
or U321 (N_321,In_28,In_469);
or U322 (N_322,In_114,In_37);
nor U323 (N_323,In_359,In_50);
nor U324 (N_324,In_212,In_362);
nor U325 (N_325,In_3,In_156);
and U326 (N_326,In_200,In_11);
nand U327 (N_327,In_276,In_410);
nand U328 (N_328,In_100,In_8);
or U329 (N_329,In_228,In_123);
or U330 (N_330,In_497,In_255);
or U331 (N_331,In_275,In_284);
or U332 (N_332,In_205,In_237);
nor U333 (N_333,In_176,In_234);
or U334 (N_334,In_288,In_150);
nor U335 (N_335,In_106,In_318);
or U336 (N_336,In_137,In_54);
and U337 (N_337,In_78,In_250);
nand U338 (N_338,In_254,In_271);
and U339 (N_339,In_424,In_202);
xor U340 (N_340,In_356,In_113);
or U341 (N_341,In_254,In_144);
nor U342 (N_342,In_144,In_379);
nand U343 (N_343,In_158,In_424);
or U344 (N_344,In_433,In_56);
or U345 (N_345,In_30,In_178);
or U346 (N_346,In_345,In_194);
and U347 (N_347,In_186,In_256);
or U348 (N_348,In_196,In_349);
nor U349 (N_349,In_423,In_437);
and U350 (N_350,In_195,In_212);
or U351 (N_351,In_367,In_264);
or U352 (N_352,In_8,In_203);
xnor U353 (N_353,In_54,In_345);
nor U354 (N_354,In_15,In_277);
or U355 (N_355,In_42,In_311);
or U356 (N_356,In_344,In_288);
or U357 (N_357,In_25,In_28);
nor U358 (N_358,In_56,In_496);
or U359 (N_359,In_69,In_233);
and U360 (N_360,In_481,In_371);
nor U361 (N_361,In_277,In_43);
nor U362 (N_362,In_80,In_13);
nand U363 (N_363,In_198,In_68);
and U364 (N_364,In_222,In_60);
or U365 (N_365,In_186,In_13);
and U366 (N_366,In_148,In_400);
nand U367 (N_367,In_454,In_174);
nor U368 (N_368,In_177,In_227);
nor U369 (N_369,In_2,In_55);
nor U370 (N_370,In_228,In_295);
and U371 (N_371,In_278,In_451);
nor U372 (N_372,In_110,In_223);
or U373 (N_373,In_322,In_212);
or U374 (N_374,In_496,In_492);
nand U375 (N_375,In_206,In_51);
nor U376 (N_376,In_467,In_202);
and U377 (N_377,In_119,In_372);
or U378 (N_378,In_458,In_265);
and U379 (N_379,In_68,In_482);
nand U380 (N_380,In_429,In_376);
or U381 (N_381,In_308,In_288);
nor U382 (N_382,In_495,In_168);
or U383 (N_383,In_51,In_226);
nor U384 (N_384,In_66,In_103);
or U385 (N_385,In_126,In_46);
and U386 (N_386,In_21,In_186);
nand U387 (N_387,In_201,In_428);
nand U388 (N_388,In_349,In_421);
nand U389 (N_389,In_149,In_58);
or U390 (N_390,In_329,In_201);
nor U391 (N_391,In_67,In_126);
nor U392 (N_392,In_42,In_138);
or U393 (N_393,In_358,In_486);
nor U394 (N_394,In_453,In_259);
or U395 (N_395,In_173,In_130);
or U396 (N_396,In_47,In_456);
nand U397 (N_397,In_475,In_210);
or U398 (N_398,In_395,In_290);
and U399 (N_399,In_7,In_230);
xor U400 (N_400,In_16,In_70);
nand U401 (N_401,In_324,In_427);
or U402 (N_402,In_492,In_343);
nor U403 (N_403,In_1,In_63);
nor U404 (N_404,In_442,In_244);
or U405 (N_405,In_320,In_340);
nand U406 (N_406,In_0,In_103);
nor U407 (N_407,In_481,In_61);
nor U408 (N_408,In_342,In_369);
nand U409 (N_409,In_416,In_354);
nor U410 (N_410,In_149,In_257);
nor U411 (N_411,In_245,In_54);
and U412 (N_412,In_459,In_224);
and U413 (N_413,In_181,In_104);
nand U414 (N_414,In_488,In_75);
and U415 (N_415,In_155,In_11);
nand U416 (N_416,In_237,In_483);
nand U417 (N_417,In_339,In_136);
and U418 (N_418,In_60,In_67);
nor U419 (N_419,In_162,In_93);
nand U420 (N_420,In_286,In_337);
or U421 (N_421,In_256,In_307);
nand U422 (N_422,In_30,In_96);
and U423 (N_423,In_237,In_350);
nor U424 (N_424,In_108,In_222);
or U425 (N_425,In_88,In_47);
or U426 (N_426,In_120,In_486);
and U427 (N_427,In_165,In_273);
or U428 (N_428,In_278,In_253);
nand U429 (N_429,In_420,In_99);
nor U430 (N_430,In_214,In_239);
and U431 (N_431,In_449,In_432);
or U432 (N_432,In_339,In_327);
nor U433 (N_433,In_298,In_456);
and U434 (N_434,In_337,In_318);
or U435 (N_435,In_25,In_379);
nand U436 (N_436,In_291,In_348);
nor U437 (N_437,In_431,In_112);
nand U438 (N_438,In_457,In_446);
and U439 (N_439,In_334,In_310);
nor U440 (N_440,In_265,In_435);
and U441 (N_441,In_24,In_220);
and U442 (N_442,In_11,In_496);
nor U443 (N_443,In_289,In_43);
nor U444 (N_444,In_302,In_234);
nor U445 (N_445,In_111,In_298);
or U446 (N_446,In_414,In_280);
nor U447 (N_447,In_49,In_298);
nand U448 (N_448,In_21,In_198);
and U449 (N_449,In_405,In_453);
nand U450 (N_450,In_224,In_328);
nor U451 (N_451,In_396,In_21);
or U452 (N_452,In_388,In_158);
nor U453 (N_453,In_343,In_490);
nand U454 (N_454,In_245,In_280);
and U455 (N_455,In_424,In_289);
or U456 (N_456,In_392,In_11);
nand U457 (N_457,In_338,In_489);
or U458 (N_458,In_34,In_237);
nand U459 (N_459,In_155,In_233);
or U460 (N_460,In_444,In_478);
and U461 (N_461,In_313,In_443);
and U462 (N_462,In_261,In_92);
and U463 (N_463,In_125,In_161);
nand U464 (N_464,In_0,In_101);
nor U465 (N_465,In_92,In_148);
nand U466 (N_466,In_220,In_311);
nand U467 (N_467,In_54,In_157);
nor U468 (N_468,In_105,In_329);
or U469 (N_469,In_426,In_44);
nand U470 (N_470,In_70,In_6);
nand U471 (N_471,In_362,In_326);
or U472 (N_472,In_439,In_323);
or U473 (N_473,In_35,In_329);
and U474 (N_474,In_374,In_261);
nand U475 (N_475,In_402,In_104);
or U476 (N_476,In_130,In_442);
and U477 (N_477,In_358,In_342);
nand U478 (N_478,In_340,In_466);
and U479 (N_479,In_92,In_374);
nor U480 (N_480,In_47,In_295);
nand U481 (N_481,In_259,In_238);
or U482 (N_482,In_291,In_7);
and U483 (N_483,In_311,In_310);
nor U484 (N_484,In_148,In_45);
or U485 (N_485,In_108,In_238);
or U486 (N_486,In_269,In_43);
and U487 (N_487,In_67,In_62);
or U488 (N_488,In_291,In_103);
nand U489 (N_489,In_106,In_254);
nor U490 (N_490,In_34,In_361);
and U491 (N_491,In_112,In_134);
or U492 (N_492,In_266,In_115);
or U493 (N_493,In_447,In_156);
or U494 (N_494,In_16,In_448);
nand U495 (N_495,In_387,In_60);
nor U496 (N_496,In_131,In_403);
or U497 (N_497,In_193,In_258);
nand U498 (N_498,In_473,In_181);
and U499 (N_499,In_254,In_408);
or U500 (N_500,In_122,In_292);
nand U501 (N_501,In_412,In_385);
or U502 (N_502,In_185,In_175);
and U503 (N_503,In_335,In_72);
or U504 (N_504,In_58,In_286);
nor U505 (N_505,In_373,In_240);
nand U506 (N_506,In_353,In_21);
or U507 (N_507,In_458,In_172);
nand U508 (N_508,In_208,In_165);
and U509 (N_509,In_240,In_100);
nor U510 (N_510,In_99,In_245);
or U511 (N_511,In_280,In_470);
or U512 (N_512,In_484,In_381);
nand U513 (N_513,In_148,In_404);
nand U514 (N_514,In_91,In_51);
or U515 (N_515,In_397,In_225);
nand U516 (N_516,In_329,In_381);
nor U517 (N_517,In_313,In_328);
nor U518 (N_518,In_205,In_341);
or U519 (N_519,In_358,In_83);
nor U520 (N_520,In_251,In_100);
or U521 (N_521,In_418,In_110);
and U522 (N_522,In_349,In_294);
nor U523 (N_523,In_118,In_232);
and U524 (N_524,In_157,In_31);
or U525 (N_525,In_472,In_240);
and U526 (N_526,In_449,In_53);
and U527 (N_527,In_427,In_475);
nand U528 (N_528,In_386,In_136);
and U529 (N_529,In_417,In_20);
or U530 (N_530,In_438,In_119);
nand U531 (N_531,In_86,In_116);
and U532 (N_532,In_472,In_159);
nand U533 (N_533,In_427,In_76);
and U534 (N_534,In_302,In_397);
and U535 (N_535,In_280,In_429);
or U536 (N_536,In_481,In_172);
and U537 (N_537,In_368,In_384);
xnor U538 (N_538,In_216,In_119);
and U539 (N_539,In_387,In_207);
or U540 (N_540,In_233,In_78);
and U541 (N_541,In_286,In_497);
nor U542 (N_542,In_182,In_176);
or U543 (N_543,In_102,In_185);
and U544 (N_544,In_315,In_281);
nor U545 (N_545,In_143,In_477);
nor U546 (N_546,In_130,In_107);
nor U547 (N_547,In_352,In_339);
nand U548 (N_548,In_184,In_421);
and U549 (N_549,In_171,In_253);
nand U550 (N_550,In_408,In_499);
xor U551 (N_551,In_142,In_252);
nor U552 (N_552,In_268,In_70);
and U553 (N_553,In_105,In_202);
nor U554 (N_554,In_393,In_398);
and U555 (N_555,In_411,In_203);
and U556 (N_556,In_53,In_81);
nor U557 (N_557,In_440,In_176);
or U558 (N_558,In_206,In_119);
nor U559 (N_559,In_420,In_263);
and U560 (N_560,In_324,In_10);
and U561 (N_561,In_442,In_204);
and U562 (N_562,In_72,In_429);
or U563 (N_563,In_348,In_86);
nor U564 (N_564,In_204,In_125);
or U565 (N_565,In_465,In_144);
or U566 (N_566,In_413,In_216);
and U567 (N_567,In_158,In_299);
and U568 (N_568,In_14,In_161);
nor U569 (N_569,In_373,In_29);
and U570 (N_570,In_31,In_481);
or U571 (N_571,In_495,In_226);
and U572 (N_572,In_239,In_243);
or U573 (N_573,In_312,In_248);
nand U574 (N_574,In_472,In_140);
and U575 (N_575,In_98,In_52);
nand U576 (N_576,In_473,In_294);
nand U577 (N_577,In_337,In_285);
nand U578 (N_578,In_185,In_165);
nand U579 (N_579,In_107,In_490);
and U580 (N_580,In_353,In_80);
and U581 (N_581,In_451,In_20);
or U582 (N_582,In_468,In_301);
or U583 (N_583,In_499,In_91);
or U584 (N_584,In_17,In_227);
nand U585 (N_585,In_216,In_496);
nor U586 (N_586,In_135,In_339);
nand U587 (N_587,In_117,In_63);
nand U588 (N_588,In_297,In_19);
nand U589 (N_589,In_372,In_440);
nor U590 (N_590,In_7,In_119);
and U591 (N_591,In_75,In_262);
nor U592 (N_592,In_336,In_239);
or U593 (N_593,In_297,In_486);
nor U594 (N_594,In_489,In_182);
nand U595 (N_595,In_342,In_421);
or U596 (N_596,In_201,In_285);
xnor U597 (N_597,In_240,In_79);
or U598 (N_598,In_365,In_11);
or U599 (N_599,In_114,In_350);
or U600 (N_600,In_52,In_266);
nor U601 (N_601,In_181,In_21);
and U602 (N_602,In_84,In_23);
and U603 (N_603,In_66,In_332);
nand U604 (N_604,In_279,In_492);
nand U605 (N_605,In_111,In_51);
nand U606 (N_606,In_132,In_351);
nor U607 (N_607,In_221,In_11);
and U608 (N_608,In_422,In_464);
nor U609 (N_609,In_92,In_141);
or U610 (N_610,In_483,In_325);
and U611 (N_611,In_289,In_487);
nand U612 (N_612,In_0,In_416);
and U613 (N_613,In_168,In_336);
or U614 (N_614,In_30,In_11);
nand U615 (N_615,In_401,In_490);
nand U616 (N_616,In_440,In_9);
nand U617 (N_617,In_229,In_464);
nand U618 (N_618,In_486,In_284);
nor U619 (N_619,In_67,In_269);
and U620 (N_620,In_424,In_448);
nand U621 (N_621,In_494,In_113);
nor U622 (N_622,In_316,In_293);
nor U623 (N_623,In_263,In_325);
nand U624 (N_624,In_247,In_209);
and U625 (N_625,In_247,In_95);
nand U626 (N_626,In_386,In_351);
or U627 (N_627,In_465,In_259);
and U628 (N_628,In_228,In_279);
nor U629 (N_629,In_234,In_137);
and U630 (N_630,In_153,In_266);
nor U631 (N_631,In_98,In_26);
and U632 (N_632,In_415,In_80);
nor U633 (N_633,In_220,In_341);
nand U634 (N_634,In_122,In_163);
or U635 (N_635,In_364,In_416);
nor U636 (N_636,In_35,In_490);
and U637 (N_637,In_168,In_173);
or U638 (N_638,In_274,In_125);
or U639 (N_639,In_448,In_187);
and U640 (N_640,In_452,In_356);
and U641 (N_641,In_90,In_248);
or U642 (N_642,In_303,In_6);
nor U643 (N_643,In_316,In_255);
nor U644 (N_644,In_78,In_2);
and U645 (N_645,In_465,In_42);
and U646 (N_646,In_327,In_186);
or U647 (N_647,In_182,In_416);
and U648 (N_648,In_80,In_338);
nand U649 (N_649,In_232,In_72);
or U650 (N_650,In_103,In_104);
nor U651 (N_651,In_162,In_115);
nand U652 (N_652,In_401,In_251);
nand U653 (N_653,In_262,In_276);
nor U654 (N_654,In_353,In_202);
and U655 (N_655,In_80,In_300);
nand U656 (N_656,In_115,In_94);
nand U657 (N_657,In_153,In_176);
nand U658 (N_658,In_186,In_411);
nor U659 (N_659,In_303,In_198);
or U660 (N_660,In_397,In_405);
or U661 (N_661,In_136,In_371);
nand U662 (N_662,In_13,In_482);
nor U663 (N_663,In_368,In_363);
or U664 (N_664,In_215,In_281);
or U665 (N_665,In_224,In_211);
nor U666 (N_666,In_424,In_425);
and U667 (N_667,In_234,In_124);
nand U668 (N_668,In_312,In_360);
or U669 (N_669,In_390,In_258);
nor U670 (N_670,In_195,In_289);
nand U671 (N_671,In_103,In_212);
or U672 (N_672,In_473,In_58);
or U673 (N_673,In_495,In_108);
and U674 (N_674,In_79,In_367);
nand U675 (N_675,In_332,In_190);
or U676 (N_676,In_79,In_366);
nor U677 (N_677,In_287,In_284);
and U678 (N_678,In_200,In_344);
nand U679 (N_679,In_410,In_379);
nor U680 (N_680,In_279,In_452);
nand U681 (N_681,In_182,In_441);
or U682 (N_682,In_408,In_275);
or U683 (N_683,In_278,In_476);
and U684 (N_684,In_67,In_397);
or U685 (N_685,In_335,In_111);
or U686 (N_686,In_362,In_430);
and U687 (N_687,In_411,In_196);
or U688 (N_688,In_383,In_319);
nor U689 (N_689,In_258,In_61);
nand U690 (N_690,In_107,In_29);
or U691 (N_691,In_170,In_213);
and U692 (N_692,In_403,In_437);
nor U693 (N_693,In_163,In_464);
nor U694 (N_694,In_140,In_390);
nor U695 (N_695,In_363,In_311);
nand U696 (N_696,In_44,In_261);
nand U697 (N_697,In_495,In_264);
nor U698 (N_698,In_494,In_157);
or U699 (N_699,In_174,In_189);
or U700 (N_700,In_456,In_204);
or U701 (N_701,In_80,In_443);
or U702 (N_702,In_136,In_124);
and U703 (N_703,In_374,In_430);
or U704 (N_704,In_218,In_477);
and U705 (N_705,In_375,In_159);
and U706 (N_706,In_472,In_172);
and U707 (N_707,In_275,In_461);
and U708 (N_708,In_482,In_249);
xor U709 (N_709,In_466,In_389);
or U710 (N_710,In_58,In_376);
nor U711 (N_711,In_85,In_138);
and U712 (N_712,In_448,In_79);
nor U713 (N_713,In_485,In_91);
or U714 (N_714,In_143,In_173);
and U715 (N_715,In_479,In_142);
and U716 (N_716,In_181,In_66);
nor U717 (N_717,In_118,In_267);
nor U718 (N_718,In_148,In_298);
nor U719 (N_719,In_420,In_160);
nor U720 (N_720,In_268,In_341);
or U721 (N_721,In_251,In_372);
or U722 (N_722,In_320,In_56);
nand U723 (N_723,In_301,In_5);
nor U724 (N_724,In_207,In_455);
and U725 (N_725,In_53,In_71);
and U726 (N_726,In_460,In_159);
or U727 (N_727,In_335,In_282);
and U728 (N_728,In_427,In_241);
and U729 (N_729,In_72,In_166);
nand U730 (N_730,In_202,In_412);
and U731 (N_731,In_474,In_424);
nand U732 (N_732,In_172,In_157);
nor U733 (N_733,In_357,In_203);
and U734 (N_734,In_61,In_458);
nand U735 (N_735,In_492,In_478);
nand U736 (N_736,In_301,In_216);
nor U737 (N_737,In_218,In_391);
nor U738 (N_738,In_220,In_458);
nor U739 (N_739,In_499,In_325);
and U740 (N_740,In_328,In_289);
nor U741 (N_741,In_6,In_397);
or U742 (N_742,In_228,In_129);
nor U743 (N_743,In_17,In_136);
or U744 (N_744,In_429,In_391);
nor U745 (N_745,In_386,In_79);
or U746 (N_746,In_251,In_144);
or U747 (N_747,In_238,In_467);
nand U748 (N_748,In_359,In_63);
or U749 (N_749,In_159,In_290);
and U750 (N_750,N_461,N_712);
and U751 (N_751,N_107,N_238);
nand U752 (N_752,N_569,N_646);
and U753 (N_753,N_674,N_410);
and U754 (N_754,N_636,N_320);
nand U755 (N_755,N_329,N_693);
nor U756 (N_756,N_348,N_376);
and U757 (N_757,N_552,N_747);
or U758 (N_758,N_33,N_384);
nand U759 (N_759,N_448,N_727);
nor U760 (N_760,N_23,N_432);
nand U761 (N_761,N_575,N_344);
nand U762 (N_762,N_709,N_204);
or U763 (N_763,N_2,N_267);
or U764 (N_764,N_434,N_295);
nor U765 (N_765,N_26,N_296);
and U766 (N_766,N_394,N_442);
nand U767 (N_767,N_585,N_37);
and U768 (N_768,N_655,N_325);
nand U769 (N_769,N_437,N_164);
nand U770 (N_770,N_639,N_579);
or U771 (N_771,N_472,N_492);
nand U772 (N_772,N_142,N_371);
or U773 (N_773,N_280,N_430);
nor U774 (N_774,N_463,N_563);
nor U775 (N_775,N_279,N_538);
nor U776 (N_776,N_270,N_484);
nand U777 (N_777,N_469,N_634);
nand U778 (N_778,N_245,N_20);
and U779 (N_779,N_124,N_653);
or U780 (N_780,N_161,N_734);
or U781 (N_781,N_205,N_741);
or U782 (N_782,N_166,N_532);
and U783 (N_783,N_548,N_573);
and U784 (N_784,N_732,N_198);
and U785 (N_785,N_108,N_698);
nand U786 (N_786,N_81,N_284);
nor U787 (N_787,N_379,N_18);
and U788 (N_788,N_455,N_711);
xor U789 (N_789,N_255,N_521);
nand U790 (N_790,N_452,N_578);
nand U791 (N_791,N_593,N_367);
or U792 (N_792,N_219,N_1);
nand U793 (N_793,N_592,N_386);
or U794 (N_794,N_433,N_475);
or U795 (N_795,N_453,N_723);
nand U796 (N_796,N_558,N_742);
and U797 (N_797,N_511,N_168);
and U798 (N_798,N_632,N_55);
or U799 (N_799,N_586,N_670);
and U800 (N_800,N_597,N_169);
nand U801 (N_801,N_252,N_607);
nand U802 (N_802,N_244,N_738);
or U803 (N_803,N_112,N_378);
nand U804 (N_804,N_617,N_272);
nor U805 (N_805,N_704,N_685);
nand U806 (N_806,N_400,N_323);
xnor U807 (N_807,N_393,N_612);
nand U808 (N_808,N_236,N_232);
nand U809 (N_809,N_675,N_293);
nand U810 (N_810,N_415,N_456);
or U811 (N_811,N_97,N_546);
or U812 (N_812,N_731,N_705);
nor U813 (N_813,N_743,N_744);
nand U814 (N_814,N_445,N_99);
or U815 (N_815,N_598,N_583);
or U816 (N_816,N_450,N_116);
or U817 (N_817,N_623,N_483);
and U818 (N_818,N_275,N_346);
or U819 (N_819,N_356,N_468);
and U820 (N_820,N_285,N_717);
or U821 (N_821,N_447,N_357);
or U822 (N_822,N_721,N_703);
nand U823 (N_823,N_663,N_604);
and U824 (N_824,N_369,N_534);
nor U825 (N_825,N_500,N_129);
and U826 (N_826,N_733,N_336);
and U827 (N_827,N_350,N_12);
and U828 (N_828,N_659,N_358);
and U829 (N_829,N_423,N_408);
or U830 (N_830,N_40,N_235);
nor U831 (N_831,N_694,N_94);
and U832 (N_832,N_404,N_611);
or U833 (N_833,N_673,N_264);
nor U834 (N_834,N_418,N_524);
and U835 (N_835,N_630,N_398);
nor U836 (N_836,N_222,N_446);
and U837 (N_837,N_80,N_218);
or U838 (N_838,N_93,N_605);
nor U839 (N_839,N_226,N_125);
or U840 (N_840,N_289,N_454);
nand U841 (N_841,N_749,N_726);
nand U842 (N_842,N_132,N_247);
nand U843 (N_843,N_419,N_626);
nand U844 (N_844,N_426,N_201);
nor U845 (N_845,N_78,N_702);
or U846 (N_846,N_555,N_460);
and U847 (N_847,N_234,N_34);
nand U848 (N_848,N_691,N_724);
nand U849 (N_849,N_57,N_126);
and U850 (N_850,N_225,N_206);
nor U851 (N_851,N_335,N_413);
nor U852 (N_852,N_391,N_601);
nor U853 (N_853,N_332,N_321);
or U854 (N_854,N_113,N_507);
nor U855 (N_855,N_17,N_103);
and U856 (N_856,N_523,N_417);
and U857 (N_857,N_317,N_220);
nor U858 (N_858,N_600,N_137);
nor U859 (N_859,N_495,N_282);
and U860 (N_860,N_428,N_9);
nand U861 (N_861,N_622,N_595);
nor U862 (N_862,N_118,N_457);
and U863 (N_863,N_82,N_259);
or U864 (N_864,N_624,N_525);
nor U865 (N_865,N_516,N_609);
nor U866 (N_866,N_75,N_41);
nand U867 (N_867,N_554,N_256);
nand U868 (N_868,N_735,N_635);
nor U869 (N_869,N_429,N_680);
xor U870 (N_870,N_53,N_499);
nor U871 (N_871,N_651,N_286);
or U872 (N_872,N_679,N_28);
nand U873 (N_873,N_505,N_50);
or U874 (N_874,N_581,N_713);
nor U875 (N_875,N_248,N_265);
nor U876 (N_876,N_362,N_130);
or U877 (N_877,N_76,N_146);
nand U878 (N_878,N_520,N_209);
nor U879 (N_879,N_402,N_677);
nand U880 (N_880,N_156,N_63);
nor U881 (N_881,N_425,N_544);
nand U882 (N_882,N_707,N_196);
nor U883 (N_883,N_261,N_21);
or U884 (N_884,N_668,N_397);
and U885 (N_885,N_551,N_628);
nor U886 (N_886,N_486,N_422);
and U887 (N_887,N_215,N_145);
and U888 (N_888,N_708,N_281);
nor U889 (N_889,N_331,N_533);
nand U890 (N_890,N_83,N_324);
and U891 (N_891,N_480,N_60);
and U892 (N_892,N_65,N_619);
or U893 (N_893,N_678,N_682);
and U894 (N_894,N_322,N_745);
and U895 (N_895,N_584,N_213);
nor U896 (N_896,N_566,N_514);
and U897 (N_897,N_288,N_599);
and U898 (N_898,N_545,N_621);
or U899 (N_899,N_517,N_643);
and U900 (N_900,N_462,N_86);
or U901 (N_901,N_687,N_494);
or U902 (N_902,N_52,N_212);
or U903 (N_903,N_590,N_158);
or U904 (N_904,N_3,N_345);
nor U905 (N_905,N_341,N_377);
and U906 (N_906,N_683,N_443);
nand U907 (N_907,N_412,N_90);
nand U908 (N_908,N_602,N_587);
or U909 (N_909,N_411,N_568);
nand U910 (N_910,N_313,N_334);
and U911 (N_911,N_233,N_572);
and U912 (N_912,N_383,N_138);
or U913 (N_913,N_135,N_706);
or U914 (N_914,N_186,N_361);
nor U915 (N_915,N_44,N_650);
and U916 (N_916,N_258,N_123);
or U917 (N_917,N_230,N_27);
xnor U918 (N_918,N_471,N_276);
and U919 (N_919,N_466,N_278);
or U920 (N_920,N_10,N_543);
nand U921 (N_921,N_441,N_686);
and U922 (N_922,N_305,N_487);
and U923 (N_923,N_510,N_243);
nor U924 (N_924,N_8,N_629);
and U925 (N_925,N_440,N_62);
nand U926 (N_926,N_239,N_211);
nor U927 (N_927,N_197,N_657);
or U928 (N_928,N_547,N_536);
and U929 (N_929,N_165,N_104);
nor U930 (N_930,N_491,N_102);
nor U931 (N_931,N_291,N_594);
or U932 (N_932,N_420,N_192);
nor U933 (N_933,N_254,N_737);
and U934 (N_934,N_656,N_436);
xor U935 (N_935,N_326,N_549);
nand U936 (N_936,N_22,N_181);
nand U937 (N_937,N_88,N_373);
nor U938 (N_938,N_477,N_613);
xnor U939 (N_939,N_620,N_527);
xor U940 (N_940,N_170,N_42);
or U941 (N_941,N_79,N_614);
or U942 (N_942,N_539,N_576);
nor U943 (N_943,N_45,N_180);
nand U944 (N_944,N_105,N_263);
and U945 (N_945,N_224,N_557);
nor U946 (N_946,N_25,N_515);
nand U947 (N_947,N_106,N_740);
or U948 (N_948,N_497,N_360);
nand U949 (N_949,N_38,N_644);
nand U950 (N_950,N_134,N_459);
nand U951 (N_951,N_661,N_242);
nand U952 (N_952,N_395,N_306);
and U953 (N_953,N_368,N_633);
nand U954 (N_954,N_228,N_338);
nand U955 (N_955,N_39,N_526);
nor U956 (N_956,N_355,N_406);
and U957 (N_957,N_262,N_6);
or U958 (N_958,N_409,N_110);
nor U959 (N_959,N_95,N_401);
and U960 (N_960,N_182,N_363);
nor U961 (N_961,N_308,N_310);
nand U962 (N_962,N_147,N_631);
and U963 (N_963,N_74,N_160);
nand U964 (N_964,N_474,N_638);
nand U965 (N_965,N_700,N_85);
nand U966 (N_966,N_115,N_35);
nand U967 (N_967,N_489,N_496);
nand U968 (N_968,N_405,N_307);
nand U969 (N_969,N_71,N_203);
nand U970 (N_970,N_444,N_519);
nand U971 (N_971,N_399,N_249);
nand U972 (N_972,N_47,N_513);
and U973 (N_973,N_427,N_59);
or U974 (N_974,N_375,N_266);
nand U975 (N_975,N_493,N_191);
and U976 (N_976,N_596,N_529);
and U977 (N_977,N_684,N_736);
or U978 (N_978,N_127,N_561);
and U979 (N_979,N_403,N_688);
and U980 (N_980,N_91,N_184);
nor U981 (N_981,N_542,N_501);
nand U982 (N_982,N_72,N_46);
or U983 (N_983,N_143,N_48);
nor U984 (N_984,N_370,N_518);
and U985 (N_985,N_68,N_385);
nand U986 (N_986,N_589,N_210);
or U987 (N_987,N_503,N_580);
and U988 (N_988,N_150,N_273);
or U989 (N_989,N_509,N_231);
or U990 (N_990,N_294,N_564);
and U991 (N_991,N_172,N_43);
nor U992 (N_992,N_64,N_642);
and U993 (N_993,N_550,N_465);
nand U994 (N_994,N_30,N_697);
or U995 (N_995,N_508,N_464);
or U996 (N_996,N_297,N_467);
or U997 (N_997,N_381,N_372);
or U998 (N_998,N_152,N_187);
nand U999 (N_999,N_163,N_227);
or U1000 (N_1000,N_562,N_627);
nand U1001 (N_1001,N_119,N_268);
and U1002 (N_1002,N_560,N_315);
nor U1003 (N_1003,N_214,N_140);
and U1004 (N_1004,N_716,N_333);
nand U1005 (N_1005,N_725,N_58);
nor U1006 (N_1006,N_476,N_535);
and U1007 (N_1007,N_4,N_32);
nor U1008 (N_1008,N_339,N_512);
and U1009 (N_1009,N_701,N_311);
and U1010 (N_1010,N_301,N_615);
or U1011 (N_1011,N_207,N_641);
nor U1012 (N_1012,N_365,N_720);
nand U1013 (N_1013,N_541,N_660);
or U1014 (N_1014,N_640,N_710);
nor U1015 (N_1015,N_208,N_390);
nand U1016 (N_1016,N_389,N_435);
nand U1017 (N_1017,N_151,N_342);
and U1018 (N_1018,N_251,N_148);
nor U1019 (N_1019,N_302,N_606);
and U1020 (N_1020,N_449,N_277);
or U1021 (N_1021,N_84,N_157);
nand U1022 (N_1022,N_531,N_200);
and U1023 (N_1023,N_176,N_567);
nor U1024 (N_1024,N_101,N_290);
nand U1025 (N_1025,N_353,N_392);
nand U1026 (N_1026,N_689,N_382);
or U1027 (N_1027,N_692,N_193);
and U1028 (N_1028,N_690,N_61);
and U1029 (N_1029,N_424,N_175);
or U1030 (N_1030,N_67,N_571);
nor U1031 (N_1031,N_359,N_177);
nand U1032 (N_1032,N_588,N_15);
nand U1033 (N_1033,N_155,N_73);
and U1034 (N_1034,N_0,N_319);
and U1035 (N_1035,N_24,N_648);
nand U1036 (N_1036,N_122,N_173);
and U1037 (N_1037,N_246,N_671);
or U1038 (N_1038,N_167,N_221);
nand U1039 (N_1039,N_292,N_714);
nand U1040 (N_1040,N_637,N_695);
nor U1041 (N_1041,N_274,N_349);
nor U1042 (N_1042,N_618,N_616);
nand U1043 (N_1043,N_504,N_318);
nor U1044 (N_1044,N_250,N_330);
nand U1045 (N_1045,N_316,N_298);
or U1046 (N_1046,N_388,N_458);
and U1047 (N_1047,N_139,N_488);
nand U1048 (N_1048,N_287,N_240);
or U1049 (N_1049,N_652,N_347);
nand U1050 (N_1050,N_387,N_216);
nand U1051 (N_1051,N_540,N_14);
or U1052 (N_1052,N_739,N_431);
or U1053 (N_1053,N_195,N_87);
and U1054 (N_1054,N_662,N_49);
and U1055 (N_1055,N_194,N_269);
nand U1056 (N_1056,N_189,N_352);
nand U1057 (N_1057,N_672,N_374);
or U1058 (N_1058,N_11,N_51);
nor U1059 (N_1059,N_625,N_153);
nor U1060 (N_1060,N_328,N_591);
nor U1061 (N_1061,N_96,N_131);
and U1062 (N_1062,N_699,N_676);
or U1063 (N_1063,N_141,N_380);
nor U1064 (N_1064,N_223,N_647);
nand U1065 (N_1065,N_128,N_610);
or U1066 (N_1066,N_77,N_715);
or U1067 (N_1067,N_482,N_414);
nor U1068 (N_1068,N_603,N_506);
nor U1069 (N_1069,N_522,N_577);
and U1070 (N_1070,N_666,N_681);
nor U1071 (N_1071,N_304,N_645);
and U1072 (N_1072,N_649,N_451);
nor U1073 (N_1073,N_730,N_7);
and U1074 (N_1074,N_29,N_343);
nand U1075 (N_1075,N_309,N_667);
or U1076 (N_1076,N_479,N_217);
nand U1077 (N_1077,N_179,N_438);
nand U1078 (N_1078,N_260,N_185);
or U1079 (N_1079,N_31,N_162);
and U1080 (N_1080,N_556,N_416);
nand U1081 (N_1081,N_188,N_149);
and U1082 (N_1082,N_364,N_574);
or U1083 (N_1083,N_237,N_565);
and U1084 (N_1084,N_111,N_229);
nor U1085 (N_1085,N_98,N_748);
nand U1086 (N_1086,N_54,N_654);
nand U1087 (N_1087,N_69,N_396);
nand U1088 (N_1088,N_354,N_89);
nand U1089 (N_1089,N_120,N_746);
nand U1090 (N_1090,N_257,N_669);
or U1091 (N_1091,N_473,N_327);
nor U1092 (N_1092,N_478,N_722);
or U1093 (N_1093,N_154,N_337);
xor U1094 (N_1094,N_582,N_481);
nand U1095 (N_1095,N_718,N_485);
and U1096 (N_1096,N_117,N_144);
nor U1097 (N_1097,N_178,N_13);
and U1098 (N_1098,N_299,N_241);
nand U1099 (N_1099,N_190,N_559);
or U1100 (N_1100,N_5,N_253);
nor U1101 (N_1101,N_199,N_439);
nor U1102 (N_1102,N_303,N_421);
nand U1103 (N_1103,N_340,N_696);
and U1104 (N_1104,N_202,N_470);
or U1105 (N_1105,N_183,N_133);
or U1106 (N_1106,N_490,N_553);
or U1107 (N_1107,N_66,N_136);
nor U1108 (N_1108,N_608,N_16);
and U1109 (N_1109,N_366,N_56);
and U1110 (N_1110,N_300,N_36);
or U1111 (N_1111,N_498,N_537);
or U1112 (N_1112,N_92,N_271);
and U1113 (N_1113,N_719,N_109);
nor U1114 (N_1114,N_19,N_283);
nor U1115 (N_1115,N_159,N_174);
or U1116 (N_1116,N_114,N_729);
and U1117 (N_1117,N_407,N_528);
and U1118 (N_1118,N_658,N_665);
or U1119 (N_1119,N_502,N_664);
nor U1120 (N_1120,N_312,N_70);
nor U1121 (N_1121,N_530,N_351);
nand U1122 (N_1122,N_570,N_314);
nand U1123 (N_1123,N_171,N_728);
and U1124 (N_1124,N_100,N_121);
or U1125 (N_1125,N_143,N_127);
nand U1126 (N_1126,N_592,N_601);
or U1127 (N_1127,N_731,N_48);
or U1128 (N_1128,N_387,N_552);
or U1129 (N_1129,N_198,N_102);
or U1130 (N_1130,N_3,N_687);
and U1131 (N_1131,N_546,N_104);
nand U1132 (N_1132,N_567,N_330);
nand U1133 (N_1133,N_560,N_312);
nor U1134 (N_1134,N_30,N_117);
or U1135 (N_1135,N_254,N_616);
nor U1136 (N_1136,N_24,N_511);
and U1137 (N_1137,N_367,N_557);
nand U1138 (N_1138,N_746,N_298);
and U1139 (N_1139,N_237,N_120);
and U1140 (N_1140,N_447,N_387);
nor U1141 (N_1141,N_79,N_61);
nand U1142 (N_1142,N_652,N_496);
and U1143 (N_1143,N_352,N_701);
or U1144 (N_1144,N_72,N_93);
and U1145 (N_1145,N_611,N_729);
nor U1146 (N_1146,N_281,N_68);
xnor U1147 (N_1147,N_550,N_710);
nand U1148 (N_1148,N_286,N_138);
nand U1149 (N_1149,N_86,N_53);
and U1150 (N_1150,N_368,N_469);
nand U1151 (N_1151,N_211,N_576);
or U1152 (N_1152,N_595,N_121);
nor U1153 (N_1153,N_540,N_562);
or U1154 (N_1154,N_440,N_119);
and U1155 (N_1155,N_705,N_200);
and U1156 (N_1156,N_635,N_441);
and U1157 (N_1157,N_60,N_590);
and U1158 (N_1158,N_123,N_695);
nand U1159 (N_1159,N_302,N_49);
and U1160 (N_1160,N_514,N_722);
nand U1161 (N_1161,N_617,N_253);
nor U1162 (N_1162,N_40,N_85);
nand U1163 (N_1163,N_640,N_601);
nand U1164 (N_1164,N_684,N_466);
and U1165 (N_1165,N_345,N_54);
nor U1166 (N_1166,N_34,N_591);
nor U1167 (N_1167,N_420,N_143);
nand U1168 (N_1168,N_650,N_712);
nor U1169 (N_1169,N_553,N_435);
nor U1170 (N_1170,N_664,N_417);
or U1171 (N_1171,N_732,N_38);
or U1172 (N_1172,N_415,N_153);
and U1173 (N_1173,N_628,N_631);
nand U1174 (N_1174,N_477,N_712);
and U1175 (N_1175,N_524,N_573);
nor U1176 (N_1176,N_609,N_31);
nand U1177 (N_1177,N_86,N_525);
nor U1178 (N_1178,N_266,N_298);
or U1179 (N_1179,N_83,N_654);
or U1180 (N_1180,N_489,N_523);
or U1181 (N_1181,N_17,N_73);
or U1182 (N_1182,N_182,N_113);
nor U1183 (N_1183,N_591,N_327);
nand U1184 (N_1184,N_563,N_704);
and U1185 (N_1185,N_644,N_544);
nor U1186 (N_1186,N_159,N_28);
and U1187 (N_1187,N_408,N_209);
nor U1188 (N_1188,N_409,N_569);
nor U1189 (N_1189,N_170,N_629);
nor U1190 (N_1190,N_466,N_377);
nor U1191 (N_1191,N_254,N_473);
or U1192 (N_1192,N_199,N_542);
or U1193 (N_1193,N_136,N_688);
or U1194 (N_1194,N_737,N_46);
nand U1195 (N_1195,N_447,N_279);
or U1196 (N_1196,N_514,N_333);
nand U1197 (N_1197,N_310,N_328);
nand U1198 (N_1198,N_642,N_46);
nand U1199 (N_1199,N_388,N_703);
and U1200 (N_1200,N_294,N_721);
or U1201 (N_1201,N_375,N_123);
nand U1202 (N_1202,N_335,N_176);
and U1203 (N_1203,N_208,N_323);
and U1204 (N_1204,N_507,N_84);
nand U1205 (N_1205,N_520,N_586);
nor U1206 (N_1206,N_735,N_4);
and U1207 (N_1207,N_238,N_395);
nand U1208 (N_1208,N_713,N_727);
or U1209 (N_1209,N_99,N_362);
nand U1210 (N_1210,N_739,N_724);
and U1211 (N_1211,N_575,N_336);
nor U1212 (N_1212,N_192,N_645);
or U1213 (N_1213,N_711,N_618);
or U1214 (N_1214,N_382,N_28);
nand U1215 (N_1215,N_185,N_329);
or U1216 (N_1216,N_534,N_118);
or U1217 (N_1217,N_735,N_493);
nand U1218 (N_1218,N_288,N_350);
and U1219 (N_1219,N_136,N_210);
nand U1220 (N_1220,N_565,N_388);
and U1221 (N_1221,N_432,N_294);
or U1222 (N_1222,N_332,N_649);
nand U1223 (N_1223,N_76,N_75);
nand U1224 (N_1224,N_700,N_367);
nand U1225 (N_1225,N_150,N_9);
and U1226 (N_1226,N_520,N_652);
nor U1227 (N_1227,N_184,N_215);
and U1228 (N_1228,N_137,N_495);
nor U1229 (N_1229,N_107,N_706);
or U1230 (N_1230,N_542,N_418);
and U1231 (N_1231,N_122,N_643);
nand U1232 (N_1232,N_698,N_613);
nand U1233 (N_1233,N_529,N_141);
or U1234 (N_1234,N_100,N_301);
or U1235 (N_1235,N_227,N_644);
and U1236 (N_1236,N_582,N_392);
nor U1237 (N_1237,N_377,N_571);
nor U1238 (N_1238,N_76,N_261);
or U1239 (N_1239,N_29,N_80);
or U1240 (N_1240,N_94,N_227);
and U1241 (N_1241,N_611,N_417);
nand U1242 (N_1242,N_57,N_351);
or U1243 (N_1243,N_454,N_467);
nor U1244 (N_1244,N_185,N_167);
nand U1245 (N_1245,N_361,N_214);
and U1246 (N_1246,N_449,N_116);
nand U1247 (N_1247,N_717,N_649);
or U1248 (N_1248,N_147,N_106);
and U1249 (N_1249,N_232,N_159);
nor U1250 (N_1250,N_549,N_381);
nor U1251 (N_1251,N_36,N_701);
and U1252 (N_1252,N_90,N_400);
nand U1253 (N_1253,N_52,N_359);
or U1254 (N_1254,N_241,N_283);
and U1255 (N_1255,N_243,N_333);
nor U1256 (N_1256,N_532,N_224);
or U1257 (N_1257,N_547,N_349);
and U1258 (N_1258,N_22,N_432);
or U1259 (N_1259,N_38,N_117);
or U1260 (N_1260,N_368,N_253);
or U1261 (N_1261,N_693,N_646);
nand U1262 (N_1262,N_143,N_300);
and U1263 (N_1263,N_390,N_107);
or U1264 (N_1264,N_184,N_519);
nor U1265 (N_1265,N_239,N_737);
and U1266 (N_1266,N_416,N_160);
or U1267 (N_1267,N_711,N_300);
and U1268 (N_1268,N_29,N_304);
and U1269 (N_1269,N_263,N_588);
nand U1270 (N_1270,N_271,N_688);
nand U1271 (N_1271,N_314,N_108);
or U1272 (N_1272,N_262,N_48);
and U1273 (N_1273,N_527,N_574);
nor U1274 (N_1274,N_591,N_250);
and U1275 (N_1275,N_417,N_321);
nand U1276 (N_1276,N_34,N_364);
xnor U1277 (N_1277,N_469,N_624);
or U1278 (N_1278,N_266,N_710);
or U1279 (N_1279,N_247,N_90);
nor U1280 (N_1280,N_398,N_443);
nor U1281 (N_1281,N_677,N_324);
and U1282 (N_1282,N_221,N_274);
and U1283 (N_1283,N_164,N_61);
or U1284 (N_1284,N_335,N_669);
xnor U1285 (N_1285,N_379,N_707);
nand U1286 (N_1286,N_582,N_71);
nand U1287 (N_1287,N_605,N_474);
nor U1288 (N_1288,N_62,N_294);
nor U1289 (N_1289,N_448,N_684);
or U1290 (N_1290,N_372,N_571);
and U1291 (N_1291,N_661,N_148);
nand U1292 (N_1292,N_667,N_3);
nand U1293 (N_1293,N_363,N_315);
and U1294 (N_1294,N_157,N_588);
or U1295 (N_1295,N_600,N_727);
or U1296 (N_1296,N_742,N_120);
or U1297 (N_1297,N_741,N_35);
nor U1298 (N_1298,N_302,N_602);
nand U1299 (N_1299,N_384,N_268);
and U1300 (N_1300,N_188,N_53);
nand U1301 (N_1301,N_419,N_582);
nand U1302 (N_1302,N_246,N_148);
and U1303 (N_1303,N_158,N_140);
or U1304 (N_1304,N_728,N_366);
nor U1305 (N_1305,N_464,N_215);
nor U1306 (N_1306,N_612,N_398);
and U1307 (N_1307,N_208,N_604);
nand U1308 (N_1308,N_87,N_170);
nand U1309 (N_1309,N_72,N_740);
or U1310 (N_1310,N_586,N_53);
nand U1311 (N_1311,N_746,N_112);
and U1312 (N_1312,N_446,N_159);
nand U1313 (N_1313,N_317,N_60);
or U1314 (N_1314,N_6,N_616);
nor U1315 (N_1315,N_194,N_696);
and U1316 (N_1316,N_297,N_292);
nand U1317 (N_1317,N_161,N_126);
nand U1318 (N_1318,N_217,N_710);
or U1319 (N_1319,N_6,N_309);
nor U1320 (N_1320,N_251,N_385);
nor U1321 (N_1321,N_524,N_407);
or U1322 (N_1322,N_97,N_424);
and U1323 (N_1323,N_407,N_628);
nor U1324 (N_1324,N_382,N_175);
and U1325 (N_1325,N_453,N_57);
nand U1326 (N_1326,N_623,N_329);
nand U1327 (N_1327,N_718,N_195);
or U1328 (N_1328,N_667,N_625);
nand U1329 (N_1329,N_239,N_3);
nor U1330 (N_1330,N_520,N_47);
nand U1331 (N_1331,N_595,N_285);
or U1332 (N_1332,N_138,N_167);
and U1333 (N_1333,N_157,N_283);
or U1334 (N_1334,N_109,N_536);
and U1335 (N_1335,N_390,N_439);
nand U1336 (N_1336,N_256,N_114);
and U1337 (N_1337,N_6,N_604);
and U1338 (N_1338,N_522,N_644);
or U1339 (N_1339,N_487,N_718);
nand U1340 (N_1340,N_293,N_267);
xor U1341 (N_1341,N_732,N_258);
nor U1342 (N_1342,N_536,N_454);
or U1343 (N_1343,N_578,N_135);
nand U1344 (N_1344,N_133,N_264);
and U1345 (N_1345,N_571,N_186);
and U1346 (N_1346,N_451,N_584);
nor U1347 (N_1347,N_357,N_285);
nor U1348 (N_1348,N_184,N_565);
nand U1349 (N_1349,N_22,N_254);
nand U1350 (N_1350,N_341,N_340);
and U1351 (N_1351,N_577,N_217);
nor U1352 (N_1352,N_318,N_492);
nand U1353 (N_1353,N_119,N_275);
or U1354 (N_1354,N_425,N_616);
xor U1355 (N_1355,N_727,N_406);
nand U1356 (N_1356,N_329,N_64);
or U1357 (N_1357,N_395,N_685);
nor U1358 (N_1358,N_58,N_331);
nor U1359 (N_1359,N_325,N_367);
or U1360 (N_1360,N_374,N_245);
and U1361 (N_1361,N_331,N_568);
and U1362 (N_1362,N_388,N_224);
and U1363 (N_1363,N_452,N_196);
nand U1364 (N_1364,N_723,N_676);
and U1365 (N_1365,N_34,N_671);
and U1366 (N_1366,N_681,N_385);
and U1367 (N_1367,N_593,N_702);
nand U1368 (N_1368,N_174,N_463);
and U1369 (N_1369,N_524,N_1);
nor U1370 (N_1370,N_95,N_334);
nor U1371 (N_1371,N_516,N_213);
or U1372 (N_1372,N_142,N_456);
nand U1373 (N_1373,N_241,N_294);
nand U1374 (N_1374,N_563,N_503);
nor U1375 (N_1375,N_657,N_687);
and U1376 (N_1376,N_719,N_225);
nor U1377 (N_1377,N_138,N_323);
nand U1378 (N_1378,N_138,N_75);
nor U1379 (N_1379,N_418,N_490);
and U1380 (N_1380,N_733,N_628);
and U1381 (N_1381,N_198,N_401);
nor U1382 (N_1382,N_286,N_216);
or U1383 (N_1383,N_541,N_462);
or U1384 (N_1384,N_88,N_136);
nand U1385 (N_1385,N_415,N_702);
nand U1386 (N_1386,N_724,N_189);
or U1387 (N_1387,N_456,N_367);
nand U1388 (N_1388,N_392,N_40);
nor U1389 (N_1389,N_254,N_104);
or U1390 (N_1390,N_96,N_191);
and U1391 (N_1391,N_577,N_680);
or U1392 (N_1392,N_50,N_533);
and U1393 (N_1393,N_481,N_357);
or U1394 (N_1394,N_378,N_497);
nand U1395 (N_1395,N_205,N_481);
and U1396 (N_1396,N_563,N_376);
nor U1397 (N_1397,N_424,N_711);
nor U1398 (N_1398,N_216,N_243);
nor U1399 (N_1399,N_626,N_58);
nand U1400 (N_1400,N_4,N_323);
nand U1401 (N_1401,N_466,N_700);
nand U1402 (N_1402,N_738,N_292);
or U1403 (N_1403,N_523,N_436);
nor U1404 (N_1404,N_346,N_566);
or U1405 (N_1405,N_117,N_368);
xor U1406 (N_1406,N_674,N_198);
nor U1407 (N_1407,N_147,N_230);
or U1408 (N_1408,N_33,N_604);
or U1409 (N_1409,N_425,N_392);
nand U1410 (N_1410,N_242,N_674);
or U1411 (N_1411,N_164,N_508);
and U1412 (N_1412,N_535,N_600);
and U1413 (N_1413,N_732,N_343);
nand U1414 (N_1414,N_154,N_419);
and U1415 (N_1415,N_89,N_594);
nand U1416 (N_1416,N_495,N_3);
or U1417 (N_1417,N_299,N_639);
nor U1418 (N_1418,N_70,N_556);
nor U1419 (N_1419,N_412,N_171);
or U1420 (N_1420,N_78,N_165);
and U1421 (N_1421,N_389,N_367);
and U1422 (N_1422,N_462,N_634);
and U1423 (N_1423,N_300,N_644);
nor U1424 (N_1424,N_22,N_398);
or U1425 (N_1425,N_515,N_437);
nand U1426 (N_1426,N_473,N_156);
or U1427 (N_1427,N_174,N_610);
or U1428 (N_1428,N_300,N_484);
nand U1429 (N_1429,N_77,N_551);
nand U1430 (N_1430,N_51,N_749);
or U1431 (N_1431,N_369,N_511);
and U1432 (N_1432,N_743,N_400);
nand U1433 (N_1433,N_40,N_221);
nand U1434 (N_1434,N_375,N_516);
and U1435 (N_1435,N_328,N_97);
nand U1436 (N_1436,N_645,N_182);
or U1437 (N_1437,N_85,N_185);
or U1438 (N_1438,N_157,N_744);
and U1439 (N_1439,N_216,N_217);
nor U1440 (N_1440,N_470,N_307);
or U1441 (N_1441,N_110,N_459);
or U1442 (N_1442,N_220,N_676);
nor U1443 (N_1443,N_258,N_192);
and U1444 (N_1444,N_84,N_578);
nand U1445 (N_1445,N_367,N_6);
nand U1446 (N_1446,N_346,N_549);
nor U1447 (N_1447,N_320,N_494);
and U1448 (N_1448,N_735,N_638);
or U1449 (N_1449,N_584,N_609);
and U1450 (N_1450,N_633,N_183);
nand U1451 (N_1451,N_269,N_738);
and U1452 (N_1452,N_568,N_705);
nand U1453 (N_1453,N_444,N_711);
or U1454 (N_1454,N_433,N_22);
and U1455 (N_1455,N_462,N_23);
nand U1456 (N_1456,N_78,N_131);
nand U1457 (N_1457,N_331,N_708);
nor U1458 (N_1458,N_378,N_379);
nand U1459 (N_1459,N_206,N_205);
nand U1460 (N_1460,N_138,N_474);
and U1461 (N_1461,N_740,N_288);
and U1462 (N_1462,N_674,N_720);
and U1463 (N_1463,N_707,N_559);
nor U1464 (N_1464,N_607,N_285);
nor U1465 (N_1465,N_121,N_450);
nand U1466 (N_1466,N_87,N_241);
xor U1467 (N_1467,N_436,N_208);
or U1468 (N_1468,N_413,N_647);
or U1469 (N_1469,N_29,N_662);
and U1470 (N_1470,N_55,N_522);
nor U1471 (N_1471,N_347,N_85);
nor U1472 (N_1472,N_574,N_360);
nor U1473 (N_1473,N_495,N_250);
and U1474 (N_1474,N_336,N_91);
nor U1475 (N_1475,N_25,N_187);
nand U1476 (N_1476,N_294,N_492);
nor U1477 (N_1477,N_89,N_31);
and U1478 (N_1478,N_264,N_280);
and U1479 (N_1479,N_540,N_512);
nor U1480 (N_1480,N_202,N_76);
nand U1481 (N_1481,N_517,N_195);
nand U1482 (N_1482,N_31,N_706);
nor U1483 (N_1483,N_168,N_407);
or U1484 (N_1484,N_667,N_257);
nor U1485 (N_1485,N_742,N_642);
nor U1486 (N_1486,N_133,N_653);
nand U1487 (N_1487,N_228,N_415);
nor U1488 (N_1488,N_621,N_132);
nand U1489 (N_1489,N_664,N_276);
nor U1490 (N_1490,N_733,N_238);
or U1491 (N_1491,N_88,N_517);
nor U1492 (N_1492,N_177,N_241);
xnor U1493 (N_1493,N_406,N_118);
nand U1494 (N_1494,N_28,N_315);
nor U1495 (N_1495,N_450,N_599);
and U1496 (N_1496,N_232,N_283);
and U1497 (N_1497,N_649,N_385);
nor U1498 (N_1498,N_399,N_722);
nand U1499 (N_1499,N_683,N_136);
or U1500 (N_1500,N_1132,N_1100);
or U1501 (N_1501,N_1400,N_1351);
and U1502 (N_1502,N_948,N_1133);
nor U1503 (N_1503,N_1181,N_1069);
and U1504 (N_1504,N_1124,N_932);
and U1505 (N_1505,N_1269,N_1194);
and U1506 (N_1506,N_1396,N_1083);
or U1507 (N_1507,N_899,N_865);
and U1508 (N_1508,N_1322,N_866);
and U1509 (N_1509,N_1496,N_851);
nor U1510 (N_1510,N_1020,N_1289);
nor U1511 (N_1511,N_1432,N_1393);
or U1512 (N_1512,N_933,N_950);
and U1513 (N_1513,N_971,N_1366);
and U1514 (N_1514,N_837,N_999);
nand U1515 (N_1515,N_773,N_965);
nor U1516 (N_1516,N_1300,N_1471);
nand U1517 (N_1517,N_1098,N_1424);
nand U1518 (N_1518,N_855,N_1097);
nand U1519 (N_1519,N_1439,N_1392);
nor U1520 (N_1520,N_1349,N_1378);
or U1521 (N_1521,N_1058,N_1105);
and U1522 (N_1522,N_1182,N_1456);
or U1523 (N_1523,N_1174,N_1332);
or U1524 (N_1524,N_990,N_1316);
nand U1525 (N_1525,N_1409,N_1075);
nand U1526 (N_1526,N_896,N_1157);
nor U1527 (N_1527,N_1281,N_1472);
or U1528 (N_1528,N_1338,N_1186);
and U1529 (N_1529,N_1175,N_1234);
and U1530 (N_1530,N_1272,N_1382);
nor U1531 (N_1531,N_1017,N_923);
nand U1532 (N_1532,N_996,N_929);
and U1533 (N_1533,N_1296,N_1379);
nor U1534 (N_1534,N_880,N_1423);
or U1535 (N_1535,N_1290,N_1141);
or U1536 (N_1536,N_1150,N_1346);
and U1537 (N_1537,N_1035,N_869);
or U1538 (N_1538,N_1421,N_856);
and U1539 (N_1539,N_1203,N_963);
nor U1540 (N_1540,N_1275,N_995);
and U1541 (N_1541,N_810,N_1023);
nor U1542 (N_1542,N_1301,N_1498);
or U1543 (N_1543,N_1119,N_1386);
nand U1544 (N_1544,N_1276,N_815);
nor U1545 (N_1545,N_1024,N_1079);
nor U1546 (N_1546,N_1266,N_821);
or U1547 (N_1547,N_883,N_1044);
nor U1548 (N_1548,N_1013,N_1220);
and U1549 (N_1549,N_926,N_889);
nor U1550 (N_1550,N_1110,N_1214);
and U1551 (N_1551,N_1031,N_1096);
or U1552 (N_1552,N_1018,N_1304);
nand U1553 (N_1553,N_1254,N_986);
and U1554 (N_1554,N_1491,N_1347);
nor U1555 (N_1555,N_1122,N_775);
nor U1556 (N_1556,N_1371,N_1000);
nand U1557 (N_1557,N_1059,N_812);
or U1558 (N_1558,N_843,N_1321);
and U1559 (N_1559,N_983,N_1412);
or U1560 (N_1560,N_788,N_1253);
and U1561 (N_1561,N_1185,N_994);
nor U1562 (N_1562,N_1232,N_1015);
nand U1563 (N_1563,N_1457,N_1162);
nor U1564 (N_1564,N_868,N_1435);
and U1565 (N_1565,N_864,N_1241);
and U1566 (N_1566,N_1206,N_1411);
nor U1567 (N_1567,N_787,N_894);
and U1568 (N_1568,N_1192,N_1052);
nand U1569 (N_1569,N_960,N_879);
or U1570 (N_1570,N_1271,N_1144);
and U1571 (N_1571,N_826,N_946);
nor U1572 (N_1572,N_1299,N_1273);
and U1573 (N_1573,N_1292,N_1065);
nand U1574 (N_1574,N_1312,N_1030);
and U1575 (N_1575,N_1309,N_840);
and U1576 (N_1576,N_819,N_1436);
nand U1577 (N_1577,N_940,N_1270);
or U1578 (N_1578,N_1198,N_874);
nand U1579 (N_1579,N_814,N_1061);
nor U1580 (N_1580,N_791,N_1111);
nor U1581 (N_1581,N_1293,N_1212);
nand U1582 (N_1582,N_1414,N_1369);
nand U1583 (N_1583,N_1437,N_1106);
and U1584 (N_1584,N_1121,N_1389);
and U1585 (N_1585,N_1342,N_786);
nand U1586 (N_1586,N_952,N_951);
or U1587 (N_1587,N_873,N_915);
nand U1588 (N_1588,N_888,N_1138);
or U1589 (N_1589,N_763,N_959);
nor U1590 (N_1590,N_800,N_1315);
nor U1591 (N_1591,N_1189,N_780);
and U1592 (N_1592,N_1323,N_799);
nand U1593 (N_1593,N_774,N_881);
and U1594 (N_1594,N_1455,N_1166);
nor U1595 (N_1595,N_1135,N_1217);
xnor U1596 (N_1596,N_887,N_809);
xor U1597 (N_1597,N_1391,N_1209);
nand U1598 (N_1598,N_1360,N_858);
or U1599 (N_1599,N_830,N_750);
nand U1600 (N_1600,N_920,N_1442);
nand U1601 (N_1601,N_1376,N_1385);
xor U1602 (N_1602,N_1464,N_1444);
nand U1603 (N_1603,N_1104,N_1359);
and U1604 (N_1604,N_1196,N_1011);
or U1605 (N_1605,N_973,N_1090);
and U1606 (N_1606,N_991,N_1427);
nor U1607 (N_1607,N_759,N_967);
and U1608 (N_1608,N_1470,N_939);
or U1609 (N_1609,N_934,N_1302);
xor U1610 (N_1610,N_975,N_1005);
nand U1611 (N_1611,N_1449,N_1026);
nand U1612 (N_1612,N_1358,N_1045);
nor U1613 (N_1613,N_901,N_1319);
nor U1614 (N_1614,N_1218,N_980);
or U1615 (N_1615,N_1226,N_878);
and U1616 (N_1616,N_1154,N_1365);
nand U1617 (N_1617,N_925,N_1481);
or U1618 (N_1618,N_1343,N_1328);
nand U1619 (N_1619,N_1043,N_779);
nor U1620 (N_1620,N_935,N_968);
nor U1621 (N_1621,N_1397,N_1229);
or U1622 (N_1622,N_798,N_1487);
or U1623 (N_1623,N_998,N_1350);
and U1624 (N_1624,N_1200,N_922);
and U1625 (N_1625,N_801,N_1329);
and U1626 (N_1626,N_957,N_941);
nor U1627 (N_1627,N_1330,N_1418);
and U1628 (N_1628,N_1048,N_1362);
nor U1629 (N_1629,N_1134,N_1327);
nand U1630 (N_1630,N_1081,N_962);
nand U1631 (N_1631,N_789,N_870);
and U1632 (N_1632,N_1443,N_1248);
or U1633 (N_1633,N_1032,N_1406);
or U1634 (N_1634,N_927,N_921);
nand U1635 (N_1635,N_909,N_1142);
nand U1636 (N_1636,N_1469,N_1477);
or U1637 (N_1637,N_877,N_1473);
and U1638 (N_1638,N_1039,N_984);
nor U1639 (N_1639,N_769,N_924);
nor U1640 (N_1640,N_958,N_1430);
or U1641 (N_1641,N_988,N_1384);
nand U1642 (N_1642,N_1148,N_1037);
nand U1643 (N_1643,N_811,N_1262);
and U1644 (N_1644,N_908,N_1102);
nor U1645 (N_1645,N_1107,N_1120);
and U1646 (N_1646,N_842,N_1419);
nor U1647 (N_1647,N_846,N_1308);
and U1648 (N_1648,N_1155,N_772);
nor U1649 (N_1649,N_1341,N_1402);
or U1650 (N_1650,N_1260,N_1067);
and U1651 (N_1651,N_1215,N_838);
nor U1652 (N_1652,N_1373,N_862);
nand U1653 (N_1653,N_832,N_1264);
nor U1654 (N_1654,N_1152,N_1036);
nor U1655 (N_1655,N_1176,N_848);
nor U1656 (N_1656,N_804,N_1465);
nor U1657 (N_1657,N_1288,N_1183);
nand U1658 (N_1658,N_1277,N_972);
nor U1659 (N_1659,N_1213,N_914);
nor U1660 (N_1660,N_1195,N_1029);
nor U1661 (N_1661,N_860,N_757);
or U1662 (N_1662,N_1094,N_1490);
or U1663 (N_1663,N_1187,N_1320);
nor U1664 (N_1664,N_1250,N_805);
nand U1665 (N_1665,N_1398,N_1497);
nand U1666 (N_1666,N_942,N_1178);
or U1667 (N_1667,N_1259,N_1025);
or U1668 (N_1668,N_847,N_1433);
nand U1669 (N_1669,N_1452,N_1261);
and U1670 (N_1670,N_1056,N_1249);
or U1671 (N_1671,N_1172,N_1165);
and U1672 (N_1672,N_793,N_824);
nand U1673 (N_1673,N_893,N_1395);
nand U1674 (N_1674,N_1388,N_1093);
or U1675 (N_1675,N_1072,N_1179);
nand U1676 (N_1676,N_1171,N_857);
or U1677 (N_1677,N_1053,N_1014);
and U1678 (N_1678,N_1480,N_1243);
nand U1679 (N_1679,N_1156,N_1231);
nand U1680 (N_1680,N_1363,N_1066);
and U1681 (N_1681,N_978,N_930);
nand U1682 (N_1682,N_977,N_974);
and U1683 (N_1683,N_1246,N_1137);
and U1684 (N_1684,N_1108,N_913);
or U1685 (N_1685,N_902,N_956);
nor U1686 (N_1686,N_1028,N_849);
nor U1687 (N_1687,N_1394,N_776);
nor U1688 (N_1688,N_1303,N_755);
or U1689 (N_1689,N_1242,N_1168);
nand U1690 (N_1690,N_756,N_820);
nand U1691 (N_1691,N_807,N_1461);
nand U1692 (N_1692,N_1230,N_1112);
nand U1693 (N_1693,N_1344,N_949);
nor U1694 (N_1694,N_1415,N_1445);
nor U1695 (N_1695,N_854,N_816);
nor U1696 (N_1696,N_1208,N_912);
or U1697 (N_1697,N_1184,N_1074);
nor U1698 (N_1698,N_1493,N_872);
or U1699 (N_1699,N_911,N_1311);
or U1700 (N_1700,N_753,N_1492);
nand U1701 (N_1701,N_936,N_1170);
nand U1702 (N_1702,N_1008,N_891);
nor U1703 (N_1703,N_1268,N_841);
nand U1704 (N_1704,N_1438,N_785);
xor U1705 (N_1705,N_1305,N_917);
and U1706 (N_1706,N_1140,N_1314);
nor U1707 (N_1707,N_985,N_1012);
and U1708 (N_1708,N_1280,N_1219);
or U1709 (N_1709,N_1339,N_953);
nor U1710 (N_1710,N_1434,N_1125);
nand U1711 (N_1711,N_795,N_1495);
nor U1712 (N_1712,N_1294,N_836);
nand U1713 (N_1713,N_1129,N_1016);
or U1714 (N_1714,N_1380,N_1127);
and U1715 (N_1715,N_1115,N_1278);
and U1716 (N_1716,N_1291,N_1282);
or U1717 (N_1717,N_989,N_1085);
and U1718 (N_1718,N_898,N_1033);
or U1719 (N_1719,N_1001,N_1286);
nor U1720 (N_1720,N_919,N_1431);
or U1721 (N_1721,N_1224,N_1190);
and U1722 (N_1722,N_876,N_803);
nand U1723 (N_1723,N_1364,N_1163);
nor U1724 (N_1724,N_931,N_1352);
or U1725 (N_1725,N_1420,N_1089);
nand U1726 (N_1726,N_1482,N_1313);
nor U1727 (N_1727,N_937,N_938);
nor U1728 (N_1728,N_1454,N_859);
nor U1729 (N_1729,N_758,N_1051);
or U1730 (N_1730,N_1310,N_1054);
nor U1731 (N_1731,N_1126,N_890);
and U1732 (N_1732,N_1007,N_1354);
or U1733 (N_1733,N_1034,N_1447);
or U1734 (N_1734,N_790,N_861);
nor U1735 (N_1735,N_863,N_1188);
and U1736 (N_1736,N_875,N_1370);
or U1737 (N_1737,N_1173,N_1381);
and U1738 (N_1738,N_1201,N_1413);
or U1739 (N_1739,N_1448,N_813);
or U1740 (N_1740,N_1216,N_1297);
nor U1741 (N_1741,N_1003,N_1486);
or U1742 (N_1742,N_1468,N_1410);
nor U1743 (N_1743,N_1467,N_976);
nand U1744 (N_1744,N_1228,N_764);
and U1745 (N_1745,N_1331,N_1145);
nand U1746 (N_1746,N_1404,N_1151);
and U1747 (N_1747,N_987,N_1084);
and U1748 (N_1748,N_1118,N_1484);
nor U1749 (N_1749,N_1210,N_1307);
or U1750 (N_1750,N_1027,N_1263);
nor U1751 (N_1751,N_1405,N_928);
nor U1752 (N_1752,N_1136,N_1284);
and U1753 (N_1753,N_1450,N_1345);
nand U1754 (N_1754,N_1479,N_794);
nand U1755 (N_1755,N_1462,N_1063);
nor U1756 (N_1756,N_1197,N_817);
or U1757 (N_1757,N_1009,N_781);
and U1758 (N_1758,N_1459,N_829);
and U1759 (N_1759,N_892,N_997);
nor U1760 (N_1760,N_1239,N_1237);
or U1761 (N_1761,N_1245,N_993);
nor U1762 (N_1762,N_1235,N_1227);
or U1763 (N_1763,N_1368,N_1222);
and U1764 (N_1764,N_1383,N_1353);
or U1765 (N_1765,N_947,N_818);
nand U1766 (N_1766,N_1440,N_1489);
nor U1767 (N_1767,N_853,N_1022);
nor U1768 (N_1768,N_1298,N_1076);
nor U1769 (N_1769,N_1367,N_882);
nor U1770 (N_1770,N_1161,N_1265);
nor U1771 (N_1771,N_1340,N_1267);
nor U1772 (N_1772,N_1086,N_1047);
and U1773 (N_1773,N_1422,N_1113);
nand U1774 (N_1774,N_1095,N_1485);
and U1775 (N_1775,N_1092,N_792);
nor U1776 (N_1776,N_916,N_903);
nand U1777 (N_1777,N_1283,N_1042);
and U1778 (N_1778,N_1101,N_981);
nand U1779 (N_1779,N_852,N_1474);
or U1780 (N_1780,N_1055,N_1207);
and U1781 (N_1781,N_1463,N_1071);
nand U1782 (N_1782,N_970,N_1451);
nand U1783 (N_1783,N_884,N_1060);
and U1784 (N_1784,N_1193,N_1416);
nand U1785 (N_1785,N_885,N_784);
and U1786 (N_1786,N_1070,N_778);
and U1787 (N_1787,N_1169,N_850);
nand U1788 (N_1788,N_1139,N_1258);
nand U1789 (N_1789,N_1287,N_897);
nor U1790 (N_1790,N_1080,N_823);
nor U1791 (N_1791,N_768,N_1478);
xnor U1792 (N_1792,N_1130,N_1116);
nand U1793 (N_1793,N_1336,N_1425);
nor U1794 (N_1794,N_833,N_762);
nand U1795 (N_1795,N_944,N_1180);
nor U1796 (N_1796,N_992,N_1091);
or U1797 (N_1797,N_1143,N_1114);
and U1798 (N_1798,N_1441,N_1046);
nor U1799 (N_1799,N_1223,N_1204);
and U1800 (N_1800,N_964,N_1401);
nor U1801 (N_1801,N_1318,N_1238);
and U1802 (N_1802,N_1361,N_754);
and U1803 (N_1803,N_777,N_907);
nand U1804 (N_1804,N_1006,N_1247);
nor U1805 (N_1805,N_765,N_1407);
nand U1806 (N_1806,N_783,N_1225);
or U1807 (N_1807,N_1333,N_1147);
and U1808 (N_1808,N_1252,N_979);
nor U1809 (N_1809,N_1167,N_1021);
nor U1810 (N_1810,N_828,N_982);
nor U1811 (N_1811,N_1233,N_796);
and U1812 (N_1812,N_1082,N_1149);
or U1813 (N_1813,N_900,N_1123);
or U1814 (N_1814,N_1335,N_1068);
nand U1815 (N_1815,N_945,N_906);
and U1816 (N_1816,N_943,N_1177);
and U1817 (N_1817,N_905,N_1199);
nor U1818 (N_1818,N_1488,N_904);
nand U1819 (N_1819,N_1244,N_761);
nand U1820 (N_1820,N_1453,N_770);
nor U1821 (N_1821,N_835,N_767);
or U1822 (N_1822,N_1357,N_1356);
or U1823 (N_1823,N_1202,N_825);
nand U1824 (N_1824,N_1274,N_1256);
and U1825 (N_1825,N_760,N_1475);
nor U1826 (N_1826,N_1164,N_1306);
and U1827 (N_1827,N_1019,N_1050);
or U1828 (N_1828,N_1251,N_1158);
nor U1829 (N_1829,N_1236,N_954);
nand U1830 (N_1830,N_1403,N_1038);
and U1831 (N_1831,N_1153,N_961);
or U1832 (N_1832,N_845,N_1257);
nand U1833 (N_1833,N_910,N_766);
nor U1834 (N_1834,N_1337,N_1375);
nand U1835 (N_1835,N_1221,N_1317);
or U1836 (N_1836,N_834,N_918);
and U1837 (N_1837,N_1041,N_808);
or U1838 (N_1838,N_1240,N_797);
xor U1839 (N_1839,N_1374,N_1446);
nor U1840 (N_1840,N_1062,N_1049);
and U1841 (N_1841,N_1146,N_1211);
nor U1842 (N_1842,N_844,N_1040);
and U1843 (N_1843,N_1460,N_1408);
nor U1844 (N_1844,N_1205,N_1426);
nor U1845 (N_1845,N_1387,N_1109);
nand U1846 (N_1846,N_1458,N_822);
xnor U1847 (N_1847,N_1004,N_1377);
nand U1848 (N_1848,N_1099,N_867);
and U1849 (N_1849,N_1494,N_1128);
or U1850 (N_1850,N_969,N_966);
xnor U1851 (N_1851,N_1131,N_1160);
or U1852 (N_1852,N_1077,N_782);
and U1853 (N_1853,N_1002,N_1103);
and U1854 (N_1854,N_871,N_1191);
or U1855 (N_1855,N_1117,N_1087);
nand U1856 (N_1856,N_886,N_1326);
or U1857 (N_1857,N_1088,N_1348);
nor U1858 (N_1858,N_1285,N_1476);
nand U1859 (N_1859,N_751,N_1428);
nor U1860 (N_1860,N_771,N_955);
xnor U1861 (N_1861,N_1355,N_1073);
nor U1862 (N_1862,N_827,N_1279);
or U1863 (N_1863,N_895,N_1324);
nor U1864 (N_1864,N_1064,N_802);
or U1865 (N_1865,N_1255,N_831);
or U1866 (N_1866,N_1372,N_752);
and U1867 (N_1867,N_1057,N_1295);
and U1868 (N_1868,N_1159,N_1417);
xnor U1869 (N_1869,N_839,N_1429);
or U1870 (N_1870,N_1325,N_1483);
and U1871 (N_1871,N_1078,N_806);
or U1872 (N_1872,N_1399,N_1499);
or U1873 (N_1873,N_1334,N_1010);
nand U1874 (N_1874,N_1466,N_1390);
and U1875 (N_1875,N_1150,N_1151);
and U1876 (N_1876,N_1128,N_1130);
nand U1877 (N_1877,N_1027,N_1448);
nand U1878 (N_1878,N_791,N_850);
and U1879 (N_1879,N_956,N_872);
or U1880 (N_1880,N_1237,N_1077);
or U1881 (N_1881,N_1202,N_756);
nand U1882 (N_1882,N_840,N_1303);
nor U1883 (N_1883,N_994,N_907);
nor U1884 (N_1884,N_1438,N_1442);
and U1885 (N_1885,N_937,N_1229);
nand U1886 (N_1886,N_1040,N_1276);
and U1887 (N_1887,N_1327,N_1151);
nor U1888 (N_1888,N_1138,N_1070);
and U1889 (N_1889,N_1121,N_899);
nor U1890 (N_1890,N_1390,N_1279);
or U1891 (N_1891,N_1238,N_1460);
nor U1892 (N_1892,N_1477,N_769);
nor U1893 (N_1893,N_1384,N_989);
and U1894 (N_1894,N_1454,N_944);
or U1895 (N_1895,N_879,N_885);
nor U1896 (N_1896,N_1364,N_880);
nor U1897 (N_1897,N_1243,N_1307);
nor U1898 (N_1898,N_1325,N_1413);
nand U1899 (N_1899,N_894,N_852);
or U1900 (N_1900,N_1087,N_1030);
nand U1901 (N_1901,N_792,N_845);
and U1902 (N_1902,N_1124,N_1442);
and U1903 (N_1903,N_1410,N_1219);
and U1904 (N_1904,N_1289,N_819);
or U1905 (N_1905,N_841,N_807);
nor U1906 (N_1906,N_800,N_843);
nor U1907 (N_1907,N_1489,N_1198);
and U1908 (N_1908,N_1268,N_995);
or U1909 (N_1909,N_1384,N_1297);
and U1910 (N_1910,N_1269,N_1017);
nand U1911 (N_1911,N_1387,N_1470);
nor U1912 (N_1912,N_1259,N_936);
nor U1913 (N_1913,N_1106,N_1267);
or U1914 (N_1914,N_1081,N_1137);
and U1915 (N_1915,N_853,N_968);
nor U1916 (N_1916,N_944,N_1281);
nand U1917 (N_1917,N_1297,N_1198);
and U1918 (N_1918,N_789,N_1294);
and U1919 (N_1919,N_889,N_1369);
nor U1920 (N_1920,N_1237,N_858);
nor U1921 (N_1921,N_922,N_1183);
nor U1922 (N_1922,N_1458,N_1375);
and U1923 (N_1923,N_762,N_1216);
and U1924 (N_1924,N_1373,N_779);
nor U1925 (N_1925,N_866,N_1390);
or U1926 (N_1926,N_911,N_1310);
and U1927 (N_1927,N_1395,N_913);
nand U1928 (N_1928,N_1014,N_1412);
nor U1929 (N_1929,N_979,N_1423);
or U1930 (N_1930,N_895,N_1398);
and U1931 (N_1931,N_827,N_1325);
nand U1932 (N_1932,N_920,N_1261);
nand U1933 (N_1933,N_1023,N_950);
and U1934 (N_1934,N_851,N_933);
and U1935 (N_1935,N_1050,N_795);
and U1936 (N_1936,N_865,N_1272);
xor U1937 (N_1937,N_856,N_1497);
and U1938 (N_1938,N_900,N_1397);
nand U1939 (N_1939,N_985,N_1264);
or U1940 (N_1940,N_767,N_866);
nand U1941 (N_1941,N_1435,N_1201);
and U1942 (N_1942,N_769,N_1271);
and U1943 (N_1943,N_1470,N_1251);
nor U1944 (N_1944,N_1230,N_889);
or U1945 (N_1945,N_987,N_1339);
and U1946 (N_1946,N_963,N_1205);
nand U1947 (N_1947,N_1155,N_1176);
nand U1948 (N_1948,N_843,N_1379);
nor U1949 (N_1949,N_891,N_754);
and U1950 (N_1950,N_871,N_1003);
nand U1951 (N_1951,N_1235,N_1376);
and U1952 (N_1952,N_1210,N_1265);
and U1953 (N_1953,N_928,N_1155);
and U1954 (N_1954,N_872,N_792);
nand U1955 (N_1955,N_828,N_1017);
or U1956 (N_1956,N_909,N_901);
nor U1957 (N_1957,N_816,N_987);
or U1958 (N_1958,N_795,N_1382);
nor U1959 (N_1959,N_1128,N_1470);
or U1960 (N_1960,N_1281,N_1095);
nor U1961 (N_1961,N_1412,N_1230);
nand U1962 (N_1962,N_1444,N_1283);
and U1963 (N_1963,N_1438,N_1038);
and U1964 (N_1964,N_782,N_1468);
nand U1965 (N_1965,N_1499,N_1190);
nand U1966 (N_1966,N_1169,N_1204);
or U1967 (N_1967,N_1316,N_1284);
and U1968 (N_1968,N_1301,N_909);
or U1969 (N_1969,N_1432,N_1434);
and U1970 (N_1970,N_1406,N_972);
nor U1971 (N_1971,N_982,N_790);
nor U1972 (N_1972,N_1071,N_1391);
nor U1973 (N_1973,N_973,N_791);
nand U1974 (N_1974,N_1137,N_916);
and U1975 (N_1975,N_1039,N_1034);
nor U1976 (N_1976,N_761,N_1038);
or U1977 (N_1977,N_1133,N_1483);
or U1978 (N_1978,N_1439,N_1199);
or U1979 (N_1979,N_1116,N_1330);
and U1980 (N_1980,N_889,N_1292);
nand U1981 (N_1981,N_1493,N_1299);
nand U1982 (N_1982,N_1459,N_1372);
nand U1983 (N_1983,N_795,N_988);
nor U1984 (N_1984,N_1451,N_763);
and U1985 (N_1985,N_1139,N_1225);
and U1986 (N_1986,N_1095,N_1183);
or U1987 (N_1987,N_1307,N_1449);
nand U1988 (N_1988,N_959,N_1344);
and U1989 (N_1989,N_1424,N_1354);
and U1990 (N_1990,N_1142,N_782);
and U1991 (N_1991,N_919,N_1261);
nand U1992 (N_1992,N_756,N_794);
nand U1993 (N_1993,N_1050,N_1029);
nand U1994 (N_1994,N_1063,N_1374);
and U1995 (N_1995,N_1259,N_852);
nand U1996 (N_1996,N_1282,N_1411);
xor U1997 (N_1997,N_1236,N_1270);
nand U1998 (N_1998,N_860,N_1117);
xnor U1999 (N_1999,N_870,N_766);
nor U2000 (N_2000,N_1193,N_816);
and U2001 (N_2001,N_1349,N_1029);
or U2002 (N_2002,N_1086,N_1207);
nand U2003 (N_2003,N_854,N_940);
and U2004 (N_2004,N_930,N_1186);
or U2005 (N_2005,N_1041,N_1434);
nor U2006 (N_2006,N_988,N_770);
nor U2007 (N_2007,N_1000,N_917);
nor U2008 (N_2008,N_832,N_1053);
nand U2009 (N_2009,N_1333,N_802);
or U2010 (N_2010,N_1142,N_930);
and U2011 (N_2011,N_1246,N_1495);
nor U2012 (N_2012,N_1178,N_1100);
and U2013 (N_2013,N_1449,N_1476);
nor U2014 (N_2014,N_1161,N_877);
nor U2015 (N_2015,N_1260,N_1074);
and U2016 (N_2016,N_1250,N_965);
nor U2017 (N_2017,N_914,N_1489);
nand U2018 (N_2018,N_1433,N_1224);
nor U2019 (N_2019,N_956,N_900);
nor U2020 (N_2020,N_771,N_919);
nor U2021 (N_2021,N_1158,N_882);
nor U2022 (N_2022,N_1428,N_1020);
and U2023 (N_2023,N_1278,N_1357);
or U2024 (N_2024,N_780,N_1297);
nand U2025 (N_2025,N_1134,N_1499);
nor U2026 (N_2026,N_1317,N_919);
nor U2027 (N_2027,N_781,N_1020);
and U2028 (N_2028,N_1324,N_1479);
or U2029 (N_2029,N_1372,N_763);
nand U2030 (N_2030,N_956,N_770);
nor U2031 (N_2031,N_920,N_847);
or U2032 (N_2032,N_1380,N_1383);
nor U2033 (N_2033,N_1006,N_1145);
or U2034 (N_2034,N_1309,N_1026);
and U2035 (N_2035,N_1452,N_891);
or U2036 (N_2036,N_1385,N_1199);
and U2037 (N_2037,N_987,N_795);
nand U2038 (N_2038,N_1015,N_1461);
nand U2039 (N_2039,N_1376,N_863);
and U2040 (N_2040,N_910,N_833);
nand U2041 (N_2041,N_816,N_775);
nor U2042 (N_2042,N_1442,N_925);
and U2043 (N_2043,N_1129,N_1009);
and U2044 (N_2044,N_1129,N_1469);
nor U2045 (N_2045,N_1471,N_1311);
nor U2046 (N_2046,N_1233,N_1288);
and U2047 (N_2047,N_913,N_1221);
and U2048 (N_2048,N_951,N_1314);
nor U2049 (N_2049,N_897,N_1429);
or U2050 (N_2050,N_1305,N_987);
nor U2051 (N_2051,N_1464,N_1006);
nand U2052 (N_2052,N_987,N_913);
nor U2053 (N_2053,N_935,N_1384);
nor U2054 (N_2054,N_1042,N_1035);
or U2055 (N_2055,N_990,N_1293);
or U2056 (N_2056,N_780,N_751);
nor U2057 (N_2057,N_1439,N_1457);
and U2058 (N_2058,N_884,N_1471);
or U2059 (N_2059,N_883,N_1303);
or U2060 (N_2060,N_1277,N_1226);
nor U2061 (N_2061,N_890,N_901);
nand U2062 (N_2062,N_1305,N_1075);
nand U2063 (N_2063,N_1405,N_1245);
nand U2064 (N_2064,N_870,N_1238);
or U2065 (N_2065,N_1405,N_1160);
and U2066 (N_2066,N_1229,N_779);
or U2067 (N_2067,N_945,N_858);
nand U2068 (N_2068,N_1381,N_1485);
nand U2069 (N_2069,N_1449,N_1039);
and U2070 (N_2070,N_1478,N_797);
and U2071 (N_2071,N_776,N_1156);
and U2072 (N_2072,N_771,N_1461);
and U2073 (N_2073,N_1127,N_1438);
nor U2074 (N_2074,N_1447,N_1470);
nor U2075 (N_2075,N_1120,N_1293);
nor U2076 (N_2076,N_1372,N_823);
nand U2077 (N_2077,N_909,N_1067);
nand U2078 (N_2078,N_887,N_1205);
and U2079 (N_2079,N_1111,N_1117);
and U2080 (N_2080,N_918,N_991);
nand U2081 (N_2081,N_883,N_1006);
and U2082 (N_2082,N_1363,N_1145);
nand U2083 (N_2083,N_923,N_803);
nand U2084 (N_2084,N_1488,N_1413);
nor U2085 (N_2085,N_820,N_1088);
or U2086 (N_2086,N_1134,N_1357);
nor U2087 (N_2087,N_1108,N_1310);
and U2088 (N_2088,N_839,N_972);
and U2089 (N_2089,N_782,N_834);
and U2090 (N_2090,N_835,N_1247);
nor U2091 (N_2091,N_778,N_1335);
or U2092 (N_2092,N_1308,N_1420);
and U2093 (N_2093,N_1041,N_1444);
and U2094 (N_2094,N_1266,N_1336);
nor U2095 (N_2095,N_849,N_1017);
nand U2096 (N_2096,N_1396,N_938);
nor U2097 (N_2097,N_943,N_1437);
nor U2098 (N_2098,N_929,N_1150);
nor U2099 (N_2099,N_1462,N_1459);
or U2100 (N_2100,N_1196,N_1159);
nand U2101 (N_2101,N_1131,N_1387);
nor U2102 (N_2102,N_1470,N_840);
nor U2103 (N_2103,N_1018,N_1495);
and U2104 (N_2104,N_1049,N_969);
nand U2105 (N_2105,N_1129,N_1396);
or U2106 (N_2106,N_1098,N_1022);
nor U2107 (N_2107,N_840,N_1077);
or U2108 (N_2108,N_1119,N_1321);
nand U2109 (N_2109,N_1280,N_1152);
nor U2110 (N_2110,N_1056,N_1296);
nor U2111 (N_2111,N_764,N_1280);
nor U2112 (N_2112,N_1101,N_864);
and U2113 (N_2113,N_1490,N_1271);
nor U2114 (N_2114,N_1264,N_801);
nor U2115 (N_2115,N_1177,N_1247);
or U2116 (N_2116,N_1125,N_1178);
nor U2117 (N_2117,N_1008,N_1382);
and U2118 (N_2118,N_1370,N_757);
or U2119 (N_2119,N_999,N_1005);
or U2120 (N_2120,N_1364,N_1453);
nand U2121 (N_2121,N_1282,N_1019);
or U2122 (N_2122,N_1354,N_930);
nand U2123 (N_2123,N_1442,N_1255);
nor U2124 (N_2124,N_1306,N_1200);
nor U2125 (N_2125,N_1389,N_1495);
nor U2126 (N_2126,N_1270,N_985);
and U2127 (N_2127,N_1437,N_1239);
nor U2128 (N_2128,N_1308,N_1184);
nand U2129 (N_2129,N_1488,N_1225);
nor U2130 (N_2130,N_946,N_1007);
nand U2131 (N_2131,N_955,N_1004);
nand U2132 (N_2132,N_986,N_787);
and U2133 (N_2133,N_878,N_993);
or U2134 (N_2134,N_916,N_930);
nor U2135 (N_2135,N_948,N_830);
nand U2136 (N_2136,N_759,N_898);
nor U2137 (N_2137,N_767,N_1451);
or U2138 (N_2138,N_1342,N_1105);
or U2139 (N_2139,N_817,N_1332);
or U2140 (N_2140,N_1162,N_1190);
and U2141 (N_2141,N_1227,N_927);
nor U2142 (N_2142,N_798,N_1076);
and U2143 (N_2143,N_1385,N_1061);
nand U2144 (N_2144,N_985,N_1086);
nor U2145 (N_2145,N_906,N_852);
nor U2146 (N_2146,N_894,N_1463);
and U2147 (N_2147,N_1146,N_983);
xnor U2148 (N_2148,N_1482,N_1375);
or U2149 (N_2149,N_1272,N_1033);
or U2150 (N_2150,N_1047,N_1125);
nand U2151 (N_2151,N_895,N_1200);
and U2152 (N_2152,N_1088,N_1209);
and U2153 (N_2153,N_1188,N_1220);
and U2154 (N_2154,N_1016,N_1487);
or U2155 (N_2155,N_894,N_812);
nor U2156 (N_2156,N_1384,N_1338);
or U2157 (N_2157,N_1434,N_1060);
and U2158 (N_2158,N_1168,N_1353);
nand U2159 (N_2159,N_917,N_1204);
and U2160 (N_2160,N_1368,N_1362);
nor U2161 (N_2161,N_1038,N_1175);
and U2162 (N_2162,N_907,N_967);
nor U2163 (N_2163,N_1167,N_1216);
and U2164 (N_2164,N_894,N_808);
nor U2165 (N_2165,N_806,N_1230);
or U2166 (N_2166,N_907,N_1295);
nor U2167 (N_2167,N_1146,N_1440);
nand U2168 (N_2168,N_1488,N_858);
nor U2169 (N_2169,N_946,N_829);
and U2170 (N_2170,N_813,N_959);
nor U2171 (N_2171,N_1454,N_997);
nand U2172 (N_2172,N_1340,N_1484);
or U2173 (N_2173,N_789,N_1384);
or U2174 (N_2174,N_1033,N_963);
and U2175 (N_2175,N_828,N_1121);
nand U2176 (N_2176,N_1360,N_1463);
nand U2177 (N_2177,N_1147,N_964);
nand U2178 (N_2178,N_1421,N_1031);
or U2179 (N_2179,N_1236,N_1445);
or U2180 (N_2180,N_1129,N_1065);
nor U2181 (N_2181,N_1043,N_1123);
nand U2182 (N_2182,N_1065,N_1355);
nor U2183 (N_2183,N_822,N_1151);
and U2184 (N_2184,N_1001,N_1483);
and U2185 (N_2185,N_1245,N_920);
nand U2186 (N_2186,N_1172,N_855);
nand U2187 (N_2187,N_915,N_1252);
and U2188 (N_2188,N_1216,N_859);
or U2189 (N_2189,N_1140,N_839);
xnor U2190 (N_2190,N_932,N_896);
nand U2191 (N_2191,N_977,N_965);
and U2192 (N_2192,N_1045,N_1039);
nor U2193 (N_2193,N_1096,N_778);
nor U2194 (N_2194,N_1190,N_1006);
and U2195 (N_2195,N_1340,N_862);
nor U2196 (N_2196,N_1470,N_1125);
nor U2197 (N_2197,N_1138,N_984);
and U2198 (N_2198,N_1244,N_1358);
or U2199 (N_2199,N_1328,N_1483);
nor U2200 (N_2200,N_1191,N_1096);
nor U2201 (N_2201,N_1380,N_1001);
nand U2202 (N_2202,N_1087,N_1032);
and U2203 (N_2203,N_1372,N_935);
nor U2204 (N_2204,N_1180,N_1025);
nand U2205 (N_2205,N_896,N_939);
or U2206 (N_2206,N_1017,N_1052);
nand U2207 (N_2207,N_1337,N_991);
or U2208 (N_2208,N_1098,N_897);
nand U2209 (N_2209,N_1133,N_1467);
or U2210 (N_2210,N_1393,N_1053);
or U2211 (N_2211,N_1075,N_985);
nand U2212 (N_2212,N_924,N_842);
xnor U2213 (N_2213,N_842,N_1161);
nor U2214 (N_2214,N_1302,N_876);
xnor U2215 (N_2215,N_1280,N_1392);
nand U2216 (N_2216,N_968,N_1406);
and U2217 (N_2217,N_1289,N_1067);
and U2218 (N_2218,N_839,N_876);
or U2219 (N_2219,N_1253,N_1052);
nand U2220 (N_2220,N_1420,N_1129);
nor U2221 (N_2221,N_1390,N_900);
or U2222 (N_2222,N_1305,N_770);
and U2223 (N_2223,N_1405,N_780);
nor U2224 (N_2224,N_1220,N_949);
nor U2225 (N_2225,N_1293,N_989);
and U2226 (N_2226,N_1165,N_1154);
nor U2227 (N_2227,N_1185,N_1440);
nand U2228 (N_2228,N_1055,N_1264);
nand U2229 (N_2229,N_881,N_1164);
and U2230 (N_2230,N_1347,N_1327);
nor U2231 (N_2231,N_1404,N_1075);
and U2232 (N_2232,N_1335,N_972);
nand U2233 (N_2233,N_1326,N_1323);
and U2234 (N_2234,N_1119,N_1103);
nor U2235 (N_2235,N_1155,N_1477);
nor U2236 (N_2236,N_991,N_1140);
nand U2237 (N_2237,N_1368,N_1119);
nor U2238 (N_2238,N_1077,N_848);
or U2239 (N_2239,N_1355,N_909);
nand U2240 (N_2240,N_1410,N_1097);
and U2241 (N_2241,N_1054,N_1360);
and U2242 (N_2242,N_836,N_1159);
nor U2243 (N_2243,N_942,N_1483);
or U2244 (N_2244,N_1329,N_1041);
or U2245 (N_2245,N_1493,N_820);
or U2246 (N_2246,N_1370,N_1213);
or U2247 (N_2247,N_836,N_1470);
nand U2248 (N_2248,N_871,N_1023);
and U2249 (N_2249,N_1416,N_1052);
and U2250 (N_2250,N_1789,N_1797);
or U2251 (N_2251,N_1810,N_1725);
and U2252 (N_2252,N_2236,N_1794);
or U2253 (N_2253,N_1770,N_2131);
nor U2254 (N_2254,N_2096,N_1537);
nand U2255 (N_2255,N_2081,N_1516);
nor U2256 (N_2256,N_2104,N_1556);
and U2257 (N_2257,N_1600,N_1615);
and U2258 (N_2258,N_1777,N_1680);
and U2259 (N_2259,N_1675,N_1742);
and U2260 (N_2260,N_1785,N_2125);
nand U2261 (N_2261,N_2127,N_1830);
or U2262 (N_2262,N_1930,N_1625);
and U2263 (N_2263,N_2205,N_1584);
or U2264 (N_2264,N_1567,N_1987);
nor U2265 (N_2265,N_2100,N_1821);
nor U2266 (N_2266,N_1815,N_1583);
nor U2267 (N_2267,N_1791,N_1884);
nor U2268 (N_2268,N_1866,N_2213);
nand U2269 (N_2269,N_1984,N_2012);
nor U2270 (N_2270,N_1874,N_2050);
and U2271 (N_2271,N_1698,N_2141);
nor U2272 (N_2272,N_1569,N_2024);
nor U2273 (N_2273,N_1669,N_1842);
nor U2274 (N_2274,N_2217,N_1934);
nand U2275 (N_2275,N_1761,N_2069);
or U2276 (N_2276,N_1955,N_1504);
or U2277 (N_2277,N_1767,N_1599);
nor U2278 (N_2278,N_2110,N_2044);
nor U2279 (N_2279,N_2155,N_1948);
and U2280 (N_2280,N_1817,N_2116);
nand U2281 (N_2281,N_1641,N_1841);
or U2282 (N_2282,N_2083,N_1697);
or U2283 (N_2283,N_1729,N_2201);
nand U2284 (N_2284,N_2071,N_1849);
nor U2285 (N_2285,N_1793,N_1885);
nand U2286 (N_2286,N_1896,N_2019);
and U2287 (N_2287,N_1564,N_1652);
or U2288 (N_2288,N_2009,N_2244);
or U2289 (N_2289,N_1524,N_2222);
or U2290 (N_2290,N_2229,N_2191);
nand U2291 (N_2291,N_1505,N_2215);
nand U2292 (N_2292,N_1883,N_1924);
nor U2293 (N_2293,N_2036,N_2247);
nor U2294 (N_2294,N_1538,N_2235);
and U2295 (N_2295,N_2159,N_2172);
and U2296 (N_2296,N_1996,N_1749);
or U2297 (N_2297,N_2147,N_1965);
or U2298 (N_2298,N_2230,N_1713);
nor U2299 (N_2299,N_1640,N_2192);
and U2300 (N_2300,N_2248,N_2175);
and U2301 (N_2301,N_1779,N_1834);
nand U2302 (N_2302,N_1756,N_1981);
or U2303 (N_2303,N_1663,N_1868);
nor U2304 (N_2304,N_1732,N_1752);
nand U2305 (N_2305,N_1637,N_1920);
nand U2306 (N_2306,N_2072,N_1977);
nor U2307 (N_2307,N_1700,N_1906);
or U2308 (N_2308,N_1903,N_1911);
nor U2309 (N_2309,N_2039,N_1501);
nand U2310 (N_2310,N_1708,N_1969);
nor U2311 (N_2311,N_1542,N_1714);
or U2312 (N_2312,N_1731,N_1835);
or U2313 (N_2313,N_1978,N_2183);
and U2314 (N_2314,N_1611,N_2207);
nor U2315 (N_2315,N_1990,N_1892);
nand U2316 (N_2316,N_1908,N_1551);
or U2317 (N_2317,N_1781,N_2087);
and U2318 (N_2318,N_1787,N_1730);
xnor U2319 (N_2319,N_1786,N_1531);
nand U2320 (N_2320,N_2045,N_1737);
or U2321 (N_2321,N_2057,N_2090);
nor U2322 (N_2322,N_2173,N_1851);
or U2323 (N_2323,N_1701,N_1915);
or U2324 (N_2324,N_1607,N_1719);
nand U2325 (N_2325,N_2133,N_1783);
nor U2326 (N_2326,N_1704,N_1820);
nand U2327 (N_2327,N_1929,N_1862);
or U2328 (N_2328,N_1836,N_1964);
nand U2329 (N_2329,N_1968,N_2170);
or U2330 (N_2330,N_1947,N_1557);
or U2331 (N_2331,N_1630,N_1943);
and U2332 (N_2332,N_1746,N_1959);
nand U2333 (N_2333,N_2000,N_1852);
or U2334 (N_2334,N_2187,N_1799);
xnor U2335 (N_2335,N_1559,N_2035);
nand U2336 (N_2336,N_1613,N_1644);
or U2337 (N_2337,N_2149,N_1878);
and U2338 (N_2338,N_2026,N_2243);
nand U2339 (N_2339,N_1952,N_2067);
or U2340 (N_2340,N_1921,N_2181);
or U2341 (N_2341,N_1745,N_1638);
nor U2342 (N_2342,N_2140,N_2156);
and U2343 (N_2343,N_1932,N_2017);
nand U2344 (N_2344,N_2003,N_1664);
nor U2345 (N_2345,N_1662,N_1762);
nor U2346 (N_2346,N_1586,N_2239);
and U2347 (N_2347,N_1561,N_1869);
or U2348 (N_2348,N_1806,N_1782);
nor U2349 (N_2349,N_2169,N_1945);
nand U2350 (N_2350,N_2080,N_1660);
nand U2351 (N_2351,N_1598,N_1506);
or U2352 (N_2352,N_1811,N_2008);
nor U2353 (N_2353,N_1617,N_2129);
or U2354 (N_2354,N_1950,N_1974);
and U2355 (N_2355,N_1728,N_1620);
and U2356 (N_2356,N_1667,N_2063);
and U2357 (N_2357,N_2148,N_2073);
nand U2358 (N_2358,N_1658,N_2174);
nor U2359 (N_2359,N_1527,N_2178);
nand U2360 (N_2360,N_2006,N_1876);
nand U2361 (N_2361,N_1766,N_2053);
nand U2362 (N_2362,N_2124,N_2059);
or U2363 (N_2363,N_1650,N_1857);
nand U2364 (N_2364,N_1925,N_1606);
nand U2365 (N_2365,N_2228,N_1702);
nand U2366 (N_2366,N_1734,N_1580);
nor U2367 (N_2367,N_2227,N_2091);
nor U2368 (N_2368,N_1988,N_1688);
and U2369 (N_2369,N_1741,N_2190);
nand U2370 (N_2370,N_2219,N_1631);
and U2371 (N_2371,N_1998,N_1581);
and U2372 (N_2372,N_1818,N_1848);
nor U2373 (N_2373,N_2068,N_1525);
nand U2374 (N_2374,N_2233,N_2030);
nand U2375 (N_2375,N_2011,N_1696);
nand U2376 (N_2376,N_1999,N_1859);
and U2377 (N_2377,N_2203,N_1914);
or U2378 (N_2378,N_2023,N_1944);
and U2379 (N_2379,N_1991,N_1568);
and U2380 (N_2380,N_2077,N_1622);
or U2381 (N_2381,N_2075,N_1926);
nor U2382 (N_2382,N_1519,N_1691);
and U2383 (N_2383,N_2218,N_1554);
or U2384 (N_2384,N_1587,N_1532);
nand U2385 (N_2385,N_1512,N_1758);
and U2386 (N_2386,N_2048,N_1549);
and U2387 (N_2387,N_2062,N_2216);
and U2388 (N_2388,N_1648,N_1877);
or U2389 (N_2389,N_1970,N_2226);
nand U2390 (N_2390,N_1595,N_1526);
and U2391 (N_2391,N_1686,N_2056);
or U2392 (N_2392,N_2099,N_1910);
nor U2393 (N_2393,N_2074,N_1891);
nor U2394 (N_2394,N_1623,N_1861);
nor U2395 (N_2395,N_1951,N_2220);
or U2396 (N_2396,N_2095,N_1536);
nor U2397 (N_2397,N_2113,N_1735);
nand U2398 (N_2398,N_2088,N_1529);
nor U2399 (N_2399,N_1773,N_2002);
nand U2400 (N_2400,N_1689,N_2163);
nand U2401 (N_2401,N_1986,N_1935);
or U2402 (N_2402,N_1802,N_1796);
and U2403 (N_2403,N_2001,N_1983);
and U2404 (N_2404,N_1601,N_1575);
or U2405 (N_2405,N_1853,N_1961);
nand U2406 (N_2406,N_1604,N_2241);
nor U2407 (N_2407,N_2120,N_1979);
or U2408 (N_2408,N_2033,N_2043);
and U2409 (N_2409,N_1808,N_2112);
or U2410 (N_2410,N_2094,N_1733);
or U2411 (N_2411,N_1678,N_2122);
nand U2412 (N_2412,N_1517,N_1744);
nand U2413 (N_2413,N_1850,N_1508);
and U2414 (N_2414,N_1743,N_2029);
or U2415 (N_2415,N_2168,N_2028);
and U2416 (N_2416,N_1739,N_1681);
nor U2417 (N_2417,N_2079,N_2142);
and U2418 (N_2418,N_1798,N_1975);
or U2419 (N_2419,N_1748,N_1847);
or U2420 (N_2420,N_1940,N_1997);
nand U2421 (N_2421,N_1923,N_1657);
or U2422 (N_2422,N_1543,N_1901);
nor U2423 (N_2423,N_2200,N_1594);
xnor U2424 (N_2424,N_1795,N_2164);
nand U2425 (N_2425,N_1771,N_2143);
nor U2426 (N_2426,N_1579,N_2249);
nand U2427 (N_2427,N_2186,N_2089);
or U2428 (N_2428,N_2126,N_2013);
and U2429 (N_2429,N_2047,N_1804);
or U2430 (N_2430,N_1654,N_1668);
nor U2431 (N_2431,N_1826,N_1683);
nor U2432 (N_2432,N_1922,N_1894);
or U2433 (N_2433,N_2020,N_1539);
and U2434 (N_2434,N_1726,N_1515);
or U2435 (N_2435,N_1647,N_1672);
nand U2436 (N_2436,N_2121,N_2064);
nand U2437 (N_2437,N_2032,N_1813);
and U2438 (N_2438,N_1502,N_2018);
nor U2439 (N_2439,N_1995,N_2225);
and U2440 (N_2440,N_1775,N_1710);
and U2441 (N_2441,N_2234,N_1546);
nor U2442 (N_2442,N_2197,N_1812);
nor U2443 (N_2443,N_2037,N_2237);
nand U2444 (N_2444,N_2211,N_2195);
nand U2445 (N_2445,N_1570,N_2042);
or U2446 (N_2446,N_1816,N_2139);
and U2447 (N_2447,N_1865,N_2171);
nand U2448 (N_2448,N_1778,N_1880);
or U2449 (N_2449,N_1838,N_2005);
nand U2450 (N_2450,N_1819,N_2084);
nor U2451 (N_2451,N_2108,N_1592);
nand U2452 (N_2452,N_1518,N_1521);
or U2453 (N_2453,N_1905,N_1523);
and U2454 (N_2454,N_1723,N_1715);
or U2455 (N_2455,N_1692,N_1938);
or U2456 (N_2456,N_2117,N_1629);
nor U2457 (N_2457,N_1655,N_1687);
nor U2458 (N_2458,N_1917,N_1801);
or U2459 (N_2459,N_1541,N_1928);
nor U2460 (N_2460,N_1949,N_1674);
and U2461 (N_2461,N_1954,N_1858);
nand U2462 (N_2462,N_2021,N_1937);
nor U2463 (N_2463,N_1608,N_1585);
and U2464 (N_2464,N_1670,N_2136);
nor U2465 (N_2465,N_1738,N_1957);
and U2466 (N_2466,N_1563,N_2086);
and U2467 (N_2467,N_1833,N_1677);
nand U2468 (N_2468,N_1552,N_1854);
or U2469 (N_2469,N_1912,N_1636);
nand U2470 (N_2470,N_1602,N_2109);
nor U2471 (N_2471,N_1902,N_1511);
nor U2472 (N_2472,N_1706,N_2180);
nand U2473 (N_2473,N_1718,N_1916);
or U2474 (N_2474,N_1814,N_1863);
or U2475 (N_2475,N_1768,N_1510);
and U2476 (N_2476,N_1805,N_2097);
nor U2477 (N_2477,N_1942,N_1673);
and U2478 (N_2478,N_1596,N_2015);
or U2479 (N_2479,N_2154,N_1900);
nand U2480 (N_2480,N_1591,N_1875);
and U2481 (N_2481,N_1764,N_1870);
nor U2482 (N_2482,N_2105,N_2016);
nand U2483 (N_2483,N_1985,N_2041);
nor U2484 (N_2484,N_2223,N_1717);
nor U2485 (N_2485,N_2093,N_1824);
nand U2486 (N_2486,N_1776,N_2092);
and U2487 (N_2487,N_1962,N_2199);
and U2488 (N_2488,N_1774,N_2027);
nand U2489 (N_2489,N_2052,N_2014);
and U2490 (N_2490,N_1844,N_2060);
or U2491 (N_2491,N_2066,N_1720);
and U2492 (N_2492,N_2137,N_1973);
nor U2493 (N_2493,N_2161,N_2204);
and U2494 (N_2494,N_2128,N_1571);
or U2495 (N_2495,N_1839,N_1855);
or U2496 (N_2496,N_2138,N_2007);
or U2497 (N_2497,N_1904,N_1809);
nor U2498 (N_2498,N_1618,N_2206);
and U2499 (N_2499,N_1966,N_2040);
nor U2500 (N_2500,N_1769,N_2132);
nand U2501 (N_2501,N_2103,N_2070);
nor U2502 (N_2502,N_2182,N_1772);
or U2503 (N_2503,N_2179,N_1649);
nand U2504 (N_2504,N_1831,N_1867);
nor U2505 (N_2505,N_2176,N_1871);
nor U2506 (N_2506,N_1893,N_1825);
or U2507 (N_2507,N_1760,N_1548);
nand U2508 (N_2508,N_1695,N_1513);
or U2509 (N_2509,N_1560,N_1707);
and U2510 (N_2510,N_1822,N_1864);
nand U2511 (N_2511,N_1890,N_1643);
nor U2512 (N_2512,N_2145,N_1624);
nand U2513 (N_2513,N_2058,N_1633);
or U2514 (N_2514,N_1530,N_2221);
nand U2515 (N_2515,N_2065,N_1544);
and U2516 (N_2516,N_1588,N_1879);
nand U2517 (N_2517,N_2146,N_1872);
and U2518 (N_2518,N_1562,N_2051);
and U2519 (N_2519,N_1653,N_1888);
nand U2520 (N_2520,N_1763,N_1898);
nor U2521 (N_2521,N_1566,N_1682);
nor U2522 (N_2522,N_1656,N_2167);
and U2523 (N_2523,N_2038,N_1590);
nor U2524 (N_2524,N_1646,N_1547);
and U2525 (N_2525,N_1626,N_1693);
or U2526 (N_2526,N_2022,N_2153);
or U2527 (N_2527,N_1757,N_1753);
nand U2528 (N_2528,N_1823,N_1972);
nand U2529 (N_2529,N_1666,N_1659);
nand U2530 (N_2530,N_1573,N_1642);
nor U2531 (N_2531,N_1558,N_2158);
or U2532 (N_2532,N_1895,N_2198);
nor U2533 (N_2533,N_1989,N_1711);
or U2534 (N_2534,N_1887,N_1827);
or U2535 (N_2535,N_1933,N_1605);
nand U2536 (N_2536,N_1829,N_1555);
nor U2537 (N_2537,N_1840,N_1553);
or U2538 (N_2538,N_1679,N_2188);
nor U2539 (N_2539,N_2189,N_1982);
or U2540 (N_2540,N_2135,N_2246);
and U2541 (N_2541,N_1792,N_1740);
and U2542 (N_2542,N_2130,N_1703);
and U2543 (N_2543,N_1994,N_1754);
xnor U2544 (N_2544,N_2004,N_1780);
and U2545 (N_2545,N_1759,N_1828);
or U2546 (N_2546,N_2185,N_1832);
and U2547 (N_2547,N_2123,N_1676);
or U2548 (N_2548,N_2055,N_1665);
or U2549 (N_2549,N_1939,N_1572);
or U2550 (N_2550,N_2160,N_1993);
or U2551 (N_2551,N_2098,N_1671);
nand U2552 (N_2552,N_2118,N_1927);
nor U2553 (N_2553,N_2076,N_1705);
nand U2554 (N_2554,N_2152,N_1550);
and U2555 (N_2555,N_2101,N_1958);
nor U2556 (N_2556,N_1634,N_1722);
or U2557 (N_2557,N_1627,N_1784);
nand U2558 (N_2558,N_1509,N_1919);
nand U2559 (N_2559,N_1540,N_1632);
nor U2560 (N_2560,N_1661,N_1712);
and U2561 (N_2561,N_2119,N_1520);
or U2562 (N_2562,N_1528,N_1960);
and U2563 (N_2563,N_1619,N_2102);
or U2564 (N_2564,N_2196,N_2157);
and U2565 (N_2565,N_2049,N_1582);
nor U2566 (N_2566,N_1845,N_1727);
or U2567 (N_2567,N_1918,N_1612);
nor U2568 (N_2568,N_2061,N_2245);
nor U2569 (N_2569,N_2114,N_1574);
or U2570 (N_2570,N_2082,N_1503);
nand U2571 (N_2571,N_2214,N_1533);
and U2572 (N_2572,N_1716,N_1946);
and U2573 (N_2573,N_2078,N_1507);
or U2574 (N_2574,N_1765,N_2242);
nor U2575 (N_2575,N_1931,N_1699);
nor U2576 (N_2576,N_1628,N_2232);
nor U2577 (N_2577,N_1614,N_1803);
or U2578 (N_2578,N_1976,N_2054);
nor U2579 (N_2579,N_1565,N_2224);
nor U2580 (N_2580,N_2165,N_1881);
nor U2581 (N_2581,N_2194,N_2010);
or U2582 (N_2582,N_1788,N_1721);
and U2583 (N_2583,N_1639,N_1936);
nor U2584 (N_2584,N_2208,N_1807);
or U2585 (N_2585,N_1800,N_1963);
or U2586 (N_2586,N_1747,N_1651);
nand U2587 (N_2587,N_2151,N_2046);
or U2588 (N_2588,N_2240,N_1755);
and U2589 (N_2589,N_1843,N_1621);
or U2590 (N_2590,N_2107,N_1897);
or U2591 (N_2591,N_1616,N_2238);
or U2592 (N_2592,N_2150,N_2025);
and U2593 (N_2593,N_1685,N_1593);
nor U2594 (N_2594,N_1909,N_1750);
or U2595 (N_2595,N_1522,N_1577);
and U2596 (N_2596,N_1992,N_2111);
nand U2597 (N_2597,N_1576,N_2162);
nor U2598 (N_2598,N_1500,N_1790);
or U2599 (N_2599,N_2209,N_2134);
nor U2600 (N_2600,N_1736,N_1535);
or U2601 (N_2601,N_2231,N_1956);
or U2602 (N_2602,N_2210,N_1941);
and U2603 (N_2603,N_1837,N_2115);
nand U2604 (N_2604,N_1967,N_2144);
nor U2605 (N_2605,N_1597,N_1907);
or U2606 (N_2606,N_1886,N_1860);
nand U2607 (N_2607,N_1578,N_2166);
or U2608 (N_2608,N_1684,N_1751);
nor U2609 (N_2609,N_1709,N_1694);
or U2610 (N_2610,N_1610,N_2085);
nand U2611 (N_2611,N_1645,N_1856);
nand U2612 (N_2612,N_1589,N_1899);
and U2613 (N_2613,N_2184,N_1980);
nand U2614 (N_2614,N_2177,N_1514);
nor U2615 (N_2615,N_1846,N_1953);
nand U2616 (N_2616,N_2212,N_1635);
nor U2617 (N_2617,N_1873,N_1724);
and U2618 (N_2618,N_2193,N_2202);
nor U2619 (N_2619,N_1889,N_1690);
nand U2620 (N_2620,N_1882,N_1545);
nor U2621 (N_2621,N_2106,N_2034);
xor U2622 (N_2622,N_1603,N_1913);
and U2623 (N_2623,N_1534,N_2031);
nand U2624 (N_2624,N_1971,N_1609);
and U2625 (N_2625,N_1991,N_1841);
nand U2626 (N_2626,N_1519,N_1534);
nor U2627 (N_2627,N_2064,N_1915);
and U2628 (N_2628,N_1920,N_2130);
nor U2629 (N_2629,N_1532,N_2168);
and U2630 (N_2630,N_1664,N_2065);
and U2631 (N_2631,N_2153,N_2170);
and U2632 (N_2632,N_1990,N_2185);
or U2633 (N_2633,N_1915,N_2234);
nor U2634 (N_2634,N_1521,N_2183);
and U2635 (N_2635,N_2168,N_1681);
nand U2636 (N_2636,N_1657,N_2093);
nor U2637 (N_2637,N_2089,N_2005);
and U2638 (N_2638,N_2146,N_2202);
or U2639 (N_2639,N_2084,N_1583);
and U2640 (N_2640,N_2108,N_1807);
and U2641 (N_2641,N_1914,N_2093);
and U2642 (N_2642,N_1976,N_2148);
nor U2643 (N_2643,N_1670,N_1605);
or U2644 (N_2644,N_2193,N_1908);
and U2645 (N_2645,N_2014,N_1834);
nand U2646 (N_2646,N_2203,N_1692);
nor U2647 (N_2647,N_1974,N_1849);
and U2648 (N_2648,N_2224,N_1883);
nand U2649 (N_2649,N_2076,N_1843);
and U2650 (N_2650,N_1971,N_1847);
nand U2651 (N_2651,N_1505,N_1851);
or U2652 (N_2652,N_2153,N_2047);
and U2653 (N_2653,N_1787,N_1744);
nor U2654 (N_2654,N_1982,N_1949);
and U2655 (N_2655,N_2139,N_1689);
or U2656 (N_2656,N_2177,N_1912);
or U2657 (N_2657,N_1877,N_1974);
and U2658 (N_2658,N_2229,N_2125);
nand U2659 (N_2659,N_1671,N_1537);
nand U2660 (N_2660,N_1501,N_1899);
nor U2661 (N_2661,N_1884,N_1923);
nand U2662 (N_2662,N_2018,N_2031);
and U2663 (N_2663,N_2068,N_1806);
and U2664 (N_2664,N_1930,N_1566);
and U2665 (N_2665,N_2133,N_1592);
nor U2666 (N_2666,N_1951,N_1592);
nor U2667 (N_2667,N_2101,N_2010);
and U2668 (N_2668,N_2206,N_1602);
or U2669 (N_2669,N_2170,N_2179);
nor U2670 (N_2670,N_1526,N_1592);
nor U2671 (N_2671,N_1858,N_1510);
or U2672 (N_2672,N_1706,N_1702);
or U2673 (N_2673,N_1714,N_1813);
nand U2674 (N_2674,N_2113,N_1987);
nand U2675 (N_2675,N_2210,N_2104);
or U2676 (N_2676,N_1755,N_2123);
and U2677 (N_2677,N_1673,N_2172);
nor U2678 (N_2678,N_1845,N_1865);
and U2679 (N_2679,N_2021,N_1918);
or U2680 (N_2680,N_1752,N_2132);
nor U2681 (N_2681,N_2183,N_1930);
nand U2682 (N_2682,N_1987,N_2199);
nand U2683 (N_2683,N_1626,N_2046);
and U2684 (N_2684,N_2231,N_1839);
nand U2685 (N_2685,N_1698,N_1563);
nand U2686 (N_2686,N_1949,N_1596);
nor U2687 (N_2687,N_1838,N_1759);
and U2688 (N_2688,N_2222,N_1681);
and U2689 (N_2689,N_1902,N_1864);
or U2690 (N_2690,N_2233,N_1573);
or U2691 (N_2691,N_2242,N_2099);
and U2692 (N_2692,N_1939,N_1686);
or U2693 (N_2693,N_2148,N_2233);
or U2694 (N_2694,N_1567,N_1618);
nand U2695 (N_2695,N_1779,N_2220);
and U2696 (N_2696,N_2047,N_2215);
nand U2697 (N_2697,N_2029,N_1865);
and U2698 (N_2698,N_2048,N_2009);
or U2699 (N_2699,N_2201,N_1980);
nor U2700 (N_2700,N_2081,N_2135);
or U2701 (N_2701,N_1853,N_2109);
and U2702 (N_2702,N_2116,N_1904);
and U2703 (N_2703,N_1983,N_1694);
and U2704 (N_2704,N_1860,N_2202);
and U2705 (N_2705,N_1966,N_1736);
nand U2706 (N_2706,N_2113,N_2209);
xor U2707 (N_2707,N_1868,N_2087);
nand U2708 (N_2708,N_1851,N_1783);
and U2709 (N_2709,N_2172,N_2203);
and U2710 (N_2710,N_2128,N_1851);
or U2711 (N_2711,N_1875,N_1683);
nor U2712 (N_2712,N_2018,N_1801);
nand U2713 (N_2713,N_2227,N_1735);
nor U2714 (N_2714,N_1984,N_1508);
and U2715 (N_2715,N_1749,N_1957);
and U2716 (N_2716,N_1538,N_1653);
or U2717 (N_2717,N_1866,N_1715);
or U2718 (N_2718,N_1568,N_1651);
and U2719 (N_2719,N_1684,N_1711);
nor U2720 (N_2720,N_1816,N_1596);
nand U2721 (N_2721,N_2152,N_1849);
and U2722 (N_2722,N_1804,N_1811);
or U2723 (N_2723,N_1783,N_2021);
nand U2724 (N_2724,N_2024,N_2167);
xor U2725 (N_2725,N_2138,N_1577);
nor U2726 (N_2726,N_1719,N_1959);
nand U2727 (N_2727,N_2108,N_1978);
and U2728 (N_2728,N_1635,N_1731);
nand U2729 (N_2729,N_1686,N_2228);
nand U2730 (N_2730,N_1610,N_1769);
nand U2731 (N_2731,N_2227,N_2215);
and U2732 (N_2732,N_1523,N_1720);
nand U2733 (N_2733,N_2029,N_1956);
nor U2734 (N_2734,N_1877,N_1823);
and U2735 (N_2735,N_2146,N_1915);
nor U2736 (N_2736,N_2246,N_2043);
nand U2737 (N_2737,N_1720,N_1952);
or U2738 (N_2738,N_2168,N_2051);
nor U2739 (N_2739,N_2046,N_1882);
nand U2740 (N_2740,N_2246,N_1686);
or U2741 (N_2741,N_1544,N_2090);
xnor U2742 (N_2742,N_2196,N_1576);
and U2743 (N_2743,N_2234,N_1660);
and U2744 (N_2744,N_1900,N_1744);
and U2745 (N_2745,N_1955,N_2004);
nor U2746 (N_2746,N_1817,N_1512);
or U2747 (N_2747,N_1944,N_1831);
or U2748 (N_2748,N_2161,N_2221);
nand U2749 (N_2749,N_2106,N_1802);
nand U2750 (N_2750,N_1653,N_1940);
and U2751 (N_2751,N_2060,N_1556);
nor U2752 (N_2752,N_2223,N_1897);
nand U2753 (N_2753,N_2101,N_2134);
or U2754 (N_2754,N_2200,N_1742);
nand U2755 (N_2755,N_1585,N_2016);
or U2756 (N_2756,N_1670,N_2181);
nand U2757 (N_2757,N_1751,N_2126);
and U2758 (N_2758,N_1922,N_1557);
or U2759 (N_2759,N_2101,N_2169);
and U2760 (N_2760,N_1500,N_2213);
nand U2761 (N_2761,N_1668,N_1682);
nor U2762 (N_2762,N_2224,N_1518);
and U2763 (N_2763,N_1991,N_2188);
or U2764 (N_2764,N_2205,N_1925);
nor U2765 (N_2765,N_2221,N_1667);
nand U2766 (N_2766,N_2211,N_2009);
nor U2767 (N_2767,N_1836,N_1887);
and U2768 (N_2768,N_1509,N_2146);
or U2769 (N_2769,N_2199,N_1526);
nand U2770 (N_2770,N_2095,N_1598);
and U2771 (N_2771,N_1774,N_1911);
nand U2772 (N_2772,N_1663,N_2179);
or U2773 (N_2773,N_1539,N_1587);
or U2774 (N_2774,N_1602,N_1619);
and U2775 (N_2775,N_1721,N_2081);
and U2776 (N_2776,N_2192,N_2045);
and U2777 (N_2777,N_1936,N_2105);
nand U2778 (N_2778,N_1718,N_1652);
nand U2779 (N_2779,N_1714,N_2211);
and U2780 (N_2780,N_1919,N_1847);
nor U2781 (N_2781,N_2179,N_1675);
and U2782 (N_2782,N_1713,N_1693);
and U2783 (N_2783,N_1752,N_2005);
and U2784 (N_2784,N_1794,N_1657);
and U2785 (N_2785,N_1577,N_1768);
or U2786 (N_2786,N_1584,N_2076);
nand U2787 (N_2787,N_1595,N_1580);
nand U2788 (N_2788,N_1608,N_2113);
nor U2789 (N_2789,N_1796,N_1775);
or U2790 (N_2790,N_1926,N_1524);
nor U2791 (N_2791,N_2146,N_2014);
or U2792 (N_2792,N_2089,N_1680);
nand U2793 (N_2793,N_1681,N_2197);
nor U2794 (N_2794,N_2239,N_2156);
and U2795 (N_2795,N_2064,N_2219);
nand U2796 (N_2796,N_2044,N_1515);
nor U2797 (N_2797,N_1988,N_1553);
or U2798 (N_2798,N_1841,N_1881);
and U2799 (N_2799,N_2038,N_2078);
and U2800 (N_2800,N_2220,N_1848);
or U2801 (N_2801,N_2094,N_2199);
nand U2802 (N_2802,N_1575,N_2090);
nand U2803 (N_2803,N_1864,N_2136);
or U2804 (N_2804,N_1920,N_1660);
and U2805 (N_2805,N_1574,N_2038);
nor U2806 (N_2806,N_1921,N_1900);
and U2807 (N_2807,N_2237,N_1897);
and U2808 (N_2808,N_1565,N_1724);
nand U2809 (N_2809,N_1993,N_1560);
nand U2810 (N_2810,N_1946,N_2144);
or U2811 (N_2811,N_1834,N_2050);
and U2812 (N_2812,N_1810,N_2164);
nor U2813 (N_2813,N_1853,N_1515);
or U2814 (N_2814,N_1514,N_2232);
or U2815 (N_2815,N_1522,N_2044);
or U2816 (N_2816,N_1685,N_2176);
and U2817 (N_2817,N_2002,N_1619);
xor U2818 (N_2818,N_1632,N_1583);
or U2819 (N_2819,N_2241,N_1833);
and U2820 (N_2820,N_2081,N_1857);
or U2821 (N_2821,N_2075,N_2051);
and U2822 (N_2822,N_1982,N_1899);
xor U2823 (N_2823,N_1666,N_2138);
nor U2824 (N_2824,N_2220,N_1830);
nor U2825 (N_2825,N_1962,N_2084);
or U2826 (N_2826,N_2126,N_2113);
nor U2827 (N_2827,N_1689,N_2129);
and U2828 (N_2828,N_1860,N_2071);
or U2829 (N_2829,N_2054,N_1902);
nor U2830 (N_2830,N_1860,N_2067);
nor U2831 (N_2831,N_1613,N_2154);
or U2832 (N_2832,N_1905,N_2131);
nand U2833 (N_2833,N_1672,N_1775);
or U2834 (N_2834,N_1713,N_2081);
and U2835 (N_2835,N_1700,N_1560);
or U2836 (N_2836,N_1854,N_1922);
or U2837 (N_2837,N_1906,N_2130);
or U2838 (N_2838,N_2133,N_2038);
and U2839 (N_2839,N_1735,N_1655);
and U2840 (N_2840,N_1698,N_1600);
nand U2841 (N_2841,N_1644,N_1924);
and U2842 (N_2842,N_2081,N_2149);
nor U2843 (N_2843,N_1919,N_1833);
nand U2844 (N_2844,N_2083,N_2093);
or U2845 (N_2845,N_1806,N_2000);
or U2846 (N_2846,N_1999,N_2174);
nand U2847 (N_2847,N_1745,N_1549);
and U2848 (N_2848,N_2219,N_1508);
and U2849 (N_2849,N_1906,N_1664);
nor U2850 (N_2850,N_1876,N_2100);
nor U2851 (N_2851,N_2152,N_1716);
or U2852 (N_2852,N_1994,N_2221);
nor U2853 (N_2853,N_1865,N_1517);
or U2854 (N_2854,N_2179,N_1994);
nand U2855 (N_2855,N_1623,N_2100);
nor U2856 (N_2856,N_1815,N_1897);
nand U2857 (N_2857,N_2084,N_2098);
nor U2858 (N_2858,N_1844,N_1746);
and U2859 (N_2859,N_2010,N_1697);
or U2860 (N_2860,N_1947,N_1531);
nor U2861 (N_2861,N_1618,N_1739);
or U2862 (N_2862,N_1836,N_2210);
or U2863 (N_2863,N_1609,N_1972);
nor U2864 (N_2864,N_1874,N_2042);
nand U2865 (N_2865,N_1579,N_2196);
nor U2866 (N_2866,N_2181,N_2173);
or U2867 (N_2867,N_1984,N_1762);
nand U2868 (N_2868,N_1852,N_1511);
and U2869 (N_2869,N_1809,N_1817);
or U2870 (N_2870,N_2076,N_2116);
nor U2871 (N_2871,N_1967,N_1525);
nor U2872 (N_2872,N_1938,N_1678);
and U2873 (N_2873,N_2013,N_1638);
nor U2874 (N_2874,N_1584,N_2214);
nor U2875 (N_2875,N_2031,N_1637);
nand U2876 (N_2876,N_1920,N_1911);
and U2877 (N_2877,N_1580,N_1513);
and U2878 (N_2878,N_1806,N_1600);
nor U2879 (N_2879,N_1618,N_1895);
nor U2880 (N_2880,N_2028,N_1585);
or U2881 (N_2881,N_2228,N_1665);
nor U2882 (N_2882,N_2056,N_2098);
nand U2883 (N_2883,N_1661,N_1681);
nor U2884 (N_2884,N_2043,N_2134);
nand U2885 (N_2885,N_1759,N_1817);
nor U2886 (N_2886,N_2249,N_2074);
and U2887 (N_2887,N_2050,N_1897);
nand U2888 (N_2888,N_1645,N_2025);
nand U2889 (N_2889,N_1726,N_1584);
nand U2890 (N_2890,N_1833,N_1976);
nand U2891 (N_2891,N_1580,N_1899);
or U2892 (N_2892,N_1617,N_1593);
or U2893 (N_2893,N_1619,N_2205);
xnor U2894 (N_2894,N_1996,N_1693);
and U2895 (N_2895,N_1502,N_1815);
or U2896 (N_2896,N_2158,N_1884);
nor U2897 (N_2897,N_1941,N_2085);
nor U2898 (N_2898,N_1687,N_1756);
or U2899 (N_2899,N_1542,N_1804);
and U2900 (N_2900,N_1899,N_2020);
nand U2901 (N_2901,N_2171,N_1795);
nand U2902 (N_2902,N_1952,N_1597);
nand U2903 (N_2903,N_2240,N_2110);
and U2904 (N_2904,N_1724,N_1543);
or U2905 (N_2905,N_2123,N_1802);
nor U2906 (N_2906,N_2137,N_1817);
or U2907 (N_2907,N_2104,N_1791);
and U2908 (N_2908,N_2214,N_1532);
nand U2909 (N_2909,N_1536,N_1699);
or U2910 (N_2910,N_1794,N_2237);
nor U2911 (N_2911,N_1890,N_1511);
nand U2912 (N_2912,N_1689,N_2060);
nand U2913 (N_2913,N_1788,N_1948);
and U2914 (N_2914,N_1737,N_2159);
nor U2915 (N_2915,N_1713,N_1964);
nor U2916 (N_2916,N_1755,N_1941);
and U2917 (N_2917,N_1644,N_2061);
nor U2918 (N_2918,N_2076,N_1777);
nand U2919 (N_2919,N_2249,N_1652);
nand U2920 (N_2920,N_2013,N_1904);
and U2921 (N_2921,N_2114,N_1633);
or U2922 (N_2922,N_1733,N_1652);
nor U2923 (N_2923,N_1888,N_1914);
nor U2924 (N_2924,N_1647,N_2217);
or U2925 (N_2925,N_1864,N_2150);
or U2926 (N_2926,N_1926,N_1701);
or U2927 (N_2927,N_1787,N_2146);
and U2928 (N_2928,N_1580,N_2164);
nand U2929 (N_2929,N_1552,N_1985);
nor U2930 (N_2930,N_1582,N_1551);
nor U2931 (N_2931,N_1699,N_1640);
and U2932 (N_2932,N_1650,N_2246);
nand U2933 (N_2933,N_2228,N_1583);
and U2934 (N_2934,N_2051,N_1630);
or U2935 (N_2935,N_1868,N_1956);
and U2936 (N_2936,N_2077,N_1512);
nand U2937 (N_2937,N_2001,N_1966);
and U2938 (N_2938,N_2100,N_1537);
or U2939 (N_2939,N_1985,N_1605);
xor U2940 (N_2940,N_1690,N_2143);
or U2941 (N_2941,N_1927,N_1732);
or U2942 (N_2942,N_2241,N_1679);
nor U2943 (N_2943,N_1521,N_2169);
nor U2944 (N_2944,N_2115,N_1517);
nor U2945 (N_2945,N_1620,N_1985);
or U2946 (N_2946,N_1685,N_1895);
or U2947 (N_2947,N_1774,N_1959);
and U2948 (N_2948,N_1702,N_1793);
or U2949 (N_2949,N_2069,N_2170);
or U2950 (N_2950,N_1664,N_2156);
nand U2951 (N_2951,N_1585,N_1517);
nor U2952 (N_2952,N_1832,N_1671);
and U2953 (N_2953,N_1821,N_1528);
or U2954 (N_2954,N_1770,N_2161);
or U2955 (N_2955,N_1789,N_2213);
nor U2956 (N_2956,N_1780,N_1604);
nor U2957 (N_2957,N_1934,N_1553);
or U2958 (N_2958,N_1594,N_1570);
and U2959 (N_2959,N_1650,N_1788);
or U2960 (N_2960,N_1618,N_1944);
nor U2961 (N_2961,N_2111,N_1815);
and U2962 (N_2962,N_1725,N_2205);
nand U2963 (N_2963,N_1684,N_1517);
or U2964 (N_2964,N_2045,N_2193);
nand U2965 (N_2965,N_1826,N_1676);
and U2966 (N_2966,N_2058,N_1672);
or U2967 (N_2967,N_1502,N_1728);
nor U2968 (N_2968,N_1652,N_1984);
nand U2969 (N_2969,N_1730,N_1708);
nand U2970 (N_2970,N_1915,N_2042);
or U2971 (N_2971,N_1918,N_2010);
and U2972 (N_2972,N_1626,N_2196);
or U2973 (N_2973,N_1968,N_2190);
or U2974 (N_2974,N_1665,N_1774);
nand U2975 (N_2975,N_2210,N_2024);
nand U2976 (N_2976,N_1658,N_1918);
nand U2977 (N_2977,N_1840,N_1861);
or U2978 (N_2978,N_1705,N_1726);
nor U2979 (N_2979,N_1687,N_1589);
nor U2980 (N_2980,N_1969,N_1603);
and U2981 (N_2981,N_1837,N_1718);
nor U2982 (N_2982,N_2154,N_1809);
xnor U2983 (N_2983,N_1918,N_1671);
nor U2984 (N_2984,N_1652,N_1828);
nand U2985 (N_2985,N_1624,N_2201);
or U2986 (N_2986,N_1917,N_1991);
nor U2987 (N_2987,N_1750,N_1997);
nand U2988 (N_2988,N_1676,N_2224);
and U2989 (N_2989,N_2144,N_1989);
or U2990 (N_2990,N_2053,N_1561);
nor U2991 (N_2991,N_1898,N_1893);
and U2992 (N_2992,N_1785,N_1761);
nor U2993 (N_2993,N_1645,N_1531);
or U2994 (N_2994,N_1713,N_1772);
nand U2995 (N_2995,N_2095,N_1776);
nor U2996 (N_2996,N_1791,N_2141);
and U2997 (N_2997,N_1683,N_1929);
or U2998 (N_2998,N_2172,N_2043);
nand U2999 (N_2999,N_1988,N_2131);
or UO_0 (O_0,N_2474,N_2995);
nor UO_1 (O_1,N_2260,N_2471);
nor UO_2 (O_2,N_2849,N_2517);
nor UO_3 (O_3,N_2923,N_2468);
or UO_4 (O_4,N_2296,N_2674);
and UO_5 (O_5,N_2637,N_2342);
nand UO_6 (O_6,N_2675,N_2437);
and UO_7 (O_7,N_2405,N_2503);
and UO_8 (O_8,N_2992,N_2444);
nor UO_9 (O_9,N_2403,N_2483);
and UO_10 (O_10,N_2857,N_2854);
nor UO_11 (O_11,N_2879,N_2753);
or UO_12 (O_12,N_2427,N_2274);
nor UO_13 (O_13,N_2316,N_2608);
and UO_14 (O_14,N_2948,N_2802);
and UO_15 (O_15,N_2304,N_2903);
or UO_16 (O_16,N_2365,N_2932);
and UO_17 (O_17,N_2817,N_2385);
nor UO_18 (O_18,N_2621,N_2616);
nand UO_19 (O_19,N_2732,N_2492);
nand UO_20 (O_20,N_2839,N_2850);
nor UO_21 (O_21,N_2863,N_2988);
nand UO_22 (O_22,N_2460,N_2320);
nand UO_23 (O_23,N_2364,N_2787);
or UO_24 (O_24,N_2480,N_2630);
or UO_25 (O_25,N_2484,N_2551);
and UO_26 (O_26,N_2671,N_2540);
and UO_27 (O_27,N_2401,N_2269);
and UO_28 (O_28,N_2459,N_2314);
and UO_29 (O_29,N_2846,N_2629);
and UO_30 (O_30,N_2951,N_2821);
or UO_31 (O_31,N_2658,N_2865);
and UO_32 (O_32,N_2457,N_2346);
or UO_33 (O_33,N_2946,N_2499);
nand UO_34 (O_34,N_2772,N_2795);
nand UO_35 (O_35,N_2765,N_2742);
nand UO_36 (O_36,N_2712,N_2347);
and UO_37 (O_37,N_2598,N_2723);
nand UO_38 (O_38,N_2644,N_2507);
nor UO_39 (O_39,N_2831,N_2315);
nor UO_40 (O_40,N_2659,N_2357);
or UO_41 (O_41,N_2733,N_2895);
or UO_42 (O_42,N_2899,N_2774);
nand UO_43 (O_43,N_2613,N_2798);
and UO_44 (O_44,N_2412,N_2328);
and UO_45 (O_45,N_2703,N_2736);
and UO_46 (O_46,N_2331,N_2423);
nand UO_47 (O_47,N_2336,N_2702);
or UO_48 (O_48,N_2757,N_2958);
nand UO_49 (O_49,N_2266,N_2668);
and UO_50 (O_50,N_2633,N_2627);
nand UO_51 (O_51,N_2333,N_2987);
or UO_52 (O_52,N_2799,N_2509);
and UO_53 (O_53,N_2332,N_2717);
nand UO_54 (O_54,N_2761,N_2436);
nand UO_55 (O_55,N_2720,N_2264);
and UO_56 (O_56,N_2651,N_2268);
nand UO_57 (O_57,N_2709,N_2773);
or UO_58 (O_58,N_2543,N_2522);
nor UO_59 (O_59,N_2599,N_2491);
or UO_60 (O_60,N_2295,N_2250);
nor UO_61 (O_61,N_2511,N_2752);
nor UO_62 (O_62,N_2607,N_2931);
and UO_63 (O_63,N_2496,N_2527);
and UO_64 (O_64,N_2366,N_2575);
nand UO_65 (O_65,N_2533,N_2940);
nand UO_66 (O_66,N_2413,N_2688);
or UO_67 (O_67,N_2794,N_2411);
or UO_68 (O_68,N_2662,N_2615);
or UO_69 (O_69,N_2263,N_2327);
nand UO_70 (O_70,N_2446,N_2354);
or UO_71 (O_71,N_2494,N_2893);
nor UO_72 (O_72,N_2525,N_2420);
and UO_73 (O_73,N_2355,N_2978);
nor UO_74 (O_74,N_2467,N_2382);
nor UO_75 (O_75,N_2909,N_2583);
and UO_76 (O_76,N_2939,N_2341);
or UO_77 (O_77,N_2843,N_2469);
or UO_78 (O_78,N_2272,N_2804);
and UO_79 (O_79,N_2816,N_2323);
or UO_80 (O_80,N_2855,N_2516);
and UO_81 (O_81,N_2618,N_2737);
or UO_82 (O_82,N_2783,N_2586);
nor UO_83 (O_83,N_2495,N_2299);
or UO_84 (O_84,N_2890,N_2252);
nor UO_85 (O_85,N_2350,N_2271);
xor UO_86 (O_86,N_2445,N_2695);
nand UO_87 (O_87,N_2955,N_2421);
nand UO_88 (O_88,N_2383,N_2470);
and UO_89 (O_89,N_2253,N_2463);
or UO_90 (O_90,N_2681,N_2769);
nor UO_91 (O_91,N_2257,N_2657);
or UO_92 (O_92,N_2465,N_2766);
or UO_93 (O_93,N_2547,N_2891);
nor UO_94 (O_94,N_2718,N_2914);
nand UO_95 (O_95,N_2941,N_2661);
and UO_96 (O_96,N_2925,N_2667);
and UO_97 (O_97,N_2727,N_2970);
nor UO_98 (O_98,N_2584,N_2319);
or UO_99 (O_99,N_2882,N_2915);
and UO_100 (O_100,N_2567,N_2281);
nor UO_101 (O_101,N_2834,N_2735);
nor UO_102 (O_102,N_2707,N_2605);
or UO_103 (O_103,N_2454,N_2532);
and UO_104 (O_104,N_2763,N_2293);
and UO_105 (O_105,N_2493,N_2847);
and UO_106 (O_106,N_2399,N_2273);
and UO_107 (O_107,N_2812,N_2801);
nand UO_108 (O_108,N_2764,N_2968);
and UO_109 (O_109,N_2410,N_2409);
nor UO_110 (O_110,N_2284,N_2580);
nand UO_111 (O_111,N_2530,N_2669);
and UO_112 (O_112,N_2784,N_2868);
nand UO_113 (O_113,N_2747,N_2571);
nand UO_114 (O_114,N_2933,N_2458);
or UO_115 (O_115,N_2639,N_2472);
and UO_116 (O_116,N_2856,N_2619);
nor UO_117 (O_117,N_2654,N_2878);
nor UO_118 (O_118,N_2957,N_2603);
nor UO_119 (O_119,N_2976,N_2577);
nand UO_120 (O_120,N_2579,N_2440);
nor UO_121 (O_121,N_2339,N_2949);
nand UO_122 (O_122,N_2259,N_2901);
nor UO_123 (O_123,N_2838,N_2340);
nand UO_124 (O_124,N_2318,N_2638);
nand UO_125 (O_125,N_2415,N_2287);
nor UO_126 (O_126,N_2922,N_2835);
nor UO_127 (O_127,N_2864,N_2521);
nor UO_128 (O_128,N_2701,N_2455);
nor UO_129 (O_129,N_2672,N_2544);
or UO_130 (O_130,N_2588,N_2452);
or UO_131 (O_131,N_2373,N_2289);
nand UO_132 (O_132,N_2930,N_2476);
or UO_133 (O_133,N_2964,N_2473);
or UO_134 (O_134,N_2929,N_2792);
and UO_135 (O_135,N_2602,N_2404);
or UO_136 (O_136,N_2449,N_2279);
nand UO_137 (O_137,N_2488,N_2622);
and UO_138 (O_138,N_2387,N_2983);
or UO_139 (O_139,N_2820,N_2510);
and UO_140 (O_140,N_2528,N_2256);
or UO_141 (O_141,N_2620,N_2686);
xnor UO_142 (O_142,N_2549,N_2282);
and UO_143 (O_143,N_2617,N_2956);
or UO_144 (O_144,N_2505,N_2700);
nor UO_145 (O_145,N_2921,N_2335);
nor UO_146 (O_146,N_2568,N_2569);
and UO_147 (O_147,N_2317,N_2866);
or UO_148 (O_148,N_2466,N_2748);
nand UO_149 (O_149,N_2380,N_2744);
and UO_150 (O_150,N_2979,N_2362);
and UO_151 (O_151,N_2640,N_2937);
or UO_152 (O_152,N_2926,N_2635);
nor UO_153 (O_153,N_2881,N_2408);
and UO_154 (O_154,N_2677,N_2837);
nor UO_155 (O_155,N_2848,N_2965);
and UO_156 (O_156,N_2400,N_2612);
nand UO_157 (O_157,N_2767,N_2725);
and UO_158 (O_158,N_2745,N_2267);
or UO_159 (O_159,N_2962,N_2938);
nand UO_160 (O_160,N_2561,N_2919);
and UO_161 (O_161,N_2434,N_2345);
nor UO_162 (O_162,N_2791,N_2486);
and UO_163 (O_163,N_2352,N_2574);
or UO_164 (O_164,N_2554,N_2953);
nand UO_165 (O_165,N_2447,N_2285);
nor UO_166 (O_166,N_2653,N_2634);
nor UO_167 (O_167,N_2916,N_2971);
and UO_168 (O_168,N_2508,N_2582);
nand UO_169 (O_169,N_2601,N_2626);
and UO_170 (O_170,N_2927,N_2322);
or UO_171 (O_171,N_2425,N_2343);
nor UO_172 (O_172,N_2556,N_2872);
and UO_173 (O_173,N_2824,N_2381);
or UO_174 (O_174,N_2487,N_2704);
nand UO_175 (O_175,N_2908,N_2311);
and UO_176 (O_176,N_2984,N_2706);
or UO_177 (O_177,N_2749,N_2578);
nor UO_178 (O_178,N_2699,N_2642);
or UO_179 (O_179,N_2697,N_2515);
nand UO_180 (O_180,N_2432,N_2572);
nor UO_181 (O_181,N_2429,N_2894);
nor UO_182 (O_182,N_2565,N_2836);
and UO_183 (O_183,N_2945,N_2682);
nand UO_184 (O_184,N_2541,N_2329);
or UO_185 (O_185,N_2779,N_2553);
nand UO_186 (O_186,N_2713,N_2740);
and UO_187 (O_187,N_2889,N_2407);
nor UO_188 (O_188,N_2665,N_2858);
nand UO_189 (O_189,N_2482,N_2972);
nor UO_190 (O_190,N_2985,N_2840);
or UO_191 (O_191,N_2648,N_2952);
nor UO_192 (O_192,N_2719,N_2456);
xnor UO_193 (O_193,N_2768,N_2873);
nand UO_194 (O_194,N_2646,N_2888);
and UO_195 (O_195,N_2593,N_2523);
and UO_196 (O_196,N_2442,N_2361);
nor UO_197 (O_197,N_2524,N_2678);
and UO_198 (O_198,N_2379,N_2762);
nand UO_199 (O_199,N_2743,N_2959);
and UO_200 (O_200,N_2441,N_2845);
nand UO_201 (O_201,N_2498,N_2770);
and UO_202 (O_202,N_2632,N_2363);
or UO_203 (O_203,N_2874,N_2375);
and UO_204 (O_204,N_2396,N_2999);
nand UO_205 (O_205,N_2321,N_2394);
nand UO_206 (O_206,N_2776,N_2852);
or UO_207 (O_207,N_2711,N_2811);
or UO_208 (O_208,N_2685,N_2679);
nor UO_209 (O_209,N_2963,N_2990);
nor UO_210 (O_210,N_2832,N_2782);
and UO_211 (O_211,N_2800,N_2907);
nand UO_212 (O_212,N_2258,N_2785);
and UO_213 (O_213,N_2803,N_2687);
or UO_214 (O_214,N_2809,N_2756);
nand UO_215 (O_215,N_2722,N_2283);
nand UO_216 (O_216,N_2924,N_2928);
and UO_217 (O_217,N_2690,N_2478);
and UO_218 (O_218,N_2934,N_2594);
nand UO_219 (O_219,N_2288,N_2708);
nor UO_220 (O_220,N_2351,N_2504);
or UO_221 (O_221,N_2418,N_2301);
nor UO_222 (O_222,N_2867,N_2649);
nor UO_223 (O_223,N_2376,N_2870);
or UO_224 (O_224,N_2676,N_2606);
nand UO_225 (O_225,N_2489,N_2998);
or UO_226 (O_226,N_2975,N_2330);
nand UO_227 (O_227,N_2325,N_2771);
or UO_228 (O_228,N_2275,N_2300);
nor UO_229 (O_229,N_2666,N_2292);
or UO_230 (O_230,N_2307,N_2414);
or UO_231 (O_231,N_2477,N_2278);
and UO_232 (O_232,N_2297,N_2374);
and UO_233 (O_233,N_2973,N_2609);
nor UO_234 (O_234,N_2398,N_2673);
nor UO_235 (O_235,N_2367,N_2969);
or UO_236 (O_236,N_2625,N_2805);
nand UO_237 (O_237,N_2650,N_2819);
nor UO_238 (O_238,N_2705,N_2276);
nor UO_239 (O_239,N_2906,N_2918);
nand UO_240 (O_240,N_2859,N_2419);
nand UO_241 (O_241,N_2754,N_2841);
nor UO_242 (O_242,N_2270,N_2596);
nand UO_243 (O_243,N_2898,N_2497);
nor UO_244 (O_244,N_2291,N_2944);
and UO_245 (O_245,N_2910,N_2546);
or UO_246 (O_246,N_2833,N_2981);
and UO_247 (O_247,N_2628,N_2326);
nand UO_248 (O_248,N_2557,N_2393);
xnor UO_249 (O_249,N_2448,N_2974);
nor UO_250 (O_250,N_2728,N_2604);
or UO_251 (O_251,N_2377,N_2698);
and UO_252 (O_252,N_2537,N_2545);
and UO_253 (O_253,N_2997,N_2844);
nor UO_254 (O_254,N_2349,N_2386);
nand UO_255 (O_255,N_2851,N_2371);
and UO_256 (O_256,N_2589,N_2853);
or UO_257 (O_257,N_2684,N_2359);
nor UO_258 (O_258,N_2693,N_2828);
or UO_259 (O_259,N_2825,N_2388);
nand UO_260 (O_260,N_2729,N_2775);
and UO_261 (O_261,N_2994,N_2254);
nor UO_262 (O_262,N_2741,N_2531);
or UO_263 (O_263,N_2778,N_2306);
or UO_264 (O_264,N_2947,N_2536);
or UO_265 (O_265,N_2520,N_2875);
nand UO_266 (O_266,N_2353,N_2416);
and UO_267 (O_267,N_2392,N_2724);
nor UO_268 (O_268,N_2538,N_2822);
and UO_269 (O_269,N_2904,N_2790);
and UO_270 (O_270,N_2348,N_2739);
nand UO_271 (O_271,N_2265,N_2892);
and UO_272 (O_272,N_2464,N_2826);
and UO_273 (O_273,N_2645,N_2255);
or UO_274 (O_274,N_2815,N_2500);
nor UO_275 (O_275,N_2310,N_2670);
and UO_276 (O_276,N_2683,N_2885);
and UO_277 (O_277,N_2424,N_2566);
or UO_278 (O_278,N_2694,N_2303);
or UO_279 (O_279,N_2797,N_2786);
or UO_280 (O_280,N_2395,N_2912);
nor UO_281 (O_281,N_2871,N_2433);
nor UO_282 (O_282,N_2308,N_2623);
nor UO_283 (O_283,N_2734,N_2902);
nor UO_284 (O_284,N_2731,N_2462);
and UO_285 (O_285,N_2960,N_2636);
nand UO_286 (O_286,N_2862,N_2417);
or UO_287 (O_287,N_2542,N_2758);
and UO_288 (O_288,N_2755,N_2451);
or UO_289 (O_289,N_2810,N_2624);
or UO_290 (O_290,N_2656,N_2738);
or UO_291 (O_291,N_2896,N_2559);
nor UO_292 (O_292,N_2986,N_2806);
nor UO_293 (O_293,N_2506,N_2550);
or UO_294 (O_294,N_2548,N_2989);
nor UO_295 (O_295,N_2360,N_2600);
nor UO_296 (O_296,N_2570,N_2555);
nand UO_297 (O_297,N_2807,N_2827);
nor UO_298 (O_298,N_2534,N_2305);
nand UO_299 (O_299,N_2581,N_2818);
and UO_300 (O_300,N_2356,N_2591);
and UO_301 (O_301,N_2780,N_2880);
and UO_302 (O_302,N_2501,N_2631);
nor UO_303 (O_303,N_2760,N_2829);
or UO_304 (O_304,N_2490,N_2730);
or UO_305 (O_305,N_2344,N_2967);
nand UO_306 (O_306,N_2502,N_2647);
and UO_307 (O_307,N_2368,N_2422);
and UO_308 (O_308,N_2913,N_2935);
or UO_309 (O_309,N_2917,N_2789);
nand UO_310 (O_310,N_2313,N_2954);
nor UO_311 (O_311,N_2384,N_2298);
nand UO_312 (O_312,N_2710,N_2714);
or UO_313 (O_313,N_2750,N_2905);
or UO_314 (O_314,N_2563,N_2312);
nand UO_315 (O_315,N_2643,N_2977);
nand UO_316 (O_316,N_2652,N_2877);
nand UO_317 (O_317,N_2781,N_2309);
nor UO_318 (O_318,N_2796,N_2813);
and UO_319 (O_319,N_2860,N_2814);
nand UO_320 (O_320,N_2991,N_2660);
nor UO_321 (O_321,N_2887,N_2261);
or UO_322 (O_322,N_2996,N_2372);
nand UO_323 (O_323,N_2519,N_2982);
and UO_324 (O_324,N_2759,N_2655);
nor UO_325 (O_325,N_2830,N_2334);
xnor UO_326 (O_326,N_2716,N_2611);
nor UO_327 (O_327,N_2842,N_2680);
or UO_328 (O_328,N_2746,N_2262);
and UO_329 (O_329,N_2438,N_2426);
nand UO_330 (O_330,N_2562,N_2869);
or UO_331 (O_331,N_2560,N_2324);
or UO_332 (O_332,N_2430,N_2861);
nand UO_333 (O_333,N_2614,N_2390);
nand UO_334 (O_334,N_2479,N_2439);
or UO_335 (O_335,N_2573,N_2378);
nor UO_336 (O_336,N_2788,N_2689);
or UO_337 (O_337,N_2290,N_2513);
nand UO_338 (O_338,N_2564,N_2942);
nand UO_339 (O_339,N_2721,N_2302);
and UO_340 (O_340,N_2397,N_2993);
nor UO_341 (O_341,N_2461,N_2966);
nor UO_342 (O_342,N_2715,N_2358);
nand UO_343 (O_343,N_2453,N_2526);
and UO_344 (O_344,N_2980,N_2696);
and UO_345 (O_345,N_2692,N_2883);
or UO_346 (O_346,N_2664,N_2443);
nand UO_347 (O_347,N_2726,N_2431);
and UO_348 (O_348,N_2402,N_2389);
or UO_349 (O_349,N_2900,N_2691);
and UO_350 (O_350,N_2406,N_2777);
or UO_351 (O_351,N_2391,N_2514);
nand UO_352 (O_352,N_2277,N_2884);
nand UO_353 (O_353,N_2529,N_2369);
or UO_354 (O_354,N_2558,N_2610);
nand UO_355 (O_355,N_2485,N_2592);
or UO_356 (O_356,N_2450,N_2595);
and UO_357 (O_357,N_2518,N_2961);
and UO_358 (O_358,N_2481,N_2539);
and UO_359 (O_359,N_2251,N_2294);
or UO_360 (O_360,N_2920,N_2535);
nor UO_361 (O_361,N_2886,N_2552);
nor UO_362 (O_362,N_2808,N_2590);
and UO_363 (O_363,N_2936,N_2663);
or UO_364 (O_364,N_2950,N_2337);
or UO_365 (O_365,N_2597,N_2793);
nand UO_366 (O_366,N_2576,N_2897);
xnor UO_367 (O_367,N_2475,N_2587);
or UO_368 (O_368,N_2751,N_2943);
and UO_369 (O_369,N_2512,N_2280);
or UO_370 (O_370,N_2435,N_2911);
nand UO_371 (O_371,N_2585,N_2286);
nand UO_372 (O_372,N_2428,N_2370);
nor UO_373 (O_373,N_2641,N_2338);
or UO_374 (O_374,N_2876,N_2823);
and UO_375 (O_375,N_2543,N_2529);
nor UO_376 (O_376,N_2520,N_2425);
or UO_377 (O_377,N_2448,N_2883);
xor UO_378 (O_378,N_2880,N_2713);
nor UO_379 (O_379,N_2691,N_2831);
nor UO_380 (O_380,N_2882,N_2476);
and UO_381 (O_381,N_2411,N_2906);
nor UO_382 (O_382,N_2292,N_2714);
and UO_383 (O_383,N_2462,N_2712);
nor UO_384 (O_384,N_2950,N_2934);
nor UO_385 (O_385,N_2915,N_2331);
or UO_386 (O_386,N_2582,N_2661);
and UO_387 (O_387,N_2571,N_2613);
nor UO_388 (O_388,N_2867,N_2846);
and UO_389 (O_389,N_2762,N_2519);
or UO_390 (O_390,N_2518,N_2290);
nand UO_391 (O_391,N_2976,N_2788);
nor UO_392 (O_392,N_2989,N_2813);
xnor UO_393 (O_393,N_2296,N_2616);
or UO_394 (O_394,N_2347,N_2979);
nor UO_395 (O_395,N_2276,N_2268);
nor UO_396 (O_396,N_2797,N_2501);
or UO_397 (O_397,N_2997,N_2776);
nand UO_398 (O_398,N_2853,N_2771);
nor UO_399 (O_399,N_2689,N_2897);
or UO_400 (O_400,N_2579,N_2727);
nor UO_401 (O_401,N_2390,N_2981);
and UO_402 (O_402,N_2890,N_2971);
nor UO_403 (O_403,N_2391,N_2534);
and UO_404 (O_404,N_2383,N_2450);
nor UO_405 (O_405,N_2721,N_2753);
nand UO_406 (O_406,N_2753,N_2814);
nor UO_407 (O_407,N_2984,N_2530);
and UO_408 (O_408,N_2715,N_2640);
or UO_409 (O_409,N_2663,N_2578);
or UO_410 (O_410,N_2300,N_2701);
nand UO_411 (O_411,N_2764,N_2541);
nand UO_412 (O_412,N_2725,N_2936);
nor UO_413 (O_413,N_2804,N_2264);
nand UO_414 (O_414,N_2965,N_2661);
nand UO_415 (O_415,N_2603,N_2832);
nor UO_416 (O_416,N_2285,N_2855);
xnor UO_417 (O_417,N_2902,N_2694);
nor UO_418 (O_418,N_2679,N_2829);
or UO_419 (O_419,N_2943,N_2631);
and UO_420 (O_420,N_2390,N_2566);
or UO_421 (O_421,N_2258,N_2313);
nand UO_422 (O_422,N_2855,N_2299);
and UO_423 (O_423,N_2644,N_2514);
nor UO_424 (O_424,N_2409,N_2547);
or UO_425 (O_425,N_2289,N_2696);
or UO_426 (O_426,N_2793,N_2872);
nor UO_427 (O_427,N_2746,N_2536);
nand UO_428 (O_428,N_2730,N_2950);
nor UO_429 (O_429,N_2371,N_2323);
or UO_430 (O_430,N_2582,N_2292);
nand UO_431 (O_431,N_2308,N_2875);
or UO_432 (O_432,N_2364,N_2402);
nor UO_433 (O_433,N_2344,N_2805);
nand UO_434 (O_434,N_2850,N_2400);
and UO_435 (O_435,N_2296,N_2464);
or UO_436 (O_436,N_2803,N_2520);
or UO_437 (O_437,N_2862,N_2584);
and UO_438 (O_438,N_2276,N_2305);
nor UO_439 (O_439,N_2250,N_2325);
nor UO_440 (O_440,N_2520,N_2985);
nand UO_441 (O_441,N_2966,N_2413);
nor UO_442 (O_442,N_2653,N_2282);
or UO_443 (O_443,N_2621,N_2689);
nor UO_444 (O_444,N_2910,N_2694);
or UO_445 (O_445,N_2887,N_2597);
or UO_446 (O_446,N_2547,N_2776);
or UO_447 (O_447,N_2475,N_2979);
or UO_448 (O_448,N_2648,N_2626);
nand UO_449 (O_449,N_2789,N_2689);
nor UO_450 (O_450,N_2513,N_2331);
or UO_451 (O_451,N_2768,N_2368);
or UO_452 (O_452,N_2903,N_2664);
and UO_453 (O_453,N_2254,N_2307);
nand UO_454 (O_454,N_2373,N_2890);
and UO_455 (O_455,N_2628,N_2275);
or UO_456 (O_456,N_2752,N_2536);
nand UO_457 (O_457,N_2609,N_2443);
nor UO_458 (O_458,N_2586,N_2772);
or UO_459 (O_459,N_2444,N_2262);
or UO_460 (O_460,N_2817,N_2818);
nand UO_461 (O_461,N_2854,N_2995);
and UO_462 (O_462,N_2357,N_2862);
nor UO_463 (O_463,N_2379,N_2365);
nor UO_464 (O_464,N_2755,N_2541);
nor UO_465 (O_465,N_2699,N_2740);
nand UO_466 (O_466,N_2910,N_2941);
or UO_467 (O_467,N_2630,N_2521);
and UO_468 (O_468,N_2429,N_2969);
or UO_469 (O_469,N_2358,N_2546);
nand UO_470 (O_470,N_2657,N_2910);
nand UO_471 (O_471,N_2790,N_2330);
or UO_472 (O_472,N_2842,N_2873);
and UO_473 (O_473,N_2355,N_2708);
or UO_474 (O_474,N_2845,N_2420);
and UO_475 (O_475,N_2790,N_2736);
nand UO_476 (O_476,N_2399,N_2749);
nor UO_477 (O_477,N_2936,N_2807);
and UO_478 (O_478,N_2265,N_2627);
and UO_479 (O_479,N_2587,N_2325);
nand UO_480 (O_480,N_2380,N_2257);
nor UO_481 (O_481,N_2442,N_2343);
nand UO_482 (O_482,N_2828,N_2449);
and UO_483 (O_483,N_2868,N_2378);
or UO_484 (O_484,N_2400,N_2689);
nand UO_485 (O_485,N_2875,N_2649);
and UO_486 (O_486,N_2321,N_2616);
nand UO_487 (O_487,N_2661,N_2285);
nor UO_488 (O_488,N_2791,N_2965);
nor UO_489 (O_489,N_2977,N_2406);
nand UO_490 (O_490,N_2405,N_2942);
and UO_491 (O_491,N_2495,N_2968);
nand UO_492 (O_492,N_2901,N_2572);
and UO_493 (O_493,N_2572,N_2935);
or UO_494 (O_494,N_2795,N_2718);
and UO_495 (O_495,N_2739,N_2391);
nor UO_496 (O_496,N_2483,N_2383);
nor UO_497 (O_497,N_2314,N_2652);
nor UO_498 (O_498,N_2877,N_2991);
or UO_499 (O_499,N_2285,N_2810);
endmodule