module basic_2000_20000_2500_50_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_784,In_1894);
xnor U1 (N_1,In_1792,In_1446);
nor U2 (N_2,In_571,In_1714);
and U3 (N_3,In_269,In_1854);
nand U4 (N_4,In_673,In_1657);
nand U5 (N_5,In_517,In_1752);
nor U6 (N_6,In_1205,In_490);
or U7 (N_7,In_1443,In_1661);
nor U8 (N_8,In_1827,In_965);
xor U9 (N_9,In_75,In_1569);
nand U10 (N_10,In_1152,In_668);
nor U11 (N_11,In_913,In_1545);
nor U12 (N_12,In_581,In_1702);
xnor U13 (N_13,In_1859,In_1946);
xor U14 (N_14,In_1779,In_37);
nand U15 (N_15,In_474,In_1422);
and U16 (N_16,In_1313,In_1666);
and U17 (N_17,In_45,In_1477);
or U18 (N_18,In_1227,In_1662);
or U19 (N_19,In_1004,In_1904);
and U20 (N_20,In_24,In_1069);
and U21 (N_21,In_1271,In_1669);
nand U22 (N_22,In_1317,In_1713);
nand U23 (N_23,In_545,In_1575);
nor U24 (N_24,In_1272,In_899);
or U25 (N_25,In_276,In_1725);
nand U26 (N_26,In_1395,In_1221);
or U27 (N_27,In_1898,In_1000);
xor U28 (N_28,In_38,In_859);
and U29 (N_29,In_1439,In_1252);
and U30 (N_30,In_535,In_1745);
nand U31 (N_31,In_752,In_369);
nand U32 (N_32,In_325,In_1768);
nand U33 (N_33,In_1112,In_1959);
xnor U34 (N_34,In_1651,In_970);
xnor U35 (N_35,In_1863,In_538);
xnor U36 (N_36,In_1468,In_737);
xor U37 (N_37,In_1947,In_1249);
xnor U38 (N_38,In_124,In_1290);
or U39 (N_39,In_487,In_1675);
and U40 (N_40,In_164,In_1358);
nor U41 (N_41,In_666,In_1993);
nor U42 (N_42,In_1254,In_1698);
xnor U43 (N_43,In_1034,In_97);
and U44 (N_44,In_1777,In_1934);
nor U45 (N_45,In_1343,In_1967);
xor U46 (N_46,In_399,In_1451);
and U47 (N_47,In_1509,In_1263);
nand U48 (N_48,In_1214,In_1849);
nor U49 (N_49,In_441,In_1593);
xor U50 (N_50,In_44,In_771);
or U51 (N_51,In_198,In_1919);
or U52 (N_52,In_173,In_161);
nor U53 (N_53,In_1082,In_1708);
nor U54 (N_54,In_1453,In_1552);
or U55 (N_55,In_36,In_1250);
xor U56 (N_56,In_215,In_914);
or U57 (N_57,In_1283,In_1142);
and U58 (N_58,In_1746,In_755);
xnor U59 (N_59,In_109,In_437);
and U60 (N_60,In_1346,In_943);
or U61 (N_61,In_34,In_1874);
nand U62 (N_62,In_575,In_808);
or U63 (N_63,In_499,In_1432);
nand U64 (N_64,In_1066,In_1711);
xor U65 (N_65,In_239,In_1473);
xor U66 (N_66,In_1915,In_507);
nand U67 (N_67,In_1872,In_1398);
xor U68 (N_68,In_1327,In_937);
and U69 (N_69,In_734,In_1630);
xor U70 (N_70,In_1587,In_66);
or U71 (N_71,In_822,In_1938);
nand U72 (N_72,In_1274,In_108);
or U73 (N_73,In_703,In_1712);
or U74 (N_74,In_1354,In_159);
nand U75 (N_75,In_1411,In_142);
nor U76 (N_76,In_848,In_193);
nor U77 (N_77,In_166,In_18);
and U78 (N_78,In_1573,In_445);
nor U79 (N_79,In_527,In_971);
xnor U80 (N_80,In_1914,In_1834);
xnor U81 (N_81,In_72,In_1005);
nor U82 (N_82,In_1828,In_426);
or U83 (N_83,In_1615,In_1355);
xnor U84 (N_84,In_1780,In_1980);
or U85 (N_85,In_254,In_1731);
or U86 (N_86,In_115,In_826);
nor U87 (N_87,In_1311,In_313);
xor U88 (N_88,In_756,In_1370);
nor U89 (N_89,In_1988,In_1588);
nand U90 (N_90,In_1627,In_1373);
nor U91 (N_91,In_990,In_1490);
xor U92 (N_92,In_1508,In_1018);
nand U93 (N_93,In_514,In_1030);
xor U94 (N_94,In_1016,In_864);
and U95 (N_95,In_1485,In_87);
xor U96 (N_96,In_1910,In_884);
xnor U97 (N_97,In_1644,In_422);
xnor U98 (N_98,In_1760,In_74);
or U99 (N_99,In_977,In_88);
and U100 (N_100,In_1676,In_840);
nor U101 (N_101,In_926,In_1164);
or U102 (N_102,In_1351,In_1368);
and U103 (N_103,In_1456,In_1562);
nor U104 (N_104,In_1907,In_631);
nor U105 (N_105,In_1510,In_1732);
nand U106 (N_106,In_1623,In_931);
nand U107 (N_107,In_434,In_238);
nand U108 (N_108,In_997,In_711);
or U109 (N_109,In_1330,In_641);
xor U110 (N_110,In_1624,In_1484);
or U111 (N_111,In_1554,In_1308);
or U112 (N_112,In_1457,In_1927);
xnor U113 (N_113,In_502,In_524);
and U114 (N_114,In_1171,In_488);
and U115 (N_115,In_518,In_1954);
xor U116 (N_116,In_176,In_1995);
or U117 (N_117,In_1729,In_760);
xnor U118 (N_118,In_1923,In_1469);
nand U119 (N_119,In_764,In_182);
or U120 (N_120,In_1160,In_1233);
or U121 (N_121,In_958,In_1754);
or U122 (N_122,In_1186,In_942);
xor U123 (N_123,In_119,In_1889);
xnor U124 (N_124,In_622,In_1957);
nand U125 (N_125,In_1204,In_1078);
nand U126 (N_126,In_1503,In_599);
nand U127 (N_127,In_579,In_1649);
xor U128 (N_128,In_1912,In_427);
or U129 (N_129,In_412,In_151);
or U130 (N_130,In_1495,In_1645);
nor U131 (N_131,In_68,In_1133);
nand U132 (N_132,In_1189,In_192);
nor U133 (N_133,In_334,In_744);
nand U134 (N_134,In_832,In_957);
xnor U135 (N_135,In_1803,In_1480);
xor U136 (N_136,In_69,In_1851);
nand U137 (N_137,In_1774,In_1929);
and U138 (N_138,In_1251,In_785);
and U139 (N_139,In_546,In_1117);
and U140 (N_140,In_1279,In_1818);
xor U141 (N_141,In_263,In_1149);
nor U142 (N_142,In_359,In_1790);
or U143 (N_143,In_1942,In_972);
and U144 (N_144,In_1194,In_1693);
nor U145 (N_145,In_681,In_1841);
or U146 (N_146,In_1656,In_1177);
and U147 (N_147,In_850,In_1951);
nor U148 (N_148,In_1408,In_1344);
or U149 (N_149,In_1489,In_1933);
and U150 (N_150,In_948,In_510);
nor U151 (N_151,In_1040,In_844);
xor U152 (N_152,In_1839,In_1688);
or U153 (N_153,In_1709,In_1414);
xor U154 (N_154,In_1917,In_758);
and U155 (N_155,In_1155,In_1478);
nand U156 (N_156,In_190,In_504);
xor U157 (N_157,In_939,In_1950);
xnor U158 (N_158,In_647,In_1814);
and U159 (N_159,In_1217,In_255);
xnor U160 (N_160,In_241,In_1629);
and U161 (N_161,In_1310,In_1643);
nor U162 (N_162,In_1418,In_1945);
nor U163 (N_163,In_409,In_978);
nand U164 (N_164,In_1442,In_1222);
or U165 (N_165,In_878,In_1539);
and U166 (N_166,In_1870,In_1765);
and U167 (N_167,In_341,In_1288);
or U168 (N_168,In_339,In_169);
and U169 (N_169,In_51,In_836);
or U170 (N_170,In_418,In_178);
and U171 (N_171,In_916,In_1819);
or U172 (N_172,In_640,In_739);
or U173 (N_173,In_1707,In_1493);
and U174 (N_174,In_491,In_573);
or U175 (N_175,In_905,In_944);
xor U176 (N_176,In_1369,In_408);
nor U177 (N_177,In_962,In_1976);
nor U178 (N_178,In_457,In_559);
nor U179 (N_179,In_251,In_1206);
nor U180 (N_180,In_649,In_479);
xnor U181 (N_181,In_245,In_104);
or U182 (N_182,In_1329,In_1810);
and U183 (N_183,In_1599,In_308);
or U184 (N_184,In_345,In_1331);
or U185 (N_185,In_894,In_588);
nor U186 (N_186,In_740,In_478);
nand U187 (N_187,In_250,In_383);
and U188 (N_188,In_1043,In_446);
or U189 (N_189,In_876,In_378);
and U190 (N_190,In_1039,In_1060);
nand U191 (N_191,In_1120,In_1672);
xor U192 (N_192,In_317,In_1055);
nor U193 (N_193,In_442,In_904);
xnor U194 (N_194,In_1958,In_1011);
nor U195 (N_195,In_1519,In_6);
xnor U196 (N_196,In_783,In_974);
or U197 (N_197,In_521,In_1491);
and U198 (N_198,In_1211,In_390);
and U199 (N_199,In_1876,In_342);
xnor U200 (N_200,In_805,In_1797);
or U201 (N_201,In_854,In_1476);
and U202 (N_202,In_1108,In_469);
or U203 (N_203,In_560,In_1234);
xnor U204 (N_204,In_881,In_1014);
nand U205 (N_205,In_654,In_1045);
xnor U206 (N_206,In_697,In_1423);
or U207 (N_207,In_168,In_1883);
or U208 (N_208,In_472,In_1538);
or U209 (N_209,In_304,In_1377);
nand U210 (N_210,In_1800,In_580);
nand U211 (N_211,In_122,In_574);
or U212 (N_212,In_1523,In_1739);
and U213 (N_213,In_1613,In_602);
and U214 (N_214,In_1890,In_572);
and U215 (N_215,In_1571,In_829);
xnor U216 (N_216,In_1524,In_1225);
nor U217 (N_217,In_1455,In_1505);
and U218 (N_218,In_1632,In_637);
xnor U219 (N_219,In_803,In_1660);
nor U220 (N_220,In_600,In_1444);
xnor U221 (N_221,In_410,In_564);
or U222 (N_222,In_246,In_1224);
nor U223 (N_223,In_1590,In_1148);
xnor U224 (N_224,In_1017,In_1276);
xnor U225 (N_225,In_233,In_1010);
and U226 (N_226,In_125,In_382);
nor U227 (N_227,In_1541,In_1174);
nand U228 (N_228,In_1685,In_1363);
xor U229 (N_229,In_1178,In_1259);
or U230 (N_230,In_716,In_1434);
and U231 (N_231,In_582,In_1861);
or U232 (N_232,In_1589,In_872);
xor U233 (N_233,In_1364,In_1269);
xor U234 (N_234,In_199,In_1982);
or U235 (N_235,In_1079,In_476);
or U236 (N_236,In_1740,In_583);
xor U237 (N_237,In_1273,In_295);
and U238 (N_238,In_1930,In_721);
and U239 (N_239,In_1678,In_1648);
nor U240 (N_240,In_1253,In_1032);
or U241 (N_241,In_1124,In_1500);
or U242 (N_242,In_1026,In_883);
nor U243 (N_243,In_1939,In_983);
or U244 (N_244,In_1081,In_306);
nor U245 (N_245,In_1943,In_1798);
and U246 (N_246,In_1692,In_968);
nor U247 (N_247,In_1223,In_1896);
nor U248 (N_248,In_433,In_847);
nor U249 (N_249,In_1603,In_1570);
and U250 (N_250,In_1689,In_249);
and U251 (N_251,In_1384,In_1459);
or U252 (N_252,In_1763,In_1071);
and U253 (N_253,In_1385,In_332);
nor U254 (N_254,In_117,In_1466);
or U255 (N_255,In_282,In_315);
nand U256 (N_256,In_424,In_1877);
xor U257 (N_257,In_1806,In_1412);
xor U258 (N_258,In_1846,In_354);
nor U259 (N_259,In_1061,In_1486);
xor U260 (N_260,In_1090,In_1925);
nor U261 (N_261,In_413,In_1909);
nand U262 (N_262,In_1835,In_1721);
xor U263 (N_263,In_252,In_1002);
nand U264 (N_264,In_83,In_430);
and U265 (N_265,In_61,In_67);
or U266 (N_266,In_1248,In_1144);
nor U267 (N_267,In_1670,In_1610);
nor U268 (N_268,In_1577,In_102);
or U269 (N_269,In_1462,In_1723);
or U270 (N_270,In_932,In_1056);
nor U271 (N_271,In_1507,In_1960);
or U272 (N_272,In_1918,In_1137);
nand U273 (N_273,In_1302,In_346);
and U274 (N_274,In_586,In_435);
xor U275 (N_275,In_1786,In_798);
or U276 (N_276,In_1212,In_1749);
and U277 (N_277,In_1558,In_1659);
or U278 (N_278,In_796,In_268);
nand U279 (N_279,In_635,In_1375);
or U280 (N_280,In_1246,In_40);
and U281 (N_281,In_186,In_1341);
xor U282 (N_282,In_1201,In_1403);
and U283 (N_283,In_189,In_1989);
nor U284 (N_284,In_776,In_886);
xnor U285 (N_285,In_406,In_961);
nor U286 (N_286,In_219,In_1852);
nor U287 (N_287,In_1686,In_492);
xor U288 (N_288,In_969,In_1064);
nand U289 (N_289,In_825,In_732);
and U290 (N_290,In_454,In_1862);
xor U291 (N_291,In_95,In_1682);
xnor U292 (N_292,In_674,In_947);
and U293 (N_293,In_1231,In_1084);
or U294 (N_294,In_78,In_952);
xnor U295 (N_295,In_456,In_526);
xnor U296 (N_296,In_1132,In_1262);
nand U297 (N_297,In_1544,In_28);
nor U298 (N_298,In_1949,In_256);
or U299 (N_299,In_1396,In_1447);
and U300 (N_300,In_1594,In_1126);
nor U301 (N_301,In_741,In_539);
xor U302 (N_302,In_860,In_429);
and U303 (N_303,In_16,In_1449);
or U304 (N_304,In_1609,In_395);
nand U305 (N_305,In_1481,In_696);
xnor U306 (N_306,In_1677,In_1219);
nor U307 (N_307,In_1235,In_1033);
nand U308 (N_308,In_296,In_1188);
or U309 (N_309,In_873,In_1401);
or U310 (N_310,In_209,In_222);
xnor U311 (N_311,In_1975,In_1802);
nor U312 (N_312,In_1604,In_1962);
nor U313 (N_313,In_1057,In_765);
or U314 (N_314,In_880,In_1277);
nand U315 (N_315,In_1793,In_795);
nand U316 (N_316,In_302,In_1463);
or U317 (N_317,In_237,In_235);
nor U318 (N_318,In_162,In_84);
nand U319 (N_319,In_498,In_554);
or U320 (N_320,In_903,In_845);
or U321 (N_321,In_1388,In_1345);
xor U322 (N_322,In_1049,In_1093);
and U323 (N_323,In_915,In_1866);
and U324 (N_324,In_662,In_1633);
nor U325 (N_325,In_889,In_266);
nor U326 (N_326,In_1323,In_1333);
and U327 (N_327,In_1673,In_781);
nand U328 (N_328,In_1409,In_1448);
nand U329 (N_329,In_46,In_1684);
and U330 (N_330,In_1361,In_22);
nor U331 (N_331,In_1320,In_455);
and U332 (N_332,In_1542,In_1095);
or U333 (N_333,In_1920,In_1758);
and U334 (N_334,In_1766,In_1244);
nand U335 (N_335,In_307,In_401);
nor U336 (N_336,In_793,In_870);
nor U337 (N_337,In_797,In_1769);
nand U338 (N_338,In_1022,In_0);
or U339 (N_339,In_534,In_4);
nor U340 (N_340,In_1129,In_1114);
and U341 (N_341,In_896,In_105);
xor U342 (N_342,In_415,In_1963);
nand U343 (N_343,In_1887,In_114);
or U344 (N_344,In_1035,In_1628);
or U345 (N_345,In_360,In_1);
and U346 (N_346,In_1840,In_1784);
or U347 (N_347,In_55,In_849);
and U348 (N_348,In_1292,In_1715);
and U349 (N_349,In_1727,In_1566);
xor U350 (N_350,In_1534,In_1820);
or U351 (N_351,In_516,In_1638);
or U352 (N_352,In_1621,In_389);
xnor U353 (N_353,In_642,In_1134);
and U354 (N_354,In_1671,In_1001);
nand U355 (N_355,In_675,In_1342);
or U356 (N_356,In_1421,In_39);
nand U357 (N_357,In_569,In_136);
nand U358 (N_358,In_1406,In_1051);
and U359 (N_359,In_901,In_1972);
or U360 (N_360,In_1156,In_766);
or U361 (N_361,In_265,In_1650);
nor U362 (N_362,In_1298,In_1619);
nand U363 (N_363,In_1717,In_1617);
or U364 (N_364,In_1815,In_1303);
nor U365 (N_365,In_1107,In_594);
xnor U366 (N_366,In_1441,In_1195);
xnor U367 (N_367,In_126,In_918);
and U368 (N_368,In_1256,In_495);
nand U369 (N_369,In_1668,In_1121);
and U370 (N_370,In_106,In_1305);
xor U371 (N_371,In_96,In_1119);
or U372 (N_372,In_1838,In_468);
xnor U373 (N_373,In_1762,In_1563);
xnor U374 (N_374,In_1606,In_1783);
xor U375 (N_375,In_388,In_570);
nor U376 (N_376,In_1190,In_1240);
nand U377 (N_377,In_1683,In_1172);
and U378 (N_378,In_1180,In_1937);
xnor U379 (N_379,In_869,In_693);
nor U380 (N_380,In_443,In_1220);
or U381 (N_381,In_1556,In_1536);
or U382 (N_382,In_1636,In_1759);
nor U383 (N_383,In_232,In_1878);
nand U384 (N_384,In_1102,In_1584);
or U385 (N_385,In_902,In_778);
xnor U386 (N_386,In_1183,In_328);
and U387 (N_387,In_1243,In_82);
or U388 (N_388,In_1540,In_1753);
nor U389 (N_389,In_361,In_1547);
xor U390 (N_390,In_1208,In_318);
nand U391 (N_391,In_685,In_394);
or U392 (N_392,In_1371,In_800);
xor U393 (N_393,In_1748,In_505);
and U394 (N_394,In_1150,In_698);
and U395 (N_395,In_458,In_7);
or U396 (N_396,In_595,In_1900);
nor U397 (N_397,In_1572,In_1626);
xnor U398 (N_398,In_107,In_365);
nand U399 (N_399,In_231,In_165);
nor U400 (N_400,In_1467,In_1809);
xnor U401 (N_401,In_181,In_373);
or U402 (N_402,In_1198,N_239);
xor U403 (N_403,In_1674,In_671);
and U404 (N_404,In_425,N_287);
nor U405 (N_405,In_123,In_688);
xor U406 (N_406,In_1215,In_812);
or U407 (N_407,N_183,In_858);
and U408 (N_408,In_1718,In_240);
nor U409 (N_409,N_120,In_644);
nor U410 (N_410,In_1831,N_128);
and U411 (N_411,In_1940,N_148);
nor U412 (N_412,N_180,In_1978);
or U413 (N_413,In_657,In_1013);
xor U414 (N_414,N_156,N_248);
or U415 (N_415,In_645,In_1282);
nor U416 (N_416,In_1535,In_1260);
xor U417 (N_417,In_1936,N_132);
nor U418 (N_418,In_1956,N_260);
or U419 (N_419,In_1297,N_79);
nand U420 (N_420,In_41,N_295);
xnor U421 (N_421,N_133,In_1379);
nor U422 (N_422,N_208,In_343);
xnor U423 (N_423,N_297,In_497);
nor U424 (N_424,In_720,In_1291);
nor U425 (N_425,In_1964,N_110);
xor U426 (N_426,In_911,In_1236);
and U427 (N_427,In_85,In_861);
and U428 (N_428,In_677,N_147);
nand U429 (N_429,In_1110,In_610);
or U430 (N_430,In_1533,In_320);
or U431 (N_431,N_75,N_225);
and U432 (N_432,In_484,In_473);
and U433 (N_433,In_1764,In_1365);
and U434 (N_434,N_194,In_385);
xor U435 (N_435,In_609,N_231);
and U436 (N_436,In_230,In_285);
nand U437 (N_437,In_171,N_173);
and U438 (N_438,N_368,In_52);
xnor U439 (N_439,In_1275,N_284);
and U440 (N_440,N_224,In_1559);
nand U441 (N_441,In_1823,In_172);
xor U442 (N_442,In_323,In_1230);
xnor U443 (N_443,In_1173,In_551);
nand U444 (N_444,In_1736,In_1359);
nor U445 (N_445,In_1724,N_366);
xor U446 (N_446,In_153,In_908);
xnor U447 (N_447,In_1435,In_585);
or U448 (N_448,In_985,In_818);
nor U449 (N_449,N_187,In_297);
and U450 (N_450,In_1226,N_271);
or U451 (N_451,N_115,In_1794);
xnor U452 (N_452,In_1270,In_120);
nor U453 (N_453,In_60,In_1109);
and U454 (N_454,In_1785,In_223);
nand U455 (N_455,N_360,In_493);
xnor U456 (N_456,In_992,N_320);
xnor U457 (N_457,In_481,In_863);
or U458 (N_458,N_313,In_810);
and U459 (N_459,In_1494,In_964);
nand U460 (N_460,In_111,In_589);
nor U461 (N_461,In_749,In_1911);
nor U462 (N_462,In_988,In_286);
nor U463 (N_463,N_269,In_1922);
and U464 (N_464,In_1127,In_1339);
nand U465 (N_465,In_541,In_397);
nand U466 (N_466,In_1548,In_29);
xor U467 (N_467,In_705,N_153);
or U468 (N_468,In_314,In_118);
nor U469 (N_469,N_243,In_376);
and U470 (N_470,N_95,N_362);
and U471 (N_471,N_168,In_719);
nand U472 (N_472,In_357,In_1031);
or U473 (N_473,In_1420,N_223);
xor U474 (N_474,In_1294,N_257);
or U475 (N_475,In_20,In_1077);
or U476 (N_476,In_1338,In_1687);
nor U477 (N_477,N_66,N_123);
nand U478 (N_478,N_386,In_1842);
nand U479 (N_479,In_871,In_1210);
nor U480 (N_480,In_58,N_292);
or U481 (N_481,In_823,In_1209);
nand U482 (N_482,In_1808,In_814);
xnor U483 (N_483,N_21,N_202);
xor U484 (N_484,In_540,In_1191);
or U485 (N_485,In_634,In_1869);
nand U486 (N_486,In_1832,In_757);
nor U487 (N_487,N_200,In_1580);
nor U488 (N_488,In_1238,In_1681);
nand U489 (N_489,In_1293,In_1665);
or U490 (N_490,In_1038,In_1387);
nand U491 (N_491,In_291,In_1799);
xor U492 (N_492,In_1985,N_47);
nand U493 (N_493,N_62,N_35);
nand U494 (N_494,In_566,In_1770);
or U495 (N_495,In_1928,In_761);
or U496 (N_496,In_509,In_960);
nand U497 (N_497,In_1965,In_1050);
nor U498 (N_498,In_80,In_1182);
nor U499 (N_499,In_922,In_287);
and U500 (N_500,In_350,N_290);
and U501 (N_501,In_310,In_1706);
nor U502 (N_502,In_489,N_141);
or U503 (N_503,In_1268,In_772);
xor U504 (N_504,In_1871,In_1161);
or U505 (N_505,In_391,N_10);
nand U506 (N_506,In_628,In_710);
nor U507 (N_507,In_258,In_620);
or U508 (N_508,N_55,In_206);
nand U509 (N_509,In_667,In_1436);
xnor U510 (N_510,N_116,N_186);
or U511 (N_511,N_142,In_1948);
xnor U512 (N_512,N_121,In_1897);
xor U513 (N_513,In_1848,N_279);
nand U514 (N_514,In_1882,In_694);
nor U515 (N_515,In_312,In_1097);
nand U516 (N_516,In_494,In_1926);
or U517 (N_517,In_718,In_130);
nand U518 (N_518,In_831,In_200);
nand U519 (N_519,In_191,N_355);
nand U520 (N_520,In_1529,In_1826);
nand U521 (N_521,In_1932,In_133);
nor U522 (N_522,In_1047,In_1372);
xor U523 (N_523,In_1125,N_262);
or U524 (N_524,In_333,In_1153);
nor U525 (N_525,N_264,N_44);
and U526 (N_526,In_553,N_155);
nand U527 (N_527,In_77,In_1007);
xnor U528 (N_528,In_244,In_1526);
and U529 (N_529,N_96,In_1295);
or U530 (N_530,N_294,In_788);
nor U531 (N_531,In_175,N_356);
and U532 (N_532,In_1596,In_1499);
nand U533 (N_533,In_874,In_1553);
xnor U534 (N_534,In_329,In_866);
xnor U535 (N_535,N_379,N_345);
nand U536 (N_536,In_607,In_1350);
or U537 (N_537,In_584,In_596);
xnor U538 (N_538,In_25,In_224);
or U539 (N_539,N_129,In_444);
or U540 (N_540,In_1321,In_824);
or U541 (N_541,In_738,N_164);
nor U542 (N_542,In_326,N_72);
or U543 (N_543,In_706,In_1895);
and U544 (N_544,In_780,In_381);
nand U545 (N_545,In_1139,In_837);
or U546 (N_546,In_533,In_146);
or U547 (N_547,In_459,In_1415);
xnor U548 (N_548,N_329,In_1100);
xor U549 (N_549,In_1560,In_821);
nand U550 (N_550,In_843,In_953);
nand U551 (N_551,In_658,N_321);
and U552 (N_552,In_53,In_909);
nand U553 (N_553,In_841,In_212);
xnor U554 (N_554,In_1163,In_149);
xnor U555 (N_555,N_193,N_254);
and U556 (N_556,In_1987,In_1048);
or U557 (N_557,In_1741,In_1696);
xnor U558 (N_558,In_128,In_272);
nor U559 (N_559,In_464,N_198);
and U560 (N_560,N_46,In_248);
or U561 (N_561,In_981,N_253);
or U562 (N_562,In_15,In_1374);
or U563 (N_563,In_727,N_102);
nor U564 (N_564,In_1788,N_60);
or U565 (N_565,In_1857,In_851);
nand U566 (N_566,In_14,In_157);
nor U567 (N_567,In_790,In_138);
nor U568 (N_568,N_238,In_1378);
xor U569 (N_569,In_1394,In_1192);
nand U570 (N_570,In_621,In_1053);
or U571 (N_571,N_54,In_1267);
nor U572 (N_572,In_1402,In_404);
nor U573 (N_573,In_1136,In_1105);
nand U574 (N_574,In_1537,N_242);
nor U575 (N_575,In_531,N_302);
nand U576 (N_576,N_22,N_337);
xor U577 (N_577,N_317,In_1203);
nand U578 (N_578,N_109,In_548);
nand U579 (N_579,In_664,N_378);
nand U580 (N_580,N_195,N_125);
nand U581 (N_581,N_14,In_1837);
and U582 (N_582,N_99,In_1655);
xor U583 (N_583,In_1245,In_229);
nor U584 (N_584,In_227,N_311);
or U585 (N_585,In_537,In_1722);
nor U586 (N_586,In_979,N_167);
nor U587 (N_587,N_259,N_58);
or U588 (N_588,In_271,N_163);
and U589 (N_589,N_89,In_436);
xor U590 (N_590,In_49,In_1289);
and U591 (N_591,In_733,N_252);
xnor U592 (N_592,In_611,N_373);
and U593 (N_593,In_767,In_1352);
and U594 (N_594,In_447,N_280);
or U595 (N_595,In_1482,In_565);
nand U596 (N_596,N_65,In_1347);
and U597 (N_597,In_643,N_82);
xnor U598 (N_598,In_1772,N_70);
or U599 (N_599,In_704,In_700);
or U600 (N_600,In_1543,In_1574);
or U601 (N_601,In_763,In_274);
and U602 (N_602,N_322,In_363);
nand U603 (N_603,In_1044,N_218);
or U604 (N_604,In_1737,In_57);
xnor U605 (N_605,N_370,In_1036);
nand U606 (N_606,In_1921,In_1116);
or U607 (N_607,In_725,N_392);
xor U608 (N_608,In_951,In_403);
or U609 (N_609,In_1019,In_11);
nor U610 (N_610,In_221,In_1020);
or U611 (N_611,N_363,In_1115);
nand U612 (N_612,In_103,In_8);
nand U613 (N_613,In_769,N_53);
and U614 (N_614,In_1492,N_255);
xor U615 (N_615,In_1935,N_272);
nor U616 (N_616,In_174,N_171);
or U617 (N_617,In_1634,In_1607);
and U618 (N_618,In_1075,In_787);
or U619 (N_619,In_1170,In_1845);
nand U620 (N_620,In_1996,N_2);
and U621 (N_621,N_13,In_995);
or U622 (N_622,In_1065,In_1450);
xnor U623 (N_623,N_256,N_296);
nor U624 (N_624,In_316,In_145);
xor U625 (N_625,In_1525,In_1601);
nor U626 (N_626,In_347,In_201);
nand U627 (N_627,N_209,N_235);
and U628 (N_628,In_1738,In_1280);
xor U629 (N_629,N_312,N_36);
nand U630 (N_630,In_1734,In_1701);
nand U631 (N_631,N_289,In_924);
nor U632 (N_632,In_1257,N_380);
or U633 (N_633,N_177,In_1652);
and U634 (N_634,In_1899,In_1498);
xor U635 (N_635,In_1356,In_1516);
nand U636 (N_636,In_1074,N_237);
nor U637 (N_637,In_1241,In_423);
nor U638 (N_638,N_185,In_1667);
xor U639 (N_639,In_1316,In_471);
nand U640 (N_640,N_5,In_1916);
nor U641 (N_641,In_1873,In_279);
xnor U642 (N_642,In_1501,In_888);
xnor U643 (N_643,N_276,In_1970);
xnor U644 (N_644,In_656,In_672);
nor U645 (N_645,N_340,In_1585);
nand U646 (N_646,In_967,In_152);
nand U647 (N_647,In_1154,N_318);
xnor U648 (N_648,In_1822,In_477);
nor U649 (N_649,In_1646,N_108);
and U650 (N_650,In_1389,In_1096);
nand U651 (N_651,In_1997,N_157);
nor U652 (N_652,In_1631,N_216);
xor U653 (N_653,In_242,In_1386);
nand U654 (N_654,N_367,In_1483);
xnor U655 (N_655,In_1605,In_775);
nor U656 (N_656,In_753,N_56);
nor U657 (N_657,N_240,In_1518);
and U658 (N_658,N_113,In_655);
nor U659 (N_659,N_326,In_195);
or U660 (N_660,In_1165,N_64);
nand U661 (N_661,In_416,In_300);
xor U662 (N_662,In_1567,In_567);
nor U663 (N_663,N_134,N_212);
or U664 (N_664,In_910,In_1080);
and U665 (N_665,In_1076,In_1886);
xnor U666 (N_666,In_1795,In_1118);
nor U667 (N_667,N_377,N_97);
xnor U668 (N_668,In_1561,In_742);
and U669 (N_669,N_285,In_1383);
or U670 (N_670,In_1111,N_6);
nor U671 (N_671,N_338,In_1789);
nor U672 (N_672,In_839,In_1184);
or U673 (N_673,N_357,In_1893);
nand U674 (N_674,In_1324,In_1416);
xor U675 (N_675,In_267,In_402);
nor U676 (N_676,In_1973,In_670);
xor U677 (N_677,N_389,In_1089);
nand U678 (N_678,In_353,In_506);
xor U679 (N_679,N_275,In_475);
or U680 (N_680,In_1419,N_274);
or U681 (N_681,In_1287,N_166);
and U682 (N_682,N_374,N_67);
nand U683 (N_683,In_1012,N_9);
xnor U684 (N_684,N_277,In_280);
nand U685 (N_685,In_236,In_608);
and U686 (N_686,In_1608,In_1296);
nand U687 (N_687,In_963,In_387);
and U688 (N_688,N_28,In_1318);
nor U689 (N_689,N_350,N_291);
nand U690 (N_690,In_1067,N_16);
xor U691 (N_691,In_1864,In_1602);
nand U692 (N_692,In_508,In_374);
nor U693 (N_693,In_451,In_1261);
nand U694 (N_694,In_465,In_19);
xor U695 (N_695,In_31,N_88);
nand U696 (N_696,In_1207,In_699);
nor U697 (N_697,In_460,In_70);
nor U698 (N_698,N_206,N_324);
or U699 (N_699,In_1787,In_627);
xnor U700 (N_700,In_605,In_99);
and U701 (N_701,N_170,In_259);
nand U702 (N_702,In_65,N_181);
nand U703 (N_703,In_1924,N_348);
nand U704 (N_704,In_542,N_172);
nand U705 (N_705,N_42,In_1856);
and U706 (N_706,N_263,In_1479);
nand U707 (N_707,In_1088,In_1106);
and U708 (N_708,In_748,In_1337);
nor U709 (N_709,In_1703,In_1391);
nor U710 (N_710,N_384,In_1860);
or U711 (N_711,In_1471,In_680);
and U712 (N_712,In_1564,In_598);
xor U713 (N_713,In_335,In_1122);
or U714 (N_714,N_201,In_262);
nor U715 (N_715,In_603,In_1242);
or U716 (N_716,In_439,In_1008);
and U717 (N_717,In_449,In_1694);
nand U718 (N_718,In_1858,In_877);
and U719 (N_719,In_1025,In_1782);
or U720 (N_720,In_218,In_2);
and U721 (N_721,In_71,In_1438);
xnor U722 (N_722,In_827,In_1986);
nand U723 (N_723,In_1513,In_1006);
and U724 (N_724,In_702,In_1690);
xor U725 (N_725,In_1255,In_1716);
nand U726 (N_726,N_309,In_906);
nand U727 (N_727,In_1098,In_528);
nand U728 (N_728,In_54,In_949);
xnor U729 (N_729,In_1658,In_1128);
and U730 (N_730,In_991,N_117);
and U731 (N_731,In_183,In_1647);
nand U732 (N_732,In_1974,In_180);
xnor U733 (N_733,In_337,In_1735);
nor U734 (N_734,N_314,N_393);
xor U735 (N_735,In_1470,In_194);
and U736 (N_736,In_1399,N_19);
and U737 (N_737,N_396,In_830);
or U738 (N_738,In_529,In_774);
and U739 (N_739,N_140,In_777);
xnor U740 (N_740,In_453,In_1622);
nand U741 (N_741,In_35,In_1381);
nor U742 (N_742,In_1968,In_555);
nor U743 (N_743,N_222,In_895);
or U744 (N_744,In_1833,N_395);
or U745 (N_745,In_1867,In_1232);
xor U746 (N_746,In_331,N_107);
and U747 (N_747,N_308,In_486);
and U748 (N_748,In_1578,In_1353);
nand U749 (N_749,In_1309,In_372);
nor U750 (N_750,In_646,In_1300);
nand U751 (N_751,In_751,In_1591);
nand U752 (N_752,In_299,In_264);
nand U753 (N_753,In_1218,In_419);
nand U754 (N_754,In_1094,In_801);
and U755 (N_755,N_387,In_513);
xor U756 (N_756,In_882,In_1884);
and U757 (N_757,N_353,In_1285);
xnor U758 (N_758,In_1952,In_519);
or U759 (N_759,In_660,In_1971);
nor U760 (N_760,In_597,In_1425);
and U761 (N_761,In_1009,In_420);
xnor U762 (N_762,In_1167,In_349);
and U763 (N_763,In_802,In_523);
nand U764 (N_764,In_503,In_557);
nor U765 (N_765,N_59,In_525);
nor U766 (N_766,In_928,In_1908);
xnor U767 (N_767,In_301,In_1620);
and U768 (N_768,N_301,In_587);
xnor U769 (N_769,In_1175,In_1773);
nor U770 (N_770,N_245,N_305);
xor U771 (N_771,N_349,In_1085);
nor U772 (N_772,N_335,In_1059);
nand U773 (N_773,In_799,In_701);
or U774 (N_774,N_101,In_1757);
or U775 (N_775,In_1131,In_893);
and U776 (N_776,In_515,In_1410);
nand U777 (N_777,In_205,N_52);
or U778 (N_778,In_1504,In_480);
xnor U779 (N_779,In_377,In_921);
nand U780 (N_780,In_651,In_817);
nor U781 (N_781,In_1576,In_724);
nor U782 (N_782,In_1522,In_204);
xnor U783 (N_783,In_1286,In_659);
or U784 (N_784,In_155,In_833);
nand U785 (N_785,In_1176,In_619);
nand U786 (N_786,In_1357,In_392);
nor U787 (N_787,In_163,In_1091);
or U788 (N_788,In_633,In_311);
or U789 (N_789,In_998,In_213);
nor U790 (N_790,In_220,In_154);
nand U791 (N_791,In_919,In_452);
nand U792 (N_792,N_197,In_370);
nor U793 (N_793,In_1023,In_1704);
nor U794 (N_794,In_1433,N_146);
nand U795 (N_795,In_1550,N_328);
or U796 (N_796,In_708,In_64);
or U797 (N_797,In_1557,N_247);
or U798 (N_798,N_48,N_234);
nor U799 (N_799,In_828,N_41);
xnor U800 (N_800,In_639,In_247);
nand U801 (N_801,N_652,N_408);
nor U802 (N_802,In_17,In_141);
or U803 (N_803,N_541,In_1742);
and U804 (N_804,N_680,In_1140);
or U805 (N_805,N_765,In_1728);
nand U806 (N_806,In_1159,In_1614);
xor U807 (N_807,N_658,N_472);
or U808 (N_808,N_273,In_1778);
xnor U809 (N_809,N_354,In_98);
nor U810 (N_810,N_410,N_574);
xor U811 (N_811,N_407,In_1581);
and U812 (N_812,N_478,In_994);
nand U813 (N_813,In_289,N_303);
or U814 (N_814,In_281,N_130);
nand U815 (N_815,N_174,N_697);
nand U816 (N_816,In_500,N_781);
nand U817 (N_817,N_660,In_1892);
xor U818 (N_818,In_820,In_1445);
or U819 (N_819,In_1464,In_1322);
nor U820 (N_820,N_449,N_528);
nor U821 (N_821,N_706,N_669);
and U822 (N_822,N_647,In_616);
and U823 (N_823,In_636,N_634);
or U824 (N_824,In_482,In_1196);
and U825 (N_825,N_798,In_1239);
nor U826 (N_826,N_152,In_687);
nand U827 (N_827,In_638,In_440);
nor U828 (N_828,In_1512,N_330);
or U829 (N_829,In_1229,In_1767);
nor U830 (N_830,In_1042,N_204);
nand U831 (N_831,In_956,N_736);
or U832 (N_832,N_161,In_807);
and U833 (N_833,N_764,In_1028);
xor U834 (N_834,N_390,N_494);
nor U835 (N_835,In_1027,In_892);
and U836 (N_836,In_982,In_625);
or U837 (N_837,N_626,N_207);
or U838 (N_838,N_91,In_131);
xor U839 (N_839,N_84,In_270);
or U840 (N_840,N_533,In_1824);
xnor U841 (N_841,In_1751,N_63);
nand U842 (N_842,In_1705,In_768);
xnor U843 (N_843,N_451,N_126);
nand U844 (N_844,N_729,In_1336);
nor U845 (N_845,In_712,N_398);
and U846 (N_846,N_244,N_154);
or U847 (N_847,N_763,N_564);
or U848 (N_848,In_298,N_138);
nor U849 (N_849,N_485,N_283);
xor U850 (N_850,N_103,N_411);
xor U851 (N_851,In_898,In_355);
and U852 (N_852,In_1977,In_789);
and U853 (N_853,N_610,In_90);
and U854 (N_854,N_268,N_601);
nand U855 (N_855,In_139,In_177);
nor U856 (N_856,N_416,In_1612);
xor U857 (N_857,N_210,In_48);
xnor U858 (N_858,N_415,In_1474);
nand U859 (N_859,N_266,N_417);
or U860 (N_860,N_3,In_214);
nand U861 (N_861,In_1151,In_1264);
nand U862 (N_862,In_1021,In_1315);
or U863 (N_863,In_1200,In_344);
and U864 (N_864,In_217,N_474);
xnor U865 (N_865,In_421,N_508);
nand U866 (N_866,N_444,N_489);
and U867 (N_867,N_213,In_144);
nor U868 (N_868,In_1905,In_1083);
nor U869 (N_869,N_76,N_717);
or U870 (N_870,N_503,N_713);
nand U871 (N_871,N_184,In_1639);
and U872 (N_872,In_1314,In_338);
nand U873 (N_873,N_439,N_104);
and U874 (N_874,In_935,N_734);
nor U875 (N_875,In_386,N_571);
or U876 (N_876,N_744,N_668);
nor U877 (N_877,In_1817,N_459);
nor U878 (N_878,N_572,N_640);
nand U879 (N_879,In_891,N_568);
xnor U880 (N_880,N_24,N_588);
xnor U881 (N_881,N_710,N_428);
nand U882 (N_882,In_1130,N_431);
nor U883 (N_883,In_623,N_114);
nor U884 (N_884,In_562,In_1319);
xnor U885 (N_885,N_457,N_700);
and U886 (N_886,N_501,In_1771);
nand U887 (N_887,In_1761,N_498);
nand U888 (N_888,N_673,In_1054);
nor U889 (N_889,N_118,N_792);
xnor U890 (N_890,N_519,N_463);
xnor U891 (N_891,In_47,In_690);
nor U892 (N_892,In_137,N_495);
nor U893 (N_893,In_134,In_352);
or U894 (N_894,In_578,In_336);
xor U895 (N_895,In_1825,N_352);
and U896 (N_896,In_1326,N_175);
and U897 (N_897,N_343,N_637);
xnor U898 (N_898,In_632,In_1546);
nand U899 (N_899,In_1029,N_136);
nor U900 (N_900,In_941,N_514);
nand U901 (N_901,N_702,N_653);
or U902 (N_902,N_573,In_613);
nor U903 (N_903,N_483,In_243);
nor U904 (N_904,N_487,N_250);
nand U905 (N_905,N_643,In_558);
or U906 (N_906,In_601,In_367);
nor U907 (N_907,In_208,In_1068);
and U908 (N_908,N_429,In_592);
or U909 (N_909,N_215,N_106);
xnor U910 (N_910,In_1424,In_1747);
nor U911 (N_911,N_100,N_74);
nor U912 (N_912,N_676,In_1487);
or U913 (N_913,N_731,N_585);
nor U914 (N_914,N_310,In_366);
nand U915 (N_915,N_538,In_1551);
nand U916 (N_916,In_1073,In_1390);
or U917 (N_917,In_1307,N_371);
and U918 (N_918,In_604,N_614);
nand U919 (N_919,N_470,N_780);
nand U920 (N_920,In_30,In_1680);
nand U921 (N_921,N_748,N_465);
or U922 (N_922,In_1348,In_1258);
nor U923 (N_923,N_677,N_582);
xor U924 (N_924,N_61,In_253);
nor U925 (N_925,N_769,In_665);
or U926 (N_926,N_176,In_879);
nor U927 (N_927,N_27,In_736);
nand U928 (N_928,N_738,In_1113);
and U929 (N_929,In_684,N_762);
xor U930 (N_930,In_1697,In_1103);
and U931 (N_931,In_284,N_445);
or U932 (N_932,N_32,N_414);
nor U933 (N_933,N_57,In_652);
or U934 (N_934,N_608,In_875);
xnor U935 (N_935,N_699,N_773);
nand U936 (N_936,N_632,In_550);
nor U937 (N_937,N_92,N_581);
and U938 (N_938,In_679,N_388);
nand U939 (N_939,N_600,In_405);
and U940 (N_940,In_396,N_430);
or U941 (N_941,In_1506,N_196);
nor U942 (N_942,In_1844,N_372);
or U943 (N_943,N_443,N_77);
nand U944 (N_944,In_865,In_779);
xor U945 (N_945,In_1237,In_143);
nand U946 (N_946,In_1299,In_27);
or U947 (N_947,In_1427,N_446);
or U948 (N_948,N_124,N_510);
xor U949 (N_949,In_1913,N_742);
nand U950 (N_950,In_407,In_448);
xnor U951 (N_951,In_393,In_996);
nor U952 (N_952,In_116,In_556);
and U953 (N_953,N_527,In_1611);
and U954 (N_954,N_565,In_862);
or U955 (N_955,In_1158,N_127);
nor U956 (N_956,N_557,In_1530);
xnor U957 (N_957,In_81,In_292);
nand U958 (N_958,N_258,In_1664);
and U959 (N_959,In_1400,In_520);
xor U960 (N_960,In_1891,In_955);
nor U961 (N_961,N_131,N_165);
and U962 (N_962,In_1247,In_1166);
and U963 (N_963,In_707,In_356);
or U964 (N_964,N_661,In_228);
nor U965 (N_965,In_290,In_1431);
and U966 (N_966,N_532,N_685);
or U967 (N_967,N_381,In_683);
nand U968 (N_968,N_657,N_405);
or U969 (N_969,N_675,N_784);
nand U970 (N_970,In_1931,N_412);
nand U971 (N_971,In_887,N_598);
xor U972 (N_972,In_13,In_1367);
nor U973 (N_973,N_606,N_655);
xor U974 (N_974,N_486,N_618);
nand U975 (N_975,In_63,N_691);
xnor U976 (N_976,In_819,N_90);
nand U977 (N_977,N_300,In_1531);
xnor U978 (N_978,N_751,In_1579);
nand U979 (N_979,N_552,N_1);
or U980 (N_980,In_1454,N_659);
and U981 (N_981,N_427,In_676);
or U982 (N_982,N_770,In_1821);
nand U983 (N_983,N_592,In_324);
nand U984 (N_984,N_786,N_315);
and U985 (N_985,In_791,In_226);
nand U986 (N_986,N_739,In_917);
xor U987 (N_987,N_746,In_467);
xnor U988 (N_988,N_774,N_467);
nand U989 (N_989,N_684,N_604);
nor U990 (N_990,N_631,In_938);
xor U991 (N_991,N_785,N_630);
nor U992 (N_992,In_1804,N_12);
nand U993 (N_993,N_78,N_730);
or U994 (N_994,N_584,In_1405);
nor U995 (N_995,In_1046,In_1981);
nor U996 (N_996,N_26,In_946);
or U997 (N_997,In_135,N_648);
nor U998 (N_998,N_404,In_148);
and U999 (N_999,In_804,N_358);
nor U1000 (N_1000,In_1216,N_8);
nor U1001 (N_1001,In_1565,In_1072);
xnor U1002 (N_1002,N_563,In_1380);
nor U1003 (N_1003,In_43,N_745);
and U1004 (N_1004,N_286,In_1961);
nor U1005 (N_1005,N_775,In_530);
xnor U1006 (N_1006,N_550,In_414);
xnor U1007 (N_1007,In_1202,N_69);
or U1008 (N_1008,In_1555,N_20);
or U1009 (N_1009,N_555,N_265);
or U1010 (N_1010,N_794,N_535);
and U1011 (N_1011,N_607,In_59);
xnor U1012 (N_1012,In_358,N_484);
nor U1013 (N_1013,N_325,N_344);
nor U1014 (N_1014,N_221,In_1984);
xnor U1015 (N_1015,In_1744,In_1417);
and U1016 (N_1016,N_613,In_615);
xnor U1017 (N_1017,N_323,N_728);
and U1018 (N_1018,N_442,N_15);
or U1019 (N_1019,In_450,In_197);
or U1020 (N_1020,N_779,In_1312);
nor U1021 (N_1021,In_1843,In_1969);
nor U1022 (N_1022,In_319,N_620);
xor U1023 (N_1023,N_635,In_1413);
and U1024 (N_1024,N_29,N_419);
nor U1025 (N_1025,In_1037,N_278);
nor U1026 (N_1026,In_380,In_438);
xnor U1027 (N_1027,N_455,N_332);
or U1028 (N_1028,In_686,In_147);
and U1029 (N_1029,In_816,N_521);
or U1030 (N_1030,N_757,N_391);
xor U1031 (N_1031,N_719,N_394);
nand U1032 (N_1032,In_735,N_43);
nand U1033 (N_1033,In_140,In_568);
nor U1034 (N_1034,N_0,N_513);
nor U1035 (N_1035,In_1999,In_1521);
and U1036 (N_1036,In_794,In_1382);
or U1037 (N_1037,N_650,N_490);
or U1038 (N_1038,N_334,In_987);
xnor U1039 (N_1039,In_463,In_501);
and U1040 (N_1040,In_1514,In_511);
or U1041 (N_1041,In_1349,N_464);
nand U1042 (N_1042,N_440,In_846);
nor U1043 (N_1043,In_512,N_462);
and U1044 (N_1044,In_1868,N_365);
nor U1045 (N_1045,N_73,In_42);
nand U1046 (N_1046,In_1475,N_229);
xnor U1047 (N_1047,N_537,N_654);
or U1048 (N_1048,In_1138,In_591);
and U1049 (N_1049,N_424,In_1193);
xnor U1050 (N_1050,N_182,In_129);
nor U1051 (N_1051,N_406,N_18);
nor U1052 (N_1052,In_1187,N_38);
xor U1053 (N_1053,N_515,N_23);
and U1054 (N_1054,N_456,In_1881);
and U1055 (N_1055,N_615,N_525);
nand U1056 (N_1056,N_536,In_852);
nor U1057 (N_1057,In_1625,N_80);
or U1058 (N_1058,N_496,N_664);
and U1059 (N_1059,N_83,N_468);
xnor U1060 (N_1060,N_737,N_293);
nand U1061 (N_1061,N_432,In_868);
and U1062 (N_1062,In_954,In_1376);
or U1063 (N_1063,In_857,N_203);
or U1064 (N_1064,In_1875,In_759);
xnor U1065 (N_1065,In_1392,In_207);
xnor U1066 (N_1066,In_746,In_782);
nor U1067 (N_1067,N_768,In_1598);
nor U1068 (N_1068,In_1816,N_576);
xnor U1069 (N_1069,N_85,In_1428);
xnor U1070 (N_1070,N_651,N_605);
and U1071 (N_1071,In_984,In_1679);
xnor U1072 (N_1072,N_232,N_551);
and U1073 (N_1073,In_629,In_1199);
nor U1074 (N_1074,In_728,N_612);
nor U1075 (N_1075,In_1941,In_273);
and U1076 (N_1076,In_933,N_87);
nor U1077 (N_1077,N_421,In_770);
and U1078 (N_1078,N_752,In_1654);
nor U1079 (N_1079,N_226,In_400);
nor U1080 (N_1080,N_505,In_532);
nand U1081 (N_1081,N_361,N_438);
nor U1082 (N_1082,N_529,N_418);
xor U1083 (N_1083,N_249,In_813);
nor U1084 (N_1084,In_663,In_986);
nand U1085 (N_1085,N_319,In_1145);
and U1086 (N_1086,N_475,In_714);
nand U1087 (N_1087,N_526,In_709);
and U1088 (N_1088,N_298,N_299);
nor U1089 (N_1089,N_788,N_520);
nand U1090 (N_1090,In_1853,In_1397);
nor U1091 (N_1091,In_1515,N_683);
xor U1092 (N_1092,N_627,N_705);
nand U1093 (N_1093,N_236,In_1169);
xnor U1094 (N_1094,In_1733,N_461);
or U1095 (N_1095,N_750,In_234);
or U1096 (N_1096,In_1791,N_665);
nor U1097 (N_1097,In_1407,N_671);
xor U1098 (N_1098,In_1162,In_678);
and U1099 (N_1099,N_543,In_216);
nand U1100 (N_1100,In_113,In_1497);
and U1101 (N_1101,In_1502,In_1440);
xor U1102 (N_1102,N_471,N_40);
nand U1103 (N_1103,In_33,In_966);
nor U1104 (N_1104,In_1520,In_1597);
or U1105 (N_1105,N_558,N_666);
or U1106 (N_1106,N_599,In_1003);
nor U1107 (N_1107,In_1568,N_523);
nor U1108 (N_1108,N_656,N_178);
xor U1109 (N_1109,In_1700,In_1888);
and U1110 (N_1110,In_210,In_618);
xnor U1111 (N_1111,In_897,In_1024);
nor U1112 (N_1112,In_1517,In_543);
nand U1113 (N_1113,In_773,In_94);
nand U1114 (N_1114,In_1743,In_834);
xor U1115 (N_1115,In_112,In_1691);
nand U1116 (N_1116,In_1360,In_743);
xnor U1117 (N_1117,In_1829,In_91);
and U1118 (N_1118,N_331,In_1879);
and U1119 (N_1119,In_1460,In_1720);
nand U1120 (N_1120,N_629,In_1496);
nand U1121 (N_1121,N_649,In_1903);
nand U1122 (N_1122,In_980,N_68);
or U1123 (N_1123,N_771,N_162);
or U1124 (N_1124,In_294,N_530);
and U1125 (N_1125,N_711,In_56);
nor U1126 (N_1126,N_787,N_560);
or U1127 (N_1127,In_202,In_293);
nor U1128 (N_1128,N_580,In_110);
and U1129 (N_1129,N_401,In_1393);
or U1130 (N_1130,N_422,In_278);
or U1131 (N_1131,N_540,In_689);
xor U1132 (N_1132,In_976,In_1135);
xnor U1133 (N_1133,N_473,N_589);
nand U1134 (N_1134,In_1583,N_714);
nand U1135 (N_1135,N_31,In_762);
xnor U1136 (N_1136,In_853,In_340);
and U1137 (N_1137,N_217,N_516);
and U1138 (N_1138,N_641,N_567);
nand U1139 (N_1139,N_482,In_890);
or U1140 (N_1140,N_733,In_10);
nand U1141 (N_1141,In_1430,In_754);
or U1142 (N_1142,In_1595,In_100);
or U1143 (N_1143,In_211,In_303);
nor U1144 (N_1144,N_81,N_33);
nand U1145 (N_1145,In_1992,N_307);
nand U1146 (N_1146,In_842,In_1141);
nand U1147 (N_1147,In_1429,N_687);
nand U1148 (N_1148,N_94,N_346);
xor U1149 (N_1149,N_701,In_5);
nor U1150 (N_1150,N_509,In_750);
nand U1151 (N_1151,In_461,N_579);
nor U1152 (N_1152,N_11,N_721);
or U1153 (N_1153,In_1653,N_261);
nor U1154 (N_1154,N_797,N_435);
or U1155 (N_1155,In_1332,In_1836);
and U1156 (N_1156,In_786,N_531);
nand U1157 (N_1157,In_1637,In_624);
and U1158 (N_1158,N_638,In_1618);
xor U1159 (N_1159,In_1663,N_351);
nor U1160 (N_1160,In_900,N_479);
xnor U1161 (N_1161,In_309,In_1197);
nand U1162 (N_1162,In_715,In_838);
nor U1163 (N_1163,N_791,In_930);
xnor U1164 (N_1164,In_590,N_105);
nand U1165 (N_1165,In_466,N_281);
and U1166 (N_1166,N_718,N_7);
nand U1167 (N_1167,In_225,N_34);
nand U1168 (N_1168,N_151,N_480);
nor U1169 (N_1169,N_436,In_187);
nand U1170 (N_1170,In_188,N_624);
nand U1171 (N_1171,N_539,N_622);
nor U1172 (N_1172,In_989,In_1058);
nand U1173 (N_1173,In_1830,In_1527);
or U1174 (N_1174,In_1092,In_428);
or U1175 (N_1175,In_1511,N_679);
nand U1176 (N_1176,N_740,N_545);
and U1177 (N_1177,N_375,In_1052);
nor U1178 (N_1178,In_923,N_4);
nand U1179 (N_1179,In_32,In_855);
and U1180 (N_1180,In_1123,In_1901);
xor U1181 (N_1181,N_616,N_112);
and U1182 (N_1182,N_709,N_399);
xnor U1183 (N_1183,In_1063,N_595);
nand U1184 (N_1184,In_1301,In_1334);
nand U1185 (N_1185,N_219,N_625);
nor U1186 (N_1186,N_670,In_417);
and U1187 (N_1187,In_648,N_400);
or U1188 (N_1188,N_192,In_1181);
and U1189 (N_1189,N_144,N_662);
and U1190 (N_1190,In_1041,In_717);
and U1191 (N_1191,N_481,N_241);
and U1192 (N_1192,N_753,N_646);
xnor U1193 (N_1193,In_1902,In_375);
nor U1194 (N_1194,In_1340,N_159);
nor U1195 (N_1195,In_167,In_975);
nor U1196 (N_1196,N_205,N_644);
and U1197 (N_1197,N_364,N_17);
xnor U1198 (N_1198,In_1281,N_754);
or U1199 (N_1199,N_502,N_681);
nor U1200 (N_1200,N_469,In_76);
or U1201 (N_1201,N_1060,N_562);
or U1202 (N_1202,N_952,N_851);
xnor U1203 (N_1203,In_1015,N_139);
xnor U1204 (N_1204,N_453,N_1116);
and U1205 (N_1205,N_1186,N_890);
xnor U1206 (N_1206,N_1114,N_1112);
and U1207 (N_1207,N_704,N_1072);
and U1208 (N_1208,N_919,N_1125);
nand U1209 (N_1209,In_158,N_93);
nor U1210 (N_1210,N_868,N_957);
xor U1211 (N_1211,N_992,N_1185);
and U1212 (N_1212,N_727,N_1018);
or U1213 (N_1213,In_650,N_849);
xor U1214 (N_1214,In_1726,N_972);
nand U1215 (N_1215,N_1001,N_819);
nand U1216 (N_1216,N_1070,In_432);
nor U1217 (N_1217,N_1034,N_1189);
nor U1218 (N_1218,In_1101,N_1055);
xor U1219 (N_1219,N_645,N_1096);
and U1220 (N_1220,N_802,N_437);
or U1221 (N_1221,N_948,N_507);
nor U1222 (N_1222,N_37,N_1180);
nand U1223 (N_1223,N_122,N_1118);
or U1224 (N_1224,N_796,N_758);
xnor U1225 (N_1225,N_45,N_403);
nor U1226 (N_1226,N_695,N_894);
or U1227 (N_1227,N_1164,In_1265);
nand U1228 (N_1228,N_871,N_993);
xnor U1229 (N_1229,In_288,In_379);
nor U1230 (N_1230,N_917,N_682);
and U1231 (N_1231,N_901,In_730);
nand U1232 (N_1232,N_1012,N_946);
nor U1233 (N_1233,N_160,N_1102);
nor U1234 (N_1234,N_884,N_932);
or U1235 (N_1235,In_179,In_1695);
and U1236 (N_1236,N_316,N_522);
or U1237 (N_1237,In_275,N_831);
nand U1238 (N_1238,N_1166,In_9);
or U1239 (N_1239,N_1195,N_847);
xnor U1240 (N_1240,N_813,N_949);
nor U1241 (N_1241,N_872,In_1979);
nor U1242 (N_1242,N_732,N_896);
nor U1243 (N_1243,In_856,N_867);
or U1244 (N_1244,N_982,In_1807);
or U1245 (N_1245,N_383,N_1076);
nor U1246 (N_1246,In_364,In_612);
and U1247 (N_1247,N_199,N_782);
nor U1248 (N_1248,N_71,In_713);
nor U1249 (N_1249,In_1641,N_1065);
nor U1250 (N_1250,N_953,N_667);
nand U1251 (N_1251,N_450,N_826);
nor U1252 (N_1252,N_789,N_1171);
nor U1253 (N_1253,N_820,N_466);
nand U1254 (N_1254,N_969,In_12);
nand U1255 (N_1255,In_945,N_609);
xnor U1256 (N_1256,In_1775,N_723);
nor U1257 (N_1257,In_745,N_866);
nand U1258 (N_1258,N_1178,In_384);
xor U1259 (N_1259,In_1998,N_1058);
nor U1260 (N_1260,N_930,N_251);
nand U1261 (N_1261,N_950,N_425);
nor U1262 (N_1262,In_62,N_995);
and U1263 (N_1263,N_693,N_996);
or U1264 (N_1264,In_1228,N_233);
xor U1265 (N_1265,N_922,N_981);
nand U1266 (N_1266,N_840,N_743);
or U1267 (N_1267,In_1781,In_73);
xor U1268 (N_1268,N_1027,In_496);
nand U1269 (N_1269,In_1532,N_1179);
nand U1270 (N_1270,N_1146,In_92);
or U1271 (N_1271,In_1805,N_845);
xnor U1272 (N_1272,In_1306,N_119);
nand U1273 (N_1273,N_282,N_1100);
xor U1274 (N_1274,N_1086,N_1005);
and U1275 (N_1275,In_1750,N_556);
nand U1276 (N_1276,N_1028,N_441);
nor U1277 (N_1277,N_1030,N_426);
nor U1278 (N_1278,N_1139,N_885);
nor U1279 (N_1279,In_723,N_793);
xor U1280 (N_1280,N_544,In_93);
nand U1281 (N_1281,N_688,N_834);
nand U1282 (N_1282,N_678,N_900);
nand U1283 (N_1283,N_409,In_1983);
or U1284 (N_1284,N_1071,N_452);
nor U1285 (N_1285,N_1098,N_1088);
nand U1286 (N_1286,N_943,N_940);
and U1287 (N_1287,N_1080,N_835);
and U1288 (N_1288,N_1092,In_1755);
xnor U1289 (N_1289,N_959,N_339);
and U1290 (N_1290,N_965,N_897);
xor U1291 (N_1291,In_1994,N_855);
nor U1292 (N_1292,N_548,In_50);
xor U1293 (N_1293,N_832,N_611);
nor U1294 (N_1294,N_1140,N_1194);
and U1295 (N_1295,N_1095,N_497);
or U1296 (N_1296,N_1187,N_978);
or U1297 (N_1297,In_371,N_1067);
nor U1298 (N_1298,N_1198,N_756);
nor U1299 (N_1299,N_1062,In_747);
or U1300 (N_1300,In_21,In_1147);
and U1301 (N_1301,N_617,N_725);
nand U1302 (N_1302,N_674,N_1050);
xnor U1303 (N_1303,N_1184,In_431);
nand U1304 (N_1304,N_694,In_1906);
nor U1305 (N_1305,In_925,In_1813);
xor U1306 (N_1306,N_1121,N_720);
nand U1307 (N_1307,In_1404,N_1053);
nor U1308 (N_1308,In_1756,In_184);
nand U1309 (N_1309,N_1167,N_517);
or U1310 (N_1310,In_912,N_596);
xnor U1311 (N_1311,N_1130,N_145);
nor U1312 (N_1312,N_1181,N_593);
and U1313 (N_1313,N_759,N_827);
xnor U1314 (N_1314,In_1179,N_270);
nand U1315 (N_1315,In_1592,N_336);
xnor U1316 (N_1316,N_970,In_606);
nor U1317 (N_1317,N_899,N_518);
or U1318 (N_1318,N_844,N_594);
nand U1319 (N_1319,N_747,In_669);
xor U1320 (N_1320,N_947,N_882);
nand U1321 (N_1321,In_1104,N_876);
and U1322 (N_1322,N_1035,N_926);
nand U1323 (N_1323,In_920,N_856);
or U1324 (N_1324,N_858,In_305);
nor U1325 (N_1325,N_306,N_811);
nor U1326 (N_1326,N_1081,N_1077);
or U1327 (N_1327,N_434,N_857);
nor U1328 (N_1328,N_1142,N_636);
or U1329 (N_1329,N_1155,N_460);
nand U1330 (N_1330,N_1097,N_1061);
nor U1331 (N_1331,N_913,N_878);
nor U1332 (N_1332,N_1003,N_755);
xor U1333 (N_1333,N_1068,N_150);
nand U1334 (N_1334,N_143,In_1366);
nor U1335 (N_1335,In_617,N_861);
nand U1336 (N_1336,N_1110,N_1010);
and U1337 (N_1337,In_1086,N_852);
nand U1338 (N_1338,In_1472,In_1710);
nor U1339 (N_1339,N_989,N_898);
nand U1340 (N_1340,In_1362,N_111);
or U1341 (N_1341,N_936,N_967);
nor U1342 (N_1342,In_470,N_1091);
and U1343 (N_1343,N_961,In_1801);
or U1344 (N_1344,N_825,N_1190);
xor U1345 (N_1345,In_1865,N_909);
and U1346 (N_1346,N_994,In_156);
nand U1347 (N_1347,In_1266,N_850);
nor U1348 (N_1348,N_939,N_954);
nand U1349 (N_1349,N_883,N_777);
xnor U1350 (N_1350,In_1966,N_893);
or U1351 (N_1351,In_1855,In_121);
and U1352 (N_1352,In_1062,N_1047);
and U1353 (N_1353,N_230,N_1032);
nor U1354 (N_1354,N_761,N_1156);
xnor U1355 (N_1355,N_135,N_955);
nand U1356 (N_1356,In_1335,N_925);
and U1357 (N_1357,N_1128,N_1014);
nand U1358 (N_1358,N_1122,N_854);
nand U1359 (N_1359,N_420,N_963);
nor U1360 (N_1360,N_988,In_1812);
and U1361 (N_1361,In_330,N_760);
xor U1362 (N_1362,N_1054,In_1600);
or U1363 (N_1363,N_1007,N_570);
or U1364 (N_1364,N_51,N_575);
nand U1365 (N_1365,In_462,N_805);
xor U1366 (N_1366,In_950,N_783);
nand U1367 (N_1367,N_931,N_342);
nor U1368 (N_1368,N_928,N_942);
and U1369 (N_1369,N_1052,N_968);
or U1370 (N_1370,In_1796,N_191);
nor U1371 (N_1371,N_937,N_1120);
nor U1372 (N_1372,In_695,N_549);
and U1373 (N_1373,N_1153,N_1066);
nor U1374 (N_1374,In_1811,N_829);
or U1375 (N_1375,N_990,In_973);
or U1376 (N_1376,N_1082,N_1165);
or U1377 (N_1377,In_722,N_803);
nor U1378 (N_1378,In_1640,N_1011);
and U1379 (N_1379,N_488,N_1057);
or U1380 (N_1380,N_1157,In_561);
or U1381 (N_1381,N_1158,N_137);
xor U1382 (N_1382,In_929,N_628);
and U1383 (N_1383,In_1528,In_150);
and U1384 (N_1384,N_220,N_1031);
or U1385 (N_1385,N_906,N_1135);
nor U1386 (N_1386,N_663,N_413);
nand U1387 (N_1387,In_691,N_817);
and U1388 (N_1388,In_170,N_228);
nand U1389 (N_1389,N_542,In_792);
nor U1390 (N_1390,N_841,N_547);
nor U1391 (N_1391,N_1108,In_1885);
or U1392 (N_1392,N_1023,N_801);
xor U1393 (N_1393,N_696,N_880);
or U1394 (N_1394,In_132,N_1124);
nor U1395 (N_1395,In_283,N_933);
and U1396 (N_1396,In_1168,N_1015);
or U1397 (N_1397,N_918,N_818);
nor U1398 (N_1398,N_887,N_951);
xnor U1399 (N_1399,N_707,N_934);
and U1400 (N_1400,N_904,N_1161);
nor U1401 (N_1401,N_839,N_1170);
nor U1402 (N_1402,In_348,N_903);
nand U1403 (N_1403,N_1131,N_511);
and U1404 (N_1404,N_158,N_1069);
and U1405 (N_1405,N_1020,N_977);
nand U1406 (N_1406,N_397,In_1284);
xnor U1407 (N_1407,In_993,N_859);
nor U1408 (N_1408,In_1586,N_1042);
nor U1409 (N_1409,In_160,N_692);
xor U1410 (N_1410,N_860,N_1133);
or U1411 (N_1411,N_838,N_1021);
nor U1412 (N_1412,N_958,N_964);
or U1413 (N_1413,N_708,N_892);
or U1414 (N_1414,In_544,N_1136);
nor U1415 (N_1415,N_865,In_593);
nand U1416 (N_1416,N_804,In_368);
xor U1417 (N_1417,In_351,N_1182);
or U1418 (N_1418,N_735,N_862);
and U1419 (N_1419,In_661,N_1079);
or U1420 (N_1420,N_726,In_1087);
and U1421 (N_1421,N_810,In_196);
or U1422 (N_1422,N_836,N_1137);
xnor U1423 (N_1423,N_776,N_1094);
or U1424 (N_1424,N_1063,N_1188);
and U1425 (N_1425,N_587,N_288);
and U1426 (N_1426,N_492,N_385);
nand U1427 (N_1427,In_1461,N_493);
nand U1428 (N_1428,N_888,N_879);
and U1429 (N_1429,N_778,N_984);
nor U1430 (N_1430,In_257,N_476);
xnor U1431 (N_1431,N_50,N_986);
nand U1432 (N_1432,N_1064,In_726);
nand U1433 (N_1433,N_941,N_1134);
nor U1434 (N_1434,N_1177,In_1616);
xnor U1435 (N_1435,N_1039,N_1090);
or U1436 (N_1436,N_39,N_1192);
xor U1437 (N_1437,N_559,In_806);
nand U1438 (N_1438,In_1944,N_902);
or U1439 (N_1439,In_1642,N_1115);
xor U1440 (N_1440,N_956,N_895);
and U1441 (N_1441,N_1176,N_1127);
and U1442 (N_1442,N_619,N_863);
xor U1443 (N_1443,N_546,N_586);
xnor U1444 (N_1444,In_398,N_382);
and U1445 (N_1445,In_1776,N_1111);
nor U1446 (N_1446,N_749,N_703);
or U1447 (N_1447,N_1147,In_1880);
or U1448 (N_1448,N_822,N_686);
nor U1449 (N_1449,In_885,N_806);
nand U1450 (N_1450,In_522,N_1099);
xor U1451 (N_1451,In_729,In_1099);
nor U1452 (N_1452,In_934,N_1148);
xor U1453 (N_1453,N_1126,In_322);
and U1454 (N_1454,In_682,N_590);
or U1455 (N_1455,N_689,N_448);
nand U1456 (N_1456,N_966,N_935);
xnor U1457 (N_1457,N_49,In_547);
or U1458 (N_1458,N_623,N_809);
nor U1459 (N_1459,N_1149,N_267);
or U1460 (N_1460,N_1009,N_1174);
xor U1461 (N_1461,N_169,In_940);
or U1462 (N_1462,In_1990,In_89);
and U1463 (N_1463,N_504,In_1635);
nand U1464 (N_1464,In_1452,N_1038);
nor U1465 (N_1465,In_483,N_1046);
nor U1466 (N_1466,N_772,N_808);
and U1467 (N_1467,In_1719,N_938);
nor U1468 (N_1468,N_975,N_211);
and U1469 (N_1469,N_915,N_1132);
xor U1470 (N_1470,In_1213,N_921);
nand U1471 (N_1471,N_1101,N_1048);
nor U1472 (N_1472,In_1549,N_846);
or U1473 (N_1473,N_962,N_1117);
and U1474 (N_1474,N_907,N_369);
and U1475 (N_1475,N_1074,In_277);
or U1476 (N_1476,N_916,N_672);
nor U1477 (N_1477,N_1073,N_1036);
xnor U1478 (N_1478,N_1026,N_179);
nor U1479 (N_1479,N_973,N_724);
or U1480 (N_1480,N_1016,N_1049);
nand U1481 (N_1481,N_1085,In_1465);
nor U1482 (N_1482,N_712,N_908);
nor U1483 (N_1483,N_1025,In_1847);
or U1484 (N_1484,In_907,N_971);
nor U1485 (N_1485,N_491,In_3);
and U1486 (N_1486,N_1056,N_828);
and U1487 (N_1487,N_1168,In_79);
and U1488 (N_1488,In_835,In_576);
and U1489 (N_1489,In_809,N_227);
nor U1490 (N_1490,N_914,N_1145);
nand U1491 (N_1491,N_991,N_1172);
nand U1492 (N_1492,N_1051,In_1304);
xor U1493 (N_1493,N_767,N_960);
xor U1494 (N_1494,In_867,N_987);
nor U1495 (N_1495,N_1045,N_814);
and U1496 (N_1496,N_423,N_976);
and U1497 (N_1497,N_1123,N_1059);
xor U1498 (N_1498,N_944,N_877);
xnor U1499 (N_1499,N_815,N_553);
nor U1500 (N_1500,N_327,N_698);
and U1501 (N_1501,N_602,N_1107);
nor U1502 (N_1502,N_433,In_23);
and U1503 (N_1503,N_554,N_1033);
nand U1504 (N_1504,N_881,In_1328);
xnor U1505 (N_1505,N_924,In_101);
or U1506 (N_1506,N_359,In_185);
nor U1507 (N_1507,N_500,N_1006);
or U1508 (N_1508,N_911,In_653);
nand U1509 (N_1509,In_692,N_848);
nand U1510 (N_1510,N_1169,N_979);
nand U1511 (N_1511,In_731,N_458);
xor U1512 (N_1512,In_1488,N_1199);
xor U1513 (N_1513,In_1730,In_1955);
nand U1514 (N_1514,N_1160,N_633);
and U1515 (N_1515,In_630,In_485);
and U1516 (N_1516,N_873,N_1078);
or U1517 (N_1517,N_621,N_1029);
xor U1518 (N_1518,In_999,N_945);
nor U1519 (N_1519,N_1089,N_1129);
xor U1520 (N_1520,N_1152,N_86);
xor U1521 (N_1521,In_552,In_936);
and U1522 (N_1522,In_1143,N_923);
nor U1523 (N_1523,In_1185,N_1138);
or U1524 (N_1524,In_1426,N_1105);
nor U1525 (N_1525,N_583,N_980);
or U1526 (N_1526,N_790,N_1087);
xor U1527 (N_1527,N_722,In_811);
or U1528 (N_1528,N_603,N_1197);
nor U1529 (N_1529,N_1022,N_1004);
and U1530 (N_1530,N_1093,N_1017);
xnor U1531 (N_1531,N_597,In_1458);
and U1532 (N_1532,In_260,In_86);
xnor U1533 (N_1533,N_578,N_889);
nand U1534 (N_1534,N_837,N_997);
nor U1535 (N_1535,N_1109,N_1106);
and U1536 (N_1536,N_715,N_910);
and U1537 (N_1537,N_30,N_875);
xnor U1538 (N_1538,N_999,N_830);
nand U1539 (N_1539,N_929,N_1193);
and U1540 (N_1540,In_1699,In_1157);
and U1541 (N_1541,N_905,In_203);
nand U1542 (N_1542,In_321,N_347);
nand U1543 (N_1543,N_1119,N_566);
nor U1544 (N_1544,N_1041,In_327);
nand U1545 (N_1545,N_920,In_1278);
nand U1546 (N_1546,N_1150,In_26);
xnor U1547 (N_1547,N_912,N_1144);
or U1548 (N_1548,N_1163,N_1175);
nand U1549 (N_1549,N_1183,N_983);
and U1550 (N_1550,N_1024,N_1196);
nor U1551 (N_1551,N_869,N_447);
or U1552 (N_1552,N_454,N_891);
xnor U1553 (N_1553,In_1953,N_998);
and U1554 (N_1554,N_477,N_1104);
nor U1555 (N_1555,N_402,N_1043);
nor U1556 (N_1556,N_690,N_843);
and U1557 (N_1557,N_1151,N_189);
or U1558 (N_1558,In_563,N_246);
and U1559 (N_1559,N_823,N_304);
xor U1560 (N_1560,N_524,N_1162);
and U1561 (N_1561,In_1850,N_833);
or U1562 (N_1562,N_341,N_985);
nor U1563 (N_1563,N_1113,In_549);
or U1564 (N_1564,N_807,N_870);
nand U1565 (N_1565,N_512,N_886);
nor U1566 (N_1566,N_506,N_499);
nand U1567 (N_1567,N_1008,N_1143);
xnor U1568 (N_1568,N_1173,N_639);
or U1569 (N_1569,N_1154,N_642);
nor U1570 (N_1570,N_1103,N_1019);
nor U1571 (N_1571,In_626,In_1437);
nor U1572 (N_1572,N_1000,In_1991);
xor U1573 (N_1573,In_1325,N_591);
nor U1574 (N_1574,N_1044,N_974);
xnor U1575 (N_1575,N_864,N_149);
xnor U1576 (N_1576,N_716,N_1002);
xnor U1577 (N_1577,N_376,In_614);
and U1578 (N_1578,In_261,In_411);
nand U1579 (N_1579,N_25,N_816);
xnor U1580 (N_1580,In_927,In_1582);
nand U1581 (N_1581,N_190,N_874);
nand U1582 (N_1582,N_799,N_333);
nor U1583 (N_1583,In_577,N_561);
and U1584 (N_1584,N_853,N_842);
or U1585 (N_1585,In_536,In_1070);
nand U1586 (N_1586,N_214,N_766);
and U1587 (N_1587,In_127,N_824);
nand U1588 (N_1588,In_1146,N_812);
nor U1589 (N_1589,N_534,N_821);
xnor U1590 (N_1590,In_959,N_98);
and U1591 (N_1591,N_1013,N_1191);
and U1592 (N_1592,N_569,N_1075);
nand U1593 (N_1593,N_1083,N_1159);
or U1594 (N_1594,In_815,N_800);
nor U1595 (N_1595,N_795,N_1084);
nor U1596 (N_1596,N_1037,N_741);
xor U1597 (N_1597,N_1141,In_362);
or U1598 (N_1598,N_1040,N_577);
or U1599 (N_1599,N_188,N_927);
or U1600 (N_1600,N_1312,N_1449);
or U1601 (N_1601,N_1250,N_1229);
nand U1602 (N_1602,N_1479,N_1364);
nand U1603 (N_1603,N_1267,N_1456);
or U1604 (N_1604,N_1290,N_1533);
xor U1605 (N_1605,N_1204,N_1462);
xor U1606 (N_1606,N_1279,N_1294);
nand U1607 (N_1607,N_1428,N_1504);
nor U1608 (N_1608,N_1383,N_1409);
nand U1609 (N_1609,N_1342,N_1548);
nor U1610 (N_1610,N_1522,N_1245);
or U1611 (N_1611,N_1315,N_1519);
xor U1612 (N_1612,N_1436,N_1272);
nor U1613 (N_1613,N_1368,N_1212);
or U1614 (N_1614,N_1230,N_1460);
nand U1615 (N_1615,N_1343,N_1202);
xnor U1616 (N_1616,N_1545,N_1553);
nand U1617 (N_1617,N_1253,N_1201);
nand U1618 (N_1618,N_1538,N_1213);
xnor U1619 (N_1619,N_1494,N_1236);
nand U1620 (N_1620,N_1340,N_1339);
nand U1621 (N_1621,N_1411,N_1405);
xnor U1622 (N_1622,N_1255,N_1510);
and U1623 (N_1623,N_1419,N_1572);
xor U1624 (N_1624,N_1222,N_1505);
and U1625 (N_1625,N_1393,N_1549);
xnor U1626 (N_1626,N_1225,N_1567);
or U1627 (N_1627,N_1521,N_1265);
and U1628 (N_1628,N_1321,N_1503);
xnor U1629 (N_1629,N_1446,N_1324);
xnor U1630 (N_1630,N_1431,N_1484);
nor U1631 (N_1631,N_1478,N_1264);
or U1632 (N_1632,N_1218,N_1260);
or U1633 (N_1633,N_1427,N_1273);
nand U1634 (N_1634,N_1248,N_1281);
or U1635 (N_1635,N_1286,N_1251);
xor U1636 (N_1636,N_1376,N_1358);
or U1637 (N_1637,N_1524,N_1475);
nor U1638 (N_1638,N_1214,N_1491);
nor U1639 (N_1639,N_1327,N_1566);
nand U1640 (N_1640,N_1313,N_1437);
or U1641 (N_1641,N_1380,N_1448);
nor U1642 (N_1642,N_1434,N_1216);
and U1643 (N_1643,N_1311,N_1473);
xnor U1644 (N_1644,N_1481,N_1283);
or U1645 (N_1645,N_1455,N_1247);
nor U1646 (N_1646,N_1599,N_1465);
nor U1647 (N_1647,N_1497,N_1374);
and U1648 (N_1648,N_1337,N_1438);
and U1649 (N_1649,N_1357,N_1464);
or U1650 (N_1650,N_1309,N_1477);
nor U1651 (N_1651,N_1583,N_1587);
nand U1652 (N_1652,N_1495,N_1317);
or U1653 (N_1653,N_1526,N_1512);
nand U1654 (N_1654,N_1386,N_1345);
xnor U1655 (N_1655,N_1378,N_1335);
or U1656 (N_1656,N_1454,N_1370);
and U1657 (N_1657,N_1365,N_1226);
and U1658 (N_1658,N_1389,N_1363);
nand U1659 (N_1659,N_1304,N_1242);
xnor U1660 (N_1660,N_1444,N_1301);
xnor U1661 (N_1661,N_1366,N_1288);
and U1662 (N_1662,N_1535,N_1221);
or U1663 (N_1663,N_1597,N_1573);
and U1664 (N_1664,N_1249,N_1332);
nand U1665 (N_1665,N_1412,N_1574);
nor U1666 (N_1666,N_1373,N_1596);
xnor U1667 (N_1667,N_1489,N_1487);
nand U1668 (N_1668,N_1447,N_1388);
and U1669 (N_1669,N_1530,N_1501);
nand U1670 (N_1670,N_1203,N_1470);
nor U1671 (N_1671,N_1275,N_1285);
xnor U1672 (N_1672,N_1562,N_1371);
nor U1673 (N_1673,N_1433,N_1341);
or U1674 (N_1674,N_1367,N_1268);
nand U1675 (N_1675,N_1308,N_1261);
nor U1676 (N_1676,N_1556,N_1537);
and U1677 (N_1677,N_1352,N_1356);
nor U1678 (N_1678,N_1550,N_1360);
and U1679 (N_1679,N_1490,N_1333);
nor U1680 (N_1680,N_1532,N_1403);
and U1681 (N_1681,N_1227,N_1557);
xor U1682 (N_1682,N_1421,N_1584);
nor U1683 (N_1683,N_1542,N_1582);
nor U1684 (N_1684,N_1554,N_1220);
nand U1685 (N_1685,N_1565,N_1392);
or U1686 (N_1686,N_1558,N_1207);
or U1687 (N_1687,N_1424,N_1257);
and U1688 (N_1688,N_1243,N_1523);
nor U1689 (N_1689,N_1420,N_1588);
and U1690 (N_1690,N_1570,N_1450);
xnor U1691 (N_1691,N_1507,N_1296);
xnor U1692 (N_1692,N_1568,N_1498);
xor U1693 (N_1693,N_1385,N_1440);
xor U1694 (N_1694,N_1458,N_1468);
nand U1695 (N_1695,N_1506,N_1509);
and U1696 (N_1696,N_1486,N_1577);
nand U1697 (N_1697,N_1406,N_1362);
nor U1698 (N_1698,N_1407,N_1298);
xor U1699 (N_1699,N_1234,N_1269);
or U1700 (N_1700,N_1502,N_1231);
and U1701 (N_1701,N_1316,N_1443);
nor U1702 (N_1702,N_1215,N_1320);
nor U1703 (N_1703,N_1598,N_1326);
nor U1704 (N_1704,N_1408,N_1330);
nor U1705 (N_1705,N_1539,N_1233);
or U1706 (N_1706,N_1461,N_1310);
nand U1707 (N_1707,N_1414,N_1520);
and U1708 (N_1708,N_1295,N_1452);
nor U1709 (N_1709,N_1280,N_1467);
or U1710 (N_1710,N_1543,N_1271);
nand U1711 (N_1711,N_1246,N_1435);
or U1712 (N_1712,N_1381,N_1476);
or U1713 (N_1713,N_1518,N_1552);
xnor U1714 (N_1714,N_1354,N_1559);
nand U1715 (N_1715,N_1235,N_1219);
nand U1716 (N_1716,N_1578,N_1463);
and U1717 (N_1717,N_1322,N_1482);
and U1718 (N_1718,N_1228,N_1353);
or U1719 (N_1719,N_1238,N_1579);
and U1720 (N_1720,N_1323,N_1571);
nand U1721 (N_1721,N_1423,N_1418);
nor U1722 (N_1722,N_1527,N_1457);
nand U1723 (N_1723,N_1529,N_1480);
xor U1724 (N_1724,N_1293,N_1355);
or U1725 (N_1725,N_1307,N_1351);
nor U1726 (N_1726,N_1391,N_1432);
nor U1727 (N_1727,N_1318,N_1282);
xor U1728 (N_1728,N_1400,N_1300);
and U1729 (N_1729,N_1511,N_1276);
nand U1730 (N_1730,N_1595,N_1241);
xnor U1731 (N_1731,N_1472,N_1387);
xor U1732 (N_1732,N_1546,N_1569);
nor U1733 (N_1733,N_1442,N_1541);
and U1734 (N_1734,N_1410,N_1211);
nor U1735 (N_1735,N_1589,N_1575);
nand U1736 (N_1736,N_1284,N_1372);
and U1737 (N_1737,N_1328,N_1302);
xor U1738 (N_1738,N_1223,N_1361);
or U1739 (N_1739,N_1397,N_1266);
and U1740 (N_1740,N_1586,N_1592);
nor U1741 (N_1741,N_1338,N_1344);
nand U1742 (N_1742,N_1451,N_1258);
and U1743 (N_1743,N_1439,N_1346);
or U1744 (N_1744,N_1534,N_1359);
or U1745 (N_1745,N_1206,N_1563);
nand U1746 (N_1746,N_1379,N_1292);
nor U1747 (N_1747,N_1237,N_1394);
nand U1748 (N_1748,N_1429,N_1398);
nand U1749 (N_1749,N_1517,N_1402);
or U1750 (N_1750,N_1453,N_1515);
nand U1751 (N_1751,N_1314,N_1287);
nor U1752 (N_1752,N_1306,N_1445);
and U1753 (N_1753,N_1240,N_1395);
nand U1754 (N_1754,N_1334,N_1263);
nand U1755 (N_1755,N_1404,N_1516);
nand U1756 (N_1756,N_1422,N_1254);
nor U1757 (N_1757,N_1580,N_1319);
and U1758 (N_1758,N_1384,N_1555);
nor U1759 (N_1759,N_1508,N_1540);
nand U1760 (N_1760,N_1401,N_1396);
nor U1761 (N_1761,N_1278,N_1547);
nor U1762 (N_1762,N_1259,N_1289);
and U1763 (N_1763,N_1349,N_1331);
nor U1764 (N_1764,N_1525,N_1270);
nor U1765 (N_1765,N_1291,N_1466);
nor U1766 (N_1766,N_1459,N_1375);
and U1767 (N_1767,N_1514,N_1277);
or U1768 (N_1768,N_1425,N_1305);
nand U1769 (N_1769,N_1413,N_1496);
or U1770 (N_1770,N_1252,N_1528);
or U1771 (N_1771,N_1585,N_1488);
and U1772 (N_1772,N_1500,N_1239);
nand U1773 (N_1773,N_1209,N_1208);
or U1774 (N_1774,N_1441,N_1594);
nand U1775 (N_1775,N_1415,N_1564);
xnor U1776 (N_1776,N_1536,N_1485);
nor U1777 (N_1777,N_1581,N_1350);
nor U1778 (N_1778,N_1329,N_1224);
nor U1779 (N_1779,N_1593,N_1205);
or U1780 (N_1780,N_1576,N_1336);
xor U1781 (N_1781,N_1303,N_1544);
xnor U1782 (N_1782,N_1347,N_1297);
and U1783 (N_1783,N_1274,N_1217);
nand U1784 (N_1784,N_1560,N_1210);
and U1785 (N_1785,N_1377,N_1426);
nor U1786 (N_1786,N_1513,N_1591);
or U1787 (N_1787,N_1232,N_1430);
xor U1788 (N_1788,N_1416,N_1493);
and U1789 (N_1789,N_1200,N_1590);
nand U1790 (N_1790,N_1299,N_1531);
nand U1791 (N_1791,N_1399,N_1474);
and U1792 (N_1792,N_1244,N_1471);
and U1793 (N_1793,N_1492,N_1551);
or U1794 (N_1794,N_1417,N_1499);
and U1795 (N_1795,N_1325,N_1390);
or U1796 (N_1796,N_1483,N_1348);
nand U1797 (N_1797,N_1262,N_1469);
nor U1798 (N_1798,N_1561,N_1256);
nand U1799 (N_1799,N_1382,N_1369);
xor U1800 (N_1800,N_1496,N_1504);
nand U1801 (N_1801,N_1417,N_1579);
nor U1802 (N_1802,N_1258,N_1456);
nand U1803 (N_1803,N_1326,N_1286);
or U1804 (N_1804,N_1304,N_1531);
nand U1805 (N_1805,N_1222,N_1343);
nand U1806 (N_1806,N_1431,N_1235);
xnor U1807 (N_1807,N_1238,N_1333);
nor U1808 (N_1808,N_1520,N_1487);
or U1809 (N_1809,N_1522,N_1561);
or U1810 (N_1810,N_1360,N_1487);
nor U1811 (N_1811,N_1325,N_1505);
and U1812 (N_1812,N_1598,N_1389);
nand U1813 (N_1813,N_1406,N_1590);
nor U1814 (N_1814,N_1246,N_1444);
xor U1815 (N_1815,N_1340,N_1525);
xor U1816 (N_1816,N_1276,N_1464);
nor U1817 (N_1817,N_1561,N_1354);
or U1818 (N_1818,N_1461,N_1272);
nand U1819 (N_1819,N_1334,N_1460);
xnor U1820 (N_1820,N_1466,N_1299);
and U1821 (N_1821,N_1478,N_1474);
and U1822 (N_1822,N_1462,N_1444);
nor U1823 (N_1823,N_1565,N_1536);
and U1824 (N_1824,N_1325,N_1343);
or U1825 (N_1825,N_1558,N_1325);
or U1826 (N_1826,N_1210,N_1216);
nor U1827 (N_1827,N_1508,N_1424);
or U1828 (N_1828,N_1280,N_1545);
or U1829 (N_1829,N_1469,N_1405);
or U1830 (N_1830,N_1567,N_1412);
nor U1831 (N_1831,N_1335,N_1216);
and U1832 (N_1832,N_1248,N_1533);
or U1833 (N_1833,N_1462,N_1453);
nor U1834 (N_1834,N_1525,N_1418);
nor U1835 (N_1835,N_1266,N_1410);
xnor U1836 (N_1836,N_1248,N_1377);
xnor U1837 (N_1837,N_1256,N_1225);
nor U1838 (N_1838,N_1234,N_1290);
nand U1839 (N_1839,N_1367,N_1208);
and U1840 (N_1840,N_1484,N_1518);
and U1841 (N_1841,N_1426,N_1406);
xnor U1842 (N_1842,N_1296,N_1391);
xnor U1843 (N_1843,N_1466,N_1221);
or U1844 (N_1844,N_1411,N_1465);
and U1845 (N_1845,N_1422,N_1565);
xor U1846 (N_1846,N_1500,N_1219);
nand U1847 (N_1847,N_1552,N_1359);
nand U1848 (N_1848,N_1543,N_1439);
or U1849 (N_1849,N_1215,N_1323);
and U1850 (N_1850,N_1565,N_1248);
and U1851 (N_1851,N_1279,N_1596);
nor U1852 (N_1852,N_1345,N_1529);
nor U1853 (N_1853,N_1265,N_1466);
or U1854 (N_1854,N_1305,N_1338);
and U1855 (N_1855,N_1554,N_1282);
nor U1856 (N_1856,N_1459,N_1215);
nor U1857 (N_1857,N_1232,N_1505);
or U1858 (N_1858,N_1485,N_1236);
xor U1859 (N_1859,N_1288,N_1313);
or U1860 (N_1860,N_1572,N_1292);
and U1861 (N_1861,N_1532,N_1285);
and U1862 (N_1862,N_1236,N_1249);
or U1863 (N_1863,N_1583,N_1236);
xor U1864 (N_1864,N_1284,N_1257);
and U1865 (N_1865,N_1281,N_1351);
or U1866 (N_1866,N_1323,N_1556);
xor U1867 (N_1867,N_1293,N_1271);
and U1868 (N_1868,N_1474,N_1235);
xor U1869 (N_1869,N_1276,N_1452);
nand U1870 (N_1870,N_1259,N_1313);
and U1871 (N_1871,N_1436,N_1510);
nand U1872 (N_1872,N_1399,N_1367);
nor U1873 (N_1873,N_1420,N_1347);
nand U1874 (N_1874,N_1342,N_1250);
nand U1875 (N_1875,N_1499,N_1528);
or U1876 (N_1876,N_1277,N_1273);
nor U1877 (N_1877,N_1315,N_1246);
xnor U1878 (N_1878,N_1390,N_1399);
or U1879 (N_1879,N_1380,N_1292);
xor U1880 (N_1880,N_1295,N_1376);
nand U1881 (N_1881,N_1262,N_1409);
or U1882 (N_1882,N_1540,N_1267);
or U1883 (N_1883,N_1320,N_1485);
xnor U1884 (N_1884,N_1474,N_1291);
xnor U1885 (N_1885,N_1563,N_1552);
and U1886 (N_1886,N_1516,N_1377);
xor U1887 (N_1887,N_1587,N_1246);
nor U1888 (N_1888,N_1483,N_1550);
xor U1889 (N_1889,N_1383,N_1489);
and U1890 (N_1890,N_1306,N_1213);
or U1891 (N_1891,N_1449,N_1280);
nor U1892 (N_1892,N_1221,N_1257);
and U1893 (N_1893,N_1598,N_1309);
or U1894 (N_1894,N_1388,N_1504);
and U1895 (N_1895,N_1495,N_1550);
nand U1896 (N_1896,N_1328,N_1238);
and U1897 (N_1897,N_1306,N_1260);
xor U1898 (N_1898,N_1517,N_1500);
xnor U1899 (N_1899,N_1305,N_1508);
or U1900 (N_1900,N_1394,N_1500);
nand U1901 (N_1901,N_1587,N_1285);
xnor U1902 (N_1902,N_1229,N_1236);
and U1903 (N_1903,N_1470,N_1456);
nor U1904 (N_1904,N_1227,N_1415);
xnor U1905 (N_1905,N_1293,N_1541);
or U1906 (N_1906,N_1499,N_1415);
or U1907 (N_1907,N_1332,N_1422);
nand U1908 (N_1908,N_1573,N_1308);
and U1909 (N_1909,N_1379,N_1374);
nor U1910 (N_1910,N_1343,N_1452);
and U1911 (N_1911,N_1526,N_1390);
nor U1912 (N_1912,N_1302,N_1375);
and U1913 (N_1913,N_1340,N_1558);
xnor U1914 (N_1914,N_1247,N_1326);
and U1915 (N_1915,N_1207,N_1215);
and U1916 (N_1916,N_1216,N_1390);
and U1917 (N_1917,N_1262,N_1561);
nand U1918 (N_1918,N_1574,N_1493);
nor U1919 (N_1919,N_1320,N_1463);
xnor U1920 (N_1920,N_1493,N_1324);
nor U1921 (N_1921,N_1525,N_1431);
or U1922 (N_1922,N_1487,N_1462);
nor U1923 (N_1923,N_1573,N_1448);
or U1924 (N_1924,N_1524,N_1564);
and U1925 (N_1925,N_1290,N_1574);
xnor U1926 (N_1926,N_1468,N_1439);
nor U1927 (N_1927,N_1420,N_1220);
nand U1928 (N_1928,N_1402,N_1295);
or U1929 (N_1929,N_1552,N_1203);
xnor U1930 (N_1930,N_1500,N_1421);
nor U1931 (N_1931,N_1295,N_1421);
nand U1932 (N_1932,N_1481,N_1566);
nor U1933 (N_1933,N_1544,N_1376);
and U1934 (N_1934,N_1290,N_1301);
or U1935 (N_1935,N_1515,N_1448);
or U1936 (N_1936,N_1250,N_1440);
xor U1937 (N_1937,N_1475,N_1247);
nor U1938 (N_1938,N_1469,N_1582);
or U1939 (N_1939,N_1260,N_1206);
and U1940 (N_1940,N_1201,N_1453);
or U1941 (N_1941,N_1241,N_1578);
or U1942 (N_1942,N_1467,N_1585);
and U1943 (N_1943,N_1303,N_1485);
or U1944 (N_1944,N_1522,N_1466);
or U1945 (N_1945,N_1574,N_1484);
xnor U1946 (N_1946,N_1300,N_1483);
xor U1947 (N_1947,N_1269,N_1238);
or U1948 (N_1948,N_1556,N_1498);
nand U1949 (N_1949,N_1387,N_1364);
xor U1950 (N_1950,N_1211,N_1342);
nor U1951 (N_1951,N_1547,N_1297);
nor U1952 (N_1952,N_1563,N_1454);
nand U1953 (N_1953,N_1333,N_1343);
or U1954 (N_1954,N_1268,N_1438);
nor U1955 (N_1955,N_1526,N_1241);
xnor U1956 (N_1956,N_1487,N_1344);
nor U1957 (N_1957,N_1435,N_1376);
nor U1958 (N_1958,N_1475,N_1245);
nor U1959 (N_1959,N_1274,N_1397);
and U1960 (N_1960,N_1537,N_1207);
and U1961 (N_1961,N_1357,N_1260);
nor U1962 (N_1962,N_1358,N_1221);
nand U1963 (N_1963,N_1432,N_1327);
nor U1964 (N_1964,N_1354,N_1401);
and U1965 (N_1965,N_1244,N_1277);
or U1966 (N_1966,N_1580,N_1236);
or U1967 (N_1967,N_1401,N_1494);
and U1968 (N_1968,N_1222,N_1455);
nand U1969 (N_1969,N_1546,N_1557);
nor U1970 (N_1970,N_1313,N_1339);
nor U1971 (N_1971,N_1320,N_1474);
nand U1972 (N_1972,N_1278,N_1517);
nor U1973 (N_1973,N_1359,N_1429);
xnor U1974 (N_1974,N_1304,N_1246);
xor U1975 (N_1975,N_1508,N_1558);
nor U1976 (N_1976,N_1534,N_1330);
xor U1977 (N_1977,N_1462,N_1253);
nor U1978 (N_1978,N_1484,N_1563);
nand U1979 (N_1979,N_1360,N_1384);
nor U1980 (N_1980,N_1260,N_1210);
nand U1981 (N_1981,N_1555,N_1589);
xnor U1982 (N_1982,N_1298,N_1325);
nor U1983 (N_1983,N_1364,N_1505);
or U1984 (N_1984,N_1559,N_1345);
nor U1985 (N_1985,N_1322,N_1457);
xor U1986 (N_1986,N_1498,N_1372);
nand U1987 (N_1987,N_1373,N_1507);
or U1988 (N_1988,N_1488,N_1247);
xor U1989 (N_1989,N_1204,N_1368);
and U1990 (N_1990,N_1443,N_1341);
nand U1991 (N_1991,N_1364,N_1325);
nand U1992 (N_1992,N_1460,N_1340);
and U1993 (N_1993,N_1280,N_1366);
and U1994 (N_1994,N_1439,N_1224);
nand U1995 (N_1995,N_1264,N_1468);
xor U1996 (N_1996,N_1455,N_1281);
and U1997 (N_1997,N_1356,N_1308);
or U1998 (N_1998,N_1338,N_1510);
nor U1999 (N_1999,N_1318,N_1488);
nand U2000 (N_2000,N_1893,N_1858);
or U2001 (N_2001,N_1660,N_1972);
or U2002 (N_2002,N_1819,N_1673);
or U2003 (N_2003,N_1759,N_1918);
nand U2004 (N_2004,N_1715,N_1605);
nor U2005 (N_2005,N_1929,N_1820);
nor U2006 (N_2006,N_1821,N_1900);
and U2007 (N_2007,N_1609,N_1762);
nand U2008 (N_2008,N_1919,N_1904);
xnor U2009 (N_2009,N_1914,N_1978);
nor U2010 (N_2010,N_1936,N_1777);
and U2011 (N_2011,N_1963,N_1780);
and U2012 (N_2012,N_1808,N_1686);
or U2013 (N_2013,N_1846,N_1903);
xor U2014 (N_2014,N_1735,N_1908);
and U2015 (N_2015,N_1922,N_1631);
or U2016 (N_2016,N_1977,N_1807);
nand U2017 (N_2017,N_1694,N_1614);
or U2018 (N_2018,N_1882,N_1770);
xor U2019 (N_2019,N_1696,N_1848);
nand U2020 (N_2020,N_1647,N_1749);
or U2021 (N_2021,N_1782,N_1776);
nor U2022 (N_2022,N_1994,N_1864);
or U2023 (N_2023,N_1991,N_1910);
nor U2024 (N_2024,N_1973,N_1716);
or U2025 (N_2025,N_1877,N_1608);
or U2026 (N_2026,N_1956,N_1729);
xor U2027 (N_2027,N_1630,N_1906);
nor U2028 (N_2028,N_1932,N_1946);
and U2029 (N_2029,N_1815,N_1911);
xor U2030 (N_2030,N_1705,N_1612);
nor U2031 (N_2031,N_1933,N_1969);
xnor U2032 (N_2032,N_1623,N_1832);
and U2033 (N_2033,N_1600,N_1618);
or U2034 (N_2034,N_1721,N_1666);
and U2035 (N_2035,N_1857,N_1624);
nand U2036 (N_2036,N_1649,N_1681);
and U2037 (N_2037,N_1615,N_1634);
nand U2038 (N_2038,N_1747,N_1785);
and U2039 (N_2039,N_1650,N_1960);
nor U2040 (N_2040,N_1632,N_1626);
xnor U2041 (N_2041,N_1713,N_1629);
and U2042 (N_2042,N_1986,N_1703);
nand U2043 (N_2043,N_1739,N_1641);
and U2044 (N_2044,N_1949,N_1720);
and U2045 (N_2045,N_1794,N_1708);
nand U2046 (N_2046,N_1635,N_1826);
nor U2047 (N_2047,N_1775,N_1921);
nand U2048 (N_2048,N_1773,N_1702);
and U2049 (N_2049,N_1855,N_1862);
xnor U2050 (N_2050,N_1841,N_1723);
nand U2051 (N_2051,N_1889,N_1913);
or U2052 (N_2052,N_1709,N_1684);
nand U2053 (N_2053,N_1825,N_1707);
nor U2054 (N_2054,N_1719,N_1627);
or U2055 (N_2055,N_1912,N_1812);
xor U2056 (N_2056,N_1831,N_1697);
or U2057 (N_2057,N_1726,N_1845);
xnor U2058 (N_2058,N_1804,N_1685);
or U2059 (N_2059,N_1766,N_1805);
or U2060 (N_2060,N_1644,N_1866);
and U2061 (N_2061,N_1669,N_1665);
and U2062 (N_2062,N_1863,N_1836);
xnor U2063 (N_2063,N_1645,N_1727);
and U2064 (N_2064,N_1730,N_1757);
and U2065 (N_2065,N_1690,N_1602);
and U2066 (N_2066,N_1606,N_1689);
or U2067 (N_2067,N_1789,N_1951);
nand U2068 (N_2068,N_1931,N_1989);
nor U2069 (N_2069,N_1851,N_1881);
and U2070 (N_2070,N_1633,N_1971);
nor U2071 (N_2071,N_1965,N_1661);
or U2072 (N_2072,N_1700,N_1979);
and U2073 (N_2073,N_1717,N_1616);
xnor U2074 (N_2074,N_1695,N_1687);
nand U2075 (N_2075,N_1983,N_1966);
or U2076 (N_2076,N_1682,N_1976);
nor U2077 (N_2077,N_1810,N_1625);
or U2078 (N_2078,N_1704,N_1842);
or U2079 (N_2079,N_1891,N_1743);
nand U2080 (N_2080,N_1651,N_1806);
and U2081 (N_2081,N_1886,N_1742);
xor U2082 (N_2082,N_1835,N_1924);
xor U2083 (N_2083,N_1763,N_1672);
or U2084 (N_2084,N_1896,N_1740);
nand U2085 (N_2085,N_1917,N_1987);
or U2086 (N_2086,N_1797,N_1993);
xnor U2087 (N_2087,N_1957,N_1788);
or U2088 (N_2088,N_1736,N_1916);
nor U2089 (N_2089,N_1679,N_1664);
or U2090 (N_2090,N_1867,N_1947);
and U2091 (N_2091,N_1668,N_1722);
nor U2092 (N_2092,N_1659,N_1756);
nand U2093 (N_2093,N_1827,N_1905);
and U2094 (N_2094,N_1646,N_1818);
and U2095 (N_2095,N_1907,N_1754);
nor U2096 (N_2096,N_1784,N_1868);
and U2097 (N_2097,N_1793,N_1823);
xor U2098 (N_2098,N_1968,N_1786);
and U2099 (N_2099,N_1676,N_1871);
nor U2100 (N_2100,N_1648,N_1699);
nand U2101 (N_2101,N_1928,N_1755);
nor U2102 (N_2102,N_1945,N_1767);
and U2103 (N_2103,N_1760,N_1996);
nor U2104 (N_2104,N_1604,N_1725);
nor U2105 (N_2105,N_1950,N_1753);
or U2106 (N_2106,N_1942,N_1887);
xor U2107 (N_2107,N_1890,N_1909);
xor U2108 (N_2108,N_1714,N_1964);
nand U2109 (N_2109,N_1779,N_1758);
nand U2110 (N_2110,N_1675,N_1860);
or U2111 (N_2111,N_1828,N_1940);
nor U2112 (N_2112,N_1761,N_1822);
nand U2113 (N_2113,N_1741,N_1601);
nand U2114 (N_2114,N_1698,N_1621);
nand U2115 (N_2115,N_1837,N_1653);
nor U2116 (N_2116,N_1856,N_1670);
xor U2117 (N_2117,N_1975,N_1892);
nor U2118 (N_2118,N_1652,N_1640);
or U2119 (N_2119,N_1674,N_1817);
nand U2120 (N_2120,N_1829,N_1952);
nand U2121 (N_2121,N_1934,N_1671);
nor U2122 (N_2122,N_1967,N_1954);
and U2123 (N_2123,N_1751,N_1944);
and U2124 (N_2124,N_1691,N_1953);
nor U2125 (N_2125,N_1875,N_1622);
nor U2126 (N_2126,N_1885,N_1998);
nor U2127 (N_2127,N_1870,N_1710);
nand U2128 (N_2128,N_1611,N_1958);
nor U2129 (N_2129,N_1738,N_1748);
or U2130 (N_2130,N_1955,N_1902);
nand U2131 (N_2131,N_1657,N_1799);
or U2132 (N_2132,N_1992,N_1915);
or U2133 (N_2133,N_1844,N_1795);
nor U2134 (N_2134,N_1658,N_1920);
xor U2135 (N_2135,N_1849,N_1667);
nor U2136 (N_2136,N_1744,N_1850);
and U2137 (N_2137,N_1617,N_1791);
nand U2138 (N_2138,N_1603,N_1880);
and U2139 (N_2139,N_1796,N_1833);
nor U2140 (N_2140,N_1637,N_1999);
and U2141 (N_2141,N_1607,N_1774);
nand U2142 (N_2142,N_1814,N_1643);
xor U2143 (N_2143,N_1701,N_1663);
nand U2144 (N_2144,N_1878,N_1772);
and U2145 (N_2145,N_1731,N_1765);
and U2146 (N_2146,N_1959,N_1824);
nand U2147 (N_2147,N_1688,N_1656);
or U2148 (N_2148,N_1980,N_1926);
and U2149 (N_2149,N_1984,N_1613);
nor U2150 (N_2150,N_1988,N_1781);
nor U2151 (N_2151,N_1840,N_1677);
or U2152 (N_2152,N_1974,N_1733);
nor U2153 (N_2153,N_1899,N_1732);
nand U2154 (N_2154,N_1771,N_1970);
xnor U2155 (N_2155,N_1941,N_1706);
nand U2156 (N_2156,N_1874,N_1962);
xnor U2157 (N_2157,N_1724,N_1752);
nor U2158 (N_2158,N_1711,N_1927);
nor U2159 (N_2159,N_1680,N_1683);
nor U2160 (N_2160,N_1873,N_1655);
nand U2161 (N_2161,N_1925,N_1990);
or U2162 (N_2162,N_1935,N_1783);
or U2163 (N_2163,N_1839,N_1838);
nand U2164 (N_2164,N_1939,N_1718);
and U2165 (N_2165,N_1662,N_1901);
and U2166 (N_2166,N_1995,N_1746);
xnor U2167 (N_2167,N_1768,N_1737);
and U2168 (N_2168,N_1619,N_1861);
nor U2169 (N_2169,N_1897,N_1865);
xor U2170 (N_2170,N_1693,N_1859);
nand U2171 (N_2171,N_1678,N_1883);
nor U2172 (N_2172,N_1830,N_1790);
nand U2173 (N_2173,N_1734,N_1620);
xnor U2174 (N_2174,N_1876,N_1778);
xnor U2175 (N_2175,N_1628,N_1801);
or U2176 (N_2176,N_1764,N_1638);
or U2177 (N_2177,N_1943,N_1692);
xor U2178 (N_2178,N_1712,N_1843);
xor U2179 (N_2179,N_1894,N_1847);
xnor U2180 (N_2180,N_1898,N_1872);
and U2181 (N_2181,N_1853,N_1800);
nand U2182 (N_2182,N_1961,N_1895);
or U2183 (N_2183,N_1639,N_1787);
nor U2184 (N_2184,N_1869,N_1982);
or U2185 (N_2185,N_1816,N_1981);
and U2186 (N_2186,N_1769,N_1923);
and U2187 (N_2187,N_1948,N_1803);
nand U2188 (N_2188,N_1834,N_1642);
nand U2189 (N_2189,N_1930,N_1728);
nor U2190 (N_2190,N_1798,N_1884);
nor U2191 (N_2191,N_1888,N_1813);
and U2192 (N_2192,N_1852,N_1636);
nand U2193 (N_2193,N_1879,N_1610);
and U2194 (N_2194,N_1985,N_1809);
nand U2195 (N_2195,N_1854,N_1811);
and U2196 (N_2196,N_1792,N_1745);
nor U2197 (N_2197,N_1654,N_1802);
nor U2198 (N_2198,N_1750,N_1997);
and U2199 (N_2199,N_1937,N_1938);
xnor U2200 (N_2200,N_1875,N_1989);
nand U2201 (N_2201,N_1819,N_1728);
nor U2202 (N_2202,N_1738,N_1693);
nor U2203 (N_2203,N_1781,N_1849);
and U2204 (N_2204,N_1711,N_1731);
xor U2205 (N_2205,N_1682,N_1979);
and U2206 (N_2206,N_1711,N_1695);
nor U2207 (N_2207,N_1845,N_1692);
nand U2208 (N_2208,N_1751,N_1788);
nand U2209 (N_2209,N_1844,N_1838);
nand U2210 (N_2210,N_1609,N_1802);
nor U2211 (N_2211,N_1738,N_1715);
and U2212 (N_2212,N_1804,N_1731);
or U2213 (N_2213,N_1615,N_1612);
nand U2214 (N_2214,N_1782,N_1932);
nor U2215 (N_2215,N_1656,N_1676);
nor U2216 (N_2216,N_1749,N_1750);
xor U2217 (N_2217,N_1782,N_1962);
or U2218 (N_2218,N_1882,N_1962);
nor U2219 (N_2219,N_1794,N_1640);
nor U2220 (N_2220,N_1746,N_1924);
xnor U2221 (N_2221,N_1959,N_1650);
nor U2222 (N_2222,N_1848,N_1907);
nor U2223 (N_2223,N_1684,N_1867);
and U2224 (N_2224,N_1844,N_1711);
nor U2225 (N_2225,N_1726,N_1832);
and U2226 (N_2226,N_1743,N_1964);
or U2227 (N_2227,N_1834,N_1765);
nor U2228 (N_2228,N_1714,N_1771);
or U2229 (N_2229,N_1946,N_1867);
or U2230 (N_2230,N_1980,N_1986);
nor U2231 (N_2231,N_1917,N_1875);
nand U2232 (N_2232,N_1856,N_1870);
nor U2233 (N_2233,N_1841,N_1684);
and U2234 (N_2234,N_1756,N_1981);
xor U2235 (N_2235,N_1763,N_1979);
xnor U2236 (N_2236,N_1958,N_1841);
and U2237 (N_2237,N_1987,N_1763);
nand U2238 (N_2238,N_1781,N_1882);
nor U2239 (N_2239,N_1965,N_1959);
nor U2240 (N_2240,N_1985,N_1764);
xnor U2241 (N_2241,N_1875,N_1758);
xor U2242 (N_2242,N_1746,N_1909);
nand U2243 (N_2243,N_1684,N_1813);
xnor U2244 (N_2244,N_1896,N_1755);
xor U2245 (N_2245,N_1915,N_1638);
nor U2246 (N_2246,N_1804,N_1713);
or U2247 (N_2247,N_1950,N_1746);
nand U2248 (N_2248,N_1766,N_1902);
or U2249 (N_2249,N_1842,N_1953);
nor U2250 (N_2250,N_1883,N_1757);
or U2251 (N_2251,N_1877,N_1657);
nand U2252 (N_2252,N_1902,N_1684);
nor U2253 (N_2253,N_1930,N_1662);
and U2254 (N_2254,N_1765,N_1686);
and U2255 (N_2255,N_1685,N_1796);
xnor U2256 (N_2256,N_1901,N_1644);
nor U2257 (N_2257,N_1982,N_1791);
xor U2258 (N_2258,N_1639,N_1960);
nor U2259 (N_2259,N_1952,N_1716);
or U2260 (N_2260,N_1645,N_1919);
or U2261 (N_2261,N_1678,N_1645);
xor U2262 (N_2262,N_1836,N_1689);
and U2263 (N_2263,N_1763,N_1743);
and U2264 (N_2264,N_1630,N_1603);
xnor U2265 (N_2265,N_1853,N_1818);
nor U2266 (N_2266,N_1618,N_1856);
nand U2267 (N_2267,N_1607,N_1801);
nor U2268 (N_2268,N_1634,N_1917);
xor U2269 (N_2269,N_1775,N_1896);
nor U2270 (N_2270,N_1629,N_1737);
nor U2271 (N_2271,N_1783,N_1721);
nand U2272 (N_2272,N_1944,N_1908);
and U2273 (N_2273,N_1641,N_1705);
xor U2274 (N_2274,N_1837,N_1620);
or U2275 (N_2275,N_1617,N_1933);
nor U2276 (N_2276,N_1724,N_1718);
or U2277 (N_2277,N_1823,N_1910);
and U2278 (N_2278,N_1731,N_1791);
or U2279 (N_2279,N_1776,N_1834);
nand U2280 (N_2280,N_1826,N_1796);
and U2281 (N_2281,N_1993,N_1628);
nand U2282 (N_2282,N_1778,N_1988);
xor U2283 (N_2283,N_1990,N_1704);
nor U2284 (N_2284,N_1779,N_1625);
xnor U2285 (N_2285,N_1615,N_1818);
nor U2286 (N_2286,N_1778,N_1744);
nor U2287 (N_2287,N_1618,N_1622);
nor U2288 (N_2288,N_1700,N_1965);
nand U2289 (N_2289,N_1922,N_1984);
nor U2290 (N_2290,N_1655,N_1937);
xor U2291 (N_2291,N_1623,N_1602);
nand U2292 (N_2292,N_1902,N_1815);
xor U2293 (N_2293,N_1620,N_1823);
and U2294 (N_2294,N_1695,N_1904);
nand U2295 (N_2295,N_1792,N_1959);
nor U2296 (N_2296,N_1792,N_1852);
xor U2297 (N_2297,N_1853,N_1785);
xor U2298 (N_2298,N_1649,N_1733);
nand U2299 (N_2299,N_1699,N_1998);
nand U2300 (N_2300,N_1608,N_1791);
and U2301 (N_2301,N_1856,N_1666);
nor U2302 (N_2302,N_1690,N_1830);
nand U2303 (N_2303,N_1955,N_1863);
or U2304 (N_2304,N_1887,N_1636);
and U2305 (N_2305,N_1976,N_1886);
xnor U2306 (N_2306,N_1825,N_1938);
xnor U2307 (N_2307,N_1718,N_1876);
nor U2308 (N_2308,N_1661,N_1671);
nand U2309 (N_2309,N_1668,N_1794);
and U2310 (N_2310,N_1985,N_1826);
nand U2311 (N_2311,N_1726,N_1696);
and U2312 (N_2312,N_1980,N_1728);
or U2313 (N_2313,N_1895,N_1600);
and U2314 (N_2314,N_1654,N_1931);
and U2315 (N_2315,N_1744,N_1722);
xor U2316 (N_2316,N_1694,N_1670);
nor U2317 (N_2317,N_1684,N_1905);
xnor U2318 (N_2318,N_1661,N_1682);
nand U2319 (N_2319,N_1611,N_1690);
nor U2320 (N_2320,N_1869,N_1694);
and U2321 (N_2321,N_1791,N_1776);
nand U2322 (N_2322,N_1686,N_1718);
nor U2323 (N_2323,N_1622,N_1769);
nand U2324 (N_2324,N_1831,N_1852);
nor U2325 (N_2325,N_1803,N_1769);
nor U2326 (N_2326,N_1851,N_1984);
nand U2327 (N_2327,N_1624,N_1667);
and U2328 (N_2328,N_1789,N_1898);
nand U2329 (N_2329,N_1946,N_1784);
and U2330 (N_2330,N_1831,N_1649);
xnor U2331 (N_2331,N_1831,N_1886);
xor U2332 (N_2332,N_1810,N_1705);
and U2333 (N_2333,N_1892,N_1639);
xnor U2334 (N_2334,N_1985,N_1842);
nand U2335 (N_2335,N_1970,N_1743);
nand U2336 (N_2336,N_1822,N_1622);
xor U2337 (N_2337,N_1989,N_1711);
xnor U2338 (N_2338,N_1767,N_1762);
or U2339 (N_2339,N_1838,N_1744);
nor U2340 (N_2340,N_1930,N_1802);
xor U2341 (N_2341,N_1825,N_1885);
nand U2342 (N_2342,N_1906,N_1965);
or U2343 (N_2343,N_1933,N_1776);
nand U2344 (N_2344,N_1609,N_1755);
nor U2345 (N_2345,N_1780,N_1662);
nor U2346 (N_2346,N_1934,N_1617);
nor U2347 (N_2347,N_1812,N_1784);
nand U2348 (N_2348,N_1909,N_1854);
xor U2349 (N_2349,N_1672,N_1928);
nor U2350 (N_2350,N_1992,N_1969);
or U2351 (N_2351,N_1730,N_1637);
nand U2352 (N_2352,N_1718,N_1911);
or U2353 (N_2353,N_1924,N_1973);
or U2354 (N_2354,N_1648,N_1732);
nand U2355 (N_2355,N_1986,N_1950);
or U2356 (N_2356,N_1701,N_1658);
or U2357 (N_2357,N_1723,N_1718);
xor U2358 (N_2358,N_1690,N_1685);
nand U2359 (N_2359,N_1809,N_1924);
xor U2360 (N_2360,N_1780,N_1658);
or U2361 (N_2361,N_1650,N_1936);
xor U2362 (N_2362,N_1780,N_1670);
nand U2363 (N_2363,N_1964,N_1961);
nor U2364 (N_2364,N_1648,N_1632);
and U2365 (N_2365,N_1884,N_1952);
and U2366 (N_2366,N_1786,N_1789);
nor U2367 (N_2367,N_1687,N_1710);
and U2368 (N_2368,N_1892,N_1685);
nand U2369 (N_2369,N_1850,N_1739);
xnor U2370 (N_2370,N_1745,N_1695);
nor U2371 (N_2371,N_1974,N_1802);
nor U2372 (N_2372,N_1866,N_1876);
xor U2373 (N_2373,N_1895,N_1938);
or U2374 (N_2374,N_1675,N_1712);
xor U2375 (N_2375,N_1995,N_1952);
nor U2376 (N_2376,N_1924,N_1860);
nor U2377 (N_2377,N_1927,N_1818);
xor U2378 (N_2378,N_1730,N_1818);
or U2379 (N_2379,N_1801,N_1985);
and U2380 (N_2380,N_1774,N_1622);
or U2381 (N_2381,N_1930,N_1678);
nand U2382 (N_2382,N_1708,N_1881);
nand U2383 (N_2383,N_1919,N_1773);
xor U2384 (N_2384,N_1784,N_1914);
or U2385 (N_2385,N_1865,N_1876);
xnor U2386 (N_2386,N_1893,N_1829);
or U2387 (N_2387,N_1874,N_1678);
nand U2388 (N_2388,N_1605,N_1891);
xor U2389 (N_2389,N_1842,N_1644);
or U2390 (N_2390,N_1981,N_1746);
nand U2391 (N_2391,N_1847,N_1783);
or U2392 (N_2392,N_1951,N_1757);
nor U2393 (N_2393,N_1788,N_1949);
nor U2394 (N_2394,N_1604,N_1713);
nor U2395 (N_2395,N_1700,N_1914);
xor U2396 (N_2396,N_1745,N_1878);
or U2397 (N_2397,N_1808,N_1747);
and U2398 (N_2398,N_1600,N_1954);
nand U2399 (N_2399,N_1926,N_1796);
nand U2400 (N_2400,N_2125,N_2291);
xnor U2401 (N_2401,N_2123,N_2287);
and U2402 (N_2402,N_2087,N_2134);
or U2403 (N_2403,N_2062,N_2336);
or U2404 (N_2404,N_2199,N_2014);
and U2405 (N_2405,N_2396,N_2360);
and U2406 (N_2406,N_2350,N_2247);
or U2407 (N_2407,N_2117,N_2207);
xor U2408 (N_2408,N_2246,N_2078);
nor U2409 (N_2409,N_2046,N_2222);
and U2410 (N_2410,N_2118,N_2235);
nor U2411 (N_2411,N_2334,N_2254);
nand U2412 (N_2412,N_2327,N_2294);
nand U2413 (N_2413,N_2156,N_2077);
xor U2414 (N_2414,N_2160,N_2065);
and U2415 (N_2415,N_2371,N_2169);
nor U2416 (N_2416,N_2231,N_2007);
or U2417 (N_2417,N_2075,N_2299);
nand U2418 (N_2418,N_2001,N_2303);
nand U2419 (N_2419,N_2094,N_2052);
nand U2420 (N_2420,N_2274,N_2086);
nand U2421 (N_2421,N_2027,N_2047);
xor U2422 (N_2422,N_2184,N_2079);
nand U2423 (N_2423,N_2127,N_2016);
xor U2424 (N_2424,N_2313,N_2102);
nor U2425 (N_2425,N_2392,N_2385);
or U2426 (N_2426,N_2120,N_2048);
or U2427 (N_2427,N_2204,N_2167);
or U2428 (N_2428,N_2149,N_2017);
xor U2429 (N_2429,N_2384,N_2076);
or U2430 (N_2430,N_2105,N_2279);
and U2431 (N_2431,N_2292,N_2059);
nor U2432 (N_2432,N_2053,N_2343);
or U2433 (N_2433,N_2122,N_2245);
nor U2434 (N_2434,N_2280,N_2262);
nor U2435 (N_2435,N_2365,N_2352);
and U2436 (N_2436,N_2181,N_2203);
and U2437 (N_2437,N_2244,N_2234);
and U2438 (N_2438,N_2057,N_2000);
and U2439 (N_2439,N_2219,N_2084);
nand U2440 (N_2440,N_2081,N_2377);
xor U2441 (N_2441,N_2172,N_2314);
nand U2442 (N_2442,N_2186,N_2183);
and U2443 (N_2443,N_2364,N_2055);
and U2444 (N_2444,N_2383,N_2178);
or U2445 (N_2445,N_2237,N_2300);
nor U2446 (N_2446,N_2323,N_2020);
nor U2447 (N_2447,N_2296,N_2273);
xnor U2448 (N_2448,N_2088,N_2345);
and U2449 (N_2449,N_2312,N_2354);
nor U2450 (N_2450,N_2180,N_2179);
xor U2451 (N_2451,N_2215,N_2265);
or U2452 (N_2452,N_2353,N_2216);
nand U2453 (N_2453,N_2316,N_2090);
nor U2454 (N_2454,N_2064,N_2010);
xor U2455 (N_2455,N_2011,N_2039);
or U2456 (N_2456,N_2286,N_2190);
and U2457 (N_2457,N_2242,N_2168);
nor U2458 (N_2458,N_2306,N_2356);
or U2459 (N_2459,N_2344,N_2259);
and U2460 (N_2460,N_2028,N_2302);
and U2461 (N_2461,N_2013,N_2326);
xnor U2462 (N_2462,N_2243,N_2285);
and U2463 (N_2463,N_2100,N_2034);
and U2464 (N_2464,N_2196,N_2391);
nor U2465 (N_2465,N_2269,N_2217);
and U2466 (N_2466,N_2171,N_2363);
and U2467 (N_2467,N_2139,N_2146);
and U2468 (N_2468,N_2157,N_2397);
or U2469 (N_2469,N_2348,N_2085);
or U2470 (N_2470,N_2281,N_2335);
or U2471 (N_2471,N_2275,N_2317);
xnor U2472 (N_2472,N_2095,N_2370);
or U2473 (N_2473,N_2188,N_2290);
nand U2474 (N_2474,N_2006,N_2126);
nor U2475 (N_2475,N_2319,N_2056);
xnor U2476 (N_2476,N_2256,N_2309);
and U2477 (N_2477,N_2250,N_2098);
xnor U2478 (N_2478,N_2096,N_2283);
and U2479 (N_2479,N_2340,N_2315);
or U2480 (N_2480,N_2241,N_2214);
nand U2481 (N_2481,N_2021,N_2266);
and U2482 (N_2482,N_2165,N_2147);
and U2483 (N_2483,N_2308,N_2240);
xor U2484 (N_2484,N_2387,N_2150);
and U2485 (N_2485,N_2282,N_2272);
nor U2486 (N_2486,N_2230,N_2136);
and U2487 (N_2487,N_2026,N_2239);
nand U2488 (N_2488,N_2128,N_2191);
nand U2489 (N_2489,N_2071,N_2398);
or U2490 (N_2490,N_2399,N_2394);
and U2491 (N_2491,N_2213,N_2012);
nand U2492 (N_2492,N_2093,N_2194);
and U2493 (N_2493,N_2263,N_2355);
and U2494 (N_2494,N_2267,N_2189);
nand U2495 (N_2495,N_2261,N_2375);
nor U2496 (N_2496,N_2025,N_2301);
xnor U2497 (N_2497,N_2103,N_2271);
and U2498 (N_2498,N_2041,N_2161);
or U2499 (N_2499,N_2163,N_2187);
xnor U2500 (N_2500,N_2320,N_2023);
nor U2501 (N_2501,N_2089,N_2101);
or U2502 (N_2502,N_2382,N_2332);
nand U2503 (N_2503,N_2192,N_2322);
or U2504 (N_2504,N_2284,N_2288);
nor U2505 (N_2505,N_2067,N_2009);
xor U2506 (N_2506,N_2257,N_2258);
xnor U2507 (N_2507,N_2137,N_2074);
nor U2508 (N_2508,N_2379,N_2307);
nor U2509 (N_2509,N_2135,N_2054);
and U2510 (N_2510,N_2200,N_2201);
xor U2511 (N_2511,N_2251,N_2174);
or U2512 (N_2512,N_2069,N_2050);
nor U2513 (N_2513,N_2182,N_2018);
xor U2514 (N_2514,N_2347,N_2226);
or U2515 (N_2515,N_2277,N_2107);
xor U2516 (N_2516,N_2121,N_2395);
nand U2517 (N_2517,N_2031,N_2212);
or U2518 (N_2518,N_2004,N_2293);
and U2519 (N_2519,N_2049,N_2115);
or U2520 (N_2520,N_2040,N_2276);
or U2521 (N_2521,N_2378,N_2268);
and U2522 (N_2522,N_2112,N_2373);
and U2523 (N_2523,N_2158,N_2130);
and U2524 (N_2524,N_2198,N_2061);
nor U2525 (N_2525,N_2119,N_2238);
or U2526 (N_2526,N_2328,N_2252);
or U2527 (N_2527,N_2386,N_2106);
and U2528 (N_2528,N_2145,N_2166);
and U2529 (N_2529,N_2357,N_2366);
or U2530 (N_2530,N_2393,N_2042);
and U2531 (N_2531,N_2232,N_2022);
and U2532 (N_2532,N_2133,N_2045);
nor U2533 (N_2533,N_2176,N_2037);
and U2534 (N_2534,N_2003,N_2109);
nand U2535 (N_2535,N_2140,N_2029);
or U2536 (N_2536,N_2083,N_2374);
nor U2537 (N_2537,N_2227,N_2051);
nand U2538 (N_2538,N_2116,N_2208);
and U2539 (N_2539,N_2082,N_2152);
xor U2540 (N_2540,N_2368,N_2177);
or U2541 (N_2541,N_2329,N_2380);
nor U2542 (N_2542,N_2361,N_2024);
nand U2543 (N_2543,N_2060,N_2058);
and U2544 (N_2544,N_2236,N_2225);
nor U2545 (N_2545,N_2249,N_2376);
nor U2546 (N_2546,N_2193,N_2185);
and U2547 (N_2547,N_2311,N_2030);
and U2548 (N_2548,N_2390,N_2143);
nand U2549 (N_2549,N_2202,N_2099);
or U2550 (N_2550,N_2164,N_2035);
xnor U2551 (N_2551,N_2223,N_2389);
or U2552 (N_2552,N_2091,N_2151);
or U2553 (N_2553,N_2295,N_2111);
or U2554 (N_2554,N_2367,N_2005);
and U2555 (N_2555,N_2297,N_2325);
nor U2556 (N_2556,N_2346,N_2142);
and U2557 (N_2557,N_2218,N_2066);
and U2558 (N_2558,N_2138,N_2233);
and U2559 (N_2559,N_2339,N_2063);
and U2560 (N_2560,N_2381,N_2369);
and U2561 (N_2561,N_2036,N_2092);
and U2562 (N_2562,N_2206,N_2362);
or U2563 (N_2563,N_2388,N_2304);
or U2564 (N_2564,N_2154,N_2337);
nor U2565 (N_2565,N_2211,N_2114);
nand U2566 (N_2566,N_2351,N_2068);
nand U2567 (N_2567,N_2072,N_2173);
nor U2568 (N_2568,N_2210,N_2110);
xor U2569 (N_2569,N_2015,N_2338);
or U2570 (N_2570,N_2175,N_2073);
or U2571 (N_2571,N_2170,N_2097);
and U2572 (N_2572,N_2318,N_2229);
xnor U2573 (N_2573,N_2321,N_2070);
xor U2574 (N_2574,N_2019,N_2108);
nor U2575 (N_2575,N_2159,N_2341);
nor U2576 (N_2576,N_2289,N_2260);
nor U2577 (N_2577,N_2298,N_2310);
nor U2578 (N_2578,N_2153,N_2221);
nand U2579 (N_2579,N_2195,N_2220);
nand U2580 (N_2580,N_2131,N_2032);
or U2581 (N_2581,N_2228,N_2129);
nand U2582 (N_2582,N_2124,N_2080);
nand U2583 (N_2583,N_2248,N_2324);
nand U2584 (N_2584,N_2038,N_2333);
and U2585 (N_2585,N_2255,N_2113);
nor U2586 (N_2586,N_2043,N_2264);
and U2587 (N_2587,N_2008,N_2342);
nor U2588 (N_2588,N_2104,N_2330);
nor U2589 (N_2589,N_2162,N_2224);
and U2590 (N_2590,N_2044,N_2358);
and U2591 (N_2591,N_2331,N_2305);
xnor U2592 (N_2592,N_2209,N_2002);
xor U2593 (N_2593,N_2253,N_2278);
nand U2594 (N_2594,N_2155,N_2197);
nor U2595 (N_2595,N_2144,N_2372);
nand U2596 (N_2596,N_2359,N_2033);
nor U2597 (N_2597,N_2148,N_2141);
or U2598 (N_2598,N_2205,N_2270);
xor U2599 (N_2599,N_2132,N_2349);
xor U2600 (N_2600,N_2264,N_2211);
and U2601 (N_2601,N_2071,N_2314);
nand U2602 (N_2602,N_2265,N_2391);
and U2603 (N_2603,N_2247,N_2105);
and U2604 (N_2604,N_2204,N_2245);
and U2605 (N_2605,N_2098,N_2125);
and U2606 (N_2606,N_2070,N_2296);
and U2607 (N_2607,N_2372,N_2054);
nand U2608 (N_2608,N_2050,N_2324);
nand U2609 (N_2609,N_2162,N_2392);
nor U2610 (N_2610,N_2088,N_2341);
nor U2611 (N_2611,N_2358,N_2180);
nor U2612 (N_2612,N_2020,N_2152);
nand U2613 (N_2613,N_2330,N_2165);
xnor U2614 (N_2614,N_2065,N_2096);
and U2615 (N_2615,N_2190,N_2355);
nand U2616 (N_2616,N_2362,N_2365);
and U2617 (N_2617,N_2048,N_2152);
xor U2618 (N_2618,N_2239,N_2010);
nor U2619 (N_2619,N_2113,N_2181);
and U2620 (N_2620,N_2152,N_2302);
nor U2621 (N_2621,N_2028,N_2290);
or U2622 (N_2622,N_2370,N_2074);
nor U2623 (N_2623,N_2161,N_2193);
and U2624 (N_2624,N_2035,N_2228);
or U2625 (N_2625,N_2087,N_2192);
and U2626 (N_2626,N_2346,N_2238);
xor U2627 (N_2627,N_2139,N_2156);
and U2628 (N_2628,N_2262,N_2111);
nor U2629 (N_2629,N_2249,N_2339);
or U2630 (N_2630,N_2049,N_2221);
nand U2631 (N_2631,N_2011,N_2275);
and U2632 (N_2632,N_2140,N_2273);
xnor U2633 (N_2633,N_2393,N_2208);
or U2634 (N_2634,N_2131,N_2041);
and U2635 (N_2635,N_2257,N_2371);
nand U2636 (N_2636,N_2107,N_2002);
xor U2637 (N_2637,N_2266,N_2090);
xor U2638 (N_2638,N_2267,N_2062);
and U2639 (N_2639,N_2253,N_2329);
nor U2640 (N_2640,N_2005,N_2153);
or U2641 (N_2641,N_2371,N_2086);
or U2642 (N_2642,N_2068,N_2273);
nand U2643 (N_2643,N_2179,N_2380);
nand U2644 (N_2644,N_2202,N_2362);
nand U2645 (N_2645,N_2393,N_2071);
xnor U2646 (N_2646,N_2268,N_2333);
and U2647 (N_2647,N_2389,N_2305);
nor U2648 (N_2648,N_2226,N_2117);
nor U2649 (N_2649,N_2244,N_2068);
nor U2650 (N_2650,N_2233,N_2137);
xnor U2651 (N_2651,N_2254,N_2377);
nand U2652 (N_2652,N_2174,N_2299);
and U2653 (N_2653,N_2395,N_2371);
nor U2654 (N_2654,N_2298,N_2038);
nand U2655 (N_2655,N_2320,N_2218);
xor U2656 (N_2656,N_2052,N_2193);
nand U2657 (N_2657,N_2343,N_2324);
or U2658 (N_2658,N_2066,N_2197);
xnor U2659 (N_2659,N_2333,N_2107);
or U2660 (N_2660,N_2351,N_2161);
and U2661 (N_2661,N_2283,N_2121);
or U2662 (N_2662,N_2076,N_2132);
and U2663 (N_2663,N_2112,N_2139);
xor U2664 (N_2664,N_2207,N_2070);
nor U2665 (N_2665,N_2095,N_2339);
xor U2666 (N_2666,N_2320,N_2268);
xnor U2667 (N_2667,N_2249,N_2395);
and U2668 (N_2668,N_2255,N_2272);
or U2669 (N_2669,N_2363,N_2368);
nor U2670 (N_2670,N_2256,N_2318);
or U2671 (N_2671,N_2343,N_2370);
xor U2672 (N_2672,N_2230,N_2357);
xnor U2673 (N_2673,N_2169,N_2297);
or U2674 (N_2674,N_2244,N_2057);
nand U2675 (N_2675,N_2395,N_2346);
nand U2676 (N_2676,N_2291,N_2296);
nand U2677 (N_2677,N_2322,N_2304);
or U2678 (N_2678,N_2291,N_2053);
xor U2679 (N_2679,N_2134,N_2126);
or U2680 (N_2680,N_2365,N_2060);
or U2681 (N_2681,N_2207,N_2076);
or U2682 (N_2682,N_2234,N_2175);
nand U2683 (N_2683,N_2066,N_2025);
or U2684 (N_2684,N_2264,N_2084);
nand U2685 (N_2685,N_2254,N_2172);
and U2686 (N_2686,N_2151,N_2087);
or U2687 (N_2687,N_2006,N_2397);
and U2688 (N_2688,N_2020,N_2147);
and U2689 (N_2689,N_2288,N_2193);
and U2690 (N_2690,N_2384,N_2285);
nand U2691 (N_2691,N_2051,N_2054);
nand U2692 (N_2692,N_2114,N_2261);
or U2693 (N_2693,N_2352,N_2276);
or U2694 (N_2694,N_2143,N_2337);
xor U2695 (N_2695,N_2174,N_2144);
nor U2696 (N_2696,N_2068,N_2306);
nand U2697 (N_2697,N_2042,N_2394);
nand U2698 (N_2698,N_2366,N_2031);
or U2699 (N_2699,N_2245,N_2263);
nand U2700 (N_2700,N_2002,N_2187);
or U2701 (N_2701,N_2392,N_2361);
or U2702 (N_2702,N_2069,N_2193);
nand U2703 (N_2703,N_2079,N_2181);
nand U2704 (N_2704,N_2350,N_2284);
nand U2705 (N_2705,N_2154,N_2348);
or U2706 (N_2706,N_2355,N_2269);
or U2707 (N_2707,N_2358,N_2331);
xor U2708 (N_2708,N_2323,N_2385);
nand U2709 (N_2709,N_2280,N_2223);
nor U2710 (N_2710,N_2352,N_2286);
nor U2711 (N_2711,N_2026,N_2110);
nor U2712 (N_2712,N_2228,N_2037);
xnor U2713 (N_2713,N_2249,N_2175);
and U2714 (N_2714,N_2336,N_2301);
or U2715 (N_2715,N_2202,N_2288);
and U2716 (N_2716,N_2385,N_2031);
xnor U2717 (N_2717,N_2262,N_2195);
or U2718 (N_2718,N_2194,N_2133);
and U2719 (N_2719,N_2320,N_2278);
and U2720 (N_2720,N_2245,N_2235);
and U2721 (N_2721,N_2291,N_2325);
nor U2722 (N_2722,N_2187,N_2016);
nand U2723 (N_2723,N_2233,N_2305);
xnor U2724 (N_2724,N_2351,N_2101);
xnor U2725 (N_2725,N_2142,N_2353);
nor U2726 (N_2726,N_2049,N_2320);
nand U2727 (N_2727,N_2133,N_2073);
or U2728 (N_2728,N_2314,N_2109);
nand U2729 (N_2729,N_2200,N_2179);
nor U2730 (N_2730,N_2125,N_2107);
xnor U2731 (N_2731,N_2128,N_2020);
xnor U2732 (N_2732,N_2103,N_2390);
or U2733 (N_2733,N_2104,N_2394);
nor U2734 (N_2734,N_2332,N_2288);
xnor U2735 (N_2735,N_2023,N_2299);
nor U2736 (N_2736,N_2049,N_2283);
nand U2737 (N_2737,N_2396,N_2203);
xnor U2738 (N_2738,N_2392,N_2195);
or U2739 (N_2739,N_2139,N_2093);
nor U2740 (N_2740,N_2144,N_2390);
nand U2741 (N_2741,N_2244,N_2166);
and U2742 (N_2742,N_2032,N_2076);
and U2743 (N_2743,N_2276,N_2348);
nor U2744 (N_2744,N_2203,N_2215);
nor U2745 (N_2745,N_2195,N_2079);
and U2746 (N_2746,N_2345,N_2387);
and U2747 (N_2747,N_2182,N_2317);
nand U2748 (N_2748,N_2136,N_2204);
nand U2749 (N_2749,N_2009,N_2369);
and U2750 (N_2750,N_2274,N_2074);
nand U2751 (N_2751,N_2292,N_2076);
xnor U2752 (N_2752,N_2303,N_2073);
xnor U2753 (N_2753,N_2169,N_2178);
nor U2754 (N_2754,N_2015,N_2309);
nand U2755 (N_2755,N_2381,N_2213);
or U2756 (N_2756,N_2121,N_2261);
nor U2757 (N_2757,N_2195,N_2173);
and U2758 (N_2758,N_2168,N_2317);
and U2759 (N_2759,N_2395,N_2399);
and U2760 (N_2760,N_2273,N_2366);
and U2761 (N_2761,N_2362,N_2285);
nand U2762 (N_2762,N_2195,N_2159);
xnor U2763 (N_2763,N_2174,N_2306);
or U2764 (N_2764,N_2353,N_2072);
and U2765 (N_2765,N_2138,N_2015);
and U2766 (N_2766,N_2305,N_2304);
or U2767 (N_2767,N_2157,N_2088);
nand U2768 (N_2768,N_2394,N_2366);
or U2769 (N_2769,N_2205,N_2101);
nand U2770 (N_2770,N_2279,N_2389);
xor U2771 (N_2771,N_2116,N_2163);
and U2772 (N_2772,N_2130,N_2238);
and U2773 (N_2773,N_2199,N_2217);
nand U2774 (N_2774,N_2111,N_2100);
or U2775 (N_2775,N_2216,N_2262);
or U2776 (N_2776,N_2376,N_2208);
nand U2777 (N_2777,N_2063,N_2135);
and U2778 (N_2778,N_2048,N_2255);
nor U2779 (N_2779,N_2053,N_2337);
nand U2780 (N_2780,N_2293,N_2097);
nand U2781 (N_2781,N_2200,N_2117);
nand U2782 (N_2782,N_2383,N_2209);
or U2783 (N_2783,N_2327,N_2080);
or U2784 (N_2784,N_2343,N_2180);
nand U2785 (N_2785,N_2260,N_2059);
and U2786 (N_2786,N_2096,N_2106);
nand U2787 (N_2787,N_2146,N_2185);
and U2788 (N_2788,N_2136,N_2167);
nand U2789 (N_2789,N_2150,N_2243);
or U2790 (N_2790,N_2279,N_2234);
nor U2791 (N_2791,N_2276,N_2083);
nor U2792 (N_2792,N_2072,N_2099);
and U2793 (N_2793,N_2392,N_2088);
xnor U2794 (N_2794,N_2045,N_2001);
and U2795 (N_2795,N_2235,N_2059);
and U2796 (N_2796,N_2357,N_2121);
and U2797 (N_2797,N_2184,N_2128);
xor U2798 (N_2798,N_2058,N_2127);
and U2799 (N_2799,N_2000,N_2294);
or U2800 (N_2800,N_2703,N_2506);
and U2801 (N_2801,N_2573,N_2538);
or U2802 (N_2802,N_2746,N_2600);
or U2803 (N_2803,N_2681,N_2599);
xnor U2804 (N_2804,N_2578,N_2477);
nand U2805 (N_2805,N_2781,N_2760);
nand U2806 (N_2806,N_2479,N_2432);
or U2807 (N_2807,N_2735,N_2523);
xnor U2808 (N_2808,N_2655,N_2639);
or U2809 (N_2809,N_2671,N_2695);
nand U2810 (N_2810,N_2789,N_2546);
nand U2811 (N_2811,N_2644,N_2463);
xor U2812 (N_2812,N_2542,N_2504);
or U2813 (N_2813,N_2541,N_2685);
nor U2814 (N_2814,N_2772,N_2441);
or U2815 (N_2815,N_2620,N_2490);
and U2816 (N_2816,N_2696,N_2783);
nand U2817 (N_2817,N_2519,N_2790);
and U2818 (N_2818,N_2420,N_2713);
xnor U2819 (N_2819,N_2635,N_2698);
nand U2820 (N_2820,N_2614,N_2739);
nand U2821 (N_2821,N_2454,N_2611);
nor U2822 (N_2822,N_2462,N_2526);
or U2823 (N_2823,N_2528,N_2427);
xor U2824 (N_2824,N_2440,N_2622);
nand U2825 (N_2825,N_2413,N_2414);
nand U2826 (N_2826,N_2785,N_2527);
nand U2827 (N_2827,N_2492,N_2687);
nand U2828 (N_2828,N_2552,N_2660);
or U2829 (N_2829,N_2792,N_2525);
and U2830 (N_2830,N_2484,N_2469);
or U2831 (N_2831,N_2710,N_2791);
nand U2832 (N_2832,N_2607,N_2457);
or U2833 (N_2833,N_2470,N_2659);
xnor U2834 (N_2834,N_2697,N_2664);
xor U2835 (N_2835,N_2627,N_2613);
nand U2836 (N_2836,N_2530,N_2582);
nor U2837 (N_2837,N_2480,N_2769);
or U2838 (N_2838,N_2483,N_2586);
nand U2839 (N_2839,N_2491,N_2505);
xor U2840 (N_2840,N_2471,N_2690);
nand U2841 (N_2841,N_2476,N_2631);
or U2842 (N_2842,N_2455,N_2422);
xnor U2843 (N_2843,N_2540,N_2517);
nand U2844 (N_2844,N_2765,N_2650);
nor U2845 (N_2845,N_2726,N_2445);
nand U2846 (N_2846,N_2515,N_2720);
xor U2847 (N_2847,N_2736,N_2674);
nor U2848 (N_2848,N_2668,N_2553);
or U2849 (N_2849,N_2705,N_2592);
nor U2850 (N_2850,N_2663,N_2562);
or U2851 (N_2851,N_2612,N_2550);
or U2852 (N_2852,N_2428,N_2782);
nand U2853 (N_2853,N_2770,N_2638);
nand U2854 (N_2854,N_2533,N_2532);
nand U2855 (N_2855,N_2495,N_2508);
or U2856 (N_2856,N_2594,N_2721);
nor U2857 (N_2857,N_2794,N_2418);
nand U2858 (N_2858,N_2590,N_2511);
xnor U2859 (N_2859,N_2482,N_2534);
xor U2860 (N_2860,N_2501,N_2725);
xnor U2861 (N_2861,N_2734,N_2684);
nor U2862 (N_2862,N_2521,N_2448);
nor U2863 (N_2863,N_2425,N_2617);
xor U2864 (N_2864,N_2507,N_2738);
nor U2865 (N_2865,N_2439,N_2412);
and U2866 (N_2866,N_2716,N_2547);
xnor U2867 (N_2867,N_2577,N_2410);
or U2868 (N_2868,N_2597,N_2580);
xor U2869 (N_2869,N_2675,N_2548);
nor U2870 (N_2870,N_2634,N_2758);
nand U2871 (N_2871,N_2679,N_2670);
xnor U2872 (N_2872,N_2767,N_2694);
nand U2873 (N_2873,N_2752,N_2688);
nand U2874 (N_2874,N_2699,N_2485);
nor U2875 (N_2875,N_2755,N_2708);
nor U2876 (N_2876,N_2610,N_2784);
nand U2877 (N_2877,N_2678,N_2615);
xnor U2878 (N_2878,N_2447,N_2754);
nor U2879 (N_2879,N_2574,N_2549);
nor U2880 (N_2880,N_2632,N_2741);
or U2881 (N_2881,N_2443,N_2561);
and U2882 (N_2882,N_2753,N_2798);
or U2883 (N_2883,N_2654,N_2619);
or U2884 (N_2884,N_2467,N_2665);
or U2885 (N_2885,N_2702,N_2570);
xor U2886 (N_2886,N_2777,N_2451);
or U2887 (N_2887,N_2700,N_2621);
or U2888 (N_2888,N_2737,N_2707);
xnor U2889 (N_2889,N_2558,N_2536);
xnor U2890 (N_2890,N_2588,N_2723);
xor U2891 (N_2891,N_2647,N_2793);
or U2892 (N_2892,N_2625,N_2453);
nor U2893 (N_2893,N_2626,N_2435);
and U2894 (N_2894,N_2421,N_2404);
or U2895 (N_2895,N_2596,N_2624);
xor U2896 (N_2896,N_2669,N_2520);
nor U2897 (N_2897,N_2569,N_2692);
nor U2898 (N_2898,N_2513,N_2572);
and U2899 (N_2899,N_2799,N_2608);
xnor U2900 (N_2900,N_2729,N_2584);
and U2901 (N_2901,N_2731,N_2740);
nor U2902 (N_2902,N_2605,N_2401);
xor U2903 (N_2903,N_2653,N_2494);
or U2904 (N_2904,N_2606,N_2510);
nand U2905 (N_2905,N_2406,N_2557);
or U2906 (N_2906,N_2604,N_2555);
or U2907 (N_2907,N_2762,N_2514);
or U2908 (N_2908,N_2633,N_2499);
and U2909 (N_2909,N_2400,N_2645);
and U2910 (N_2910,N_2556,N_2779);
nor U2911 (N_2911,N_2727,N_2748);
nor U2912 (N_2912,N_2623,N_2539);
nor U2913 (N_2913,N_2717,N_2486);
nor U2914 (N_2914,N_2518,N_2651);
nor U2915 (N_2915,N_2787,N_2661);
or U2916 (N_2916,N_2648,N_2459);
or U2917 (N_2917,N_2630,N_2641);
xor U2918 (N_2918,N_2642,N_2442);
and U2919 (N_2919,N_2656,N_2559);
or U2920 (N_2920,N_2689,N_2461);
nor U2921 (N_2921,N_2543,N_2408);
or U2922 (N_2922,N_2747,N_2643);
nor U2923 (N_2923,N_2683,N_2657);
or U2924 (N_2924,N_2693,N_2497);
nor U2925 (N_2925,N_2468,N_2718);
and U2926 (N_2926,N_2402,N_2452);
and U2927 (N_2927,N_2637,N_2728);
or U2928 (N_2928,N_2714,N_2446);
nand U2929 (N_2929,N_2733,N_2424);
xor U2930 (N_2930,N_2576,N_2593);
xnor U2931 (N_2931,N_2512,N_2436);
nor U2932 (N_2932,N_2666,N_2481);
or U2933 (N_2933,N_2750,N_2583);
or U2934 (N_2934,N_2776,N_2545);
or U2935 (N_2935,N_2475,N_2673);
nor U2936 (N_2936,N_2730,N_2431);
or U2937 (N_2937,N_2509,N_2672);
nor U2938 (N_2938,N_2773,N_2701);
and U2939 (N_2939,N_2759,N_2778);
nor U2940 (N_2940,N_2761,N_2680);
nor U2941 (N_2941,N_2745,N_2749);
xor U2942 (N_2942,N_2722,N_2568);
or U2943 (N_2943,N_2602,N_2551);
or U2944 (N_2944,N_2496,N_2591);
or U2945 (N_2945,N_2628,N_2516);
nand U2946 (N_2946,N_2662,N_2598);
and U2947 (N_2947,N_2712,N_2775);
nand U2948 (N_2948,N_2658,N_2649);
nor U2949 (N_2949,N_2601,N_2544);
xor U2950 (N_2950,N_2724,N_2488);
nor U2951 (N_2951,N_2732,N_2757);
and U2952 (N_2952,N_2751,N_2585);
nand U2953 (N_2953,N_2711,N_2438);
and U2954 (N_2954,N_2609,N_2640);
nor U2955 (N_2955,N_2756,N_2429);
xor U2956 (N_2956,N_2524,N_2560);
and U2957 (N_2957,N_2458,N_2682);
and U2958 (N_2958,N_2629,N_2780);
or U2959 (N_2959,N_2763,N_2567);
nor U2960 (N_2960,N_2786,N_2691);
and U2961 (N_2961,N_2487,N_2709);
or U2962 (N_2962,N_2575,N_2473);
or U2963 (N_2963,N_2677,N_2449);
and U2964 (N_2964,N_2407,N_2416);
or U2965 (N_2965,N_2704,N_2478);
or U2966 (N_2966,N_2405,N_2464);
nand U2967 (N_2967,N_2456,N_2566);
xor U2968 (N_2968,N_2676,N_2581);
and U2969 (N_2969,N_2686,N_2616);
nor U2970 (N_2970,N_2474,N_2502);
nor U2971 (N_2971,N_2423,N_2667);
and U2972 (N_2972,N_2433,N_2465);
and U2973 (N_2973,N_2719,N_2764);
xnor U2974 (N_2974,N_2564,N_2706);
or U2975 (N_2975,N_2409,N_2489);
and U2976 (N_2976,N_2472,N_2715);
nand U2977 (N_2977,N_2411,N_2646);
and U2978 (N_2978,N_2537,N_2795);
nor U2979 (N_2979,N_2768,N_2603);
or U2980 (N_2980,N_2535,N_2493);
xnor U2981 (N_2981,N_2563,N_2743);
and U2982 (N_2982,N_2788,N_2797);
or U2983 (N_2983,N_2652,N_2403);
nor U2984 (N_2984,N_2766,N_2571);
xor U2985 (N_2985,N_2531,N_2434);
xor U2986 (N_2986,N_2774,N_2589);
and U2987 (N_2987,N_2636,N_2450);
nor U2988 (N_2988,N_2554,N_2796);
nor U2989 (N_2989,N_2595,N_2742);
nor U2990 (N_2990,N_2444,N_2419);
nor U2991 (N_2991,N_2503,N_2771);
nand U2992 (N_2992,N_2430,N_2500);
or U2993 (N_2993,N_2460,N_2529);
nand U2994 (N_2994,N_2744,N_2417);
or U2995 (N_2995,N_2522,N_2579);
nand U2996 (N_2996,N_2415,N_2466);
nand U2997 (N_2997,N_2437,N_2498);
or U2998 (N_2998,N_2587,N_2426);
nor U2999 (N_2999,N_2565,N_2618);
nand U3000 (N_3000,N_2641,N_2665);
nand U3001 (N_3001,N_2621,N_2475);
nand U3002 (N_3002,N_2439,N_2492);
nor U3003 (N_3003,N_2704,N_2715);
xor U3004 (N_3004,N_2771,N_2623);
nand U3005 (N_3005,N_2633,N_2757);
nand U3006 (N_3006,N_2776,N_2510);
xor U3007 (N_3007,N_2613,N_2596);
or U3008 (N_3008,N_2692,N_2626);
or U3009 (N_3009,N_2517,N_2650);
nor U3010 (N_3010,N_2542,N_2688);
nor U3011 (N_3011,N_2786,N_2444);
nand U3012 (N_3012,N_2782,N_2552);
xor U3013 (N_3013,N_2532,N_2542);
nor U3014 (N_3014,N_2537,N_2568);
nor U3015 (N_3015,N_2521,N_2760);
and U3016 (N_3016,N_2609,N_2617);
nor U3017 (N_3017,N_2784,N_2492);
nand U3018 (N_3018,N_2657,N_2567);
nor U3019 (N_3019,N_2480,N_2788);
nor U3020 (N_3020,N_2659,N_2611);
or U3021 (N_3021,N_2654,N_2744);
nand U3022 (N_3022,N_2610,N_2629);
or U3023 (N_3023,N_2613,N_2785);
nand U3024 (N_3024,N_2500,N_2436);
or U3025 (N_3025,N_2648,N_2688);
or U3026 (N_3026,N_2675,N_2479);
or U3027 (N_3027,N_2462,N_2714);
and U3028 (N_3028,N_2593,N_2502);
nand U3029 (N_3029,N_2526,N_2633);
nor U3030 (N_3030,N_2552,N_2790);
nand U3031 (N_3031,N_2531,N_2572);
and U3032 (N_3032,N_2566,N_2671);
and U3033 (N_3033,N_2552,N_2450);
or U3034 (N_3034,N_2427,N_2607);
nor U3035 (N_3035,N_2430,N_2720);
and U3036 (N_3036,N_2452,N_2598);
nor U3037 (N_3037,N_2482,N_2635);
nor U3038 (N_3038,N_2427,N_2777);
and U3039 (N_3039,N_2687,N_2609);
or U3040 (N_3040,N_2446,N_2462);
or U3041 (N_3041,N_2422,N_2714);
and U3042 (N_3042,N_2726,N_2469);
xnor U3043 (N_3043,N_2646,N_2465);
or U3044 (N_3044,N_2645,N_2429);
xnor U3045 (N_3045,N_2574,N_2502);
or U3046 (N_3046,N_2427,N_2616);
nor U3047 (N_3047,N_2785,N_2620);
or U3048 (N_3048,N_2666,N_2678);
or U3049 (N_3049,N_2629,N_2754);
nand U3050 (N_3050,N_2545,N_2416);
xnor U3051 (N_3051,N_2777,N_2737);
and U3052 (N_3052,N_2598,N_2417);
or U3053 (N_3053,N_2500,N_2632);
and U3054 (N_3054,N_2446,N_2493);
nand U3055 (N_3055,N_2422,N_2586);
or U3056 (N_3056,N_2773,N_2635);
or U3057 (N_3057,N_2450,N_2726);
xnor U3058 (N_3058,N_2560,N_2718);
nor U3059 (N_3059,N_2629,N_2778);
xor U3060 (N_3060,N_2758,N_2690);
and U3061 (N_3061,N_2463,N_2704);
nand U3062 (N_3062,N_2409,N_2672);
nor U3063 (N_3063,N_2491,N_2716);
and U3064 (N_3064,N_2534,N_2738);
nor U3065 (N_3065,N_2528,N_2505);
or U3066 (N_3066,N_2515,N_2427);
or U3067 (N_3067,N_2538,N_2532);
or U3068 (N_3068,N_2747,N_2645);
or U3069 (N_3069,N_2596,N_2725);
and U3070 (N_3070,N_2773,N_2696);
xor U3071 (N_3071,N_2482,N_2745);
and U3072 (N_3072,N_2431,N_2642);
nand U3073 (N_3073,N_2573,N_2772);
nor U3074 (N_3074,N_2559,N_2561);
xnor U3075 (N_3075,N_2746,N_2647);
or U3076 (N_3076,N_2550,N_2589);
and U3077 (N_3077,N_2555,N_2764);
xnor U3078 (N_3078,N_2559,N_2604);
nor U3079 (N_3079,N_2751,N_2767);
xor U3080 (N_3080,N_2680,N_2618);
xor U3081 (N_3081,N_2670,N_2462);
xnor U3082 (N_3082,N_2714,N_2674);
nor U3083 (N_3083,N_2521,N_2626);
nor U3084 (N_3084,N_2406,N_2506);
or U3085 (N_3085,N_2430,N_2687);
or U3086 (N_3086,N_2697,N_2548);
and U3087 (N_3087,N_2718,N_2570);
and U3088 (N_3088,N_2783,N_2640);
nand U3089 (N_3089,N_2759,N_2733);
xor U3090 (N_3090,N_2601,N_2772);
xnor U3091 (N_3091,N_2473,N_2463);
nor U3092 (N_3092,N_2472,N_2751);
xnor U3093 (N_3093,N_2794,N_2699);
or U3094 (N_3094,N_2690,N_2565);
nand U3095 (N_3095,N_2774,N_2590);
xnor U3096 (N_3096,N_2494,N_2404);
xor U3097 (N_3097,N_2704,N_2454);
or U3098 (N_3098,N_2607,N_2779);
nand U3099 (N_3099,N_2791,N_2602);
xnor U3100 (N_3100,N_2692,N_2632);
or U3101 (N_3101,N_2561,N_2508);
xor U3102 (N_3102,N_2659,N_2728);
and U3103 (N_3103,N_2688,N_2428);
xnor U3104 (N_3104,N_2745,N_2590);
xor U3105 (N_3105,N_2565,N_2788);
and U3106 (N_3106,N_2409,N_2744);
or U3107 (N_3107,N_2685,N_2642);
nor U3108 (N_3108,N_2698,N_2734);
nand U3109 (N_3109,N_2581,N_2766);
nand U3110 (N_3110,N_2404,N_2679);
and U3111 (N_3111,N_2547,N_2536);
and U3112 (N_3112,N_2618,N_2536);
xor U3113 (N_3113,N_2769,N_2497);
xor U3114 (N_3114,N_2472,N_2407);
and U3115 (N_3115,N_2558,N_2765);
nand U3116 (N_3116,N_2474,N_2418);
or U3117 (N_3117,N_2652,N_2402);
nor U3118 (N_3118,N_2470,N_2518);
or U3119 (N_3119,N_2446,N_2706);
and U3120 (N_3120,N_2554,N_2502);
nand U3121 (N_3121,N_2440,N_2659);
xor U3122 (N_3122,N_2612,N_2585);
xor U3123 (N_3123,N_2768,N_2566);
or U3124 (N_3124,N_2473,N_2712);
or U3125 (N_3125,N_2470,N_2666);
or U3126 (N_3126,N_2461,N_2555);
xor U3127 (N_3127,N_2659,N_2594);
and U3128 (N_3128,N_2702,N_2532);
xor U3129 (N_3129,N_2632,N_2525);
xor U3130 (N_3130,N_2497,N_2786);
and U3131 (N_3131,N_2622,N_2443);
nor U3132 (N_3132,N_2651,N_2458);
and U3133 (N_3133,N_2569,N_2715);
or U3134 (N_3134,N_2561,N_2647);
and U3135 (N_3135,N_2694,N_2697);
and U3136 (N_3136,N_2622,N_2789);
nand U3137 (N_3137,N_2629,N_2424);
xnor U3138 (N_3138,N_2558,N_2456);
and U3139 (N_3139,N_2472,N_2508);
nor U3140 (N_3140,N_2555,N_2556);
xnor U3141 (N_3141,N_2619,N_2578);
nor U3142 (N_3142,N_2719,N_2572);
nand U3143 (N_3143,N_2516,N_2654);
or U3144 (N_3144,N_2648,N_2526);
nand U3145 (N_3145,N_2461,N_2489);
nand U3146 (N_3146,N_2755,N_2614);
nand U3147 (N_3147,N_2558,N_2464);
nand U3148 (N_3148,N_2516,N_2538);
xor U3149 (N_3149,N_2628,N_2653);
nand U3150 (N_3150,N_2510,N_2757);
nand U3151 (N_3151,N_2736,N_2416);
xnor U3152 (N_3152,N_2645,N_2761);
nor U3153 (N_3153,N_2622,N_2480);
nor U3154 (N_3154,N_2740,N_2497);
and U3155 (N_3155,N_2753,N_2730);
nor U3156 (N_3156,N_2631,N_2512);
nor U3157 (N_3157,N_2656,N_2686);
and U3158 (N_3158,N_2771,N_2500);
and U3159 (N_3159,N_2734,N_2456);
nor U3160 (N_3160,N_2473,N_2435);
xnor U3161 (N_3161,N_2584,N_2599);
nor U3162 (N_3162,N_2691,N_2417);
or U3163 (N_3163,N_2488,N_2454);
nand U3164 (N_3164,N_2467,N_2637);
and U3165 (N_3165,N_2756,N_2555);
nor U3166 (N_3166,N_2450,N_2697);
or U3167 (N_3167,N_2448,N_2597);
xnor U3168 (N_3168,N_2582,N_2503);
nand U3169 (N_3169,N_2611,N_2525);
nand U3170 (N_3170,N_2404,N_2682);
xnor U3171 (N_3171,N_2664,N_2786);
nor U3172 (N_3172,N_2472,N_2686);
xor U3173 (N_3173,N_2580,N_2663);
and U3174 (N_3174,N_2764,N_2492);
xor U3175 (N_3175,N_2772,N_2718);
nand U3176 (N_3176,N_2738,N_2779);
and U3177 (N_3177,N_2532,N_2731);
xor U3178 (N_3178,N_2577,N_2658);
nand U3179 (N_3179,N_2442,N_2650);
nor U3180 (N_3180,N_2490,N_2538);
xnor U3181 (N_3181,N_2563,N_2625);
xnor U3182 (N_3182,N_2473,N_2636);
nand U3183 (N_3183,N_2663,N_2536);
nand U3184 (N_3184,N_2784,N_2762);
or U3185 (N_3185,N_2758,N_2603);
xor U3186 (N_3186,N_2438,N_2449);
nor U3187 (N_3187,N_2716,N_2509);
and U3188 (N_3188,N_2419,N_2630);
nand U3189 (N_3189,N_2734,N_2794);
xor U3190 (N_3190,N_2614,N_2665);
or U3191 (N_3191,N_2454,N_2477);
nand U3192 (N_3192,N_2638,N_2664);
nand U3193 (N_3193,N_2761,N_2624);
nor U3194 (N_3194,N_2660,N_2753);
xor U3195 (N_3195,N_2730,N_2787);
xnor U3196 (N_3196,N_2695,N_2561);
or U3197 (N_3197,N_2525,N_2529);
nand U3198 (N_3198,N_2597,N_2434);
nor U3199 (N_3199,N_2712,N_2495);
xor U3200 (N_3200,N_3139,N_3175);
xnor U3201 (N_3201,N_3011,N_2952);
and U3202 (N_3202,N_3158,N_3198);
or U3203 (N_3203,N_2938,N_3087);
nand U3204 (N_3204,N_2898,N_3150);
or U3205 (N_3205,N_3193,N_2890);
nand U3206 (N_3206,N_3016,N_3069);
xnor U3207 (N_3207,N_3199,N_2936);
and U3208 (N_3208,N_2904,N_3141);
and U3209 (N_3209,N_3051,N_3177);
nand U3210 (N_3210,N_2980,N_2993);
nand U3211 (N_3211,N_3037,N_3106);
nor U3212 (N_3212,N_2970,N_2876);
or U3213 (N_3213,N_2974,N_2918);
or U3214 (N_3214,N_3161,N_3067);
and U3215 (N_3215,N_3008,N_3024);
nand U3216 (N_3216,N_3181,N_3187);
nor U3217 (N_3217,N_2839,N_2841);
or U3218 (N_3218,N_2831,N_3033);
or U3219 (N_3219,N_2911,N_2947);
or U3220 (N_3220,N_3032,N_3107);
nand U3221 (N_3221,N_3125,N_2910);
nor U3222 (N_3222,N_2805,N_2972);
nor U3223 (N_3223,N_2885,N_3034);
nor U3224 (N_3224,N_3006,N_2930);
and U3225 (N_3225,N_2887,N_3116);
xor U3226 (N_3226,N_2833,N_2946);
xor U3227 (N_3227,N_2867,N_3164);
nor U3228 (N_3228,N_3036,N_3010);
or U3229 (N_3229,N_2921,N_3059);
xor U3230 (N_3230,N_3159,N_3062);
nor U3231 (N_3231,N_3196,N_3121);
nor U3232 (N_3232,N_3080,N_3029);
or U3233 (N_3233,N_3140,N_2807);
nand U3234 (N_3234,N_3179,N_3003);
or U3235 (N_3235,N_2934,N_2979);
and U3236 (N_3236,N_2826,N_2956);
or U3237 (N_3237,N_3044,N_3194);
and U3238 (N_3238,N_2883,N_3054);
xor U3239 (N_3239,N_3035,N_2865);
or U3240 (N_3240,N_3174,N_3082);
xnor U3241 (N_3241,N_3073,N_3004);
or U3242 (N_3242,N_3163,N_2895);
or U3243 (N_3243,N_3137,N_2933);
xnor U3244 (N_3244,N_3064,N_3048);
nor U3245 (N_3245,N_2837,N_2940);
and U3246 (N_3246,N_2968,N_3025);
nand U3247 (N_3247,N_2822,N_2861);
and U3248 (N_3248,N_2873,N_3118);
or U3249 (N_3249,N_3105,N_2815);
nor U3250 (N_3250,N_2958,N_2897);
nand U3251 (N_3251,N_3111,N_2830);
or U3252 (N_3252,N_3104,N_2962);
nand U3253 (N_3253,N_3076,N_3056);
and U3254 (N_3254,N_2998,N_2814);
and U3255 (N_3255,N_2823,N_2996);
nor U3256 (N_3256,N_3023,N_3001);
or U3257 (N_3257,N_2960,N_2955);
nor U3258 (N_3258,N_2913,N_3017);
nand U3259 (N_3259,N_3167,N_2868);
or U3260 (N_3260,N_3108,N_2824);
and U3261 (N_3261,N_2808,N_2984);
and U3262 (N_3262,N_3109,N_3114);
and U3263 (N_3263,N_2886,N_2893);
nand U3264 (N_3264,N_2848,N_3027);
nand U3265 (N_3265,N_2928,N_2959);
nand U3266 (N_3266,N_2879,N_3086);
nor U3267 (N_3267,N_2931,N_3135);
xnor U3268 (N_3268,N_2922,N_2969);
or U3269 (N_3269,N_3160,N_3147);
and U3270 (N_3270,N_2894,N_2994);
xnor U3271 (N_3271,N_3088,N_2812);
or U3272 (N_3272,N_2948,N_3055);
and U3273 (N_3273,N_2860,N_3012);
xnor U3274 (N_3274,N_2884,N_2908);
nand U3275 (N_3275,N_2821,N_3152);
nor U3276 (N_3276,N_2896,N_3026);
nand U3277 (N_3277,N_2877,N_2991);
xor U3278 (N_3278,N_2803,N_3149);
nor U3279 (N_3279,N_3074,N_3170);
and U3280 (N_3280,N_2920,N_2945);
or U3281 (N_3281,N_2929,N_3042);
nand U3282 (N_3282,N_2827,N_2977);
or U3283 (N_3283,N_2976,N_2872);
and U3284 (N_3284,N_3022,N_3113);
nand U3285 (N_3285,N_3090,N_2975);
nor U3286 (N_3286,N_2825,N_3182);
nor U3287 (N_3287,N_3058,N_2971);
and U3288 (N_3288,N_2995,N_2853);
and U3289 (N_3289,N_3095,N_2878);
xor U3290 (N_3290,N_3045,N_2942);
and U3291 (N_3291,N_3101,N_3039);
xnor U3292 (N_3292,N_3078,N_3171);
or U3293 (N_3293,N_2819,N_2862);
nor U3294 (N_3294,N_3180,N_3097);
or U3295 (N_3295,N_2909,N_2811);
nand U3296 (N_3296,N_3041,N_3100);
and U3297 (N_3297,N_3053,N_3191);
nand U3298 (N_3298,N_3183,N_2874);
xnor U3299 (N_3299,N_3112,N_2989);
or U3300 (N_3300,N_2801,N_3178);
xor U3301 (N_3301,N_3009,N_3168);
nand U3302 (N_3302,N_2927,N_2966);
nor U3303 (N_3303,N_3084,N_3070);
xor U3304 (N_3304,N_2905,N_3122);
nand U3305 (N_3305,N_3021,N_2828);
nor U3306 (N_3306,N_3065,N_3154);
or U3307 (N_3307,N_2817,N_3052);
and U3308 (N_3308,N_3134,N_2965);
xor U3309 (N_3309,N_2949,N_2809);
nor U3310 (N_3310,N_2856,N_3098);
xnor U3311 (N_3311,N_2900,N_2882);
or U3312 (N_3312,N_2846,N_3085);
and U3313 (N_3313,N_2914,N_2838);
xnor U3314 (N_3314,N_2891,N_3057);
nand U3315 (N_3315,N_2963,N_2802);
xnor U3316 (N_3316,N_2939,N_2985);
or U3317 (N_3317,N_2906,N_3192);
nand U3318 (N_3318,N_3145,N_2943);
xnor U3319 (N_3319,N_3172,N_2888);
and U3320 (N_3320,N_3068,N_3148);
nor U3321 (N_3321,N_3132,N_2849);
and U3322 (N_3322,N_3190,N_3103);
nor U3323 (N_3323,N_3131,N_3126);
nor U3324 (N_3324,N_3144,N_2875);
and U3325 (N_3325,N_2944,N_3020);
nor U3326 (N_3326,N_2997,N_3110);
or U3327 (N_3327,N_2820,N_2932);
nand U3328 (N_3328,N_2951,N_3093);
nor U3329 (N_3329,N_2912,N_3184);
or U3330 (N_3330,N_2973,N_3066);
nand U3331 (N_3331,N_3060,N_3138);
or U3332 (N_3332,N_3173,N_2840);
and U3333 (N_3333,N_3136,N_3153);
nand U3334 (N_3334,N_2859,N_2961);
or U3335 (N_3335,N_2889,N_3197);
nand U3336 (N_3336,N_3063,N_2845);
and U3337 (N_3337,N_3165,N_2983);
nand U3338 (N_3338,N_2901,N_3043);
nand U3339 (N_3339,N_2899,N_3030);
or U3340 (N_3340,N_3157,N_3089);
nor U3341 (N_3341,N_2880,N_3099);
and U3342 (N_3342,N_3083,N_2804);
or U3343 (N_3343,N_2843,N_2916);
nand U3344 (N_3344,N_3133,N_3130);
nor U3345 (N_3345,N_2902,N_3007);
and U3346 (N_3346,N_2937,N_3015);
or U3347 (N_3347,N_2818,N_2835);
xnor U3348 (N_3348,N_2816,N_2800);
xnor U3349 (N_3349,N_3014,N_3127);
nor U3350 (N_3350,N_2847,N_2954);
and U3351 (N_3351,N_3195,N_2806);
and U3352 (N_3352,N_3072,N_2829);
and U3353 (N_3353,N_3117,N_2836);
nand U3354 (N_3354,N_3156,N_3094);
and U3355 (N_3355,N_3000,N_2850);
nor U3356 (N_3356,N_3189,N_2844);
and U3357 (N_3357,N_2881,N_3146);
and U3358 (N_3358,N_3142,N_2967);
nor U3359 (N_3359,N_3049,N_2919);
or U3360 (N_3360,N_3129,N_2981);
or U3361 (N_3361,N_3013,N_3071);
xor U3362 (N_3362,N_2957,N_2857);
nand U3363 (N_3363,N_3115,N_2869);
xor U3364 (N_3364,N_2926,N_3151);
and U3365 (N_3365,N_2982,N_3028);
xor U3366 (N_3366,N_2852,N_2903);
or U3367 (N_3367,N_3061,N_3102);
or U3368 (N_3368,N_3040,N_3077);
and U3369 (N_3369,N_3050,N_2986);
xor U3370 (N_3370,N_2923,N_2950);
or U3371 (N_3371,N_2832,N_2813);
nand U3372 (N_3372,N_3005,N_2892);
or U3373 (N_3373,N_2854,N_2858);
nor U3374 (N_3374,N_3096,N_2925);
nor U3375 (N_3375,N_2978,N_2924);
and U3376 (N_3376,N_3018,N_3162);
or U3377 (N_3377,N_2935,N_3038);
or U3378 (N_3378,N_3188,N_3124);
or U3379 (N_3379,N_3169,N_2987);
nor U3380 (N_3380,N_3019,N_3031);
xor U3381 (N_3381,N_3176,N_2917);
or U3382 (N_3382,N_3185,N_2907);
or U3383 (N_3383,N_2941,N_2863);
and U3384 (N_3384,N_3002,N_2851);
nor U3385 (N_3385,N_3128,N_3120);
or U3386 (N_3386,N_2864,N_2988);
or U3387 (N_3387,N_2855,N_2953);
nand U3388 (N_3388,N_3155,N_2810);
nor U3389 (N_3389,N_3123,N_3166);
and U3390 (N_3390,N_2871,N_2992);
or U3391 (N_3391,N_2866,N_3079);
nand U3392 (N_3392,N_2964,N_2915);
nand U3393 (N_3393,N_3186,N_3075);
xor U3394 (N_3394,N_3047,N_3143);
nor U3395 (N_3395,N_2870,N_3081);
or U3396 (N_3396,N_2990,N_3091);
or U3397 (N_3397,N_3119,N_2842);
xor U3398 (N_3398,N_3092,N_2834);
or U3399 (N_3399,N_2999,N_3046);
nand U3400 (N_3400,N_2952,N_2948);
xor U3401 (N_3401,N_2958,N_2986);
xnor U3402 (N_3402,N_3138,N_2954);
xnor U3403 (N_3403,N_3033,N_2890);
nand U3404 (N_3404,N_3039,N_3090);
or U3405 (N_3405,N_2925,N_2804);
nand U3406 (N_3406,N_2929,N_2911);
or U3407 (N_3407,N_3004,N_3152);
nand U3408 (N_3408,N_2970,N_2982);
nand U3409 (N_3409,N_3129,N_3161);
or U3410 (N_3410,N_3060,N_2954);
and U3411 (N_3411,N_3091,N_2994);
and U3412 (N_3412,N_3156,N_3185);
nor U3413 (N_3413,N_3133,N_2941);
nor U3414 (N_3414,N_3050,N_3001);
or U3415 (N_3415,N_3056,N_2898);
xor U3416 (N_3416,N_3097,N_3044);
or U3417 (N_3417,N_2897,N_3163);
or U3418 (N_3418,N_2953,N_2993);
and U3419 (N_3419,N_3167,N_3112);
and U3420 (N_3420,N_2860,N_3079);
and U3421 (N_3421,N_3079,N_2984);
or U3422 (N_3422,N_3199,N_2876);
xor U3423 (N_3423,N_2870,N_2979);
and U3424 (N_3424,N_2940,N_2960);
nand U3425 (N_3425,N_2851,N_3017);
nor U3426 (N_3426,N_3016,N_3101);
nor U3427 (N_3427,N_2945,N_3075);
nand U3428 (N_3428,N_3154,N_2974);
nand U3429 (N_3429,N_2847,N_2816);
and U3430 (N_3430,N_3117,N_3005);
nand U3431 (N_3431,N_3095,N_3000);
xor U3432 (N_3432,N_3102,N_2856);
and U3433 (N_3433,N_2998,N_2880);
xnor U3434 (N_3434,N_3005,N_2900);
nand U3435 (N_3435,N_3111,N_2982);
xor U3436 (N_3436,N_3081,N_3090);
xnor U3437 (N_3437,N_2973,N_3019);
and U3438 (N_3438,N_3033,N_2851);
xnor U3439 (N_3439,N_3197,N_3020);
xnor U3440 (N_3440,N_2939,N_3080);
nand U3441 (N_3441,N_3030,N_2999);
or U3442 (N_3442,N_3158,N_2916);
nand U3443 (N_3443,N_2934,N_2852);
nor U3444 (N_3444,N_3128,N_3039);
or U3445 (N_3445,N_2885,N_2996);
and U3446 (N_3446,N_3152,N_2935);
and U3447 (N_3447,N_2906,N_2996);
nand U3448 (N_3448,N_3092,N_3161);
or U3449 (N_3449,N_2940,N_3127);
nor U3450 (N_3450,N_2924,N_2936);
and U3451 (N_3451,N_2841,N_3151);
and U3452 (N_3452,N_2988,N_3147);
and U3453 (N_3453,N_2857,N_3044);
nand U3454 (N_3454,N_2849,N_3131);
xor U3455 (N_3455,N_2823,N_2956);
nand U3456 (N_3456,N_3149,N_3096);
and U3457 (N_3457,N_2895,N_3139);
nor U3458 (N_3458,N_2884,N_2834);
xnor U3459 (N_3459,N_2917,N_3137);
nand U3460 (N_3460,N_3140,N_3181);
and U3461 (N_3461,N_2807,N_2877);
xnor U3462 (N_3462,N_3043,N_2808);
nand U3463 (N_3463,N_2832,N_3170);
or U3464 (N_3464,N_2995,N_2971);
and U3465 (N_3465,N_3129,N_3068);
or U3466 (N_3466,N_2894,N_3053);
or U3467 (N_3467,N_3118,N_3158);
nor U3468 (N_3468,N_3152,N_3138);
and U3469 (N_3469,N_3050,N_2824);
and U3470 (N_3470,N_2892,N_2914);
nand U3471 (N_3471,N_3126,N_3162);
and U3472 (N_3472,N_2853,N_3065);
nor U3473 (N_3473,N_2953,N_2818);
nor U3474 (N_3474,N_2970,N_2905);
or U3475 (N_3475,N_2887,N_2877);
or U3476 (N_3476,N_2918,N_3020);
and U3477 (N_3477,N_2867,N_3024);
and U3478 (N_3478,N_2882,N_2892);
nand U3479 (N_3479,N_2870,N_2997);
xor U3480 (N_3480,N_2955,N_3103);
and U3481 (N_3481,N_3183,N_2891);
nor U3482 (N_3482,N_3014,N_2906);
nor U3483 (N_3483,N_3134,N_2828);
xor U3484 (N_3484,N_2815,N_2825);
or U3485 (N_3485,N_2916,N_3121);
xor U3486 (N_3486,N_2922,N_2994);
nor U3487 (N_3487,N_3011,N_2996);
xor U3488 (N_3488,N_2910,N_2825);
xnor U3489 (N_3489,N_3015,N_2824);
or U3490 (N_3490,N_3187,N_3168);
and U3491 (N_3491,N_2950,N_2927);
or U3492 (N_3492,N_3113,N_2984);
and U3493 (N_3493,N_2820,N_2804);
nor U3494 (N_3494,N_2955,N_2845);
nand U3495 (N_3495,N_3159,N_2997);
nand U3496 (N_3496,N_2898,N_2835);
nor U3497 (N_3497,N_2972,N_2942);
xnor U3498 (N_3498,N_3092,N_2824);
and U3499 (N_3499,N_3091,N_2841);
xnor U3500 (N_3500,N_2854,N_3062);
nor U3501 (N_3501,N_2827,N_3125);
nor U3502 (N_3502,N_2858,N_3177);
nand U3503 (N_3503,N_3021,N_3172);
nor U3504 (N_3504,N_3124,N_2913);
nand U3505 (N_3505,N_2941,N_2840);
nand U3506 (N_3506,N_2967,N_2902);
or U3507 (N_3507,N_2823,N_3088);
nor U3508 (N_3508,N_2933,N_3169);
nor U3509 (N_3509,N_3081,N_2965);
xnor U3510 (N_3510,N_3171,N_2876);
xor U3511 (N_3511,N_2947,N_2884);
or U3512 (N_3512,N_3031,N_2965);
or U3513 (N_3513,N_3010,N_3019);
nand U3514 (N_3514,N_2905,N_3043);
nand U3515 (N_3515,N_2876,N_3075);
nor U3516 (N_3516,N_3185,N_3173);
and U3517 (N_3517,N_2858,N_3048);
xor U3518 (N_3518,N_2926,N_2912);
nor U3519 (N_3519,N_2951,N_2846);
and U3520 (N_3520,N_3048,N_3112);
nand U3521 (N_3521,N_2917,N_2814);
nand U3522 (N_3522,N_3158,N_2864);
nand U3523 (N_3523,N_3154,N_3096);
and U3524 (N_3524,N_3084,N_2917);
and U3525 (N_3525,N_2916,N_3167);
or U3526 (N_3526,N_3122,N_2957);
xnor U3527 (N_3527,N_3139,N_2901);
nand U3528 (N_3528,N_3199,N_2939);
nor U3529 (N_3529,N_3149,N_3080);
or U3530 (N_3530,N_2992,N_3109);
or U3531 (N_3531,N_2952,N_3197);
and U3532 (N_3532,N_2862,N_2810);
and U3533 (N_3533,N_3116,N_2895);
and U3534 (N_3534,N_3194,N_2909);
and U3535 (N_3535,N_2877,N_3064);
nand U3536 (N_3536,N_3105,N_3150);
nand U3537 (N_3537,N_3197,N_3097);
and U3538 (N_3538,N_3028,N_3090);
and U3539 (N_3539,N_3048,N_2912);
or U3540 (N_3540,N_2808,N_3108);
or U3541 (N_3541,N_3167,N_3048);
xnor U3542 (N_3542,N_3147,N_2877);
and U3543 (N_3543,N_2945,N_2987);
and U3544 (N_3544,N_2969,N_2937);
and U3545 (N_3545,N_3186,N_2871);
xor U3546 (N_3546,N_3016,N_3094);
nand U3547 (N_3547,N_3074,N_2920);
and U3548 (N_3548,N_2969,N_2959);
xnor U3549 (N_3549,N_2804,N_2957);
nor U3550 (N_3550,N_3050,N_2839);
or U3551 (N_3551,N_2887,N_3176);
nand U3552 (N_3552,N_2995,N_2813);
nand U3553 (N_3553,N_3047,N_3178);
and U3554 (N_3554,N_2800,N_2860);
nand U3555 (N_3555,N_3092,N_2823);
or U3556 (N_3556,N_2802,N_3132);
nand U3557 (N_3557,N_2810,N_2819);
or U3558 (N_3558,N_3058,N_3022);
xnor U3559 (N_3559,N_3059,N_2913);
or U3560 (N_3560,N_2957,N_3004);
xor U3561 (N_3561,N_3157,N_2840);
and U3562 (N_3562,N_3128,N_2974);
and U3563 (N_3563,N_2965,N_2856);
nor U3564 (N_3564,N_2930,N_3068);
and U3565 (N_3565,N_3077,N_3099);
or U3566 (N_3566,N_3125,N_2954);
xor U3567 (N_3567,N_2917,N_2875);
xor U3568 (N_3568,N_3016,N_3079);
nand U3569 (N_3569,N_3186,N_2842);
and U3570 (N_3570,N_3021,N_2839);
xor U3571 (N_3571,N_3114,N_2861);
nor U3572 (N_3572,N_2935,N_3016);
nor U3573 (N_3573,N_2895,N_2845);
xor U3574 (N_3574,N_2938,N_2997);
or U3575 (N_3575,N_2887,N_3077);
xnor U3576 (N_3576,N_2842,N_2829);
nand U3577 (N_3577,N_2870,N_3102);
and U3578 (N_3578,N_2936,N_2903);
nand U3579 (N_3579,N_2972,N_2893);
nand U3580 (N_3580,N_2812,N_2991);
nand U3581 (N_3581,N_3192,N_2931);
nor U3582 (N_3582,N_2878,N_3142);
xor U3583 (N_3583,N_2939,N_3156);
and U3584 (N_3584,N_2832,N_2837);
and U3585 (N_3585,N_3175,N_2841);
nor U3586 (N_3586,N_3080,N_3164);
xnor U3587 (N_3587,N_2932,N_3136);
nand U3588 (N_3588,N_3186,N_3132);
xnor U3589 (N_3589,N_2998,N_2953);
nand U3590 (N_3590,N_3186,N_3135);
xnor U3591 (N_3591,N_3061,N_2830);
and U3592 (N_3592,N_3016,N_3062);
nand U3593 (N_3593,N_3181,N_3041);
or U3594 (N_3594,N_3174,N_2997);
xnor U3595 (N_3595,N_2914,N_3174);
or U3596 (N_3596,N_2941,N_2834);
xor U3597 (N_3597,N_3146,N_3170);
or U3598 (N_3598,N_2901,N_2888);
or U3599 (N_3599,N_3057,N_2941);
or U3600 (N_3600,N_3570,N_3433);
nand U3601 (N_3601,N_3521,N_3306);
nand U3602 (N_3602,N_3445,N_3204);
and U3603 (N_3603,N_3435,N_3232);
nor U3604 (N_3604,N_3289,N_3505);
nor U3605 (N_3605,N_3368,N_3497);
and U3606 (N_3606,N_3288,N_3251);
nand U3607 (N_3607,N_3346,N_3567);
or U3608 (N_3608,N_3278,N_3331);
nor U3609 (N_3609,N_3579,N_3285);
or U3610 (N_3610,N_3245,N_3396);
and U3611 (N_3611,N_3320,N_3226);
nor U3612 (N_3612,N_3248,N_3498);
and U3613 (N_3613,N_3523,N_3566);
xor U3614 (N_3614,N_3373,N_3574);
and U3615 (N_3615,N_3565,N_3587);
and U3616 (N_3616,N_3543,N_3214);
xor U3617 (N_3617,N_3514,N_3427);
nand U3618 (N_3618,N_3321,N_3267);
nand U3619 (N_3619,N_3479,N_3298);
xor U3620 (N_3620,N_3504,N_3469);
nand U3621 (N_3621,N_3531,N_3360);
or U3622 (N_3622,N_3268,N_3413);
nor U3623 (N_3623,N_3483,N_3467);
or U3624 (N_3624,N_3317,N_3557);
xnor U3625 (N_3625,N_3376,N_3481);
nand U3626 (N_3626,N_3492,N_3548);
nand U3627 (N_3627,N_3243,N_3271);
nand U3628 (N_3628,N_3502,N_3474);
or U3629 (N_3629,N_3560,N_3593);
nor U3630 (N_3630,N_3582,N_3381);
and U3631 (N_3631,N_3430,N_3541);
nor U3632 (N_3632,N_3225,N_3510);
xor U3633 (N_3633,N_3244,N_3356);
nor U3634 (N_3634,N_3301,N_3403);
and U3635 (N_3635,N_3350,N_3341);
and U3636 (N_3636,N_3366,N_3219);
nor U3637 (N_3637,N_3429,N_3363);
xnor U3638 (N_3638,N_3280,N_3416);
or U3639 (N_3639,N_3349,N_3563);
or U3640 (N_3640,N_3421,N_3372);
nor U3641 (N_3641,N_3554,N_3410);
nand U3642 (N_3642,N_3409,N_3438);
or U3643 (N_3643,N_3526,N_3583);
or U3644 (N_3644,N_3432,N_3369);
xnor U3645 (N_3645,N_3542,N_3463);
nor U3646 (N_3646,N_3466,N_3335);
nor U3647 (N_3647,N_3499,N_3462);
nor U3648 (N_3648,N_3273,N_3391);
nand U3649 (N_3649,N_3539,N_3407);
nand U3650 (N_3650,N_3338,N_3522);
and U3651 (N_3651,N_3578,N_3465);
nor U3652 (N_3652,N_3247,N_3476);
nor U3653 (N_3653,N_3549,N_3309);
nand U3654 (N_3654,N_3353,N_3382);
nor U3655 (N_3655,N_3405,N_3550);
xor U3656 (N_3656,N_3540,N_3297);
nor U3657 (N_3657,N_3461,N_3241);
or U3658 (N_3658,N_3294,N_3420);
nand U3659 (N_3659,N_3580,N_3236);
nor U3660 (N_3660,N_3229,N_3326);
or U3661 (N_3661,N_3491,N_3392);
nand U3662 (N_3662,N_3544,N_3304);
nand U3663 (N_3663,N_3450,N_3324);
or U3664 (N_3664,N_3446,N_3328);
and U3665 (N_3665,N_3584,N_3380);
xnor U3666 (N_3666,N_3203,N_3595);
and U3667 (N_3667,N_3507,N_3598);
and U3668 (N_3668,N_3210,N_3454);
and U3669 (N_3669,N_3312,N_3254);
nor U3670 (N_3670,N_3387,N_3200);
xnor U3671 (N_3671,N_3443,N_3493);
nor U3672 (N_3672,N_3555,N_3212);
xnor U3673 (N_3673,N_3528,N_3250);
or U3674 (N_3674,N_3276,N_3313);
and U3675 (N_3675,N_3252,N_3242);
xnor U3676 (N_3676,N_3322,N_3515);
xor U3677 (N_3677,N_3290,N_3553);
nand U3678 (N_3678,N_3558,N_3472);
nand U3679 (N_3679,N_3569,N_3423);
nor U3680 (N_3680,N_3546,N_3451);
and U3681 (N_3681,N_3277,N_3470);
and U3682 (N_3682,N_3456,N_3508);
nor U3683 (N_3683,N_3545,N_3484);
or U3684 (N_3684,N_3586,N_3240);
nand U3685 (N_3685,N_3293,N_3437);
or U3686 (N_3686,N_3585,N_3547);
or U3687 (N_3687,N_3354,N_3434);
xor U3688 (N_3688,N_3340,N_3314);
or U3689 (N_3689,N_3308,N_3556);
and U3690 (N_3690,N_3424,N_3258);
xnor U3691 (N_3691,N_3230,N_3577);
and U3692 (N_3692,N_3417,N_3255);
nor U3693 (N_3693,N_3562,N_3530);
nand U3694 (N_3694,N_3342,N_3249);
and U3695 (N_3695,N_3216,N_3319);
and U3696 (N_3696,N_3404,N_3329);
nor U3697 (N_3697,N_3339,N_3383);
nand U3698 (N_3698,N_3516,N_3253);
nor U3699 (N_3699,N_3362,N_3496);
nand U3700 (N_3700,N_3415,N_3302);
nand U3701 (N_3701,N_3334,N_3345);
or U3702 (N_3702,N_3374,N_3524);
nand U3703 (N_3703,N_3468,N_3535);
nand U3704 (N_3704,N_3398,N_3482);
nand U3705 (N_3705,N_3385,N_3581);
xnor U3706 (N_3706,N_3220,N_3412);
or U3707 (N_3707,N_3457,N_3389);
and U3708 (N_3708,N_3575,N_3459);
and U3709 (N_3709,N_3263,N_3519);
and U3710 (N_3710,N_3488,N_3272);
nand U3711 (N_3711,N_3453,N_3259);
and U3712 (N_3712,N_3370,N_3239);
or U3713 (N_3713,N_3561,N_3233);
nand U3714 (N_3714,N_3591,N_3213);
nand U3715 (N_3715,N_3439,N_3441);
nand U3716 (N_3716,N_3422,N_3206);
nand U3717 (N_3717,N_3495,N_3379);
and U3718 (N_3718,N_3332,N_3477);
nand U3719 (N_3719,N_3310,N_3573);
and U3720 (N_3720,N_3596,N_3390);
nand U3721 (N_3721,N_3274,N_3300);
nand U3722 (N_3722,N_3411,N_3330);
xor U3723 (N_3723,N_3358,N_3414);
nor U3724 (N_3724,N_3221,N_3533);
nor U3725 (N_3725,N_3336,N_3395);
xnor U3726 (N_3726,N_3448,N_3426);
nand U3727 (N_3727,N_3269,N_3384);
xnor U3728 (N_3728,N_3375,N_3344);
and U3729 (N_3729,N_3568,N_3460);
nand U3730 (N_3730,N_3256,N_3223);
nand U3731 (N_3731,N_3597,N_3286);
nor U3732 (N_3732,N_3217,N_3501);
nor U3733 (N_3733,N_3265,N_3590);
or U3734 (N_3734,N_3490,N_3449);
or U3735 (N_3735,N_3231,N_3386);
or U3736 (N_3736,N_3257,N_3473);
nand U3737 (N_3737,N_3589,N_3408);
or U3738 (N_3738,N_3295,N_3208);
and U3739 (N_3739,N_3337,N_3347);
nand U3740 (N_3740,N_3287,N_3215);
nor U3741 (N_3741,N_3211,N_3537);
nor U3742 (N_3742,N_3475,N_3393);
or U3743 (N_3743,N_3348,N_3209);
xnor U3744 (N_3744,N_3487,N_3471);
or U3745 (N_3745,N_3486,N_3224);
or U3746 (N_3746,N_3520,N_3343);
or U3747 (N_3747,N_3532,N_3235);
xor U3748 (N_3748,N_3291,N_3576);
nand U3749 (N_3749,N_3361,N_3536);
nand U3750 (N_3750,N_3513,N_3359);
nor U3751 (N_3751,N_3260,N_3357);
nor U3752 (N_3752,N_3455,N_3303);
and U3753 (N_3753,N_3512,N_3351);
and U3754 (N_3754,N_3237,N_3318);
nand U3755 (N_3755,N_3447,N_3572);
and U3756 (N_3756,N_3205,N_3325);
xnor U3757 (N_3757,N_3296,N_3365);
or U3758 (N_3758,N_3305,N_3246);
and U3759 (N_3759,N_3367,N_3552);
nor U3760 (N_3760,N_3400,N_3440);
nand U3761 (N_3761,N_3262,N_3559);
xor U3762 (N_3762,N_3234,N_3480);
or U3763 (N_3763,N_3264,N_3281);
xnor U3764 (N_3764,N_3238,N_3364);
nor U3765 (N_3765,N_3444,N_3517);
nand U3766 (N_3766,N_3311,N_3592);
xnor U3767 (N_3767,N_3315,N_3352);
nand U3768 (N_3768,N_3551,N_3594);
nor U3769 (N_3769,N_3222,N_3316);
nand U3770 (N_3770,N_3292,N_3511);
and U3771 (N_3771,N_3355,N_3202);
nor U3772 (N_3772,N_3323,N_3428);
xnor U3773 (N_3773,N_3494,N_3518);
xor U3774 (N_3774,N_3378,N_3458);
xnor U3775 (N_3775,N_3436,N_3500);
and U3776 (N_3776,N_3485,N_3571);
nor U3777 (N_3777,N_3266,N_3503);
nand U3778 (N_3778,N_3425,N_3442);
or U3779 (N_3779,N_3201,N_3418);
or U3780 (N_3780,N_3283,N_3394);
nand U3781 (N_3781,N_3527,N_3529);
nand U3782 (N_3782,N_3599,N_3207);
nor U3783 (N_3783,N_3402,N_3534);
xor U3784 (N_3784,N_3588,N_3401);
nand U3785 (N_3785,N_3228,N_3227);
xnor U3786 (N_3786,N_3282,N_3464);
nand U3787 (N_3787,N_3489,N_3509);
nor U3788 (N_3788,N_3388,N_3218);
nand U3789 (N_3789,N_3419,N_3564);
nor U3790 (N_3790,N_3275,N_3284);
or U3791 (N_3791,N_3399,N_3377);
nor U3792 (N_3792,N_3431,N_3506);
nand U3793 (N_3793,N_3279,N_3261);
or U3794 (N_3794,N_3406,N_3538);
nor U3795 (N_3795,N_3299,N_3525);
nand U3796 (N_3796,N_3327,N_3371);
and U3797 (N_3797,N_3452,N_3333);
xor U3798 (N_3798,N_3270,N_3307);
and U3799 (N_3799,N_3397,N_3478);
or U3800 (N_3800,N_3412,N_3265);
nand U3801 (N_3801,N_3559,N_3230);
nand U3802 (N_3802,N_3524,N_3428);
and U3803 (N_3803,N_3326,N_3494);
nand U3804 (N_3804,N_3432,N_3218);
xor U3805 (N_3805,N_3298,N_3362);
nand U3806 (N_3806,N_3501,N_3482);
xnor U3807 (N_3807,N_3432,N_3499);
nor U3808 (N_3808,N_3438,N_3260);
nand U3809 (N_3809,N_3349,N_3345);
or U3810 (N_3810,N_3570,N_3473);
and U3811 (N_3811,N_3415,N_3207);
or U3812 (N_3812,N_3562,N_3244);
nor U3813 (N_3813,N_3408,N_3416);
or U3814 (N_3814,N_3559,N_3265);
xnor U3815 (N_3815,N_3511,N_3253);
or U3816 (N_3816,N_3562,N_3524);
nor U3817 (N_3817,N_3214,N_3383);
or U3818 (N_3818,N_3499,N_3545);
nand U3819 (N_3819,N_3556,N_3453);
nand U3820 (N_3820,N_3239,N_3340);
nand U3821 (N_3821,N_3444,N_3501);
and U3822 (N_3822,N_3283,N_3292);
nor U3823 (N_3823,N_3344,N_3220);
or U3824 (N_3824,N_3202,N_3339);
xnor U3825 (N_3825,N_3520,N_3525);
nor U3826 (N_3826,N_3257,N_3374);
nor U3827 (N_3827,N_3546,N_3307);
nor U3828 (N_3828,N_3301,N_3479);
nand U3829 (N_3829,N_3279,N_3339);
nor U3830 (N_3830,N_3597,N_3574);
nand U3831 (N_3831,N_3450,N_3473);
nand U3832 (N_3832,N_3453,N_3369);
nor U3833 (N_3833,N_3423,N_3471);
and U3834 (N_3834,N_3272,N_3441);
nand U3835 (N_3835,N_3346,N_3377);
nand U3836 (N_3836,N_3399,N_3287);
xor U3837 (N_3837,N_3519,N_3318);
xnor U3838 (N_3838,N_3212,N_3324);
nand U3839 (N_3839,N_3495,N_3573);
nand U3840 (N_3840,N_3401,N_3234);
or U3841 (N_3841,N_3495,N_3420);
nor U3842 (N_3842,N_3456,N_3569);
xnor U3843 (N_3843,N_3595,N_3586);
nand U3844 (N_3844,N_3582,N_3251);
and U3845 (N_3845,N_3525,N_3426);
and U3846 (N_3846,N_3443,N_3300);
nand U3847 (N_3847,N_3533,N_3235);
nand U3848 (N_3848,N_3265,N_3304);
and U3849 (N_3849,N_3486,N_3289);
and U3850 (N_3850,N_3389,N_3286);
xnor U3851 (N_3851,N_3348,N_3471);
or U3852 (N_3852,N_3589,N_3376);
xnor U3853 (N_3853,N_3293,N_3414);
nor U3854 (N_3854,N_3334,N_3401);
nor U3855 (N_3855,N_3234,N_3231);
nor U3856 (N_3856,N_3328,N_3300);
nor U3857 (N_3857,N_3575,N_3208);
xor U3858 (N_3858,N_3369,N_3252);
xor U3859 (N_3859,N_3586,N_3474);
nand U3860 (N_3860,N_3442,N_3259);
nand U3861 (N_3861,N_3473,N_3384);
nor U3862 (N_3862,N_3437,N_3404);
or U3863 (N_3863,N_3363,N_3472);
xor U3864 (N_3864,N_3379,N_3304);
and U3865 (N_3865,N_3495,N_3305);
and U3866 (N_3866,N_3490,N_3342);
nand U3867 (N_3867,N_3529,N_3485);
and U3868 (N_3868,N_3479,N_3557);
and U3869 (N_3869,N_3551,N_3348);
or U3870 (N_3870,N_3349,N_3461);
xnor U3871 (N_3871,N_3355,N_3292);
nand U3872 (N_3872,N_3363,N_3413);
or U3873 (N_3873,N_3291,N_3574);
or U3874 (N_3874,N_3291,N_3376);
and U3875 (N_3875,N_3594,N_3422);
nand U3876 (N_3876,N_3500,N_3512);
xnor U3877 (N_3877,N_3208,N_3269);
and U3878 (N_3878,N_3477,N_3554);
nor U3879 (N_3879,N_3391,N_3551);
nand U3880 (N_3880,N_3523,N_3588);
xor U3881 (N_3881,N_3525,N_3380);
or U3882 (N_3882,N_3579,N_3560);
nor U3883 (N_3883,N_3437,N_3469);
and U3884 (N_3884,N_3318,N_3305);
or U3885 (N_3885,N_3505,N_3532);
or U3886 (N_3886,N_3268,N_3340);
nor U3887 (N_3887,N_3424,N_3457);
or U3888 (N_3888,N_3266,N_3430);
or U3889 (N_3889,N_3402,N_3274);
nor U3890 (N_3890,N_3544,N_3459);
nor U3891 (N_3891,N_3380,N_3555);
nand U3892 (N_3892,N_3291,N_3308);
or U3893 (N_3893,N_3321,N_3431);
and U3894 (N_3894,N_3368,N_3224);
or U3895 (N_3895,N_3435,N_3592);
xnor U3896 (N_3896,N_3480,N_3460);
nand U3897 (N_3897,N_3410,N_3213);
xor U3898 (N_3898,N_3443,N_3426);
or U3899 (N_3899,N_3579,N_3583);
nand U3900 (N_3900,N_3296,N_3382);
nand U3901 (N_3901,N_3417,N_3403);
and U3902 (N_3902,N_3453,N_3330);
or U3903 (N_3903,N_3506,N_3418);
or U3904 (N_3904,N_3400,N_3346);
xor U3905 (N_3905,N_3577,N_3374);
xor U3906 (N_3906,N_3481,N_3403);
nand U3907 (N_3907,N_3445,N_3597);
or U3908 (N_3908,N_3315,N_3360);
or U3909 (N_3909,N_3231,N_3503);
nor U3910 (N_3910,N_3524,N_3222);
xor U3911 (N_3911,N_3526,N_3382);
and U3912 (N_3912,N_3350,N_3311);
or U3913 (N_3913,N_3533,N_3284);
and U3914 (N_3914,N_3492,N_3568);
nand U3915 (N_3915,N_3495,N_3529);
nor U3916 (N_3916,N_3495,N_3348);
or U3917 (N_3917,N_3571,N_3378);
xnor U3918 (N_3918,N_3497,N_3344);
nor U3919 (N_3919,N_3579,N_3425);
nor U3920 (N_3920,N_3326,N_3201);
or U3921 (N_3921,N_3394,N_3440);
or U3922 (N_3922,N_3532,N_3306);
xor U3923 (N_3923,N_3314,N_3356);
xor U3924 (N_3924,N_3481,N_3423);
nand U3925 (N_3925,N_3391,N_3207);
and U3926 (N_3926,N_3229,N_3218);
and U3927 (N_3927,N_3222,N_3452);
nand U3928 (N_3928,N_3375,N_3580);
nand U3929 (N_3929,N_3333,N_3360);
and U3930 (N_3930,N_3482,N_3366);
nor U3931 (N_3931,N_3368,N_3518);
and U3932 (N_3932,N_3445,N_3574);
xnor U3933 (N_3933,N_3528,N_3251);
nor U3934 (N_3934,N_3423,N_3298);
nor U3935 (N_3935,N_3341,N_3280);
xor U3936 (N_3936,N_3299,N_3206);
nand U3937 (N_3937,N_3225,N_3485);
or U3938 (N_3938,N_3554,N_3205);
xor U3939 (N_3939,N_3565,N_3483);
and U3940 (N_3940,N_3230,N_3328);
or U3941 (N_3941,N_3506,N_3368);
or U3942 (N_3942,N_3221,N_3398);
or U3943 (N_3943,N_3223,N_3294);
nor U3944 (N_3944,N_3412,N_3598);
nor U3945 (N_3945,N_3316,N_3501);
nand U3946 (N_3946,N_3556,N_3413);
and U3947 (N_3947,N_3395,N_3509);
or U3948 (N_3948,N_3286,N_3344);
nor U3949 (N_3949,N_3371,N_3307);
nand U3950 (N_3950,N_3598,N_3433);
nor U3951 (N_3951,N_3428,N_3223);
and U3952 (N_3952,N_3368,N_3537);
and U3953 (N_3953,N_3365,N_3210);
or U3954 (N_3954,N_3429,N_3273);
and U3955 (N_3955,N_3242,N_3417);
xnor U3956 (N_3956,N_3414,N_3277);
nor U3957 (N_3957,N_3465,N_3413);
or U3958 (N_3958,N_3392,N_3234);
nand U3959 (N_3959,N_3326,N_3538);
and U3960 (N_3960,N_3544,N_3508);
nand U3961 (N_3961,N_3373,N_3369);
and U3962 (N_3962,N_3370,N_3574);
or U3963 (N_3963,N_3473,N_3530);
and U3964 (N_3964,N_3507,N_3380);
nand U3965 (N_3965,N_3338,N_3320);
or U3966 (N_3966,N_3432,N_3494);
nand U3967 (N_3967,N_3453,N_3438);
nand U3968 (N_3968,N_3459,N_3408);
or U3969 (N_3969,N_3258,N_3206);
or U3970 (N_3970,N_3414,N_3566);
and U3971 (N_3971,N_3419,N_3280);
nand U3972 (N_3972,N_3548,N_3317);
or U3973 (N_3973,N_3293,N_3230);
xnor U3974 (N_3974,N_3377,N_3395);
nand U3975 (N_3975,N_3264,N_3207);
nor U3976 (N_3976,N_3413,N_3502);
nand U3977 (N_3977,N_3360,N_3353);
and U3978 (N_3978,N_3572,N_3379);
nor U3979 (N_3979,N_3493,N_3363);
nand U3980 (N_3980,N_3242,N_3517);
xnor U3981 (N_3981,N_3456,N_3442);
nor U3982 (N_3982,N_3211,N_3290);
xnor U3983 (N_3983,N_3288,N_3257);
and U3984 (N_3984,N_3349,N_3209);
or U3985 (N_3985,N_3239,N_3420);
nor U3986 (N_3986,N_3259,N_3398);
or U3987 (N_3987,N_3464,N_3556);
and U3988 (N_3988,N_3228,N_3307);
nor U3989 (N_3989,N_3546,N_3441);
nor U3990 (N_3990,N_3338,N_3456);
xor U3991 (N_3991,N_3513,N_3595);
nand U3992 (N_3992,N_3232,N_3553);
xnor U3993 (N_3993,N_3224,N_3357);
xor U3994 (N_3994,N_3349,N_3595);
xor U3995 (N_3995,N_3448,N_3547);
and U3996 (N_3996,N_3534,N_3438);
nor U3997 (N_3997,N_3408,N_3561);
xnor U3998 (N_3998,N_3563,N_3424);
or U3999 (N_3999,N_3203,N_3366);
nand U4000 (N_4000,N_3644,N_3875);
nor U4001 (N_4001,N_3901,N_3630);
nor U4002 (N_4002,N_3740,N_3694);
xor U4003 (N_4003,N_3874,N_3671);
or U4004 (N_4004,N_3910,N_3773);
and U4005 (N_4005,N_3873,N_3878);
xnor U4006 (N_4006,N_3943,N_3746);
nand U4007 (N_4007,N_3906,N_3655);
xnor U4008 (N_4008,N_3974,N_3652);
or U4009 (N_4009,N_3650,N_3712);
xnor U4010 (N_4010,N_3839,N_3780);
xnor U4011 (N_4011,N_3790,N_3675);
xor U4012 (N_4012,N_3733,N_3997);
xor U4013 (N_4013,N_3880,N_3635);
or U4014 (N_4014,N_3982,N_3653);
xnor U4015 (N_4015,N_3944,N_3604);
xor U4016 (N_4016,N_3667,N_3926);
or U4017 (N_4017,N_3656,N_3639);
nand U4018 (N_4018,N_3781,N_3841);
or U4019 (N_4019,N_3817,N_3867);
and U4020 (N_4020,N_3939,N_3826);
xor U4021 (N_4021,N_3664,N_3627);
xnor U4022 (N_4022,N_3835,N_3614);
xnor U4023 (N_4023,N_3897,N_3849);
nand U4024 (N_4024,N_3800,N_3603);
or U4025 (N_4025,N_3732,N_3699);
nand U4026 (N_4026,N_3634,N_3757);
nand U4027 (N_4027,N_3845,N_3713);
or U4028 (N_4028,N_3886,N_3807);
and U4029 (N_4029,N_3723,N_3809);
or U4030 (N_4030,N_3979,N_3850);
nand U4031 (N_4031,N_3913,N_3775);
nor U4032 (N_4032,N_3904,N_3629);
and U4033 (N_4033,N_3605,N_3969);
nand U4034 (N_4034,N_3611,N_3861);
or U4035 (N_4035,N_3988,N_3619);
xnor U4036 (N_4036,N_3762,N_3754);
or U4037 (N_4037,N_3753,N_3922);
nor U4038 (N_4038,N_3719,N_3683);
and U4039 (N_4039,N_3882,N_3900);
and U4040 (N_4040,N_3632,N_3899);
and U4041 (N_4041,N_3661,N_3711);
nor U4042 (N_4042,N_3784,N_3721);
and U4043 (N_4043,N_3726,N_3881);
or U4044 (N_4044,N_3698,N_3638);
nand U4045 (N_4045,N_3785,N_3720);
nor U4046 (N_4046,N_3637,N_3797);
nor U4047 (N_4047,N_3854,N_3853);
xor U4048 (N_4048,N_3991,N_3973);
nand U4049 (N_4049,N_3708,N_3654);
xnor U4050 (N_4050,N_3776,N_3600);
and U4051 (N_4051,N_3987,N_3774);
and U4052 (N_4052,N_3620,N_3858);
nand U4053 (N_4053,N_3860,N_3802);
or U4054 (N_4054,N_3617,N_3765);
nand U4055 (N_4055,N_3792,N_3889);
and U4056 (N_4056,N_3616,N_3716);
nor U4057 (N_4057,N_3633,N_3872);
or U4058 (N_4058,N_3651,N_3962);
nor U4059 (N_4059,N_3706,N_3859);
nor U4060 (N_4060,N_3981,N_3879);
nand U4061 (N_4061,N_3662,N_3688);
xor U4062 (N_4062,N_3751,N_3942);
xor U4063 (N_4063,N_3812,N_3779);
xor U4064 (N_4064,N_3609,N_3682);
nand U4065 (N_4065,N_3885,N_3978);
nand U4066 (N_4066,N_3862,N_3642);
or U4067 (N_4067,N_3813,N_3610);
nand U4068 (N_4068,N_3932,N_3980);
nand U4069 (N_4069,N_3677,N_3976);
nor U4070 (N_4070,N_3837,N_3704);
xnor U4071 (N_4071,N_3782,N_3748);
nor U4072 (N_4072,N_3832,N_3766);
or U4073 (N_4073,N_3940,N_3947);
or U4074 (N_4074,N_3703,N_3709);
nand U4075 (N_4075,N_3710,N_3787);
nand U4076 (N_4076,N_3814,N_3950);
xnor U4077 (N_4077,N_3631,N_3791);
and U4078 (N_4078,N_3657,N_3865);
and U4079 (N_4079,N_3798,N_3685);
nand U4080 (N_4080,N_3663,N_3788);
nor U4081 (N_4081,N_3640,N_3915);
and U4082 (N_4082,N_3938,N_3952);
nand U4083 (N_4083,N_3917,N_3998);
or U4084 (N_4084,N_3896,N_3730);
nor U4085 (N_4085,N_3624,N_3838);
xnor U4086 (N_4086,N_3894,N_3890);
xor U4087 (N_4087,N_3935,N_3856);
or U4088 (N_4088,N_3916,N_3953);
nand U4089 (N_4089,N_3739,N_3934);
and U4090 (N_4090,N_3876,N_3747);
and U4091 (N_4091,N_3755,N_3923);
and U4092 (N_4092,N_3696,N_3804);
nand U4093 (N_4093,N_3911,N_3602);
and U4094 (N_4094,N_3819,N_3672);
nand U4095 (N_4095,N_3618,N_3705);
and U4096 (N_4096,N_3745,N_3707);
nor U4097 (N_4097,N_3613,N_3673);
or U4098 (N_4098,N_3697,N_3684);
nand U4099 (N_4099,N_3606,N_3735);
and U4100 (N_4100,N_3975,N_3990);
or U4101 (N_4101,N_3737,N_3718);
xor U4102 (N_4102,N_3866,N_3729);
and U4103 (N_4103,N_3680,N_3808);
and U4104 (N_4104,N_3985,N_3725);
xor U4105 (N_4105,N_3972,N_3636);
nand U4106 (N_4106,N_3763,N_3670);
nand U4107 (N_4107,N_3898,N_3892);
or U4108 (N_4108,N_3601,N_3722);
or U4109 (N_4109,N_3928,N_3959);
nand U4110 (N_4110,N_3815,N_3831);
or U4111 (N_4111,N_3967,N_3818);
nand U4112 (N_4112,N_3918,N_3786);
or U4113 (N_4113,N_3921,N_3877);
or U4114 (N_4114,N_3772,N_3919);
nor U4115 (N_4115,N_3768,N_3648);
or U4116 (N_4116,N_3693,N_3803);
and U4117 (N_4117,N_3778,N_3948);
or U4118 (N_4118,N_3869,N_3727);
and U4119 (N_4119,N_3659,N_3796);
nor U4120 (N_4120,N_3895,N_3686);
nor U4121 (N_4121,N_3806,N_3700);
xnor U4122 (N_4122,N_3863,N_3647);
or U4123 (N_4123,N_3843,N_3666);
and U4124 (N_4124,N_3678,N_3759);
or U4125 (N_4125,N_3717,N_3658);
nand U4126 (N_4126,N_3825,N_3771);
xnor U4127 (N_4127,N_3665,N_3783);
nand U4128 (N_4128,N_3743,N_3714);
nor U4129 (N_4129,N_3701,N_3758);
and U4130 (N_4130,N_3914,N_3994);
and U4131 (N_4131,N_3993,N_3607);
nor U4132 (N_4132,N_3954,N_3968);
and U4133 (N_4133,N_3871,N_3695);
or U4134 (N_4134,N_3820,N_3828);
or U4135 (N_4135,N_3668,N_3902);
and U4136 (N_4136,N_3852,N_3626);
xnor U4137 (N_4137,N_3830,N_3687);
xnor U4138 (N_4138,N_3794,N_3681);
nor U4139 (N_4139,N_3690,N_3805);
and U4140 (N_4140,N_3977,N_3649);
or U4141 (N_4141,N_3761,N_3833);
or U4142 (N_4142,N_3736,N_3801);
xnor U4143 (N_4143,N_3756,N_3963);
or U4144 (N_4144,N_3933,N_3937);
nand U4145 (N_4145,N_3752,N_3789);
and U4146 (N_4146,N_3621,N_3927);
nor U4147 (N_4147,N_3957,N_3941);
or U4148 (N_4148,N_3731,N_3971);
and U4149 (N_4149,N_3692,N_3907);
or U4150 (N_4150,N_3912,N_3844);
xnor U4151 (N_4151,N_3623,N_3908);
or U4152 (N_4152,N_3965,N_3888);
or U4153 (N_4153,N_3984,N_3999);
xor U4154 (N_4154,N_3827,N_3930);
and U4155 (N_4155,N_3870,N_3691);
nand U4156 (N_4156,N_3795,N_3641);
xnor U4157 (N_4157,N_3961,N_3760);
or U4158 (N_4158,N_3864,N_3992);
or U4159 (N_4159,N_3689,N_3728);
xnor U4160 (N_4160,N_3715,N_3868);
and U4161 (N_4161,N_3986,N_3669);
or U4162 (N_4162,N_3851,N_3767);
and U4163 (N_4163,N_3738,N_3946);
and U4164 (N_4164,N_3793,N_3883);
nand U4165 (N_4165,N_3777,N_3741);
nor U4166 (N_4166,N_3966,N_3924);
and U4167 (N_4167,N_3769,N_3884);
or U4168 (N_4168,N_3960,N_3811);
or U4169 (N_4169,N_3945,N_3920);
or U4170 (N_4170,N_3983,N_3964);
nand U4171 (N_4171,N_3829,N_3949);
nor U4172 (N_4172,N_3887,N_3679);
or U4173 (N_4173,N_3742,N_3958);
and U4174 (N_4174,N_3951,N_3816);
nand U4175 (N_4175,N_3836,N_3848);
xor U4176 (N_4176,N_3847,N_3608);
nand U4177 (N_4177,N_3770,N_3615);
and U4178 (N_4178,N_3643,N_3810);
or U4179 (N_4179,N_3936,N_3749);
xnor U4180 (N_4180,N_3855,N_3646);
and U4181 (N_4181,N_3744,N_3799);
and U4182 (N_4182,N_3612,N_3625);
and U4183 (N_4183,N_3903,N_3842);
nor U4184 (N_4184,N_3724,N_3764);
nor U4185 (N_4185,N_3734,N_3840);
nor U4186 (N_4186,N_3676,N_3893);
or U4187 (N_4187,N_3970,N_3645);
nand U4188 (N_4188,N_3702,N_3857);
and U4189 (N_4189,N_3834,N_3823);
xnor U4190 (N_4190,N_3750,N_3931);
nor U4191 (N_4191,N_3824,N_3996);
nand U4192 (N_4192,N_3955,N_3925);
or U4193 (N_4193,N_3628,N_3622);
nand U4194 (N_4194,N_3891,N_3929);
nand U4195 (N_4195,N_3956,N_3846);
or U4196 (N_4196,N_3660,N_3674);
nor U4197 (N_4197,N_3909,N_3905);
nor U4198 (N_4198,N_3989,N_3822);
and U4199 (N_4199,N_3995,N_3821);
or U4200 (N_4200,N_3742,N_3707);
xnor U4201 (N_4201,N_3749,N_3646);
or U4202 (N_4202,N_3981,N_3707);
nor U4203 (N_4203,N_3648,N_3601);
and U4204 (N_4204,N_3975,N_3681);
and U4205 (N_4205,N_3717,N_3842);
xnor U4206 (N_4206,N_3710,N_3910);
xnor U4207 (N_4207,N_3721,N_3947);
or U4208 (N_4208,N_3990,N_3861);
nor U4209 (N_4209,N_3783,N_3782);
nor U4210 (N_4210,N_3696,N_3602);
nand U4211 (N_4211,N_3649,N_3783);
nand U4212 (N_4212,N_3661,N_3951);
nand U4213 (N_4213,N_3976,N_3957);
nand U4214 (N_4214,N_3666,N_3810);
xnor U4215 (N_4215,N_3890,N_3991);
xnor U4216 (N_4216,N_3871,N_3718);
nor U4217 (N_4217,N_3664,N_3862);
and U4218 (N_4218,N_3630,N_3686);
xnor U4219 (N_4219,N_3601,N_3765);
nand U4220 (N_4220,N_3709,N_3762);
nand U4221 (N_4221,N_3716,N_3638);
and U4222 (N_4222,N_3808,N_3682);
and U4223 (N_4223,N_3660,N_3760);
nand U4224 (N_4224,N_3992,N_3721);
nor U4225 (N_4225,N_3970,N_3809);
nand U4226 (N_4226,N_3981,N_3724);
xor U4227 (N_4227,N_3929,N_3868);
or U4228 (N_4228,N_3626,N_3942);
or U4229 (N_4229,N_3643,N_3682);
nand U4230 (N_4230,N_3631,N_3851);
nand U4231 (N_4231,N_3965,N_3901);
and U4232 (N_4232,N_3863,N_3858);
and U4233 (N_4233,N_3813,N_3978);
nand U4234 (N_4234,N_3985,N_3722);
and U4235 (N_4235,N_3681,N_3949);
nor U4236 (N_4236,N_3857,N_3832);
or U4237 (N_4237,N_3823,N_3656);
nor U4238 (N_4238,N_3667,N_3846);
nand U4239 (N_4239,N_3915,N_3879);
or U4240 (N_4240,N_3947,N_3749);
nor U4241 (N_4241,N_3627,N_3794);
nand U4242 (N_4242,N_3631,N_3944);
nand U4243 (N_4243,N_3918,N_3846);
and U4244 (N_4244,N_3757,N_3703);
nand U4245 (N_4245,N_3788,N_3967);
nand U4246 (N_4246,N_3728,N_3818);
and U4247 (N_4247,N_3662,N_3944);
xnor U4248 (N_4248,N_3880,N_3639);
nand U4249 (N_4249,N_3658,N_3746);
xor U4250 (N_4250,N_3828,N_3646);
xor U4251 (N_4251,N_3719,N_3656);
or U4252 (N_4252,N_3694,N_3890);
nand U4253 (N_4253,N_3807,N_3721);
and U4254 (N_4254,N_3890,N_3620);
nor U4255 (N_4255,N_3921,N_3915);
xor U4256 (N_4256,N_3623,N_3976);
xor U4257 (N_4257,N_3932,N_3610);
nand U4258 (N_4258,N_3926,N_3973);
or U4259 (N_4259,N_3626,N_3932);
or U4260 (N_4260,N_3756,N_3931);
or U4261 (N_4261,N_3909,N_3831);
nand U4262 (N_4262,N_3866,N_3976);
xor U4263 (N_4263,N_3940,N_3851);
xor U4264 (N_4264,N_3622,N_3727);
and U4265 (N_4265,N_3991,N_3618);
and U4266 (N_4266,N_3673,N_3704);
or U4267 (N_4267,N_3742,N_3951);
xnor U4268 (N_4268,N_3725,N_3967);
nand U4269 (N_4269,N_3634,N_3849);
xnor U4270 (N_4270,N_3610,N_3691);
nand U4271 (N_4271,N_3920,N_3958);
and U4272 (N_4272,N_3636,N_3601);
nor U4273 (N_4273,N_3720,N_3866);
nor U4274 (N_4274,N_3859,N_3718);
nand U4275 (N_4275,N_3946,N_3804);
nand U4276 (N_4276,N_3919,N_3707);
nand U4277 (N_4277,N_3944,N_3878);
or U4278 (N_4278,N_3666,N_3693);
xnor U4279 (N_4279,N_3960,N_3732);
xor U4280 (N_4280,N_3629,N_3923);
nor U4281 (N_4281,N_3970,N_3873);
or U4282 (N_4282,N_3680,N_3728);
nor U4283 (N_4283,N_3772,N_3748);
and U4284 (N_4284,N_3769,N_3964);
or U4285 (N_4285,N_3919,N_3848);
nor U4286 (N_4286,N_3687,N_3734);
xnor U4287 (N_4287,N_3685,N_3810);
nor U4288 (N_4288,N_3981,N_3719);
nand U4289 (N_4289,N_3804,N_3644);
or U4290 (N_4290,N_3736,N_3735);
nor U4291 (N_4291,N_3703,N_3621);
xor U4292 (N_4292,N_3681,N_3900);
and U4293 (N_4293,N_3722,N_3650);
xor U4294 (N_4294,N_3733,N_3693);
xnor U4295 (N_4295,N_3848,N_3967);
and U4296 (N_4296,N_3798,N_3710);
or U4297 (N_4297,N_3854,N_3980);
and U4298 (N_4298,N_3940,N_3910);
nor U4299 (N_4299,N_3765,N_3759);
or U4300 (N_4300,N_3759,N_3619);
and U4301 (N_4301,N_3786,N_3694);
and U4302 (N_4302,N_3728,N_3885);
or U4303 (N_4303,N_3956,N_3737);
or U4304 (N_4304,N_3854,N_3779);
nand U4305 (N_4305,N_3906,N_3915);
and U4306 (N_4306,N_3670,N_3711);
nor U4307 (N_4307,N_3902,N_3891);
and U4308 (N_4308,N_3606,N_3974);
nand U4309 (N_4309,N_3871,N_3884);
and U4310 (N_4310,N_3940,N_3673);
nand U4311 (N_4311,N_3844,N_3814);
nand U4312 (N_4312,N_3845,N_3825);
nand U4313 (N_4313,N_3825,N_3624);
nor U4314 (N_4314,N_3861,N_3747);
and U4315 (N_4315,N_3925,N_3655);
or U4316 (N_4316,N_3838,N_3753);
xnor U4317 (N_4317,N_3950,N_3614);
xnor U4318 (N_4318,N_3832,N_3803);
nand U4319 (N_4319,N_3911,N_3638);
nor U4320 (N_4320,N_3748,N_3718);
nor U4321 (N_4321,N_3914,N_3877);
nor U4322 (N_4322,N_3752,N_3919);
or U4323 (N_4323,N_3737,N_3920);
or U4324 (N_4324,N_3782,N_3726);
nor U4325 (N_4325,N_3870,N_3694);
or U4326 (N_4326,N_3946,N_3608);
or U4327 (N_4327,N_3807,N_3976);
nor U4328 (N_4328,N_3613,N_3670);
xor U4329 (N_4329,N_3654,N_3782);
or U4330 (N_4330,N_3974,N_3954);
xnor U4331 (N_4331,N_3670,N_3975);
xor U4332 (N_4332,N_3796,N_3621);
xnor U4333 (N_4333,N_3721,N_3789);
xor U4334 (N_4334,N_3788,N_3680);
nor U4335 (N_4335,N_3675,N_3997);
xnor U4336 (N_4336,N_3886,N_3847);
nor U4337 (N_4337,N_3853,N_3962);
and U4338 (N_4338,N_3698,N_3684);
or U4339 (N_4339,N_3643,N_3786);
nor U4340 (N_4340,N_3912,N_3952);
nand U4341 (N_4341,N_3774,N_3824);
or U4342 (N_4342,N_3792,N_3604);
nor U4343 (N_4343,N_3625,N_3904);
and U4344 (N_4344,N_3860,N_3973);
nor U4345 (N_4345,N_3642,N_3705);
and U4346 (N_4346,N_3604,N_3657);
nor U4347 (N_4347,N_3742,N_3902);
xor U4348 (N_4348,N_3865,N_3889);
nand U4349 (N_4349,N_3642,N_3734);
nand U4350 (N_4350,N_3980,N_3961);
or U4351 (N_4351,N_3640,N_3824);
nand U4352 (N_4352,N_3813,N_3877);
nand U4353 (N_4353,N_3848,N_3761);
nand U4354 (N_4354,N_3887,N_3991);
xor U4355 (N_4355,N_3988,N_3723);
or U4356 (N_4356,N_3730,N_3732);
and U4357 (N_4357,N_3975,N_3655);
nor U4358 (N_4358,N_3729,N_3855);
nor U4359 (N_4359,N_3832,N_3631);
nand U4360 (N_4360,N_3999,N_3780);
or U4361 (N_4361,N_3897,N_3951);
nor U4362 (N_4362,N_3629,N_3935);
or U4363 (N_4363,N_3712,N_3898);
nand U4364 (N_4364,N_3905,N_3734);
nand U4365 (N_4365,N_3649,N_3727);
nor U4366 (N_4366,N_3778,N_3752);
nand U4367 (N_4367,N_3862,N_3650);
and U4368 (N_4368,N_3669,N_3974);
xnor U4369 (N_4369,N_3869,N_3725);
and U4370 (N_4370,N_3672,N_3783);
nor U4371 (N_4371,N_3700,N_3725);
xnor U4372 (N_4372,N_3884,N_3961);
nor U4373 (N_4373,N_3986,N_3845);
nand U4374 (N_4374,N_3842,N_3910);
xor U4375 (N_4375,N_3918,N_3924);
or U4376 (N_4376,N_3895,N_3771);
nand U4377 (N_4377,N_3805,N_3621);
nor U4378 (N_4378,N_3916,N_3862);
and U4379 (N_4379,N_3947,N_3981);
nor U4380 (N_4380,N_3606,N_3916);
nand U4381 (N_4381,N_3911,N_3684);
nor U4382 (N_4382,N_3720,N_3754);
and U4383 (N_4383,N_3962,N_3754);
or U4384 (N_4384,N_3971,N_3807);
and U4385 (N_4385,N_3667,N_3648);
and U4386 (N_4386,N_3755,N_3685);
nor U4387 (N_4387,N_3824,N_3709);
nor U4388 (N_4388,N_3806,N_3664);
nor U4389 (N_4389,N_3933,N_3766);
and U4390 (N_4390,N_3964,N_3934);
nor U4391 (N_4391,N_3884,N_3669);
or U4392 (N_4392,N_3932,N_3851);
xnor U4393 (N_4393,N_3973,N_3909);
or U4394 (N_4394,N_3945,N_3950);
nand U4395 (N_4395,N_3690,N_3960);
xor U4396 (N_4396,N_3827,N_3794);
nand U4397 (N_4397,N_3900,N_3828);
xnor U4398 (N_4398,N_3845,N_3835);
nor U4399 (N_4399,N_3706,N_3923);
nand U4400 (N_4400,N_4274,N_4105);
nand U4401 (N_4401,N_4334,N_4313);
xnor U4402 (N_4402,N_4170,N_4277);
and U4403 (N_4403,N_4039,N_4162);
and U4404 (N_4404,N_4373,N_4174);
and U4405 (N_4405,N_4305,N_4267);
and U4406 (N_4406,N_4380,N_4086);
and U4407 (N_4407,N_4252,N_4003);
nand U4408 (N_4408,N_4154,N_4257);
or U4409 (N_4409,N_4331,N_4110);
nand U4410 (N_4410,N_4125,N_4289);
xor U4411 (N_4411,N_4290,N_4349);
nand U4412 (N_4412,N_4200,N_4220);
or U4413 (N_4413,N_4061,N_4320);
xnor U4414 (N_4414,N_4202,N_4332);
and U4415 (N_4415,N_4369,N_4384);
or U4416 (N_4416,N_4306,N_4047);
or U4417 (N_4417,N_4326,N_4073);
nand U4418 (N_4418,N_4315,N_4312);
xor U4419 (N_4419,N_4211,N_4316);
or U4420 (N_4420,N_4241,N_4339);
xor U4421 (N_4421,N_4067,N_4228);
nand U4422 (N_4422,N_4256,N_4194);
and U4423 (N_4423,N_4197,N_4008);
nand U4424 (N_4424,N_4282,N_4040);
nor U4425 (N_4425,N_4034,N_4084);
or U4426 (N_4426,N_4358,N_4029);
nand U4427 (N_4427,N_4063,N_4167);
xor U4428 (N_4428,N_4210,N_4002);
nor U4429 (N_4429,N_4226,N_4178);
xnor U4430 (N_4430,N_4215,N_4160);
and U4431 (N_4431,N_4307,N_4318);
and U4432 (N_4432,N_4183,N_4328);
or U4433 (N_4433,N_4177,N_4381);
or U4434 (N_4434,N_4189,N_4341);
or U4435 (N_4435,N_4106,N_4046);
and U4436 (N_4436,N_4020,N_4234);
nand U4437 (N_4437,N_4078,N_4066);
or U4438 (N_4438,N_4119,N_4043);
xor U4439 (N_4439,N_4023,N_4236);
or U4440 (N_4440,N_4145,N_4379);
nor U4441 (N_4441,N_4348,N_4155);
nor U4442 (N_4442,N_4222,N_4227);
nand U4443 (N_4443,N_4111,N_4301);
and U4444 (N_4444,N_4122,N_4135);
and U4445 (N_4445,N_4322,N_4054);
and U4446 (N_4446,N_4325,N_4346);
nor U4447 (N_4447,N_4057,N_4180);
or U4448 (N_4448,N_4157,N_4244);
nand U4449 (N_4449,N_4156,N_4038);
nor U4450 (N_4450,N_4131,N_4389);
or U4451 (N_4451,N_4016,N_4191);
or U4452 (N_4452,N_4100,N_4265);
xnor U4453 (N_4453,N_4143,N_4351);
and U4454 (N_4454,N_4260,N_4338);
or U4455 (N_4455,N_4209,N_4262);
xor U4456 (N_4456,N_4233,N_4030);
or U4457 (N_4457,N_4127,N_4015);
and U4458 (N_4458,N_4288,N_4044);
or U4459 (N_4459,N_4103,N_4272);
xor U4460 (N_4460,N_4092,N_4330);
and U4461 (N_4461,N_4059,N_4198);
and U4462 (N_4462,N_4161,N_4093);
xor U4463 (N_4463,N_4268,N_4163);
nor U4464 (N_4464,N_4229,N_4079);
nor U4465 (N_4465,N_4245,N_4012);
nor U4466 (N_4466,N_4120,N_4152);
and U4467 (N_4467,N_4058,N_4035);
xor U4468 (N_4468,N_4094,N_4324);
xor U4469 (N_4469,N_4190,N_4321);
xnor U4470 (N_4470,N_4327,N_4367);
and U4471 (N_4471,N_4371,N_4006);
and U4472 (N_4472,N_4344,N_4129);
xnor U4473 (N_4473,N_4336,N_4049);
and U4474 (N_4474,N_4001,N_4254);
xnor U4475 (N_4475,N_4353,N_4337);
nor U4476 (N_4476,N_4231,N_4273);
xor U4477 (N_4477,N_4062,N_4014);
or U4478 (N_4478,N_4212,N_4025);
nand U4479 (N_4479,N_4098,N_4284);
nor U4480 (N_4480,N_4181,N_4009);
nand U4481 (N_4481,N_4335,N_4219);
nand U4482 (N_4482,N_4088,N_4102);
nor U4483 (N_4483,N_4109,N_4390);
or U4484 (N_4484,N_4304,N_4045);
or U4485 (N_4485,N_4294,N_4146);
xnor U4486 (N_4486,N_4216,N_4280);
xnor U4487 (N_4487,N_4206,N_4101);
or U4488 (N_4488,N_4107,N_4080);
nor U4489 (N_4489,N_4286,N_4218);
nand U4490 (N_4490,N_4083,N_4354);
xor U4491 (N_4491,N_4074,N_4378);
xnor U4492 (N_4492,N_4176,N_4342);
and U4493 (N_4493,N_4214,N_4310);
xor U4494 (N_4494,N_4225,N_4293);
and U4495 (N_4495,N_4037,N_4366);
nor U4496 (N_4496,N_4395,N_4077);
nand U4497 (N_4497,N_4147,N_4171);
xor U4498 (N_4498,N_4150,N_4018);
nand U4499 (N_4499,N_4221,N_4287);
xor U4500 (N_4500,N_4246,N_4345);
nand U4501 (N_4501,N_4165,N_4064);
and U4502 (N_4502,N_4028,N_4271);
xnor U4503 (N_4503,N_4269,N_4114);
nor U4504 (N_4504,N_4208,N_4375);
or U4505 (N_4505,N_4255,N_4082);
or U4506 (N_4506,N_4319,N_4340);
nand U4507 (N_4507,N_4087,N_4270);
and U4508 (N_4508,N_4394,N_4139);
nand U4509 (N_4509,N_4377,N_4142);
nand U4510 (N_4510,N_4179,N_4075);
nor U4511 (N_4511,N_4311,N_4302);
nor U4512 (N_4512,N_4253,N_4050);
and U4513 (N_4513,N_4153,N_4070);
nand U4514 (N_4514,N_4130,N_4048);
xor U4515 (N_4515,N_4223,N_4115);
xnor U4516 (N_4516,N_4372,N_4007);
or U4517 (N_4517,N_4350,N_4362);
nor U4518 (N_4518,N_4356,N_4343);
nand U4519 (N_4519,N_4232,N_4297);
and U4520 (N_4520,N_4298,N_4141);
nand U4521 (N_4521,N_4385,N_4213);
nor U4522 (N_4522,N_4091,N_4169);
or U4523 (N_4523,N_4149,N_4329);
nor U4524 (N_4524,N_4053,N_4359);
or U4525 (N_4525,N_4242,N_4089);
or U4526 (N_4526,N_4168,N_4113);
xnor U4527 (N_4527,N_4132,N_4323);
nand U4528 (N_4528,N_4076,N_4185);
xnor U4529 (N_4529,N_4238,N_4134);
xor U4530 (N_4530,N_4317,N_4081);
xor U4531 (N_4531,N_4388,N_4104);
and U4532 (N_4532,N_4291,N_4108);
and U4533 (N_4533,N_4387,N_4022);
nand U4534 (N_4534,N_4243,N_4224);
nand U4535 (N_4535,N_4071,N_4032);
nor U4536 (N_4536,N_4195,N_4249);
nor U4537 (N_4537,N_4261,N_4173);
and U4538 (N_4538,N_4397,N_4042);
and U4539 (N_4539,N_4391,N_4392);
or U4540 (N_4540,N_4138,N_4186);
or U4541 (N_4541,N_4137,N_4203);
or U4542 (N_4542,N_4121,N_4056);
or U4543 (N_4543,N_4357,N_4279);
nand U4544 (N_4544,N_4248,N_4123);
nor U4545 (N_4545,N_4013,N_4347);
nand U4546 (N_4546,N_4299,N_4296);
and U4547 (N_4547,N_4205,N_4193);
nor U4548 (N_4548,N_4097,N_4027);
nand U4549 (N_4549,N_4264,N_4295);
or U4550 (N_4550,N_4052,N_4148);
nor U4551 (N_4551,N_4386,N_4383);
nand U4552 (N_4552,N_4204,N_4360);
or U4553 (N_4553,N_4182,N_4060);
nor U4554 (N_4554,N_4376,N_4128);
nor U4555 (N_4555,N_4283,N_4116);
or U4556 (N_4556,N_4368,N_4026);
nor U4557 (N_4557,N_4396,N_4237);
or U4558 (N_4558,N_4158,N_4352);
nor U4559 (N_4559,N_4207,N_4399);
or U4560 (N_4560,N_4055,N_4051);
nand U4561 (N_4561,N_4364,N_4144);
and U4562 (N_4562,N_4258,N_4068);
xnor U4563 (N_4563,N_4187,N_4024);
nand U4564 (N_4564,N_4117,N_4247);
nand U4565 (N_4565,N_4361,N_4309);
nand U4566 (N_4566,N_4393,N_4276);
and U4567 (N_4567,N_4259,N_4124);
or U4568 (N_4568,N_4314,N_4292);
nand U4569 (N_4569,N_4275,N_4230);
xor U4570 (N_4570,N_4065,N_4151);
xnor U4571 (N_4571,N_4099,N_4184);
nand U4572 (N_4572,N_4365,N_4370);
xnor U4573 (N_4573,N_4041,N_4036);
or U4574 (N_4574,N_4019,N_4235);
nand U4575 (N_4575,N_4239,N_4159);
nor U4576 (N_4576,N_4251,N_4300);
and U4577 (N_4577,N_4363,N_4175);
xor U4578 (N_4578,N_4201,N_4382);
nand U4579 (N_4579,N_4118,N_4285);
xor U4580 (N_4580,N_4266,N_4021);
nand U4581 (N_4581,N_4011,N_4398);
and U4582 (N_4582,N_4281,N_4090);
and U4583 (N_4583,N_4000,N_4196);
nor U4584 (N_4584,N_4126,N_4005);
nand U4585 (N_4585,N_4303,N_4263);
and U4586 (N_4586,N_4031,N_4192);
nand U4587 (N_4587,N_4240,N_4199);
nor U4588 (N_4588,N_4188,N_4095);
nor U4589 (N_4589,N_4033,N_4355);
nor U4590 (N_4590,N_4112,N_4374);
or U4591 (N_4591,N_4166,N_4172);
xnor U4592 (N_4592,N_4250,N_4140);
nor U4593 (N_4593,N_4333,N_4096);
and U4594 (N_4594,N_4164,N_4017);
and U4595 (N_4595,N_4278,N_4010);
nor U4596 (N_4596,N_4004,N_4217);
nor U4597 (N_4597,N_4085,N_4136);
or U4598 (N_4598,N_4072,N_4069);
nand U4599 (N_4599,N_4133,N_4308);
xnor U4600 (N_4600,N_4175,N_4127);
xnor U4601 (N_4601,N_4069,N_4336);
or U4602 (N_4602,N_4084,N_4087);
nand U4603 (N_4603,N_4141,N_4070);
nor U4604 (N_4604,N_4091,N_4307);
and U4605 (N_4605,N_4118,N_4135);
nand U4606 (N_4606,N_4094,N_4089);
and U4607 (N_4607,N_4046,N_4386);
nand U4608 (N_4608,N_4280,N_4188);
nand U4609 (N_4609,N_4077,N_4037);
nand U4610 (N_4610,N_4173,N_4319);
nor U4611 (N_4611,N_4394,N_4090);
and U4612 (N_4612,N_4051,N_4247);
nand U4613 (N_4613,N_4128,N_4285);
xnor U4614 (N_4614,N_4010,N_4059);
xor U4615 (N_4615,N_4159,N_4035);
nand U4616 (N_4616,N_4189,N_4052);
nand U4617 (N_4617,N_4118,N_4105);
xnor U4618 (N_4618,N_4166,N_4140);
or U4619 (N_4619,N_4059,N_4037);
nor U4620 (N_4620,N_4147,N_4060);
and U4621 (N_4621,N_4047,N_4387);
and U4622 (N_4622,N_4000,N_4089);
or U4623 (N_4623,N_4393,N_4399);
or U4624 (N_4624,N_4143,N_4121);
xnor U4625 (N_4625,N_4002,N_4246);
xnor U4626 (N_4626,N_4104,N_4250);
nand U4627 (N_4627,N_4024,N_4020);
or U4628 (N_4628,N_4292,N_4324);
or U4629 (N_4629,N_4017,N_4156);
nor U4630 (N_4630,N_4086,N_4324);
nand U4631 (N_4631,N_4323,N_4160);
nand U4632 (N_4632,N_4102,N_4398);
or U4633 (N_4633,N_4162,N_4008);
nor U4634 (N_4634,N_4288,N_4014);
and U4635 (N_4635,N_4149,N_4167);
or U4636 (N_4636,N_4236,N_4130);
or U4637 (N_4637,N_4321,N_4229);
nor U4638 (N_4638,N_4210,N_4252);
nand U4639 (N_4639,N_4194,N_4276);
and U4640 (N_4640,N_4008,N_4226);
and U4641 (N_4641,N_4319,N_4043);
xor U4642 (N_4642,N_4153,N_4108);
nor U4643 (N_4643,N_4374,N_4020);
xnor U4644 (N_4644,N_4054,N_4159);
or U4645 (N_4645,N_4214,N_4128);
nand U4646 (N_4646,N_4215,N_4034);
and U4647 (N_4647,N_4330,N_4015);
nand U4648 (N_4648,N_4330,N_4162);
or U4649 (N_4649,N_4084,N_4092);
xnor U4650 (N_4650,N_4274,N_4305);
nor U4651 (N_4651,N_4032,N_4382);
xnor U4652 (N_4652,N_4331,N_4239);
nor U4653 (N_4653,N_4335,N_4220);
or U4654 (N_4654,N_4324,N_4305);
xnor U4655 (N_4655,N_4393,N_4342);
xor U4656 (N_4656,N_4194,N_4254);
xnor U4657 (N_4657,N_4002,N_4056);
or U4658 (N_4658,N_4313,N_4018);
xnor U4659 (N_4659,N_4351,N_4365);
nand U4660 (N_4660,N_4027,N_4077);
or U4661 (N_4661,N_4238,N_4053);
and U4662 (N_4662,N_4005,N_4110);
nor U4663 (N_4663,N_4119,N_4013);
and U4664 (N_4664,N_4078,N_4316);
nand U4665 (N_4665,N_4230,N_4148);
and U4666 (N_4666,N_4395,N_4267);
xor U4667 (N_4667,N_4354,N_4190);
or U4668 (N_4668,N_4255,N_4044);
and U4669 (N_4669,N_4337,N_4066);
and U4670 (N_4670,N_4232,N_4333);
xor U4671 (N_4671,N_4292,N_4193);
xnor U4672 (N_4672,N_4028,N_4202);
or U4673 (N_4673,N_4334,N_4051);
nor U4674 (N_4674,N_4287,N_4258);
nand U4675 (N_4675,N_4232,N_4236);
nand U4676 (N_4676,N_4190,N_4377);
and U4677 (N_4677,N_4215,N_4135);
nor U4678 (N_4678,N_4034,N_4047);
nor U4679 (N_4679,N_4302,N_4368);
nand U4680 (N_4680,N_4062,N_4361);
xnor U4681 (N_4681,N_4219,N_4088);
nor U4682 (N_4682,N_4277,N_4392);
xor U4683 (N_4683,N_4384,N_4078);
nor U4684 (N_4684,N_4204,N_4119);
xor U4685 (N_4685,N_4034,N_4061);
or U4686 (N_4686,N_4109,N_4270);
nor U4687 (N_4687,N_4393,N_4206);
and U4688 (N_4688,N_4204,N_4379);
nor U4689 (N_4689,N_4297,N_4264);
xor U4690 (N_4690,N_4353,N_4071);
nor U4691 (N_4691,N_4053,N_4324);
and U4692 (N_4692,N_4276,N_4362);
nor U4693 (N_4693,N_4361,N_4038);
nand U4694 (N_4694,N_4010,N_4161);
nor U4695 (N_4695,N_4211,N_4146);
xnor U4696 (N_4696,N_4397,N_4083);
and U4697 (N_4697,N_4321,N_4137);
xor U4698 (N_4698,N_4136,N_4108);
nor U4699 (N_4699,N_4186,N_4335);
nand U4700 (N_4700,N_4322,N_4038);
and U4701 (N_4701,N_4154,N_4077);
or U4702 (N_4702,N_4388,N_4320);
xor U4703 (N_4703,N_4005,N_4382);
xor U4704 (N_4704,N_4143,N_4372);
and U4705 (N_4705,N_4008,N_4384);
nand U4706 (N_4706,N_4308,N_4033);
nand U4707 (N_4707,N_4000,N_4091);
and U4708 (N_4708,N_4014,N_4363);
and U4709 (N_4709,N_4168,N_4007);
nor U4710 (N_4710,N_4111,N_4085);
nor U4711 (N_4711,N_4279,N_4391);
xnor U4712 (N_4712,N_4314,N_4029);
nor U4713 (N_4713,N_4287,N_4139);
xor U4714 (N_4714,N_4052,N_4085);
nor U4715 (N_4715,N_4088,N_4071);
or U4716 (N_4716,N_4372,N_4171);
nor U4717 (N_4717,N_4038,N_4386);
nor U4718 (N_4718,N_4192,N_4220);
xor U4719 (N_4719,N_4111,N_4011);
or U4720 (N_4720,N_4094,N_4354);
nand U4721 (N_4721,N_4120,N_4250);
and U4722 (N_4722,N_4390,N_4025);
and U4723 (N_4723,N_4362,N_4139);
nor U4724 (N_4724,N_4327,N_4267);
or U4725 (N_4725,N_4072,N_4192);
and U4726 (N_4726,N_4363,N_4151);
nor U4727 (N_4727,N_4183,N_4107);
xor U4728 (N_4728,N_4202,N_4090);
nand U4729 (N_4729,N_4222,N_4095);
or U4730 (N_4730,N_4125,N_4334);
and U4731 (N_4731,N_4010,N_4123);
nand U4732 (N_4732,N_4302,N_4087);
and U4733 (N_4733,N_4304,N_4384);
xor U4734 (N_4734,N_4358,N_4185);
nor U4735 (N_4735,N_4148,N_4006);
or U4736 (N_4736,N_4276,N_4033);
nor U4737 (N_4737,N_4122,N_4316);
and U4738 (N_4738,N_4103,N_4006);
xor U4739 (N_4739,N_4315,N_4260);
and U4740 (N_4740,N_4007,N_4304);
nor U4741 (N_4741,N_4139,N_4036);
and U4742 (N_4742,N_4357,N_4330);
nor U4743 (N_4743,N_4202,N_4064);
and U4744 (N_4744,N_4364,N_4216);
xor U4745 (N_4745,N_4392,N_4299);
nand U4746 (N_4746,N_4152,N_4142);
nand U4747 (N_4747,N_4384,N_4070);
nand U4748 (N_4748,N_4273,N_4279);
or U4749 (N_4749,N_4045,N_4142);
and U4750 (N_4750,N_4178,N_4218);
xor U4751 (N_4751,N_4177,N_4232);
and U4752 (N_4752,N_4350,N_4213);
nor U4753 (N_4753,N_4133,N_4271);
xor U4754 (N_4754,N_4360,N_4093);
or U4755 (N_4755,N_4135,N_4076);
or U4756 (N_4756,N_4225,N_4193);
and U4757 (N_4757,N_4360,N_4172);
nor U4758 (N_4758,N_4255,N_4025);
xnor U4759 (N_4759,N_4064,N_4139);
or U4760 (N_4760,N_4257,N_4080);
nor U4761 (N_4761,N_4209,N_4367);
and U4762 (N_4762,N_4388,N_4015);
and U4763 (N_4763,N_4167,N_4211);
nand U4764 (N_4764,N_4377,N_4386);
and U4765 (N_4765,N_4267,N_4175);
xor U4766 (N_4766,N_4065,N_4093);
nor U4767 (N_4767,N_4172,N_4136);
and U4768 (N_4768,N_4017,N_4391);
xnor U4769 (N_4769,N_4117,N_4150);
nand U4770 (N_4770,N_4374,N_4008);
and U4771 (N_4771,N_4159,N_4399);
or U4772 (N_4772,N_4180,N_4117);
nor U4773 (N_4773,N_4357,N_4022);
nand U4774 (N_4774,N_4208,N_4089);
nor U4775 (N_4775,N_4268,N_4190);
nor U4776 (N_4776,N_4069,N_4068);
nand U4777 (N_4777,N_4311,N_4291);
xor U4778 (N_4778,N_4291,N_4191);
or U4779 (N_4779,N_4125,N_4244);
nand U4780 (N_4780,N_4134,N_4219);
and U4781 (N_4781,N_4380,N_4227);
xnor U4782 (N_4782,N_4147,N_4221);
xnor U4783 (N_4783,N_4159,N_4095);
or U4784 (N_4784,N_4053,N_4132);
or U4785 (N_4785,N_4117,N_4258);
and U4786 (N_4786,N_4087,N_4043);
nor U4787 (N_4787,N_4120,N_4067);
and U4788 (N_4788,N_4171,N_4140);
nor U4789 (N_4789,N_4339,N_4076);
nand U4790 (N_4790,N_4141,N_4394);
nand U4791 (N_4791,N_4204,N_4395);
or U4792 (N_4792,N_4328,N_4387);
nand U4793 (N_4793,N_4346,N_4097);
or U4794 (N_4794,N_4137,N_4196);
xor U4795 (N_4795,N_4391,N_4289);
and U4796 (N_4796,N_4024,N_4132);
or U4797 (N_4797,N_4078,N_4349);
and U4798 (N_4798,N_4290,N_4110);
or U4799 (N_4799,N_4348,N_4133);
nand U4800 (N_4800,N_4721,N_4714);
nor U4801 (N_4801,N_4660,N_4519);
and U4802 (N_4802,N_4743,N_4467);
nor U4803 (N_4803,N_4567,N_4754);
and U4804 (N_4804,N_4546,N_4544);
or U4805 (N_4805,N_4736,N_4453);
nand U4806 (N_4806,N_4563,N_4663);
and U4807 (N_4807,N_4592,N_4430);
or U4808 (N_4808,N_4596,N_4445);
xnor U4809 (N_4809,N_4530,N_4724);
nand U4810 (N_4810,N_4580,N_4585);
xor U4811 (N_4811,N_4441,N_4521);
xor U4812 (N_4812,N_4422,N_4507);
nand U4813 (N_4813,N_4644,N_4656);
nand U4814 (N_4814,N_4685,N_4751);
nor U4815 (N_4815,N_4602,N_4409);
and U4816 (N_4816,N_4742,N_4509);
or U4817 (N_4817,N_4790,N_4650);
nand U4818 (N_4818,N_4505,N_4462);
or U4819 (N_4819,N_4691,N_4683);
nand U4820 (N_4820,N_4799,N_4680);
nor U4821 (N_4821,N_4485,N_4463);
xnor U4822 (N_4822,N_4594,N_4610);
nand U4823 (N_4823,N_4551,N_4667);
and U4824 (N_4824,N_4541,N_4454);
nand U4825 (N_4825,N_4762,N_4728);
xor U4826 (N_4826,N_4695,N_4746);
nor U4827 (N_4827,N_4568,N_4452);
xor U4828 (N_4828,N_4711,N_4489);
or U4829 (N_4829,N_4536,N_4664);
xor U4830 (N_4830,N_4496,N_4626);
xnor U4831 (N_4831,N_4523,N_4584);
and U4832 (N_4832,N_4778,N_4690);
nor U4833 (N_4833,N_4624,N_4710);
or U4834 (N_4834,N_4630,N_4620);
and U4835 (N_4835,N_4439,N_4446);
nand U4836 (N_4836,N_4456,N_4730);
xnor U4837 (N_4837,N_4529,N_4460);
nand U4838 (N_4838,N_4646,N_4435);
nand U4839 (N_4839,N_4517,N_4566);
or U4840 (N_4840,N_4688,N_4639);
nand U4841 (N_4841,N_4766,N_4535);
nor U4842 (N_4842,N_4699,N_4632);
xnor U4843 (N_4843,N_4769,N_4410);
and U4844 (N_4844,N_4773,N_4638);
and U4845 (N_4845,N_4574,N_4586);
xor U4846 (N_4846,N_4666,N_4765);
and U4847 (N_4847,N_4513,N_4692);
nand U4848 (N_4848,N_4673,N_4403);
nand U4849 (N_4849,N_4508,N_4733);
xnor U4850 (N_4850,N_4616,N_4590);
or U4851 (N_4851,N_4474,N_4674);
and U4852 (N_4852,N_4793,N_4504);
nor U4853 (N_4853,N_4725,N_4526);
xor U4854 (N_4854,N_4515,N_4412);
nand U4855 (N_4855,N_4708,N_4687);
nand U4856 (N_4856,N_4482,N_4494);
or U4857 (N_4857,N_4752,N_4545);
xnor U4858 (N_4858,N_4654,N_4423);
nor U4859 (N_4859,N_4770,N_4682);
nand U4860 (N_4860,N_4753,N_4424);
or U4861 (N_4861,N_4481,N_4684);
and U4862 (N_4862,N_4777,N_4548);
nor U4863 (N_4863,N_4605,N_4514);
xnor U4864 (N_4864,N_4491,N_4716);
or U4865 (N_4865,N_4500,N_4552);
or U4866 (N_4866,N_4537,N_4681);
nand U4867 (N_4867,N_4693,N_4791);
xnor U4868 (N_4868,N_4720,N_4479);
nand U4869 (N_4869,N_4755,N_4533);
nand U4870 (N_4870,N_4640,N_4631);
or U4871 (N_4871,N_4641,N_4623);
or U4872 (N_4872,N_4516,N_4476);
nor U4873 (N_4873,N_4732,N_4598);
and U4874 (N_4874,N_4562,N_4670);
xor U4875 (N_4875,N_4502,N_4749);
and U4876 (N_4876,N_4741,N_4712);
and U4877 (N_4877,N_4459,N_4643);
nor U4878 (N_4878,N_4417,N_4540);
and U4879 (N_4879,N_4577,N_4557);
xor U4880 (N_4880,N_4661,N_4745);
xnor U4881 (N_4881,N_4652,N_4442);
or U4882 (N_4882,N_4414,N_4560);
nor U4883 (N_4883,N_4676,N_4490);
nand U4884 (N_4884,N_4703,N_4492);
nor U4885 (N_4885,N_4635,N_4555);
nand U4886 (N_4886,N_4748,N_4582);
or U4887 (N_4887,N_4416,N_4431);
xor U4888 (N_4888,N_4539,N_4653);
nand U4889 (N_4889,N_4677,N_4478);
xor U4890 (N_4890,N_4468,N_4565);
and U4891 (N_4891,N_4591,N_4633);
or U4892 (N_4892,N_4727,N_4651);
and U4893 (N_4893,N_4600,N_4700);
nand U4894 (N_4894,N_4455,N_4538);
and U4895 (N_4895,N_4593,N_4675);
and U4896 (N_4896,N_4495,N_4512);
xor U4897 (N_4897,N_4419,N_4451);
and U4898 (N_4898,N_4744,N_4718);
nand U4899 (N_4899,N_4776,N_4606);
or U4900 (N_4900,N_4797,N_4415);
and U4901 (N_4901,N_4556,N_4464);
nand U4902 (N_4902,N_4614,N_4740);
nor U4903 (N_4903,N_4411,N_4449);
nor U4904 (N_4904,N_4406,N_4483);
xor U4905 (N_4905,N_4796,N_4480);
xor U4906 (N_4906,N_4629,N_4707);
and U4907 (N_4907,N_4785,N_4611);
nor U4908 (N_4908,N_4501,N_4433);
nor U4909 (N_4909,N_4665,N_4561);
nand U4910 (N_4910,N_4783,N_4534);
nand U4911 (N_4911,N_4472,N_4617);
and U4912 (N_4912,N_4434,N_4771);
and U4913 (N_4913,N_4671,N_4607);
nand U4914 (N_4914,N_4627,N_4625);
xnor U4915 (N_4915,N_4789,N_4447);
or U4916 (N_4916,N_4589,N_4443);
nor U4917 (N_4917,N_4525,N_4679);
nand U4918 (N_4918,N_4713,N_4759);
nor U4919 (N_4919,N_4575,N_4609);
nor U4920 (N_4920,N_4738,N_4405);
xor U4921 (N_4921,N_4510,N_4780);
nand U4922 (N_4922,N_4787,N_4628);
and U4923 (N_4923,N_4484,N_4599);
xor U4924 (N_4924,N_4798,N_4524);
nor U4925 (N_4925,N_4788,N_4794);
nor U4926 (N_4926,N_4466,N_4553);
xor U4927 (N_4927,N_4702,N_4781);
xnor U4928 (N_4928,N_4709,N_4698);
and U4929 (N_4929,N_4413,N_4706);
nor U4930 (N_4930,N_4701,N_4764);
nor U4931 (N_4931,N_4572,N_4795);
xor U4932 (N_4932,N_4694,N_4475);
or U4933 (N_4933,N_4717,N_4613);
and U4934 (N_4934,N_4722,N_4618);
nand U4935 (N_4935,N_4457,N_4658);
xnor U4936 (N_4936,N_4772,N_4668);
nor U4937 (N_4937,N_4404,N_4615);
and U4938 (N_4938,N_4437,N_4686);
and U4939 (N_4939,N_4608,N_4470);
or U4940 (N_4940,N_4657,N_4655);
nand U4941 (N_4941,N_4554,N_4418);
and U4942 (N_4942,N_4786,N_4486);
or U4943 (N_4943,N_4542,N_4550);
and U4944 (N_4944,N_4723,N_4767);
and U4945 (N_4945,N_4579,N_4719);
xnor U4946 (N_4946,N_4637,N_4757);
and U4947 (N_4947,N_4648,N_4581);
nor U4948 (N_4948,N_4473,N_4729);
or U4949 (N_4949,N_4761,N_4436);
nand U4950 (N_4950,N_4522,N_4649);
nand U4951 (N_4951,N_4559,N_4739);
nor U4952 (N_4952,N_4527,N_4726);
and U4953 (N_4953,N_4571,N_4493);
and U4954 (N_4954,N_4401,N_4428);
nor U4955 (N_4955,N_4715,N_4775);
xor U4956 (N_4956,N_4488,N_4779);
and U4957 (N_4957,N_4645,N_4774);
nand U4958 (N_4958,N_4603,N_4497);
nor U4959 (N_4959,N_4543,N_4531);
xor U4960 (N_4960,N_4421,N_4426);
xnor U4961 (N_4961,N_4465,N_4407);
nor U4962 (N_4962,N_4578,N_4420);
nand U4963 (N_4963,N_4469,N_4621);
nor U4964 (N_4964,N_4471,N_4458);
xor U4965 (N_4965,N_4400,N_4642);
or U4966 (N_4966,N_4601,N_4438);
nor U4967 (N_4967,N_4669,N_4763);
nor U4968 (N_4968,N_4503,N_4532);
nand U4969 (N_4969,N_4784,N_4782);
nand U4970 (N_4970,N_4672,N_4734);
nand U4971 (N_4971,N_4558,N_4549);
or U4972 (N_4972,N_4768,N_4612);
nor U4973 (N_4973,N_4570,N_4518);
and U4974 (N_4974,N_4737,N_4689);
nand U4975 (N_4975,N_4520,N_4750);
and U4976 (N_4976,N_4647,N_4432);
or U4977 (N_4977,N_4498,N_4588);
nor U4978 (N_4978,N_4487,N_4634);
nor U4979 (N_4979,N_4747,N_4547);
nor U4980 (N_4980,N_4696,N_4659);
xnor U4981 (N_4981,N_4569,N_4705);
xor U4982 (N_4982,N_4499,N_4528);
nand U4983 (N_4983,N_4444,N_4704);
xnor U4984 (N_4984,N_4576,N_4619);
nor U4985 (N_4985,N_4573,N_4511);
nor U4986 (N_4986,N_4429,N_4450);
nand U4987 (N_4987,N_4402,N_4583);
nor U4988 (N_4988,N_4408,N_4756);
xor U4989 (N_4989,N_4440,N_4595);
nand U4990 (N_4990,N_4731,N_4760);
nor U4991 (N_4991,N_4597,N_4425);
xnor U4992 (N_4992,N_4636,N_4678);
xnor U4993 (N_4993,N_4792,N_4662);
nor U4994 (N_4994,N_4427,N_4448);
nor U4995 (N_4995,N_4587,N_4564);
or U4996 (N_4996,N_4477,N_4622);
nor U4997 (N_4997,N_4697,N_4604);
or U4998 (N_4998,N_4735,N_4506);
xor U4999 (N_4999,N_4461,N_4758);
xor U5000 (N_5000,N_4706,N_4567);
or U5001 (N_5001,N_4797,N_4643);
nor U5002 (N_5002,N_4496,N_4468);
and U5003 (N_5003,N_4655,N_4590);
nand U5004 (N_5004,N_4748,N_4559);
or U5005 (N_5005,N_4640,N_4471);
nand U5006 (N_5006,N_4464,N_4423);
nor U5007 (N_5007,N_4544,N_4616);
nor U5008 (N_5008,N_4577,N_4468);
xnor U5009 (N_5009,N_4597,N_4591);
nand U5010 (N_5010,N_4794,N_4709);
and U5011 (N_5011,N_4454,N_4437);
xor U5012 (N_5012,N_4563,N_4708);
and U5013 (N_5013,N_4670,N_4564);
and U5014 (N_5014,N_4454,N_4719);
or U5015 (N_5015,N_4799,N_4473);
xor U5016 (N_5016,N_4428,N_4505);
nand U5017 (N_5017,N_4653,N_4727);
or U5018 (N_5018,N_4581,N_4691);
or U5019 (N_5019,N_4548,N_4582);
xnor U5020 (N_5020,N_4615,N_4700);
nor U5021 (N_5021,N_4537,N_4525);
xor U5022 (N_5022,N_4485,N_4486);
nand U5023 (N_5023,N_4581,N_4628);
or U5024 (N_5024,N_4478,N_4763);
and U5025 (N_5025,N_4562,N_4744);
nand U5026 (N_5026,N_4493,N_4451);
nor U5027 (N_5027,N_4502,N_4527);
nand U5028 (N_5028,N_4570,N_4502);
xnor U5029 (N_5029,N_4690,N_4554);
nand U5030 (N_5030,N_4541,N_4750);
or U5031 (N_5031,N_4738,N_4729);
xnor U5032 (N_5032,N_4504,N_4715);
nand U5033 (N_5033,N_4791,N_4747);
nand U5034 (N_5034,N_4788,N_4596);
nand U5035 (N_5035,N_4767,N_4430);
xor U5036 (N_5036,N_4421,N_4787);
xnor U5037 (N_5037,N_4746,N_4450);
and U5038 (N_5038,N_4512,N_4494);
nor U5039 (N_5039,N_4694,N_4547);
nor U5040 (N_5040,N_4720,N_4632);
and U5041 (N_5041,N_4627,N_4728);
and U5042 (N_5042,N_4719,N_4611);
and U5043 (N_5043,N_4539,N_4647);
or U5044 (N_5044,N_4597,N_4453);
or U5045 (N_5045,N_4456,N_4608);
nor U5046 (N_5046,N_4627,N_4662);
nor U5047 (N_5047,N_4517,N_4450);
and U5048 (N_5048,N_4790,N_4738);
xnor U5049 (N_5049,N_4777,N_4415);
nor U5050 (N_5050,N_4536,N_4610);
nor U5051 (N_5051,N_4440,N_4614);
and U5052 (N_5052,N_4645,N_4743);
nand U5053 (N_5053,N_4657,N_4591);
nand U5054 (N_5054,N_4611,N_4484);
nor U5055 (N_5055,N_4518,N_4596);
and U5056 (N_5056,N_4691,N_4576);
or U5057 (N_5057,N_4403,N_4496);
xnor U5058 (N_5058,N_4706,N_4662);
nand U5059 (N_5059,N_4514,N_4769);
and U5060 (N_5060,N_4498,N_4759);
xor U5061 (N_5061,N_4629,N_4409);
and U5062 (N_5062,N_4633,N_4520);
and U5063 (N_5063,N_4526,N_4442);
nand U5064 (N_5064,N_4720,N_4701);
nand U5065 (N_5065,N_4729,N_4566);
nand U5066 (N_5066,N_4712,N_4691);
nor U5067 (N_5067,N_4441,N_4777);
xnor U5068 (N_5068,N_4795,N_4773);
nor U5069 (N_5069,N_4531,N_4505);
xor U5070 (N_5070,N_4551,N_4425);
or U5071 (N_5071,N_4553,N_4640);
or U5072 (N_5072,N_4598,N_4757);
or U5073 (N_5073,N_4542,N_4761);
and U5074 (N_5074,N_4587,N_4574);
or U5075 (N_5075,N_4696,N_4587);
and U5076 (N_5076,N_4452,N_4573);
or U5077 (N_5077,N_4525,N_4449);
nor U5078 (N_5078,N_4405,N_4468);
xnor U5079 (N_5079,N_4666,N_4432);
nor U5080 (N_5080,N_4691,N_4787);
and U5081 (N_5081,N_4786,N_4439);
or U5082 (N_5082,N_4497,N_4582);
nand U5083 (N_5083,N_4789,N_4632);
xor U5084 (N_5084,N_4621,N_4577);
and U5085 (N_5085,N_4649,N_4406);
xor U5086 (N_5086,N_4617,N_4611);
xor U5087 (N_5087,N_4574,N_4731);
nor U5088 (N_5088,N_4593,N_4547);
nor U5089 (N_5089,N_4611,N_4576);
and U5090 (N_5090,N_4643,N_4521);
nor U5091 (N_5091,N_4642,N_4675);
nand U5092 (N_5092,N_4450,N_4561);
and U5093 (N_5093,N_4449,N_4489);
and U5094 (N_5094,N_4521,N_4450);
or U5095 (N_5095,N_4446,N_4432);
xor U5096 (N_5096,N_4488,N_4454);
nand U5097 (N_5097,N_4608,N_4525);
nor U5098 (N_5098,N_4655,N_4709);
nor U5099 (N_5099,N_4728,N_4759);
or U5100 (N_5100,N_4708,N_4727);
and U5101 (N_5101,N_4466,N_4616);
nor U5102 (N_5102,N_4458,N_4775);
and U5103 (N_5103,N_4799,N_4720);
xnor U5104 (N_5104,N_4626,N_4696);
nor U5105 (N_5105,N_4520,N_4540);
and U5106 (N_5106,N_4665,N_4511);
and U5107 (N_5107,N_4735,N_4523);
or U5108 (N_5108,N_4790,N_4563);
nor U5109 (N_5109,N_4683,N_4692);
xor U5110 (N_5110,N_4423,N_4608);
nor U5111 (N_5111,N_4670,N_4759);
nor U5112 (N_5112,N_4660,N_4658);
nor U5113 (N_5113,N_4551,N_4539);
or U5114 (N_5114,N_4627,N_4535);
and U5115 (N_5115,N_4489,N_4700);
or U5116 (N_5116,N_4509,N_4723);
and U5117 (N_5117,N_4472,N_4507);
or U5118 (N_5118,N_4482,N_4449);
nor U5119 (N_5119,N_4414,N_4503);
nor U5120 (N_5120,N_4639,N_4664);
nor U5121 (N_5121,N_4767,N_4545);
nand U5122 (N_5122,N_4642,N_4626);
nand U5123 (N_5123,N_4545,N_4486);
or U5124 (N_5124,N_4578,N_4681);
nand U5125 (N_5125,N_4487,N_4775);
nor U5126 (N_5126,N_4413,N_4798);
nor U5127 (N_5127,N_4589,N_4472);
nand U5128 (N_5128,N_4527,N_4737);
nor U5129 (N_5129,N_4414,N_4794);
nand U5130 (N_5130,N_4758,N_4644);
and U5131 (N_5131,N_4635,N_4538);
and U5132 (N_5132,N_4618,N_4576);
xnor U5133 (N_5133,N_4403,N_4407);
nand U5134 (N_5134,N_4443,N_4735);
or U5135 (N_5135,N_4730,N_4479);
xor U5136 (N_5136,N_4684,N_4712);
and U5137 (N_5137,N_4484,N_4742);
and U5138 (N_5138,N_4679,N_4717);
and U5139 (N_5139,N_4697,N_4429);
and U5140 (N_5140,N_4519,N_4676);
or U5141 (N_5141,N_4680,N_4728);
xnor U5142 (N_5142,N_4787,N_4702);
nand U5143 (N_5143,N_4417,N_4693);
and U5144 (N_5144,N_4749,N_4401);
xor U5145 (N_5145,N_4418,N_4516);
nor U5146 (N_5146,N_4643,N_4602);
or U5147 (N_5147,N_4476,N_4764);
nor U5148 (N_5148,N_4678,N_4664);
or U5149 (N_5149,N_4537,N_4773);
and U5150 (N_5150,N_4774,N_4640);
nor U5151 (N_5151,N_4563,N_4487);
and U5152 (N_5152,N_4690,N_4436);
nand U5153 (N_5153,N_4607,N_4562);
or U5154 (N_5154,N_4760,N_4438);
nand U5155 (N_5155,N_4740,N_4556);
and U5156 (N_5156,N_4715,N_4555);
and U5157 (N_5157,N_4503,N_4545);
and U5158 (N_5158,N_4599,N_4460);
nor U5159 (N_5159,N_4698,N_4560);
or U5160 (N_5160,N_4703,N_4772);
and U5161 (N_5161,N_4705,N_4782);
nand U5162 (N_5162,N_4635,N_4607);
xor U5163 (N_5163,N_4626,N_4689);
xor U5164 (N_5164,N_4774,N_4627);
nor U5165 (N_5165,N_4637,N_4483);
nor U5166 (N_5166,N_4634,N_4759);
xnor U5167 (N_5167,N_4463,N_4493);
nand U5168 (N_5168,N_4651,N_4646);
or U5169 (N_5169,N_4536,N_4611);
nand U5170 (N_5170,N_4403,N_4678);
or U5171 (N_5171,N_4653,N_4744);
or U5172 (N_5172,N_4441,N_4482);
nand U5173 (N_5173,N_4688,N_4722);
or U5174 (N_5174,N_4573,N_4474);
and U5175 (N_5175,N_4598,N_4743);
and U5176 (N_5176,N_4698,N_4591);
and U5177 (N_5177,N_4446,N_4643);
and U5178 (N_5178,N_4648,N_4640);
or U5179 (N_5179,N_4786,N_4487);
or U5180 (N_5180,N_4577,N_4690);
and U5181 (N_5181,N_4570,N_4514);
nand U5182 (N_5182,N_4595,N_4455);
nand U5183 (N_5183,N_4486,N_4441);
nand U5184 (N_5184,N_4530,N_4429);
nand U5185 (N_5185,N_4423,N_4731);
nor U5186 (N_5186,N_4757,N_4623);
or U5187 (N_5187,N_4702,N_4710);
nor U5188 (N_5188,N_4665,N_4504);
xnor U5189 (N_5189,N_4786,N_4534);
or U5190 (N_5190,N_4451,N_4567);
nand U5191 (N_5191,N_4691,N_4690);
nand U5192 (N_5192,N_4550,N_4562);
or U5193 (N_5193,N_4751,N_4460);
or U5194 (N_5194,N_4532,N_4595);
nand U5195 (N_5195,N_4429,N_4730);
nand U5196 (N_5196,N_4747,N_4632);
or U5197 (N_5197,N_4609,N_4434);
or U5198 (N_5198,N_4646,N_4488);
and U5199 (N_5199,N_4636,N_4702);
or U5200 (N_5200,N_5091,N_4880);
nand U5201 (N_5201,N_5110,N_4984);
xnor U5202 (N_5202,N_4967,N_4914);
nand U5203 (N_5203,N_4834,N_4823);
nand U5204 (N_5204,N_4839,N_5192);
or U5205 (N_5205,N_5171,N_4923);
nand U5206 (N_5206,N_4864,N_4850);
or U5207 (N_5207,N_4819,N_4995);
and U5208 (N_5208,N_4884,N_5198);
nand U5209 (N_5209,N_4997,N_5071);
and U5210 (N_5210,N_4887,N_5056);
or U5211 (N_5211,N_4856,N_5082);
nor U5212 (N_5212,N_4961,N_4820);
or U5213 (N_5213,N_5008,N_4872);
and U5214 (N_5214,N_4845,N_4902);
xnor U5215 (N_5215,N_4917,N_5013);
nor U5216 (N_5216,N_5190,N_4949);
and U5217 (N_5217,N_4915,N_4951);
xnor U5218 (N_5218,N_4958,N_5048);
nor U5219 (N_5219,N_4867,N_4925);
nor U5220 (N_5220,N_5009,N_4855);
or U5221 (N_5221,N_4927,N_5076);
and U5222 (N_5222,N_5191,N_4810);
xor U5223 (N_5223,N_4806,N_5124);
and U5224 (N_5224,N_5093,N_5040);
or U5225 (N_5225,N_4905,N_4965);
xor U5226 (N_5226,N_5141,N_5011);
and U5227 (N_5227,N_4975,N_5032);
nand U5228 (N_5228,N_4926,N_5080);
nor U5229 (N_5229,N_5084,N_4950);
xor U5230 (N_5230,N_5025,N_5033);
nor U5231 (N_5231,N_5142,N_5024);
and U5232 (N_5232,N_5151,N_5144);
nor U5233 (N_5233,N_4874,N_4896);
xnor U5234 (N_5234,N_4893,N_5061);
xnor U5235 (N_5235,N_5128,N_5062);
xor U5236 (N_5236,N_4817,N_5022);
nor U5237 (N_5237,N_5012,N_5030);
and U5238 (N_5238,N_5006,N_5098);
nor U5239 (N_5239,N_5027,N_4921);
or U5240 (N_5240,N_4930,N_5109);
and U5241 (N_5241,N_4828,N_4957);
and U5242 (N_5242,N_5114,N_5175);
or U5243 (N_5243,N_5156,N_4999);
and U5244 (N_5244,N_5010,N_4912);
nor U5245 (N_5245,N_4816,N_4898);
nand U5246 (N_5246,N_4968,N_5193);
nand U5247 (N_5247,N_5060,N_4919);
xor U5248 (N_5248,N_4899,N_4888);
xor U5249 (N_5249,N_4844,N_4897);
and U5250 (N_5250,N_5150,N_4859);
nand U5251 (N_5251,N_4939,N_4871);
or U5252 (N_5252,N_5184,N_5072);
and U5253 (N_5253,N_4849,N_5137);
nand U5254 (N_5254,N_4824,N_5070);
or U5255 (N_5255,N_5099,N_4848);
nor U5256 (N_5256,N_5196,N_5058);
nand U5257 (N_5257,N_5169,N_4895);
nor U5258 (N_5258,N_4945,N_5115);
xor U5259 (N_5259,N_5105,N_4983);
xnor U5260 (N_5260,N_5131,N_4916);
xnor U5261 (N_5261,N_4875,N_4885);
and U5262 (N_5262,N_5152,N_4970);
or U5263 (N_5263,N_5102,N_4838);
or U5264 (N_5264,N_4802,N_5026);
or U5265 (N_5265,N_4944,N_5132);
xnor U5266 (N_5266,N_5019,N_5155);
and U5267 (N_5267,N_5185,N_5118);
and U5268 (N_5268,N_4803,N_5077);
and U5269 (N_5269,N_4988,N_5004);
xor U5270 (N_5270,N_5090,N_5135);
xor U5271 (N_5271,N_5016,N_4931);
or U5272 (N_5272,N_5015,N_4842);
nor U5273 (N_5273,N_4989,N_4889);
xnor U5274 (N_5274,N_5199,N_4811);
nor U5275 (N_5275,N_5020,N_4805);
and U5276 (N_5276,N_5126,N_5074);
nand U5277 (N_5277,N_4869,N_5167);
nand U5278 (N_5278,N_5069,N_4966);
and U5279 (N_5279,N_4994,N_4807);
and U5280 (N_5280,N_4815,N_4801);
or U5281 (N_5281,N_5139,N_5174);
or U5282 (N_5282,N_4933,N_4960);
xor U5283 (N_5283,N_5063,N_5170);
or U5284 (N_5284,N_4809,N_4831);
xor U5285 (N_5285,N_4863,N_4808);
nand U5286 (N_5286,N_4892,N_4920);
nand U5287 (N_5287,N_4903,N_5089);
xnor U5288 (N_5288,N_4913,N_5017);
xor U5289 (N_5289,N_5112,N_4821);
or U5290 (N_5290,N_4936,N_5168);
nand U5291 (N_5291,N_4929,N_4907);
nor U5292 (N_5292,N_5140,N_4846);
nor U5293 (N_5293,N_5014,N_4900);
nand U5294 (N_5294,N_4977,N_5050);
or U5295 (N_5295,N_5057,N_4964);
and U5296 (N_5296,N_5172,N_4861);
or U5297 (N_5297,N_5041,N_4987);
and U5298 (N_5298,N_5001,N_4868);
nor U5299 (N_5299,N_5146,N_4878);
nand U5300 (N_5300,N_4934,N_4942);
xnor U5301 (N_5301,N_5038,N_5195);
xnor U5302 (N_5302,N_4948,N_5085);
and U5303 (N_5303,N_5134,N_5127);
nand U5304 (N_5304,N_4873,N_4937);
nand U5305 (N_5305,N_4904,N_5037);
and U5306 (N_5306,N_5163,N_5073);
xor U5307 (N_5307,N_5164,N_5103);
nand U5308 (N_5308,N_5104,N_5176);
xor U5309 (N_5309,N_4996,N_4860);
nor U5310 (N_5310,N_5180,N_4857);
xnor U5311 (N_5311,N_5194,N_5097);
and U5312 (N_5312,N_5083,N_4865);
or U5313 (N_5313,N_5181,N_4827);
xnor U5314 (N_5314,N_5122,N_4911);
and U5315 (N_5315,N_4890,N_4894);
or U5316 (N_5316,N_4955,N_5160);
or U5317 (N_5317,N_4883,N_5094);
xnor U5318 (N_5318,N_5107,N_4974);
nand U5319 (N_5319,N_5149,N_4947);
nor U5320 (N_5320,N_5120,N_4851);
nand U5321 (N_5321,N_4969,N_5079);
nor U5322 (N_5322,N_4858,N_4829);
or U5323 (N_5323,N_5054,N_5148);
nand U5324 (N_5324,N_5125,N_4998);
or U5325 (N_5325,N_5007,N_4876);
and U5326 (N_5326,N_5049,N_5052);
nand U5327 (N_5327,N_5034,N_4990);
nor U5328 (N_5328,N_4836,N_5035);
nand U5329 (N_5329,N_5182,N_4901);
and U5330 (N_5330,N_5162,N_5119);
xor U5331 (N_5331,N_4918,N_5096);
nand U5332 (N_5332,N_5117,N_4832);
nand U5333 (N_5333,N_4826,N_4908);
xnor U5334 (N_5334,N_5130,N_5183);
and U5335 (N_5335,N_4813,N_5088);
or U5336 (N_5336,N_4870,N_5045);
nor U5337 (N_5337,N_5157,N_4910);
nand U5338 (N_5338,N_4954,N_5095);
and U5339 (N_5339,N_5147,N_5179);
or U5340 (N_5340,N_5039,N_4976);
xor U5341 (N_5341,N_5101,N_5018);
nand U5342 (N_5342,N_4979,N_5068);
xnor U5343 (N_5343,N_5100,N_5047);
xnor U5344 (N_5344,N_4978,N_4959);
nor U5345 (N_5345,N_5121,N_5178);
xor U5346 (N_5346,N_4924,N_5087);
or U5347 (N_5347,N_4822,N_4804);
nand U5348 (N_5348,N_4941,N_5166);
xor U5349 (N_5349,N_4991,N_4835);
xor U5350 (N_5350,N_4818,N_5031);
nor U5351 (N_5351,N_4843,N_5066);
xor U5352 (N_5352,N_5055,N_5002);
nand U5353 (N_5353,N_4963,N_4891);
xor U5354 (N_5354,N_5189,N_5108);
and U5355 (N_5355,N_5078,N_4812);
nor U5356 (N_5356,N_5106,N_4922);
or U5357 (N_5357,N_5092,N_4962);
and U5358 (N_5358,N_5029,N_4886);
and U5359 (N_5359,N_4993,N_5116);
or U5360 (N_5360,N_5043,N_5005);
or U5361 (N_5361,N_5123,N_5161);
nor U5362 (N_5362,N_5133,N_5138);
nand U5363 (N_5363,N_4909,N_4986);
nor U5364 (N_5364,N_5044,N_5197);
or U5365 (N_5365,N_5053,N_5111);
nor U5366 (N_5366,N_4980,N_4877);
xnor U5367 (N_5367,N_5075,N_5143);
nand U5368 (N_5368,N_4847,N_4938);
nor U5369 (N_5369,N_4830,N_5046);
nand U5370 (N_5370,N_4862,N_5021);
and U5371 (N_5371,N_5136,N_4932);
or U5372 (N_5372,N_5113,N_5036);
and U5373 (N_5373,N_5000,N_4935);
or U5374 (N_5374,N_5177,N_5186);
and U5375 (N_5375,N_5188,N_4956);
xor U5376 (N_5376,N_5165,N_5158);
or U5377 (N_5377,N_4800,N_5064);
nand U5378 (N_5378,N_5051,N_4854);
nand U5379 (N_5379,N_4981,N_4866);
nor U5380 (N_5380,N_5153,N_4833);
and U5381 (N_5381,N_4940,N_4837);
nand U5382 (N_5382,N_5159,N_5028);
xor U5383 (N_5383,N_4992,N_5086);
xor U5384 (N_5384,N_5067,N_5154);
or U5385 (N_5385,N_5145,N_4879);
or U5386 (N_5386,N_4953,N_4982);
or U5387 (N_5387,N_4946,N_5003);
nand U5388 (N_5388,N_4852,N_4985);
xnor U5389 (N_5389,N_4973,N_4971);
and U5390 (N_5390,N_4825,N_4972);
xnor U5391 (N_5391,N_4841,N_4928);
or U5392 (N_5392,N_5173,N_5023);
nor U5393 (N_5393,N_4840,N_5081);
nor U5394 (N_5394,N_4906,N_4943);
nor U5395 (N_5395,N_4814,N_4952);
and U5396 (N_5396,N_5129,N_4881);
or U5397 (N_5397,N_5059,N_4882);
xnor U5398 (N_5398,N_5042,N_5187);
xnor U5399 (N_5399,N_4853,N_5065);
xnor U5400 (N_5400,N_4987,N_4970);
or U5401 (N_5401,N_4907,N_5162);
xor U5402 (N_5402,N_4988,N_5106);
and U5403 (N_5403,N_4966,N_4897);
nor U5404 (N_5404,N_5053,N_5147);
nand U5405 (N_5405,N_4970,N_4852);
nor U5406 (N_5406,N_4878,N_4867);
nor U5407 (N_5407,N_5188,N_4832);
nor U5408 (N_5408,N_5025,N_5197);
nand U5409 (N_5409,N_4984,N_5101);
or U5410 (N_5410,N_4842,N_4844);
or U5411 (N_5411,N_4834,N_5065);
and U5412 (N_5412,N_5160,N_5085);
and U5413 (N_5413,N_4872,N_4851);
nor U5414 (N_5414,N_4960,N_4852);
xor U5415 (N_5415,N_5072,N_4828);
or U5416 (N_5416,N_5010,N_4885);
xor U5417 (N_5417,N_4895,N_5111);
nand U5418 (N_5418,N_5042,N_4848);
nor U5419 (N_5419,N_5012,N_5190);
or U5420 (N_5420,N_4898,N_4894);
nor U5421 (N_5421,N_4825,N_4839);
nand U5422 (N_5422,N_4829,N_5119);
nor U5423 (N_5423,N_4867,N_5122);
and U5424 (N_5424,N_4932,N_5079);
and U5425 (N_5425,N_5059,N_5034);
and U5426 (N_5426,N_5174,N_4805);
nor U5427 (N_5427,N_4892,N_4976);
xnor U5428 (N_5428,N_5117,N_4987);
xnor U5429 (N_5429,N_4977,N_5100);
and U5430 (N_5430,N_5177,N_5192);
or U5431 (N_5431,N_4974,N_4983);
xnor U5432 (N_5432,N_4990,N_4846);
nand U5433 (N_5433,N_5009,N_4969);
nor U5434 (N_5434,N_4990,N_5169);
nor U5435 (N_5435,N_4860,N_4941);
nand U5436 (N_5436,N_4948,N_5077);
or U5437 (N_5437,N_4942,N_5173);
nand U5438 (N_5438,N_5171,N_5089);
or U5439 (N_5439,N_4802,N_5104);
or U5440 (N_5440,N_5166,N_5087);
or U5441 (N_5441,N_4899,N_5077);
and U5442 (N_5442,N_5165,N_5013);
nand U5443 (N_5443,N_5071,N_4815);
and U5444 (N_5444,N_4960,N_4943);
nor U5445 (N_5445,N_4947,N_5021);
or U5446 (N_5446,N_5079,N_4971);
nand U5447 (N_5447,N_5048,N_4902);
nand U5448 (N_5448,N_4941,N_4969);
or U5449 (N_5449,N_4997,N_5039);
or U5450 (N_5450,N_5181,N_5174);
nor U5451 (N_5451,N_5062,N_5071);
or U5452 (N_5452,N_5185,N_4942);
nand U5453 (N_5453,N_5090,N_5071);
or U5454 (N_5454,N_5020,N_4950);
nor U5455 (N_5455,N_5111,N_4807);
nor U5456 (N_5456,N_4801,N_5036);
or U5457 (N_5457,N_5108,N_4904);
xor U5458 (N_5458,N_4820,N_5142);
and U5459 (N_5459,N_5131,N_5196);
xnor U5460 (N_5460,N_5007,N_4990);
or U5461 (N_5461,N_4810,N_5137);
xnor U5462 (N_5462,N_4891,N_5115);
nand U5463 (N_5463,N_4901,N_5147);
or U5464 (N_5464,N_5020,N_5048);
nor U5465 (N_5465,N_5055,N_5080);
xnor U5466 (N_5466,N_5010,N_5065);
nor U5467 (N_5467,N_4847,N_4822);
and U5468 (N_5468,N_4873,N_5035);
nor U5469 (N_5469,N_4813,N_5058);
and U5470 (N_5470,N_5057,N_4978);
xor U5471 (N_5471,N_5107,N_4868);
nor U5472 (N_5472,N_5012,N_4981);
nand U5473 (N_5473,N_4905,N_5164);
nor U5474 (N_5474,N_4969,N_5176);
and U5475 (N_5475,N_5144,N_5052);
nor U5476 (N_5476,N_5118,N_4872);
xnor U5477 (N_5477,N_4927,N_4959);
or U5478 (N_5478,N_5151,N_5116);
nor U5479 (N_5479,N_4974,N_5124);
or U5480 (N_5480,N_5100,N_5108);
or U5481 (N_5481,N_4940,N_4926);
nor U5482 (N_5482,N_4960,N_5163);
nor U5483 (N_5483,N_5095,N_5052);
nor U5484 (N_5484,N_4847,N_4805);
or U5485 (N_5485,N_5151,N_4805);
xor U5486 (N_5486,N_4891,N_5040);
nor U5487 (N_5487,N_4978,N_5152);
nand U5488 (N_5488,N_4887,N_5157);
nor U5489 (N_5489,N_5016,N_5095);
nand U5490 (N_5490,N_5160,N_5028);
xnor U5491 (N_5491,N_5082,N_4860);
xnor U5492 (N_5492,N_5063,N_4960);
xnor U5493 (N_5493,N_4970,N_4892);
or U5494 (N_5494,N_4838,N_5035);
or U5495 (N_5495,N_5078,N_4806);
xor U5496 (N_5496,N_4931,N_4934);
or U5497 (N_5497,N_5145,N_5100);
nor U5498 (N_5498,N_5076,N_4865);
and U5499 (N_5499,N_5112,N_4893);
and U5500 (N_5500,N_4814,N_5012);
nor U5501 (N_5501,N_5136,N_5038);
nand U5502 (N_5502,N_4912,N_5070);
nor U5503 (N_5503,N_5115,N_5021);
nand U5504 (N_5504,N_5129,N_5139);
or U5505 (N_5505,N_4945,N_4937);
and U5506 (N_5506,N_4907,N_4928);
xor U5507 (N_5507,N_4958,N_5029);
xnor U5508 (N_5508,N_4846,N_4887);
nand U5509 (N_5509,N_4839,N_5101);
nor U5510 (N_5510,N_5108,N_4970);
or U5511 (N_5511,N_5177,N_5176);
nand U5512 (N_5512,N_4917,N_4817);
xor U5513 (N_5513,N_5068,N_5051);
nand U5514 (N_5514,N_5190,N_4986);
nor U5515 (N_5515,N_5127,N_4880);
nor U5516 (N_5516,N_5178,N_4866);
nand U5517 (N_5517,N_5011,N_4870);
xnor U5518 (N_5518,N_5007,N_4921);
and U5519 (N_5519,N_4850,N_5147);
and U5520 (N_5520,N_5024,N_5041);
nor U5521 (N_5521,N_5052,N_4975);
xor U5522 (N_5522,N_5088,N_4905);
nand U5523 (N_5523,N_4936,N_5024);
xnor U5524 (N_5524,N_5126,N_4981);
nor U5525 (N_5525,N_5191,N_5162);
nand U5526 (N_5526,N_5024,N_4946);
nor U5527 (N_5527,N_5095,N_4962);
xor U5528 (N_5528,N_4824,N_4959);
nor U5529 (N_5529,N_4870,N_5085);
xnor U5530 (N_5530,N_4974,N_4829);
xnor U5531 (N_5531,N_5193,N_5058);
nor U5532 (N_5532,N_4876,N_4889);
and U5533 (N_5533,N_5172,N_5005);
nand U5534 (N_5534,N_5183,N_4944);
xor U5535 (N_5535,N_5195,N_4899);
and U5536 (N_5536,N_5005,N_5114);
or U5537 (N_5537,N_5119,N_5165);
xnor U5538 (N_5538,N_4968,N_4999);
or U5539 (N_5539,N_5044,N_5146);
and U5540 (N_5540,N_5129,N_5188);
nand U5541 (N_5541,N_5193,N_4975);
nand U5542 (N_5542,N_5139,N_4941);
and U5543 (N_5543,N_5161,N_5158);
and U5544 (N_5544,N_5051,N_4885);
xor U5545 (N_5545,N_5114,N_5025);
or U5546 (N_5546,N_5002,N_5110);
xor U5547 (N_5547,N_4923,N_5022);
or U5548 (N_5548,N_4901,N_5157);
or U5549 (N_5549,N_4810,N_5030);
nor U5550 (N_5550,N_4847,N_4802);
or U5551 (N_5551,N_4902,N_4945);
and U5552 (N_5552,N_5152,N_5111);
nand U5553 (N_5553,N_5002,N_4972);
nand U5554 (N_5554,N_4979,N_5028);
nand U5555 (N_5555,N_5033,N_4834);
or U5556 (N_5556,N_4888,N_4986);
and U5557 (N_5557,N_5182,N_4871);
nand U5558 (N_5558,N_4808,N_4999);
or U5559 (N_5559,N_5042,N_4835);
nor U5560 (N_5560,N_5067,N_4890);
nor U5561 (N_5561,N_5071,N_5196);
or U5562 (N_5562,N_5140,N_4890);
nor U5563 (N_5563,N_4880,N_4841);
or U5564 (N_5564,N_5199,N_4901);
xnor U5565 (N_5565,N_4993,N_5030);
and U5566 (N_5566,N_4980,N_4974);
and U5567 (N_5567,N_4840,N_5106);
and U5568 (N_5568,N_5143,N_4813);
and U5569 (N_5569,N_4832,N_4924);
xnor U5570 (N_5570,N_5066,N_5116);
xnor U5571 (N_5571,N_5004,N_5097);
and U5572 (N_5572,N_5025,N_5171);
nand U5573 (N_5573,N_4936,N_4950);
or U5574 (N_5574,N_5122,N_4843);
or U5575 (N_5575,N_4809,N_5108);
xnor U5576 (N_5576,N_4903,N_5132);
or U5577 (N_5577,N_4835,N_4918);
nor U5578 (N_5578,N_5014,N_4811);
nand U5579 (N_5579,N_4959,N_5051);
nor U5580 (N_5580,N_4890,N_4995);
or U5581 (N_5581,N_5186,N_4866);
or U5582 (N_5582,N_4925,N_5038);
and U5583 (N_5583,N_4853,N_5012);
xor U5584 (N_5584,N_4878,N_5119);
xor U5585 (N_5585,N_4969,N_4905);
nor U5586 (N_5586,N_4962,N_5056);
xor U5587 (N_5587,N_5162,N_4833);
nor U5588 (N_5588,N_5182,N_5093);
xor U5589 (N_5589,N_5077,N_4980);
nor U5590 (N_5590,N_4910,N_5015);
nand U5591 (N_5591,N_5157,N_4927);
and U5592 (N_5592,N_5060,N_5080);
nor U5593 (N_5593,N_4845,N_4975);
xnor U5594 (N_5594,N_5161,N_5034);
or U5595 (N_5595,N_5159,N_4979);
nand U5596 (N_5596,N_4828,N_4988);
xnor U5597 (N_5597,N_4995,N_4892);
or U5598 (N_5598,N_5004,N_5123);
and U5599 (N_5599,N_4874,N_4969);
and U5600 (N_5600,N_5228,N_5386);
xor U5601 (N_5601,N_5227,N_5316);
xnor U5602 (N_5602,N_5575,N_5354);
nor U5603 (N_5603,N_5296,N_5422);
nand U5604 (N_5604,N_5405,N_5390);
and U5605 (N_5605,N_5303,N_5500);
nor U5606 (N_5606,N_5557,N_5524);
nand U5607 (N_5607,N_5495,N_5514);
or U5608 (N_5608,N_5361,N_5291);
or U5609 (N_5609,N_5398,N_5211);
and U5610 (N_5610,N_5200,N_5219);
xor U5611 (N_5611,N_5490,N_5574);
or U5612 (N_5612,N_5353,N_5203);
and U5613 (N_5613,N_5262,N_5502);
xnor U5614 (N_5614,N_5310,N_5389);
xnor U5615 (N_5615,N_5275,N_5463);
nor U5616 (N_5616,N_5446,N_5244);
nor U5617 (N_5617,N_5335,N_5285);
nand U5618 (N_5618,N_5309,N_5538);
nand U5619 (N_5619,N_5572,N_5481);
nand U5620 (N_5620,N_5434,N_5245);
and U5621 (N_5621,N_5284,N_5237);
nand U5622 (N_5622,N_5480,N_5469);
nor U5623 (N_5623,N_5512,N_5370);
and U5624 (N_5624,N_5213,N_5358);
or U5625 (N_5625,N_5451,N_5475);
nor U5626 (N_5626,N_5493,N_5421);
or U5627 (N_5627,N_5461,N_5295);
and U5628 (N_5628,N_5242,N_5371);
and U5629 (N_5629,N_5334,N_5224);
xor U5630 (N_5630,N_5388,N_5263);
nor U5631 (N_5631,N_5553,N_5207);
nor U5632 (N_5632,N_5438,N_5464);
nor U5633 (N_5633,N_5444,N_5397);
xnor U5634 (N_5634,N_5276,N_5594);
nor U5635 (N_5635,N_5513,N_5328);
nor U5636 (N_5636,N_5202,N_5487);
xor U5637 (N_5637,N_5235,N_5427);
and U5638 (N_5638,N_5544,N_5445);
nand U5639 (N_5639,N_5570,N_5364);
or U5640 (N_5640,N_5217,N_5474);
xnor U5641 (N_5641,N_5406,N_5453);
nand U5642 (N_5642,N_5356,N_5560);
nand U5643 (N_5643,N_5431,N_5530);
nor U5644 (N_5644,N_5561,N_5322);
xnor U5645 (N_5645,N_5331,N_5515);
or U5646 (N_5646,N_5349,N_5404);
and U5647 (N_5647,N_5230,N_5326);
nor U5648 (N_5648,N_5441,N_5576);
nor U5649 (N_5649,N_5551,N_5332);
nor U5650 (N_5650,N_5343,N_5344);
or U5651 (N_5651,N_5348,N_5563);
or U5652 (N_5652,N_5411,N_5271);
nor U5653 (N_5653,N_5267,N_5206);
nor U5654 (N_5654,N_5457,N_5430);
xor U5655 (N_5655,N_5279,N_5414);
xor U5656 (N_5656,N_5496,N_5266);
nor U5657 (N_5657,N_5450,N_5379);
xnor U5658 (N_5658,N_5392,N_5257);
nor U5659 (N_5659,N_5545,N_5448);
and U5660 (N_5660,N_5467,N_5523);
xnor U5661 (N_5661,N_5247,N_5240);
or U5662 (N_5662,N_5525,N_5598);
xor U5663 (N_5663,N_5297,N_5208);
or U5664 (N_5664,N_5582,N_5304);
nand U5665 (N_5665,N_5527,N_5290);
xnor U5666 (N_5666,N_5306,N_5340);
and U5667 (N_5667,N_5516,N_5375);
nand U5668 (N_5668,N_5483,N_5599);
or U5669 (N_5669,N_5373,N_5568);
nor U5670 (N_5670,N_5540,N_5505);
nor U5671 (N_5671,N_5550,N_5565);
nor U5672 (N_5672,N_5229,N_5471);
or U5673 (N_5673,N_5204,N_5320);
or U5674 (N_5674,N_5201,N_5314);
or U5675 (N_5675,N_5250,N_5269);
nor U5676 (N_5676,N_5393,N_5399);
nand U5677 (N_5677,N_5577,N_5278);
nor U5678 (N_5678,N_5462,N_5417);
and U5679 (N_5679,N_5341,N_5590);
xor U5680 (N_5680,N_5367,N_5368);
or U5681 (N_5681,N_5221,N_5564);
or U5682 (N_5682,N_5491,N_5531);
xor U5683 (N_5683,N_5482,N_5503);
nor U5684 (N_5684,N_5347,N_5433);
xnor U5685 (N_5685,N_5486,N_5508);
nor U5686 (N_5686,N_5336,N_5258);
or U5687 (N_5687,N_5330,N_5359);
and U5688 (N_5688,N_5401,N_5528);
nand U5689 (N_5689,N_5232,N_5289);
nand U5690 (N_5690,N_5272,N_5579);
nand U5691 (N_5691,N_5324,N_5350);
nand U5692 (N_5692,N_5548,N_5473);
and U5693 (N_5693,N_5281,N_5223);
xor U5694 (N_5694,N_5466,N_5408);
nand U5695 (N_5695,N_5246,N_5562);
xor U5696 (N_5696,N_5585,N_5479);
nand U5697 (N_5697,N_5308,N_5292);
and U5698 (N_5698,N_5384,N_5209);
nand U5699 (N_5699,N_5345,N_5311);
nand U5700 (N_5700,N_5249,N_5225);
nand U5701 (N_5701,N_5355,N_5552);
xnor U5702 (N_5702,N_5442,N_5363);
nor U5703 (N_5703,N_5299,N_5456);
xnor U5704 (N_5704,N_5301,N_5534);
xor U5705 (N_5705,N_5239,N_5243);
or U5706 (N_5706,N_5597,N_5477);
nor U5707 (N_5707,N_5520,N_5254);
nor U5708 (N_5708,N_5317,N_5425);
nor U5709 (N_5709,N_5423,N_5259);
nor U5710 (N_5710,N_5333,N_5318);
or U5711 (N_5711,N_5468,N_5584);
and U5712 (N_5712,N_5327,N_5329);
and U5713 (N_5713,N_5380,N_5220);
nand U5714 (N_5714,N_5573,N_5248);
nor U5715 (N_5715,N_5378,N_5218);
nor U5716 (N_5716,N_5286,N_5385);
and U5717 (N_5717,N_5455,N_5492);
and U5718 (N_5718,N_5436,N_5494);
nor U5719 (N_5719,N_5537,N_5415);
xnor U5720 (N_5720,N_5287,N_5533);
and U5721 (N_5721,N_5305,N_5539);
xnor U5722 (N_5722,N_5460,N_5409);
or U5723 (N_5723,N_5578,N_5268);
nand U5724 (N_5724,N_5592,N_5391);
or U5725 (N_5725,N_5546,N_5300);
nor U5726 (N_5726,N_5352,N_5591);
xor U5727 (N_5727,N_5497,N_5382);
or U5728 (N_5728,N_5458,N_5569);
or U5729 (N_5729,N_5499,N_5261);
nor U5730 (N_5730,N_5360,N_5319);
or U5731 (N_5731,N_5396,N_5222);
nor U5732 (N_5732,N_5383,N_5435);
xnor U5733 (N_5733,N_5325,N_5315);
and U5734 (N_5734,N_5419,N_5372);
or U5735 (N_5735,N_5412,N_5264);
nand U5736 (N_5736,N_5559,N_5484);
xnor U5737 (N_5737,N_5277,N_5472);
or U5738 (N_5738,N_5443,N_5426);
xor U5739 (N_5739,N_5231,N_5233);
and U5740 (N_5740,N_5596,N_5357);
nand U5741 (N_5741,N_5588,N_5234);
nor U5742 (N_5742,N_5216,N_5407);
or U5743 (N_5743,N_5519,N_5256);
nand U5744 (N_5744,N_5459,N_5418);
xor U5745 (N_5745,N_5449,N_5470);
nor U5746 (N_5746,N_5205,N_5252);
and U5747 (N_5747,N_5273,N_5294);
or U5748 (N_5748,N_5529,N_5581);
or U5749 (N_5749,N_5589,N_5571);
nor U5750 (N_5750,N_5447,N_5413);
and U5751 (N_5751,N_5346,N_5476);
nand U5752 (N_5752,N_5509,N_5593);
xnor U5753 (N_5753,N_5238,N_5526);
and U5754 (N_5754,N_5511,N_5362);
nor U5755 (N_5755,N_5270,N_5283);
nand U5756 (N_5756,N_5416,N_5226);
nor U5757 (N_5757,N_5339,N_5323);
or U5758 (N_5758,N_5387,N_5522);
xnor U5759 (N_5759,N_5432,N_5517);
or U5760 (N_5760,N_5440,N_5549);
nand U5761 (N_5761,N_5376,N_5452);
nand U5762 (N_5762,N_5583,N_5402);
nor U5763 (N_5763,N_5410,N_5282);
xor U5764 (N_5764,N_5595,N_5394);
xor U5765 (N_5765,N_5420,N_5307);
nor U5766 (N_5766,N_5542,N_5321);
xnor U5767 (N_5767,N_5381,N_5337);
and U5768 (N_5768,N_5554,N_5251);
and U5769 (N_5769,N_5365,N_5506);
and U5770 (N_5770,N_5543,N_5260);
or U5771 (N_5771,N_5501,N_5498);
nand U5772 (N_5772,N_5338,N_5567);
nor U5773 (N_5773,N_5555,N_5236);
and U5774 (N_5774,N_5439,N_5510);
nand U5775 (N_5775,N_5265,N_5424);
nor U5776 (N_5776,N_5366,N_5298);
or U5777 (N_5777,N_5429,N_5478);
xnor U5778 (N_5778,N_5288,N_5465);
xnor U5779 (N_5779,N_5566,N_5403);
xor U5780 (N_5780,N_5302,N_5255);
xnor U5781 (N_5781,N_5374,N_5536);
nor U5782 (N_5782,N_5437,N_5241);
nand U5783 (N_5783,N_5586,N_5587);
nor U5784 (N_5784,N_5312,N_5580);
xor U5785 (N_5785,N_5504,N_5313);
and U5786 (N_5786,N_5369,N_5215);
xor U5787 (N_5787,N_5280,N_5210);
or U5788 (N_5788,N_5395,N_5377);
nand U5789 (N_5789,N_5351,N_5214);
nand U5790 (N_5790,N_5507,N_5454);
or U5791 (N_5791,N_5342,N_5488);
nor U5792 (N_5792,N_5253,N_5485);
nand U5793 (N_5793,N_5547,N_5541);
and U5794 (N_5794,N_5489,N_5518);
and U5795 (N_5795,N_5293,N_5274);
xnor U5796 (N_5796,N_5535,N_5558);
and U5797 (N_5797,N_5556,N_5428);
xor U5798 (N_5798,N_5400,N_5521);
xnor U5799 (N_5799,N_5212,N_5532);
nand U5800 (N_5800,N_5447,N_5572);
nand U5801 (N_5801,N_5552,N_5527);
xnor U5802 (N_5802,N_5303,N_5475);
nor U5803 (N_5803,N_5475,N_5382);
nand U5804 (N_5804,N_5261,N_5568);
and U5805 (N_5805,N_5527,N_5239);
nand U5806 (N_5806,N_5395,N_5355);
and U5807 (N_5807,N_5588,N_5514);
nor U5808 (N_5808,N_5427,N_5370);
nand U5809 (N_5809,N_5572,N_5501);
nor U5810 (N_5810,N_5405,N_5268);
nor U5811 (N_5811,N_5383,N_5379);
and U5812 (N_5812,N_5590,N_5294);
nor U5813 (N_5813,N_5444,N_5322);
or U5814 (N_5814,N_5409,N_5221);
nand U5815 (N_5815,N_5585,N_5448);
nor U5816 (N_5816,N_5520,N_5305);
nand U5817 (N_5817,N_5407,N_5432);
nand U5818 (N_5818,N_5538,N_5583);
and U5819 (N_5819,N_5265,N_5302);
xnor U5820 (N_5820,N_5567,N_5550);
xor U5821 (N_5821,N_5385,N_5452);
nand U5822 (N_5822,N_5564,N_5230);
xnor U5823 (N_5823,N_5332,N_5369);
xnor U5824 (N_5824,N_5489,N_5202);
or U5825 (N_5825,N_5288,N_5244);
and U5826 (N_5826,N_5384,N_5217);
xor U5827 (N_5827,N_5569,N_5251);
nor U5828 (N_5828,N_5596,N_5381);
nor U5829 (N_5829,N_5561,N_5245);
and U5830 (N_5830,N_5246,N_5474);
and U5831 (N_5831,N_5518,N_5229);
and U5832 (N_5832,N_5200,N_5218);
or U5833 (N_5833,N_5567,N_5523);
nor U5834 (N_5834,N_5334,N_5388);
and U5835 (N_5835,N_5436,N_5552);
nand U5836 (N_5836,N_5205,N_5450);
or U5837 (N_5837,N_5397,N_5565);
nand U5838 (N_5838,N_5596,N_5251);
nor U5839 (N_5839,N_5329,N_5201);
or U5840 (N_5840,N_5218,N_5206);
and U5841 (N_5841,N_5523,N_5566);
nor U5842 (N_5842,N_5248,N_5531);
nand U5843 (N_5843,N_5204,N_5488);
nor U5844 (N_5844,N_5369,N_5465);
xor U5845 (N_5845,N_5598,N_5415);
and U5846 (N_5846,N_5448,N_5497);
or U5847 (N_5847,N_5381,N_5561);
and U5848 (N_5848,N_5223,N_5383);
nor U5849 (N_5849,N_5486,N_5419);
and U5850 (N_5850,N_5298,N_5386);
nor U5851 (N_5851,N_5507,N_5276);
and U5852 (N_5852,N_5583,N_5251);
or U5853 (N_5853,N_5385,N_5372);
nor U5854 (N_5854,N_5412,N_5329);
or U5855 (N_5855,N_5544,N_5378);
or U5856 (N_5856,N_5474,N_5441);
or U5857 (N_5857,N_5242,N_5391);
nor U5858 (N_5858,N_5476,N_5556);
and U5859 (N_5859,N_5552,N_5385);
xnor U5860 (N_5860,N_5572,N_5471);
nor U5861 (N_5861,N_5397,N_5552);
nor U5862 (N_5862,N_5534,N_5549);
xnor U5863 (N_5863,N_5526,N_5593);
or U5864 (N_5864,N_5346,N_5588);
nor U5865 (N_5865,N_5311,N_5575);
nor U5866 (N_5866,N_5285,N_5337);
or U5867 (N_5867,N_5580,N_5285);
nand U5868 (N_5868,N_5227,N_5235);
and U5869 (N_5869,N_5489,N_5280);
nand U5870 (N_5870,N_5567,N_5202);
nand U5871 (N_5871,N_5483,N_5397);
nand U5872 (N_5872,N_5400,N_5209);
or U5873 (N_5873,N_5306,N_5253);
and U5874 (N_5874,N_5240,N_5558);
or U5875 (N_5875,N_5548,N_5459);
nand U5876 (N_5876,N_5440,N_5414);
xor U5877 (N_5877,N_5368,N_5563);
xor U5878 (N_5878,N_5570,N_5210);
and U5879 (N_5879,N_5577,N_5392);
xnor U5880 (N_5880,N_5419,N_5327);
or U5881 (N_5881,N_5434,N_5483);
nand U5882 (N_5882,N_5440,N_5401);
nor U5883 (N_5883,N_5389,N_5254);
xnor U5884 (N_5884,N_5420,N_5488);
nor U5885 (N_5885,N_5370,N_5305);
nor U5886 (N_5886,N_5486,N_5577);
or U5887 (N_5887,N_5554,N_5401);
and U5888 (N_5888,N_5329,N_5433);
nor U5889 (N_5889,N_5246,N_5493);
nor U5890 (N_5890,N_5494,N_5310);
and U5891 (N_5891,N_5446,N_5300);
nand U5892 (N_5892,N_5434,N_5269);
nand U5893 (N_5893,N_5452,N_5295);
xnor U5894 (N_5894,N_5512,N_5514);
nand U5895 (N_5895,N_5565,N_5523);
or U5896 (N_5896,N_5341,N_5266);
xor U5897 (N_5897,N_5514,N_5483);
and U5898 (N_5898,N_5297,N_5571);
nand U5899 (N_5899,N_5582,N_5289);
or U5900 (N_5900,N_5221,N_5494);
nand U5901 (N_5901,N_5481,N_5526);
xnor U5902 (N_5902,N_5202,N_5383);
or U5903 (N_5903,N_5211,N_5409);
nor U5904 (N_5904,N_5385,N_5429);
and U5905 (N_5905,N_5234,N_5490);
and U5906 (N_5906,N_5364,N_5437);
xnor U5907 (N_5907,N_5464,N_5473);
xnor U5908 (N_5908,N_5334,N_5564);
nand U5909 (N_5909,N_5240,N_5450);
and U5910 (N_5910,N_5344,N_5549);
or U5911 (N_5911,N_5256,N_5338);
or U5912 (N_5912,N_5413,N_5393);
and U5913 (N_5913,N_5470,N_5586);
nand U5914 (N_5914,N_5277,N_5426);
nor U5915 (N_5915,N_5242,N_5447);
and U5916 (N_5916,N_5273,N_5572);
xnor U5917 (N_5917,N_5344,N_5496);
or U5918 (N_5918,N_5251,N_5430);
nor U5919 (N_5919,N_5380,N_5431);
nand U5920 (N_5920,N_5392,N_5422);
nand U5921 (N_5921,N_5260,N_5401);
nand U5922 (N_5922,N_5507,N_5492);
and U5923 (N_5923,N_5223,N_5449);
xor U5924 (N_5924,N_5430,N_5591);
or U5925 (N_5925,N_5278,N_5519);
nand U5926 (N_5926,N_5494,N_5235);
xnor U5927 (N_5927,N_5482,N_5478);
xor U5928 (N_5928,N_5215,N_5431);
or U5929 (N_5929,N_5481,N_5395);
and U5930 (N_5930,N_5321,N_5328);
or U5931 (N_5931,N_5562,N_5464);
or U5932 (N_5932,N_5423,N_5459);
nor U5933 (N_5933,N_5467,N_5359);
or U5934 (N_5934,N_5428,N_5593);
xnor U5935 (N_5935,N_5543,N_5513);
nor U5936 (N_5936,N_5243,N_5218);
nand U5937 (N_5937,N_5295,N_5522);
or U5938 (N_5938,N_5335,N_5299);
or U5939 (N_5939,N_5482,N_5455);
and U5940 (N_5940,N_5458,N_5236);
or U5941 (N_5941,N_5376,N_5491);
and U5942 (N_5942,N_5367,N_5207);
or U5943 (N_5943,N_5276,N_5260);
nor U5944 (N_5944,N_5529,N_5563);
nand U5945 (N_5945,N_5444,N_5574);
and U5946 (N_5946,N_5440,N_5584);
nor U5947 (N_5947,N_5490,N_5397);
and U5948 (N_5948,N_5266,N_5449);
xor U5949 (N_5949,N_5489,N_5497);
or U5950 (N_5950,N_5433,N_5216);
or U5951 (N_5951,N_5559,N_5435);
xor U5952 (N_5952,N_5539,N_5252);
nor U5953 (N_5953,N_5432,N_5501);
xor U5954 (N_5954,N_5310,N_5400);
or U5955 (N_5955,N_5406,N_5366);
nand U5956 (N_5956,N_5210,N_5490);
or U5957 (N_5957,N_5581,N_5407);
xor U5958 (N_5958,N_5527,N_5483);
nor U5959 (N_5959,N_5220,N_5222);
and U5960 (N_5960,N_5504,N_5451);
xnor U5961 (N_5961,N_5544,N_5335);
and U5962 (N_5962,N_5526,N_5479);
and U5963 (N_5963,N_5225,N_5333);
xnor U5964 (N_5964,N_5267,N_5232);
or U5965 (N_5965,N_5387,N_5234);
nand U5966 (N_5966,N_5586,N_5424);
or U5967 (N_5967,N_5415,N_5211);
nor U5968 (N_5968,N_5593,N_5576);
xnor U5969 (N_5969,N_5316,N_5416);
and U5970 (N_5970,N_5463,N_5367);
nand U5971 (N_5971,N_5326,N_5392);
xnor U5972 (N_5972,N_5209,N_5524);
and U5973 (N_5973,N_5328,N_5547);
xor U5974 (N_5974,N_5568,N_5244);
nor U5975 (N_5975,N_5400,N_5402);
nor U5976 (N_5976,N_5545,N_5267);
and U5977 (N_5977,N_5595,N_5332);
and U5978 (N_5978,N_5202,N_5478);
nor U5979 (N_5979,N_5396,N_5541);
xor U5980 (N_5980,N_5576,N_5523);
nand U5981 (N_5981,N_5568,N_5300);
or U5982 (N_5982,N_5472,N_5230);
nor U5983 (N_5983,N_5538,N_5311);
nand U5984 (N_5984,N_5505,N_5354);
xnor U5985 (N_5985,N_5381,N_5493);
nand U5986 (N_5986,N_5592,N_5499);
nor U5987 (N_5987,N_5440,N_5492);
xor U5988 (N_5988,N_5265,N_5238);
and U5989 (N_5989,N_5270,N_5460);
xor U5990 (N_5990,N_5582,N_5499);
and U5991 (N_5991,N_5346,N_5553);
nand U5992 (N_5992,N_5569,N_5438);
xor U5993 (N_5993,N_5449,N_5376);
xor U5994 (N_5994,N_5222,N_5305);
or U5995 (N_5995,N_5502,N_5587);
nand U5996 (N_5996,N_5577,N_5315);
and U5997 (N_5997,N_5510,N_5433);
nor U5998 (N_5998,N_5553,N_5219);
xor U5999 (N_5999,N_5536,N_5291);
nor U6000 (N_6000,N_5712,N_5785);
or U6001 (N_6001,N_5704,N_5972);
nand U6002 (N_6002,N_5695,N_5786);
and U6003 (N_6003,N_5825,N_5870);
and U6004 (N_6004,N_5781,N_5846);
or U6005 (N_6005,N_5634,N_5606);
or U6006 (N_6006,N_5741,N_5642);
or U6007 (N_6007,N_5663,N_5819);
or U6008 (N_6008,N_5960,N_5768);
xnor U6009 (N_6009,N_5985,N_5787);
nor U6010 (N_6010,N_5766,N_5650);
nor U6011 (N_6011,N_5660,N_5603);
nor U6012 (N_6012,N_5818,N_5667);
nor U6013 (N_6013,N_5969,N_5738);
and U6014 (N_6014,N_5607,N_5792);
xor U6015 (N_6015,N_5814,N_5841);
nand U6016 (N_6016,N_5821,N_5622);
and U6017 (N_6017,N_5611,N_5823);
and U6018 (N_6018,N_5891,N_5955);
nand U6019 (N_6019,N_5772,N_5793);
xnor U6020 (N_6020,N_5703,N_5850);
or U6021 (N_6021,N_5829,N_5817);
xor U6022 (N_6022,N_5859,N_5919);
and U6023 (N_6023,N_5689,N_5815);
nand U6024 (N_6024,N_5938,N_5945);
xnor U6025 (N_6025,N_5675,N_5615);
and U6026 (N_6026,N_5926,N_5849);
xnor U6027 (N_6027,N_5964,N_5636);
xnor U6028 (N_6028,N_5681,N_5726);
or U6029 (N_6029,N_5759,N_5720);
nand U6030 (N_6030,N_5897,N_5933);
nor U6031 (N_6031,N_5764,N_5628);
nor U6032 (N_6032,N_5807,N_5736);
nor U6033 (N_6033,N_5635,N_5899);
and U6034 (N_6034,N_5629,N_5837);
nand U6035 (N_6035,N_5905,N_5674);
nand U6036 (N_6036,N_5789,N_5929);
nor U6037 (N_6037,N_5924,N_5653);
nor U6038 (N_6038,N_5991,N_5902);
nand U6039 (N_6039,N_5760,N_5932);
nor U6040 (N_6040,N_5980,N_5946);
nand U6041 (N_6041,N_5649,N_5655);
nor U6042 (N_6042,N_5942,N_5680);
nor U6043 (N_6043,N_5769,N_5887);
and U6044 (N_6044,N_5647,N_5844);
xnor U6045 (N_6045,N_5971,N_5696);
and U6046 (N_6046,N_5913,N_5914);
and U6047 (N_6047,N_5739,N_5728);
nor U6048 (N_6048,N_5927,N_5996);
or U6049 (N_6049,N_5828,N_5882);
xnor U6050 (N_6050,N_5612,N_5697);
nand U6051 (N_6051,N_5659,N_5824);
and U6052 (N_6052,N_5874,N_5725);
or U6053 (N_6053,N_5722,N_5701);
or U6054 (N_6054,N_5977,N_5868);
nand U6055 (N_6055,N_5613,N_5808);
nor U6056 (N_6056,N_5630,N_5620);
xnor U6057 (N_6057,N_5830,N_5707);
nor U6058 (N_6058,N_5752,N_5956);
nand U6059 (N_6059,N_5958,N_5835);
nor U6060 (N_6060,N_5831,N_5621);
nor U6061 (N_6061,N_5867,N_5862);
or U6062 (N_6062,N_5788,N_5627);
and U6063 (N_6063,N_5918,N_5940);
and U6064 (N_6064,N_5753,N_5638);
and U6065 (N_6065,N_5967,N_5797);
nand U6066 (N_6066,N_5686,N_5845);
and U6067 (N_6067,N_5757,N_5842);
nand U6068 (N_6068,N_5840,N_5664);
or U6069 (N_6069,N_5883,N_5966);
or U6070 (N_6070,N_5911,N_5648);
and U6071 (N_6071,N_5915,N_5806);
nor U6072 (N_6072,N_5656,N_5672);
xnor U6073 (N_6073,N_5602,N_5671);
nand U6074 (N_6074,N_5761,N_5652);
and U6075 (N_6075,N_5799,N_5685);
and U6076 (N_6076,N_5605,N_5993);
and U6077 (N_6077,N_5646,N_5921);
and U6078 (N_6078,N_5639,N_5865);
or U6079 (N_6079,N_5857,N_5645);
and U6080 (N_6080,N_5771,N_5986);
xnor U6081 (N_6081,N_5812,N_5898);
or U6082 (N_6082,N_5715,N_5763);
or U6083 (N_6083,N_5978,N_5893);
nand U6084 (N_6084,N_5661,N_5767);
and U6085 (N_6085,N_5983,N_5988);
nor U6086 (N_6086,N_5907,N_5925);
or U6087 (N_6087,N_5890,N_5894);
nor U6088 (N_6088,N_5952,N_5953);
nand U6089 (N_6089,N_5944,N_5827);
nand U6090 (N_6090,N_5832,N_5801);
xor U6091 (N_6091,N_5614,N_5719);
nor U6092 (N_6092,N_5608,N_5724);
xnor U6093 (N_6093,N_5854,N_5903);
nor U6094 (N_6094,N_5856,N_5888);
xor U6095 (N_6095,N_5884,N_5886);
or U6096 (N_6096,N_5916,N_5755);
or U6097 (N_6097,N_5651,N_5745);
nand U6098 (N_6098,N_5692,N_5880);
or U6099 (N_6099,N_5843,N_5976);
and U6100 (N_6100,N_5970,N_5709);
or U6101 (N_6101,N_5737,N_5896);
xnor U6102 (N_6102,N_5676,N_5705);
nand U6103 (N_6103,N_5826,N_5904);
and U6104 (N_6104,N_5878,N_5873);
nand U6105 (N_6105,N_5943,N_5791);
xnor U6106 (N_6106,N_5750,N_5941);
and U6107 (N_6107,N_5864,N_5858);
nor U6108 (N_6108,N_5816,N_5780);
nand U6109 (N_6109,N_5910,N_5776);
nor U6110 (N_6110,N_5892,N_5782);
nand U6111 (N_6111,N_5775,N_5637);
xnor U6112 (N_6112,N_5917,N_5673);
nor U6113 (N_6113,N_5730,N_5889);
or U6114 (N_6114,N_5810,N_5798);
and U6115 (N_6115,N_5901,N_5935);
nor U6116 (N_6116,N_5802,N_5982);
and U6117 (N_6117,N_5743,N_5803);
nor U6118 (N_6118,N_5618,N_5997);
and U6119 (N_6119,N_5879,N_5694);
and U6120 (N_6120,N_5625,N_5770);
xor U6121 (N_6121,N_5633,N_5989);
or U6122 (N_6122,N_5654,N_5968);
and U6123 (N_6123,N_5965,N_5714);
nor U6124 (N_6124,N_5912,N_5658);
or U6125 (N_6125,N_5794,N_5700);
nand U6126 (N_6126,N_5934,N_5687);
nor U6127 (N_6127,N_5833,N_5979);
nor U6128 (N_6128,N_5740,N_5616);
nand U6129 (N_6129,N_5800,N_5895);
nand U6130 (N_6130,N_5747,N_5702);
nand U6131 (N_6131,N_5626,N_5847);
xnor U6132 (N_6132,N_5604,N_5721);
nor U6133 (N_6133,N_5682,N_5951);
and U6134 (N_6134,N_5669,N_5711);
and U6135 (N_6135,N_5959,N_5718);
and U6136 (N_6136,N_5754,N_5640);
or U6137 (N_6137,N_5733,N_5632);
nand U6138 (N_6138,N_5691,N_5838);
nor U6139 (N_6139,N_5872,N_5954);
and U6140 (N_6140,N_5729,N_5662);
nor U6141 (N_6141,N_5748,N_5973);
nor U6142 (N_6142,N_5601,N_5665);
nor U6143 (N_6143,N_5949,N_5852);
xnor U6144 (N_6144,N_5804,N_5744);
or U6145 (N_6145,N_5688,N_5937);
and U6146 (N_6146,N_5751,N_5906);
and U6147 (N_6147,N_5778,N_5994);
or U6148 (N_6148,N_5641,N_5666);
nand U6149 (N_6149,N_5939,N_5683);
and U6150 (N_6150,N_5670,N_5813);
nand U6151 (N_6151,N_5936,N_5773);
and U6152 (N_6152,N_5962,N_5848);
and U6153 (N_6153,N_5657,N_5875);
and U6154 (N_6154,N_5928,N_5995);
or U6155 (N_6155,N_5668,N_5610);
xnor U6156 (N_6156,N_5922,N_5836);
or U6157 (N_6157,N_5866,N_5909);
and U6158 (N_6158,N_5617,N_5758);
nor U6159 (N_6159,N_5619,N_5795);
xor U6160 (N_6160,N_5881,N_5713);
nor U6161 (N_6161,N_5699,N_5885);
nor U6162 (N_6162,N_5623,N_5974);
nand U6163 (N_6163,N_5990,N_5999);
or U6164 (N_6164,N_5853,N_5877);
nor U6165 (N_6165,N_5742,N_5624);
nor U6166 (N_6166,N_5805,N_5957);
nor U6167 (N_6167,N_5600,N_5930);
nor U6168 (N_6168,N_5834,N_5947);
xnor U6169 (N_6169,N_5631,N_5790);
nor U6170 (N_6170,N_5809,N_5820);
nand U6171 (N_6171,N_5679,N_5677);
or U6172 (N_6172,N_5609,N_5734);
xor U6173 (N_6173,N_5987,N_5746);
and U6174 (N_6174,N_5861,N_5710);
and U6175 (N_6175,N_5860,N_5950);
xnor U6176 (N_6176,N_5811,N_5863);
xnor U6177 (N_6177,N_5735,N_5920);
and U6178 (N_6178,N_5908,N_5644);
nor U6179 (N_6179,N_5871,N_5774);
nand U6180 (N_6180,N_5869,N_5756);
xnor U6181 (N_6181,N_5693,N_5975);
or U6182 (N_6182,N_5855,N_5717);
nand U6183 (N_6183,N_5762,N_5732);
or U6184 (N_6184,N_5783,N_5784);
nand U6185 (N_6185,N_5777,N_5984);
xnor U6186 (N_6186,N_5749,N_5765);
nor U6187 (N_6187,N_5839,N_5981);
or U6188 (N_6188,N_5716,N_5727);
nor U6189 (N_6189,N_5684,N_5923);
nand U6190 (N_6190,N_5822,N_5690);
nor U6191 (N_6191,N_5900,N_5643);
or U6192 (N_6192,N_5931,N_5706);
nor U6193 (N_6193,N_5678,N_5708);
xnor U6194 (N_6194,N_5779,N_5851);
nor U6195 (N_6195,N_5961,N_5731);
nand U6196 (N_6196,N_5698,N_5948);
or U6197 (N_6197,N_5796,N_5876);
or U6198 (N_6198,N_5992,N_5998);
xor U6199 (N_6199,N_5963,N_5723);
nand U6200 (N_6200,N_5964,N_5771);
xor U6201 (N_6201,N_5980,N_5856);
and U6202 (N_6202,N_5954,N_5692);
and U6203 (N_6203,N_5652,N_5810);
nand U6204 (N_6204,N_5720,N_5908);
nand U6205 (N_6205,N_5923,N_5928);
or U6206 (N_6206,N_5750,N_5984);
nand U6207 (N_6207,N_5626,N_5963);
xor U6208 (N_6208,N_5971,N_5804);
nor U6209 (N_6209,N_5982,N_5668);
and U6210 (N_6210,N_5815,N_5900);
nor U6211 (N_6211,N_5660,N_5705);
and U6212 (N_6212,N_5919,N_5869);
or U6213 (N_6213,N_5916,N_5682);
xor U6214 (N_6214,N_5950,N_5839);
nand U6215 (N_6215,N_5738,N_5886);
nand U6216 (N_6216,N_5754,N_5992);
nand U6217 (N_6217,N_5826,N_5725);
xor U6218 (N_6218,N_5606,N_5930);
or U6219 (N_6219,N_5904,N_5828);
and U6220 (N_6220,N_5952,N_5633);
xor U6221 (N_6221,N_5992,N_5883);
and U6222 (N_6222,N_5684,N_5933);
nand U6223 (N_6223,N_5970,N_5999);
nor U6224 (N_6224,N_5863,N_5788);
nor U6225 (N_6225,N_5973,N_5999);
nand U6226 (N_6226,N_5840,N_5676);
and U6227 (N_6227,N_5646,N_5917);
or U6228 (N_6228,N_5868,N_5751);
and U6229 (N_6229,N_5648,N_5663);
and U6230 (N_6230,N_5632,N_5636);
and U6231 (N_6231,N_5705,N_5988);
xor U6232 (N_6232,N_5892,N_5678);
and U6233 (N_6233,N_5944,N_5960);
or U6234 (N_6234,N_5768,N_5644);
and U6235 (N_6235,N_5601,N_5681);
nand U6236 (N_6236,N_5999,N_5687);
and U6237 (N_6237,N_5791,N_5682);
xnor U6238 (N_6238,N_5813,N_5930);
or U6239 (N_6239,N_5762,N_5831);
nor U6240 (N_6240,N_5998,N_5652);
xor U6241 (N_6241,N_5902,N_5712);
nand U6242 (N_6242,N_5924,N_5762);
and U6243 (N_6243,N_5947,N_5832);
or U6244 (N_6244,N_5718,N_5934);
and U6245 (N_6245,N_5806,N_5903);
nand U6246 (N_6246,N_5723,N_5770);
or U6247 (N_6247,N_5842,N_5923);
and U6248 (N_6248,N_5989,N_5960);
or U6249 (N_6249,N_5735,N_5750);
and U6250 (N_6250,N_5660,N_5600);
and U6251 (N_6251,N_5673,N_5625);
nand U6252 (N_6252,N_5946,N_5904);
and U6253 (N_6253,N_5913,N_5938);
nand U6254 (N_6254,N_5896,N_5683);
or U6255 (N_6255,N_5644,N_5792);
nand U6256 (N_6256,N_5677,N_5616);
xnor U6257 (N_6257,N_5601,N_5815);
and U6258 (N_6258,N_5989,N_5858);
xor U6259 (N_6259,N_5816,N_5772);
nor U6260 (N_6260,N_5781,N_5654);
and U6261 (N_6261,N_5912,N_5762);
and U6262 (N_6262,N_5649,N_5630);
nand U6263 (N_6263,N_5971,N_5699);
and U6264 (N_6264,N_5617,N_5837);
nor U6265 (N_6265,N_5618,N_5945);
nor U6266 (N_6266,N_5708,N_5627);
and U6267 (N_6267,N_5764,N_5617);
nand U6268 (N_6268,N_5921,N_5831);
xor U6269 (N_6269,N_5804,N_5803);
and U6270 (N_6270,N_5673,N_5620);
or U6271 (N_6271,N_5993,N_5639);
and U6272 (N_6272,N_5962,N_5934);
and U6273 (N_6273,N_5720,N_5816);
nand U6274 (N_6274,N_5636,N_5789);
xor U6275 (N_6275,N_5766,N_5891);
nor U6276 (N_6276,N_5761,N_5819);
or U6277 (N_6277,N_5626,N_5744);
and U6278 (N_6278,N_5959,N_5603);
and U6279 (N_6279,N_5926,N_5831);
and U6280 (N_6280,N_5609,N_5899);
and U6281 (N_6281,N_5732,N_5824);
or U6282 (N_6282,N_5928,N_5745);
and U6283 (N_6283,N_5834,N_5607);
xnor U6284 (N_6284,N_5970,N_5720);
nand U6285 (N_6285,N_5940,N_5899);
xor U6286 (N_6286,N_5625,N_5921);
nor U6287 (N_6287,N_5875,N_5957);
xor U6288 (N_6288,N_5778,N_5985);
and U6289 (N_6289,N_5680,N_5794);
xor U6290 (N_6290,N_5787,N_5864);
nand U6291 (N_6291,N_5922,N_5603);
and U6292 (N_6292,N_5630,N_5713);
xor U6293 (N_6293,N_5788,N_5743);
or U6294 (N_6294,N_5916,N_5934);
nand U6295 (N_6295,N_5905,N_5887);
nand U6296 (N_6296,N_5949,N_5773);
xor U6297 (N_6297,N_5732,N_5785);
or U6298 (N_6298,N_5876,N_5621);
nand U6299 (N_6299,N_5931,N_5918);
or U6300 (N_6300,N_5731,N_5626);
xor U6301 (N_6301,N_5761,N_5681);
xnor U6302 (N_6302,N_5636,N_5962);
and U6303 (N_6303,N_5639,N_5656);
or U6304 (N_6304,N_5630,N_5856);
and U6305 (N_6305,N_5685,N_5962);
nand U6306 (N_6306,N_5693,N_5996);
or U6307 (N_6307,N_5835,N_5714);
xor U6308 (N_6308,N_5801,N_5739);
nor U6309 (N_6309,N_5960,N_5761);
nand U6310 (N_6310,N_5785,N_5998);
nor U6311 (N_6311,N_5600,N_5780);
nand U6312 (N_6312,N_5912,N_5933);
nor U6313 (N_6313,N_5927,N_5770);
nor U6314 (N_6314,N_5729,N_5862);
and U6315 (N_6315,N_5824,N_5977);
and U6316 (N_6316,N_5864,N_5733);
nor U6317 (N_6317,N_5925,N_5956);
nor U6318 (N_6318,N_5819,N_5654);
xor U6319 (N_6319,N_5852,N_5837);
nand U6320 (N_6320,N_5667,N_5905);
or U6321 (N_6321,N_5671,N_5768);
nand U6322 (N_6322,N_5813,N_5651);
nor U6323 (N_6323,N_5641,N_5801);
nand U6324 (N_6324,N_5760,N_5731);
or U6325 (N_6325,N_5754,N_5906);
xor U6326 (N_6326,N_5602,N_5682);
nor U6327 (N_6327,N_5950,N_5739);
nor U6328 (N_6328,N_5795,N_5629);
xor U6329 (N_6329,N_5931,N_5615);
nand U6330 (N_6330,N_5840,N_5857);
nand U6331 (N_6331,N_5824,N_5740);
nand U6332 (N_6332,N_5793,N_5713);
nor U6333 (N_6333,N_5904,N_5701);
xor U6334 (N_6334,N_5720,N_5709);
and U6335 (N_6335,N_5617,N_5621);
and U6336 (N_6336,N_5961,N_5729);
or U6337 (N_6337,N_5626,N_5789);
xnor U6338 (N_6338,N_5755,N_5746);
and U6339 (N_6339,N_5937,N_5707);
nor U6340 (N_6340,N_5813,N_5765);
and U6341 (N_6341,N_5808,N_5615);
and U6342 (N_6342,N_5995,N_5641);
or U6343 (N_6343,N_5799,N_5732);
and U6344 (N_6344,N_5961,N_5822);
and U6345 (N_6345,N_5668,N_5609);
nand U6346 (N_6346,N_5721,N_5917);
or U6347 (N_6347,N_5706,N_5717);
xor U6348 (N_6348,N_5786,N_5720);
nand U6349 (N_6349,N_5850,N_5796);
and U6350 (N_6350,N_5906,N_5847);
nand U6351 (N_6351,N_5967,N_5811);
nand U6352 (N_6352,N_5623,N_5806);
xnor U6353 (N_6353,N_5631,N_5617);
nand U6354 (N_6354,N_5651,N_5689);
nand U6355 (N_6355,N_5862,N_5818);
or U6356 (N_6356,N_5749,N_5655);
nor U6357 (N_6357,N_5968,N_5923);
nor U6358 (N_6358,N_5767,N_5917);
or U6359 (N_6359,N_5919,N_5888);
nor U6360 (N_6360,N_5978,N_5648);
xor U6361 (N_6361,N_5660,N_5625);
or U6362 (N_6362,N_5949,N_5901);
and U6363 (N_6363,N_5767,N_5872);
nor U6364 (N_6364,N_5938,N_5677);
xor U6365 (N_6365,N_5633,N_5789);
xor U6366 (N_6366,N_5768,N_5937);
nor U6367 (N_6367,N_5777,N_5686);
nor U6368 (N_6368,N_5787,N_5602);
nor U6369 (N_6369,N_5676,N_5716);
or U6370 (N_6370,N_5715,N_5814);
nor U6371 (N_6371,N_5886,N_5726);
nand U6372 (N_6372,N_5942,N_5884);
or U6373 (N_6373,N_5628,N_5775);
or U6374 (N_6374,N_5848,N_5639);
xor U6375 (N_6375,N_5760,N_5624);
and U6376 (N_6376,N_5805,N_5729);
and U6377 (N_6377,N_5659,N_5661);
or U6378 (N_6378,N_5975,N_5946);
and U6379 (N_6379,N_5871,N_5697);
and U6380 (N_6380,N_5835,N_5653);
and U6381 (N_6381,N_5801,N_5970);
and U6382 (N_6382,N_5714,N_5855);
nand U6383 (N_6383,N_5626,N_5845);
nand U6384 (N_6384,N_5800,N_5883);
xnor U6385 (N_6385,N_5918,N_5620);
nor U6386 (N_6386,N_5747,N_5882);
nand U6387 (N_6387,N_5761,N_5779);
nand U6388 (N_6388,N_5927,N_5955);
xor U6389 (N_6389,N_5795,N_5955);
nor U6390 (N_6390,N_5787,N_5732);
or U6391 (N_6391,N_5786,N_5819);
nor U6392 (N_6392,N_5991,N_5663);
or U6393 (N_6393,N_5620,N_5978);
xnor U6394 (N_6394,N_5824,N_5940);
or U6395 (N_6395,N_5930,N_5862);
nand U6396 (N_6396,N_5947,N_5906);
or U6397 (N_6397,N_5845,N_5762);
nor U6398 (N_6398,N_5663,N_5688);
nand U6399 (N_6399,N_5782,N_5972);
nand U6400 (N_6400,N_6073,N_6253);
nand U6401 (N_6401,N_6258,N_6078);
or U6402 (N_6402,N_6291,N_6210);
or U6403 (N_6403,N_6230,N_6184);
xnor U6404 (N_6404,N_6372,N_6166);
or U6405 (N_6405,N_6333,N_6032);
or U6406 (N_6406,N_6099,N_6292);
xor U6407 (N_6407,N_6239,N_6397);
nor U6408 (N_6408,N_6118,N_6286);
nor U6409 (N_6409,N_6116,N_6182);
xor U6410 (N_6410,N_6074,N_6080);
nand U6411 (N_6411,N_6389,N_6186);
and U6412 (N_6412,N_6146,N_6161);
nor U6413 (N_6413,N_6367,N_6029);
nor U6414 (N_6414,N_6172,N_6115);
and U6415 (N_6415,N_6297,N_6361);
xor U6416 (N_6416,N_6298,N_6196);
nor U6417 (N_6417,N_6380,N_6165);
nor U6418 (N_6418,N_6202,N_6315);
nand U6419 (N_6419,N_6133,N_6224);
nand U6420 (N_6420,N_6132,N_6143);
or U6421 (N_6421,N_6303,N_6157);
nor U6422 (N_6422,N_6122,N_6136);
or U6423 (N_6423,N_6378,N_6283);
xor U6424 (N_6424,N_6047,N_6265);
and U6425 (N_6425,N_6288,N_6294);
or U6426 (N_6426,N_6362,N_6038);
or U6427 (N_6427,N_6162,N_6335);
or U6428 (N_6428,N_6042,N_6190);
xnor U6429 (N_6429,N_6175,N_6026);
nand U6430 (N_6430,N_6383,N_6109);
xnor U6431 (N_6431,N_6075,N_6130);
xor U6432 (N_6432,N_6251,N_6226);
nor U6433 (N_6433,N_6147,N_6189);
nand U6434 (N_6434,N_6227,N_6219);
and U6435 (N_6435,N_6002,N_6369);
nor U6436 (N_6436,N_6097,N_6174);
or U6437 (N_6437,N_6326,N_6151);
nor U6438 (N_6438,N_6101,N_6120);
nor U6439 (N_6439,N_6160,N_6168);
nor U6440 (N_6440,N_6246,N_6373);
and U6441 (N_6441,N_6039,N_6338);
nor U6442 (N_6442,N_6142,N_6170);
or U6443 (N_6443,N_6067,N_6191);
or U6444 (N_6444,N_6276,N_6313);
or U6445 (N_6445,N_6134,N_6054);
nand U6446 (N_6446,N_6332,N_6187);
nor U6447 (N_6447,N_6200,N_6035);
nor U6448 (N_6448,N_6153,N_6365);
and U6449 (N_6449,N_6155,N_6236);
nand U6450 (N_6450,N_6261,N_6302);
and U6451 (N_6451,N_6144,N_6106);
xnor U6452 (N_6452,N_6030,N_6152);
nand U6453 (N_6453,N_6237,N_6388);
xnor U6454 (N_6454,N_6204,N_6090);
or U6455 (N_6455,N_6164,N_6371);
or U6456 (N_6456,N_6211,N_6242);
nand U6457 (N_6457,N_6323,N_6346);
nor U6458 (N_6458,N_6308,N_6129);
and U6459 (N_6459,N_6064,N_6299);
and U6460 (N_6460,N_6334,N_6125);
nor U6461 (N_6461,N_6353,N_6275);
nand U6462 (N_6462,N_6018,N_6310);
or U6463 (N_6463,N_6138,N_6317);
nand U6464 (N_6464,N_6354,N_6216);
xnor U6465 (N_6465,N_6025,N_6231);
nand U6466 (N_6466,N_6278,N_6086);
or U6467 (N_6467,N_6398,N_6010);
and U6468 (N_6468,N_6069,N_6094);
and U6469 (N_6469,N_6046,N_6245);
and U6470 (N_6470,N_6004,N_6104);
or U6471 (N_6471,N_6045,N_6267);
xor U6472 (N_6472,N_6240,N_6021);
xnor U6473 (N_6473,N_6093,N_6033);
and U6474 (N_6474,N_6287,N_6041);
or U6475 (N_6475,N_6169,N_6177);
nand U6476 (N_6476,N_6014,N_6306);
nor U6477 (N_6477,N_6314,N_6357);
nor U6478 (N_6478,N_6220,N_6135);
nand U6479 (N_6479,N_6229,N_6259);
or U6480 (N_6480,N_6309,N_6344);
and U6481 (N_6481,N_6111,N_6096);
nand U6482 (N_6482,N_6206,N_6049);
and U6483 (N_6483,N_6279,N_6195);
or U6484 (N_6484,N_6301,N_6312);
nor U6485 (N_6485,N_6053,N_6063);
and U6486 (N_6486,N_6062,N_6137);
or U6487 (N_6487,N_6040,N_6325);
xnor U6488 (N_6488,N_6359,N_6342);
or U6489 (N_6489,N_6052,N_6149);
and U6490 (N_6490,N_6396,N_6254);
or U6491 (N_6491,N_6262,N_6375);
xor U6492 (N_6492,N_6000,N_6320);
nor U6493 (N_6493,N_6188,N_6065);
xnor U6494 (N_6494,N_6159,N_6167);
nor U6495 (N_6495,N_6023,N_6390);
xor U6496 (N_6496,N_6296,N_6207);
and U6497 (N_6497,N_6154,N_6260);
nand U6498 (N_6498,N_6285,N_6201);
nor U6499 (N_6499,N_6368,N_6011);
or U6500 (N_6500,N_6257,N_6197);
or U6501 (N_6501,N_6095,N_6060);
nor U6502 (N_6502,N_6392,N_6381);
and U6503 (N_6503,N_6300,N_6247);
or U6504 (N_6504,N_6061,N_6356);
xor U6505 (N_6505,N_6171,N_6072);
or U6506 (N_6506,N_6056,N_6268);
xor U6507 (N_6507,N_6345,N_6307);
xor U6508 (N_6508,N_6100,N_6319);
xnor U6509 (N_6509,N_6222,N_6295);
or U6510 (N_6510,N_6327,N_6007);
nand U6511 (N_6511,N_6214,N_6077);
nor U6512 (N_6512,N_6213,N_6178);
nand U6513 (N_6513,N_6238,N_6181);
nor U6514 (N_6514,N_6043,N_6385);
nor U6515 (N_6515,N_6360,N_6048);
nor U6516 (N_6516,N_6193,N_6079);
nor U6517 (N_6517,N_6016,N_6330);
nand U6518 (N_6518,N_6103,N_6350);
xnor U6519 (N_6519,N_6290,N_6318);
xor U6520 (N_6520,N_6255,N_6266);
or U6521 (N_6521,N_6244,N_6006);
nor U6522 (N_6522,N_6374,N_6399);
or U6523 (N_6523,N_6321,N_6176);
nor U6524 (N_6524,N_6013,N_6036);
nand U6525 (N_6525,N_6092,N_6119);
nor U6526 (N_6526,N_6156,N_6008);
nor U6527 (N_6527,N_6059,N_6347);
or U6528 (N_6528,N_6233,N_6185);
nand U6529 (N_6529,N_6228,N_6234);
nor U6530 (N_6530,N_6068,N_6370);
and U6531 (N_6531,N_6249,N_6324);
or U6532 (N_6532,N_6284,N_6012);
nor U6533 (N_6533,N_6293,N_6387);
or U6534 (N_6534,N_6091,N_6089);
nor U6535 (N_6535,N_6180,N_6280);
nor U6536 (N_6536,N_6364,N_6150);
nand U6537 (N_6537,N_6085,N_6179);
xnor U6538 (N_6538,N_6336,N_6393);
nor U6539 (N_6539,N_6084,N_6055);
nand U6540 (N_6540,N_6376,N_6215);
nor U6541 (N_6541,N_6117,N_6001);
or U6542 (N_6542,N_6145,N_6027);
or U6543 (N_6543,N_6256,N_6140);
and U6544 (N_6544,N_6395,N_6348);
and U6545 (N_6545,N_6102,N_6087);
nand U6546 (N_6546,N_6250,N_6269);
and U6547 (N_6547,N_6289,N_6391);
and U6548 (N_6548,N_6329,N_6281);
nand U6549 (N_6549,N_6082,N_6126);
and U6550 (N_6550,N_6105,N_6127);
nor U6551 (N_6551,N_6355,N_6304);
and U6552 (N_6552,N_6305,N_6208);
or U6553 (N_6553,N_6225,N_6339);
nand U6554 (N_6554,N_6358,N_6163);
and U6555 (N_6555,N_6384,N_6199);
nand U6556 (N_6556,N_6366,N_6217);
xor U6557 (N_6557,N_6070,N_6205);
nor U6558 (N_6558,N_6352,N_6194);
and U6559 (N_6559,N_6098,N_6066);
and U6560 (N_6560,N_6209,N_6263);
nand U6561 (N_6561,N_6377,N_6110);
or U6562 (N_6562,N_6218,N_6277);
xor U6563 (N_6563,N_6271,N_6340);
nand U6564 (N_6564,N_6003,N_6337);
nor U6565 (N_6565,N_6316,N_6131);
nor U6566 (N_6566,N_6341,N_6235);
and U6567 (N_6567,N_6024,N_6343);
xnor U6568 (N_6568,N_6273,N_6071);
and U6569 (N_6569,N_6020,N_6123);
nand U6570 (N_6570,N_6113,N_6124);
or U6571 (N_6571,N_6121,N_6274);
nand U6572 (N_6572,N_6028,N_6044);
nand U6573 (N_6573,N_6272,N_6221);
nor U6574 (N_6574,N_6248,N_6241);
nand U6575 (N_6575,N_6051,N_6019);
nand U6576 (N_6576,N_6386,N_6252);
xnor U6577 (N_6577,N_6232,N_6005);
nand U6578 (N_6578,N_6076,N_6264);
or U6579 (N_6579,N_6282,N_6328);
xnor U6580 (N_6580,N_6107,N_6139);
nand U6581 (N_6581,N_6363,N_6088);
and U6582 (N_6582,N_6322,N_6158);
nor U6583 (N_6583,N_6108,N_6243);
and U6584 (N_6584,N_6349,N_6081);
xor U6585 (N_6585,N_6331,N_6112);
or U6586 (N_6586,N_6009,N_6141);
and U6587 (N_6587,N_6148,N_6017);
or U6588 (N_6588,N_6034,N_6031);
nor U6589 (N_6589,N_6128,N_6015);
nor U6590 (N_6590,N_6050,N_6083);
xor U6591 (N_6591,N_6311,N_6022);
nand U6592 (N_6592,N_6212,N_6058);
nand U6593 (N_6593,N_6203,N_6382);
nor U6594 (N_6594,N_6057,N_6037);
xor U6595 (N_6595,N_6183,N_6351);
or U6596 (N_6596,N_6379,N_6270);
xor U6597 (N_6597,N_6114,N_6394);
and U6598 (N_6598,N_6192,N_6223);
or U6599 (N_6599,N_6198,N_6173);
or U6600 (N_6600,N_6140,N_6313);
xor U6601 (N_6601,N_6204,N_6305);
nand U6602 (N_6602,N_6291,N_6217);
xnor U6603 (N_6603,N_6193,N_6177);
and U6604 (N_6604,N_6071,N_6216);
nand U6605 (N_6605,N_6261,N_6247);
nand U6606 (N_6606,N_6155,N_6069);
or U6607 (N_6607,N_6018,N_6139);
nor U6608 (N_6608,N_6125,N_6194);
or U6609 (N_6609,N_6170,N_6069);
or U6610 (N_6610,N_6286,N_6214);
nor U6611 (N_6611,N_6210,N_6052);
and U6612 (N_6612,N_6240,N_6195);
nand U6613 (N_6613,N_6293,N_6332);
or U6614 (N_6614,N_6365,N_6114);
or U6615 (N_6615,N_6252,N_6378);
or U6616 (N_6616,N_6154,N_6232);
xnor U6617 (N_6617,N_6203,N_6061);
nor U6618 (N_6618,N_6376,N_6107);
and U6619 (N_6619,N_6329,N_6316);
nand U6620 (N_6620,N_6328,N_6323);
nand U6621 (N_6621,N_6004,N_6056);
xnor U6622 (N_6622,N_6255,N_6189);
nand U6623 (N_6623,N_6147,N_6331);
nand U6624 (N_6624,N_6359,N_6029);
nand U6625 (N_6625,N_6149,N_6276);
or U6626 (N_6626,N_6283,N_6318);
and U6627 (N_6627,N_6382,N_6015);
or U6628 (N_6628,N_6386,N_6290);
nand U6629 (N_6629,N_6332,N_6063);
nor U6630 (N_6630,N_6368,N_6348);
nor U6631 (N_6631,N_6137,N_6036);
or U6632 (N_6632,N_6152,N_6370);
xnor U6633 (N_6633,N_6310,N_6238);
nand U6634 (N_6634,N_6214,N_6396);
or U6635 (N_6635,N_6336,N_6029);
nor U6636 (N_6636,N_6195,N_6140);
and U6637 (N_6637,N_6089,N_6386);
or U6638 (N_6638,N_6167,N_6203);
or U6639 (N_6639,N_6357,N_6300);
or U6640 (N_6640,N_6162,N_6079);
xor U6641 (N_6641,N_6356,N_6130);
or U6642 (N_6642,N_6016,N_6020);
nor U6643 (N_6643,N_6112,N_6240);
nor U6644 (N_6644,N_6041,N_6201);
or U6645 (N_6645,N_6356,N_6185);
nor U6646 (N_6646,N_6026,N_6225);
and U6647 (N_6647,N_6197,N_6252);
and U6648 (N_6648,N_6064,N_6250);
xnor U6649 (N_6649,N_6322,N_6044);
or U6650 (N_6650,N_6059,N_6106);
nor U6651 (N_6651,N_6227,N_6243);
nand U6652 (N_6652,N_6263,N_6102);
nand U6653 (N_6653,N_6023,N_6011);
nor U6654 (N_6654,N_6385,N_6137);
xor U6655 (N_6655,N_6017,N_6156);
nand U6656 (N_6656,N_6231,N_6353);
nand U6657 (N_6657,N_6014,N_6272);
and U6658 (N_6658,N_6049,N_6277);
and U6659 (N_6659,N_6146,N_6077);
nand U6660 (N_6660,N_6223,N_6379);
or U6661 (N_6661,N_6091,N_6014);
xor U6662 (N_6662,N_6252,N_6349);
xor U6663 (N_6663,N_6246,N_6011);
nor U6664 (N_6664,N_6284,N_6111);
xnor U6665 (N_6665,N_6248,N_6064);
nor U6666 (N_6666,N_6387,N_6273);
xnor U6667 (N_6667,N_6061,N_6035);
xnor U6668 (N_6668,N_6144,N_6185);
xnor U6669 (N_6669,N_6345,N_6358);
xnor U6670 (N_6670,N_6225,N_6147);
or U6671 (N_6671,N_6033,N_6192);
nor U6672 (N_6672,N_6333,N_6116);
nor U6673 (N_6673,N_6375,N_6108);
or U6674 (N_6674,N_6007,N_6102);
nor U6675 (N_6675,N_6266,N_6128);
xor U6676 (N_6676,N_6067,N_6105);
xnor U6677 (N_6677,N_6188,N_6165);
nand U6678 (N_6678,N_6040,N_6105);
and U6679 (N_6679,N_6281,N_6397);
or U6680 (N_6680,N_6077,N_6055);
and U6681 (N_6681,N_6260,N_6003);
nor U6682 (N_6682,N_6172,N_6149);
or U6683 (N_6683,N_6291,N_6303);
xnor U6684 (N_6684,N_6130,N_6094);
or U6685 (N_6685,N_6046,N_6167);
and U6686 (N_6686,N_6224,N_6064);
nor U6687 (N_6687,N_6228,N_6070);
and U6688 (N_6688,N_6041,N_6024);
and U6689 (N_6689,N_6292,N_6072);
nand U6690 (N_6690,N_6023,N_6092);
xor U6691 (N_6691,N_6335,N_6074);
or U6692 (N_6692,N_6231,N_6295);
and U6693 (N_6693,N_6397,N_6034);
xnor U6694 (N_6694,N_6111,N_6215);
nand U6695 (N_6695,N_6012,N_6142);
and U6696 (N_6696,N_6166,N_6004);
xor U6697 (N_6697,N_6297,N_6223);
xnor U6698 (N_6698,N_6209,N_6110);
and U6699 (N_6699,N_6220,N_6067);
or U6700 (N_6700,N_6384,N_6209);
and U6701 (N_6701,N_6188,N_6227);
or U6702 (N_6702,N_6340,N_6246);
xnor U6703 (N_6703,N_6125,N_6247);
nor U6704 (N_6704,N_6256,N_6388);
nor U6705 (N_6705,N_6159,N_6375);
nand U6706 (N_6706,N_6184,N_6339);
xnor U6707 (N_6707,N_6360,N_6195);
xor U6708 (N_6708,N_6188,N_6232);
nor U6709 (N_6709,N_6395,N_6205);
xor U6710 (N_6710,N_6300,N_6232);
and U6711 (N_6711,N_6331,N_6271);
xor U6712 (N_6712,N_6074,N_6165);
xnor U6713 (N_6713,N_6386,N_6095);
nor U6714 (N_6714,N_6136,N_6205);
nor U6715 (N_6715,N_6259,N_6349);
nand U6716 (N_6716,N_6282,N_6053);
xor U6717 (N_6717,N_6284,N_6218);
and U6718 (N_6718,N_6023,N_6106);
nor U6719 (N_6719,N_6202,N_6298);
nor U6720 (N_6720,N_6032,N_6008);
nor U6721 (N_6721,N_6004,N_6271);
nand U6722 (N_6722,N_6223,N_6258);
xnor U6723 (N_6723,N_6184,N_6164);
and U6724 (N_6724,N_6097,N_6080);
nand U6725 (N_6725,N_6373,N_6237);
xor U6726 (N_6726,N_6223,N_6308);
nor U6727 (N_6727,N_6223,N_6183);
nand U6728 (N_6728,N_6176,N_6155);
or U6729 (N_6729,N_6321,N_6122);
xor U6730 (N_6730,N_6050,N_6194);
nand U6731 (N_6731,N_6188,N_6051);
or U6732 (N_6732,N_6345,N_6063);
nand U6733 (N_6733,N_6259,N_6244);
nor U6734 (N_6734,N_6247,N_6096);
or U6735 (N_6735,N_6265,N_6213);
nor U6736 (N_6736,N_6264,N_6227);
nand U6737 (N_6737,N_6034,N_6315);
nor U6738 (N_6738,N_6031,N_6018);
or U6739 (N_6739,N_6044,N_6282);
nor U6740 (N_6740,N_6161,N_6268);
and U6741 (N_6741,N_6108,N_6011);
and U6742 (N_6742,N_6127,N_6092);
or U6743 (N_6743,N_6012,N_6038);
xor U6744 (N_6744,N_6350,N_6327);
nor U6745 (N_6745,N_6395,N_6065);
nand U6746 (N_6746,N_6032,N_6150);
or U6747 (N_6747,N_6337,N_6232);
xnor U6748 (N_6748,N_6118,N_6322);
nor U6749 (N_6749,N_6017,N_6177);
nor U6750 (N_6750,N_6088,N_6173);
nand U6751 (N_6751,N_6391,N_6116);
nand U6752 (N_6752,N_6336,N_6117);
nand U6753 (N_6753,N_6088,N_6319);
xnor U6754 (N_6754,N_6249,N_6101);
nand U6755 (N_6755,N_6284,N_6046);
nand U6756 (N_6756,N_6195,N_6131);
or U6757 (N_6757,N_6105,N_6367);
and U6758 (N_6758,N_6234,N_6316);
or U6759 (N_6759,N_6344,N_6188);
xor U6760 (N_6760,N_6382,N_6325);
or U6761 (N_6761,N_6258,N_6393);
and U6762 (N_6762,N_6074,N_6304);
xor U6763 (N_6763,N_6212,N_6340);
nand U6764 (N_6764,N_6089,N_6336);
or U6765 (N_6765,N_6245,N_6187);
and U6766 (N_6766,N_6135,N_6012);
and U6767 (N_6767,N_6245,N_6293);
or U6768 (N_6768,N_6272,N_6060);
and U6769 (N_6769,N_6278,N_6332);
nand U6770 (N_6770,N_6257,N_6244);
and U6771 (N_6771,N_6214,N_6074);
nor U6772 (N_6772,N_6289,N_6089);
nor U6773 (N_6773,N_6244,N_6192);
or U6774 (N_6774,N_6038,N_6087);
and U6775 (N_6775,N_6164,N_6055);
xor U6776 (N_6776,N_6270,N_6010);
nand U6777 (N_6777,N_6165,N_6066);
nand U6778 (N_6778,N_6196,N_6072);
or U6779 (N_6779,N_6331,N_6267);
and U6780 (N_6780,N_6201,N_6330);
nand U6781 (N_6781,N_6099,N_6355);
and U6782 (N_6782,N_6306,N_6349);
and U6783 (N_6783,N_6342,N_6239);
nor U6784 (N_6784,N_6176,N_6219);
or U6785 (N_6785,N_6339,N_6204);
xor U6786 (N_6786,N_6193,N_6242);
or U6787 (N_6787,N_6221,N_6079);
xnor U6788 (N_6788,N_6118,N_6166);
nand U6789 (N_6789,N_6286,N_6018);
nor U6790 (N_6790,N_6191,N_6018);
or U6791 (N_6791,N_6306,N_6105);
nor U6792 (N_6792,N_6398,N_6266);
and U6793 (N_6793,N_6251,N_6337);
xnor U6794 (N_6794,N_6057,N_6217);
xor U6795 (N_6795,N_6298,N_6157);
and U6796 (N_6796,N_6195,N_6254);
xor U6797 (N_6797,N_6104,N_6143);
or U6798 (N_6798,N_6264,N_6126);
and U6799 (N_6799,N_6218,N_6216);
xor U6800 (N_6800,N_6626,N_6417);
nand U6801 (N_6801,N_6554,N_6536);
xor U6802 (N_6802,N_6443,N_6753);
xnor U6803 (N_6803,N_6691,N_6513);
or U6804 (N_6804,N_6501,N_6579);
xnor U6805 (N_6805,N_6498,N_6438);
and U6806 (N_6806,N_6724,N_6707);
xor U6807 (N_6807,N_6401,N_6407);
xnor U6808 (N_6808,N_6439,N_6721);
xor U6809 (N_6809,N_6575,N_6675);
and U6810 (N_6810,N_6486,N_6733);
xnor U6811 (N_6811,N_6732,N_6740);
or U6812 (N_6812,N_6549,N_6709);
nand U6813 (N_6813,N_6465,N_6510);
xor U6814 (N_6814,N_6539,N_6754);
or U6815 (N_6815,N_6661,N_6516);
and U6816 (N_6816,N_6553,N_6734);
and U6817 (N_6817,N_6424,N_6455);
or U6818 (N_6818,N_6777,N_6674);
xnor U6819 (N_6819,N_6520,N_6503);
xnor U6820 (N_6820,N_6766,N_6795);
nand U6821 (N_6821,N_6568,N_6489);
and U6822 (N_6822,N_6507,N_6454);
and U6823 (N_6823,N_6610,N_6594);
xor U6824 (N_6824,N_6739,N_6676);
nand U6825 (N_6825,N_6637,N_6776);
xnor U6826 (N_6826,N_6402,N_6673);
or U6827 (N_6827,N_6615,N_6548);
xnor U6828 (N_6828,N_6569,N_6587);
or U6829 (N_6829,N_6490,N_6537);
xnor U6830 (N_6830,N_6680,N_6755);
xnor U6831 (N_6831,N_6614,N_6480);
xor U6832 (N_6832,N_6589,N_6749);
and U6833 (N_6833,N_6640,N_6412);
nand U6834 (N_6834,N_6664,N_6584);
and U6835 (N_6835,N_6727,N_6542);
or U6836 (N_6836,N_6530,N_6759);
or U6837 (N_6837,N_6440,N_6582);
or U6838 (N_6838,N_6572,N_6798);
nor U6839 (N_6839,N_6476,N_6748);
xnor U6840 (N_6840,N_6634,N_6599);
nor U6841 (N_6841,N_6606,N_6478);
and U6842 (N_6842,N_6552,N_6526);
xnor U6843 (N_6843,N_6598,N_6481);
or U6844 (N_6844,N_6566,N_6446);
and U6845 (N_6845,N_6469,N_6484);
or U6846 (N_6846,N_6604,N_6525);
nand U6847 (N_6847,N_6714,N_6595);
nor U6848 (N_6848,N_6585,N_6430);
or U6849 (N_6849,N_6411,N_6785);
or U6850 (N_6850,N_6467,N_6658);
or U6851 (N_6851,N_6767,N_6408);
xnor U6852 (N_6852,N_6656,N_6725);
xor U6853 (N_6853,N_6508,N_6699);
xor U6854 (N_6854,N_6462,N_6442);
or U6855 (N_6855,N_6414,N_6609);
xnor U6856 (N_6856,N_6563,N_6752);
nor U6857 (N_6857,N_6635,N_6485);
nor U6858 (N_6858,N_6743,N_6760);
or U6859 (N_6859,N_6715,N_6444);
nor U6860 (N_6860,N_6698,N_6405);
xor U6861 (N_6861,N_6791,N_6527);
nand U6862 (N_6862,N_6550,N_6722);
nand U6863 (N_6863,N_6729,N_6796);
xnor U6864 (N_6864,N_6705,N_6792);
xnor U6865 (N_6865,N_6421,N_6448);
and U6866 (N_6866,N_6670,N_6639);
xnor U6867 (N_6867,N_6689,N_6644);
nand U6868 (N_6868,N_6578,N_6735);
nor U6869 (N_6869,N_6617,N_6782);
or U6870 (N_6870,N_6746,N_6741);
or U6871 (N_6871,N_6681,N_6757);
nand U6872 (N_6872,N_6713,N_6780);
and U6873 (N_6873,N_6645,N_6535);
nor U6874 (N_6874,N_6738,N_6627);
xor U6875 (N_6875,N_6684,N_6437);
or U6876 (N_6876,N_6660,N_6493);
and U6877 (N_6877,N_6747,N_6488);
xor U6878 (N_6878,N_6601,N_6559);
nand U6879 (N_6879,N_6678,N_6758);
and U6880 (N_6880,N_6642,N_6499);
xor U6881 (N_6881,N_6630,N_6596);
and U6882 (N_6882,N_6477,N_6663);
or U6883 (N_6883,N_6558,N_6666);
and U6884 (N_6884,N_6400,N_6761);
nand U6885 (N_6885,N_6685,N_6571);
xnor U6886 (N_6886,N_6564,N_6768);
xnor U6887 (N_6887,N_6745,N_6471);
nor U6888 (N_6888,N_6463,N_6742);
nor U6889 (N_6889,N_6788,N_6551);
or U6890 (N_6890,N_6441,N_6461);
and U6891 (N_6891,N_6688,N_6410);
nand U6892 (N_6892,N_6718,N_6750);
nor U6893 (N_6893,N_6719,N_6545);
nand U6894 (N_6894,N_6413,N_6669);
or U6895 (N_6895,N_6631,N_6653);
nand U6896 (N_6896,N_6581,N_6435);
nand U6897 (N_6897,N_6693,N_6602);
nor U6898 (N_6898,N_6576,N_6771);
nand U6899 (N_6899,N_6641,N_6547);
or U6900 (N_6900,N_6638,N_6731);
xnor U6901 (N_6901,N_6473,N_6612);
and U6902 (N_6902,N_6712,N_6655);
or U6903 (N_6903,N_6770,N_6555);
or U6904 (N_6904,N_6623,N_6577);
or U6905 (N_6905,N_6562,N_6586);
nor U6906 (N_6906,N_6540,N_6483);
nand U6907 (N_6907,N_6774,N_6522);
nor U6908 (N_6908,N_6528,N_6418);
nor U6909 (N_6909,N_6667,N_6662);
or U6910 (N_6910,N_6646,N_6671);
and U6911 (N_6911,N_6521,N_6686);
nor U6912 (N_6912,N_6544,N_6511);
and U6913 (N_6913,N_6696,N_6452);
or U6914 (N_6914,N_6565,N_6702);
or U6915 (N_6915,N_6629,N_6497);
xnor U6916 (N_6916,N_6450,N_6532);
and U6917 (N_6917,N_6538,N_6457);
or U6918 (N_6918,N_6573,N_6711);
nand U6919 (N_6919,N_6561,N_6625);
xnor U6920 (N_6920,N_6460,N_6464);
and U6921 (N_6921,N_6636,N_6657);
nand U6922 (N_6922,N_6431,N_6672);
xnor U6923 (N_6923,N_6619,N_6781);
nor U6924 (N_6924,N_6580,N_6519);
or U6925 (N_6925,N_6423,N_6787);
nor U6926 (N_6926,N_6404,N_6487);
and U6927 (N_6927,N_6514,N_6769);
xor U6928 (N_6928,N_6425,N_6406);
or U6929 (N_6929,N_6495,N_6679);
nor U6930 (N_6930,N_6756,N_6677);
nor U6931 (N_6931,N_6683,N_6482);
and U6932 (N_6932,N_6533,N_6474);
and U6933 (N_6933,N_6434,N_6593);
xor U6934 (N_6934,N_6415,N_6736);
or U6935 (N_6935,N_6567,N_6591);
and U6936 (N_6936,N_6730,N_6650);
nand U6937 (N_6937,N_6794,N_6772);
or U6938 (N_6938,N_6574,N_6728);
nor U6939 (N_6939,N_6506,N_6509);
nand U6940 (N_6940,N_6496,N_6436);
nor U6941 (N_6941,N_6737,N_6654);
xnor U6942 (N_6942,N_6659,N_6603);
or U6943 (N_6943,N_6611,N_6695);
and U6944 (N_6944,N_6668,N_6797);
or U6945 (N_6945,N_6647,N_6557);
or U6946 (N_6946,N_6700,N_6518);
nand U6947 (N_6947,N_6583,N_6445);
nor U6948 (N_6948,N_6783,N_6720);
nor U6949 (N_6949,N_6628,N_6652);
nand U6950 (N_6950,N_6793,N_6723);
or U6951 (N_6951,N_6687,N_6590);
and U6952 (N_6952,N_6529,N_6523);
nand U6953 (N_6953,N_6790,N_6502);
xor U6954 (N_6954,N_6762,N_6618);
and U6955 (N_6955,N_6447,N_6690);
nor U6956 (N_6956,N_6512,N_6570);
xor U6957 (N_6957,N_6475,N_6697);
or U6958 (N_6958,N_6608,N_6763);
or U6959 (N_6959,N_6409,N_6643);
and U6960 (N_6960,N_6624,N_6607);
and U6961 (N_6961,N_6710,N_6459);
and U6962 (N_6962,N_6491,N_6426);
and U6963 (N_6963,N_6786,N_6648);
nor U6964 (N_6964,N_6744,N_6546);
xor U6965 (N_6965,N_6500,N_6682);
nand U6966 (N_6966,N_6494,N_6779);
or U6967 (N_6967,N_6706,N_6492);
nand U6968 (N_6968,N_6616,N_6420);
xnor U6969 (N_6969,N_6543,N_6458);
xor U6970 (N_6970,N_6751,N_6504);
nand U6971 (N_6971,N_6472,N_6704);
or U6972 (N_6972,N_6622,N_6427);
nand U6973 (N_6973,N_6556,N_6403);
nor U6974 (N_6974,N_6541,N_6778);
xnor U6975 (N_6975,N_6775,N_6620);
or U6976 (N_6976,N_6717,N_6428);
nor U6977 (N_6977,N_6517,N_6466);
nor U6978 (N_6978,N_6694,N_6505);
or U6979 (N_6979,N_6665,N_6456);
nand U6980 (N_6980,N_6453,N_6524);
nor U6981 (N_6981,N_6600,N_6799);
nor U6982 (N_6982,N_6605,N_6765);
and U6983 (N_6983,N_6633,N_6432);
nand U6984 (N_6984,N_6651,N_6560);
nand U6985 (N_6985,N_6708,N_6433);
nor U6986 (N_6986,N_6592,N_6422);
nand U6987 (N_6987,N_6649,N_6531);
xor U6988 (N_6988,N_6419,N_6416);
nand U6989 (N_6989,N_6468,N_6621);
xnor U6990 (N_6990,N_6632,N_6703);
nand U6991 (N_6991,N_6726,N_6716);
or U6992 (N_6992,N_6515,N_6773);
and U6993 (N_6993,N_6534,N_6588);
or U6994 (N_6994,N_6692,N_6429);
nor U6995 (N_6995,N_6764,N_6451);
and U6996 (N_6996,N_6597,N_6613);
nor U6997 (N_6997,N_6479,N_6784);
nand U6998 (N_6998,N_6470,N_6789);
xor U6999 (N_6999,N_6449,N_6701);
or U7000 (N_7000,N_6704,N_6483);
and U7001 (N_7001,N_6590,N_6570);
nor U7002 (N_7002,N_6665,N_6563);
nor U7003 (N_7003,N_6599,N_6467);
nor U7004 (N_7004,N_6583,N_6472);
and U7005 (N_7005,N_6799,N_6669);
nor U7006 (N_7006,N_6717,N_6579);
or U7007 (N_7007,N_6491,N_6598);
xnor U7008 (N_7008,N_6725,N_6702);
nand U7009 (N_7009,N_6726,N_6403);
nor U7010 (N_7010,N_6519,N_6510);
and U7011 (N_7011,N_6497,N_6479);
nand U7012 (N_7012,N_6570,N_6531);
nor U7013 (N_7013,N_6404,N_6418);
or U7014 (N_7014,N_6476,N_6778);
or U7015 (N_7015,N_6540,N_6556);
nand U7016 (N_7016,N_6437,N_6434);
nand U7017 (N_7017,N_6590,N_6497);
and U7018 (N_7018,N_6540,N_6529);
or U7019 (N_7019,N_6572,N_6401);
nand U7020 (N_7020,N_6636,N_6704);
xor U7021 (N_7021,N_6545,N_6751);
or U7022 (N_7022,N_6496,N_6761);
nand U7023 (N_7023,N_6609,N_6776);
nand U7024 (N_7024,N_6519,N_6593);
nand U7025 (N_7025,N_6406,N_6671);
or U7026 (N_7026,N_6433,N_6686);
xnor U7027 (N_7027,N_6418,N_6703);
nand U7028 (N_7028,N_6648,N_6431);
nor U7029 (N_7029,N_6472,N_6434);
and U7030 (N_7030,N_6458,N_6746);
or U7031 (N_7031,N_6544,N_6632);
nor U7032 (N_7032,N_6557,N_6432);
nor U7033 (N_7033,N_6601,N_6620);
xor U7034 (N_7034,N_6665,N_6572);
xor U7035 (N_7035,N_6756,N_6778);
or U7036 (N_7036,N_6697,N_6651);
nor U7037 (N_7037,N_6459,N_6787);
or U7038 (N_7038,N_6619,N_6567);
xor U7039 (N_7039,N_6749,N_6450);
nor U7040 (N_7040,N_6683,N_6498);
xor U7041 (N_7041,N_6467,N_6483);
nor U7042 (N_7042,N_6763,N_6546);
xnor U7043 (N_7043,N_6480,N_6675);
or U7044 (N_7044,N_6517,N_6681);
xnor U7045 (N_7045,N_6635,N_6721);
and U7046 (N_7046,N_6686,N_6596);
nand U7047 (N_7047,N_6546,N_6465);
nand U7048 (N_7048,N_6572,N_6685);
xor U7049 (N_7049,N_6467,N_6568);
xor U7050 (N_7050,N_6726,N_6703);
nor U7051 (N_7051,N_6603,N_6781);
nor U7052 (N_7052,N_6701,N_6799);
or U7053 (N_7053,N_6426,N_6541);
nand U7054 (N_7054,N_6756,N_6796);
nand U7055 (N_7055,N_6538,N_6500);
and U7056 (N_7056,N_6609,N_6449);
or U7057 (N_7057,N_6649,N_6500);
xor U7058 (N_7058,N_6509,N_6657);
nand U7059 (N_7059,N_6756,N_6431);
and U7060 (N_7060,N_6416,N_6482);
nand U7061 (N_7061,N_6590,N_6449);
and U7062 (N_7062,N_6424,N_6787);
and U7063 (N_7063,N_6579,N_6624);
or U7064 (N_7064,N_6670,N_6796);
and U7065 (N_7065,N_6515,N_6659);
nand U7066 (N_7066,N_6547,N_6780);
nand U7067 (N_7067,N_6520,N_6641);
nand U7068 (N_7068,N_6468,N_6493);
xnor U7069 (N_7069,N_6622,N_6545);
or U7070 (N_7070,N_6630,N_6626);
xnor U7071 (N_7071,N_6462,N_6524);
xnor U7072 (N_7072,N_6579,N_6669);
nand U7073 (N_7073,N_6542,N_6712);
and U7074 (N_7074,N_6499,N_6736);
nor U7075 (N_7075,N_6524,N_6473);
xor U7076 (N_7076,N_6539,N_6737);
xnor U7077 (N_7077,N_6678,N_6517);
nand U7078 (N_7078,N_6473,N_6559);
or U7079 (N_7079,N_6605,N_6489);
xor U7080 (N_7080,N_6450,N_6700);
and U7081 (N_7081,N_6737,N_6764);
and U7082 (N_7082,N_6721,N_6592);
xnor U7083 (N_7083,N_6530,N_6700);
and U7084 (N_7084,N_6766,N_6466);
nand U7085 (N_7085,N_6690,N_6468);
nor U7086 (N_7086,N_6484,N_6711);
and U7087 (N_7087,N_6770,N_6629);
nor U7088 (N_7088,N_6766,N_6722);
or U7089 (N_7089,N_6735,N_6743);
nand U7090 (N_7090,N_6715,N_6571);
or U7091 (N_7091,N_6462,N_6452);
nand U7092 (N_7092,N_6772,N_6594);
xnor U7093 (N_7093,N_6788,N_6620);
nor U7094 (N_7094,N_6441,N_6594);
xor U7095 (N_7095,N_6579,N_6703);
and U7096 (N_7096,N_6718,N_6513);
xor U7097 (N_7097,N_6767,N_6608);
nand U7098 (N_7098,N_6708,N_6627);
and U7099 (N_7099,N_6669,N_6498);
nor U7100 (N_7100,N_6492,N_6447);
nor U7101 (N_7101,N_6407,N_6477);
nand U7102 (N_7102,N_6674,N_6488);
nand U7103 (N_7103,N_6674,N_6678);
xor U7104 (N_7104,N_6788,N_6428);
or U7105 (N_7105,N_6594,N_6589);
xnor U7106 (N_7106,N_6709,N_6485);
nor U7107 (N_7107,N_6551,N_6681);
and U7108 (N_7108,N_6658,N_6464);
or U7109 (N_7109,N_6713,N_6732);
nor U7110 (N_7110,N_6781,N_6483);
and U7111 (N_7111,N_6615,N_6584);
and U7112 (N_7112,N_6708,N_6795);
nand U7113 (N_7113,N_6621,N_6678);
nor U7114 (N_7114,N_6707,N_6720);
nand U7115 (N_7115,N_6681,N_6663);
nand U7116 (N_7116,N_6440,N_6611);
and U7117 (N_7117,N_6702,N_6790);
or U7118 (N_7118,N_6626,N_6663);
nor U7119 (N_7119,N_6721,N_6486);
and U7120 (N_7120,N_6706,N_6743);
nand U7121 (N_7121,N_6601,N_6420);
nor U7122 (N_7122,N_6501,N_6606);
or U7123 (N_7123,N_6716,N_6684);
nor U7124 (N_7124,N_6673,N_6735);
and U7125 (N_7125,N_6623,N_6544);
xnor U7126 (N_7126,N_6655,N_6678);
or U7127 (N_7127,N_6509,N_6540);
and U7128 (N_7128,N_6753,N_6774);
xor U7129 (N_7129,N_6469,N_6503);
xor U7130 (N_7130,N_6485,N_6741);
xnor U7131 (N_7131,N_6409,N_6734);
nor U7132 (N_7132,N_6669,N_6777);
or U7133 (N_7133,N_6736,N_6605);
xnor U7134 (N_7134,N_6489,N_6704);
nor U7135 (N_7135,N_6746,N_6520);
or U7136 (N_7136,N_6642,N_6495);
nand U7137 (N_7137,N_6743,N_6793);
nand U7138 (N_7138,N_6710,N_6402);
or U7139 (N_7139,N_6508,N_6770);
nor U7140 (N_7140,N_6657,N_6488);
and U7141 (N_7141,N_6646,N_6755);
or U7142 (N_7142,N_6553,N_6766);
xor U7143 (N_7143,N_6526,N_6740);
or U7144 (N_7144,N_6732,N_6549);
nand U7145 (N_7145,N_6748,N_6794);
nor U7146 (N_7146,N_6735,N_6712);
nor U7147 (N_7147,N_6556,N_6671);
nor U7148 (N_7148,N_6538,N_6707);
xnor U7149 (N_7149,N_6764,N_6664);
nand U7150 (N_7150,N_6508,N_6658);
xor U7151 (N_7151,N_6706,N_6604);
and U7152 (N_7152,N_6711,N_6743);
or U7153 (N_7153,N_6723,N_6441);
and U7154 (N_7154,N_6538,N_6459);
nor U7155 (N_7155,N_6736,N_6467);
xor U7156 (N_7156,N_6798,N_6472);
nor U7157 (N_7157,N_6647,N_6525);
and U7158 (N_7158,N_6480,N_6463);
xor U7159 (N_7159,N_6429,N_6439);
xor U7160 (N_7160,N_6628,N_6705);
xnor U7161 (N_7161,N_6465,N_6716);
xnor U7162 (N_7162,N_6447,N_6664);
nor U7163 (N_7163,N_6434,N_6684);
or U7164 (N_7164,N_6485,N_6488);
nor U7165 (N_7165,N_6618,N_6768);
and U7166 (N_7166,N_6517,N_6685);
and U7167 (N_7167,N_6713,N_6599);
or U7168 (N_7168,N_6463,N_6599);
nor U7169 (N_7169,N_6784,N_6639);
xnor U7170 (N_7170,N_6473,N_6601);
and U7171 (N_7171,N_6758,N_6608);
nand U7172 (N_7172,N_6633,N_6479);
and U7173 (N_7173,N_6644,N_6643);
nand U7174 (N_7174,N_6795,N_6791);
or U7175 (N_7175,N_6467,N_6468);
xnor U7176 (N_7176,N_6725,N_6643);
or U7177 (N_7177,N_6659,N_6720);
nor U7178 (N_7178,N_6657,N_6593);
xnor U7179 (N_7179,N_6755,N_6403);
nor U7180 (N_7180,N_6748,N_6553);
and U7181 (N_7181,N_6667,N_6547);
and U7182 (N_7182,N_6620,N_6709);
nand U7183 (N_7183,N_6751,N_6604);
and U7184 (N_7184,N_6728,N_6444);
or U7185 (N_7185,N_6618,N_6542);
nor U7186 (N_7186,N_6768,N_6639);
nand U7187 (N_7187,N_6541,N_6572);
nand U7188 (N_7188,N_6402,N_6737);
nor U7189 (N_7189,N_6468,N_6785);
xor U7190 (N_7190,N_6693,N_6738);
nor U7191 (N_7191,N_6505,N_6647);
xor U7192 (N_7192,N_6534,N_6475);
and U7193 (N_7193,N_6747,N_6686);
or U7194 (N_7194,N_6481,N_6429);
and U7195 (N_7195,N_6722,N_6656);
xnor U7196 (N_7196,N_6419,N_6400);
xor U7197 (N_7197,N_6709,N_6451);
or U7198 (N_7198,N_6731,N_6534);
and U7199 (N_7199,N_6405,N_6403);
nand U7200 (N_7200,N_6805,N_7034);
and U7201 (N_7201,N_6982,N_6954);
or U7202 (N_7202,N_6886,N_6952);
nor U7203 (N_7203,N_6955,N_7058);
nand U7204 (N_7204,N_6896,N_6822);
and U7205 (N_7205,N_6826,N_6844);
and U7206 (N_7206,N_6997,N_6861);
or U7207 (N_7207,N_6972,N_6808);
xor U7208 (N_7208,N_6813,N_6841);
nor U7209 (N_7209,N_6857,N_7155);
and U7210 (N_7210,N_7071,N_6869);
and U7211 (N_7211,N_6996,N_6807);
nor U7212 (N_7212,N_6817,N_6838);
nand U7213 (N_7213,N_6986,N_7054);
xnor U7214 (N_7214,N_6919,N_7135);
nand U7215 (N_7215,N_6821,N_6984);
and U7216 (N_7216,N_6883,N_6932);
xor U7217 (N_7217,N_6943,N_7077);
and U7218 (N_7218,N_6944,N_6905);
and U7219 (N_7219,N_7009,N_6999);
and U7220 (N_7220,N_7117,N_7067);
xnor U7221 (N_7221,N_6866,N_7037);
nand U7222 (N_7222,N_7146,N_6918);
or U7223 (N_7223,N_6985,N_6819);
or U7224 (N_7224,N_6892,N_6978);
and U7225 (N_7225,N_7191,N_7196);
nand U7226 (N_7226,N_6897,N_7113);
nor U7227 (N_7227,N_7199,N_7049);
nand U7228 (N_7228,N_7073,N_7131);
nor U7229 (N_7229,N_7072,N_6827);
and U7230 (N_7230,N_7013,N_7129);
and U7231 (N_7231,N_7019,N_7087);
nor U7232 (N_7232,N_7064,N_6882);
nand U7233 (N_7233,N_7176,N_6872);
and U7234 (N_7234,N_6811,N_7099);
nand U7235 (N_7235,N_7024,N_7151);
xor U7236 (N_7236,N_7132,N_7125);
xor U7237 (N_7237,N_6967,N_7080);
or U7238 (N_7238,N_7090,N_7189);
nor U7239 (N_7239,N_6823,N_7123);
xnor U7240 (N_7240,N_7011,N_6963);
nand U7241 (N_7241,N_6814,N_7041);
or U7242 (N_7242,N_6878,N_7102);
nand U7243 (N_7243,N_6865,N_6829);
nand U7244 (N_7244,N_6847,N_7078);
nor U7245 (N_7245,N_6895,N_7120);
nand U7246 (N_7246,N_7053,N_6891);
and U7247 (N_7247,N_7181,N_7167);
nor U7248 (N_7248,N_7021,N_7086);
nor U7249 (N_7249,N_7142,N_6816);
and U7250 (N_7250,N_7192,N_7154);
and U7251 (N_7251,N_7153,N_6924);
xnor U7252 (N_7252,N_7098,N_7145);
xnor U7253 (N_7253,N_7180,N_7114);
and U7254 (N_7254,N_7187,N_6949);
and U7255 (N_7255,N_6854,N_7140);
or U7256 (N_7256,N_7137,N_6917);
or U7257 (N_7257,N_7081,N_7124);
or U7258 (N_7258,N_7036,N_6804);
and U7259 (N_7259,N_7101,N_6965);
nor U7260 (N_7260,N_7110,N_6968);
or U7261 (N_7261,N_7195,N_7052);
xnor U7262 (N_7262,N_6927,N_6910);
nor U7263 (N_7263,N_7109,N_6842);
and U7264 (N_7264,N_7055,N_7068);
nand U7265 (N_7265,N_6818,N_6975);
nor U7266 (N_7266,N_6906,N_7126);
or U7267 (N_7267,N_7043,N_6974);
and U7268 (N_7268,N_6911,N_7027);
and U7269 (N_7269,N_7118,N_6947);
nand U7270 (N_7270,N_6843,N_6929);
xor U7271 (N_7271,N_6830,N_7088);
xor U7272 (N_7272,N_7143,N_7062);
and U7273 (N_7273,N_7119,N_7133);
nand U7274 (N_7274,N_6839,N_6976);
and U7275 (N_7275,N_6942,N_6907);
nor U7276 (N_7276,N_6858,N_7121);
xnor U7277 (N_7277,N_7075,N_6991);
nor U7278 (N_7278,N_6931,N_7008);
xor U7279 (N_7279,N_7168,N_7048);
xor U7280 (N_7280,N_6980,N_6928);
or U7281 (N_7281,N_7004,N_7023);
and U7282 (N_7282,N_6935,N_7045);
nand U7283 (N_7283,N_7104,N_6983);
nor U7284 (N_7284,N_6998,N_6902);
or U7285 (N_7285,N_6930,N_7061);
xnor U7286 (N_7286,N_7163,N_7093);
nor U7287 (N_7287,N_7046,N_6990);
nor U7288 (N_7288,N_7177,N_6912);
nand U7289 (N_7289,N_6987,N_6870);
or U7290 (N_7290,N_7183,N_6874);
and U7291 (N_7291,N_7094,N_7148);
nor U7292 (N_7292,N_7175,N_7158);
xnor U7293 (N_7293,N_7018,N_7105);
xor U7294 (N_7294,N_7091,N_7127);
nor U7295 (N_7295,N_6994,N_6936);
and U7296 (N_7296,N_6938,N_6853);
nand U7297 (N_7297,N_6840,N_6939);
or U7298 (N_7298,N_7122,N_6846);
and U7299 (N_7299,N_7097,N_7178);
nand U7300 (N_7300,N_6849,N_6899);
nand U7301 (N_7301,N_7152,N_7005);
and U7302 (N_7302,N_6989,N_6873);
and U7303 (N_7303,N_6877,N_7160);
nor U7304 (N_7304,N_6966,N_6964);
or U7305 (N_7305,N_7107,N_7128);
xnor U7306 (N_7306,N_7059,N_6973);
nand U7307 (N_7307,N_6923,N_7063);
nor U7308 (N_7308,N_7111,N_6950);
nand U7309 (N_7309,N_6979,N_7001);
nor U7310 (N_7310,N_7016,N_7115);
and U7311 (N_7311,N_7002,N_7050);
nand U7312 (N_7312,N_6914,N_6926);
nand U7313 (N_7313,N_7116,N_6925);
nor U7314 (N_7314,N_6993,N_7159);
xnor U7315 (N_7315,N_7079,N_6806);
nand U7316 (N_7316,N_7188,N_7056);
nor U7317 (N_7317,N_7022,N_6888);
and U7318 (N_7318,N_6836,N_6981);
nand U7319 (N_7319,N_6995,N_7170);
and U7320 (N_7320,N_7136,N_6800);
or U7321 (N_7321,N_7095,N_6848);
xnor U7322 (N_7322,N_6958,N_7190);
nor U7323 (N_7323,N_6894,N_7179);
nor U7324 (N_7324,N_6832,N_7156);
xnor U7325 (N_7325,N_7089,N_6835);
nand U7326 (N_7326,N_7103,N_7134);
and U7327 (N_7327,N_6833,N_6922);
and U7328 (N_7328,N_7051,N_6890);
nor U7329 (N_7329,N_6864,N_6916);
nand U7330 (N_7330,N_7042,N_6862);
or U7331 (N_7331,N_7014,N_6940);
nand U7332 (N_7332,N_7000,N_7017);
or U7333 (N_7333,N_7185,N_7029);
xnor U7334 (N_7334,N_7007,N_7169);
nor U7335 (N_7335,N_7040,N_6957);
and U7336 (N_7336,N_6837,N_6937);
nor U7337 (N_7337,N_7174,N_6915);
nand U7338 (N_7338,N_6815,N_7039);
nor U7339 (N_7339,N_7084,N_6856);
and U7340 (N_7340,N_7096,N_6810);
and U7341 (N_7341,N_7070,N_6908);
nor U7342 (N_7342,N_6956,N_6850);
or U7343 (N_7343,N_7038,N_7066);
and U7344 (N_7344,N_6884,N_7069);
or U7345 (N_7345,N_7065,N_6992);
nor U7346 (N_7346,N_7161,N_6901);
nor U7347 (N_7347,N_6904,N_7197);
and U7348 (N_7348,N_7141,N_6988);
nor U7349 (N_7349,N_7182,N_6977);
xnor U7350 (N_7350,N_7157,N_6880);
or U7351 (N_7351,N_6825,N_7060);
nand U7352 (N_7352,N_6852,N_7082);
and U7353 (N_7353,N_6860,N_7076);
xor U7354 (N_7354,N_7150,N_7130);
nor U7355 (N_7355,N_6969,N_7020);
nor U7356 (N_7356,N_6898,N_6933);
nor U7357 (N_7357,N_6868,N_7044);
or U7358 (N_7358,N_6831,N_6953);
and U7359 (N_7359,N_7172,N_6889);
nand U7360 (N_7360,N_6941,N_6970);
nand U7361 (N_7361,N_7144,N_7012);
and U7362 (N_7362,N_7186,N_7166);
nand U7363 (N_7363,N_6961,N_7171);
nand U7364 (N_7364,N_7164,N_6900);
or U7365 (N_7365,N_7083,N_7147);
nand U7366 (N_7366,N_6863,N_6802);
xor U7367 (N_7367,N_7106,N_7085);
nor U7368 (N_7368,N_6909,N_7162);
or U7369 (N_7369,N_6920,N_6879);
or U7370 (N_7370,N_6934,N_7165);
or U7371 (N_7371,N_7194,N_6828);
nand U7372 (N_7372,N_7057,N_6820);
xor U7373 (N_7373,N_6845,N_6948);
and U7374 (N_7374,N_7112,N_6824);
or U7375 (N_7375,N_7047,N_7028);
nand U7376 (N_7376,N_6959,N_7032);
or U7377 (N_7377,N_7138,N_7026);
or U7378 (N_7378,N_7184,N_7173);
nand U7379 (N_7379,N_6809,N_7025);
nand U7380 (N_7380,N_6859,N_7074);
nand U7381 (N_7381,N_6885,N_6875);
or U7382 (N_7382,N_6851,N_6855);
nor U7383 (N_7383,N_6876,N_7149);
and U7384 (N_7384,N_6971,N_6946);
nand U7385 (N_7385,N_7035,N_6834);
or U7386 (N_7386,N_6962,N_6867);
nor U7387 (N_7387,N_6801,N_7193);
nand U7388 (N_7388,N_6887,N_7010);
and U7389 (N_7389,N_6871,N_7198);
nor U7390 (N_7390,N_6960,N_6881);
or U7391 (N_7391,N_6945,N_7092);
nand U7392 (N_7392,N_7139,N_7030);
nor U7393 (N_7393,N_7100,N_6951);
xnor U7394 (N_7394,N_7006,N_7031);
xnor U7395 (N_7395,N_6893,N_7108);
xor U7396 (N_7396,N_6803,N_6903);
or U7397 (N_7397,N_7015,N_7003);
nand U7398 (N_7398,N_6812,N_6913);
nand U7399 (N_7399,N_6921,N_7033);
and U7400 (N_7400,N_7104,N_6911);
nor U7401 (N_7401,N_7143,N_7018);
xnor U7402 (N_7402,N_7163,N_7140);
xor U7403 (N_7403,N_6844,N_7103);
or U7404 (N_7404,N_6817,N_6803);
or U7405 (N_7405,N_7124,N_6839);
and U7406 (N_7406,N_6878,N_6928);
and U7407 (N_7407,N_7032,N_6985);
xnor U7408 (N_7408,N_7186,N_6922);
and U7409 (N_7409,N_6880,N_7080);
or U7410 (N_7410,N_7085,N_7108);
and U7411 (N_7411,N_6949,N_7082);
nand U7412 (N_7412,N_7109,N_6972);
and U7413 (N_7413,N_7011,N_6979);
and U7414 (N_7414,N_6900,N_6911);
or U7415 (N_7415,N_6981,N_7026);
nand U7416 (N_7416,N_7002,N_7106);
and U7417 (N_7417,N_7179,N_6800);
and U7418 (N_7418,N_6928,N_6844);
nand U7419 (N_7419,N_7028,N_7139);
nand U7420 (N_7420,N_7069,N_7048);
nor U7421 (N_7421,N_6865,N_6991);
nand U7422 (N_7422,N_6860,N_7110);
xor U7423 (N_7423,N_6952,N_6927);
nand U7424 (N_7424,N_6982,N_6852);
or U7425 (N_7425,N_7190,N_6881);
nand U7426 (N_7426,N_6997,N_7126);
nor U7427 (N_7427,N_7007,N_7087);
nor U7428 (N_7428,N_7104,N_7116);
nand U7429 (N_7429,N_7011,N_7055);
nand U7430 (N_7430,N_7038,N_6998);
xnor U7431 (N_7431,N_7199,N_7162);
nor U7432 (N_7432,N_6984,N_6935);
and U7433 (N_7433,N_6866,N_7118);
or U7434 (N_7434,N_7091,N_6838);
nand U7435 (N_7435,N_7057,N_7091);
and U7436 (N_7436,N_6990,N_7188);
or U7437 (N_7437,N_7180,N_6941);
nand U7438 (N_7438,N_7183,N_7165);
or U7439 (N_7439,N_7002,N_7090);
and U7440 (N_7440,N_7074,N_7038);
nor U7441 (N_7441,N_6927,N_6999);
xnor U7442 (N_7442,N_7115,N_6948);
nor U7443 (N_7443,N_6845,N_6935);
xor U7444 (N_7444,N_6985,N_6975);
and U7445 (N_7445,N_6994,N_6824);
xor U7446 (N_7446,N_7171,N_6817);
nand U7447 (N_7447,N_7095,N_7092);
nor U7448 (N_7448,N_7188,N_6822);
xnor U7449 (N_7449,N_7125,N_6995);
xor U7450 (N_7450,N_7020,N_7170);
nand U7451 (N_7451,N_7021,N_7194);
and U7452 (N_7452,N_6817,N_6993);
nor U7453 (N_7453,N_7175,N_7008);
or U7454 (N_7454,N_7142,N_7009);
and U7455 (N_7455,N_7021,N_7158);
and U7456 (N_7456,N_6836,N_7018);
nand U7457 (N_7457,N_6923,N_6803);
nand U7458 (N_7458,N_6985,N_7044);
or U7459 (N_7459,N_7190,N_6827);
xnor U7460 (N_7460,N_7053,N_6979);
and U7461 (N_7461,N_6914,N_6944);
nor U7462 (N_7462,N_7153,N_6841);
and U7463 (N_7463,N_7070,N_7163);
or U7464 (N_7464,N_7170,N_6847);
nor U7465 (N_7465,N_6801,N_7009);
xor U7466 (N_7466,N_6981,N_6921);
nand U7467 (N_7467,N_7036,N_6835);
nor U7468 (N_7468,N_7161,N_6899);
and U7469 (N_7469,N_6949,N_7058);
nor U7470 (N_7470,N_7086,N_7133);
and U7471 (N_7471,N_7102,N_6831);
and U7472 (N_7472,N_6916,N_7078);
xor U7473 (N_7473,N_6833,N_7053);
and U7474 (N_7474,N_7098,N_7118);
or U7475 (N_7475,N_7029,N_7187);
nand U7476 (N_7476,N_6932,N_6833);
and U7477 (N_7477,N_6998,N_7135);
and U7478 (N_7478,N_6918,N_7190);
xor U7479 (N_7479,N_7052,N_7051);
xor U7480 (N_7480,N_7098,N_6949);
and U7481 (N_7481,N_6846,N_7084);
nor U7482 (N_7482,N_7125,N_6896);
nor U7483 (N_7483,N_6946,N_7031);
nor U7484 (N_7484,N_7192,N_6926);
xor U7485 (N_7485,N_7148,N_7067);
xnor U7486 (N_7486,N_6828,N_6958);
nand U7487 (N_7487,N_6816,N_7062);
and U7488 (N_7488,N_6958,N_7182);
or U7489 (N_7489,N_6982,N_6824);
xnor U7490 (N_7490,N_6896,N_6919);
and U7491 (N_7491,N_7051,N_7187);
and U7492 (N_7492,N_6953,N_6913);
xnor U7493 (N_7493,N_7061,N_6959);
nor U7494 (N_7494,N_6932,N_7183);
xor U7495 (N_7495,N_7129,N_7091);
or U7496 (N_7496,N_6898,N_7085);
or U7497 (N_7497,N_7171,N_7019);
xnor U7498 (N_7498,N_6886,N_7170);
xor U7499 (N_7499,N_6812,N_7108);
xor U7500 (N_7500,N_7075,N_7189);
or U7501 (N_7501,N_7077,N_6992);
nand U7502 (N_7502,N_7112,N_6919);
nor U7503 (N_7503,N_6870,N_7116);
nor U7504 (N_7504,N_6891,N_6978);
nand U7505 (N_7505,N_7178,N_6931);
or U7506 (N_7506,N_6870,N_6972);
or U7507 (N_7507,N_6988,N_6830);
xnor U7508 (N_7508,N_6942,N_7147);
xor U7509 (N_7509,N_6933,N_7148);
nand U7510 (N_7510,N_6917,N_6965);
xnor U7511 (N_7511,N_7084,N_6841);
and U7512 (N_7512,N_6903,N_6800);
or U7513 (N_7513,N_6926,N_6924);
nor U7514 (N_7514,N_7112,N_7179);
nand U7515 (N_7515,N_7047,N_6961);
nand U7516 (N_7516,N_6890,N_6912);
and U7517 (N_7517,N_6847,N_7179);
nand U7518 (N_7518,N_7067,N_7022);
or U7519 (N_7519,N_7087,N_7017);
xnor U7520 (N_7520,N_7194,N_7171);
or U7521 (N_7521,N_6856,N_6810);
and U7522 (N_7522,N_6848,N_7100);
and U7523 (N_7523,N_6832,N_6921);
and U7524 (N_7524,N_7142,N_6814);
or U7525 (N_7525,N_6890,N_6901);
nand U7526 (N_7526,N_7123,N_6853);
nand U7527 (N_7527,N_7173,N_6999);
nor U7528 (N_7528,N_7062,N_7186);
nand U7529 (N_7529,N_7068,N_7043);
nand U7530 (N_7530,N_6840,N_7047);
or U7531 (N_7531,N_7006,N_7190);
and U7532 (N_7532,N_6949,N_6955);
nand U7533 (N_7533,N_7187,N_6817);
nor U7534 (N_7534,N_6941,N_6890);
nor U7535 (N_7535,N_6906,N_7032);
or U7536 (N_7536,N_6957,N_6947);
and U7537 (N_7537,N_7023,N_6979);
nand U7538 (N_7538,N_6807,N_6825);
nand U7539 (N_7539,N_6947,N_7097);
and U7540 (N_7540,N_6899,N_6983);
or U7541 (N_7541,N_7120,N_7005);
xor U7542 (N_7542,N_7192,N_6852);
and U7543 (N_7543,N_6983,N_6829);
nand U7544 (N_7544,N_7008,N_7138);
and U7545 (N_7545,N_7121,N_6842);
nand U7546 (N_7546,N_6984,N_6828);
xor U7547 (N_7547,N_6958,N_7003);
nor U7548 (N_7548,N_7100,N_6834);
xnor U7549 (N_7549,N_7031,N_6912);
xnor U7550 (N_7550,N_6859,N_7050);
nand U7551 (N_7551,N_7089,N_6984);
or U7552 (N_7552,N_7184,N_6804);
nand U7553 (N_7553,N_6862,N_7143);
nor U7554 (N_7554,N_6940,N_7196);
or U7555 (N_7555,N_7034,N_6982);
xnor U7556 (N_7556,N_6927,N_7170);
and U7557 (N_7557,N_6957,N_6825);
nor U7558 (N_7558,N_7044,N_7060);
nand U7559 (N_7559,N_6921,N_6879);
and U7560 (N_7560,N_7170,N_6889);
and U7561 (N_7561,N_6894,N_7036);
nand U7562 (N_7562,N_6910,N_6878);
nor U7563 (N_7563,N_7034,N_7172);
nand U7564 (N_7564,N_6855,N_6863);
nand U7565 (N_7565,N_7030,N_7170);
and U7566 (N_7566,N_6922,N_7085);
nand U7567 (N_7567,N_7056,N_6988);
xnor U7568 (N_7568,N_6859,N_6903);
and U7569 (N_7569,N_7018,N_7057);
xnor U7570 (N_7570,N_6843,N_6859);
and U7571 (N_7571,N_6802,N_6824);
or U7572 (N_7572,N_6998,N_7043);
and U7573 (N_7573,N_6825,N_6939);
nand U7574 (N_7574,N_6894,N_7081);
nor U7575 (N_7575,N_7152,N_6822);
nor U7576 (N_7576,N_6991,N_7080);
or U7577 (N_7577,N_7020,N_7160);
or U7578 (N_7578,N_6933,N_7079);
nor U7579 (N_7579,N_7064,N_7074);
nand U7580 (N_7580,N_7134,N_7004);
nor U7581 (N_7581,N_7010,N_7059);
nand U7582 (N_7582,N_6944,N_6886);
nor U7583 (N_7583,N_6841,N_6837);
nor U7584 (N_7584,N_6823,N_6809);
xnor U7585 (N_7585,N_7031,N_6889);
or U7586 (N_7586,N_6834,N_6902);
or U7587 (N_7587,N_7146,N_7179);
xor U7588 (N_7588,N_6895,N_6885);
nor U7589 (N_7589,N_6998,N_6936);
xnor U7590 (N_7590,N_7101,N_7056);
and U7591 (N_7591,N_7169,N_7126);
nor U7592 (N_7592,N_7087,N_6816);
nor U7593 (N_7593,N_7180,N_7149);
xor U7594 (N_7594,N_6987,N_6854);
nand U7595 (N_7595,N_7007,N_7079);
nor U7596 (N_7596,N_6932,N_6904);
nand U7597 (N_7597,N_7105,N_6815);
or U7598 (N_7598,N_7191,N_6925);
and U7599 (N_7599,N_7064,N_6916);
nand U7600 (N_7600,N_7492,N_7263);
and U7601 (N_7601,N_7562,N_7389);
nand U7602 (N_7602,N_7307,N_7418);
xor U7603 (N_7603,N_7211,N_7279);
nand U7604 (N_7604,N_7590,N_7358);
nand U7605 (N_7605,N_7564,N_7527);
nor U7606 (N_7606,N_7469,N_7282);
and U7607 (N_7607,N_7368,N_7526);
nand U7608 (N_7608,N_7322,N_7258);
or U7609 (N_7609,N_7437,N_7490);
nand U7610 (N_7610,N_7364,N_7424);
nand U7611 (N_7611,N_7524,N_7550);
nor U7612 (N_7612,N_7503,N_7331);
or U7613 (N_7613,N_7433,N_7381);
nor U7614 (N_7614,N_7598,N_7295);
nor U7615 (N_7615,N_7445,N_7241);
nand U7616 (N_7616,N_7391,N_7560);
nor U7617 (N_7617,N_7595,N_7313);
xnor U7618 (N_7618,N_7430,N_7372);
and U7619 (N_7619,N_7464,N_7229);
xnor U7620 (N_7620,N_7513,N_7544);
and U7621 (N_7621,N_7559,N_7403);
or U7622 (N_7622,N_7380,N_7537);
nor U7623 (N_7623,N_7556,N_7435);
nor U7624 (N_7624,N_7300,N_7589);
nand U7625 (N_7625,N_7554,N_7382);
nand U7626 (N_7626,N_7428,N_7592);
and U7627 (N_7627,N_7470,N_7512);
and U7628 (N_7628,N_7579,N_7432);
xor U7629 (N_7629,N_7434,N_7213);
or U7630 (N_7630,N_7359,N_7305);
and U7631 (N_7631,N_7581,N_7265);
nand U7632 (N_7632,N_7309,N_7580);
nor U7633 (N_7633,N_7320,N_7422);
xnor U7634 (N_7634,N_7293,N_7427);
nor U7635 (N_7635,N_7509,N_7318);
xnor U7636 (N_7636,N_7269,N_7489);
and U7637 (N_7637,N_7262,N_7543);
xor U7638 (N_7638,N_7458,N_7573);
xor U7639 (N_7639,N_7499,N_7374);
or U7640 (N_7640,N_7249,N_7370);
or U7641 (N_7641,N_7316,N_7412);
nor U7642 (N_7642,N_7261,N_7367);
xor U7643 (N_7643,N_7467,N_7463);
nor U7644 (N_7644,N_7586,N_7376);
or U7645 (N_7645,N_7506,N_7485);
and U7646 (N_7646,N_7563,N_7337);
nand U7647 (N_7647,N_7207,N_7245);
and U7648 (N_7648,N_7284,N_7341);
and U7649 (N_7649,N_7253,N_7288);
nor U7650 (N_7650,N_7471,N_7399);
nor U7651 (N_7651,N_7466,N_7294);
nor U7652 (N_7652,N_7345,N_7408);
nor U7653 (N_7653,N_7244,N_7203);
xor U7654 (N_7654,N_7461,N_7395);
xor U7655 (N_7655,N_7232,N_7326);
nor U7656 (N_7656,N_7344,N_7465);
and U7657 (N_7657,N_7250,N_7377);
nand U7658 (N_7658,N_7439,N_7555);
nand U7659 (N_7659,N_7501,N_7247);
or U7660 (N_7660,N_7327,N_7353);
and U7661 (N_7661,N_7330,N_7361);
and U7662 (N_7662,N_7311,N_7278);
nand U7663 (N_7663,N_7477,N_7453);
or U7664 (N_7664,N_7219,N_7301);
or U7665 (N_7665,N_7240,N_7446);
or U7666 (N_7666,N_7267,N_7396);
and U7667 (N_7667,N_7498,N_7587);
nand U7668 (N_7668,N_7285,N_7574);
and U7669 (N_7669,N_7291,N_7483);
or U7670 (N_7670,N_7457,N_7354);
or U7671 (N_7671,N_7576,N_7378);
xnor U7672 (N_7672,N_7369,N_7302);
and U7673 (N_7673,N_7541,N_7460);
nor U7674 (N_7674,N_7516,N_7243);
xor U7675 (N_7675,N_7222,N_7390);
nor U7676 (N_7676,N_7292,N_7238);
and U7677 (N_7677,N_7549,N_7406);
xnor U7678 (N_7678,N_7475,N_7518);
nand U7679 (N_7679,N_7546,N_7479);
and U7680 (N_7680,N_7228,N_7522);
and U7681 (N_7681,N_7597,N_7591);
nor U7682 (N_7682,N_7450,N_7454);
nor U7683 (N_7683,N_7443,N_7266);
and U7684 (N_7684,N_7405,N_7514);
or U7685 (N_7685,N_7568,N_7552);
and U7686 (N_7686,N_7303,N_7317);
nor U7687 (N_7687,N_7565,N_7478);
nand U7688 (N_7688,N_7264,N_7411);
xnor U7689 (N_7689,N_7515,N_7342);
and U7690 (N_7690,N_7414,N_7335);
nand U7691 (N_7691,N_7304,N_7500);
and U7692 (N_7692,N_7504,N_7472);
or U7693 (N_7693,N_7388,N_7336);
or U7694 (N_7694,N_7480,N_7398);
or U7695 (N_7695,N_7575,N_7363);
xor U7696 (N_7696,N_7206,N_7417);
and U7697 (N_7697,N_7255,N_7277);
nor U7698 (N_7698,N_7375,N_7507);
or U7699 (N_7699,N_7547,N_7481);
nor U7700 (N_7700,N_7431,N_7231);
or U7701 (N_7701,N_7553,N_7223);
and U7702 (N_7702,N_7462,N_7404);
xnor U7703 (N_7703,N_7355,N_7334);
xor U7704 (N_7704,N_7421,N_7594);
nand U7705 (N_7705,N_7349,N_7494);
nor U7706 (N_7706,N_7415,N_7227);
nand U7707 (N_7707,N_7209,N_7347);
or U7708 (N_7708,N_7217,N_7438);
or U7709 (N_7709,N_7281,N_7324);
or U7710 (N_7710,N_7360,N_7257);
and U7711 (N_7711,N_7224,N_7254);
nor U7712 (N_7712,N_7202,N_7436);
xor U7713 (N_7713,N_7452,N_7319);
or U7714 (N_7714,N_7387,N_7413);
xnor U7715 (N_7715,N_7487,N_7429);
or U7716 (N_7716,N_7416,N_7280);
xor U7717 (N_7717,N_7212,N_7273);
and U7718 (N_7718,N_7205,N_7409);
xnor U7719 (N_7719,N_7521,N_7297);
xor U7720 (N_7720,N_7299,N_7315);
nand U7721 (N_7721,N_7572,N_7239);
xnor U7722 (N_7722,N_7286,N_7508);
or U7723 (N_7723,N_7287,N_7225);
and U7724 (N_7724,N_7571,N_7296);
or U7725 (N_7725,N_7351,N_7226);
and U7726 (N_7726,N_7531,N_7407);
or U7727 (N_7727,N_7365,N_7237);
nor U7728 (N_7728,N_7270,N_7420);
nand U7729 (N_7729,N_7523,N_7567);
or U7730 (N_7730,N_7423,N_7449);
or U7731 (N_7731,N_7338,N_7511);
xnor U7732 (N_7732,N_7519,N_7275);
or U7733 (N_7733,N_7333,N_7566);
nor U7734 (N_7734,N_7548,N_7357);
or U7735 (N_7735,N_7397,N_7384);
and U7736 (N_7736,N_7383,N_7259);
xnor U7737 (N_7737,N_7393,N_7283);
or U7738 (N_7738,N_7584,N_7312);
nand U7739 (N_7739,N_7473,N_7352);
nand U7740 (N_7740,N_7234,N_7588);
nor U7741 (N_7741,N_7538,N_7529);
and U7742 (N_7742,N_7385,N_7379);
or U7743 (N_7743,N_7310,N_7290);
or U7744 (N_7744,N_7525,N_7271);
xnor U7745 (N_7745,N_7235,N_7208);
nand U7746 (N_7746,N_7289,N_7426);
nand U7747 (N_7747,N_7323,N_7496);
and U7748 (N_7748,N_7371,N_7356);
xor U7749 (N_7749,N_7468,N_7419);
xor U7750 (N_7750,N_7339,N_7491);
and U7751 (N_7751,N_7488,N_7325);
nand U7752 (N_7752,N_7201,N_7348);
and U7753 (N_7753,N_7248,N_7459);
and U7754 (N_7754,N_7394,N_7332);
or U7755 (N_7755,N_7210,N_7321);
nor U7756 (N_7756,N_7246,N_7570);
or U7757 (N_7757,N_7272,N_7366);
xnor U7758 (N_7758,N_7493,N_7593);
nand U7759 (N_7759,N_7536,N_7447);
nor U7760 (N_7760,N_7328,N_7252);
or U7761 (N_7761,N_7410,N_7340);
or U7762 (N_7762,N_7204,N_7596);
nor U7763 (N_7763,N_7441,N_7242);
nor U7764 (N_7764,N_7578,N_7401);
or U7765 (N_7765,N_7535,N_7551);
nand U7766 (N_7766,N_7442,N_7215);
xor U7767 (N_7767,N_7482,N_7214);
or U7768 (N_7768,N_7534,N_7599);
nor U7769 (N_7769,N_7392,N_7569);
nor U7770 (N_7770,N_7505,N_7425);
or U7771 (N_7771,N_7484,N_7533);
or U7772 (N_7772,N_7510,N_7274);
nor U7773 (N_7773,N_7350,N_7542);
nor U7774 (N_7774,N_7540,N_7545);
xor U7775 (N_7775,N_7308,N_7520);
xnor U7776 (N_7776,N_7220,N_7557);
or U7777 (N_7777,N_7362,N_7455);
nand U7778 (N_7778,N_7440,N_7517);
xor U7779 (N_7779,N_7476,N_7268);
or U7780 (N_7780,N_7233,N_7314);
nor U7781 (N_7781,N_7251,N_7386);
nor U7782 (N_7782,N_7306,N_7528);
nand U7783 (N_7783,N_7346,N_7276);
and U7784 (N_7784,N_7495,N_7402);
nand U7785 (N_7785,N_7236,N_7530);
nand U7786 (N_7786,N_7343,N_7577);
and U7787 (N_7787,N_7474,N_7329);
nand U7788 (N_7788,N_7400,N_7582);
nor U7789 (N_7789,N_7585,N_7502);
or U7790 (N_7790,N_7221,N_7558);
xor U7791 (N_7791,N_7218,N_7497);
nor U7792 (N_7792,N_7230,N_7486);
and U7793 (N_7793,N_7298,N_7200);
or U7794 (N_7794,N_7256,N_7583);
xnor U7795 (N_7795,N_7260,N_7539);
and U7796 (N_7796,N_7373,N_7532);
nand U7797 (N_7797,N_7448,N_7216);
nand U7798 (N_7798,N_7444,N_7456);
nor U7799 (N_7799,N_7451,N_7561);
or U7800 (N_7800,N_7297,N_7523);
xnor U7801 (N_7801,N_7513,N_7242);
and U7802 (N_7802,N_7379,N_7260);
or U7803 (N_7803,N_7321,N_7533);
nor U7804 (N_7804,N_7545,N_7351);
xor U7805 (N_7805,N_7393,N_7429);
or U7806 (N_7806,N_7347,N_7338);
nor U7807 (N_7807,N_7511,N_7464);
nor U7808 (N_7808,N_7273,N_7393);
nand U7809 (N_7809,N_7450,N_7458);
nor U7810 (N_7810,N_7378,N_7260);
xnor U7811 (N_7811,N_7538,N_7480);
xor U7812 (N_7812,N_7356,N_7203);
nor U7813 (N_7813,N_7597,N_7316);
nand U7814 (N_7814,N_7377,N_7285);
nor U7815 (N_7815,N_7274,N_7269);
or U7816 (N_7816,N_7595,N_7552);
nor U7817 (N_7817,N_7443,N_7465);
xnor U7818 (N_7818,N_7525,N_7449);
or U7819 (N_7819,N_7280,N_7203);
nor U7820 (N_7820,N_7346,N_7347);
and U7821 (N_7821,N_7255,N_7397);
and U7822 (N_7822,N_7330,N_7540);
xnor U7823 (N_7823,N_7529,N_7413);
nor U7824 (N_7824,N_7596,N_7460);
nand U7825 (N_7825,N_7451,N_7557);
xnor U7826 (N_7826,N_7495,N_7485);
nor U7827 (N_7827,N_7219,N_7481);
nor U7828 (N_7828,N_7485,N_7416);
xor U7829 (N_7829,N_7325,N_7476);
nand U7830 (N_7830,N_7358,N_7291);
nand U7831 (N_7831,N_7375,N_7565);
nor U7832 (N_7832,N_7583,N_7508);
nor U7833 (N_7833,N_7478,N_7347);
and U7834 (N_7834,N_7456,N_7324);
or U7835 (N_7835,N_7247,N_7409);
nor U7836 (N_7836,N_7219,N_7316);
or U7837 (N_7837,N_7539,N_7409);
xnor U7838 (N_7838,N_7266,N_7263);
or U7839 (N_7839,N_7312,N_7500);
or U7840 (N_7840,N_7593,N_7347);
and U7841 (N_7841,N_7496,N_7563);
and U7842 (N_7842,N_7224,N_7210);
xor U7843 (N_7843,N_7435,N_7507);
and U7844 (N_7844,N_7362,N_7565);
or U7845 (N_7845,N_7401,N_7484);
xnor U7846 (N_7846,N_7522,N_7318);
or U7847 (N_7847,N_7447,N_7213);
xor U7848 (N_7848,N_7541,N_7254);
and U7849 (N_7849,N_7368,N_7577);
or U7850 (N_7850,N_7524,N_7288);
and U7851 (N_7851,N_7213,N_7561);
nand U7852 (N_7852,N_7323,N_7286);
xnor U7853 (N_7853,N_7561,N_7554);
and U7854 (N_7854,N_7343,N_7233);
nor U7855 (N_7855,N_7532,N_7272);
nand U7856 (N_7856,N_7542,N_7424);
and U7857 (N_7857,N_7212,N_7241);
nor U7858 (N_7858,N_7396,N_7319);
nor U7859 (N_7859,N_7512,N_7518);
nor U7860 (N_7860,N_7438,N_7576);
nor U7861 (N_7861,N_7320,N_7529);
or U7862 (N_7862,N_7576,N_7441);
nor U7863 (N_7863,N_7478,N_7284);
xor U7864 (N_7864,N_7287,N_7224);
nor U7865 (N_7865,N_7208,N_7340);
xor U7866 (N_7866,N_7344,N_7591);
nand U7867 (N_7867,N_7560,N_7531);
nor U7868 (N_7868,N_7228,N_7239);
xnor U7869 (N_7869,N_7310,N_7554);
nand U7870 (N_7870,N_7383,N_7468);
xor U7871 (N_7871,N_7322,N_7214);
and U7872 (N_7872,N_7363,N_7582);
xnor U7873 (N_7873,N_7412,N_7591);
or U7874 (N_7874,N_7260,N_7300);
and U7875 (N_7875,N_7310,N_7584);
nor U7876 (N_7876,N_7533,N_7264);
xnor U7877 (N_7877,N_7255,N_7355);
nand U7878 (N_7878,N_7237,N_7256);
and U7879 (N_7879,N_7470,N_7249);
or U7880 (N_7880,N_7575,N_7527);
nor U7881 (N_7881,N_7478,N_7316);
xnor U7882 (N_7882,N_7453,N_7222);
nor U7883 (N_7883,N_7505,N_7419);
or U7884 (N_7884,N_7474,N_7360);
or U7885 (N_7885,N_7518,N_7466);
xnor U7886 (N_7886,N_7566,N_7331);
xor U7887 (N_7887,N_7406,N_7341);
nor U7888 (N_7888,N_7371,N_7224);
nor U7889 (N_7889,N_7514,N_7375);
nand U7890 (N_7890,N_7405,N_7517);
nand U7891 (N_7891,N_7295,N_7442);
or U7892 (N_7892,N_7363,N_7423);
and U7893 (N_7893,N_7349,N_7268);
or U7894 (N_7894,N_7585,N_7570);
nor U7895 (N_7895,N_7293,N_7342);
nand U7896 (N_7896,N_7280,N_7580);
and U7897 (N_7897,N_7516,N_7283);
nor U7898 (N_7898,N_7277,N_7437);
nor U7899 (N_7899,N_7547,N_7498);
and U7900 (N_7900,N_7232,N_7559);
nand U7901 (N_7901,N_7573,N_7563);
nand U7902 (N_7902,N_7484,N_7529);
nor U7903 (N_7903,N_7282,N_7260);
xor U7904 (N_7904,N_7575,N_7222);
or U7905 (N_7905,N_7498,N_7265);
nand U7906 (N_7906,N_7463,N_7263);
nor U7907 (N_7907,N_7480,N_7304);
nand U7908 (N_7908,N_7265,N_7575);
or U7909 (N_7909,N_7317,N_7548);
nand U7910 (N_7910,N_7380,N_7239);
nor U7911 (N_7911,N_7346,N_7351);
nand U7912 (N_7912,N_7203,N_7366);
nor U7913 (N_7913,N_7551,N_7362);
or U7914 (N_7914,N_7578,N_7251);
or U7915 (N_7915,N_7204,N_7484);
nand U7916 (N_7916,N_7471,N_7475);
and U7917 (N_7917,N_7517,N_7504);
and U7918 (N_7918,N_7587,N_7303);
xor U7919 (N_7919,N_7349,N_7498);
and U7920 (N_7920,N_7416,N_7341);
nand U7921 (N_7921,N_7201,N_7264);
or U7922 (N_7922,N_7580,N_7589);
xor U7923 (N_7923,N_7214,N_7349);
or U7924 (N_7924,N_7520,N_7310);
or U7925 (N_7925,N_7449,N_7329);
nand U7926 (N_7926,N_7391,N_7416);
nor U7927 (N_7927,N_7377,N_7463);
nand U7928 (N_7928,N_7349,N_7216);
and U7929 (N_7929,N_7281,N_7273);
nor U7930 (N_7930,N_7352,N_7355);
or U7931 (N_7931,N_7464,N_7518);
nor U7932 (N_7932,N_7553,N_7360);
xor U7933 (N_7933,N_7381,N_7594);
nor U7934 (N_7934,N_7367,N_7520);
and U7935 (N_7935,N_7373,N_7371);
nand U7936 (N_7936,N_7551,N_7494);
xor U7937 (N_7937,N_7308,N_7357);
nor U7938 (N_7938,N_7453,N_7237);
nand U7939 (N_7939,N_7404,N_7319);
and U7940 (N_7940,N_7501,N_7432);
xnor U7941 (N_7941,N_7436,N_7520);
nand U7942 (N_7942,N_7203,N_7331);
nand U7943 (N_7943,N_7423,N_7462);
nor U7944 (N_7944,N_7492,N_7316);
nand U7945 (N_7945,N_7549,N_7456);
and U7946 (N_7946,N_7488,N_7435);
or U7947 (N_7947,N_7410,N_7263);
and U7948 (N_7948,N_7209,N_7503);
xnor U7949 (N_7949,N_7513,N_7226);
or U7950 (N_7950,N_7269,N_7508);
xnor U7951 (N_7951,N_7457,N_7559);
and U7952 (N_7952,N_7407,N_7414);
nand U7953 (N_7953,N_7552,N_7495);
or U7954 (N_7954,N_7281,N_7598);
or U7955 (N_7955,N_7598,N_7420);
nor U7956 (N_7956,N_7273,N_7270);
or U7957 (N_7957,N_7514,N_7537);
and U7958 (N_7958,N_7246,N_7435);
and U7959 (N_7959,N_7208,N_7238);
or U7960 (N_7960,N_7361,N_7344);
nor U7961 (N_7961,N_7430,N_7494);
xnor U7962 (N_7962,N_7505,N_7267);
nand U7963 (N_7963,N_7435,N_7220);
or U7964 (N_7964,N_7463,N_7480);
or U7965 (N_7965,N_7317,N_7409);
and U7966 (N_7966,N_7202,N_7299);
and U7967 (N_7967,N_7224,N_7214);
nor U7968 (N_7968,N_7501,N_7591);
and U7969 (N_7969,N_7526,N_7201);
or U7970 (N_7970,N_7283,N_7460);
and U7971 (N_7971,N_7523,N_7501);
and U7972 (N_7972,N_7363,N_7551);
or U7973 (N_7973,N_7466,N_7428);
xor U7974 (N_7974,N_7548,N_7558);
xor U7975 (N_7975,N_7235,N_7272);
nand U7976 (N_7976,N_7547,N_7511);
nor U7977 (N_7977,N_7259,N_7340);
and U7978 (N_7978,N_7521,N_7206);
and U7979 (N_7979,N_7413,N_7419);
or U7980 (N_7980,N_7441,N_7385);
and U7981 (N_7981,N_7519,N_7397);
xnor U7982 (N_7982,N_7569,N_7376);
and U7983 (N_7983,N_7307,N_7357);
xor U7984 (N_7984,N_7304,N_7577);
and U7985 (N_7985,N_7419,N_7393);
nand U7986 (N_7986,N_7210,N_7463);
nand U7987 (N_7987,N_7314,N_7560);
nand U7988 (N_7988,N_7526,N_7466);
nor U7989 (N_7989,N_7573,N_7362);
xor U7990 (N_7990,N_7559,N_7523);
nor U7991 (N_7991,N_7290,N_7321);
nor U7992 (N_7992,N_7348,N_7370);
nand U7993 (N_7993,N_7365,N_7434);
nor U7994 (N_7994,N_7429,N_7205);
and U7995 (N_7995,N_7242,N_7444);
or U7996 (N_7996,N_7420,N_7494);
nand U7997 (N_7997,N_7557,N_7571);
and U7998 (N_7998,N_7548,N_7396);
xor U7999 (N_7999,N_7426,N_7240);
nand U8000 (N_8000,N_7675,N_7963);
nand U8001 (N_8001,N_7663,N_7689);
nor U8002 (N_8002,N_7834,N_7729);
nor U8003 (N_8003,N_7617,N_7662);
nor U8004 (N_8004,N_7779,N_7700);
nor U8005 (N_8005,N_7873,N_7616);
and U8006 (N_8006,N_7864,N_7913);
nor U8007 (N_8007,N_7870,N_7695);
or U8008 (N_8008,N_7709,N_7904);
and U8009 (N_8009,N_7838,N_7799);
or U8010 (N_8010,N_7882,N_7981);
or U8011 (N_8011,N_7612,N_7766);
nand U8012 (N_8012,N_7807,N_7814);
nor U8013 (N_8013,N_7697,N_7982);
or U8014 (N_8014,N_7725,N_7891);
nor U8015 (N_8015,N_7713,N_7998);
and U8016 (N_8016,N_7993,N_7845);
nand U8017 (N_8017,N_7907,N_7658);
and U8018 (N_8018,N_7951,N_7678);
or U8019 (N_8019,N_7990,N_7996);
and U8020 (N_8020,N_7723,N_7622);
nand U8021 (N_8021,N_7965,N_7832);
xnor U8022 (N_8022,N_7641,N_7906);
nand U8023 (N_8023,N_7682,N_7738);
or U8024 (N_8024,N_7960,N_7936);
or U8025 (N_8025,N_7966,N_7625);
or U8026 (N_8026,N_7929,N_7946);
or U8027 (N_8027,N_7626,N_7915);
and U8028 (N_8028,N_7822,N_7941);
and U8029 (N_8029,N_7706,N_7911);
xor U8030 (N_8030,N_7782,N_7744);
and U8031 (N_8031,N_7645,N_7735);
nor U8032 (N_8032,N_7619,N_7787);
or U8033 (N_8033,N_7773,N_7840);
xnor U8034 (N_8034,N_7847,N_7969);
or U8035 (N_8035,N_7861,N_7742);
or U8036 (N_8036,N_7863,N_7989);
and U8037 (N_8037,N_7755,N_7874);
and U8038 (N_8038,N_7868,N_7602);
and U8039 (N_8039,N_7710,N_7869);
xor U8040 (N_8040,N_7821,N_7705);
nand U8041 (N_8041,N_7659,N_7791);
or U8042 (N_8042,N_7968,N_7926);
nand U8043 (N_8043,N_7778,N_7718);
nand U8044 (N_8044,N_7912,N_7944);
and U8045 (N_8045,N_7885,N_7953);
and U8046 (N_8046,N_7858,N_7649);
xor U8047 (N_8047,N_7698,N_7991);
or U8048 (N_8048,N_7806,N_7740);
and U8049 (N_8049,N_7841,N_7643);
nor U8050 (N_8050,N_7792,N_7939);
nor U8051 (N_8051,N_7974,N_7614);
nor U8052 (N_8052,N_7670,N_7867);
and U8053 (N_8053,N_7727,N_7691);
xnor U8054 (N_8054,N_7642,N_7843);
nand U8055 (N_8055,N_7985,N_7648);
nand U8056 (N_8056,N_7699,N_7788);
and U8057 (N_8057,N_7837,N_7910);
or U8058 (N_8058,N_7997,N_7650);
xor U8059 (N_8059,N_7654,N_7604);
and U8060 (N_8060,N_7608,N_7736);
xnor U8061 (N_8061,N_7835,N_7759);
and U8062 (N_8062,N_7896,N_7784);
or U8063 (N_8063,N_7775,N_7986);
nor U8064 (N_8064,N_7731,N_7655);
xor U8065 (N_8065,N_7620,N_7681);
and U8066 (N_8066,N_7628,N_7739);
or U8067 (N_8067,N_7763,N_7627);
nor U8068 (N_8068,N_7880,N_7865);
nand U8069 (N_8069,N_7859,N_7635);
xnor U8070 (N_8070,N_7828,N_7803);
nor U8071 (N_8071,N_7857,N_7934);
xnor U8072 (N_8072,N_7769,N_7666);
nand U8073 (N_8073,N_7603,N_7606);
or U8074 (N_8074,N_7640,N_7850);
nor U8075 (N_8075,N_7973,N_7937);
and U8076 (N_8076,N_7853,N_7917);
or U8077 (N_8077,N_7632,N_7909);
nor U8078 (N_8078,N_7657,N_7844);
nand U8079 (N_8079,N_7932,N_7730);
nand U8080 (N_8080,N_7772,N_7719);
nor U8081 (N_8081,N_7901,N_7607);
or U8082 (N_8082,N_7902,N_7781);
nor U8083 (N_8083,N_7668,N_7783);
or U8084 (N_8084,N_7667,N_7688);
and U8085 (N_8085,N_7879,N_7983);
or U8086 (N_8086,N_7651,N_7726);
xnor U8087 (N_8087,N_7900,N_7704);
nand U8088 (N_8088,N_7748,N_7754);
nand U8089 (N_8089,N_7961,N_7930);
nor U8090 (N_8090,N_7609,N_7647);
and U8091 (N_8091,N_7798,N_7777);
xor U8092 (N_8092,N_7638,N_7600);
xnor U8093 (N_8093,N_7646,N_7734);
nor U8094 (N_8094,N_7686,N_7800);
nor U8095 (N_8095,N_7976,N_7898);
nand U8096 (N_8096,N_7690,N_7970);
nor U8097 (N_8097,N_7980,N_7862);
or U8098 (N_8098,N_7919,N_7842);
xnor U8099 (N_8099,N_7888,N_7890);
nand U8100 (N_8100,N_7671,N_7673);
nor U8101 (N_8101,N_7825,N_7829);
nor U8102 (N_8102,N_7680,N_7967);
nand U8103 (N_8103,N_7819,N_7687);
nor U8104 (N_8104,N_7899,N_7875);
or U8105 (N_8105,N_7809,N_7639);
and U8106 (N_8106,N_7728,N_7743);
nor U8107 (N_8107,N_7920,N_7786);
xnor U8108 (N_8108,N_7644,N_7872);
or U8109 (N_8109,N_7925,N_7694);
and U8110 (N_8110,N_7979,N_7764);
nand U8111 (N_8111,N_7836,N_7717);
or U8112 (N_8112,N_7672,N_7708);
or U8113 (N_8113,N_7745,N_7988);
nand U8114 (N_8114,N_7685,N_7889);
and U8115 (N_8115,N_7724,N_7751);
or U8116 (N_8116,N_7733,N_7774);
xor U8117 (N_8117,N_7928,N_7796);
xnor U8118 (N_8118,N_7860,N_7707);
xor U8119 (N_8119,N_7720,N_7765);
and U8120 (N_8120,N_7922,N_7992);
nor U8121 (N_8121,N_7601,N_7897);
or U8122 (N_8122,N_7972,N_7737);
nand U8123 (N_8123,N_7802,N_7818);
or U8124 (N_8124,N_7877,N_7676);
xor U8125 (N_8125,N_7615,N_7984);
or U8126 (N_8126,N_7839,N_7940);
and U8127 (N_8127,N_7793,N_7652);
nor U8128 (N_8128,N_7795,N_7831);
nor U8129 (N_8129,N_7701,N_7833);
and U8130 (N_8130,N_7756,N_7947);
and U8131 (N_8131,N_7664,N_7933);
and U8132 (N_8132,N_7894,N_7905);
nand U8133 (N_8133,N_7964,N_7805);
xnor U8134 (N_8134,N_7813,N_7634);
xnor U8135 (N_8135,N_7696,N_7794);
nand U8136 (N_8136,N_7914,N_7752);
nand U8137 (N_8137,N_7624,N_7886);
nand U8138 (N_8138,N_7732,N_7958);
nand U8139 (N_8139,N_7848,N_7661);
nor U8140 (N_8140,N_7776,N_7801);
nand U8141 (N_8141,N_7714,N_7815);
nand U8142 (N_8142,N_7816,N_7811);
xnor U8143 (N_8143,N_7753,N_7820);
and U8144 (N_8144,N_7653,N_7952);
xor U8145 (N_8145,N_7871,N_7935);
nor U8146 (N_8146,N_7780,N_7962);
or U8147 (N_8147,N_7948,N_7679);
nor U8148 (N_8148,N_7903,N_7975);
nand U8149 (N_8149,N_7943,N_7866);
and U8150 (N_8150,N_7804,N_7684);
xnor U8151 (N_8151,N_7895,N_7823);
nor U8152 (N_8152,N_7757,N_7945);
nand U8153 (N_8153,N_7712,N_7767);
or U8154 (N_8154,N_7760,N_7856);
or U8155 (N_8155,N_7750,N_7938);
nand U8156 (N_8156,N_7855,N_7878);
nand U8157 (N_8157,N_7949,N_7851);
or U8158 (N_8158,N_7876,N_7761);
xor U8159 (N_8159,N_7610,N_7630);
and U8160 (N_8160,N_7631,N_7987);
nand U8161 (N_8161,N_7715,N_7605);
xor U8162 (N_8162,N_7824,N_7942);
and U8163 (N_8163,N_7716,N_7722);
and U8164 (N_8164,N_7741,N_7916);
nand U8165 (N_8165,N_7884,N_7956);
xnor U8166 (N_8166,N_7893,N_7995);
nand U8167 (N_8167,N_7827,N_7892);
nand U8168 (N_8168,N_7918,N_7629);
or U8169 (N_8169,N_7817,N_7637);
xor U8170 (N_8170,N_7971,N_7994);
xor U8171 (N_8171,N_7950,N_7957);
xnor U8172 (N_8172,N_7826,N_7613);
nor U8173 (N_8173,N_7618,N_7703);
nand U8174 (N_8174,N_7768,N_7854);
nor U8175 (N_8175,N_7954,N_7623);
nand U8176 (N_8176,N_7746,N_7883);
nand U8177 (N_8177,N_7785,N_7702);
xnor U8178 (N_8178,N_7721,N_7808);
xnor U8179 (N_8179,N_7924,N_7692);
nand U8180 (N_8180,N_7887,N_7611);
or U8181 (N_8181,N_7955,N_7674);
and U8182 (N_8182,N_7849,N_7959);
xor U8183 (N_8183,N_7999,N_7921);
xor U8184 (N_8184,N_7923,N_7830);
or U8185 (N_8185,N_7846,N_7669);
and U8186 (N_8186,N_7977,N_7812);
xnor U8187 (N_8187,N_7656,N_7789);
xor U8188 (N_8188,N_7683,N_7797);
xor U8189 (N_8189,N_7758,N_7749);
and U8190 (N_8190,N_7677,N_7665);
nor U8191 (N_8191,N_7711,N_7762);
nor U8192 (N_8192,N_7931,N_7633);
or U8193 (N_8193,N_7908,N_7771);
nor U8194 (N_8194,N_7770,N_7881);
nand U8195 (N_8195,N_7747,N_7636);
and U8196 (N_8196,N_7978,N_7927);
nor U8197 (N_8197,N_7621,N_7852);
xor U8198 (N_8198,N_7693,N_7810);
nand U8199 (N_8199,N_7660,N_7790);
nor U8200 (N_8200,N_7651,N_7679);
nand U8201 (N_8201,N_7608,N_7893);
and U8202 (N_8202,N_7817,N_7780);
nand U8203 (N_8203,N_7607,N_7627);
nand U8204 (N_8204,N_7982,N_7894);
and U8205 (N_8205,N_7965,N_7850);
xor U8206 (N_8206,N_7644,N_7984);
nor U8207 (N_8207,N_7742,N_7762);
and U8208 (N_8208,N_7822,N_7694);
nor U8209 (N_8209,N_7922,N_7669);
xor U8210 (N_8210,N_7901,N_7853);
xor U8211 (N_8211,N_7656,N_7768);
nor U8212 (N_8212,N_7792,N_7669);
xnor U8213 (N_8213,N_7909,N_7610);
or U8214 (N_8214,N_7621,N_7758);
xnor U8215 (N_8215,N_7635,N_7958);
nand U8216 (N_8216,N_7775,N_7756);
and U8217 (N_8217,N_7696,N_7884);
xnor U8218 (N_8218,N_7785,N_7947);
or U8219 (N_8219,N_7644,N_7737);
nor U8220 (N_8220,N_7609,N_7891);
nand U8221 (N_8221,N_7916,N_7647);
or U8222 (N_8222,N_7677,N_7604);
and U8223 (N_8223,N_7707,N_7970);
nand U8224 (N_8224,N_7684,N_7773);
nand U8225 (N_8225,N_7795,N_7916);
nand U8226 (N_8226,N_7886,N_7964);
xor U8227 (N_8227,N_7653,N_7789);
or U8228 (N_8228,N_7634,N_7760);
and U8229 (N_8229,N_7784,N_7787);
and U8230 (N_8230,N_7713,N_7927);
or U8231 (N_8231,N_7740,N_7757);
or U8232 (N_8232,N_7853,N_7779);
xnor U8233 (N_8233,N_7732,N_7830);
nand U8234 (N_8234,N_7960,N_7644);
xnor U8235 (N_8235,N_7747,N_7773);
nor U8236 (N_8236,N_7965,N_7600);
nand U8237 (N_8237,N_7827,N_7641);
or U8238 (N_8238,N_7936,N_7654);
nand U8239 (N_8239,N_7919,N_7927);
and U8240 (N_8240,N_7948,N_7933);
nand U8241 (N_8241,N_7745,N_7843);
xor U8242 (N_8242,N_7784,N_7800);
xor U8243 (N_8243,N_7667,N_7800);
xnor U8244 (N_8244,N_7716,N_7721);
nor U8245 (N_8245,N_7824,N_7787);
nor U8246 (N_8246,N_7807,N_7911);
xnor U8247 (N_8247,N_7981,N_7726);
or U8248 (N_8248,N_7910,N_7665);
nand U8249 (N_8249,N_7685,N_7832);
nor U8250 (N_8250,N_7879,N_7666);
or U8251 (N_8251,N_7704,N_7713);
or U8252 (N_8252,N_7971,N_7832);
xor U8253 (N_8253,N_7976,N_7870);
or U8254 (N_8254,N_7679,N_7641);
nand U8255 (N_8255,N_7856,N_7652);
nand U8256 (N_8256,N_7658,N_7982);
nand U8257 (N_8257,N_7709,N_7638);
nor U8258 (N_8258,N_7803,N_7988);
nor U8259 (N_8259,N_7990,N_7965);
and U8260 (N_8260,N_7663,N_7613);
or U8261 (N_8261,N_7617,N_7775);
nand U8262 (N_8262,N_7821,N_7718);
or U8263 (N_8263,N_7745,N_7932);
nand U8264 (N_8264,N_7677,N_7800);
or U8265 (N_8265,N_7843,N_7818);
xor U8266 (N_8266,N_7863,N_7789);
or U8267 (N_8267,N_7609,N_7742);
or U8268 (N_8268,N_7644,N_7702);
and U8269 (N_8269,N_7621,N_7960);
or U8270 (N_8270,N_7740,N_7818);
xnor U8271 (N_8271,N_7602,N_7839);
and U8272 (N_8272,N_7601,N_7658);
or U8273 (N_8273,N_7828,N_7714);
nor U8274 (N_8274,N_7755,N_7926);
nand U8275 (N_8275,N_7689,N_7990);
or U8276 (N_8276,N_7828,N_7995);
nor U8277 (N_8277,N_7610,N_7871);
nand U8278 (N_8278,N_7878,N_7786);
nand U8279 (N_8279,N_7908,N_7681);
xnor U8280 (N_8280,N_7921,N_7956);
and U8281 (N_8281,N_7723,N_7727);
and U8282 (N_8282,N_7815,N_7646);
or U8283 (N_8283,N_7822,N_7668);
or U8284 (N_8284,N_7898,N_7711);
nor U8285 (N_8285,N_7833,N_7868);
or U8286 (N_8286,N_7612,N_7678);
or U8287 (N_8287,N_7893,N_7717);
nand U8288 (N_8288,N_7963,N_7735);
xnor U8289 (N_8289,N_7862,N_7764);
xor U8290 (N_8290,N_7713,N_7617);
nor U8291 (N_8291,N_7865,N_7791);
nand U8292 (N_8292,N_7943,N_7823);
nand U8293 (N_8293,N_7851,N_7933);
nor U8294 (N_8294,N_7646,N_7988);
xnor U8295 (N_8295,N_7621,N_7862);
or U8296 (N_8296,N_7885,N_7956);
nor U8297 (N_8297,N_7820,N_7986);
and U8298 (N_8298,N_7721,N_7789);
nor U8299 (N_8299,N_7603,N_7773);
or U8300 (N_8300,N_7703,N_7867);
xnor U8301 (N_8301,N_7732,N_7859);
and U8302 (N_8302,N_7799,N_7852);
nand U8303 (N_8303,N_7969,N_7967);
nand U8304 (N_8304,N_7889,N_7879);
nor U8305 (N_8305,N_7924,N_7953);
or U8306 (N_8306,N_7666,N_7710);
nor U8307 (N_8307,N_7826,N_7752);
nor U8308 (N_8308,N_7961,N_7711);
nor U8309 (N_8309,N_7790,N_7829);
or U8310 (N_8310,N_7616,N_7604);
or U8311 (N_8311,N_7811,N_7772);
xor U8312 (N_8312,N_7696,N_7858);
nor U8313 (N_8313,N_7688,N_7696);
nand U8314 (N_8314,N_7943,N_7904);
nand U8315 (N_8315,N_7772,N_7831);
and U8316 (N_8316,N_7948,N_7628);
xor U8317 (N_8317,N_7901,N_7916);
xnor U8318 (N_8318,N_7854,N_7960);
and U8319 (N_8319,N_7696,N_7713);
and U8320 (N_8320,N_7691,N_7736);
xnor U8321 (N_8321,N_7743,N_7984);
nor U8322 (N_8322,N_7769,N_7892);
nand U8323 (N_8323,N_7918,N_7965);
xor U8324 (N_8324,N_7734,N_7650);
xor U8325 (N_8325,N_7752,N_7667);
and U8326 (N_8326,N_7712,N_7891);
and U8327 (N_8327,N_7843,N_7846);
and U8328 (N_8328,N_7951,N_7829);
and U8329 (N_8329,N_7697,N_7741);
and U8330 (N_8330,N_7753,N_7602);
nor U8331 (N_8331,N_7875,N_7712);
xor U8332 (N_8332,N_7991,N_7665);
xor U8333 (N_8333,N_7601,N_7800);
or U8334 (N_8334,N_7757,N_7886);
and U8335 (N_8335,N_7770,N_7601);
nand U8336 (N_8336,N_7681,N_7790);
nor U8337 (N_8337,N_7829,N_7629);
and U8338 (N_8338,N_7842,N_7728);
or U8339 (N_8339,N_7884,N_7756);
nor U8340 (N_8340,N_7875,N_7843);
nor U8341 (N_8341,N_7990,N_7648);
or U8342 (N_8342,N_7952,N_7976);
or U8343 (N_8343,N_7973,N_7673);
nor U8344 (N_8344,N_7930,N_7886);
or U8345 (N_8345,N_7729,N_7631);
and U8346 (N_8346,N_7646,N_7620);
xnor U8347 (N_8347,N_7724,N_7787);
nor U8348 (N_8348,N_7716,N_7940);
nand U8349 (N_8349,N_7961,N_7695);
or U8350 (N_8350,N_7617,N_7945);
or U8351 (N_8351,N_7647,N_7773);
or U8352 (N_8352,N_7820,N_7620);
nor U8353 (N_8353,N_7627,N_7897);
or U8354 (N_8354,N_7679,N_7984);
nand U8355 (N_8355,N_7715,N_7876);
and U8356 (N_8356,N_7921,N_7828);
or U8357 (N_8357,N_7887,N_7818);
nand U8358 (N_8358,N_7650,N_7848);
and U8359 (N_8359,N_7852,N_7905);
nor U8360 (N_8360,N_7651,N_7805);
and U8361 (N_8361,N_7996,N_7708);
nor U8362 (N_8362,N_7820,N_7958);
nand U8363 (N_8363,N_7605,N_7858);
or U8364 (N_8364,N_7757,N_7658);
xor U8365 (N_8365,N_7709,N_7748);
and U8366 (N_8366,N_7707,N_7810);
nor U8367 (N_8367,N_7679,N_7823);
or U8368 (N_8368,N_7870,N_7974);
nor U8369 (N_8369,N_7748,N_7703);
or U8370 (N_8370,N_7710,N_7920);
nand U8371 (N_8371,N_7658,N_7876);
nor U8372 (N_8372,N_7768,N_7881);
nand U8373 (N_8373,N_7750,N_7890);
nand U8374 (N_8374,N_7738,N_7910);
or U8375 (N_8375,N_7733,N_7855);
nor U8376 (N_8376,N_7695,N_7935);
nor U8377 (N_8377,N_7847,N_7901);
and U8378 (N_8378,N_7608,N_7829);
or U8379 (N_8379,N_7781,N_7799);
nand U8380 (N_8380,N_7793,N_7843);
and U8381 (N_8381,N_7923,N_7959);
or U8382 (N_8382,N_7861,N_7973);
nand U8383 (N_8383,N_7759,N_7650);
nor U8384 (N_8384,N_7794,N_7810);
or U8385 (N_8385,N_7884,N_7827);
or U8386 (N_8386,N_7628,N_7939);
nor U8387 (N_8387,N_7624,N_7841);
and U8388 (N_8388,N_7856,N_7872);
xnor U8389 (N_8389,N_7901,N_7884);
or U8390 (N_8390,N_7658,N_7622);
nor U8391 (N_8391,N_7824,N_7880);
nand U8392 (N_8392,N_7999,N_7852);
nand U8393 (N_8393,N_7650,N_7761);
nand U8394 (N_8394,N_7651,N_7671);
xnor U8395 (N_8395,N_7807,N_7955);
nand U8396 (N_8396,N_7985,N_7708);
xor U8397 (N_8397,N_7821,N_7603);
and U8398 (N_8398,N_7923,N_7833);
nor U8399 (N_8399,N_7773,N_7861);
xnor U8400 (N_8400,N_8367,N_8059);
or U8401 (N_8401,N_8150,N_8183);
nand U8402 (N_8402,N_8247,N_8284);
nand U8403 (N_8403,N_8331,N_8342);
and U8404 (N_8404,N_8161,N_8220);
xor U8405 (N_8405,N_8072,N_8135);
xnor U8406 (N_8406,N_8002,N_8116);
xor U8407 (N_8407,N_8381,N_8211);
xnor U8408 (N_8408,N_8227,N_8393);
or U8409 (N_8409,N_8197,N_8269);
nor U8410 (N_8410,N_8217,N_8365);
xnor U8411 (N_8411,N_8131,N_8222);
nand U8412 (N_8412,N_8094,N_8314);
nor U8413 (N_8413,N_8056,N_8387);
xor U8414 (N_8414,N_8016,N_8057);
xnor U8415 (N_8415,N_8065,N_8190);
xnor U8416 (N_8416,N_8321,N_8088);
nand U8417 (N_8417,N_8117,N_8375);
or U8418 (N_8418,N_8020,N_8185);
nand U8419 (N_8419,N_8276,N_8148);
or U8420 (N_8420,N_8015,N_8089);
nand U8421 (N_8421,N_8093,N_8206);
or U8422 (N_8422,N_8353,N_8319);
nand U8423 (N_8423,N_8005,N_8001);
nor U8424 (N_8424,N_8007,N_8237);
nand U8425 (N_8425,N_8386,N_8310);
nand U8426 (N_8426,N_8109,N_8244);
xnor U8427 (N_8427,N_8078,N_8274);
xnor U8428 (N_8428,N_8344,N_8070);
nor U8429 (N_8429,N_8398,N_8293);
or U8430 (N_8430,N_8242,N_8263);
and U8431 (N_8431,N_8108,N_8379);
xnor U8432 (N_8432,N_8008,N_8160);
and U8433 (N_8433,N_8125,N_8046);
nor U8434 (N_8434,N_8081,N_8324);
nor U8435 (N_8435,N_8282,N_8102);
or U8436 (N_8436,N_8168,N_8045);
xor U8437 (N_8437,N_8240,N_8285);
nor U8438 (N_8438,N_8212,N_8303);
and U8439 (N_8439,N_8066,N_8335);
or U8440 (N_8440,N_8145,N_8171);
or U8441 (N_8441,N_8097,N_8030);
nor U8442 (N_8442,N_8100,N_8062);
nand U8443 (N_8443,N_8351,N_8060);
xor U8444 (N_8444,N_8238,N_8149);
nor U8445 (N_8445,N_8096,N_8166);
nor U8446 (N_8446,N_8343,N_8028);
or U8447 (N_8447,N_8291,N_8076);
nor U8448 (N_8448,N_8064,N_8152);
or U8449 (N_8449,N_8069,N_8235);
xnor U8450 (N_8450,N_8306,N_8083);
xnor U8451 (N_8451,N_8010,N_8213);
or U8452 (N_8452,N_8019,N_8243);
xor U8453 (N_8453,N_8360,N_8195);
xnor U8454 (N_8454,N_8165,N_8281);
and U8455 (N_8455,N_8397,N_8164);
xnor U8456 (N_8456,N_8372,N_8156);
and U8457 (N_8457,N_8175,N_8223);
xor U8458 (N_8458,N_8355,N_8074);
and U8459 (N_8459,N_8170,N_8278);
and U8460 (N_8460,N_8210,N_8399);
or U8461 (N_8461,N_8270,N_8196);
nand U8462 (N_8462,N_8308,N_8391);
and U8463 (N_8463,N_8080,N_8251);
nand U8464 (N_8464,N_8265,N_8396);
or U8465 (N_8465,N_8024,N_8390);
and U8466 (N_8466,N_8043,N_8051);
xnor U8467 (N_8467,N_8176,N_8289);
and U8468 (N_8468,N_8358,N_8252);
and U8469 (N_8469,N_8337,N_8157);
and U8470 (N_8470,N_8249,N_8011);
and U8471 (N_8471,N_8384,N_8328);
nand U8472 (N_8472,N_8132,N_8141);
xnor U8473 (N_8473,N_8086,N_8385);
nor U8474 (N_8474,N_8298,N_8194);
and U8475 (N_8475,N_8061,N_8296);
nor U8476 (N_8476,N_8233,N_8111);
xor U8477 (N_8477,N_8272,N_8101);
nor U8478 (N_8478,N_8262,N_8147);
xor U8479 (N_8479,N_8257,N_8041);
and U8480 (N_8480,N_8120,N_8198);
nand U8481 (N_8481,N_8241,N_8144);
and U8482 (N_8482,N_8146,N_8133);
xnor U8483 (N_8483,N_8162,N_8032);
nand U8484 (N_8484,N_8022,N_8092);
nor U8485 (N_8485,N_8258,N_8373);
or U8486 (N_8486,N_8173,N_8359);
nand U8487 (N_8487,N_8079,N_8026);
and U8488 (N_8488,N_8042,N_8317);
nor U8489 (N_8489,N_8153,N_8394);
nand U8490 (N_8490,N_8049,N_8099);
nor U8491 (N_8491,N_8134,N_8260);
xor U8492 (N_8492,N_8126,N_8169);
and U8493 (N_8493,N_8221,N_8055);
or U8494 (N_8494,N_8151,N_8119);
nand U8495 (N_8495,N_8268,N_8122);
xnor U8496 (N_8496,N_8297,N_8329);
nand U8497 (N_8497,N_8369,N_8186);
and U8498 (N_8498,N_8294,N_8047);
nand U8499 (N_8499,N_8229,N_8259);
nand U8500 (N_8500,N_8128,N_8137);
xnor U8501 (N_8501,N_8143,N_8364);
and U8502 (N_8502,N_8199,N_8366);
nor U8503 (N_8503,N_8037,N_8200);
and U8504 (N_8504,N_8085,N_8218);
or U8505 (N_8505,N_8067,N_8389);
nand U8506 (N_8506,N_8129,N_8036);
and U8507 (N_8507,N_8163,N_8136);
and U8508 (N_8508,N_8280,N_8191);
or U8509 (N_8509,N_8232,N_8215);
nor U8510 (N_8510,N_8225,N_8054);
xnor U8511 (N_8511,N_8264,N_8301);
xor U8512 (N_8512,N_8334,N_8338);
or U8513 (N_8513,N_8124,N_8356);
nand U8514 (N_8514,N_8246,N_8357);
xnor U8515 (N_8515,N_8371,N_8184);
nor U8516 (N_8516,N_8179,N_8346);
or U8517 (N_8517,N_8058,N_8339);
and U8518 (N_8518,N_8110,N_8159);
and U8519 (N_8519,N_8340,N_8350);
xor U8520 (N_8520,N_8003,N_8118);
or U8521 (N_8521,N_8154,N_8341);
xor U8522 (N_8522,N_8138,N_8256);
nor U8523 (N_8523,N_8140,N_8277);
or U8524 (N_8524,N_8300,N_8228);
nand U8525 (N_8525,N_8239,N_8107);
nand U8526 (N_8526,N_8354,N_8031);
or U8527 (N_8527,N_8311,N_8139);
or U8528 (N_8528,N_8320,N_8231);
xor U8529 (N_8529,N_8383,N_8009);
nor U8530 (N_8530,N_8348,N_8382);
and U8531 (N_8531,N_8377,N_8039);
xor U8532 (N_8532,N_8018,N_8236);
and U8533 (N_8533,N_8044,N_8155);
and U8534 (N_8534,N_8035,N_8172);
xor U8535 (N_8535,N_8362,N_8192);
nand U8536 (N_8536,N_8033,N_8275);
or U8537 (N_8537,N_8352,N_8053);
or U8538 (N_8538,N_8370,N_8226);
and U8539 (N_8539,N_8392,N_8267);
xor U8540 (N_8540,N_8112,N_8034);
and U8541 (N_8541,N_8038,N_8273);
and U8542 (N_8542,N_8087,N_8071);
and U8543 (N_8543,N_8084,N_8021);
or U8544 (N_8544,N_8261,N_8177);
nor U8545 (N_8545,N_8204,N_8180);
xnor U8546 (N_8546,N_8368,N_8201);
nor U8547 (N_8547,N_8322,N_8279);
xor U8548 (N_8548,N_8347,N_8315);
xnor U8549 (N_8549,N_8023,N_8349);
and U8550 (N_8550,N_8114,N_8327);
xor U8551 (N_8551,N_8219,N_8063);
xnor U8552 (N_8552,N_8336,N_8295);
or U8553 (N_8553,N_8006,N_8073);
or U8554 (N_8554,N_8013,N_8115);
xor U8555 (N_8555,N_8290,N_8224);
nand U8556 (N_8556,N_8376,N_8316);
xnor U8557 (N_8557,N_8254,N_8181);
nand U8558 (N_8558,N_8105,N_8189);
nor U8559 (N_8559,N_8216,N_8326);
and U8560 (N_8560,N_8325,N_8205);
or U8561 (N_8561,N_8098,N_8253);
or U8562 (N_8562,N_8208,N_8305);
xnor U8563 (N_8563,N_8323,N_8203);
nand U8564 (N_8564,N_8082,N_8130);
xor U8565 (N_8565,N_8017,N_8245);
or U8566 (N_8566,N_8052,N_8178);
or U8567 (N_8567,N_8193,N_8202);
nand U8568 (N_8568,N_8012,N_8075);
nor U8569 (N_8569,N_8266,N_8304);
xor U8570 (N_8570,N_8068,N_8004);
and U8571 (N_8571,N_8127,N_8167);
nand U8572 (N_8572,N_8380,N_8345);
xor U8573 (N_8573,N_8318,N_8332);
xnor U8574 (N_8574,N_8271,N_8174);
and U8575 (N_8575,N_8378,N_8286);
or U8576 (N_8576,N_8374,N_8103);
or U8577 (N_8577,N_8027,N_8299);
nand U8578 (N_8578,N_8248,N_8309);
or U8579 (N_8579,N_8014,N_8029);
xnor U8580 (N_8580,N_8142,N_8307);
nand U8581 (N_8581,N_8361,N_8104);
nand U8582 (N_8582,N_8207,N_8230);
and U8583 (N_8583,N_8312,N_8313);
or U8584 (N_8584,N_8395,N_8214);
xor U8585 (N_8585,N_8000,N_8106);
or U8586 (N_8586,N_8077,N_8090);
nor U8587 (N_8587,N_8388,N_8182);
nand U8588 (N_8588,N_8123,N_8188);
xnor U8589 (N_8589,N_8091,N_8283);
and U8590 (N_8590,N_8025,N_8250);
and U8591 (N_8591,N_8287,N_8288);
nand U8592 (N_8592,N_8040,N_8113);
and U8593 (N_8593,N_8048,N_8363);
xor U8594 (N_8594,N_8209,N_8333);
and U8595 (N_8595,N_8187,N_8158);
nor U8596 (N_8596,N_8121,N_8302);
and U8597 (N_8597,N_8255,N_8330);
nand U8598 (N_8598,N_8292,N_8095);
xor U8599 (N_8599,N_8234,N_8050);
xnor U8600 (N_8600,N_8220,N_8009);
or U8601 (N_8601,N_8366,N_8026);
nor U8602 (N_8602,N_8120,N_8256);
xor U8603 (N_8603,N_8012,N_8019);
nor U8604 (N_8604,N_8241,N_8136);
nand U8605 (N_8605,N_8277,N_8285);
nand U8606 (N_8606,N_8087,N_8229);
xnor U8607 (N_8607,N_8018,N_8119);
xnor U8608 (N_8608,N_8382,N_8190);
xnor U8609 (N_8609,N_8112,N_8382);
and U8610 (N_8610,N_8107,N_8042);
and U8611 (N_8611,N_8019,N_8397);
or U8612 (N_8612,N_8173,N_8213);
and U8613 (N_8613,N_8387,N_8371);
nor U8614 (N_8614,N_8225,N_8386);
xnor U8615 (N_8615,N_8214,N_8056);
xnor U8616 (N_8616,N_8355,N_8159);
and U8617 (N_8617,N_8386,N_8038);
xor U8618 (N_8618,N_8209,N_8240);
and U8619 (N_8619,N_8375,N_8361);
and U8620 (N_8620,N_8266,N_8105);
xnor U8621 (N_8621,N_8312,N_8291);
or U8622 (N_8622,N_8030,N_8275);
nand U8623 (N_8623,N_8108,N_8376);
or U8624 (N_8624,N_8109,N_8270);
nand U8625 (N_8625,N_8086,N_8223);
and U8626 (N_8626,N_8186,N_8247);
xnor U8627 (N_8627,N_8037,N_8031);
nand U8628 (N_8628,N_8061,N_8226);
or U8629 (N_8629,N_8191,N_8338);
nand U8630 (N_8630,N_8167,N_8051);
and U8631 (N_8631,N_8120,N_8389);
nand U8632 (N_8632,N_8179,N_8022);
or U8633 (N_8633,N_8274,N_8380);
xnor U8634 (N_8634,N_8380,N_8212);
xnor U8635 (N_8635,N_8285,N_8148);
xor U8636 (N_8636,N_8103,N_8340);
nand U8637 (N_8637,N_8020,N_8275);
or U8638 (N_8638,N_8072,N_8276);
xor U8639 (N_8639,N_8264,N_8298);
nand U8640 (N_8640,N_8284,N_8050);
nor U8641 (N_8641,N_8109,N_8121);
or U8642 (N_8642,N_8369,N_8394);
nor U8643 (N_8643,N_8152,N_8001);
nand U8644 (N_8644,N_8038,N_8087);
nand U8645 (N_8645,N_8277,N_8074);
or U8646 (N_8646,N_8034,N_8257);
nor U8647 (N_8647,N_8075,N_8065);
nand U8648 (N_8648,N_8028,N_8185);
nand U8649 (N_8649,N_8313,N_8256);
and U8650 (N_8650,N_8337,N_8302);
nand U8651 (N_8651,N_8071,N_8052);
nand U8652 (N_8652,N_8395,N_8223);
nor U8653 (N_8653,N_8209,N_8270);
xor U8654 (N_8654,N_8078,N_8226);
nor U8655 (N_8655,N_8031,N_8212);
xnor U8656 (N_8656,N_8237,N_8329);
xnor U8657 (N_8657,N_8254,N_8048);
or U8658 (N_8658,N_8268,N_8381);
nand U8659 (N_8659,N_8000,N_8107);
nor U8660 (N_8660,N_8166,N_8347);
xnor U8661 (N_8661,N_8275,N_8013);
and U8662 (N_8662,N_8162,N_8241);
and U8663 (N_8663,N_8325,N_8121);
or U8664 (N_8664,N_8247,N_8036);
nand U8665 (N_8665,N_8390,N_8240);
nand U8666 (N_8666,N_8041,N_8211);
or U8667 (N_8667,N_8223,N_8264);
and U8668 (N_8668,N_8358,N_8056);
xor U8669 (N_8669,N_8339,N_8260);
nand U8670 (N_8670,N_8308,N_8321);
and U8671 (N_8671,N_8224,N_8208);
or U8672 (N_8672,N_8224,N_8354);
xor U8673 (N_8673,N_8128,N_8178);
and U8674 (N_8674,N_8002,N_8080);
and U8675 (N_8675,N_8222,N_8136);
nor U8676 (N_8676,N_8358,N_8305);
nor U8677 (N_8677,N_8224,N_8057);
xnor U8678 (N_8678,N_8215,N_8078);
or U8679 (N_8679,N_8172,N_8268);
nor U8680 (N_8680,N_8168,N_8359);
xor U8681 (N_8681,N_8332,N_8178);
nor U8682 (N_8682,N_8238,N_8192);
nor U8683 (N_8683,N_8031,N_8352);
and U8684 (N_8684,N_8061,N_8294);
and U8685 (N_8685,N_8049,N_8392);
and U8686 (N_8686,N_8206,N_8039);
or U8687 (N_8687,N_8007,N_8058);
nor U8688 (N_8688,N_8145,N_8059);
or U8689 (N_8689,N_8144,N_8157);
or U8690 (N_8690,N_8141,N_8386);
or U8691 (N_8691,N_8227,N_8086);
nor U8692 (N_8692,N_8032,N_8098);
xnor U8693 (N_8693,N_8167,N_8272);
or U8694 (N_8694,N_8081,N_8301);
nor U8695 (N_8695,N_8180,N_8399);
xnor U8696 (N_8696,N_8194,N_8301);
nor U8697 (N_8697,N_8248,N_8396);
and U8698 (N_8698,N_8371,N_8102);
or U8699 (N_8699,N_8090,N_8314);
or U8700 (N_8700,N_8206,N_8041);
and U8701 (N_8701,N_8298,N_8209);
nor U8702 (N_8702,N_8229,N_8108);
xnor U8703 (N_8703,N_8233,N_8083);
nor U8704 (N_8704,N_8201,N_8077);
nor U8705 (N_8705,N_8263,N_8373);
or U8706 (N_8706,N_8138,N_8252);
nor U8707 (N_8707,N_8299,N_8319);
and U8708 (N_8708,N_8037,N_8215);
nand U8709 (N_8709,N_8338,N_8380);
nor U8710 (N_8710,N_8399,N_8310);
nor U8711 (N_8711,N_8009,N_8253);
nor U8712 (N_8712,N_8006,N_8207);
nand U8713 (N_8713,N_8007,N_8083);
or U8714 (N_8714,N_8149,N_8177);
or U8715 (N_8715,N_8234,N_8397);
nand U8716 (N_8716,N_8081,N_8003);
nand U8717 (N_8717,N_8195,N_8155);
or U8718 (N_8718,N_8033,N_8280);
or U8719 (N_8719,N_8070,N_8243);
nand U8720 (N_8720,N_8389,N_8125);
nor U8721 (N_8721,N_8295,N_8000);
xnor U8722 (N_8722,N_8016,N_8055);
or U8723 (N_8723,N_8371,N_8131);
xnor U8724 (N_8724,N_8257,N_8149);
nand U8725 (N_8725,N_8146,N_8396);
or U8726 (N_8726,N_8325,N_8213);
and U8727 (N_8727,N_8290,N_8035);
or U8728 (N_8728,N_8009,N_8000);
and U8729 (N_8729,N_8245,N_8322);
and U8730 (N_8730,N_8382,N_8305);
and U8731 (N_8731,N_8271,N_8051);
nor U8732 (N_8732,N_8232,N_8089);
nand U8733 (N_8733,N_8281,N_8144);
nand U8734 (N_8734,N_8214,N_8200);
and U8735 (N_8735,N_8379,N_8261);
xnor U8736 (N_8736,N_8107,N_8035);
nand U8737 (N_8737,N_8033,N_8372);
nand U8738 (N_8738,N_8228,N_8222);
nor U8739 (N_8739,N_8185,N_8070);
or U8740 (N_8740,N_8093,N_8134);
xor U8741 (N_8741,N_8052,N_8244);
or U8742 (N_8742,N_8381,N_8223);
nor U8743 (N_8743,N_8056,N_8075);
or U8744 (N_8744,N_8357,N_8331);
xor U8745 (N_8745,N_8208,N_8014);
nand U8746 (N_8746,N_8295,N_8029);
xnor U8747 (N_8747,N_8049,N_8026);
nor U8748 (N_8748,N_8362,N_8026);
and U8749 (N_8749,N_8327,N_8091);
xnor U8750 (N_8750,N_8201,N_8004);
and U8751 (N_8751,N_8008,N_8076);
or U8752 (N_8752,N_8259,N_8357);
and U8753 (N_8753,N_8380,N_8275);
and U8754 (N_8754,N_8343,N_8023);
or U8755 (N_8755,N_8359,N_8160);
or U8756 (N_8756,N_8133,N_8362);
or U8757 (N_8757,N_8343,N_8317);
and U8758 (N_8758,N_8337,N_8085);
nor U8759 (N_8759,N_8300,N_8129);
xor U8760 (N_8760,N_8140,N_8398);
or U8761 (N_8761,N_8130,N_8076);
xor U8762 (N_8762,N_8349,N_8088);
or U8763 (N_8763,N_8299,N_8042);
and U8764 (N_8764,N_8299,N_8392);
nand U8765 (N_8765,N_8127,N_8113);
nor U8766 (N_8766,N_8195,N_8044);
xnor U8767 (N_8767,N_8329,N_8044);
or U8768 (N_8768,N_8073,N_8163);
or U8769 (N_8769,N_8187,N_8175);
and U8770 (N_8770,N_8380,N_8283);
and U8771 (N_8771,N_8324,N_8322);
and U8772 (N_8772,N_8028,N_8252);
nor U8773 (N_8773,N_8197,N_8059);
nand U8774 (N_8774,N_8282,N_8199);
xnor U8775 (N_8775,N_8389,N_8318);
nand U8776 (N_8776,N_8244,N_8082);
nor U8777 (N_8777,N_8240,N_8015);
xor U8778 (N_8778,N_8026,N_8190);
or U8779 (N_8779,N_8099,N_8392);
xnor U8780 (N_8780,N_8091,N_8070);
or U8781 (N_8781,N_8288,N_8281);
and U8782 (N_8782,N_8214,N_8226);
nand U8783 (N_8783,N_8040,N_8016);
nor U8784 (N_8784,N_8021,N_8367);
nor U8785 (N_8785,N_8204,N_8010);
and U8786 (N_8786,N_8060,N_8365);
nand U8787 (N_8787,N_8247,N_8275);
or U8788 (N_8788,N_8305,N_8019);
and U8789 (N_8789,N_8135,N_8388);
xnor U8790 (N_8790,N_8093,N_8255);
xor U8791 (N_8791,N_8008,N_8001);
nor U8792 (N_8792,N_8113,N_8072);
xor U8793 (N_8793,N_8291,N_8077);
nor U8794 (N_8794,N_8131,N_8057);
nand U8795 (N_8795,N_8109,N_8184);
and U8796 (N_8796,N_8247,N_8027);
xor U8797 (N_8797,N_8068,N_8218);
and U8798 (N_8798,N_8123,N_8315);
nor U8799 (N_8799,N_8302,N_8005);
and U8800 (N_8800,N_8573,N_8443);
and U8801 (N_8801,N_8625,N_8407);
xor U8802 (N_8802,N_8642,N_8627);
nand U8803 (N_8803,N_8638,N_8452);
xnor U8804 (N_8804,N_8605,N_8763);
and U8805 (N_8805,N_8715,N_8676);
nor U8806 (N_8806,N_8457,N_8487);
or U8807 (N_8807,N_8532,N_8453);
xor U8808 (N_8808,N_8510,N_8546);
nor U8809 (N_8809,N_8542,N_8795);
or U8810 (N_8810,N_8619,N_8661);
nor U8811 (N_8811,N_8680,N_8583);
nand U8812 (N_8812,N_8408,N_8495);
and U8813 (N_8813,N_8631,N_8422);
and U8814 (N_8814,N_8640,N_8548);
or U8815 (N_8815,N_8691,N_8591);
nand U8816 (N_8816,N_8561,N_8569);
and U8817 (N_8817,N_8481,N_8737);
xor U8818 (N_8818,N_8797,N_8716);
xnor U8819 (N_8819,N_8770,N_8724);
nor U8820 (N_8820,N_8456,N_8576);
xnor U8821 (N_8821,N_8773,N_8506);
nand U8822 (N_8822,N_8632,N_8460);
or U8823 (N_8823,N_8678,N_8410);
and U8824 (N_8824,N_8768,N_8679);
or U8825 (N_8825,N_8504,N_8694);
xor U8826 (N_8826,N_8554,N_8553);
or U8827 (N_8827,N_8497,N_8741);
nor U8828 (N_8828,N_8692,N_8611);
nor U8829 (N_8829,N_8687,N_8586);
nand U8830 (N_8830,N_8693,N_8491);
nand U8831 (N_8831,N_8609,N_8484);
xnor U8832 (N_8832,N_8549,N_8784);
nor U8833 (N_8833,N_8745,N_8656);
nor U8834 (N_8834,N_8430,N_8596);
or U8835 (N_8835,N_8449,N_8507);
and U8836 (N_8836,N_8539,N_8788);
nand U8837 (N_8837,N_8501,N_8413);
nor U8838 (N_8838,N_8525,N_8697);
xor U8839 (N_8839,N_8608,N_8787);
nand U8840 (N_8840,N_8646,N_8555);
and U8841 (N_8841,N_8673,N_8579);
or U8842 (N_8842,N_8782,N_8502);
and U8843 (N_8843,N_8494,N_8550);
nor U8844 (N_8844,N_8654,N_8657);
and U8845 (N_8845,N_8567,N_8723);
or U8846 (N_8846,N_8478,N_8432);
nor U8847 (N_8847,N_8752,N_8755);
xor U8848 (N_8848,N_8485,N_8473);
nand U8849 (N_8849,N_8659,N_8747);
nor U8850 (N_8850,N_8469,N_8614);
or U8851 (N_8851,N_8566,N_8786);
or U8852 (N_8852,N_8447,N_8582);
or U8853 (N_8853,N_8400,N_8604);
or U8854 (N_8854,N_8401,N_8698);
and U8855 (N_8855,N_8645,N_8547);
xnor U8856 (N_8856,N_8695,N_8749);
or U8857 (N_8857,N_8417,N_8533);
and U8858 (N_8858,N_8439,N_8793);
nor U8859 (N_8859,N_8746,N_8492);
or U8860 (N_8860,N_8479,N_8796);
nand U8861 (N_8861,N_8743,N_8458);
and U8862 (N_8862,N_8738,N_8707);
nor U8863 (N_8863,N_8756,N_8498);
nor U8864 (N_8864,N_8534,N_8589);
xor U8865 (N_8865,N_8653,N_8409);
nand U8866 (N_8866,N_8511,N_8489);
nor U8867 (N_8867,N_8736,N_8722);
nor U8868 (N_8868,N_8564,N_8704);
nand U8869 (N_8869,N_8785,N_8674);
xnor U8870 (N_8870,N_8446,N_8617);
and U8871 (N_8871,N_8411,N_8538);
xor U8872 (N_8872,N_8629,N_8558);
xnor U8873 (N_8873,N_8744,N_8630);
xnor U8874 (N_8874,N_8474,N_8414);
and U8875 (N_8875,N_8471,N_8623);
nand U8876 (N_8876,N_8610,N_8593);
nand U8877 (N_8877,N_8717,N_8513);
and U8878 (N_8878,N_8578,N_8696);
and U8879 (N_8879,N_8701,N_8750);
or U8880 (N_8880,N_8650,N_8509);
and U8881 (N_8881,N_8423,N_8636);
nand U8882 (N_8882,N_8733,N_8622);
xor U8883 (N_8883,N_8480,N_8445);
xnor U8884 (N_8884,N_8544,N_8754);
nor U8885 (N_8885,N_8799,N_8767);
and U8886 (N_8886,N_8467,N_8590);
nor U8887 (N_8887,N_8758,N_8455);
nor U8888 (N_8888,N_8552,N_8714);
nand U8889 (N_8889,N_8517,N_8448);
nor U8890 (N_8890,N_8603,N_8644);
and U8891 (N_8891,N_8710,N_8718);
nand U8892 (N_8892,N_8667,N_8626);
and U8893 (N_8893,N_8568,N_8421);
xor U8894 (N_8894,N_8402,N_8519);
and U8895 (N_8895,N_8496,N_8418);
or U8896 (N_8896,N_8686,N_8427);
nand U8897 (N_8897,N_8798,N_8420);
and U8898 (N_8898,N_8643,N_8514);
and U8899 (N_8899,N_8404,N_8442);
nor U8900 (N_8900,N_8634,N_8535);
nor U8901 (N_8901,N_8726,N_8515);
and U8902 (N_8902,N_8669,N_8735);
and U8903 (N_8903,N_8577,N_8776);
and U8904 (N_8904,N_8556,N_8601);
or U8905 (N_8905,N_8599,N_8753);
nand U8906 (N_8906,N_8571,N_8475);
nor U8907 (N_8907,N_8765,N_8703);
and U8908 (N_8908,N_8725,N_8597);
nor U8909 (N_8909,N_8523,N_8477);
or U8910 (N_8910,N_8731,N_8688);
nand U8911 (N_8911,N_8431,N_8563);
and U8912 (N_8912,N_8575,N_8450);
nor U8913 (N_8913,N_8594,N_8434);
and U8914 (N_8914,N_8760,N_8762);
nor U8915 (N_8915,N_8732,N_8468);
and U8916 (N_8916,N_8483,N_8436);
nand U8917 (N_8917,N_8551,N_8665);
nand U8918 (N_8918,N_8499,N_8618);
nor U8919 (N_8919,N_8781,N_8761);
nor U8920 (N_8920,N_8454,N_8406);
and U8921 (N_8921,N_8598,N_8766);
xnor U8922 (N_8922,N_8742,N_8664);
or U8923 (N_8923,N_8412,N_8602);
nor U8924 (N_8924,N_8462,N_8500);
and U8925 (N_8925,N_8764,N_8470);
nand U8926 (N_8926,N_8606,N_8639);
nand U8927 (N_8927,N_8488,N_8588);
and U8928 (N_8928,N_8730,N_8713);
xor U8929 (N_8929,N_8652,N_8415);
and U8930 (N_8930,N_8528,N_8429);
nand U8931 (N_8931,N_8403,N_8647);
or U8932 (N_8932,N_8682,N_8405);
xnor U8933 (N_8933,N_8437,N_8592);
nand U8934 (N_8934,N_8670,N_8702);
or U8935 (N_8935,N_8521,N_8572);
xor U8936 (N_8936,N_8790,N_8655);
and U8937 (N_8937,N_8651,N_8426);
xnor U8938 (N_8938,N_8684,N_8503);
and U8939 (N_8939,N_8791,N_8727);
nand U8940 (N_8940,N_8461,N_8416);
nor U8941 (N_8941,N_8607,N_8672);
xor U8942 (N_8942,N_8600,N_8493);
and U8943 (N_8943,N_8721,N_8775);
nand U8944 (N_8944,N_8574,N_8595);
nor U8945 (N_8945,N_8438,N_8441);
nor U8946 (N_8946,N_8512,N_8621);
nand U8947 (N_8947,N_8587,N_8757);
and U8948 (N_8948,N_8465,N_8641);
nor U8949 (N_8949,N_8580,N_8585);
or U8950 (N_8950,N_8435,N_8671);
and U8951 (N_8951,N_8490,N_8463);
nand U8952 (N_8952,N_8734,N_8581);
xnor U8953 (N_8953,N_8616,N_8508);
xnor U8954 (N_8954,N_8633,N_8759);
xnor U8955 (N_8955,N_8541,N_8543);
and U8956 (N_8956,N_8728,N_8751);
and U8957 (N_8957,N_8482,N_8712);
or U8958 (N_8958,N_8683,N_8648);
nand U8959 (N_8959,N_8557,N_8668);
or U8960 (N_8960,N_8771,N_8425);
nor U8961 (N_8961,N_8689,N_8472);
xnor U8962 (N_8962,N_8560,N_8464);
nor U8963 (N_8963,N_8628,N_8681);
nor U8964 (N_8964,N_8748,N_8565);
nor U8965 (N_8965,N_8615,N_8739);
nor U8966 (N_8966,N_8778,N_8451);
xnor U8967 (N_8967,N_8620,N_8476);
nor U8968 (N_8968,N_8706,N_8537);
xnor U8969 (N_8969,N_8709,N_8531);
xnor U8970 (N_8970,N_8433,N_8675);
nor U8971 (N_8971,N_8624,N_8486);
nor U8972 (N_8972,N_8522,N_8708);
and U8973 (N_8973,N_8792,N_8459);
nand U8974 (N_8974,N_8530,N_8705);
or U8975 (N_8975,N_8777,N_8690);
nand U8976 (N_8976,N_8570,N_8505);
nand U8977 (N_8977,N_8428,N_8562);
and U8978 (N_8978,N_8440,N_8637);
or U8979 (N_8979,N_8779,N_8780);
or U8980 (N_8980,N_8518,N_8584);
and U8981 (N_8981,N_8612,N_8419);
or U8982 (N_8982,N_8444,N_8662);
or U8983 (N_8983,N_8529,N_8666);
nand U8984 (N_8984,N_8729,N_8769);
nand U8985 (N_8985,N_8794,N_8545);
nor U8986 (N_8986,N_8540,N_8719);
nor U8987 (N_8987,N_8649,N_8527);
or U8988 (N_8988,N_8711,N_8524);
xor U8989 (N_8989,N_8613,N_8466);
nand U8990 (N_8990,N_8774,N_8677);
nor U8991 (N_8991,N_8658,N_8699);
xnor U8992 (N_8992,N_8740,N_8424);
xnor U8993 (N_8993,N_8559,N_8783);
xnor U8994 (N_8994,N_8772,N_8789);
and U8995 (N_8995,N_8520,N_8660);
nand U8996 (N_8996,N_8536,N_8635);
or U8997 (N_8997,N_8663,N_8685);
and U8998 (N_8998,N_8526,N_8720);
and U8999 (N_8999,N_8516,N_8700);
nand U9000 (N_9000,N_8532,N_8615);
and U9001 (N_9001,N_8517,N_8648);
or U9002 (N_9002,N_8418,N_8786);
nor U9003 (N_9003,N_8772,N_8723);
or U9004 (N_9004,N_8456,N_8402);
or U9005 (N_9005,N_8663,N_8797);
and U9006 (N_9006,N_8591,N_8746);
xor U9007 (N_9007,N_8656,N_8487);
xnor U9008 (N_9008,N_8631,N_8598);
and U9009 (N_9009,N_8762,N_8528);
and U9010 (N_9010,N_8590,N_8541);
nand U9011 (N_9011,N_8433,N_8670);
xor U9012 (N_9012,N_8634,N_8703);
xor U9013 (N_9013,N_8783,N_8527);
and U9014 (N_9014,N_8412,N_8655);
nand U9015 (N_9015,N_8536,N_8720);
or U9016 (N_9016,N_8451,N_8749);
nor U9017 (N_9017,N_8475,N_8773);
or U9018 (N_9018,N_8616,N_8422);
xor U9019 (N_9019,N_8574,N_8675);
nand U9020 (N_9020,N_8611,N_8735);
and U9021 (N_9021,N_8782,N_8771);
nand U9022 (N_9022,N_8706,N_8541);
and U9023 (N_9023,N_8647,N_8405);
xor U9024 (N_9024,N_8664,N_8504);
or U9025 (N_9025,N_8698,N_8625);
or U9026 (N_9026,N_8707,N_8446);
nor U9027 (N_9027,N_8501,N_8629);
xor U9028 (N_9028,N_8794,N_8479);
nand U9029 (N_9029,N_8527,N_8656);
or U9030 (N_9030,N_8429,N_8645);
nor U9031 (N_9031,N_8701,N_8636);
nor U9032 (N_9032,N_8763,N_8447);
or U9033 (N_9033,N_8712,N_8793);
nand U9034 (N_9034,N_8593,N_8540);
nor U9035 (N_9035,N_8672,N_8591);
nand U9036 (N_9036,N_8586,N_8431);
or U9037 (N_9037,N_8425,N_8794);
nand U9038 (N_9038,N_8434,N_8526);
nor U9039 (N_9039,N_8540,N_8657);
nor U9040 (N_9040,N_8489,N_8669);
nand U9041 (N_9041,N_8553,N_8791);
nand U9042 (N_9042,N_8676,N_8552);
nor U9043 (N_9043,N_8789,N_8794);
and U9044 (N_9044,N_8646,N_8734);
or U9045 (N_9045,N_8673,N_8742);
nand U9046 (N_9046,N_8799,N_8543);
and U9047 (N_9047,N_8791,N_8494);
xor U9048 (N_9048,N_8771,N_8474);
and U9049 (N_9049,N_8649,N_8567);
and U9050 (N_9050,N_8700,N_8576);
nand U9051 (N_9051,N_8466,N_8561);
xor U9052 (N_9052,N_8761,N_8772);
or U9053 (N_9053,N_8558,N_8765);
nor U9054 (N_9054,N_8541,N_8658);
nor U9055 (N_9055,N_8554,N_8617);
and U9056 (N_9056,N_8791,N_8718);
xor U9057 (N_9057,N_8770,N_8651);
and U9058 (N_9058,N_8695,N_8726);
nor U9059 (N_9059,N_8596,N_8746);
xnor U9060 (N_9060,N_8483,N_8504);
or U9061 (N_9061,N_8739,N_8574);
nor U9062 (N_9062,N_8507,N_8755);
nor U9063 (N_9063,N_8575,N_8404);
nand U9064 (N_9064,N_8573,N_8697);
or U9065 (N_9065,N_8631,N_8480);
nor U9066 (N_9066,N_8432,N_8430);
and U9067 (N_9067,N_8548,N_8606);
nor U9068 (N_9068,N_8649,N_8407);
nor U9069 (N_9069,N_8584,N_8753);
xnor U9070 (N_9070,N_8462,N_8472);
or U9071 (N_9071,N_8799,N_8592);
or U9072 (N_9072,N_8453,N_8772);
nor U9073 (N_9073,N_8710,N_8722);
nand U9074 (N_9074,N_8598,N_8574);
nor U9075 (N_9075,N_8727,N_8691);
nor U9076 (N_9076,N_8769,N_8585);
or U9077 (N_9077,N_8427,N_8641);
or U9078 (N_9078,N_8671,N_8734);
nor U9079 (N_9079,N_8445,N_8703);
xor U9080 (N_9080,N_8425,N_8738);
or U9081 (N_9081,N_8697,N_8487);
or U9082 (N_9082,N_8462,N_8547);
nor U9083 (N_9083,N_8452,N_8581);
or U9084 (N_9084,N_8749,N_8477);
or U9085 (N_9085,N_8447,N_8757);
nor U9086 (N_9086,N_8576,N_8643);
nand U9087 (N_9087,N_8707,N_8626);
and U9088 (N_9088,N_8767,N_8535);
nor U9089 (N_9089,N_8695,N_8743);
or U9090 (N_9090,N_8467,N_8780);
and U9091 (N_9091,N_8717,N_8673);
xnor U9092 (N_9092,N_8578,N_8724);
and U9093 (N_9093,N_8537,N_8607);
and U9094 (N_9094,N_8715,N_8707);
and U9095 (N_9095,N_8465,N_8722);
or U9096 (N_9096,N_8719,N_8544);
nand U9097 (N_9097,N_8567,N_8484);
nand U9098 (N_9098,N_8535,N_8697);
xor U9099 (N_9099,N_8658,N_8490);
or U9100 (N_9100,N_8703,N_8741);
or U9101 (N_9101,N_8751,N_8731);
or U9102 (N_9102,N_8584,N_8543);
and U9103 (N_9103,N_8739,N_8549);
nand U9104 (N_9104,N_8761,N_8480);
nand U9105 (N_9105,N_8678,N_8787);
xnor U9106 (N_9106,N_8776,N_8490);
xor U9107 (N_9107,N_8697,N_8467);
or U9108 (N_9108,N_8706,N_8598);
nand U9109 (N_9109,N_8485,N_8655);
and U9110 (N_9110,N_8558,N_8791);
xnor U9111 (N_9111,N_8537,N_8604);
and U9112 (N_9112,N_8556,N_8745);
nand U9113 (N_9113,N_8705,N_8721);
and U9114 (N_9114,N_8615,N_8569);
nor U9115 (N_9115,N_8636,N_8453);
nand U9116 (N_9116,N_8648,N_8401);
and U9117 (N_9117,N_8620,N_8429);
nand U9118 (N_9118,N_8754,N_8641);
nand U9119 (N_9119,N_8636,N_8458);
and U9120 (N_9120,N_8543,N_8572);
or U9121 (N_9121,N_8462,N_8607);
nand U9122 (N_9122,N_8665,N_8492);
or U9123 (N_9123,N_8691,N_8431);
xor U9124 (N_9124,N_8643,N_8461);
xnor U9125 (N_9125,N_8645,N_8721);
xor U9126 (N_9126,N_8618,N_8630);
and U9127 (N_9127,N_8733,N_8453);
and U9128 (N_9128,N_8407,N_8696);
nor U9129 (N_9129,N_8796,N_8456);
or U9130 (N_9130,N_8684,N_8632);
and U9131 (N_9131,N_8513,N_8403);
and U9132 (N_9132,N_8656,N_8766);
nand U9133 (N_9133,N_8664,N_8764);
and U9134 (N_9134,N_8475,N_8750);
nand U9135 (N_9135,N_8775,N_8566);
and U9136 (N_9136,N_8612,N_8697);
and U9137 (N_9137,N_8532,N_8671);
nand U9138 (N_9138,N_8572,N_8402);
nand U9139 (N_9139,N_8576,N_8738);
nor U9140 (N_9140,N_8735,N_8523);
nor U9141 (N_9141,N_8661,N_8797);
and U9142 (N_9142,N_8737,N_8763);
or U9143 (N_9143,N_8461,N_8535);
or U9144 (N_9144,N_8516,N_8717);
nor U9145 (N_9145,N_8668,N_8535);
nand U9146 (N_9146,N_8755,N_8630);
and U9147 (N_9147,N_8765,N_8771);
and U9148 (N_9148,N_8799,N_8716);
nand U9149 (N_9149,N_8650,N_8643);
nand U9150 (N_9150,N_8631,N_8507);
nor U9151 (N_9151,N_8770,N_8700);
xnor U9152 (N_9152,N_8502,N_8463);
and U9153 (N_9153,N_8460,N_8438);
xnor U9154 (N_9154,N_8658,N_8647);
and U9155 (N_9155,N_8630,N_8648);
xor U9156 (N_9156,N_8503,N_8708);
and U9157 (N_9157,N_8792,N_8506);
xor U9158 (N_9158,N_8778,N_8615);
nand U9159 (N_9159,N_8760,N_8778);
nor U9160 (N_9160,N_8402,N_8487);
nand U9161 (N_9161,N_8791,N_8654);
nand U9162 (N_9162,N_8771,N_8720);
or U9163 (N_9163,N_8629,N_8500);
nand U9164 (N_9164,N_8783,N_8647);
and U9165 (N_9165,N_8446,N_8672);
and U9166 (N_9166,N_8525,N_8550);
nand U9167 (N_9167,N_8586,N_8452);
and U9168 (N_9168,N_8560,N_8510);
nor U9169 (N_9169,N_8544,N_8716);
nor U9170 (N_9170,N_8625,N_8436);
and U9171 (N_9171,N_8436,N_8506);
and U9172 (N_9172,N_8709,N_8590);
or U9173 (N_9173,N_8625,N_8788);
nand U9174 (N_9174,N_8468,N_8583);
or U9175 (N_9175,N_8544,N_8758);
nand U9176 (N_9176,N_8472,N_8427);
and U9177 (N_9177,N_8482,N_8543);
or U9178 (N_9178,N_8478,N_8599);
nor U9179 (N_9179,N_8564,N_8566);
and U9180 (N_9180,N_8602,N_8459);
xor U9181 (N_9181,N_8542,N_8712);
nor U9182 (N_9182,N_8428,N_8523);
nor U9183 (N_9183,N_8421,N_8707);
xnor U9184 (N_9184,N_8443,N_8655);
nand U9185 (N_9185,N_8505,N_8713);
or U9186 (N_9186,N_8769,N_8619);
or U9187 (N_9187,N_8706,N_8435);
nor U9188 (N_9188,N_8622,N_8586);
or U9189 (N_9189,N_8423,N_8710);
or U9190 (N_9190,N_8430,N_8534);
xnor U9191 (N_9191,N_8782,N_8451);
nand U9192 (N_9192,N_8483,N_8493);
or U9193 (N_9193,N_8644,N_8740);
and U9194 (N_9194,N_8465,N_8536);
or U9195 (N_9195,N_8694,N_8568);
nor U9196 (N_9196,N_8772,N_8726);
nand U9197 (N_9197,N_8521,N_8771);
or U9198 (N_9198,N_8414,N_8610);
xor U9199 (N_9199,N_8532,N_8603);
nor U9200 (N_9200,N_8815,N_9119);
or U9201 (N_9201,N_8987,N_8816);
or U9202 (N_9202,N_9123,N_8938);
nand U9203 (N_9203,N_9001,N_8963);
xnor U9204 (N_9204,N_8923,N_8983);
and U9205 (N_9205,N_9192,N_9029);
xnor U9206 (N_9206,N_8859,N_8839);
nor U9207 (N_9207,N_9083,N_9188);
and U9208 (N_9208,N_9132,N_9103);
or U9209 (N_9209,N_9072,N_9044);
or U9210 (N_9210,N_9109,N_9085);
or U9211 (N_9211,N_8908,N_8984);
or U9212 (N_9212,N_8971,N_8933);
xor U9213 (N_9213,N_9171,N_9098);
and U9214 (N_9214,N_8862,N_9020);
xnor U9215 (N_9215,N_9035,N_8861);
xnor U9216 (N_9216,N_9059,N_8980);
xnor U9217 (N_9217,N_8865,N_8880);
nor U9218 (N_9218,N_9148,N_8823);
nor U9219 (N_9219,N_9181,N_9011);
nand U9220 (N_9220,N_8836,N_8900);
or U9221 (N_9221,N_8818,N_8927);
nand U9222 (N_9222,N_9061,N_9038);
nor U9223 (N_9223,N_9045,N_8848);
or U9224 (N_9224,N_9092,N_8896);
xnor U9225 (N_9225,N_8962,N_9015);
nor U9226 (N_9226,N_9099,N_9164);
xnor U9227 (N_9227,N_9010,N_8849);
or U9228 (N_9228,N_9151,N_9016);
nand U9229 (N_9229,N_9182,N_9195);
or U9230 (N_9230,N_9081,N_9165);
or U9231 (N_9231,N_8960,N_9024);
nor U9232 (N_9232,N_8954,N_8990);
nor U9233 (N_9233,N_9169,N_8835);
nor U9234 (N_9234,N_8926,N_8846);
xor U9235 (N_9235,N_8998,N_9189);
nor U9236 (N_9236,N_8915,N_8871);
xnor U9237 (N_9237,N_9000,N_9068);
nor U9238 (N_9238,N_8901,N_8813);
nand U9239 (N_9239,N_9037,N_8945);
or U9240 (N_9240,N_8810,N_9088);
or U9241 (N_9241,N_8904,N_9117);
xor U9242 (N_9242,N_8934,N_8910);
nor U9243 (N_9243,N_9082,N_8999);
or U9244 (N_9244,N_9086,N_9196);
and U9245 (N_9245,N_8852,N_9153);
nand U9246 (N_9246,N_9003,N_8937);
or U9247 (N_9247,N_8970,N_9198);
nor U9248 (N_9248,N_8988,N_9193);
and U9249 (N_9249,N_8883,N_9091);
xnor U9250 (N_9250,N_9071,N_8834);
and U9251 (N_9251,N_9019,N_8845);
or U9252 (N_9252,N_9107,N_9175);
or U9253 (N_9253,N_9112,N_8966);
xnor U9254 (N_9254,N_8866,N_8858);
xor U9255 (N_9255,N_8891,N_9187);
and U9256 (N_9256,N_8958,N_9069);
nor U9257 (N_9257,N_8807,N_9194);
or U9258 (N_9258,N_9154,N_9040);
xnor U9259 (N_9259,N_9130,N_8826);
or U9260 (N_9260,N_8832,N_9073);
and U9261 (N_9261,N_8869,N_8916);
nor U9262 (N_9262,N_8804,N_9190);
nand U9263 (N_9263,N_9006,N_8847);
or U9264 (N_9264,N_9066,N_8913);
xnor U9265 (N_9265,N_9070,N_9147);
xor U9266 (N_9266,N_8867,N_8905);
or U9267 (N_9267,N_8973,N_8802);
xor U9268 (N_9268,N_8975,N_9026);
nand U9269 (N_9269,N_8894,N_8922);
or U9270 (N_9270,N_8912,N_9178);
xor U9271 (N_9271,N_9022,N_8873);
and U9272 (N_9272,N_9105,N_8886);
xnor U9273 (N_9273,N_8967,N_8976);
xnor U9274 (N_9274,N_9067,N_8814);
or U9275 (N_9275,N_8947,N_8997);
nand U9276 (N_9276,N_8877,N_9111);
nor U9277 (N_9277,N_9156,N_9186);
nand U9278 (N_9278,N_8870,N_9143);
nor U9279 (N_9279,N_9096,N_9179);
and U9280 (N_9280,N_8925,N_9118);
xnor U9281 (N_9281,N_8949,N_8931);
nand U9282 (N_9282,N_9155,N_9162);
xnor U9283 (N_9283,N_9173,N_9050);
nand U9284 (N_9284,N_8838,N_8981);
nor U9285 (N_9285,N_8892,N_8898);
and U9286 (N_9286,N_9184,N_8935);
xor U9287 (N_9287,N_8932,N_9036);
or U9288 (N_9288,N_8860,N_8879);
xor U9289 (N_9289,N_8830,N_9102);
nor U9290 (N_9290,N_8985,N_8827);
nand U9291 (N_9291,N_9149,N_8924);
and U9292 (N_9292,N_8889,N_9141);
nor U9293 (N_9293,N_9077,N_9057);
xnor U9294 (N_9294,N_8993,N_8895);
nand U9295 (N_9295,N_9052,N_8864);
or U9296 (N_9296,N_9089,N_9018);
or U9297 (N_9297,N_8897,N_9025);
nand U9298 (N_9298,N_9041,N_9104);
or U9299 (N_9299,N_9058,N_9163);
nand U9300 (N_9300,N_8822,N_9176);
xnor U9301 (N_9301,N_9028,N_9063);
nand U9302 (N_9302,N_9122,N_9060);
or U9303 (N_9303,N_9116,N_8868);
and U9304 (N_9304,N_9080,N_9007);
nand U9305 (N_9305,N_8805,N_9013);
and U9306 (N_9306,N_9168,N_9177);
or U9307 (N_9307,N_8817,N_9101);
xnor U9308 (N_9308,N_8946,N_8831);
or U9309 (N_9309,N_9146,N_8928);
nand U9310 (N_9310,N_8909,N_9160);
or U9311 (N_9311,N_8801,N_9076);
and U9312 (N_9312,N_9124,N_8914);
or U9313 (N_9313,N_8800,N_9157);
or U9314 (N_9314,N_9197,N_8874);
nand U9315 (N_9315,N_8930,N_8875);
nor U9316 (N_9316,N_8977,N_9137);
nor U9317 (N_9317,N_8829,N_8863);
xnor U9318 (N_9318,N_8943,N_9095);
nand U9319 (N_9319,N_8821,N_9114);
or U9320 (N_9320,N_8942,N_9199);
or U9321 (N_9321,N_9185,N_9051);
and U9322 (N_9322,N_8828,N_9043);
nand U9323 (N_9323,N_8899,N_8837);
or U9324 (N_9324,N_9002,N_9139);
nor U9325 (N_9325,N_8906,N_8979);
xor U9326 (N_9326,N_9134,N_9138);
or U9327 (N_9327,N_8940,N_8978);
or U9328 (N_9328,N_9031,N_9140);
xor U9329 (N_9329,N_8887,N_9133);
or U9330 (N_9330,N_8974,N_8878);
nor U9331 (N_9331,N_8882,N_9167);
nand U9332 (N_9332,N_9027,N_9030);
or U9333 (N_9333,N_8918,N_9097);
and U9334 (N_9334,N_9090,N_8808);
nand U9335 (N_9335,N_8920,N_8986);
and U9336 (N_9336,N_9056,N_8811);
nor U9337 (N_9337,N_9023,N_9150);
nor U9338 (N_9338,N_9014,N_8996);
and U9339 (N_9339,N_8855,N_8995);
xor U9340 (N_9340,N_9049,N_9144);
nand U9341 (N_9341,N_8941,N_8956);
xnor U9342 (N_9342,N_9048,N_9159);
xor U9343 (N_9343,N_8969,N_9180);
nor U9344 (N_9344,N_9170,N_9034);
and U9345 (N_9345,N_9172,N_8825);
nand U9346 (N_9346,N_9074,N_8957);
and U9347 (N_9347,N_9062,N_9127);
or U9348 (N_9348,N_8992,N_8885);
xnor U9349 (N_9349,N_8853,N_9166);
xnor U9350 (N_9350,N_8840,N_8953);
and U9351 (N_9351,N_8812,N_8921);
and U9352 (N_9352,N_8952,N_8917);
and U9353 (N_9353,N_8890,N_9053);
or U9354 (N_9354,N_9183,N_8948);
or U9355 (N_9355,N_8893,N_8833);
nor U9356 (N_9356,N_8955,N_8944);
nand U9357 (N_9357,N_8907,N_8959);
and U9358 (N_9358,N_9129,N_9087);
nor U9359 (N_9359,N_8857,N_8911);
and U9360 (N_9360,N_9131,N_8972);
xor U9361 (N_9361,N_8851,N_8876);
nand U9362 (N_9362,N_9110,N_9106);
and U9363 (N_9363,N_9012,N_9115);
xor U9364 (N_9364,N_9017,N_8850);
and U9365 (N_9365,N_9046,N_8961);
or U9366 (N_9366,N_8803,N_8929);
nor U9367 (N_9367,N_8844,N_9064);
xor U9368 (N_9368,N_9142,N_9055);
and U9369 (N_9369,N_8991,N_8824);
xnor U9370 (N_9370,N_9125,N_9120);
and U9371 (N_9371,N_8809,N_8881);
and U9372 (N_9372,N_8951,N_9004);
and U9373 (N_9373,N_9039,N_9113);
and U9374 (N_9374,N_9005,N_8854);
or U9375 (N_9375,N_8842,N_9075);
and U9376 (N_9376,N_8964,N_9084);
or U9377 (N_9377,N_8965,N_8903);
xor U9378 (N_9378,N_8820,N_9128);
nand U9379 (N_9379,N_8819,N_9054);
nand U9380 (N_9380,N_9174,N_9126);
nand U9381 (N_9381,N_9079,N_9158);
xor U9382 (N_9382,N_9094,N_8884);
nand U9383 (N_9383,N_9065,N_9108);
or U9384 (N_9384,N_8989,N_9136);
nand U9385 (N_9385,N_9032,N_9009);
nand U9386 (N_9386,N_9100,N_8939);
xnor U9387 (N_9387,N_9135,N_8888);
nor U9388 (N_9388,N_9008,N_9093);
nor U9389 (N_9389,N_9033,N_9121);
and U9390 (N_9390,N_8950,N_8968);
nand U9391 (N_9391,N_8919,N_9078);
nand U9392 (N_9392,N_9161,N_9047);
and U9393 (N_9393,N_9042,N_8841);
nand U9394 (N_9394,N_8936,N_8843);
xor U9395 (N_9395,N_9021,N_8806);
or U9396 (N_9396,N_9191,N_9145);
and U9397 (N_9397,N_8902,N_8872);
nor U9398 (N_9398,N_8856,N_9152);
nand U9399 (N_9399,N_8982,N_8994);
nor U9400 (N_9400,N_9065,N_9198);
or U9401 (N_9401,N_8862,N_9100);
or U9402 (N_9402,N_8811,N_9121);
xor U9403 (N_9403,N_9136,N_8981);
and U9404 (N_9404,N_9089,N_9167);
nand U9405 (N_9405,N_8839,N_9197);
or U9406 (N_9406,N_9180,N_9146);
or U9407 (N_9407,N_8813,N_8903);
or U9408 (N_9408,N_9154,N_8873);
xor U9409 (N_9409,N_8831,N_9144);
nand U9410 (N_9410,N_8940,N_8986);
xnor U9411 (N_9411,N_8804,N_9159);
nand U9412 (N_9412,N_8914,N_8862);
nor U9413 (N_9413,N_9115,N_8909);
or U9414 (N_9414,N_8984,N_8980);
nor U9415 (N_9415,N_9198,N_8955);
xnor U9416 (N_9416,N_8853,N_8979);
and U9417 (N_9417,N_9125,N_9084);
nor U9418 (N_9418,N_9115,N_8977);
xnor U9419 (N_9419,N_8819,N_8829);
xor U9420 (N_9420,N_9074,N_9160);
nor U9421 (N_9421,N_8909,N_9080);
xor U9422 (N_9422,N_8800,N_9000);
nand U9423 (N_9423,N_8884,N_9060);
xnor U9424 (N_9424,N_8920,N_8821);
nand U9425 (N_9425,N_9121,N_9125);
xnor U9426 (N_9426,N_8804,N_9095);
xor U9427 (N_9427,N_9188,N_8975);
or U9428 (N_9428,N_9135,N_9185);
and U9429 (N_9429,N_8999,N_8882);
nand U9430 (N_9430,N_8880,N_9116);
xnor U9431 (N_9431,N_9013,N_9019);
or U9432 (N_9432,N_8906,N_8899);
xor U9433 (N_9433,N_8962,N_8908);
nand U9434 (N_9434,N_8818,N_8832);
and U9435 (N_9435,N_8868,N_8999);
xnor U9436 (N_9436,N_8911,N_9039);
nand U9437 (N_9437,N_8813,N_9034);
or U9438 (N_9438,N_8876,N_9046);
nand U9439 (N_9439,N_9141,N_9057);
xor U9440 (N_9440,N_8931,N_9190);
nand U9441 (N_9441,N_9120,N_9020);
and U9442 (N_9442,N_9153,N_9046);
nor U9443 (N_9443,N_9062,N_8884);
and U9444 (N_9444,N_8810,N_9119);
nor U9445 (N_9445,N_9170,N_9123);
and U9446 (N_9446,N_9144,N_8892);
nand U9447 (N_9447,N_9197,N_9055);
nor U9448 (N_9448,N_8836,N_8953);
or U9449 (N_9449,N_8879,N_9014);
and U9450 (N_9450,N_8880,N_8855);
nor U9451 (N_9451,N_8851,N_9084);
or U9452 (N_9452,N_9039,N_9130);
xor U9453 (N_9453,N_8930,N_8998);
or U9454 (N_9454,N_9082,N_8978);
nand U9455 (N_9455,N_9185,N_8893);
nor U9456 (N_9456,N_8981,N_8942);
or U9457 (N_9457,N_8906,N_8891);
nand U9458 (N_9458,N_8862,N_9094);
or U9459 (N_9459,N_9062,N_9051);
and U9460 (N_9460,N_8842,N_8976);
and U9461 (N_9461,N_9062,N_9008);
nand U9462 (N_9462,N_8948,N_8882);
and U9463 (N_9463,N_8967,N_9111);
xor U9464 (N_9464,N_8834,N_8820);
and U9465 (N_9465,N_8849,N_9114);
or U9466 (N_9466,N_9076,N_9013);
xor U9467 (N_9467,N_9139,N_9061);
nor U9468 (N_9468,N_8844,N_8934);
and U9469 (N_9469,N_8825,N_9077);
or U9470 (N_9470,N_8806,N_9058);
nor U9471 (N_9471,N_8854,N_8979);
and U9472 (N_9472,N_9173,N_8819);
and U9473 (N_9473,N_9181,N_8959);
nor U9474 (N_9474,N_9183,N_9072);
nor U9475 (N_9475,N_9173,N_9067);
and U9476 (N_9476,N_9135,N_8988);
or U9477 (N_9477,N_9000,N_8813);
nand U9478 (N_9478,N_9181,N_8982);
nor U9479 (N_9479,N_9095,N_8923);
nand U9480 (N_9480,N_9168,N_8993);
nor U9481 (N_9481,N_9179,N_9095);
or U9482 (N_9482,N_9166,N_9077);
and U9483 (N_9483,N_9109,N_9045);
or U9484 (N_9484,N_8820,N_9099);
and U9485 (N_9485,N_9105,N_9110);
nand U9486 (N_9486,N_8919,N_8912);
xnor U9487 (N_9487,N_8921,N_9031);
xnor U9488 (N_9488,N_8848,N_8847);
nor U9489 (N_9489,N_8967,N_9170);
nor U9490 (N_9490,N_9155,N_9159);
and U9491 (N_9491,N_8837,N_8949);
or U9492 (N_9492,N_9190,N_8944);
xor U9493 (N_9493,N_8870,N_8806);
or U9494 (N_9494,N_8909,N_9082);
nand U9495 (N_9495,N_8924,N_8939);
nand U9496 (N_9496,N_9099,N_8990);
nand U9497 (N_9497,N_8931,N_8925);
or U9498 (N_9498,N_8993,N_8873);
nand U9499 (N_9499,N_9108,N_9115);
nand U9500 (N_9500,N_9009,N_9061);
and U9501 (N_9501,N_9030,N_8805);
nor U9502 (N_9502,N_8946,N_9047);
xnor U9503 (N_9503,N_9080,N_9140);
nor U9504 (N_9504,N_9099,N_9177);
and U9505 (N_9505,N_8865,N_8807);
or U9506 (N_9506,N_9071,N_8828);
nor U9507 (N_9507,N_9065,N_8865);
nand U9508 (N_9508,N_9111,N_8960);
xor U9509 (N_9509,N_8961,N_9035);
and U9510 (N_9510,N_9010,N_9136);
nor U9511 (N_9511,N_8856,N_9198);
nand U9512 (N_9512,N_9029,N_8889);
or U9513 (N_9513,N_9170,N_8848);
and U9514 (N_9514,N_8850,N_8876);
or U9515 (N_9515,N_8902,N_8897);
and U9516 (N_9516,N_9186,N_9113);
xnor U9517 (N_9517,N_9171,N_9097);
nand U9518 (N_9518,N_8932,N_9163);
nor U9519 (N_9519,N_9085,N_8938);
or U9520 (N_9520,N_8966,N_9076);
or U9521 (N_9521,N_8874,N_8809);
nor U9522 (N_9522,N_8967,N_9137);
or U9523 (N_9523,N_9160,N_9128);
xor U9524 (N_9524,N_8884,N_9033);
xor U9525 (N_9525,N_9065,N_9005);
or U9526 (N_9526,N_9140,N_8816);
nand U9527 (N_9527,N_8800,N_8804);
nand U9528 (N_9528,N_8816,N_8968);
or U9529 (N_9529,N_9029,N_8990);
or U9530 (N_9530,N_9035,N_9181);
nor U9531 (N_9531,N_8807,N_9067);
or U9532 (N_9532,N_9077,N_9034);
or U9533 (N_9533,N_9123,N_8986);
nand U9534 (N_9534,N_8801,N_8930);
nor U9535 (N_9535,N_9097,N_9083);
nor U9536 (N_9536,N_8914,N_9019);
nand U9537 (N_9537,N_9052,N_9189);
nor U9538 (N_9538,N_9151,N_9012);
or U9539 (N_9539,N_8914,N_8802);
nand U9540 (N_9540,N_8849,N_8935);
and U9541 (N_9541,N_8906,N_9001);
xnor U9542 (N_9542,N_9090,N_8986);
and U9543 (N_9543,N_8814,N_8820);
and U9544 (N_9544,N_8997,N_9184);
nor U9545 (N_9545,N_9183,N_8811);
or U9546 (N_9546,N_8883,N_8826);
nor U9547 (N_9547,N_8811,N_8904);
nand U9548 (N_9548,N_8916,N_9190);
nand U9549 (N_9549,N_8842,N_8871);
nand U9550 (N_9550,N_9127,N_9135);
or U9551 (N_9551,N_8900,N_9131);
or U9552 (N_9552,N_8903,N_9190);
or U9553 (N_9553,N_9012,N_8958);
and U9554 (N_9554,N_8970,N_9165);
nor U9555 (N_9555,N_9123,N_8968);
nor U9556 (N_9556,N_8885,N_8923);
and U9557 (N_9557,N_8911,N_9020);
or U9558 (N_9558,N_8852,N_8814);
and U9559 (N_9559,N_8802,N_8872);
nand U9560 (N_9560,N_8875,N_9114);
and U9561 (N_9561,N_8895,N_8809);
nor U9562 (N_9562,N_9193,N_8860);
and U9563 (N_9563,N_9055,N_9065);
nor U9564 (N_9564,N_8907,N_9061);
or U9565 (N_9565,N_8850,N_9167);
xor U9566 (N_9566,N_8820,N_8888);
and U9567 (N_9567,N_9084,N_8984);
xnor U9568 (N_9568,N_8868,N_9004);
and U9569 (N_9569,N_8982,N_8836);
nor U9570 (N_9570,N_9094,N_8928);
nor U9571 (N_9571,N_8911,N_9017);
xnor U9572 (N_9572,N_9122,N_9046);
nand U9573 (N_9573,N_9193,N_8925);
or U9574 (N_9574,N_8911,N_9058);
xnor U9575 (N_9575,N_8979,N_8987);
nand U9576 (N_9576,N_8984,N_9127);
nor U9577 (N_9577,N_9078,N_8926);
or U9578 (N_9578,N_9156,N_8942);
nand U9579 (N_9579,N_8827,N_8800);
nand U9580 (N_9580,N_8869,N_8940);
nor U9581 (N_9581,N_8846,N_9118);
xor U9582 (N_9582,N_8897,N_9133);
and U9583 (N_9583,N_9145,N_9114);
and U9584 (N_9584,N_9129,N_8996);
and U9585 (N_9585,N_9013,N_9066);
xor U9586 (N_9586,N_8980,N_9005);
or U9587 (N_9587,N_9040,N_9182);
and U9588 (N_9588,N_8872,N_8864);
xnor U9589 (N_9589,N_8821,N_9136);
xnor U9590 (N_9590,N_8851,N_8990);
xor U9591 (N_9591,N_8917,N_8868);
nor U9592 (N_9592,N_8986,N_9082);
or U9593 (N_9593,N_8957,N_8988);
or U9594 (N_9594,N_8928,N_9093);
and U9595 (N_9595,N_8843,N_8924);
or U9596 (N_9596,N_8987,N_8867);
nor U9597 (N_9597,N_8846,N_8828);
xnor U9598 (N_9598,N_8874,N_8855);
nor U9599 (N_9599,N_8934,N_8971);
or U9600 (N_9600,N_9450,N_9528);
xnor U9601 (N_9601,N_9505,N_9326);
nor U9602 (N_9602,N_9423,N_9487);
and U9603 (N_9603,N_9314,N_9271);
xnor U9604 (N_9604,N_9529,N_9418);
or U9605 (N_9605,N_9325,N_9376);
nor U9606 (N_9606,N_9303,N_9208);
xnor U9607 (N_9607,N_9552,N_9293);
or U9608 (N_9608,N_9512,N_9234);
and U9609 (N_9609,N_9232,N_9224);
and U9610 (N_9610,N_9467,N_9394);
and U9611 (N_9611,N_9367,N_9488);
xor U9612 (N_9612,N_9546,N_9279);
nor U9613 (N_9613,N_9395,N_9273);
or U9614 (N_9614,N_9490,N_9594);
or U9615 (N_9615,N_9245,N_9496);
and U9616 (N_9616,N_9346,N_9242);
nor U9617 (N_9617,N_9441,N_9448);
xor U9618 (N_9618,N_9350,N_9391);
nand U9619 (N_9619,N_9447,N_9432);
nor U9620 (N_9620,N_9520,N_9433);
xnor U9621 (N_9621,N_9577,N_9553);
nor U9622 (N_9622,N_9464,N_9525);
nor U9623 (N_9623,N_9304,N_9492);
nor U9624 (N_9624,N_9579,N_9456);
xnor U9625 (N_9625,N_9408,N_9468);
xnor U9626 (N_9626,N_9352,N_9584);
nand U9627 (N_9627,N_9483,N_9309);
xor U9628 (N_9628,N_9585,N_9244);
and U9629 (N_9629,N_9272,N_9473);
nand U9630 (N_9630,N_9207,N_9205);
nor U9631 (N_9631,N_9401,N_9516);
nand U9632 (N_9632,N_9549,N_9344);
xor U9633 (N_9633,N_9562,N_9491);
xnor U9634 (N_9634,N_9231,N_9316);
xor U9635 (N_9635,N_9550,N_9533);
xor U9636 (N_9636,N_9308,N_9489);
xor U9637 (N_9637,N_9377,N_9247);
or U9638 (N_9638,N_9416,N_9343);
nor U9639 (N_9639,N_9386,N_9503);
xor U9640 (N_9640,N_9479,N_9311);
or U9641 (N_9641,N_9385,N_9522);
nand U9642 (N_9642,N_9331,N_9354);
xor U9643 (N_9643,N_9502,N_9313);
xnor U9644 (N_9644,N_9268,N_9518);
nand U9645 (N_9645,N_9220,N_9364);
xor U9646 (N_9646,N_9587,N_9335);
and U9647 (N_9647,N_9438,N_9451);
and U9648 (N_9648,N_9414,N_9428);
xnor U9649 (N_9649,N_9222,N_9319);
and U9650 (N_9650,N_9590,N_9274);
or U9651 (N_9651,N_9390,N_9499);
or U9652 (N_9652,N_9534,N_9286);
xnor U9653 (N_9653,N_9466,N_9586);
nand U9654 (N_9654,N_9332,N_9403);
and U9655 (N_9655,N_9453,N_9212);
or U9656 (N_9656,N_9383,N_9446);
or U9657 (N_9657,N_9570,N_9320);
xor U9658 (N_9658,N_9591,N_9569);
or U9659 (N_9659,N_9480,N_9530);
and U9660 (N_9660,N_9258,N_9485);
or U9661 (N_9661,N_9227,N_9351);
nand U9662 (N_9662,N_9458,N_9201);
xor U9663 (N_9663,N_9327,N_9238);
or U9664 (N_9664,N_9397,N_9353);
and U9665 (N_9665,N_9437,N_9495);
and U9666 (N_9666,N_9270,N_9300);
and U9667 (N_9667,N_9519,N_9429);
nand U9668 (N_9668,N_9475,N_9555);
or U9669 (N_9669,N_9213,N_9405);
xor U9670 (N_9670,N_9444,N_9223);
and U9671 (N_9671,N_9547,N_9366);
or U9672 (N_9672,N_9581,N_9260);
nor U9673 (N_9673,N_9578,N_9471);
nand U9674 (N_9674,N_9336,N_9424);
or U9675 (N_9675,N_9399,N_9506);
or U9676 (N_9676,N_9239,N_9233);
xnor U9677 (N_9677,N_9393,N_9589);
nand U9678 (N_9678,N_9531,N_9426);
xnor U9679 (N_9679,N_9265,N_9412);
xor U9680 (N_9680,N_9257,N_9306);
or U9681 (N_9681,N_9415,N_9497);
or U9682 (N_9682,N_9215,N_9461);
xnor U9683 (N_9683,N_9371,N_9538);
nor U9684 (N_9684,N_9463,N_9482);
nor U9685 (N_9685,N_9543,N_9430);
xnor U9686 (N_9686,N_9210,N_9524);
and U9687 (N_9687,N_9413,N_9375);
nor U9688 (N_9688,N_9254,N_9246);
nor U9689 (N_9689,N_9278,N_9540);
xnor U9690 (N_9690,N_9301,N_9334);
nand U9691 (N_9691,N_9501,N_9435);
nor U9692 (N_9692,N_9409,N_9442);
or U9693 (N_9693,N_9249,N_9598);
or U9694 (N_9694,N_9417,N_9348);
and U9695 (N_9695,N_9342,N_9443);
or U9696 (N_9696,N_9545,N_9514);
or U9697 (N_9697,N_9203,N_9284);
nand U9698 (N_9698,N_9544,N_9200);
or U9699 (N_9699,N_9291,N_9240);
xor U9700 (N_9700,N_9370,N_9330);
or U9701 (N_9701,N_9536,N_9276);
nand U9702 (N_9702,N_9400,N_9361);
or U9703 (N_9703,N_9478,N_9288);
xnor U9704 (N_9704,N_9329,N_9362);
nand U9705 (N_9705,N_9572,N_9554);
and U9706 (N_9706,N_9472,N_9476);
nand U9707 (N_9707,N_9431,N_9532);
and U9708 (N_9708,N_9388,N_9504);
or U9709 (N_9709,N_9228,N_9216);
nand U9710 (N_9710,N_9420,N_9369);
or U9711 (N_9711,N_9597,N_9317);
nor U9712 (N_9712,N_9527,N_9449);
xnor U9713 (N_9713,N_9481,N_9323);
nor U9714 (N_9714,N_9292,N_9470);
nand U9715 (N_9715,N_9324,N_9551);
and U9716 (N_9716,N_9455,N_9445);
or U9717 (N_9717,N_9297,N_9262);
xnor U9718 (N_9718,N_9379,N_9382);
nor U9719 (N_9719,N_9407,N_9287);
nor U9720 (N_9720,N_9237,N_9425);
nor U9721 (N_9721,N_9474,N_9338);
and U9722 (N_9722,N_9592,N_9381);
or U9723 (N_9723,N_9460,N_9267);
nor U9724 (N_9724,N_9225,N_9290);
nor U9725 (N_9725,N_9202,N_9571);
xnor U9726 (N_9726,N_9241,N_9368);
nand U9727 (N_9727,N_9500,N_9358);
xor U9728 (N_9728,N_9298,N_9515);
xor U9729 (N_9729,N_9517,N_9365);
nand U9730 (N_9730,N_9498,N_9347);
xor U9731 (N_9731,N_9266,N_9363);
nand U9732 (N_9732,N_9263,N_9484);
nor U9733 (N_9733,N_9356,N_9218);
nor U9734 (N_9734,N_9567,N_9560);
or U9735 (N_9735,N_9387,N_9582);
xnor U9736 (N_9736,N_9462,N_9235);
or U9737 (N_9737,N_9411,N_9384);
xnor U9738 (N_9738,N_9339,N_9250);
and U9739 (N_9739,N_9389,N_9565);
nor U9740 (N_9740,N_9539,N_9542);
nand U9741 (N_9741,N_9219,N_9568);
xnor U9742 (N_9742,N_9322,N_9226);
and U9743 (N_9743,N_9564,N_9236);
nand U9744 (N_9744,N_9340,N_9526);
nor U9745 (N_9745,N_9333,N_9596);
and U9746 (N_9746,N_9493,N_9294);
xnor U9747 (N_9747,N_9573,N_9277);
xnor U9748 (N_9748,N_9422,N_9477);
or U9749 (N_9749,N_9204,N_9452);
or U9750 (N_9750,N_9580,N_9427);
and U9751 (N_9751,N_9373,N_9217);
xnor U9752 (N_9752,N_9345,N_9251);
nand U9753 (N_9753,N_9558,N_9588);
nor U9754 (N_9754,N_9599,N_9253);
nor U9755 (N_9755,N_9380,N_9209);
and U9756 (N_9756,N_9289,N_9230);
nand U9757 (N_9757,N_9341,N_9318);
or U9758 (N_9758,N_9583,N_9252);
or U9759 (N_9759,N_9229,N_9372);
xnor U9760 (N_9760,N_9282,N_9440);
nand U9761 (N_9761,N_9259,N_9563);
or U9762 (N_9762,N_9315,N_9511);
xor U9763 (N_9763,N_9256,N_9402);
nor U9764 (N_9764,N_9269,N_9439);
xor U9765 (N_9765,N_9593,N_9378);
and U9766 (N_9766,N_9307,N_9494);
nand U9767 (N_9767,N_9537,N_9295);
xor U9768 (N_9768,N_9310,N_9321);
and U9769 (N_9769,N_9457,N_9404);
nand U9770 (N_9770,N_9357,N_9296);
nor U9771 (N_9771,N_9328,N_9283);
and U9772 (N_9772,N_9264,N_9285);
xnor U9773 (N_9773,N_9299,N_9548);
nor U9774 (N_9774,N_9576,N_9281);
nor U9775 (N_9775,N_9398,N_9566);
nand U9776 (N_9776,N_9434,N_9459);
nand U9777 (N_9777,N_9374,N_9535);
nor U9778 (N_9778,N_9243,N_9561);
and U9779 (N_9779,N_9510,N_9465);
nand U9780 (N_9780,N_9454,N_9221);
nor U9781 (N_9781,N_9406,N_9513);
nand U9782 (N_9782,N_9211,N_9556);
nand U9783 (N_9783,N_9421,N_9248);
and U9784 (N_9784,N_9523,N_9302);
xor U9785 (N_9785,N_9559,N_9575);
or U9786 (N_9786,N_9255,N_9541);
and U9787 (N_9787,N_9521,N_9280);
or U9788 (N_9788,N_9410,N_9275);
nand U9789 (N_9789,N_9312,N_9214);
xor U9790 (N_9790,N_9508,N_9436);
or U9791 (N_9791,N_9509,N_9206);
or U9792 (N_9792,N_9469,N_9595);
nor U9793 (N_9793,N_9396,N_9337);
nor U9794 (N_9794,N_9507,N_9392);
or U9795 (N_9795,N_9349,N_9305);
xor U9796 (N_9796,N_9261,N_9557);
xnor U9797 (N_9797,N_9359,N_9486);
xnor U9798 (N_9798,N_9574,N_9419);
and U9799 (N_9799,N_9355,N_9360);
and U9800 (N_9800,N_9323,N_9531);
nor U9801 (N_9801,N_9452,N_9315);
nand U9802 (N_9802,N_9333,N_9358);
nor U9803 (N_9803,N_9564,N_9466);
and U9804 (N_9804,N_9216,N_9521);
nor U9805 (N_9805,N_9236,N_9457);
nor U9806 (N_9806,N_9570,N_9556);
and U9807 (N_9807,N_9577,N_9410);
xnor U9808 (N_9808,N_9485,N_9400);
or U9809 (N_9809,N_9551,N_9570);
and U9810 (N_9810,N_9342,N_9438);
or U9811 (N_9811,N_9425,N_9437);
or U9812 (N_9812,N_9312,N_9454);
or U9813 (N_9813,N_9326,N_9592);
or U9814 (N_9814,N_9409,N_9592);
or U9815 (N_9815,N_9474,N_9295);
or U9816 (N_9816,N_9244,N_9446);
nor U9817 (N_9817,N_9496,N_9422);
nand U9818 (N_9818,N_9310,N_9323);
nor U9819 (N_9819,N_9386,N_9228);
and U9820 (N_9820,N_9420,N_9288);
or U9821 (N_9821,N_9474,N_9545);
and U9822 (N_9822,N_9458,N_9467);
xnor U9823 (N_9823,N_9520,N_9242);
xor U9824 (N_9824,N_9366,N_9292);
nor U9825 (N_9825,N_9313,N_9252);
nand U9826 (N_9826,N_9389,N_9593);
or U9827 (N_9827,N_9303,N_9394);
xor U9828 (N_9828,N_9239,N_9599);
nand U9829 (N_9829,N_9200,N_9404);
nand U9830 (N_9830,N_9212,N_9247);
nor U9831 (N_9831,N_9381,N_9253);
and U9832 (N_9832,N_9389,N_9235);
or U9833 (N_9833,N_9461,N_9378);
xor U9834 (N_9834,N_9520,N_9574);
xnor U9835 (N_9835,N_9583,N_9434);
and U9836 (N_9836,N_9453,N_9268);
or U9837 (N_9837,N_9357,N_9316);
nor U9838 (N_9838,N_9324,N_9472);
and U9839 (N_9839,N_9527,N_9447);
nor U9840 (N_9840,N_9580,N_9235);
xnor U9841 (N_9841,N_9213,N_9283);
or U9842 (N_9842,N_9267,N_9289);
xor U9843 (N_9843,N_9305,N_9386);
and U9844 (N_9844,N_9251,N_9249);
and U9845 (N_9845,N_9212,N_9565);
and U9846 (N_9846,N_9375,N_9336);
or U9847 (N_9847,N_9256,N_9501);
or U9848 (N_9848,N_9546,N_9438);
and U9849 (N_9849,N_9345,N_9436);
nor U9850 (N_9850,N_9501,N_9318);
xor U9851 (N_9851,N_9339,N_9592);
or U9852 (N_9852,N_9339,N_9480);
nand U9853 (N_9853,N_9230,N_9257);
nor U9854 (N_9854,N_9378,N_9516);
and U9855 (N_9855,N_9495,N_9200);
nand U9856 (N_9856,N_9443,N_9561);
or U9857 (N_9857,N_9333,N_9376);
xor U9858 (N_9858,N_9449,N_9537);
nand U9859 (N_9859,N_9560,N_9222);
nor U9860 (N_9860,N_9469,N_9507);
xor U9861 (N_9861,N_9324,N_9467);
and U9862 (N_9862,N_9513,N_9232);
xnor U9863 (N_9863,N_9587,N_9361);
nand U9864 (N_9864,N_9305,N_9358);
nor U9865 (N_9865,N_9451,N_9355);
nor U9866 (N_9866,N_9262,N_9211);
xnor U9867 (N_9867,N_9544,N_9490);
xnor U9868 (N_9868,N_9437,N_9573);
nand U9869 (N_9869,N_9345,N_9567);
xor U9870 (N_9870,N_9315,N_9563);
or U9871 (N_9871,N_9212,N_9402);
xnor U9872 (N_9872,N_9465,N_9224);
nor U9873 (N_9873,N_9523,N_9388);
nor U9874 (N_9874,N_9375,N_9215);
or U9875 (N_9875,N_9272,N_9437);
xor U9876 (N_9876,N_9594,N_9439);
and U9877 (N_9877,N_9328,N_9597);
nand U9878 (N_9878,N_9506,N_9280);
nor U9879 (N_9879,N_9594,N_9263);
or U9880 (N_9880,N_9283,N_9528);
nand U9881 (N_9881,N_9407,N_9325);
nand U9882 (N_9882,N_9284,N_9391);
or U9883 (N_9883,N_9432,N_9439);
nand U9884 (N_9884,N_9398,N_9281);
and U9885 (N_9885,N_9376,N_9462);
xnor U9886 (N_9886,N_9272,N_9517);
or U9887 (N_9887,N_9357,N_9465);
nor U9888 (N_9888,N_9363,N_9350);
and U9889 (N_9889,N_9570,N_9591);
nor U9890 (N_9890,N_9584,N_9258);
nor U9891 (N_9891,N_9516,N_9531);
nand U9892 (N_9892,N_9299,N_9401);
and U9893 (N_9893,N_9534,N_9271);
xor U9894 (N_9894,N_9321,N_9294);
and U9895 (N_9895,N_9317,N_9461);
xor U9896 (N_9896,N_9291,N_9567);
and U9897 (N_9897,N_9478,N_9558);
nand U9898 (N_9898,N_9245,N_9543);
xnor U9899 (N_9899,N_9586,N_9266);
nand U9900 (N_9900,N_9320,N_9256);
or U9901 (N_9901,N_9232,N_9218);
xnor U9902 (N_9902,N_9303,N_9393);
or U9903 (N_9903,N_9285,N_9441);
and U9904 (N_9904,N_9343,N_9279);
xnor U9905 (N_9905,N_9539,N_9577);
nor U9906 (N_9906,N_9453,N_9420);
nand U9907 (N_9907,N_9215,N_9526);
nor U9908 (N_9908,N_9486,N_9411);
xnor U9909 (N_9909,N_9256,N_9539);
and U9910 (N_9910,N_9265,N_9406);
or U9911 (N_9911,N_9311,N_9267);
and U9912 (N_9912,N_9331,N_9337);
nor U9913 (N_9913,N_9493,N_9374);
nor U9914 (N_9914,N_9582,N_9416);
nor U9915 (N_9915,N_9599,N_9353);
nand U9916 (N_9916,N_9468,N_9518);
xor U9917 (N_9917,N_9274,N_9305);
and U9918 (N_9918,N_9336,N_9257);
xnor U9919 (N_9919,N_9320,N_9418);
xor U9920 (N_9920,N_9334,N_9352);
nor U9921 (N_9921,N_9523,N_9389);
and U9922 (N_9922,N_9314,N_9474);
xnor U9923 (N_9923,N_9300,N_9388);
nor U9924 (N_9924,N_9451,N_9228);
or U9925 (N_9925,N_9355,N_9486);
nor U9926 (N_9926,N_9457,N_9233);
or U9927 (N_9927,N_9552,N_9588);
or U9928 (N_9928,N_9401,N_9333);
or U9929 (N_9929,N_9415,N_9349);
nand U9930 (N_9930,N_9572,N_9239);
nor U9931 (N_9931,N_9455,N_9366);
nand U9932 (N_9932,N_9551,N_9520);
nand U9933 (N_9933,N_9554,N_9226);
and U9934 (N_9934,N_9458,N_9373);
and U9935 (N_9935,N_9418,N_9257);
and U9936 (N_9936,N_9423,N_9558);
xor U9937 (N_9937,N_9366,N_9561);
and U9938 (N_9938,N_9361,N_9423);
xor U9939 (N_9939,N_9205,N_9242);
and U9940 (N_9940,N_9256,N_9210);
or U9941 (N_9941,N_9444,N_9525);
nand U9942 (N_9942,N_9275,N_9521);
xor U9943 (N_9943,N_9289,N_9385);
or U9944 (N_9944,N_9356,N_9475);
nor U9945 (N_9945,N_9458,N_9597);
nor U9946 (N_9946,N_9471,N_9257);
nand U9947 (N_9947,N_9438,N_9539);
or U9948 (N_9948,N_9455,N_9212);
nand U9949 (N_9949,N_9522,N_9369);
or U9950 (N_9950,N_9596,N_9578);
and U9951 (N_9951,N_9297,N_9495);
or U9952 (N_9952,N_9382,N_9210);
xor U9953 (N_9953,N_9395,N_9254);
and U9954 (N_9954,N_9588,N_9575);
nand U9955 (N_9955,N_9381,N_9282);
nand U9956 (N_9956,N_9240,N_9578);
and U9957 (N_9957,N_9469,N_9382);
nand U9958 (N_9958,N_9311,N_9348);
or U9959 (N_9959,N_9456,N_9283);
xor U9960 (N_9960,N_9574,N_9437);
or U9961 (N_9961,N_9387,N_9288);
nor U9962 (N_9962,N_9417,N_9221);
nand U9963 (N_9963,N_9581,N_9375);
nand U9964 (N_9964,N_9454,N_9319);
xor U9965 (N_9965,N_9580,N_9463);
nand U9966 (N_9966,N_9307,N_9329);
nor U9967 (N_9967,N_9356,N_9473);
nor U9968 (N_9968,N_9481,N_9562);
or U9969 (N_9969,N_9409,N_9300);
nor U9970 (N_9970,N_9425,N_9241);
and U9971 (N_9971,N_9373,N_9555);
or U9972 (N_9972,N_9584,N_9594);
nor U9973 (N_9973,N_9417,N_9414);
nand U9974 (N_9974,N_9276,N_9493);
nand U9975 (N_9975,N_9475,N_9222);
nand U9976 (N_9976,N_9532,N_9206);
or U9977 (N_9977,N_9500,N_9210);
nor U9978 (N_9978,N_9509,N_9241);
nand U9979 (N_9979,N_9524,N_9482);
and U9980 (N_9980,N_9213,N_9220);
or U9981 (N_9981,N_9321,N_9312);
xor U9982 (N_9982,N_9376,N_9485);
and U9983 (N_9983,N_9440,N_9315);
and U9984 (N_9984,N_9582,N_9268);
nand U9985 (N_9985,N_9331,N_9372);
nand U9986 (N_9986,N_9529,N_9411);
xnor U9987 (N_9987,N_9532,N_9252);
nor U9988 (N_9988,N_9297,N_9219);
and U9989 (N_9989,N_9366,N_9599);
xor U9990 (N_9990,N_9496,N_9446);
or U9991 (N_9991,N_9421,N_9565);
or U9992 (N_9992,N_9352,N_9495);
or U9993 (N_9993,N_9386,N_9205);
and U9994 (N_9994,N_9374,N_9574);
nor U9995 (N_9995,N_9527,N_9578);
xnor U9996 (N_9996,N_9501,N_9523);
or U9997 (N_9997,N_9504,N_9590);
and U9998 (N_9998,N_9241,N_9358);
nor U9999 (N_9999,N_9374,N_9297);
nand U10000 (N_10000,N_9780,N_9618);
xor U10001 (N_10001,N_9905,N_9972);
xnor U10002 (N_10002,N_9878,N_9638);
xnor U10003 (N_10003,N_9975,N_9977);
nand U10004 (N_10004,N_9758,N_9919);
nand U10005 (N_10005,N_9818,N_9898);
and U10006 (N_10006,N_9856,N_9640);
nor U10007 (N_10007,N_9921,N_9808);
nand U10008 (N_10008,N_9994,N_9860);
xnor U10009 (N_10009,N_9614,N_9723);
or U10010 (N_10010,N_9846,N_9785);
nor U10011 (N_10011,N_9991,N_9658);
xnor U10012 (N_10012,N_9872,N_9828);
nor U10013 (N_10013,N_9830,N_9945);
and U10014 (N_10014,N_9955,N_9939);
xor U10015 (N_10015,N_9601,N_9980);
and U10016 (N_10016,N_9622,N_9967);
xor U10017 (N_10017,N_9678,N_9854);
or U10018 (N_10018,N_9679,N_9687);
and U10019 (N_10019,N_9888,N_9716);
nand U10020 (N_10020,N_9677,N_9989);
and U10021 (N_10021,N_9913,N_9613);
xnor U10022 (N_10022,N_9793,N_9660);
or U10023 (N_10023,N_9901,N_9603);
nor U10024 (N_10024,N_9739,N_9686);
xnor U10025 (N_10025,N_9670,N_9762);
nand U10026 (N_10026,N_9949,N_9766);
and U10027 (N_10027,N_9884,N_9639);
nor U10028 (N_10028,N_9784,N_9732);
or U10029 (N_10029,N_9769,N_9862);
or U10030 (N_10030,N_9733,N_9692);
nand U10031 (N_10031,N_9998,N_9761);
nor U10032 (N_10032,N_9688,N_9729);
or U10033 (N_10033,N_9942,N_9805);
and U10034 (N_10034,N_9668,N_9944);
nand U10035 (N_10035,N_9834,N_9709);
xnor U10036 (N_10036,N_9877,N_9705);
and U10037 (N_10037,N_9671,N_9615);
or U10038 (N_10038,N_9985,N_9701);
or U10039 (N_10039,N_9867,N_9801);
nand U10040 (N_10040,N_9861,N_9753);
nor U10041 (N_10041,N_9796,N_9759);
and U10042 (N_10042,N_9683,N_9857);
and U10043 (N_10043,N_9804,N_9864);
and U10044 (N_10044,N_9620,N_9868);
xor U10045 (N_10045,N_9858,N_9950);
nand U10046 (N_10046,N_9772,N_9715);
xnor U10047 (N_10047,N_9912,N_9737);
nor U10048 (N_10048,N_9958,N_9665);
xnor U10049 (N_10049,N_9866,N_9629);
nand U10050 (N_10050,N_9681,N_9782);
xor U10051 (N_10051,N_9617,N_9875);
nor U10052 (N_10052,N_9833,N_9806);
and U10053 (N_10053,N_9891,N_9979);
nor U10054 (N_10054,N_9881,N_9676);
or U10055 (N_10055,N_9797,N_9844);
and U10056 (N_10056,N_9771,N_9812);
and U10057 (N_10057,N_9814,N_9837);
nor U10058 (N_10058,N_9633,N_9829);
nand U10059 (N_10059,N_9963,N_9971);
or U10060 (N_10060,N_9654,N_9611);
and U10061 (N_10061,N_9662,N_9917);
nor U10062 (N_10062,N_9841,N_9689);
nor U10063 (N_10063,N_9685,N_9885);
xor U10064 (N_10064,N_9970,N_9648);
and U10065 (N_10065,N_9775,N_9938);
or U10066 (N_10066,N_9840,N_9672);
nor U10067 (N_10067,N_9653,N_9988);
xor U10068 (N_10068,N_9634,N_9798);
nor U10069 (N_10069,N_9932,N_9961);
nand U10070 (N_10070,N_9920,N_9876);
nor U10071 (N_10071,N_9787,N_9616);
nor U10072 (N_10072,N_9974,N_9722);
and U10073 (N_10073,N_9773,N_9986);
nor U10074 (N_10074,N_9643,N_9711);
or U10075 (N_10075,N_9790,N_9734);
xnor U10076 (N_10076,N_9951,N_9776);
and U10077 (N_10077,N_9800,N_9838);
nor U10078 (N_10078,N_9853,N_9900);
xor U10079 (N_10079,N_9702,N_9887);
and U10080 (N_10080,N_9730,N_9821);
nor U10081 (N_10081,N_9667,N_9946);
nor U10082 (N_10082,N_9778,N_9751);
xor U10083 (N_10083,N_9843,N_9628);
nand U10084 (N_10084,N_9682,N_9695);
xor U10085 (N_10085,N_9926,N_9902);
nand U10086 (N_10086,N_9948,N_9930);
or U10087 (N_10087,N_9605,N_9707);
or U10088 (N_10088,N_9981,N_9791);
nor U10089 (N_10089,N_9726,N_9630);
nor U10090 (N_10090,N_9893,N_9959);
xor U10091 (N_10091,N_9720,N_9934);
nor U10092 (N_10092,N_9673,N_9651);
or U10093 (N_10093,N_9799,N_9916);
nand U10094 (N_10094,N_9906,N_9604);
nor U10095 (N_10095,N_9624,N_9774);
nor U10096 (N_10096,N_9755,N_9703);
nand U10097 (N_10097,N_9815,N_9742);
nand U10098 (N_10098,N_9645,N_9823);
nand U10099 (N_10099,N_9767,N_9915);
nor U10100 (N_10100,N_9849,N_9623);
xor U10101 (N_10101,N_9817,N_9928);
nand U10102 (N_10102,N_9855,N_9714);
and U10103 (N_10103,N_9704,N_9770);
nand U10104 (N_10104,N_9941,N_9822);
nand U10105 (N_10105,N_9914,N_9612);
or U10106 (N_10106,N_9978,N_9803);
nand U10107 (N_10107,N_9721,N_9600);
xor U10108 (N_10108,N_9680,N_9710);
and U10109 (N_10109,N_9847,N_9674);
nand U10110 (N_10110,N_9819,N_9727);
xnor U10111 (N_10111,N_9691,N_9659);
or U10112 (N_10112,N_9883,N_9957);
nand U10113 (N_10113,N_9807,N_9728);
or U10114 (N_10114,N_9954,N_9811);
xor U10115 (N_10115,N_9777,N_9999);
or U10116 (N_10116,N_9863,N_9700);
and U10117 (N_10117,N_9602,N_9927);
xor U10118 (N_10118,N_9698,N_9735);
or U10119 (N_10119,N_9896,N_9925);
and U10120 (N_10120,N_9663,N_9936);
and U10121 (N_10121,N_9990,N_9907);
nor U10122 (N_10122,N_9717,N_9610);
nor U10123 (N_10123,N_9779,N_9874);
nand U10124 (N_10124,N_9749,N_9783);
or U10125 (N_10125,N_9724,N_9836);
or U10126 (N_10126,N_9696,N_9897);
and U10127 (N_10127,N_9831,N_9652);
and U10128 (N_10128,N_9606,N_9940);
nor U10129 (N_10129,N_9816,N_9802);
xor U10130 (N_10130,N_9746,N_9657);
nor U10131 (N_10131,N_9738,N_9669);
xor U10132 (N_10132,N_9982,N_9983);
and U10133 (N_10133,N_9655,N_9992);
or U10134 (N_10134,N_9786,N_9664);
or U10135 (N_10135,N_9924,N_9873);
and U10136 (N_10136,N_9943,N_9824);
and U10137 (N_10137,N_9731,N_9996);
and U10138 (N_10138,N_9973,N_9952);
nand U10139 (N_10139,N_9923,N_9956);
xnor U10140 (N_10140,N_9747,N_9741);
and U10141 (N_10141,N_9642,N_9666);
and U10142 (N_10142,N_9910,N_9997);
xnor U10143 (N_10143,N_9851,N_9607);
xnor U10144 (N_10144,N_9865,N_9756);
or U10145 (N_10145,N_9810,N_9719);
and U10146 (N_10146,N_9895,N_9764);
xnor U10147 (N_10147,N_9889,N_9627);
nand U10148 (N_10148,N_9760,N_9641);
or U10149 (N_10149,N_9933,N_9969);
and U10150 (N_10150,N_9694,N_9965);
xor U10151 (N_10151,N_9995,N_9706);
nand U10152 (N_10152,N_9647,N_9937);
xnor U10153 (N_10153,N_9632,N_9725);
xor U10154 (N_10154,N_9795,N_9832);
xor U10155 (N_10155,N_9820,N_9848);
and U10156 (N_10156,N_9792,N_9609);
or U10157 (N_10157,N_9740,N_9768);
nor U10158 (N_10158,N_9646,N_9964);
nand U10159 (N_10159,N_9908,N_9636);
nand U10160 (N_10160,N_9931,N_9835);
and U10161 (N_10161,N_9649,N_9635);
or U10162 (N_10162,N_9839,N_9870);
or U10163 (N_10163,N_9693,N_9929);
nand U10164 (N_10164,N_9637,N_9650);
and U10165 (N_10165,N_9765,N_9718);
and U10166 (N_10166,N_9763,N_9621);
nand U10167 (N_10167,N_9656,N_9743);
or U10168 (N_10168,N_9966,N_9744);
xor U10169 (N_10169,N_9947,N_9911);
or U10170 (N_10170,N_9697,N_9745);
nor U10171 (N_10171,N_9788,N_9619);
or U10172 (N_10172,N_9750,N_9984);
nand U10173 (N_10173,N_9752,N_9713);
nand U10174 (N_10174,N_9626,N_9842);
nand U10175 (N_10175,N_9850,N_9754);
nand U10176 (N_10176,N_9890,N_9880);
xor U10177 (N_10177,N_9882,N_9661);
nand U10178 (N_10178,N_9625,N_9899);
nand U10179 (N_10179,N_9826,N_9675);
nand U10180 (N_10180,N_9871,N_9886);
nand U10181 (N_10181,N_9904,N_9976);
nand U10182 (N_10182,N_9794,N_9993);
xnor U10183 (N_10183,N_9953,N_9922);
or U10184 (N_10184,N_9644,N_9892);
or U10185 (N_10185,N_9869,N_9894);
xnor U10186 (N_10186,N_9748,N_9879);
or U10187 (N_10187,N_9960,N_9903);
and U10188 (N_10188,N_9781,N_9813);
nand U10189 (N_10189,N_9757,N_9708);
nor U10190 (N_10190,N_9859,N_9935);
and U10191 (N_10191,N_9712,N_9968);
and U10192 (N_10192,N_9789,N_9684);
nand U10193 (N_10193,N_9987,N_9909);
nor U10194 (N_10194,N_9852,N_9918);
xnor U10195 (N_10195,N_9690,N_9825);
nor U10196 (N_10196,N_9827,N_9845);
xor U10197 (N_10197,N_9962,N_9736);
and U10198 (N_10198,N_9608,N_9631);
xor U10199 (N_10199,N_9699,N_9809);
or U10200 (N_10200,N_9655,N_9952);
nand U10201 (N_10201,N_9878,N_9796);
xor U10202 (N_10202,N_9949,N_9953);
nand U10203 (N_10203,N_9823,N_9847);
xor U10204 (N_10204,N_9716,N_9799);
nand U10205 (N_10205,N_9941,N_9993);
and U10206 (N_10206,N_9857,N_9729);
xor U10207 (N_10207,N_9741,N_9607);
nor U10208 (N_10208,N_9933,N_9627);
nor U10209 (N_10209,N_9997,N_9816);
nor U10210 (N_10210,N_9871,N_9876);
nor U10211 (N_10211,N_9642,N_9716);
and U10212 (N_10212,N_9786,N_9629);
nand U10213 (N_10213,N_9702,N_9683);
xnor U10214 (N_10214,N_9877,N_9913);
and U10215 (N_10215,N_9829,N_9851);
or U10216 (N_10216,N_9780,N_9608);
or U10217 (N_10217,N_9902,N_9704);
nand U10218 (N_10218,N_9667,N_9962);
xor U10219 (N_10219,N_9994,N_9686);
nand U10220 (N_10220,N_9659,N_9901);
nand U10221 (N_10221,N_9741,N_9601);
xnor U10222 (N_10222,N_9650,N_9785);
nand U10223 (N_10223,N_9745,N_9978);
nor U10224 (N_10224,N_9748,N_9967);
nand U10225 (N_10225,N_9915,N_9829);
nand U10226 (N_10226,N_9928,N_9903);
nand U10227 (N_10227,N_9806,N_9624);
nand U10228 (N_10228,N_9644,N_9780);
or U10229 (N_10229,N_9696,N_9869);
and U10230 (N_10230,N_9896,N_9667);
nor U10231 (N_10231,N_9801,N_9968);
nor U10232 (N_10232,N_9905,N_9644);
or U10233 (N_10233,N_9713,N_9662);
nor U10234 (N_10234,N_9751,N_9925);
nor U10235 (N_10235,N_9967,N_9738);
and U10236 (N_10236,N_9677,N_9927);
xnor U10237 (N_10237,N_9605,N_9681);
and U10238 (N_10238,N_9969,N_9691);
xor U10239 (N_10239,N_9906,N_9644);
nor U10240 (N_10240,N_9601,N_9872);
nor U10241 (N_10241,N_9693,N_9931);
or U10242 (N_10242,N_9611,N_9959);
and U10243 (N_10243,N_9817,N_9797);
or U10244 (N_10244,N_9844,N_9649);
nand U10245 (N_10245,N_9738,N_9910);
nand U10246 (N_10246,N_9994,N_9905);
nor U10247 (N_10247,N_9911,N_9865);
and U10248 (N_10248,N_9989,N_9794);
or U10249 (N_10249,N_9794,N_9766);
xor U10250 (N_10250,N_9983,N_9699);
and U10251 (N_10251,N_9630,N_9756);
nor U10252 (N_10252,N_9800,N_9791);
nand U10253 (N_10253,N_9663,N_9853);
nor U10254 (N_10254,N_9648,N_9702);
or U10255 (N_10255,N_9627,N_9789);
or U10256 (N_10256,N_9677,N_9753);
nand U10257 (N_10257,N_9697,N_9739);
nor U10258 (N_10258,N_9877,N_9988);
nand U10259 (N_10259,N_9987,N_9965);
and U10260 (N_10260,N_9718,N_9819);
nand U10261 (N_10261,N_9818,N_9656);
xor U10262 (N_10262,N_9791,N_9744);
and U10263 (N_10263,N_9720,N_9600);
and U10264 (N_10264,N_9779,N_9995);
and U10265 (N_10265,N_9991,N_9788);
nor U10266 (N_10266,N_9864,N_9679);
xor U10267 (N_10267,N_9687,N_9911);
and U10268 (N_10268,N_9945,N_9842);
nand U10269 (N_10269,N_9676,N_9927);
nor U10270 (N_10270,N_9605,N_9774);
xor U10271 (N_10271,N_9911,N_9739);
and U10272 (N_10272,N_9722,N_9940);
nor U10273 (N_10273,N_9642,N_9628);
and U10274 (N_10274,N_9805,N_9939);
or U10275 (N_10275,N_9861,N_9755);
or U10276 (N_10276,N_9793,N_9619);
or U10277 (N_10277,N_9908,N_9795);
or U10278 (N_10278,N_9806,N_9761);
nor U10279 (N_10279,N_9938,N_9955);
or U10280 (N_10280,N_9909,N_9895);
nor U10281 (N_10281,N_9942,N_9630);
nor U10282 (N_10282,N_9983,N_9763);
or U10283 (N_10283,N_9753,N_9999);
or U10284 (N_10284,N_9857,N_9829);
nor U10285 (N_10285,N_9728,N_9892);
nand U10286 (N_10286,N_9634,N_9839);
nand U10287 (N_10287,N_9652,N_9827);
nor U10288 (N_10288,N_9895,N_9631);
or U10289 (N_10289,N_9747,N_9854);
nand U10290 (N_10290,N_9611,N_9610);
and U10291 (N_10291,N_9756,N_9694);
or U10292 (N_10292,N_9887,N_9750);
nand U10293 (N_10293,N_9635,N_9941);
and U10294 (N_10294,N_9637,N_9762);
nand U10295 (N_10295,N_9737,N_9730);
nand U10296 (N_10296,N_9804,N_9741);
nor U10297 (N_10297,N_9729,N_9691);
nor U10298 (N_10298,N_9796,N_9731);
nor U10299 (N_10299,N_9682,N_9790);
nand U10300 (N_10300,N_9824,N_9774);
and U10301 (N_10301,N_9642,N_9896);
nand U10302 (N_10302,N_9907,N_9731);
nor U10303 (N_10303,N_9682,N_9759);
nor U10304 (N_10304,N_9602,N_9616);
nand U10305 (N_10305,N_9835,N_9651);
xnor U10306 (N_10306,N_9846,N_9880);
nor U10307 (N_10307,N_9995,N_9608);
nor U10308 (N_10308,N_9946,N_9694);
or U10309 (N_10309,N_9685,N_9998);
or U10310 (N_10310,N_9951,N_9866);
xnor U10311 (N_10311,N_9671,N_9738);
nand U10312 (N_10312,N_9690,N_9923);
xor U10313 (N_10313,N_9629,N_9792);
or U10314 (N_10314,N_9698,N_9830);
nor U10315 (N_10315,N_9826,N_9961);
or U10316 (N_10316,N_9645,N_9615);
nand U10317 (N_10317,N_9910,N_9687);
xnor U10318 (N_10318,N_9740,N_9848);
nand U10319 (N_10319,N_9759,N_9819);
and U10320 (N_10320,N_9659,N_9987);
and U10321 (N_10321,N_9906,N_9683);
nor U10322 (N_10322,N_9831,N_9713);
nand U10323 (N_10323,N_9916,N_9800);
nor U10324 (N_10324,N_9858,N_9911);
or U10325 (N_10325,N_9662,N_9600);
nand U10326 (N_10326,N_9977,N_9735);
or U10327 (N_10327,N_9914,N_9823);
xnor U10328 (N_10328,N_9663,N_9998);
nand U10329 (N_10329,N_9889,N_9905);
or U10330 (N_10330,N_9797,N_9970);
nand U10331 (N_10331,N_9683,N_9860);
nand U10332 (N_10332,N_9643,N_9737);
and U10333 (N_10333,N_9857,N_9949);
xor U10334 (N_10334,N_9891,N_9801);
nor U10335 (N_10335,N_9612,N_9907);
or U10336 (N_10336,N_9797,N_9798);
xor U10337 (N_10337,N_9967,N_9855);
xor U10338 (N_10338,N_9873,N_9996);
xnor U10339 (N_10339,N_9833,N_9861);
nor U10340 (N_10340,N_9991,N_9969);
and U10341 (N_10341,N_9861,N_9846);
nor U10342 (N_10342,N_9846,N_9691);
nand U10343 (N_10343,N_9961,N_9708);
and U10344 (N_10344,N_9696,N_9653);
and U10345 (N_10345,N_9627,N_9852);
and U10346 (N_10346,N_9826,N_9788);
xnor U10347 (N_10347,N_9716,N_9620);
or U10348 (N_10348,N_9646,N_9979);
xor U10349 (N_10349,N_9777,N_9768);
nand U10350 (N_10350,N_9750,N_9944);
xor U10351 (N_10351,N_9830,N_9994);
xor U10352 (N_10352,N_9706,N_9972);
nor U10353 (N_10353,N_9988,N_9989);
xnor U10354 (N_10354,N_9928,N_9628);
xor U10355 (N_10355,N_9843,N_9734);
and U10356 (N_10356,N_9972,N_9620);
or U10357 (N_10357,N_9848,N_9771);
nand U10358 (N_10358,N_9893,N_9710);
or U10359 (N_10359,N_9891,N_9992);
xnor U10360 (N_10360,N_9727,N_9680);
and U10361 (N_10361,N_9646,N_9694);
or U10362 (N_10362,N_9877,N_9996);
xor U10363 (N_10363,N_9726,N_9811);
and U10364 (N_10364,N_9840,N_9890);
and U10365 (N_10365,N_9728,N_9623);
nand U10366 (N_10366,N_9961,N_9971);
nor U10367 (N_10367,N_9656,N_9788);
nand U10368 (N_10368,N_9718,N_9632);
or U10369 (N_10369,N_9630,N_9982);
nand U10370 (N_10370,N_9669,N_9664);
nand U10371 (N_10371,N_9748,N_9810);
nand U10372 (N_10372,N_9679,N_9995);
and U10373 (N_10373,N_9830,N_9886);
xor U10374 (N_10374,N_9600,N_9950);
nor U10375 (N_10375,N_9743,N_9912);
and U10376 (N_10376,N_9603,N_9634);
xnor U10377 (N_10377,N_9833,N_9615);
and U10378 (N_10378,N_9735,N_9782);
or U10379 (N_10379,N_9748,N_9935);
or U10380 (N_10380,N_9966,N_9631);
nor U10381 (N_10381,N_9782,N_9824);
nand U10382 (N_10382,N_9602,N_9686);
nand U10383 (N_10383,N_9886,N_9842);
and U10384 (N_10384,N_9664,N_9828);
nor U10385 (N_10385,N_9745,N_9924);
nor U10386 (N_10386,N_9617,N_9784);
and U10387 (N_10387,N_9760,N_9683);
nand U10388 (N_10388,N_9793,N_9750);
and U10389 (N_10389,N_9972,N_9700);
nand U10390 (N_10390,N_9920,N_9633);
nand U10391 (N_10391,N_9663,N_9691);
xnor U10392 (N_10392,N_9909,N_9705);
and U10393 (N_10393,N_9746,N_9834);
and U10394 (N_10394,N_9752,N_9771);
xor U10395 (N_10395,N_9915,N_9792);
xnor U10396 (N_10396,N_9992,N_9881);
xor U10397 (N_10397,N_9899,N_9758);
and U10398 (N_10398,N_9874,N_9899);
or U10399 (N_10399,N_9895,N_9698);
or U10400 (N_10400,N_10106,N_10278);
or U10401 (N_10401,N_10337,N_10009);
nor U10402 (N_10402,N_10262,N_10343);
or U10403 (N_10403,N_10230,N_10390);
nand U10404 (N_10404,N_10370,N_10158);
nor U10405 (N_10405,N_10076,N_10237);
nor U10406 (N_10406,N_10312,N_10268);
or U10407 (N_10407,N_10177,N_10305);
or U10408 (N_10408,N_10124,N_10293);
or U10409 (N_10409,N_10236,N_10347);
xnor U10410 (N_10410,N_10214,N_10064);
nor U10411 (N_10411,N_10067,N_10189);
and U10412 (N_10412,N_10297,N_10166);
xor U10413 (N_10413,N_10099,N_10168);
and U10414 (N_10414,N_10093,N_10160);
and U10415 (N_10415,N_10211,N_10386);
xor U10416 (N_10416,N_10169,N_10101);
xnor U10417 (N_10417,N_10216,N_10391);
xnor U10418 (N_10418,N_10273,N_10152);
nor U10419 (N_10419,N_10342,N_10065);
or U10420 (N_10420,N_10136,N_10366);
and U10421 (N_10421,N_10069,N_10353);
and U10422 (N_10422,N_10143,N_10284);
nor U10423 (N_10423,N_10203,N_10084);
nand U10424 (N_10424,N_10181,N_10039);
nand U10425 (N_10425,N_10184,N_10311);
or U10426 (N_10426,N_10049,N_10033);
and U10427 (N_10427,N_10030,N_10204);
nor U10428 (N_10428,N_10345,N_10005);
or U10429 (N_10429,N_10012,N_10326);
xor U10430 (N_10430,N_10397,N_10265);
nand U10431 (N_10431,N_10062,N_10376);
nor U10432 (N_10432,N_10144,N_10306);
nand U10433 (N_10433,N_10162,N_10250);
xnor U10434 (N_10434,N_10307,N_10344);
nand U10435 (N_10435,N_10229,N_10220);
nor U10436 (N_10436,N_10255,N_10154);
nor U10437 (N_10437,N_10015,N_10314);
nor U10438 (N_10438,N_10209,N_10113);
nand U10439 (N_10439,N_10210,N_10227);
nor U10440 (N_10440,N_10118,N_10339);
xnor U10441 (N_10441,N_10226,N_10096);
or U10442 (N_10442,N_10318,N_10327);
nor U10443 (N_10443,N_10087,N_10240);
nand U10444 (N_10444,N_10358,N_10291);
nor U10445 (N_10445,N_10129,N_10008);
nor U10446 (N_10446,N_10175,N_10384);
and U10447 (N_10447,N_10336,N_10253);
and U10448 (N_10448,N_10092,N_10023);
xnor U10449 (N_10449,N_10040,N_10356);
nand U10450 (N_10450,N_10082,N_10334);
xnor U10451 (N_10451,N_10288,N_10200);
nor U10452 (N_10452,N_10222,N_10324);
xor U10453 (N_10453,N_10004,N_10287);
and U10454 (N_10454,N_10285,N_10019);
nand U10455 (N_10455,N_10219,N_10246);
nor U10456 (N_10456,N_10025,N_10252);
and U10457 (N_10457,N_10244,N_10059);
nor U10458 (N_10458,N_10289,N_10257);
nor U10459 (N_10459,N_10322,N_10385);
nand U10460 (N_10460,N_10186,N_10316);
nor U10461 (N_10461,N_10080,N_10223);
xnor U10462 (N_10462,N_10134,N_10215);
nor U10463 (N_10463,N_10302,N_10125);
or U10464 (N_10464,N_10061,N_10355);
nand U10465 (N_10465,N_10224,N_10021);
xnor U10466 (N_10466,N_10114,N_10310);
nand U10467 (N_10467,N_10034,N_10392);
xor U10468 (N_10468,N_10235,N_10340);
nand U10469 (N_10469,N_10298,N_10281);
nand U10470 (N_10470,N_10380,N_10041);
nor U10471 (N_10471,N_10266,N_10196);
and U10472 (N_10472,N_10116,N_10123);
xnor U10473 (N_10473,N_10270,N_10044);
or U10474 (N_10474,N_10017,N_10170);
xor U10475 (N_10475,N_10301,N_10072);
nand U10476 (N_10476,N_10313,N_10395);
or U10477 (N_10477,N_10037,N_10263);
nand U10478 (N_10478,N_10042,N_10098);
and U10479 (N_10479,N_10102,N_10052);
nand U10480 (N_10480,N_10055,N_10243);
nand U10481 (N_10481,N_10117,N_10028);
nor U10482 (N_10482,N_10317,N_10173);
and U10483 (N_10483,N_10018,N_10225);
nor U10484 (N_10484,N_10001,N_10259);
and U10485 (N_10485,N_10232,N_10105);
and U10486 (N_10486,N_10341,N_10373);
xor U10487 (N_10487,N_10060,N_10205);
nand U10488 (N_10488,N_10176,N_10103);
nand U10489 (N_10489,N_10132,N_10047);
nor U10490 (N_10490,N_10145,N_10038);
or U10491 (N_10491,N_10085,N_10212);
nand U10492 (N_10492,N_10011,N_10365);
or U10493 (N_10493,N_10182,N_10398);
nand U10494 (N_10494,N_10321,N_10007);
nand U10495 (N_10495,N_10024,N_10388);
and U10496 (N_10496,N_10187,N_10239);
nor U10497 (N_10497,N_10354,N_10066);
nand U10498 (N_10498,N_10165,N_10126);
nor U10499 (N_10499,N_10112,N_10379);
and U10500 (N_10500,N_10050,N_10248);
and U10501 (N_10501,N_10382,N_10375);
nand U10502 (N_10502,N_10381,N_10083);
xor U10503 (N_10503,N_10120,N_10071);
or U10504 (N_10504,N_10371,N_10190);
nor U10505 (N_10505,N_10128,N_10241);
and U10506 (N_10506,N_10221,N_10127);
and U10507 (N_10507,N_10014,N_10027);
xnor U10508 (N_10508,N_10256,N_10146);
xnor U10509 (N_10509,N_10058,N_10111);
nand U10510 (N_10510,N_10308,N_10079);
and U10511 (N_10511,N_10264,N_10006);
xor U10512 (N_10512,N_10100,N_10197);
and U10513 (N_10513,N_10218,N_10156);
or U10514 (N_10514,N_10303,N_10258);
or U10515 (N_10515,N_10192,N_10247);
nand U10516 (N_10516,N_10315,N_10164);
or U10517 (N_10517,N_10150,N_10013);
nand U10518 (N_10518,N_10329,N_10022);
and U10519 (N_10519,N_10360,N_10290);
nand U10520 (N_10520,N_10333,N_10213);
or U10521 (N_10521,N_10323,N_10167);
or U10522 (N_10522,N_10346,N_10350);
or U10523 (N_10523,N_10286,N_10148);
xor U10524 (N_10524,N_10238,N_10073);
and U10525 (N_10525,N_10074,N_10130);
nand U10526 (N_10526,N_10294,N_10359);
nor U10527 (N_10527,N_10097,N_10026);
nand U10528 (N_10528,N_10399,N_10280);
or U10529 (N_10529,N_10029,N_10000);
nor U10530 (N_10530,N_10319,N_10367);
nor U10531 (N_10531,N_10279,N_10325);
and U10532 (N_10532,N_10078,N_10107);
nor U10533 (N_10533,N_10185,N_10335);
nand U10534 (N_10534,N_10003,N_10140);
xor U10535 (N_10535,N_10198,N_10194);
and U10536 (N_10536,N_10332,N_10063);
or U10537 (N_10537,N_10271,N_10174);
and U10538 (N_10538,N_10094,N_10108);
or U10539 (N_10539,N_10245,N_10031);
and U10540 (N_10540,N_10191,N_10352);
and U10541 (N_10541,N_10155,N_10233);
and U10542 (N_10542,N_10057,N_10163);
xnor U10543 (N_10543,N_10095,N_10172);
nor U10544 (N_10544,N_10141,N_10208);
xor U10545 (N_10545,N_10304,N_10161);
and U10546 (N_10546,N_10394,N_10153);
nor U10547 (N_10547,N_10299,N_10300);
or U10548 (N_10548,N_10374,N_10362);
or U10549 (N_10549,N_10193,N_10046);
xor U10550 (N_10550,N_10231,N_10296);
nor U10551 (N_10551,N_10396,N_10179);
nand U10552 (N_10552,N_10051,N_10089);
nand U10553 (N_10553,N_10151,N_10357);
nor U10554 (N_10554,N_10070,N_10201);
nor U10555 (N_10555,N_10045,N_10122);
and U10556 (N_10556,N_10274,N_10251);
nand U10557 (N_10557,N_10242,N_10135);
or U10558 (N_10558,N_10282,N_10010);
or U10559 (N_10559,N_10207,N_10183);
xnor U10560 (N_10560,N_10292,N_10088);
and U10561 (N_10561,N_10199,N_10036);
or U10562 (N_10562,N_10149,N_10142);
nor U10563 (N_10563,N_10138,N_10228);
or U10564 (N_10564,N_10171,N_10147);
nor U10565 (N_10565,N_10188,N_10378);
nor U10566 (N_10566,N_10159,N_10269);
xor U10567 (N_10567,N_10202,N_10331);
and U10568 (N_10568,N_10260,N_10090);
xnor U10569 (N_10569,N_10368,N_10234);
nor U10570 (N_10570,N_10081,N_10275);
and U10571 (N_10571,N_10309,N_10115);
and U10572 (N_10572,N_10020,N_10377);
and U10573 (N_10573,N_10283,N_10261);
nand U10574 (N_10574,N_10389,N_10217);
xnor U10575 (N_10575,N_10075,N_10056);
nand U10576 (N_10576,N_10387,N_10338);
nor U10577 (N_10577,N_10077,N_10104);
nand U10578 (N_10578,N_10137,N_10295);
xnor U10579 (N_10579,N_10180,N_10393);
nand U10580 (N_10580,N_10043,N_10048);
and U10581 (N_10581,N_10249,N_10016);
xnor U10582 (N_10582,N_10277,N_10320);
and U10583 (N_10583,N_10035,N_10276);
nand U10584 (N_10584,N_10178,N_10267);
or U10585 (N_10585,N_10121,N_10119);
nand U10586 (N_10586,N_10133,N_10002);
nor U10587 (N_10587,N_10109,N_10372);
or U10588 (N_10588,N_10351,N_10054);
or U10589 (N_10589,N_10157,N_10364);
and U10590 (N_10590,N_10131,N_10369);
xor U10591 (N_10591,N_10139,N_10330);
and U10592 (N_10592,N_10383,N_10068);
or U10593 (N_10593,N_10348,N_10110);
or U10594 (N_10594,N_10349,N_10032);
nand U10595 (N_10595,N_10195,N_10206);
or U10596 (N_10596,N_10272,N_10328);
nor U10597 (N_10597,N_10254,N_10086);
and U10598 (N_10598,N_10363,N_10361);
nor U10599 (N_10599,N_10091,N_10053);
and U10600 (N_10600,N_10016,N_10178);
or U10601 (N_10601,N_10275,N_10291);
nand U10602 (N_10602,N_10223,N_10376);
xor U10603 (N_10603,N_10383,N_10070);
nor U10604 (N_10604,N_10110,N_10231);
nor U10605 (N_10605,N_10139,N_10255);
nand U10606 (N_10606,N_10255,N_10064);
or U10607 (N_10607,N_10299,N_10161);
xor U10608 (N_10608,N_10100,N_10046);
and U10609 (N_10609,N_10007,N_10030);
nand U10610 (N_10610,N_10395,N_10087);
xor U10611 (N_10611,N_10212,N_10217);
nor U10612 (N_10612,N_10304,N_10128);
and U10613 (N_10613,N_10245,N_10087);
nand U10614 (N_10614,N_10321,N_10206);
and U10615 (N_10615,N_10394,N_10082);
and U10616 (N_10616,N_10396,N_10342);
and U10617 (N_10617,N_10291,N_10143);
nor U10618 (N_10618,N_10167,N_10182);
nand U10619 (N_10619,N_10067,N_10160);
xor U10620 (N_10620,N_10342,N_10146);
nor U10621 (N_10621,N_10129,N_10362);
and U10622 (N_10622,N_10016,N_10043);
nand U10623 (N_10623,N_10219,N_10094);
nand U10624 (N_10624,N_10032,N_10071);
nand U10625 (N_10625,N_10228,N_10215);
xnor U10626 (N_10626,N_10054,N_10276);
or U10627 (N_10627,N_10052,N_10154);
xor U10628 (N_10628,N_10297,N_10084);
nand U10629 (N_10629,N_10042,N_10318);
nand U10630 (N_10630,N_10090,N_10191);
xor U10631 (N_10631,N_10231,N_10008);
xnor U10632 (N_10632,N_10170,N_10325);
nand U10633 (N_10633,N_10202,N_10064);
or U10634 (N_10634,N_10331,N_10284);
xor U10635 (N_10635,N_10238,N_10222);
nand U10636 (N_10636,N_10138,N_10264);
or U10637 (N_10637,N_10272,N_10398);
and U10638 (N_10638,N_10002,N_10163);
nand U10639 (N_10639,N_10220,N_10044);
xor U10640 (N_10640,N_10249,N_10133);
nand U10641 (N_10641,N_10078,N_10013);
nand U10642 (N_10642,N_10335,N_10385);
xnor U10643 (N_10643,N_10322,N_10323);
nand U10644 (N_10644,N_10363,N_10133);
and U10645 (N_10645,N_10193,N_10399);
or U10646 (N_10646,N_10136,N_10290);
nor U10647 (N_10647,N_10192,N_10287);
nor U10648 (N_10648,N_10284,N_10261);
nand U10649 (N_10649,N_10105,N_10240);
xor U10650 (N_10650,N_10004,N_10385);
or U10651 (N_10651,N_10051,N_10171);
or U10652 (N_10652,N_10276,N_10306);
or U10653 (N_10653,N_10136,N_10167);
nor U10654 (N_10654,N_10098,N_10176);
nor U10655 (N_10655,N_10354,N_10396);
nor U10656 (N_10656,N_10193,N_10268);
nor U10657 (N_10657,N_10310,N_10122);
or U10658 (N_10658,N_10234,N_10184);
nand U10659 (N_10659,N_10192,N_10001);
nand U10660 (N_10660,N_10360,N_10152);
and U10661 (N_10661,N_10234,N_10319);
nand U10662 (N_10662,N_10118,N_10310);
xnor U10663 (N_10663,N_10191,N_10189);
or U10664 (N_10664,N_10358,N_10082);
nor U10665 (N_10665,N_10329,N_10345);
xnor U10666 (N_10666,N_10203,N_10198);
xnor U10667 (N_10667,N_10358,N_10296);
or U10668 (N_10668,N_10089,N_10170);
xor U10669 (N_10669,N_10132,N_10070);
and U10670 (N_10670,N_10130,N_10179);
xor U10671 (N_10671,N_10034,N_10004);
nor U10672 (N_10672,N_10344,N_10366);
or U10673 (N_10673,N_10324,N_10011);
nand U10674 (N_10674,N_10279,N_10091);
nor U10675 (N_10675,N_10169,N_10174);
nor U10676 (N_10676,N_10121,N_10058);
and U10677 (N_10677,N_10346,N_10103);
or U10678 (N_10678,N_10255,N_10332);
xnor U10679 (N_10679,N_10030,N_10130);
or U10680 (N_10680,N_10165,N_10208);
xnor U10681 (N_10681,N_10186,N_10029);
or U10682 (N_10682,N_10344,N_10365);
nand U10683 (N_10683,N_10148,N_10107);
xnor U10684 (N_10684,N_10153,N_10081);
or U10685 (N_10685,N_10209,N_10337);
or U10686 (N_10686,N_10244,N_10336);
or U10687 (N_10687,N_10192,N_10299);
nor U10688 (N_10688,N_10333,N_10259);
and U10689 (N_10689,N_10282,N_10228);
or U10690 (N_10690,N_10026,N_10128);
or U10691 (N_10691,N_10184,N_10318);
or U10692 (N_10692,N_10189,N_10351);
nor U10693 (N_10693,N_10293,N_10113);
nand U10694 (N_10694,N_10319,N_10064);
and U10695 (N_10695,N_10195,N_10341);
or U10696 (N_10696,N_10020,N_10051);
nor U10697 (N_10697,N_10097,N_10159);
nor U10698 (N_10698,N_10340,N_10398);
nand U10699 (N_10699,N_10100,N_10056);
nor U10700 (N_10700,N_10023,N_10201);
or U10701 (N_10701,N_10066,N_10209);
nor U10702 (N_10702,N_10006,N_10097);
and U10703 (N_10703,N_10381,N_10384);
or U10704 (N_10704,N_10064,N_10007);
and U10705 (N_10705,N_10032,N_10391);
and U10706 (N_10706,N_10158,N_10200);
nand U10707 (N_10707,N_10319,N_10018);
nand U10708 (N_10708,N_10178,N_10199);
xor U10709 (N_10709,N_10285,N_10388);
or U10710 (N_10710,N_10098,N_10026);
nand U10711 (N_10711,N_10189,N_10235);
nand U10712 (N_10712,N_10158,N_10354);
nand U10713 (N_10713,N_10244,N_10046);
and U10714 (N_10714,N_10104,N_10044);
and U10715 (N_10715,N_10355,N_10378);
xor U10716 (N_10716,N_10357,N_10065);
xnor U10717 (N_10717,N_10072,N_10119);
xnor U10718 (N_10718,N_10193,N_10316);
nor U10719 (N_10719,N_10241,N_10064);
nand U10720 (N_10720,N_10034,N_10151);
or U10721 (N_10721,N_10136,N_10016);
or U10722 (N_10722,N_10060,N_10070);
and U10723 (N_10723,N_10251,N_10238);
xnor U10724 (N_10724,N_10087,N_10148);
nand U10725 (N_10725,N_10243,N_10023);
nand U10726 (N_10726,N_10047,N_10274);
nand U10727 (N_10727,N_10074,N_10068);
or U10728 (N_10728,N_10318,N_10349);
xnor U10729 (N_10729,N_10127,N_10194);
and U10730 (N_10730,N_10201,N_10242);
nor U10731 (N_10731,N_10288,N_10199);
and U10732 (N_10732,N_10122,N_10274);
and U10733 (N_10733,N_10157,N_10128);
nor U10734 (N_10734,N_10110,N_10038);
xor U10735 (N_10735,N_10045,N_10380);
or U10736 (N_10736,N_10085,N_10366);
nor U10737 (N_10737,N_10361,N_10279);
xnor U10738 (N_10738,N_10348,N_10202);
nand U10739 (N_10739,N_10117,N_10148);
nand U10740 (N_10740,N_10055,N_10244);
nor U10741 (N_10741,N_10096,N_10057);
or U10742 (N_10742,N_10266,N_10134);
nand U10743 (N_10743,N_10011,N_10133);
or U10744 (N_10744,N_10070,N_10384);
and U10745 (N_10745,N_10397,N_10050);
nor U10746 (N_10746,N_10227,N_10228);
and U10747 (N_10747,N_10125,N_10210);
nor U10748 (N_10748,N_10201,N_10016);
nand U10749 (N_10749,N_10196,N_10083);
nand U10750 (N_10750,N_10052,N_10032);
and U10751 (N_10751,N_10372,N_10180);
xor U10752 (N_10752,N_10274,N_10031);
and U10753 (N_10753,N_10162,N_10180);
nor U10754 (N_10754,N_10078,N_10209);
nand U10755 (N_10755,N_10341,N_10190);
and U10756 (N_10756,N_10124,N_10222);
and U10757 (N_10757,N_10092,N_10364);
xor U10758 (N_10758,N_10375,N_10369);
xnor U10759 (N_10759,N_10287,N_10238);
xor U10760 (N_10760,N_10261,N_10260);
or U10761 (N_10761,N_10085,N_10290);
nor U10762 (N_10762,N_10251,N_10258);
nand U10763 (N_10763,N_10225,N_10250);
xor U10764 (N_10764,N_10331,N_10049);
nand U10765 (N_10765,N_10083,N_10171);
and U10766 (N_10766,N_10376,N_10178);
xor U10767 (N_10767,N_10388,N_10023);
nor U10768 (N_10768,N_10041,N_10190);
or U10769 (N_10769,N_10220,N_10124);
or U10770 (N_10770,N_10318,N_10236);
or U10771 (N_10771,N_10062,N_10160);
nor U10772 (N_10772,N_10276,N_10329);
or U10773 (N_10773,N_10183,N_10038);
nand U10774 (N_10774,N_10145,N_10185);
nor U10775 (N_10775,N_10268,N_10124);
nand U10776 (N_10776,N_10207,N_10275);
xnor U10777 (N_10777,N_10293,N_10268);
nor U10778 (N_10778,N_10380,N_10309);
xor U10779 (N_10779,N_10071,N_10315);
nor U10780 (N_10780,N_10218,N_10166);
nor U10781 (N_10781,N_10014,N_10164);
nand U10782 (N_10782,N_10035,N_10109);
nor U10783 (N_10783,N_10384,N_10246);
xor U10784 (N_10784,N_10084,N_10334);
nor U10785 (N_10785,N_10355,N_10354);
xnor U10786 (N_10786,N_10354,N_10264);
nand U10787 (N_10787,N_10328,N_10340);
nor U10788 (N_10788,N_10021,N_10131);
nor U10789 (N_10789,N_10224,N_10117);
or U10790 (N_10790,N_10305,N_10068);
nor U10791 (N_10791,N_10180,N_10172);
nand U10792 (N_10792,N_10150,N_10108);
nor U10793 (N_10793,N_10395,N_10273);
and U10794 (N_10794,N_10031,N_10351);
nand U10795 (N_10795,N_10352,N_10006);
and U10796 (N_10796,N_10215,N_10326);
or U10797 (N_10797,N_10284,N_10236);
xor U10798 (N_10798,N_10172,N_10047);
or U10799 (N_10799,N_10055,N_10156);
xor U10800 (N_10800,N_10796,N_10660);
or U10801 (N_10801,N_10700,N_10505);
and U10802 (N_10802,N_10637,N_10754);
or U10803 (N_10803,N_10669,N_10748);
or U10804 (N_10804,N_10607,N_10483);
or U10805 (N_10805,N_10516,N_10632);
and U10806 (N_10806,N_10639,N_10477);
or U10807 (N_10807,N_10690,N_10560);
xnor U10808 (N_10808,N_10545,N_10712);
and U10809 (N_10809,N_10458,N_10586);
xnor U10810 (N_10810,N_10565,N_10664);
nand U10811 (N_10811,N_10523,N_10490);
and U10812 (N_10812,N_10487,N_10645);
or U10813 (N_10813,N_10503,N_10549);
nor U10814 (N_10814,N_10631,N_10504);
nor U10815 (N_10815,N_10750,N_10581);
and U10816 (N_10816,N_10555,N_10563);
nor U10817 (N_10817,N_10696,N_10622);
xnor U10818 (N_10818,N_10770,N_10451);
or U10819 (N_10819,N_10765,N_10780);
and U10820 (N_10820,N_10649,N_10550);
xor U10821 (N_10821,N_10764,N_10432);
nor U10822 (N_10822,N_10424,N_10492);
xnor U10823 (N_10823,N_10556,N_10615);
nor U10824 (N_10824,N_10528,N_10566);
nand U10825 (N_10825,N_10464,N_10459);
nor U10826 (N_10826,N_10575,N_10657);
and U10827 (N_10827,N_10489,N_10533);
or U10828 (N_10828,N_10418,N_10595);
xor U10829 (N_10829,N_10731,N_10784);
and U10830 (N_10830,N_10618,N_10701);
xor U10831 (N_10831,N_10732,N_10559);
xor U10832 (N_10832,N_10496,N_10501);
or U10833 (N_10833,N_10768,N_10538);
nand U10834 (N_10834,N_10561,N_10756);
xnor U10835 (N_10835,N_10469,N_10456);
nand U10836 (N_10836,N_10776,N_10710);
nor U10837 (N_10837,N_10769,N_10402);
or U10838 (N_10838,N_10414,N_10602);
nand U10839 (N_10839,N_10715,N_10479);
nand U10840 (N_10840,N_10447,N_10634);
and U10841 (N_10841,N_10584,N_10659);
or U10842 (N_10842,N_10423,N_10761);
and U10843 (N_10843,N_10546,N_10400);
nor U10844 (N_10844,N_10404,N_10544);
nand U10845 (N_10845,N_10497,N_10653);
xnor U10846 (N_10846,N_10431,N_10727);
nor U10847 (N_10847,N_10564,N_10789);
or U10848 (N_10848,N_10486,N_10795);
nor U10849 (N_10849,N_10623,N_10766);
nor U10850 (N_10850,N_10798,N_10510);
xor U10851 (N_10851,N_10612,N_10594);
or U10852 (N_10852,N_10788,N_10433);
xnor U10853 (N_10853,N_10472,N_10635);
nor U10854 (N_10854,N_10774,N_10707);
nand U10855 (N_10855,N_10452,N_10482);
or U10856 (N_10856,N_10587,N_10751);
and U10857 (N_10857,N_10576,N_10790);
nor U10858 (N_10858,N_10512,N_10427);
nor U10859 (N_10859,N_10743,N_10408);
nor U10860 (N_10860,N_10684,N_10573);
nand U10861 (N_10861,N_10666,N_10763);
nand U10862 (N_10862,N_10711,N_10735);
and U10863 (N_10863,N_10643,N_10668);
and U10864 (N_10864,N_10494,N_10797);
nor U10865 (N_10865,N_10597,N_10692);
and U10866 (N_10866,N_10683,N_10685);
nor U10867 (N_10867,N_10500,N_10702);
xnor U10868 (N_10868,N_10740,N_10484);
xor U10869 (N_10869,N_10542,N_10686);
nor U10870 (N_10870,N_10552,N_10524);
nor U10871 (N_10871,N_10613,N_10722);
nor U10872 (N_10872,N_10579,N_10536);
and U10873 (N_10873,N_10688,N_10445);
nand U10874 (N_10874,N_10694,N_10428);
xnor U10875 (N_10875,N_10415,N_10409);
xnor U10876 (N_10876,N_10728,N_10589);
or U10877 (N_10877,N_10583,N_10434);
and U10878 (N_10878,N_10629,N_10453);
nand U10879 (N_10879,N_10411,N_10729);
and U10880 (N_10880,N_10440,N_10437);
nand U10881 (N_10881,N_10407,N_10718);
nand U10882 (N_10882,N_10651,N_10435);
and U10883 (N_10883,N_10470,N_10706);
xnor U10884 (N_10884,N_10616,N_10717);
and U10885 (N_10885,N_10682,N_10778);
nor U10886 (N_10886,N_10703,N_10713);
xor U10887 (N_10887,N_10695,N_10534);
or U10888 (N_10888,N_10783,N_10614);
and U10889 (N_10889,N_10760,N_10572);
or U10890 (N_10890,N_10767,N_10509);
nor U10891 (N_10891,N_10526,N_10689);
xnor U10892 (N_10892,N_10539,N_10551);
xnor U10893 (N_10893,N_10599,N_10749);
and U10894 (N_10894,N_10596,N_10633);
xor U10895 (N_10895,N_10498,N_10481);
nand U10896 (N_10896,N_10515,N_10541);
nand U10897 (N_10897,N_10513,N_10792);
xor U10898 (N_10898,N_10465,N_10720);
xnor U10899 (N_10899,N_10442,N_10582);
nand U10900 (N_10900,N_10678,N_10600);
and U10901 (N_10901,N_10708,N_10590);
or U10902 (N_10902,N_10744,N_10671);
or U10903 (N_10903,N_10741,N_10777);
and U10904 (N_10904,N_10719,N_10450);
and U10905 (N_10905,N_10518,N_10532);
nor U10906 (N_10906,N_10604,N_10517);
nand U10907 (N_10907,N_10454,N_10785);
nor U10908 (N_10908,N_10775,N_10473);
nand U10909 (N_10909,N_10709,N_10675);
nand U10910 (N_10910,N_10679,N_10755);
nand U10911 (N_10911,N_10762,N_10488);
xnor U10912 (N_10912,N_10401,N_10606);
nand U10913 (N_10913,N_10624,N_10562);
or U10914 (N_10914,N_10665,N_10648);
nand U10915 (N_10915,N_10733,N_10508);
nor U10916 (N_10916,N_10530,N_10738);
nor U10917 (N_10917,N_10422,N_10406);
xor U10918 (N_10918,N_10621,N_10674);
nor U10919 (N_10919,N_10759,N_10593);
and U10920 (N_10920,N_10598,N_10568);
or U10921 (N_10921,N_10742,N_10673);
nand U10922 (N_10922,N_10499,N_10519);
nor U10923 (N_10923,N_10571,N_10646);
and U10924 (N_10924,N_10667,N_10485);
xor U10925 (N_10925,N_10570,N_10609);
xor U10926 (N_10926,N_10529,N_10724);
or U10927 (N_10927,N_10662,N_10480);
nand U10928 (N_10928,N_10537,N_10558);
xnor U10929 (N_10929,N_10478,N_10620);
nand U10930 (N_10930,N_10677,N_10627);
xnor U10931 (N_10931,N_10676,N_10577);
or U10932 (N_10932,N_10641,N_10467);
or U10933 (N_10933,N_10421,N_10787);
xor U10934 (N_10934,N_10672,N_10753);
nor U10935 (N_10935,N_10691,N_10548);
nand U10936 (N_10936,N_10611,N_10468);
and U10937 (N_10937,N_10547,N_10757);
and U10938 (N_10938,N_10791,N_10773);
nand U10939 (N_10939,N_10495,N_10779);
xor U10940 (N_10940,N_10725,N_10557);
nand U10941 (N_10941,N_10507,N_10772);
xor U10942 (N_10942,N_10697,N_10540);
nand U10943 (N_10943,N_10580,N_10739);
or U10944 (N_10944,N_10543,N_10723);
nand U10945 (N_10945,N_10412,N_10567);
xnor U10946 (N_10946,N_10578,N_10799);
or U10947 (N_10947,N_10475,N_10603);
nor U10948 (N_10948,N_10569,N_10736);
or U10949 (N_10949,N_10658,N_10535);
xor U10950 (N_10950,N_10655,N_10636);
nor U10951 (N_10951,N_10714,N_10721);
or U10952 (N_10952,N_10680,N_10640);
xor U10953 (N_10953,N_10514,N_10413);
or U10954 (N_10954,N_10608,N_10446);
nor U10955 (N_10955,N_10617,N_10610);
and U10956 (N_10956,N_10444,N_10511);
nand U10957 (N_10957,N_10420,N_10416);
nand U10958 (N_10958,N_10786,N_10705);
or U10959 (N_10959,N_10730,N_10782);
and U10960 (N_10960,N_10471,N_10661);
nand U10961 (N_10961,N_10687,N_10531);
nor U10962 (N_10962,N_10455,N_10430);
xor U10963 (N_10963,N_10476,N_10448);
or U10964 (N_10964,N_10436,N_10502);
nand U10965 (N_10965,N_10463,N_10734);
and U10966 (N_10966,N_10793,N_10588);
nand U10967 (N_10967,N_10474,N_10461);
xnor U10968 (N_10968,N_10522,N_10747);
nand U10969 (N_10969,N_10726,N_10520);
nor U10970 (N_10970,N_10745,N_10650);
nand U10971 (N_10971,N_10425,N_10521);
or U10972 (N_10972,N_10405,N_10601);
nor U10973 (N_10973,N_10626,N_10628);
xnor U10974 (N_10974,N_10449,N_10716);
nand U10975 (N_10975,N_10457,N_10527);
nor U10976 (N_10976,N_10781,N_10506);
nand U10977 (N_10977,N_10642,N_10758);
nor U10978 (N_10978,N_10652,N_10746);
or U10979 (N_10979,N_10698,N_10663);
and U10980 (N_10980,N_10605,N_10443);
nor U10981 (N_10981,N_10439,N_10466);
nor U10982 (N_10982,N_10419,N_10554);
xnor U10983 (N_10983,N_10647,N_10681);
and U10984 (N_10984,N_10462,N_10670);
nor U10985 (N_10985,N_10625,N_10619);
xnor U10986 (N_10986,N_10460,N_10429);
nand U10987 (N_10987,N_10630,N_10553);
nand U10988 (N_10988,N_10654,N_10441);
xnor U10989 (N_10989,N_10794,N_10704);
nor U10990 (N_10990,N_10403,N_10656);
nor U10991 (N_10991,N_10771,N_10491);
xnor U10992 (N_10992,N_10693,N_10426);
and U10993 (N_10993,N_10410,N_10737);
or U10994 (N_10994,N_10591,N_10417);
xor U10995 (N_10995,N_10438,N_10574);
nor U10996 (N_10996,N_10644,N_10493);
xor U10997 (N_10997,N_10699,N_10525);
nand U10998 (N_10998,N_10752,N_10592);
nand U10999 (N_10999,N_10638,N_10585);
nand U11000 (N_11000,N_10490,N_10615);
and U11001 (N_11001,N_10719,N_10773);
xor U11002 (N_11002,N_10755,N_10592);
xor U11003 (N_11003,N_10507,N_10400);
nor U11004 (N_11004,N_10451,N_10620);
or U11005 (N_11005,N_10481,N_10548);
or U11006 (N_11006,N_10443,N_10455);
xor U11007 (N_11007,N_10524,N_10571);
xnor U11008 (N_11008,N_10760,N_10518);
or U11009 (N_11009,N_10424,N_10693);
xor U11010 (N_11010,N_10549,N_10622);
and U11011 (N_11011,N_10408,N_10616);
or U11012 (N_11012,N_10652,N_10487);
or U11013 (N_11013,N_10614,N_10672);
nor U11014 (N_11014,N_10624,N_10791);
xnor U11015 (N_11015,N_10784,N_10595);
or U11016 (N_11016,N_10585,N_10620);
xnor U11017 (N_11017,N_10546,N_10620);
or U11018 (N_11018,N_10687,N_10543);
nor U11019 (N_11019,N_10664,N_10728);
nor U11020 (N_11020,N_10527,N_10501);
nor U11021 (N_11021,N_10703,N_10649);
xor U11022 (N_11022,N_10747,N_10455);
xor U11023 (N_11023,N_10774,N_10596);
nor U11024 (N_11024,N_10516,N_10432);
nor U11025 (N_11025,N_10658,N_10714);
xor U11026 (N_11026,N_10743,N_10567);
or U11027 (N_11027,N_10700,N_10661);
and U11028 (N_11028,N_10602,N_10410);
xnor U11029 (N_11029,N_10448,N_10569);
nand U11030 (N_11030,N_10739,N_10755);
and U11031 (N_11031,N_10583,N_10522);
or U11032 (N_11032,N_10451,N_10669);
xor U11033 (N_11033,N_10504,N_10617);
nor U11034 (N_11034,N_10467,N_10660);
xor U11035 (N_11035,N_10732,N_10582);
xor U11036 (N_11036,N_10565,N_10542);
nand U11037 (N_11037,N_10484,N_10762);
nand U11038 (N_11038,N_10570,N_10782);
nand U11039 (N_11039,N_10701,N_10620);
and U11040 (N_11040,N_10724,N_10774);
or U11041 (N_11041,N_10496,N_10602);
xnor U11042 (N_11042,N_10419,N_10417);
nand U11043 (N_11043,N_10490,N_10416);
nor U11044 (N_11044,N_10715,N_10581);
xnor U11045 (N_11045,N_10601,N_10798);
or U11046 (N_11046,N_10673,N_10409);
nor U11047 (N_11047,N_10472,N_10776);
nand U11048 (N_11048,N_10701,N_10581);
or U11049 (N_11049,N_10651,N_10699);
nor U11050 (N_11050,N_10517,N_10426);
and U11051 (N_11051,N_10453,N_10754);
xnor U11052 (N_11052,N_10546,N_10739);
nand U11053 (N_11053,N_10784,N_10531);
xnor U11054 (N_11054,N_10518,N_10783);
or U11055 (N_11055,N_10604,N_10636);
nand U11056 (N_11056,N_10733,N_10749);
and U11057 (N_11057,N_10612,N_10572);
or U11058 (N_11058,N_10486,N_10768);
and U11059 (N_11059,N_10718,N_10736);
nor U11060 (N_11060,N_10784,N_10710);
xnor U11061 (N_11061,N_10760,N_10491);
nand U11062 (N_11062,N_10479,N_10695);
xor U11063 (N_11063,N_10758,N_10727);
and U11064 (N_11064,N_10583,N_10664);
nor U11065 (N_11065,N_10548,N_10547);
nor U11066 (N_11066,N_10486,N_10773);
nand U11067 (N_11067,N_10513,N_10613);
xnor U11068 (N_11068,N_10609,N_10644);
nand U11069 (N_11069,N_10462,N_10476);
or U11070 (N_11070,N_10772,N_10552);
nand U11071 (N_11071,N_10422,N_10457);
nor U11072 (N_11072,N_10603,N_10439);
nand U11073 (N_11073,N_10522,N_10505);
and U11074 (N_11074,N_10477,N_10498);
nand U11075 (N_11075,N_10604,N_10439);
nand U11076 (N_11076,N_10477,N_10685);
or U11077 (N_11077,N_10765,N_10511);
nand U11078 (N_11078,N_10654,N_10706);
xnor U11079 (N_11079,N_10487,N_10525);
or U11080 (N_11080,N_10618,N_10762);
or U11081 (N_11081,N_10644,N_10555);
xor U11082 (N_11082,N_10769,N_10527);
xnor U11083 (N_11083,N_10490,N_10646);
and U11084 (N_11084,N_10467,N_10764);
nor U11085 (N_11085,N_10526,N_10494);
nand U11086 (N_11086,N_10419,N_10618);
nor U11087 (N_11087,N_10420,N_10624);
and U11088 (N_11088,N_10595,N_10443);
and U11089 (N_11089,N_10680,N_10418);
or U11090 (N_11090,N_10404,N_10508);
or U11091 (N_11091,N_10425,N_10748);
nand U11092 (N_11092,N_10754,N_10593);
and U11093 (N_11093,N_10583,N_10518);
xor U11094 (N_11094,N_10622,N_10625);
nand U11095 (N_11095,N_10570,N_10439);
nor U11096 (N_11096,N_10489,N_10544);
xnor U11097 (N_11097,N_10741,N_10426);
or U11098 (N_11098,N_10679,N_10458);
or U11099 (N_11099,N_10610,N_10657);
xnor U11100 (N_11100,N_10581,N_10604);
and U11101 (N_11101,N_10686,N_10407);
or U11102 (N_11102,N_10682,N_10690);
nor U11103 (N_11103,N_10644,N_10623);
or U11104 (N_11104,N_10785,N_10537);
nor U11105 (N_11105,N_10694,N_10686);
nor U11106 (N_11106,N_10519,N_10448);
and U11107 (N_11107,N_10495,N_10660);
and U11108 (N_11108,N_10749,N_10583);
or U11109 (N_11109,N_10542,N_10728);
and U11110 (N_11110,N_10462,N_10514);
nand U11111 (N_11111,N_10746,N_10500);
nand U11112 (N_11112,N_10549,N_10612);
nand U11113 (N_11113,N_10421,N_10789);
or U11114 (N_11114,N_10688,N_10665);
xor U11115 (N_11115,N_10585,N_10671);
nor U11116 (N_11116,N_10493,N_10448);
xnor U11117 (N_11117,N_10684,N_10743);
or U11118 (N_11118,N_10492,N_10758);
nand U11119 (N_11119,N_10449,N_10794);
or U11120 (N_11120,N_10759,N_10474);
or U11121 (N_11121,N_10788,N_10635);
and U11122 (N_11122,N_10585,N_10792);
and U11123 (N_11123,N_10531,N_10655);
nand U11124 (N_11124,N_10769,N_10553);
or U11125 (N_11125,N_10734,N_10437);
or U11126 (N_11126,N_10646,N_10758);
and U11127 (N_11127,N_10746,N_10695);
or U11128 (N_11128,N_10713,N_10711);
nor U11129 (N_11129,N_10436,N_10511);
xor U11130 (N_11130,N_10610,N_10559);
or U11131 (N_11131,N_10508,N_10485);
nor U11132 (N_11132,N_10798,N_10796);
xor U11133 (N_11133,N_10455,N_10453);
nand U11134 (N_11134,N_10799,N_10656);
and U11135 (N_11135,N_10637,N_10682);
nor U11136 (N_11136,N_10748,N_10698);
xnor U11137 (N_11137,N_10517,N_10676);
or U11138 (N_11138,N_10499,N_10737);
xor U11139 (N_11139,N_10685,N_10468);
xor U11140 (N_11140,N_10405,N_10600);
xnor U11141 (N_11141,N_10502,N_10696);
nand U11142 (N_11142,N_10419,N_10575);
or U11143 (N_11143,N_10792,N_10688);
or U11144 (N_11144,N_10708,N_10498);
and U11145 (N_11145,N_10602,N_10585);
and U11146 (N_11146,N_10418,N_10600);
and U11147 (N_11147,N_10668,N_10431);
nor U11148 (N_11148,N_10507,N_10706);
xor U11149 (N_11149,N_10653,N_10509);
nand U11150 (N_11150,N_10644,N_10434);
and U11151 (N_11151,N_10449,N_10645);
xnor U11152 (N_11152,N_10729,N_10678);
xnor U11153 (N_11153,N_10537,N_10559);
xnor U11154 (N_11154,N_10586,N_10521);
and U11155 (N_11155,N_10724,N_10570);
or U11156 (N_11156,N_10725,N_10615);
or U11157 (N_11157,N_10673,N_10565);
xnor U11158 (N_11158,N_10636,N_10787);
and U11159 (N_11159,N_10629,N_10448);
nand U11160 (N_11160,N_10702,N_10677);
nor U11161 (N_11161,N_10540,N_10525);
nor U11162 (N_11162,N_10655,N_10411);
nand U11163 (N_11163,N_10551,N_10795);
xnor U11164 (N_11164,N_10567,N_10533);
nor U11165 (N_11165,N_10412,N_10782);
nor U11166 (N_11166,N_10579,N_10696);
nand U11167 (N_11167,N_10757,N_10743);
nor U11168 (N_11168,N_10626,N_10410);
xnor U11169 (N_11169,N_10686,N_10541);
xnor U11170 (N_11170,N_10711,N_10607);
nor U11171 (N_11171,N_10412,N_10602);
xnor U11172 (N_11172,N_10637,N_10763);
nor U11173 (N_11173,N_10471,N_10784);
and U11174 (N_11174,N_10775,N_10430);
and U11175 (N_11175,N_10475,N_10448);
xnor U11176 (N_11176,N_10741,N_10780);
or U11177 (N_11177,N_10591,N_10506);
and U11178 (N_11178,N_10741,N_10408);
and U11179 (N_11179,N_10671,N_10662);
xnor U11180 (N_11180,N_10665,N_10792);
nor U11181 (N_11181,N_10428,N_10511);
xnor U11182 (N_11182,N_10568,N_10457);
or U11183 (N_11183,N_10791,N_10744);
xnor U11184 (N_11184,N_10579,N_10655);
nand U11185 (N_11185,N_10404,N_10786);
xor U11186 (N_11186,N_10593,N_10529);
and U11187 (N_11187,N_10733,N_10678);
or U11188 (N_11188,N_10737,N_10669);
or U11189 (N_11189,N_10753,N_10739);
nand U11190 (N_11190,N_10595,N_10629);
xnor U11191 (N_11191,N_10568,N_10737);
or U11192 (N_11192,N_10504,N_10621);
nor U11193 (N_11193,N_10549,N_10585);
xnor U11194 (N_11194,N_10703,N_10619);
nand U11195 (N_11195,N_10681,N_10773);
and U11196 (N_11196,N_10643,N_10468);
nand U11197 (N_11197,N_10403,N_10558);
and U11198 (N_11198,N_10795,N_10495);
and U11199 (N_11199,N_10624,N_10548);
nor U11200 (N_11200,N_10846,N_11095);
and U11201 (N_11201,N_10954,N_10810);
or U11202 (N_11202,N_11016,N_10977);
xor U11203 (N_11203,N_11085,N_10880);
or U11204 (N_11204,N_11093,N_10816);
nor U11205 (N_11205,N_10902,N_10866);
nor U11206 (N_11206,N_10979,N_10921);
nor U11207 (N_11207,N_10886,N_11104);
nor U11208 (N_11208,N_11120,N_11133);
or U11209 (N_11209,N_10829,N_10917);
xnor U11210 (N_11210,N_11025,N_11186);
xor U11211 (N_11211,N_10830,N_11000);
and U11212 (N_11212,N_10833,N_11043);
nand U11213 (N_11213,N_11013,N_10962);
and U11214 (N_11214,N_11007,N_10950);
nand U11215 (N_11215,N_11144,N_11111);
or U11216 (N_11216,N_11166,N_10865);
nor U11217 (N_11217,N_11114,N_10906);
nand U11218 (N_11218,N_11102,N_11097);
nand U11219 (N_11219,N_11056,N_10915);
nand U11220 (N_11220,N_10879,N_11146);
and U11221 (N_11221,N_10802,N_10847);
nor U11222 (N_11222,N_11059,N_11149);
or U11223 (N_11223,N_10965,N_10956);
nand U11224 (N_11224,N_11193,N_11198);
or U11225 (N_11225,N_11130,N_10986);
and U11226 (N_11226,N_10887,N_11073);
xor U11227 (N_11227,N_11018,N_10985);
xnor U11228 (N_11228,N_10849,N_11113);
nand U11229 (N_11229,N_10836,N_10850);
and U11230 (N_11230,N_10938,N_10934);
xnor U11231 (N_11231,N_10852,N_11152);
xor U11232 (N_11232,N_10868,N_10825);
nand U11233 (N_11233,N_11068,N_11036);
and U11234 (N_11234,N_10922,N_11080);
and U11235 (N_11235,N_10894,N_10871);
and U11236 (N_11236,N_11042,N_10885);
nand U11237 (N_11237,N_10939,N_11086);
nand U11238 (N_11238,N_11127,N_11094);
nand U11239 (N_11239,N_10893,N_11026);
nor U11240 (N_11240,N_11183,N_11090);
and U11241 (N_11241,N_11039,N_11185);
xnor U11242 (N_11242,N_11063,N_11033);
or U11243 (N_11243,N_11184,N_10867);
nor U11244 (N_11244,N_11199,N_11099);
xnor U11245 (N_11245,N_11157,N_11156);
nor U11246 (N_11246,N_11066,N_11053);
and U11247 (N_11247,N_10976,N_10980);
nor U11248 (N_11248,N_11055,N_10820);
nor U11249 (N_11249,N_10856,N_10914);
nand U11250 (N_11250,N_10883,N_11048);
nor U11251 (N_11251,N_11164,N_10996);
xnor U11252 (N_11252,N_11159,N_10933);
nor U11253 (N_11253,N_11139,N_10990);
nor U11254 (N_11254,N_11151,N_11006);
nor U11255 (N_11255,N_11100,N_11058);
nand U11256 (N_11256,N_11008,N_10862);
or U11257 (N_11257,N_10801,N_10839);
or U11258 (N_11258,N_11150,N_10978);
or U11259 (N_11259,N_10834,N_10910);
or U11260 (N_11260,N_10875,N_10814);
nor U11261 (N_11261,N_11037,N_10890);
and U11262 (N_11262,N_11004,N_11024);
nor U11263 (N_11263,N_10824,N_10972);
and U11264 (N_11264,N_10861,N_11019);
or U11265 (N_11265,N_11163,N_11119);
nand U11266 (N_11266,N_11064,N_11060);
nand U11267 (N_11267,N_11088,N_10928);
xor U11268 (N_11268,N_11027,N_10940);
and U11269 (N_11269,N_11129,N_11096);
nor U11270 (N_11270,N_10907,N_10878);
or U11271 (N_11271,N_10998,N_11167);
nand U11272 (N_11272,N_10805,N_11194);
and U11273 (N_11273,N_11049,N_10817);
nor U11274 (N_11274,N_11170,N_11112);
nor U11275 (N_11275,N_11136,N_10935);
nor U11276 (N_11276,N_10903,N_11030);
or U11277 (N_11277,N_10900,N_10920);
and U11278 (N_11278,N_11128,N_11158);
nor U11279 (N_11279,N_11069,N_11134);
and U11280 (N_11280,N_11040,N_11074);
nor U11281 (N_11281,N_11161,N_11190);
or U11282 (N_11282,N_10995,N_10813);
or U11283 (N_11283,N_10970,N_11118);
nor U11284 (N_11284,N_10869,N_11179);
nand U11285 (N_11285,N_11005,N_11177);
or U11286 (N_11286,N_11022,N_11014);
nor U11287 (N_11287,N_11017,N_10819);
and U11288 (N_11288,N_11105,N_10924);
nand U11289 (N_11289,N_10835,N_11141);
and U11290 (N_11290,N_10993,N_10831);
nor U11291 (N_11291,N_10844,N_10937);
nand U11292 (N_11292,N_10851,N_11192);
nor U11293 (N_11293,N_10930,N_10947);
and U11294 (N_11294,N_11160,N_11154);
nand U11295 (N_11295,N_11123,N_11155);
or U11296 (N_11296,N_11009,N_11142);
xor U11297 (N_11297,N_11181,N_11138);
xor U11298 (N_11298,N_11089,N_10895);
xnor U11299 (N_11299,N_11083,N_10911);
xnor U11300 (N_11300,N_11173,N_10842);
nor U11301 (N_11301,N_10918,N_11145);
or U11302 (N_11302,N_10859,N_10872);
nand U11303 (N_11303,N_11122,N_11046);
and U11304 (N_11304,N_10973,N_11050);
and U11305 (N_11305,N_10806,N_10837);
nand U11306 (N_11306,N_11125,N_10888);
nand U11307 (N_11307,N_10951,N_10864);
or U11308 (N_11308,N_11067,N_10845);
nor U11309 (N_11309,N_11035,N_10964);
or U11310 (N_11310,N_10919,N_10955);
xor U11311 (N_11311,N_10901,N_10969);
nor U11312 (N_11312,N_10984,N_10828);
xor U11313 (N_11313,N_10958,N_10876);
xor U11314 (N_11314,N_10891,N_10925);
xnor U11315 (N_11315,N_11041,N_11061);
xor U11316 (N_11316,N_10800,N_10988);
or U11317 (N_11317,N_10932,N_10812);
or U11318 (N_11318,N_10853,N_11098);
xor U11319 (N_11319,N_10943,N_10912);
xnor U11320 (N_11320,N_10841,N_11121);
and U11321 (N_11321,N_10981,N_10823);
and U11322 (N_11322,N_10874,N_10909);
nand U11323 (N_11323,N_11011,N_11110);
nand U11324 (N_11324,N_11168,N_11148);
nor U11325 (N_11325,N_11126,N_10863);
xor U11326 (N_11326,N_11010,N_10960);
nor U11327 (N_11327,N_11002,N_10929);
nor U11328 (N_11328,N_11180,N_10804);
nor U11329 (N_11329,N_10884,N_11051);
nand U11330 (N_11330,N_11197,N_10822);
or U11331 (N_11331,N_10961,N_10897);
and U11332 (N_11332,N_11103,N_11078);
and U11333 (N_11333,N_11143,N_10987);
nand U11334 (N_11334,N_10923,N_10811);
nand U11335 (N_11335,N_10968,N_10899);
nor U11336 (N_11336,N_10966,N_10873);
or U11337 (N_11337,N_10854,N_11003);
xor U11338 (N_11338,N_11188,N_10881);
xor U11339 (N_11339,N_10963,N_11191);
xnor U11340 (N_11340,N_10971,N_11189);
or U11341 (N_11341,N_11165,N_10944);
or U11342 (N_11342,N_10858,N_10832);
or U11343 (N_11343,N_10848,N_11172);
or U11344 (N_11344,N_10967,N_10941);
and U11345 (N_11345,N_11052,N_10908);
and U11346 (N_11346,N_10889,N_11115);
nor U11347 (N_11347,N_10843,N_11109);
or U11348 (N_11348,N_11087,N_10931);
xnor U11349 (N_11349,N_11081,N_11101);
and U11350 (N_11350,N_11029,N_10855);
nand U11351 (N_11351,N_10815,N_10926);
and U11352 (N_11352,N_11171,N_10936);
nand U11353 (N_11353,N_10945,N_10989);
and U11354 (N_11354,N_11031,N_11107);
nor U11355 (N_11355,N_10991,N_11178);
nand U11356 (N_11356,N_11015,N_10857);
and U11357 (N_11357,N_11038,N_10826);
nand U11358 (N_11358,N_11117,N_11072);
and U11359 (N_11359,N_11108,N_10896);
and U11360 (N_11360,N_10953,N_10949);
and U11361 (N_11361,N_10860,N_10840);
nand U11362 (N_11362,N_10808,N_11076);
nand U11363 (N_11363,N_10999,N_11169);
nor U11364 (N_11364,N_10974,N_11196);
nor U11365 (N_11365,N_11131,N_11054);
and U11366 (N_11366,N_11023,N_10892);
and U11367 (N_11367,N_10946,N_11092);
and U11368 (N_11368,N_10904,N_11045);
nand U11369 (N_11369,N_11187,N_10959);
or U11370 (N_11370,N_10838,N_10913);
and U11371 (N_11371,N_11075,N_11047);
nand U11372 (N_11372,N_11124,N_11001);
or U11373 (N_11373,N_10992,N_11071);
nand U11374 (N_11374,N_11084,N_10983);
or U11375 (N_11375,N_11091,N_10898);
and U11376 (N_11376,N_10818,N_11028);
xor U11377 (N_11377,N_11147,N_10927);
and U11378 (N_11378,N_11176,N_11065);
xor U11379 (N_11379,N_11153,N_11062);
nor U11380 (N_11380,N_10975,N_10957);
xnor U11381 (N_11381,N_11182,N_10807);
xnor U11382 (N_11382,N_10905,N_10942);
xnor U11383 (N_11383,N_11032,N_10882);
nor U11384 (N_11384,N_11057,N_11195);
and U11385 (N_11385,N_10809,N_11140);
or U11386 (N_11386,N_10821,N_10827);
nand U11387 (N_11387,N_11044,N_10994);
and U11388 (N_11388,N_11137,N_10948);
nand U11389 (N_11389,N_10982,N_11116);
or U11390 (N_11390,N_11021,N_11034);
and U11391 (N_11391,N_11132,N_10916);
nor U11392 (N_11392,N_11162,N_10952);
nor U11393 (N_11393,N_11020,N_11106);
and U11394 (N_11394,N_10803,N_11077);
and U11395 (N_11395,N_11135,N_11082);
and U11396 (N_11396,N_10997,N_11012);
or U11397 (N_11397,N_11175,N_11070);
or U11398 (N_11398,N_10870,N_10877);
nand U11399 (N_11399,N_11174,N_11079);
nand U11400 (N_11400,N_10974,N_10801);
xor U11401 (N_11401,N_10842,N_11109);
xor U11402 (N_11402,N_10910,N_11100);
and U11403 (N_11403,N_11159,N_10894);
or U11404 (N_11404,N_11191,N_10990);
xnor U11405 (N_11405,N_10827,N_10874);
and U11406 (N_11406,N_10987,N_11010);
nor U11407 (N_11407,N_11110,N_10824);
nor U11408 (N_11408,N_10844,N_10955);
and U11409 (N_11409,N_10844,N_11061);
and U11410 (N_11410,N_10826,N_10904);
xor U11411 (N_11411,N_11065,N_10884);
nor U11412 (N_11412,N_11108,N_11084);
and U11413 (N_11413,N_11119,N_10821);
or U11414 (N_11414,N_11172,N_10972);
nor U11415 (N_11415,N_10868,N_10961);
and U11416 (N_11416,N_11184,N_10847);
nand U11417 (N_11417,N_10950,N_11184);
xor U11418 (N_11418,N_10948,N_11079);
or U11419 (N_11419,N_10899,N_11190);
nor U11420 (N_11420,N_10809,N_11060);
nor U11421 (N_11421,N_11108,N_11058);
and U11422 (N_11422,N_10828,N_10940);
or U11423 (N_11423,N_11170,N_11063);
xor U11424 (N_11424,N_10892,N_10846);
nand U11425 (N_11425,N_11117,N_11148);
nand U11426 (N_11426,N_10963,N_11163);
nand U11427 (N_11427,N_10849,N_10898);
or U11428 (N_11428,N_10868,N_10939);
and U11429 (N_11429,N_10984,N_11017);
xor U11430 (N_11430,N_11130,N_11003);
and U11431 (N_11431,N_11197,N_11079);
and U11432 (N_11432,N_11110,N_10916);
nor U11433 (N_11433,N_10930,N_11129);
nand U11434 (N_11434,N_11112,N_10900);
nand U11435 (N_11435,N_11132,N_11101);
nand U11436 (N_11436,N_10965,N_10882);
nand U11437 (N_11437,N_10801,N_10972);
nor U11438 (N_11438,N_11187,N_11094);
or U11439 (N_11439,N_11074,N_11103);
or U11440 (N_11440,N_10974,N_10926);
xnor U11441 (N_11441,N_11144,N_11124);
or U11442 (N_11442,N_11067,N_10887);
nand U11443 (N_11443,N_10983,N_10864);
or U11444 (N_11444,N_11153,N_10939);
xor U11445 (N_11445,N_10805,N_11010);
or U11446 (N_11446,N_10864,N_10883);
and U11447 (N_11447,N_10990,N_11192);
or U11448 (N_11448,N_11056,N_10970);
nor U11449 (N_11449,N_10810,N_10808);
nand U11450 (N_11450,N_10804,N_11027);
nand U11451 (N_11451,N_10828,N_10963);
nand U11452 (N_11452,N_11156,N_11071);
nor U11453 (N_11453,N_11096,N_10869);
or U11454 (N_11454,N_10974,N_10863);
nor U11455 (N_11455,N_11040,N_11131);
xor U11456 (N_11456,N_10852,N_11131);
and U11457 (N_11457,N_11166,N_10952);
xor U11458 (N_11458,N_10949,N_11174);
nand U11459 (N_11459,N_11184,N_10908);
xor U11460 (N_11460,N_11132,N_11127);
nand U11461 (N_11461,N_11132,N_11146);
nor U11462 (N_11462,N_10875,N_11120);
or U11463 (N_11463,N_10850,N_11055);
xnor U11464 (N_11464,N_10966,N_11039);
xor U11465 (N_11465,N_11165,N_10995);
and U11466 (N_11466,N_10960,N_11130);
and U11467 (N_11467,N_11182,N_11147);
nand U11468 (N_11468,N_11126,N_11155);
nor U11469 (N_11469,N_10897,N_10815);
xnor U11470 (N_11470,N_10807,N_11174);
xnor U11471 (N_11471,N_10927,N_10953);
or U11472 (N_11472,N_11012,N_10917);
nor U11473 (N_11473,N_11190,N_10859);
nand U11474 (N_11474,N_10803,N_11010);
or U11475 (N_11475,N_10887,N_10912);
nor U11476 (N_11476,N_10855,N_10810);
or U11477 (N_11477,N_11150,N_10851);
nand U11478 (N_11478,N_11121,N_11110);
or U11479 (N_11479,N_11112,N_11174);
xnor U11480 (N_11480,N_11170,N_10970);
or U11481 (N_11481,N_10961,N_11127);
or U11482 (N_11482,N_11055,N_10903);
or U11483 (N_11483,N_10865,N_11170);
nand U11484 (N_11484,N_10867,N_10821);
nor U11485 (N_11485,N_10836,N_10936);
nor U11486 (N_11486,N_10996,N_11167);
nand U11487 (N_11487,N_11135,N_10940);
nor U11488 (N_11488,N_11181,N_11044);
or U11489 (N_11489,N_10899,N_11183);
nor U11490 (N_11490,N_11089,N_10922);
xor U11491 (N_11491,N_11065,N_10826);
and U11492 (N_11492,N_11145,N_10839);
nand U11493 (N_11493,N_10843,N_11111);
nand U11494 (N_11494,N_10926,N_10888);
xnor U11495 (N_11495,N_10847,N_10803);
and U11496 (N_11496,N_10864,N_11198);
or U11497 (N_11497,N_10810,N_11066);
nand U11498 (N_11498,N_10999,N_11019);
nor U11499 (N_11499,N_10947,N_10995);
xor U11500 (N_11500,N_10891,N_10880);
nand U11501 (N_11501,N_11087,N_10956);
and U11502 (N_11502,N_11028,N_11100);
nand U11503 (N_11503,N_10895,N_10943);
or U11504 (N_11504,N_10922,N_11023);
nand U11505 (N_11505,N_10861,N_11157);
nand U11506 (N_11506,N_11170,N_10987);
and U11507 (N_11507,N_11107,N_11064);
nand U11508 (N_11508,N_10987,N_10861);
nand U11509 (N_11509,N_10927,N_10855);
or U11510 (N_11510,N_11138,N_11024);
or U11511 (N_11511,N_10922,N_11170);
xor U11512 (N_11512,N_11061,N_11010);
and U11513 (N_11513,N_10965,N_11050);
xnor U11514 (N_11514,N_10945,N_10920);
and U11515 (N_11515,N_10811,N_10901);
nand U11516 (N_11516,N_10981,N_11114);
xor U11517 (N_11517,N_10809,N_10947);
or U11518 (N_11518,N_10861,N_10967);
nor U11519 (N_11519,N_11105,N_10871);
nor U11520 (N_11520,N_11077,N_10805);
and U11521 (N_11521,N_10815,N_11082);
or U11522 (N_11522,N_11152,N_10931);
or U11523 (N_11523,N_10900,N_10808);
nand U11524 (N_11524,N_10934,N_10848);
or U11525 (N_11525,N_10808,N_11048);
nor U11526 (N_11526,N_11040,N_10842);
xnor U11527 (N_11527,N_10970,N_11023);
nor U11528 (N_11528,N_10832,N_11195);
or U11529 (N_11529,N_11075,N_11094);
or U11530 (N_11530,N_10919,N_11099);
xnor U11531 (N_11531,N_11044,N_10911);
nor U11532 (N_11532,N_10886,N_10977);
and U11533 (N_11533,N_11020,N_11071);
nor U11534 (N_11534,N_10939,N_11023);
or U11535 (N_11535,N_10836,N_11155);
and U11536 (N_11536,N_10979,N_11109);
and U11537 (N_11537,N_11066,N_10970);
nand U11538 (N_11538,N_10868,N_11169);
xor U11539 (N_11539,N_10956,N_11017);
nand U11540 (N_11540,N_10943,N_10873);
xnor U11541 (N_11541,N_11075,N_10949);
nor U11542 (N_11542,N_10940,N_10954);
xnor U11543 (N_11543,N_11041,N_10804);
xnor U11544 (N_11544,N_11119,N_10801);
xor U11545 (N_11545,N_10851,N_11008);
nor U11546 (N_11546,N_11139,N_10899);
and U11547 (N_11547,N_11146,N_10903);
nor U11548 (N_11548,N_11120,N_10910);
nor U11549 (N_11549,N_11047,N_10844);
or U11550 (N_11550,N_10945,N_10952);
or U11551 (N_11551,N_11058,N_11021);
nand U11552 (N_11552,N_11079,N_11082);
nor U11553 (N_11553,N_10906,N_10892);
or U11554 (N_11554,N_10989,N_10881);
and U11555 (N_11555,N_11079,N_11156);
or U11556 (N_11556,N_10893,N_11117);
xor U11557 (N_11557,N_11018,N_10944);
nor U11558 (N_11558,N_11103,N_11014);
or U11559 (N_11559,N_10899,N_10850);
nand U11560 (N_11560,N_11002,N_11143);
nand U11561 (N_11561,N_11039,N_11195);
nor U11562 (N_11562,N_11013,N_10887);
nor U11563 (N_11563,N_11058,N_10842);
nand U11564 (N_11564,N_11076,N_10871);
or U11565 (N_11565,N_10924,N_10907);
nand U11566 (N_11566,N_11148,N_11196);
nand U11567 (N_11567,N_10874,N_10850);
nand U11568 (N_11568,N_10963,N_10942);
and U11569 (N_11569,N_10948,N_10995);
nand U11570 (N_11570,N_10925,N_10824);
or U11571 (N_11571,N_10902,N_11024);
or U11572 (N_11572,N_10838,N_11001);
xor U11573 (N_11573,N_10927,N_10894);
and U11574 (N_11574,N_10880,N_10951);
xnor U11575 (N_11575,N_10981,N_10942);
nor U11576 (N_11576,N_11008,N_11081);
or U11577 (N_11577,N_11160,N_11120);
xor U11578 (N_11578,N_10871,N_10914);
or U11579 (N_11579,N_11121,N_11067);
nor U11580 (N_11580,N_10872,N_10960);
and U11581 (N_11581,N_11178,N_11082);
and U11582 (N_11582,N_11016,N_11149);
or U11583 (N_11583,N_11139,N_11145);
xnor U11584 (N_11584,N_11085,N_10834);
or U11585 (N_11585,N_11063,N_11015);
nand U11586 (N_11586,N_11199,N_10893);
nand U11587 (N_11587,N_10860,N_11180);
xor U11588 (N_11588,N_10972,N_11092);
and U11589 (N_11589,N_11012,N_10935);
xor U11590 (N_11590,N_10834,N_10840);
nand U11591 (N_11591,N_10989,N_11086);
or U11592 (N_11592,N_11167,N_11033);
nand U11593 (N_11593,N_11061,N_11121);
or U11594 (N_11594,N_11022,N_11055);
xor U11595 (N_11595,N_11070,N_10844);
and U11596 (N_11596,N_10969,N_10877);
xor U11597 (N_11597,N_10810,N_10986);
and U11598 (N_11598,N_11072,N_10922);
nor U11599 (N_11599,N_11076,N_10863);
nor U11600 (N_11600,N_11310,N_11207);
or U11601 (N_11601,N_11576,N_11364);
xnor U11602 (N_11602,N_11373,N_11340);
and U11603 (N_11603,N_11468,N_11586);
and U11604 (N_11604,N_11551,N_11553);
nand U11605 (N_11605,N_11360,N_11477);
nand U11606 (N_11606,N_11270,N_11287);
nor U11607 (N_11607,N_11429,N_11495);
and U11608 (N_11608,N_11474,N_11302);
and U11609 (N_11609,N_11434,N_11314);
and U11610 (N_11610,N_11325,N_11408);
nor U11611 (N_11611,N_11463,N_11464);
or U11612 (N_11612,N_11331,N_11417);
nor U11613 (N_11613,N_11354,N_11459);
and U11614 (N_11614,N_11515,N_11562);
or U11615 (N_11615,N_11232,N_11220);
xnor U11616 (N_11616,N_11432,N_11573);
nand U11617 (N_11617,N_11279,N_11595);
and U11618 (N_11618,N_11560,N_11520);
and U11619 (N_11619,N_11358,N_11554);
and U11620 (N_11620,N_11561,N_11473);
or U11621 (N_11621,N_11536,N_11484);
or U11622 (N_11622,N_11469,N_11456);
nor U11623 (N_11623,N_11260,N_11206);
and U11624 (N_11624,N_11221,N_11276);
nand U11625 (N_11625,N_11457,N_11303);
nand U11626 (N_11626,N_11203,N_11443);
or U11627 (N_11627,N_11513,N_11357);
nand U11628 (N_11628,N_11581,N_11308);
nand U11629 (N_11629,N_11394,N_11215);
and U11630 (N_11630,N_11379,N_11284);
nand U11631 (N_11631,N_11478,N_11324);
nand U11632 (N_11632,N_11508,N_11346);
xnor U11633 (N_11633,N_11307,N_11524);
or U11634 (N_11634,N_11568,N_11572);
and U11635 (N_11635,N_11589,N_11280);
or U11636 (N_11636,N_11476,N_11413);
and U11637 (N_11637,N_11248,N_11363);
nand U11638 (N_11638,N_11405,N_11541);
nand U11639 (N_11639,N_11272,N_11306);
nand U11640 (N_11640,N_11555,N_11202);
nor U11641 (N_11641,N_11522,N_11317);
nor U11642 (N_11642,N_11288,N_11256);
or U11643 (N_11643,N_11311,N_11483);
or U11644 (N_11644,N_11503,N_11448);
or U11645 (N_11645,N_11367,N_11506);
or U11646 (N_11646,N_11492,N_11430);
nor U11647 (N_11647,N_11359,N_11226);
nor U11648 (N_11648,N_11374,N_11205);
xor U11649 (N_11649,N_11519,N_11234);
nand U11650 (N_11650,N_11332,N_11337);
or U11651 (N_11651,N_11537,N_11558);
nor U11652 (N_11652,N_11548,N_11438);
or U11653 (N_11653,N_11444,N_11209);
and U11654 (N_11654,N_11592,N_11404);
xor U11655 (N_11655,N_11428,N_11542);
xnor U11656 (N_11656,N_11339,N_11391);
nor U11657 (N_11657,N_11538,N_11570);
or U11658 (N_11658,N_11333,N_11222);
nand U11659 (N_11659,N_11294,N_11588);
xor U11660 (N_11660,N_11285,N_11265);
xor U11661 (N_11661,N_11295,N_11275);
or U11662 (N_11662,N_11262,N_11435);
nand U11663 (N_11663,N_11267,N_11253);
or U11664 (N_11664,N_11535,N_11461);
xor U11665 (N_11665,N_11403,N_11458);
or U11666 (N_11666,N_11312,N_11296);
xnor U11667 (N_11667,N_11216,N_11552);
xnor U11668 (N_11668,N_11425,N_11351);
or U11669 (N_11669,N_11406,N_11534);
nand U11670 (N_11670,N_11224,N_11309);
or U11671 (N_11671,N_11366,N_11300);
or U11672 (N_11672,N_11349,N_11517);
xor U11673 (N_11673,N_11590,N_11439);
nand U11674 (N_11674,N_11424,N_11345);
or U11675 (N_11675,N_11482,N_11236);
and U11676 (N_11676,N_11584,N_11489);
nand U11677 (N_11677,N_11242,N_11328);
nor U11678 (N_11678,N_11329,N_11286);
xor U11679 (N_11679,N_11200,N_11269);
xnor U11680 (N_11680,N_11578,N_11436);
or U11681 (N_11681,N_11460,N_11211);
xor U11682 (N_11682,N_11263,N_11399);
nand U11683 (N_11683,N_11250,N_11208);
nor U11684 (N_11684,N_11481,N_11420);
nand U11685 (N_11685,N_11575,N_11313);
or U11686 (N_11686,N_11237,N_11227);
nor U11687 (N_11687,N_11433,N_11490);
nor U11688 (N_11688,N_11598,N_11247);
xnor U11689 (N_11689,N_11543,N_11368);
nor U11690 (N_11690,N_11421,N_11496);
xor U11691 (N_11691,N_11377,N_11529);
nor U11692 (N_11692,N_11422,N_11545);
or U11693 (N_11693,N_11334,N_11344);
nor U11694 (N_11694,N_11471,N_11264);
nand U11695 (N_11695,N_11564,N_11240);
and U11696 (N_11696,N_11229,N_11501);
and U11697 (N_11697,N_11557,N_11283);
xor U11698 (N_11698,N_11450,N_11365);
and U11699 (N_11699,N_11383,N_11585);
or U11700 (N_11700,N_11418,N_11583);
xor U11701 (N_11701,N_11494,N_11566);
nand U11702 (N_11702,N_11382,N_11277);
xor U11703 (N_11703,N_11293,N_11204);
and U11704 (N_11704,N_11423,N_11480);
nand U11705 (N_11705,N_11514,N_11335);
xor U11706 (N_11706,N_11577,N_11245);
or U11707 (N_11707,N_11441,N_11225);
nand U11708 (N_11708,N_11518,N_11390);
and U11709 (N_11709,N_11510,N_11246);
or U11710 (N_11710,N_11531,N_11466);
or U11711 (N_11711,N_11493,N_11449);
nand U11712 (N_11712,N_11350,N_11451);
and U11713 (N_11713,N_11526,N_11402);
or U11714 (N_11714,N_11321,N_11305);
or U11715 (N_11715,N_11252,N_11453);
nor U11716 (N_11716,N_11559,N_11378);
xnor U11717 (N_11717,N_11393,N_11580);
or U11718 (N_11718,N_11292,N_11231);
nand U11719 (N_11719,N_11330,N_11593);
or U11720 (N_11720,N_11352,N_11411);
or U11721 (N_11721,N_11326,N_11223);
nor U11722 (N_11722,N_11348,N_11228);
xor U11723 (N_11723,N_11485,N_11255);
nor U11724 (N_11724,N_11249,N_11319);
and U11725 (N_11725,N_11271,N_11426);
nand U11726 (N_11726,N_11392,N_11497);
xnor U11727 (N_11727,N_11230,N_11353);
or U11728 (N_11728,N_11452,N_11546);
nor U11729 (N_11729,N_11504,N_11338);
or U11730 (N_11730,N_11597,N_11210);
nor U11731 (N_11731,N_11596,N_11316);
xnor U11732 (N_11732,N_11437,N_11251);
and U11733 (N_11733,N_11266,N_11454);
or U11734 (N_11734,N_11407,N_11574);
and U11735 (N_11735,N_11387,N_11530);
and U11736 (N_11736,N_11419,N_11445);
and U11737 (N_11737,N_11475,N_11516);
nand U11738 (N_11738,N_11258,N_11239);
xnor U11739 (N_11739,N_11376,N_11487);
and U11740 (N_11740,N_11395,N_11582);
nand U11741 (N_11741,N_11509,N_11323);
nor U11742 (N_11742,N_11362,N_11322);
and U11743 (N_11743,N_11278,N_11488);
and U11744 (N_11744,N_11217,N_11442);
nor U11745 (N_11745,N_11401,N_11289);
or U11746 (N_11746,N_11355,N_11571);
nand U11747 (N_11747,N_11298,N_11533);
nor U11748 (N_11748,N_11290,N_11261);
nand U11749 (N_11749,N_11274,N_11369);
nand U11750 (N_11750,N_11385,N_11455);
nor U11751 (N_11751,N_11505,N_11491);
nand U11752 (N_11752,N_11238,N_11257);
or U11753 (N_11753,N_11507,N_11268);
nand U11754 (N_11754,N_11465,N_11315);
or U11755 (N_11755,N_11472,N_11549);
xor U11756 (N_11756,N_11372,N_11587);
or U11757 (N_11757,N_11414,N_11281);
or U11758 (N_11758,N_11219,N_11569);
nor U11759 (N_11759,N_11381,N_11591);
xor U11760 (N_11760,N_11299,N_11389);
xor U11761 (N_11761,N_11400,N_11282);
nand U11762 (N_11762,N_11525,N_11498);
xnor U11763 (N_11763,N_11579,N_11427);
or U11764 (N_11764,N_11336,N_11341);
xnor U11765 (N_11765,N_11233,N_11467);
or U11766 (N_11766,N_11447,N_11327);
nor U11767 (N_11767,N_11479,N_11599);
or U11768 (N_11768,N_11241,N_11567);
nand U11769 (N_11769,N_11214,N_11556);
or U11770 (N_11770,N_11547,N_11540);
nor U11771 (N_11771,N_11462,N_11244);
or U11772 (N_11772,N_11259,N_11254);
nor U11773 (N_11773,N_11396,N_11410);
nor U11774 (N_11774,N_11297,N_11386);
or U11775 (N_11775,N_11502,N_11594);
nand U11776 (N_11776,N_11235,N_11342);
or U11777 (N_11777,N_11565,N_11213);
and U11778 (N_11778,N_11500,N_11415);
xor U11779 (N_11779,N_11212,N_11243);
or U11780 (N_11780,N_11370,N_11563);
or U11781 (N_11781,N_11440,N_11318);
nor U11782 (N_11782,N_11550,N_11347);
nand U11783 (N_11783,N_11539,N_11343);
or U11784 (N_11784,N_11416,N_11499);
nor U11785 (N_11785,N_11320,N_11397);
xor U11786 (N_11786,N_11528,N_11201);
xnor U11787 (N_11787,N_11356,N_11523);
nor U11788 (N_11788,N_11511,N_11521);
or U11789 (N_11789,N_11375,N_11512);
nand U11790 (N_11790,N_11361,N_11527);
nand U11791 (N_11791,N_11398,N_11384);
and U11792 (N_11792,N_11301,N_11486);
nand U11793 (N_11793,N_11380,N_11446);
nand U11794 (N_11794,N_11218,N_11291);
or U11795 (N_11795,N_11388,N_11544);
xor U11796 (N_11796,N_11470,N_11409);
nor U11797 (N_11797,N_11273,N_11371);
nand U11798 (N_11798,N_11431,N_11532);
nor U11799 (N_11799,N_11412,N_11304);
or U11800 (N_11800,N_11468,N_11476);
nor U11801 (N_11801,N_11360,N_11314);
nand U11802 (N_11802,N_11561,N_11528);
xnor U11803 (N_11803,N_11241,N_11381);
xnor U11804 (N_11804,N_11328,N_11577);
and U11805 (N_11805,N_11549,N_11338);
and U11806 (N_11806,N_11327,N_11528);
or U11807 (N_11807,N_11291,N_11585);
or U11808 (N_11808,N_11541,N_11576);
nand U11809 (N_11809,N_11304,N_11597);
nor U11810 (N_11810,N_11455,N_11237);
or U11811 (N_11811,N_11563,N_11545);
xnor U11812 (N_11812,N_11224,N_11263);
and U11813 (N_11813,N_11546,N_11369);
nand U11814 (N_11814,N_11240,N_11238);
xor U11815 (N_11815,N_11432,N_11277);
and U11816 (N_11816,N_11501,N_11398);
xor U11817 (N_11817,N_11320,N_11500);
or U11818 (N_11818,N_11586,N_11487);
nand U11819 (N_11819,N_11244,N_11214);
and U11820 (N_11820,N_11340,N_11284);
nor U11821 (N_11821,N_11506,N_11411);
nor U11822 (N_11822,N_11434,N_11514);
xor U11823 (N_11823,N_11451,N_11473);
and U11824 (N_11824,N_11293,N_11350);
nor U11825 (N_11825,N_11353,N_11452);
and U11826 (N_11826,N_11474,N_11563);
or U11827 (N_11827,N_11347,N_11395);
or U11828 (N_11828,N_11355,N_11540);
or U11829 (N_11829,N_11305,N_11275);
and U11830 (N_11830,N_11416,N_11236);
xnor U11831 (N_11831,N_11252,N_11541);
and U11832 (N_11832,N_11509,N_11248);
xor U11833 (N_11833,N_11558,N_11241);
nor U11834 (N_11834,N_11394,N_11450);
nand U11835 (N_11835,N_11527,N_11596);
nand U11836 (N_11836,N_11200,N_11399);
or U11837 (N_11837,N_11363,N_11204);
nor U11838 (N_11838,N_11357,N_11294);
or U11839 (N_11839,N_11260,N_11453);
or U11840 (N_11840,N_11567,N_11476);
nand U11841 (N_11841,N_11490,N_11210);
and U11842 (N_11842,N_11446,N_11213);
xnor U11843 (N_11843,N_11524,N_11563);
nor U11844 (N_11844,N_11581,N_11240);
xor U11845 (N_11845,N_11436,N_11569);
nor U11846 (N_11846,N_11504,N_11254);
or U11847 (N_11847,N_11263,N_11221);
nor U11848 (N_11848,N_11411,N_11536);
and U11849 (N_11849,N_11549,N_11548);
nor U11850 (N_11850,N_11586,N_11429);
nor U11851 (N_11851,N_11434,N_11443);
or U11852 (N_11852,N_11291,N_11409);
or U11853 (N_11853,N_11272,N_11508);
or U11854 (N_11854,N_11205,N_11254);
nor U11855 (N_11855,N_11419,N_11214);
nor U11856 (N_11856,N_11485,N_11233);
nor U11857 (N_11857,N_11343,N_11395);
and U11858 (N_11858,N_11235,N_11307);
or U11859 (N_11859,N_11459,N_11311);
xor U11860 (N_11860,N_11404,N_11584);
xnor U11861 (N_11861,N_11424,N_11582);
nor U11862 (N_11862,N_11375,N_11344);
xor U11863 (N_11863,N_11247,N_11483);
nor U11864 (N_11864,N_11512,N_11580);
nand U11865 (N_11865,N_11202,N_11551);
nand U11866 (N_11866,N_11238,N_11232);
nor U11867 (N_11867,N_11487,N_11288);
or U11868 (N_11868,N_11404,N_11272);
or U11869 (N_11869,N_11392,N_11268);
nand U11870 (N_11870,N_11514,N_11294);
and U11871 (N_11871,N_11390,N_11294);
and U11872 (N_11872,N_11537,N_11361);
nor U11873 (N_11873,N_11454,N_11432);
nor U11874 (N_11874,N_11593,N_11578);
xor U11875 (N_11875,N_11214,N_11243);
xnor U11876 (N_11876,N_11384,N_11578);
nor U11877 (N_11877,N_11559,N_11514);
nand U11878 (N_11878,N_11431,N_11566);
or U11879 (N_11879,N_11479,N_11398);
or U11880 (N_11880,N_11294,N_11274);
nand U11881 (N_11881,N_11240,N_11475);
xor U11882 (N_11882,N_11492,N_11270);
nor U11883 (N_11883,N_11483,N_11538);
xor U11884 (N_11884,N_11550,N_11407);
nor U11885 (N_11885,N_11512,N_11503);
and U11886 (N_11886,N_11400,N_11268);
nand U11887 (N_11887,N_11437,N_11431);
nor U11888 (N_11888,N_11504,N_11284);
nand U11889 (N_11889,N_11350,N_11461);
and U11890 (N_11890,N_11301,N_11227);
or U11891 (N_11891,N_11494,N_11241);
nand U11892 (N_11892,N_11446,N_11241);
nand U11893 (N_11893,N_11324,N_11415);
and U11894 (N_11894,N_11368,N_11557);
nand U11895 (N_11895,N_11336,N_11474);
nor U11896 (N_11896,N_11360,N_11320);
xnor U11897 (N_11897,N_11383,N_11319);
nand U11898 (N_11898,N_11274,N_11523);
nor U11899 (N_11899,N_11273,N_11292);
xor U11900 (N_11900,N_11273,N_11468);
xnor U11901 (N_11901,N_11267,N_11264);
or U11902 (N_11902,N_11597,N_11301);
or U11903 (N_11903,N_11460,N_11429);
nor U11904 (N_11904,N_11369,N_11440);
and U11905 (N_11905,N_11468,N_11404);
xor U11906 (N_11906,N_11409,N_11205);
nand U11907 (N_11907,N_11330,N_11546);
and U11908 (N_11908,N_11315,N_11473);
or U11909 (N_11909,N_11543,N_11362);
and U11910 (N_11910,N_11346,N_11398);
nand U11911 (N_11911,N_11354,N_11222);
and U11912 (N_11912,N_11314,N_11553);
nand U11913 (N_11913,N_11562,N_11307);
nand U11914 (N_11914,N_11566,N_11564);
nor U11915 (N_11915,N_11453,N_11470);
xnor U11916 (N_11916,N_11420,N_11472);
or U11917 (N_11917,N_11338,N_11410);
nand U11918 (N_11918,N_11328,N_11390);
nand U11919 (N_11919,N_11453,N_11265);
xor U11920 (N_11920,N_11255,N_11274);
nor U11921 (N_11921,N_11220,N_11329);
nand U11922 (N_11922,N_11211,N_11221);
nand U11923 (N_11923,N_11433,N_11370);
nand U11924 (N_11924,N_11285,N_11453);
nor U11925 (N_11925,N_11484,N_11317);
or U11926 (N_11926,N_11589,N_11424);
xor U11927 (N_11927,N_11392,N_11482);
xor U11928 (N_11928,N_11313,N_11478);
nand U11929 (N_11929,N_11260,N_11310);
nand U11930 (N_11930,N_11462,N_11429);
nand U11931 (N_11931,N_11299,N_11388);
nor U11932 (N_11932,N_11583,N_11386);
nand U11933 (N_11933,N_11394,N_11281);
xor U11934 (N_11934,N_11553,N_11273);
xor U11935 (N_11935,N_11459,N_11370);
nor U11936 (N_11936,N_11336,N_11268);
nand U11937 (N_11937,N_11516,N_11514);
nor U11938 (N_11938,N_11342,N_11272);
nor U11939 (N_11939,N_11522,N_11431);
and U11940 (N_11940,N_11342,N_11460);
or U11941 (N_11941,N_11537,N_11329);
nor U11942 (N_11942,N_11335,N_11431);
nor U11943 (N_11943,N_11409,N_11222);
nor U11944 (N_11944,N_11446,N_11455);
xor U11945 (N_11945,N_11418,N_11448);
xnor U11946 (N_11946,N_11576,N_11334);
xor U11947 (N_11947,N_11540,N_11557);
nor U11948 (N_11948,N_11286,N_11455);
or U11949 (N_11949,N_11480,N_11333);
or U11950 (N_11950,N_11226,N_11347);
or U11951 (N_11951,N_11503,N_11584);
nand U11952 (N_11952,N_11310,N_11599);
nand U11953 (N_11953,N_11229,N_11584);
xor U11954 (N_11954,N_11363,N_11509);
nand U11955 (N_11955,N_11312,N_11574);
xnor U11956 (N_11956,N_11214,N_11346);
nand U11957 (N_11957,N_11246,N_11406);
or U11958 (N_11958,N_11591,N_11222);
and U11959 (N_11959,N_11303,N_11284);
nand U11960 (N_11960,N_11405,N_11287);
and U11961 (N_11961,N_11524,N_11522);
xnor U11962 (N_11962,N_11435,N_11388);
xor U11963 (N_11963,N_11447,N_11232);
xnor U11964 (N_11964,N_11443,N_11401);
or U11965 (N_11965,N_11565,N_11575);
and U11966 (N_11966,N_11266,N_11317);
xor U11967 (N_11967,N_11279,N_11319);
xnor U11968 (N_11968,N_11325,N_11238);
nand U11969 (N_11969,N_11346,N_11334);
nand U11970 (N_11970,N_11381,N_11454);
and U11971 (N_11971,N_11525,N_11489);
nor U11972 (N_11972,N_11341,N_11322);
or U11973 (N_11973,N_11395,N_11541);
or U11974 (N_11974,N_11341,N_11580);
nand U11975 (N_11975,N_11477,N_11224);
nand U11976 (N_11976,N_11265,N_11537);
xor U11977 (N_11977,N_11446,N_11457);
xnor U11978 (N_11978,N_11323,N_11246);
or U11979 (N_11979,N_11210,N_11295);
nor U11980 (N_11980,N_11504,N_11239);
and U11981 (N_11981,N_11421,N_11491);
xnor U11982 (N_11982,N_11527,N_11417);
nor U11983 (N_11983,N_11213,N_11539);
nor U11984 (N_11984,N_11599,N_11278);
nor U11985 (N_11985,N_11303,N_11578);
xnor U11986 (N_11986,N_11524,N_11575);
nor U11987 (N_11987,N_11463,N_11551);
or U11988 (N_11988,N_11339,N_11555);
nand U11989 (N_11989,N_11240,N_11297);
and U11990 (N_11990,N_11415,N_11389);
nor U11991 (N_11991,N_11469,N_11246);
nand U11992 (N_11992,N_11397,N_11469);
xnor U11993 (N_11993,N_11279,N_11529);
or U11994 (N_11994,N_11468,N_11446);
xnor U11995 (N_11995,N_11523,N_11520);
nand U11996 (N_11996,N_11424,N_11231);
or U11997 (N_11997,N_11385,N_11592);
or U11998 (N_11998,N_11592,N_11595);
and U11999 (N_11999,N_11337,N_11382);
and U12000 (N_12000,N_11658,N_11681);
xor U12001 (N_12001,N_11627,N_11939);
nand U12002 (N_12002,N_11840,N_11867);
nand U12003 (N_12003,N_11978,N_11736);
xor U12004 (N_12004,N_11609,N_11755);
or U12005 (N_12005,N_11733,N_11885);
or U12006 (N_12006,N_11941,N_11706);
and U12007 (N_12007,N_11969,N_11710);
nor U12008 (N_12008,N_11955,N_11954);
nor U12009 (N_12009,N_11964,N_11783);
and U12010 (N_12010,N_11652,N_11817);
nand U12011 (N_12011,N_11811,N_11704);
or U12012 (N_12012,N_11945,N_11775);
nor U12013 (N_12013,N_11953,N_11604);
nor U12014 (N_12014,N_11639,N_11768);
xor U12015 (N_12015,N_11937,N_11661);
or U12016 (N_12016,N_11654,N_11726);
and U12017 (N_12017,N_11801,N_11684);
xor U12018 (N_12018,N_11715,N_11643);
and U12019 (N_12019,N_11624,N_11669);
and U12020 (N_12020,N_11679,N_11788);
nand U12021 (N_12021,N_11838,N_11961);
or U12022 (N_12022,N_11799,N_11952);
or U12023 (N_12023,N_11901,N_11996);
nor U12024 (N_12024,N_11816,N_11724);
and U12025 (N_12025,N_11997,N_11748);
nor U12026 (N_12026,N_11687,N_11855);
nand U12027 (N_12027,N_11921,N_11957);
and U12028 (N_12028,N_11730,N_11894);
nand U12029 (N_12029,N_11820,N_11908);
or U12030 (N_12030,N_11998,N_11888);
or U12031 (N_12031,N_11649,N_11686);
xor U12032 (N_12032,N_11739,N_11932);
nand U12033 (N_12033,N_11902,N_11980);
xor U12034 (N_12034,N_11823,N_11930);
nand U12035 (N_12035,N_11727,N_11712);
xor U12036 (N_12036,N_11662,N_11965);
or U12037 (N_12037,N_11707,N_11640);
nand U12038 (N_12038,N_11812,N_11729);
xor U12039 (N_12039,N_11903,N_11814);
nor U12040 (N_12040,N_11762,N_11860);
or U12041 (N_12041,N_11815,N_11972);
and U12042 (N_12042,N_11784,N_11803);
and U12043 (N_12043,N_11914,N_11895);
nand U12044 (N_12044,N_11950,N_11942);
nor U12045 (N_12045,N_11636,N_11844);
nor U12046 (N_12046,N_11725,N_11990);
xnor U12047 (N_12047,N_11847,N_11618);
xor U12048 (N_12048,N_11878,N_11805);
xnor U12049 (N_12049,N_11738,N_11906);
or U12050 (N_12050,N_11656,N_11674);
or U12051 (N_12051,N_11882,N_11778);
nor U12052 (N_12052,N_11787,N_11759);
nand U12053 (N_12053,N_11833,N_11923);
or U12054 (N_12054,N_11832,N_11623);
nor U12055 (N_12055,N_11920,N_11830);
nor U12056 (N_12056,N_11771,N_11826);
and U12057 (N_12057,N_11737,N_11743);
nor U12058 (N_12058,N_11837,N_11986);
xnor U12059 (N_12059,N_11602,N_11863);
nor U12060 (N_12060,N_11880,N_11796);
or U12061 (N_12061,N_11849,N_11819);
or U12062 (N_12062,N_11946,N_11963);
xnor U12063 (N_12063,N_11936,N_11807);
nor U12064 (N_12064,N_11716,N_11827);
nor U12065 (N_12065,N_11657,N_11971);
nand U12066 (N_12066,N_11696,N_11790);
nand U12067 (N_12067,N_11839,N_11958);
and U12068 (N_12068,N_11747,N_11977);
and U12069 (N_12069,N_11646,N_11852);
and U12070 (N_12070,N_11678,N_11776);
and U12071 (N_12071,N_11718,N_11723);
or U12072 (N_12072,N_11612,N_11850);
nand U12073 (N_12073,N_11644,N_11795);
nand U12074 (N_12074,N_11813,N_11667);
or U12075 (N_12075,N_11872,N_11992);
nand U12076 (N_12076,N_11810,N_11608);
nor U12077 (N_12077,N_11959,N_11628);
or U12078 (N_12078,N_11632,N_11853);
nor U12079 (N_12079,N_11831,N_11884);
and U12080 (N_12080,N_11846,N_11637);
xnor U12081 (N_12081,N_11960,N_11913);
nand U12082 (N_12082,N_11793,N_11650);
or U12083 (N_12083,N_11655,N_11900);
nand U12084 (N_12084,N_11728,N_11638);
nand U12085 (N_12085,N_11751,N_11754);
or U12086 (N_12086,N_11693,N_11862);
and U12087 (N_12087,N_11717,N_11781);
nor U12088 (N_12088,N_11982,N_11976);
and U12089 (N_12089,N_11621,N_11605);
and U12090 (N_12090,N_11911,N_11734);
xor U12091 (N_12091,N_11848,N_11617);
and U12092 (N_12092,N_11721,N_11917);
and U12093 (N_12093,N_11808,N_11800);
nand U12094 (N_12094,N_11886,N_11794);
xor U12095 (N_12095,N_11896,N_11858);
or U12096 (N_12096,N_11873,N_11987);
or U12097 (N_12097,N_11660,N_11806);
or U12098 (N_12098,N_11984,N_11694);
xnor U12099 (N_12099,N_11635,N_11714);
nor U12100 (N_12100,N_11703,N_11909);
xor U12101 (N_12101,N_11851,N_11887);
nand U12102 (N_12102,N_11782,N_11891);
xnor U12103 (N_12103,N_11672,N_11688);
nand U12104 (N_12104,N_11633,N_11843);
nor U12105 (N_12105,N_11770,N_11933);
and U12106 (N_12106,N_11876,N_11854);
xnor U12107 (N_12107,N_11870,N_11841);
nor U12108 (N_12108,N_11702,N_11857);
and U12109 (N_12109,N_11760,N_11682);
and U12110 (N_12110,N_11993,N_11809);
xor U12111 (N_12111,N_11845,N_11626);
or U12112 (N_12112,N_11645,N_11935);
nand U12113 (N_12113,N_11974,N_11735);
or U12114 (N_12114,N_11699,N_11700);
xnor U12115 (N_12115,N_11777,N_11742);
or U12116 (N_12116,N_11789,N_11629);
xor U12117 (N_12117,N_11619,N_11695);
nand U12118 (N_12118,N_11786,N_11868);
nor U12119 (N_12119,N_11975,N_11666);
nor U12120 (N_12120,N_11692,N_11979);
xnor U12121 (N_12121,N_11607,N_11701);
and U12122 (N_12122,N_11685,N_11916);
and U12123 (N_12123,N_11651,N_11741);
nor U12124 (N_12124,N_11792,N_11749);
and U12125 (N_12125,N_11989,N_11836);
nor U12126 (N_12126,N_11879,N_11865);
nor U12127 (N_12127,N_11670,N_11927);
nor U12128 (N_12128,N_11705,N_11797);
nand U12129 (N_12129,N_11613,N_11708);
or U12130 (N_12130,N_11779,N_11925);
and U12131 (N_12131,N_11606,N_11631);
and U12132 (N_12132,N_11898,N_11664);
xnor U12133 (N_12133,N_11821,N_11892);
nand U12134 (N_12134,N_11949,N_11804);
xnor U12135 (N_12135,N_11859,N_11673);
xnor U12136 (N_12136,N_11765,N_11713);
nand U12137 (N_12137,N_11711,N_11745);
or U12138 (N_12138,N_11889,N_11828);
xor U12139 (N_12139,N_11802,N_11780);
or U12140 (N_12140,N_11610,N_11966);
nand U12141 (N_12141,N_11910,N_11634);
or U12142 (N_12142,N_11983,N_11835);
xor U12143 (N_12143,N_11740,N_11934);
and U12144 (N_12144,N_11697,N_11834);
and U12145 (N_12145,N_11970,N_11616);
or U12146 (N_12146,N_11668,N_11648);
xnor U12147 (N_12147,N_11915,N_11962);
xor U12148 (N_12148,N_11973,N_11818);
or U12149 (N_12149,N_11912,N_11625);
nor U12150 (N_12150,N_11985,N_11659);
nor U12151 (N_12151,N_11791,N_11919);
nor U12152 (N_12152,N_11722,N_11746);
xor U12153 (N_12153,N_11871,N_11922);
nor U12154 (N_12154,N_11647,N_11615);
and U12155 (N_12155,N_11689,N_11956);
nand U12156 (N_12156,N_11905,N_11981);
nand U12157 (N_12157,N_11622,N_11758);
xor U12158 (N_12158,N_11785,N_11603);
or U12159 (N_12159,N_11675,N_11967);
and U12160 (N_12160,N_11928,N_11991);
nand U12161 (N_12161,N_11671,N_11753);
nor U12162 (N_12162,N_11856,N_11732);
xnor U12163 (N_12163,N_11874,N_11774);
xnor U12164 (N_12164,N_11720,N_11630);
nand U12165 (N_12165,N_11951,N_11918);
or U12166 (N_12166,N_11824,N_11829);
or U12167 (N_12167,N_11940,N_11907);
and U12168 (N_12168,N_11798,N_11766);
nor U12169 (N_12169,N_11744,N_11929);
nor U12170 (N_12170,N_11709,N_11769);
or U12171 (N_12171,N_11764,N_11752);
xnor U12172 (N_12172,N_11620,N_11680);
or U12173 (N_12173,N_11881,N_11864);
and U12174 (N_12174,N_11944,N_11825);
nand U12175 (N_12175,N_11676,N_11683);
nand U12176 (N_12176,N_11995,N_11663);
or U12177 (N_12177,N_11968,N_11904);
nand U12178 (N_12178,N_11665,N_11600);
nor U12179 (N_12179,N_11731,N_11877);
nand U12180 (N_12180,N_11822,N_11947);
nor U12181 (N_12181,N_11999,N_11866);
nor U12182 (N_12182,N_11938,N_11767);
xnor U12183 (N_12183,N_11924,N_11948);
xor U12184 (N_12184,N_11601,N_11773);
nand U12185 (N_12185,N_11691,N_11943);
and U12186 (N_12186,N_11890,N_11994);
and U12187 (N_12187,N_11642,N_11750);
xnor U12188 (N_12188,N_11641,N_11861);
or U12189 (N_12189,N_11869,N_11931);
xor U12190 (N_12190,N_11763,N_11897);
and U12191 (N_12191,N_11757,N_11756);
nand U12192 (N_12192,N_11677,N_11719);
nor U12193 (N_12193,N_11772,N_11614);
xor U12194 (N_12194,N_11926,N_11842);
and U12195 (N_12195,N_11883,N_11611);
nand U12196 (N_12196,N_11653,N_11899);
nor U12197 (N_12197,N_11893,N_11761);
and U12198 (N_12198,N_11875,N_11698);
nand U12199 (N_12199,N_11690,N_11988);
xor U12200 (N_12200,N_11743,N_11847);
xnor U12201 (N_12201,N_11780,N_11885);
nand U12202 (N_12202,N_11918,N_11911);
xor U12203 (N_12203,N_11879,N_11823);
nor U12204 (N_12204,N_11650,N_11921);
and U12205 (N_12205,N_11834,N_11947);
or U12206 (N_12206,N_11738,N_11893);
or U12207 (N_12207,N_11814,N_11661);
nand U12208 (N_12208,N_11605,N_11990);
and U12209 (N_12209,N_11791,N_11722);
or U12210 (N_12210,N_11860,N_11792);
nor U12211 (N_12211,N_11777,N_11631);
nor U12212 (N_12212,N_11701,N_11700);
and U12213 (N_12213,N_11987,N_11989);
nand U12214 (N_12214,N_11671,N_11648);
xor U12215 (N_12215,N_11916,N_11721);
and U12216 (N_12216,N_11643,N_11753);
xor U12217 (N_12217,N_11790,N_11700);
or U12218 (N_12218,N_11833,N_11659);
xor U12219 (N_12219,N_11879,N_11971);
or U12220 (N_12220,N_11855,N_11930);
nand U12221 (N_12221,N_11749,N_11686);
xor U12222 (N_12222,N_11889,N_11742);
or U12223 (N_12223,N_11997,N_11623);
xnor U12224 (N_12224,N_11966,N_11699);
or U12225 (N_12225,N_11834,N_11747);
xnor U12226 (N_12226,N_11618,N_11955);
and U12227 (N_12227,N_11895,N_11873);
or U12228 (N_12228,N_11881,N_11823);
nand U12229 (N_12229,N_11642,N_11675);
nand U12230 (N_12230,N_11988,N_11700);
or U12231 (N_12231,N_11847,N_11633);
xnor U12232 (N_12232,N_11610,N_11964);
nor U12233 (N_12233,N_11654,N_11828);
xor U12234 (N_12234,N_11923,N_11691);
or U12235 (N_12235,N_11904,N_11737);
nand U12236 (N_12236,N_11783,N_11729);
nor U12237 (N_12237,N_11948,N_11682);
nor U12238 (N_12238,N_11777,N_11752);
xnor U12239 (N_12239,N_11926,N_11884);
nand U12240 (N_12240,N_11955,N_11720);
xor U12241 (N_12241,N_11682,N_11883);
and U12242 (N_12242,N_11767,N_11890);
or U12243 (N_12243,N_11899,N_11986);
and U12244 (N_12244,N_11829,N_11600);
nor U12245 (N_12245,N_11927,N_11770);
or U12246 (N_12246,N_11987,N_11805);
and U12247 (N_12247,N_11998,N_11844);
and U12248 (N_12248,N_11935,N_11995);
xnor U12249 (N_12249,N_11971,N_11671);
nor U12250 (N_12250,N_11771,N_11618);
nor U12251 (N_12251,N_11609,N_11828);
and U12252 (N_12252,N_11966,N_11934);
nand U12253 (N_12253,N_11827,N_11898);
xnor U12254 (N_12254,N_11813,N_11830);
or U12255 (N_12255,N_11732,N_11726);
nand U12256 (N_12256,N_11832,N_11772);
or U12257 (N_12257,N_11836,N_11840);
or U12258 (N_12258,N_11882,N_11772);
nand U12259 (N_12259,N_11605,N_11678);
xor U12260 (N_12260,N_11832,N_11723);
xnor U12261 (N_12261,N_11951,N_11730);
xnor U12262 (N_12262,N_11979,N_11866);
nand U12263 (N_12263,N_11648,N_11926);
or U12264 (N_12264,N_11751,N_11859);
nand U12265 (N_12265,N_11768,N_11646);
xor U12266 (N_12266,N_11744,N_11885);
or U12267 (N_12267,N_11860,N_11715);
xnor U12268 (N_12268,N_11774,N_11948);
and U12269 (N_12269,N_11954,N_11681);
nor U12270 (N_12270,N_11793,N_11601);
or U12271 (N_12271,N_11804,N_11691);
xor U12272 (N_12272,N_11644,N_11933);
nand U12273 (N_12273,N_11960,N_11901);
and U12274 (N_12274,N_11971,N_11821);
and U12275 (N_12275,N_11877,N_11803);
and U12276 (N_12276,N_11759,N_11778);
xnor U12277 (N_12277,N_11861,N_11954);
or U12278 (N_12278,N_11745,N_11901);
nor U12279 (N_12279,N_11954,N_11948);
and U12280 (N_12280,N_11893,N_11990);
and U12281 (N_12281,N_11602,N_11727);
or U12282 (N_12282,N_11900,N_11777);
nor U12283 (N_12283,N_11860,N_11882);
xor U12284 (N_12284,N_11975,N_11605);
nand U12285 (N_12285,N_11707,N_11663);
or U12286 (N_12286,N_11950,N_11979);
xnor U12287 (N_12287,N_11807,N_11820);
nor U12288 (N_12288,N_11958,N_11933);
xor U12289 (N_12289,N_11732,N_11889);
nor U12290 (N_12290,N_11988,N_11882);
or U12291 (N_12291,N_11656,N_11770);
or U12292 (N_12292,N_11846,N_11819);
or U12293 (N_12293,N_11970,N_11885);
nor U12294 (N_12294,N_11603,N_11934);
xnor U12295 (N_12295,N_11672,N_11703);
xor U12296 (N_12296,N_11689,N_11640);
xnor U12297 (N_12297,N_11840,N_11658);
nand U12298 (N_12298,N_11776,N_11808);
and U12299 (N_12299,N_11846,N_11874);
nand U12300 (N_12300,N_11913,N_11832);
nand U12301 (N_12301,N_11843,N_11815);
or U12302 (N_12302,N_11874,N_11931);
nand U12303 (N_12303,N_11768,N_11701);
xor U12304 (N_12304,N_11899,N_11707);
nor U12305 (N_12305,N_11652,N_11991);
or U12306 (N_12306,N_11733,N_11964);
nand U12307 (N_12307,N_11801,N_11939);
and U12308 (N_12308,N_11771,N_11837);
nand U12309 (N_12309,N_11801,N_11911);
and U12310 (N_12310,N_11974,N_11888);
nand U12311 (N_12311,N_11713,N_11927);
nor U12312 (N_12312,N_11722,N_11676);
or U12313 (N_12313,N_11711,N_11790);
nand U12314 (N_12314,N_11907,N_11800);
or U12315 (N_12315,N_11728,N_11652);
xor U12316 (N_12316,N_11926,N_11814);
or U12317 (N_12317,N_11944,N_11993);
xor U12318 (N_12318,N_11894,N_11967);
nand U12319 (N_12319,N_11830,N_11780);
xnor U12320 (N_12320,N_11990,N_11673);
xnor U12321 (N_12321,N_11905,N_11929);
xnor U12322 (N_12322,N_11720,N_11613);
xor U12323 (N_12323,N_11713,N_11986);
or U12324 (N_12324,N_11803,N_11790);
or U12325 (N_12325,N_11737,N_11908);
and U12326 (N_12326,N_11924,N_11748);
nor U12327 (N_12327,N_11629,N_11732);
and U12328 (N_12328,N_11749,N_11737);
and U12329 (N_12329,N_11834,N_11864);
xnor U12330 (N_12330,N_11684,N_11761);
or U12331 (N_12331,N_11988,N_11954);
xnor U12332 (N_12332,N_11689,N_11936);
nand U12333 (N_12333,N_11899,N_11869);
nand U12334 (N_12334,N_11849,N_11978);
or U12335 (N_12335,N_11905,N_11855);
nand U12336 (N_12336,N_11881,N_11714);
and U12337 (N_12337,N_11777,N_11888);
nor U12338 (N_12338,N_11666,N_11949);
nand U12339 (N_12339,N_11742,N_11935);
nand U12340 (N_12340,N_11809,N_11815);
nor U12341 (N_12341,N_11624,N_11705);
and U12342 (N_12342,N_11843,N_11789);
nor U12343 (N_12343,N_11621,N_11771);
nor U12344 (N_12344,N_11935,N_11776);
nand U12345 (N_12345,N_11624,N_11911);
nand U12346 (N_12346,N_11915,N_11989);
xnor U12347 (N_12347,N_11933,N_11887);
and U12348 (N_12348,N_11941,N_11757);
or U12349 (N_12349,N_11784,N_11958);
nand U12350 (N_12350,N_11666,N_11718);
nor U12351 (N_12351,N_11721,N_11911);
nand U12352 (N_12352,N_11891,N_11884);
and U12353 (N_12353,N_11721,N_11623);
and U12354 (N_12354,N_11961,N_11904);
nand U12355 (N_12355,N_11915,N_11902);
and U12356 (N_12356,N_11739,N_11952);
nand U12357 (N_12357,N_11929,N_11805);
xor U12358 (N_12358,N_11862,N_11776);
xor U12359 (N_12359,N_11786,N_11760);
nor U12360 (N_12360,N_11764,N_11665);
or U12361 (N_12361,N_11781,N_11670);
nand U12362 (N_12362,N_11991,N_11732);
nor U12363 (N_12363,N_11658,N_11732);
nand U12364 (N_12364,N_11600,N_11788);
nor U12365 (N_12365,N_11759,N_11672);
nand U12366 (N_12366,N_11902,N_11950);
and U12367 (N_12367,N_11982,N_11721);
or U12368 (N_12368,N_11640,N_11643);
nor U12369 (N_12369,N_11657,N_11614);
or U12370 (N_12370,N_11835,N_11803);
or U12371 (N_12371,N_11953,N_11723);
or U12372 (N_12372,N_11961,N_11723);
xor U12373 (N_12373,N_11609,N_11996);
xor U12374 (N_12374,N_11810,N_11794);
or U12375 (N_12375,N_11967,N_11781);
and U12376 (N_12376,N_11711,N_11956);
nand U12377 (N_12377,N_11869,N_11704);
nor U12378 (N_12378,N_11907,N_11791);
nor U12379 (N_12379,N_11994,N_11893);
xor U12380 (N_12380,N_11785,N_11635);
nand U12381 (N_12381,N_11678,N_11729);
nor U12382 (N_12382,N_11990,N_11710);
xor U12383 (N_12383,N_11921,N_11604);
xor U12384 (N_12384,N_11915,N_11859);
and U12385 (N_12385,N_11724,N_11997);
and U12386 (N_12386,N_11661,N_11822);
nor U12387 (N_12387,N_11748,N_11834);
nand U12388 (N_12388,N_11973,N_11916);
or U12389 (N_12389,N_11897,N_11627);
nor U12390 (N_12390,N_11897,N_11736);
nand U12391 (N_12391,N_11911,N_11862);
or U12392 (N_12392,N_11966,N_11768);
nand U12393 (N_12393,N_11821,N_11943);
nor U12394 (N_12394,N_11620,N_11709);
nor U12395 (N_12395,N_11855,N_11836);
nand U12396 (N_12396,N_11781,N_11736);
or U12397 (N_12397,N_11672,N_11741);
or U12398 (N_12398,N_11895,N_11642);
nor U12399 (N_12399,N_11657,N_11611);
and U12400 (N_12400,N_12298,N_12261);
nor U12401 (N_12401,N_12061,N_12060);
xor U12402 (N_12402,N_12195,N_12150);
xor U12403 (N_12403,N_12319,N_12218);
nand U12404 (N_12404,N_12334,N_12239);
or U12405 (N_12405,N_12209,N_12048);
nor U12406 (N_12406,N_12127,N_12305);
or U12407 (N_12407,N_12238,N_12352);
or U12408 (N_12408,N_12354,N_12052);
nand U12409 (N_12409,N_12384,N_12093);
nand U12410 (N_12410,N_12234,N_12389);
and U12411 (N_12411,N_12081,N_12024);
nand U12412 (N_12412,N_12097,N_12376);
nor U12413 (N_12413,N_12147,N_12193);
nor U12414 (N_12414,N_12091,N_12278);
nor U12415 (N_12415,N_12217,N_12031);
xnor U12416 (N_12416,N_12009,N_12332);
and U12417 (N_12417,N_12275,N_12341);
xnor U12418 (N_12418,N_12223,N_12393);
and U12419 (N_12419,N_12314,N_12100);
nor U12420 (N_12420,N_12006,N_12324);
nand U12421 (N_12421,N_12382,N_12379);
nand U12422 (N_12422,N_12329,N_12161);
nand U12423 (N_12423,N_12317,N_12152);
nor U12424 (N_12424,N_12023,N_12321);
nor U12425 (N_12425,N_12371,N_12098);
nand U12426 (N_12426,N_12142,N_12342);
and U12427 (N_12427,N_12364,N_12350);
xnor U12428 (N_12428,N_12349,N_12078);
nand U12429 (N_12429,N_12284,N_12079);
xor U12430 (N_12430,N_12102,N_12216);
and U12431 (N_12431,N_12155,N_12337);
xnor U12432 (N_12432,N_12072,N_12309);
xnor U12433 (N_12433,N_12368,N_12140);
or U12434 (N_12434,N_12211,N_12041);
and U12435 (N_12435,N_12158,N_12181);
and U12436 (N_12436,N_12355,N_12221);
nor U12437 (N_12437,N_12119,N_12044);
nand U12438 (N_12438,N_12124,N_12300);
xor U12439 (N_12439,N_12200,N_12062);
nor U12440 (N_12440,N_12328,N_12088);
or U12441 (N_12441,N_12028,N_12299);
and U12442 (N_12442,N_12173,N_12346);
or U12443 (N_12443,N_12198,N_12069);
or U12444 (N_12444,N_12189,N_12000);
and U12445 (N_12445,N_12067,N_12359);
and U12446 (N_12446,N_12361,N_12144);
nor U12447 (N_12447,N_12037,N_12212);
nor U12448 (N_12448,N_12229,N_12270);
and U12449 (N_12449,N_12340,N_12282);
nor U12450 (N_12450,N_12291,N_12071);
xnor U12451 (N_12451,N_12076,N_12104);
and U12452 (N_12452,N_12237,N_12267);
and U12453 (N_12453,N_12146,N_12174);
nor U12454 (N_12454,N_12316,N_12043);
nand U12455 (N_12455,N_12260,N_12378);
nor U12456 (N_12456,N_12369,N_12117);
nor U12457 (N_12457,N_12153,N_12143);
or U12458 (N_12458,N_12265,N_12356);
or U12459 (N_12459,N_12005,N_12049);
nor U12460 (N_12460,N_12302,N_12018);
or U12461 (N_12461,N_12258,N_12344);
xnor U12462 (N_12462,N_12343,N_12345);
xor U12463 (N_12463,N_12053,N_12283);
or U12464 (N_12464,N_12027,N_12003);
nand U12465 (N_12465,N_12370,N_12141);
or U12466 (N_12466,N_12017,N_12279);
xnor U12467 (N_12467,N_12199,N_12290);
or U12468 (N_12468,N_12089,N_12132);
nand U12469 (N_12469,N_12171,N_12177);
nand U12470 (N_12470,N_12358,N_12225);
nor U12471 (N_12471,N_12073,N_12264);
nand U12472 (N_12472,N_12035,N_12013);
xnor U12473 (N_12473,N_12294,N_12263);
or U12474 (N_12474,N_12387,N_12175);
or U12475 (N_12475,N_12289,N_12271);
or U12476 (N_12476,N_12253,N_12327);
nor U12477 (N_12477,N_12019,N_12220);
and U12478 (N_12478,N_12136,N_12054);
or U12479 (N_12479,N_12026,N_12208);
nand U12480 (N_12480,N_12236,N_12178);
xor U12481 (N_12481,N_12310,N_12231);
xnor U12482 (N_12482,N_12167,N_12245);
or U12483 (N_12483,N_12257,N_12168);
and U12484 (N_12484,N_12285,N_12166);
nor U12485 (N_12485,N_12066,N_12107);
nand U12486 (N_12486,N_12111,N_12213);
and U12487 (N_12487,N_12113,N_12274);
and U12488 (N_12488,N_12096,N_12086);
nor U12489 (N_12489,N_12312,N_12391);
and U12490 (N_12490,N_12162,N_12094);
and U12491 (N_12491,N_12247,N_12396);
and U12492 (N_12492,N_12042,N_12046);
xor U12493 (N_12493,N_12183,N_12307);
nand U12494 (N_12494,N_12311,N_12347);
nand U12495 (N_12495,N_12272,N_12135);
and U12496 (N_12496,N_12130,N_12323);
and U12497 (N_12497,N_12115,N_12008);
or U12498 (N_12498,N_12090,N_12256);
xor U12499 (N_12499,N_12151,N_12373);
xnor U12500 (N_12500,N_12118,N_12172);
and U12501 (N_12501,N_12249,N_12095);
or U12502 (N_12502,N_12165,N_12058);
or U12503 (N_12503,N_12110,N_12395);
nand U12504 (N_12504,N_12149,N_12268);
or U12505 (N_12505,N_12084,N_12050);
and U12506 (N_12506,N_12133,N_12336);
xor U12507 (N_12507,N_12390,N_12080);
or U12508 (N_12508,N_12194,N_12301);
and U12509 (N_12509,N_12292,N_12156);
nor U12510 (N_12510,N_12381,N_12039);
nor U12511 (N_12511,N_12322,N_12318);
xor U12512 (N_12512,N_12367,N_12126);
or U12513 (N_12513,N_12365,N_12248);
and U12514 (N_12514,N_12230,N_12068);
or U12515 (N_12515,N_12002,N_12219);
xnor U12516 (N_12516,N_12123,N_12030);
nand U12517 (N_12517,N_12383,N_12269);
and U12518 (N_12518,N_12012,N_12056);
nor U12519 (N_12519,N_12331,N_12295);
nor U12520 (N_12520,N_12197,N_12187);
xnor U12521 (N_12521,N_12250,N_12004);
xnor U12522 (N_12522,N_12109,N_12137);
xnor U12523 (N_12523,N_12235,N_12335);
nor U12524 (N_12524,N_12015,N_12025);
nor U12525 (N_12525,N_12296,N_12159);
nand U12526 (N_12526,N_12085,N_12348);
or U12527 (N_12527,N_12021,N_12108);
or U12528 (N_12528,N_12074,N_12202);
nor U12529 (N_12529,N_12210,N_12164);
nand U12530 (N_12530,N_12315,N_12372);
nor U12531 (N_12531,N_12059,N_12179);
or U12532 (N_12532,N_12385,N_12330);
or U12533 (N_12533,N_12184,N_12160);
nand U12534 (N_12534,N_12105,N_12032);
or U12535 (N_12535,N_12063,N_12033);
nand U12536 (N_12536,N_12047,N_12134);
nor U12537 (N_12537,N_12016,N_12106);
or U12538 (N_12538,N_12287,N_12351);
xor U12539 (N_12539,N_12304,N_12207);
nand U12540 (N_12540,N_12014,N_12240);
nand U12541 (N_12541,N_12399,N_12320);
nor U12542 (N_12542,N_12145,N_12129);
or U12543 (N_12543,N_12333,N_12262);
nand U12544 (N_12544,N_12259,N_12154);
nor U12545 (N_12545,N_12128,N_12297);
and U12546 (N_12546,N_12280,N_12306);
nor U12547 (N_12547,N_12185,N_12040);
nand U12548 (N_12548,N_12246,N_12170);
xor U12549 (N_12549,N_12254,N_12186);
xnor U12550 (N_12550,N_12169,N_12007);
nor U12551 (N_12551,N_12380,N_12397);
nand U12552 (N_12552,N_12339,N_12255);
and U12553 (N_12553,N_12029,N_12363);
xnor U12554 (N_12554,N_12131,N_12308);
or U12555 (N_12555,N_12022,N_12020);
nor U12556 (N_12556,N_12157,N_12176);
nand U12557 (N_12557,N_12051,N_12120);
nor U12558 (N_12558,N_12075,N_12366);
or U12559 (N_12559,N_12163,N_12139);
or U12560 (N_12560,N_12215,N_12055);
nand U12561 (N_12561,N_12057,N_12099);
and U12562 (N_12562,N_12010,N_12293);
nand U12563 (N_12563,N_12011,N_12392);
xor U12564 (N_12564,N_12377,N_12214);
xor U12565 (N_12565,N_12116,N_12325);
and U12566 (N_12566,N_12148,N_12277);
or U12567 (N_12567,N_12243,N_12241);
nor U12568 (N_12568,N_12034,N_12182);
and U12569 (N_12569,N_12190,N_12273);
nor U12570 (N_12570,N_12070,N_12394);
or U12571 (N_12571,N_12303,N_12001);
nor U12572 (N_12572,N_12252,N_12125);
xnor U12573 (N_12573,N_12038,N_12122);
or U12574 (N_12574,N_12188,N_12233);
nor U12575 (N_12575,N_12092,N_12338);
xor U12576 (N_12576,N_12226,N_12045);
or U12577 (N_12577,N_12196,N_12077);
nor U12578 (N_12578,N_12398,N_12374);
and U12579 (N_12579,N_12064,N_12201);
or U12580 (N_12580,N_12083,N_12375);
nor U12581 (N_12581,N_12101,N_12222);
or U12582 (N_12582,N_12286,N_12244);
nand U12583 (N_12583,N_12180,N_12266);
or U12584 (N_12584,N_12065,N_12326);
and U12585 (N_12585,N_12313,N_12386);
xor U12586 (N_12586,N_12288,N_12205);
and U12587 (N_12587,N_12036,N_12276);
and U12588 (N_12588,N_12138,N_12082);
and U12589 (N_12589,N_12242,N_12360);
nor U12590 (N_12590,N_12191,N_12227);
or U12591 (N_12591,N_12281,N_12087);
nor U12592 (N_12592,N_12192,N_12357);
xor U12593 (N_12593,N_12362,N_12203);
or U12594 (N_12594,N_12112,N_12353);
nand U12595 (N_12595,N_12206,N_12232);
or U12596 (N_12596,N_12228,N_12388);
nor U12597 (N_12597,N_12103,N_12121);
or U12598 (N_12598,N_12204,N_12224);
nand U12599 (N_12599,N_12114,N_12251);
nand U12600 (N_12600,N_12154,N_12086);
nand U12601 (N_12601,N_12244,N_12092);
or U12602 (N_12602,N_12334,N_12066);
or U12603 (N_12603,N_12040,N_12127);
nand U12604 (N_12604,N_12331,N_12191);
xnor U12605 (N_12605,N_12240,N_12090);
or U12606 (N_12606,N_12322,N_12068);
and U12607 (N_12607,N_12136,N_12187);
and U12608 (N_12608,N_12079,N_12264);
xnor U12609 (N_12609,N_12102,N_12387);
xor U12610 (N_12610,N_12215,N_12247);
nand U12611 (N_12611,N_12320,N_12280);
nand U12612 (N_12612,N_12397,N_12138);
nand U12613 (N_12613,N_12027,N_12121);
xor U12614 (N_12614,N_12151,N_12351);
and U12615 (N_12615,N_12113,N_12278);
or U12616 (N_12616,N_12155,N_12015);
nand U12617 (N_12617,N_12020,N_12254);
nand U12618 (N_12618,N_12216,N_12269);
xnor U12619 (N_12619,N_12214,N_12374);
xor U12620 (N_12620,N_12023,N_12282);
xor U12621 (N_12621,N_12307,N_12049);
or U12622 (N_12622,N_12283,N_12302);
nand U12623 (N_12623,N_12344,N_12078);
and U12624 (N_12624,N_12119,N_12207);
nor U12625 (N_12625,N_12341,N_12015);
nand U12626 (N_12626,N_12162,N_12282);
nor U12627 (N_12627,N_12023,N_12228);
and U12628 (N_12628,N_12318,N_12269);
nand U12629 (N_12629,N_12126,N_12101);
nor U12630 (N_12630,N_12373,N_12212);
nand U12631 (N_12631,N_12022,N_12228);
xnor U12632 (N_12632,N_12311,N_12286);
nor U12633 (N_12633,N_12138,N_12324);
or U12634 (N_12634,N_12363,N_12263);
or U12635 (N_12635,N_12092,N_12161);
and U12636 (N_12636,N_12050,N_12365);
and U12637 (N_12637,N_12035,N_12190);
xnor U12638 (N_12638,N_12347,N_12232);
or U12639 (N_12639,N_12203,N_12285);
nand U12640 (N_12640,N_12090,N_12234);
and U12641 (N_12641,N_12212,N_12123);
nor U12642 (N_12642,N_12058,N_12329);
nor U12643 (N_12643,N_12014,N_12148);
and U12644 (N_12644,N_12248,N_12217);
nand U12645 (N_12645,N_12361,N_12097);
and U12646 (N_12646,N_12101,N_12062);
nor U12647 (N_12647,N_12113,N_12164);
xor U12648 (N_12648,N_12242,N_12070);
xor U12649 (N_12649,N_12128,N_12298);
or U12650 (N_12650,N_12186,N_12006);
nor U12651 (N_12651,N_12229,N_12303);
nand U12652 (N_12652,N_12275,N_12362);
nor U12653 (N_12653,N_12199,N_12191);
or U12654 (N_12654,N_12100,N_12069);
nor U12655 (N_12655,N_12130,N_12175);
or U12656 (N_12656,N_12032,N_12269);
nand U12657 (N_12657,N_12014,N_12123);
or U12658 (N_12658,N_12377,N_12018);
nand U12659 (N_12659,N_12368,N_12300);
nand U12660 (N_12660,N_12281,N_12373);
and U12661 (N_12661,N_12216,N_12022);
xnor U12662 (N_12662,N_12377,N_12392);
nor U12663 (N_12663,N_12261,N_12119);
and U12664 (N_12664,N_12017,N_12025);
nor U12665 (N_12665,N_12291,N_12239);
or U12666 (N_12666,N_12122,N_12095);
nor U12667 (N_12667,N_12174,N_12090);
and U12668 (N_12668,N_12191,N_12183);
and U12669 (N_12669,N_12375,N_12354);
and U12670 (N_12670,N_12204,N_12133);
or U12671 (N_12671,N_12277,N_12035);
nor U12672 (N_12672,N_12035,N_12017);
or U12673 (N_12673,N_12107,N_12213);
nand U12674 (N_12674,N_12213,N_12014);
and U12675 (N_12675,N_12322,N_12053);
nor U12676 (N_12676,N_12202,N_12153);
nor U12677 (N_12677,N_12245,N_12013);
nand U12678 (N_12678,N_12012,N_12347);
nand U12679 (N_12679,N_12068,N_12298);
and U12680 (N_12680,N_12371,N_12249);
nand U12681 (N_12681,N_12030,N_12343);
and U12682 (N_12682,N_12107,N_12033);
nand U12683 (N_12683,N_12025,N_12075);
xnor U12684 (N_12684,N_12347,N_12188);
nand U12685 (N_12685,N_12078,N_12038);
and U12686 (N_12686,N_12245,N_12182);
and U12687 (N_12687,N_12147,N_12251);
or U12688 (N_12688,N_12367,N_12068);
nor U12689 (N_12689,N_12125,N_12171);
and U12690 (N_12690,N_12346,N_12115);
xor U12691 (N_12691,N_12386,N_12029);
xnor U12692 (N_12692,N_12280,N_12239);
nor U12693 (N_12693,N_12397,N_12037);
or U12694 (N_12694,N_12189,N_12319);
nand U12695 (N_12695,N_12282,N_12145);
nor U12696 (N_12696,N_12103,N_12057);
and U12697 (N_12697,N_12050,N_12211);
or U12698 (N_12698,N_12385,N_12353);
xor U12699 (N_12699,N_12246,N_12193);
or U12700 (N_12700,N_12004,N_12017);
nand U12701 (N_12701,N_12030,N_12166);
or U12702 (N_12702,N_12357,N_12366);
xnor U12703 (N_12703,N_12147,N_12214);
and U12704 (N_12704,N_12204,N_12339);
and U12705 (N_12705,N_12223,N_12309);
nand U12706 (N_12706,N_12361,N_12304);
nand U12707 (N_12707,N_12004,N_12342);
and U12708 (N_12708,N_12058,N_12098);
xnor U12709 (N_12709,N_12062,N_12213);
xnor U12710 (N_12710,N_12233,N_12111);
xor U12711 (N_12711,N_12046,N_12320);
xnor U12712 (N_12712,N_12017,N_12348);
nand U12713 (N_12713,N_12327,N_12008);
and U12714 (N_12714,N_12041,N_12353);
or U12715 (N_12715,N_12161,N_12306);
and U12716 (N_12716,N_12341,N_12325);
and U12717 (N_12717,N_12120,N_12199);
xor U12718 (N_12718,N_12207,N_12274);
xnor U12719 (N_12719,N_12270,N_12320);
and U12720 (N_12720,N_12363,N_12241);
nor U12721 (N_12721,N_12198,N_12369);
and U12722 (N_12722,N_12227,N_12086);
nor U12723 (N_12723,N_12100,N_12140);
and U12724 (N_12724,N_12140,N_12337);
nand U12725 (N_12725,N_12074,N_12283);
xnor U12726 (N_12726,N_12109,N_12201);
and U12727 (N_12727,N_12375,N_12374);
xor U12728 (N_12728,N_12361,N_12303);
nor U12729 (N_12729,N_12198,N_12145);
nand U12730 (N_12730,N_12113,N_12092);
and U12731 (N_12731,N_12273,N_12047);
nor U12732 (N_12732,N_12215,N_12365);
or U12733 (N_12733,N_12380,N_12060);
or U12734 (N_12734,N_12099,N_12282);
or U12735 (N_12735,N_12135,N_12185);
or U12736 (N_12736,N_12030,N_12046);
xor U12737 (N_12737,N_12309,N_12195);
xnor U12738 (N_12738,N_12201,N_12393);
and U12739 (N_12739,N_12392,N_12326);
and U12740 (N_12740,N_12146,N_12375);
nand U12741 (N_12741,N_12058,N_12247);
or U12742 (N_12742,N_12034,N_12269);
xnor U12743 (N_12743,N_12185,N_12331);
xnor U12744 (N_12744,N_12064,N_12397);
xnor U12745 (N_12745,N_12329,N_12114);
nor U12746 (N_12746,N_12229,N_12390);
or U12747 (N_12747,N_12247,N_12056);
nand U12748 (N_12748,N_12035,N_12133);
or U12749 (N_12749,N_12243,N_12276);
and U12750 (N_12750,N_12157,N_12205);
and U12751 (N_12751,N_12249,N_12384);
or U12752 (N_12752,N_12274,N_12159);
nor U12753 (N_12753,N_12021,N_12381);
or U12754 (N_12754,N_12310,N_12054);
and U12755 (N_12755,N_12213,N_12328);
or U12756 (N_12756,N_12228,N_12062);
nor U12757 (N_12757,N_12044,N_12286);
and U12758 (N_12758,N_12059,N_12132);
or U12759 (N_12759,N_12031,N_12232);
or U12760 (N_12760,N_12204,N_12125);
or U12761 (N_12761,N_12308,N_12003);
xnor U12762 (N_12762,N_12270,N_12070);
nor U12763 (N_12763,N_12111,N_12207);
or U12764 (N_12764,N_12216,N_12015);
or U12765 (N_12765,N_12265,N_12231);
or U12766 (N_12766,N_12304,N_12038);
nor U12767 (N_12767,N_12333,N_12392);
nor U12768 (N_12768,N_12272,N_12233);
nor U12769 (N_12769,N_12127,N_12146);
nor U12770 (N_12770,N_12016,N_12192);
xor U12771 (N_12771,N_12358,N_12084);
and U12772 (N_12772,N_12249,N_12210);
nor U12773 (N_12773,N_12356,N_12396);
nand U12774 (N_12774,N_12178,N_12169);
xnor U12775 (N_12775,N_12272,N_12070);
or U12776 (N_12776,N_12202,N_12098);
or U12777 (N_12777,N_12162,N_12072);
or U12778 (N_12778,N_12238,N_12312);
nor U12779 (N_12779,N_12257,N_12234);
nor U12780 (N_12780,N_12219,N_12054);
xnor U12781 (N_12781,N_12145,N_12030);
nand U12782 (N_12782,N_12378,N_12214);
nor U12783 (N_12783,N_12294,N_12250);
xor U12784 (N_12784,N_12292,N_12296);
or U12785 (N_12785,N_12017,N_12281);
and U12786 (N_12786,N_12149,N_12355);
or U12787 (N_12787,N_12070,N_12153);
nor U12788 (N_12788,N_12259,N_12069);
and U12789 (N_12789,N_12077,N_12387);
or U12790 (N_12790,N_12243,N_12129);
and U12791 (N_12791,N_12186,N_12060);
nor U12792 (N_12792,N_12307,N_12172);
and U12793 (N_12793,N_12057,N_12338);
or U12794 (N_12794,N_12281,N_12001);
and U12795 (N_12795,N_12191,N_12067);
nor U12796 (N_12796,N_12087,N_12193);
and U12797 (N_12797,N_12143,N_12083);
xor U12798 (N_12798,N_12382,N_12272);
nor U12799 (N_12799,N_12045,N_12320);
nand U12800 (N_12800,N_12584,N_12736);
nand U12801 (N_12801,N_12442,N_12580);
nand U12802 (N_12802,N_12737,N_12415);
nand U12803 (N_12803,N_12441,N_12431);
or U12804 (N_12804,N_12590,N_12739);
nor U12805 (N_12805,N_12464,N_12401);
or U12806 (N_12806,N_12466,N_12643);
nor U12807 (N_12807,N_12793,N_12731);
nor U12808 (N_12808,N_12542,N_12747);
or U12809 (N_12809,N_12788,N_12512);
nor U12810 (N_12810,N_12404,N_12735);
nand U12811 (N_12811,N_12725,N_12754);
nor U12812 (N_12812,N_12429,N_12406);
or U12813 (N_12813,N_12541,N_12785);
xnor U12814 (N_12814,N_12412,N_12701);
nor U12815 (N_12815,N_12524,N_12496);
or U12816 (N_12816,N_12543,N_12684);
nor U12817 (N_12817,N_12640,N_12717);
xnor U12818 (N_12818,N_12636,N_12795);
xor U12819 (N_12819,N_12693,N_12723);
xor U12820 (N_12820,N_12528,N_12417);
xnor U12821 (N_12821,N_12764,N_12500);
nor U12822 (N_12822,N_12772,N_12545);
and U12823 (N_12823,N_12537,N_12771);
nand U12824 (N_12824,N_12597,N_12465);
and U12825 (N_12825,N_12573,N_12539);
nor U12826 (N_12826,N_12400,N_12756);
or U12827 (N_12827,N_12435,N_12471);
xor U12828 (N_12828,N_12484,N_12741);
nor U12829 (N_12829,N_12689,N_12522);
or U12830 (N_12830,N_12463,N_12687);
nor U12831 (N_12831,N_12549,N_12581);
nor U12832 (N_12832,N_12599,N_12683);
nand U12833 (N_12833,N_12787,N_12510);
and U12834 (N_12834,N_12458,N_12715);
xor U12835 (N_12835,N_12409,N_12613);
and U12836 (N_12836,N_12630,N_12553);
or U12837 (N_12837,N_12713,N_12662);
and U12838 (N_12838,N_12766,N_12637);
nand U12839 (N_12839,N_12418,N_12420);
xor U12840 (N_12840,N_12469,N_12746);
and U12841 (N_12841,N_12798,N_12668);
nor U12842 (N_12842,N_12428,N_12563);
xor U12843 (N_12843,N_12661,N_12583);
and U12844 (N_12844,N_12680,N_12436);
or U12845 (N_12845,N_12757,N_12538);
nand U12846 (N_12846,N_12489,N_12686);
nand U12847 (N_12847,N_12732,N_12624);
nor U12848 (N_12848,N_12425,N_12718);
xnor U12849 (N_12849,N_12501,N_12726);
xor U12850 (N_12850,N_12768,N_12742);
nor U12851 (N_12851,N_12738,N_12504);
nor U12852 (N_12852,N_12438,N_12492);
nor U12853 (N_12853,N_12454,N_12432);
and U12854 (N_12854,N_12797,N_12440);
nand U12855 (N_12855,N_12632,N_12555);
nor U12856 (N_12856,N_12600,N_12786);
xor U12857 (N_12857,N_12696,N_12799);
and U12858 (N_12858,N_12499,N_12403);
nor U12859 (N_12859,N_12470,N_12473);
nand U12860 (N_12860,N_12783,N_12426);
or U12861 (N_12861,N_12607,N_12618);
nand U12862 (N_12862,N_12678,N_12519);
xnor U12863 (N_12863,N_12535,N_12646);
nand U12864 (N_12864,N_12762,N_12720);
and U12865 (N_12865,N_12494,N_12421);
xor U12866 (N_12866,N_12777,N_12459);
xnor U12867 (N_12867,N_12423,N_12532);
nor U12868 (N_12868,N_12571,N_12413);
xor U12869 (N_12869,N_12617,N_12619);
and U12870 (N_12870,N_12478,N_12633);
nand U12871 (N_12871,N_12449,N_12759);
xor U12872 (N_12872,N_12775,N_12482);
or U12873 (N_12873,N_12779,N_12782);
or U12874 (N_12874,N_12550,N_12536);
nor U12875 (N_12875,N_12649,N_12416);
nand U12876 (N_12876,N_12576,N_12620);
nor U12877 (N_12877,N_12530,N_12758);
xnor U12878 (N_12878,N_12452,N_12751);
and U12879 (N_12879,N_12491,N_12712);
nand U12880 (N_12880,N_12657,N_12424);
or U12881 (N_12881,N_12695,N_12439);
or U12882 (N_12882,N_12707,N_12628);
and U12883 (N_12883,N_12750,N_12774);
xnor U12884 (N_12884,N_12513,N_12767);
and U12885 (N_12885,N_12655,N_12548);
nor U12886 (N_12886,N_12588,N_12658);
and U12887 (N_12887,N_12733,N_12704);
xor U12888 (N_12888,N_12517,N_12722);
and U12889 (N_12889,N_12527,N_12670);
xnor U12890 (N_12890,N_12601,N_12564);
xnor U12891 (N_12891,N_12534,N_12474);
and U12892 (N_12892,N_12461,N_12688);
and U12893 (N_12893,N_12450,N_12457);
nand U12894 (N_12894,N_12690,N_12647);
and U12895 (N_12895,N_12546,N_12748);
or U12896 (N_12896,N_12521,N_12638);
nand U12897 (N_12897,N_12652,N_12559);
or U12898 (N_12898,N_12790,N_12666);
nor U12899 (N_12899,N_12488,N_12744);
or U12900 (N_12900,N_12639,N_12664);
xor U12901 (N_12901,N_12631,N_12634);
xnor U12902 (N_12902,N_12414,N_12547);
or U12903 (N_12903,N_12586,N_12481);
nand U12904 (N_12904,N_12650,N_12453);
or U12905 (N_12905,N_12674,N_12616);
and U12906 (N_12906,N_12653,N_12468);
nand U12907 (N_12907,N_12752,N_12677);
nor U12908 (N_12908,N_12502,N_12503);
or U12909 (N_12909,N_12525,N_12780);
or U12910 (N_12910,N_12515,N_12427);
and U12911 (N_12911,N_12663,N_12497);
or U12912 (N_12912,N_12595,N_12511);
xor U12913 (N_12913,N_12598,N_12681);
and U12914 (N_12914,N_12740,N_12665);
or U12915 (N_12915,N_12669,N_12794);
nor U12916 (N_12916,N_12654,N_12721);
nor U12917 (N_12917,N_12765,N_12611);
nand U12918 (N_12918,N_12572,N_12671);
nand U12919 (N_12919,N_12627,N_12667);
xnor U12920 (N_12920,N_12480,N_12596);
nor U12921 (N_12921,N_12609,N_12694);
nand U12922 (N_12922,N_12495,N_12753);
or U12923 (N_12923,N_12685,N_12743);
nand U12924 (N_12924,N_12791,N_12789);
nor U12925 (N_12925,N_12778,N_12625);
or U12926 (N_12926,N_12760,N_12621);
and U12927 (N_12927,N_12579,N_12734);
or U12928 (N_12928,N_12716,N_12410);
nor U12929 (N_12929,N_12703,N_12591);
nor U12930 (N_12930,N_12659,N_12648);
xor U12931 (N_12931,N_12635,N_12516);
xnor U12932 (N_12932,N_12592,N_12566);
or U12933 (N_12933,N_12518,N_12577);
or U12934 (N_12934,N_12477,N_12444);
xnor U12935 (N_12935,N_12569,N_12498);
xnor U12936 (N_12936,N_12508,N_12606);
nor U12937 (N_12937,N_12608,N_12682);
nand U12938 (N_12938,N_12675,N_12514);
nor U12939 (N_12939,N_12434,N_12673);
or U12940 (N_12940,N_12552,N_12763);
and U12941 (N_12941,N_12520,N_12603);
or U12942 (N_12942,N_12781,N_12448);
nor U12943 (N_12943,N_12587,N_12557);
or U12944 (N_12944,N_12724,N_12589);
nor U12945 (N_12945,N_12565,N_12460);
or U12946 (N_12946,N_12604,N_12651);
nor U12947 (N_12947,N_12411,N_12697);
nand U12948 (N_12948,N_12728,N_12554);
nand U12949 (N_12949,N_12614,N_12551);
nand U12950 (N_12950,N_12472,N_12476);
xnor U12951 (N_12951,N_12594,N_12729);
or U12952 (N_12952,N_12691,N_12506);
nand U12953 (N_12953,N_12433,N_12405);
nor U12954 (N_12954,N_12575,N_12509);
nand U12955 (N_12955,N_12479,N_12582);
nand U12956 (N_12956,N_12578,N_12711);
and U12957 (N_12957,N_12602,N_12702);
and U12958 (N_12958,N_12408,N_12523);
or U12959 (N_12959,N_12419,N_12612);
and U12960 (N_12960,N_12487,N_12483);
nor U12961 (N_12961,N_12706,N_12585);
nand U12962 (N_12962,N_12531,N_12769);
or U12963 (N_12963,N_12610,N_12773);
nand U12964 (N_12964,N_12570,N_12644);
and U12965 (N_12965,N_12709,N_12490);
or U12966 (N_12966,N_12462,N_12719);
nor U12967 (N_12967,N_12792,N_12761);
and U12968 (N_12968,N_12467,N_12402);
and U12969 (N_12969,N_12698,N_12770);
or U12970 (N_12970,N_12708,N_12562);
or U12971 (N_12971,N_12533,N_12642);
and U12972 (N_12972,N_12446,N_12561);
and U12973 (N_12973,N_12456,N_12507);
or U12974 (N_12974,N_12796,N_12676);
and U12975 (N_12975,N_12486,N_12623);
and U12976 (N_12976,N_12730,N_12422);
nor U12977 (N_12977,N_12710,N_12540);
or U12978 (N_12978,N_12645,N_12749);
xor U12979 (N_12979,N_12672,N_12451);
and U12980 (N_12980,N_12656,N_12443);
and U12981 (N_12981,N_12679,N_12556);
xor U12982 (N_12982,N_12475,N_12529);
nand U12983 (N_12983,N_12692,N_12437);
or U12984 (N_12984,N_12447,N_12784);
nand U12985 (N_12985,N_12745,N_12605);
nand U12986 (N_12986,N_12705,N_12544);
or U12987 (N_12987,N_12593,N_12641);
nand U12988 (N_12988,N_12700,N_12615);
nor U12989 (N_12989,N_12714,N_12430);
nor U12990 (N_12990,N_12574,N_12560);
or U12991 (N_12991,N_12568,N_12505);
and U12992 (N_12992,N_12445,N_12493);
and U12993 (N_12993,N_12407,N_12626);
nand U12994 (N_12994,N_12629,N_12622);
xnor U12995 (N_12995,N_12526,N_12776);
and U12996 (N_12996,N_12727,N_12755);
and U12997 (N_12997,N_12455,N_12485);
nand U12998 (N_12998,N_12699,N_12558);
or U12999 (N_12999,N_12660,N_12567);
xor U13000 (N_13000,N_12548,N_12789);
nor U13001 (N_13001,N_12774,N_12475);
nand U13002 (N_13002,N_12536,N_12620);
xnor U13003 (N_13003,N_12569,N_12784);
nor U13004 (N_13004,N_12452,N_12647);
xor U13005 (N_13005,N_12493,N_12739);
and U13006 (N_13006,N_12506,N_12581);
and U13007 (N_13007,N_12457,N_12591);
and U13008 (N_13008,N_12422,N_12577);
or U13009 (N_13009,N_12646,N_12706);
nor U13010 (N_13010,N_12644,N_12442);
nor U13011 (N_13011,N_12498,N_12559);
and U13012 (N_13012,N_12717,N_12447);
or U13013 (N_13013,N_12690,N_12449);
nand U13014 (N_13014,N_12551,N_12589);
or U13015 (N_13015,N_12504,N_12654);
nand U13016 (N_13016,N_12589,N_12609);
and U13017 (N_13017,N_12531,N_12740);
nand U13018 (N_13018,N_12645,N_12405);
xor U13019 (N_13019,N_12756,N_12536);
and U13020 (N_13020,N_12643,N_12690);
nor U13021 (N_13021,N_12625,N_12604);
or U13022 (N_13022,N_12712,N_12713);
xor U13023 (N_13023,N_12748,N_12658);
or U13024 (N_13024,N_12434,N_12540);
xnor U13025 (N_13025,N_12657,N_12730);
and U13026 (N_13026,N_12652,N_12506);
nor U13027 (N_13027,N_12606,N_12542);
or U13028 (N_13028,N_12545,N_12635);
or U13029 (N_13029,N_12564,N_12738);
and U13030 (N_13030,N_12710,N_12743);
nand U13031 (N_13031,N_12404,N_12712);
and U13032 (N_13032,N_12428,N_12790);
or U13033 (N_13033,N_12500,N_12450);
nand U13034 (N_13034,N_12729,N_12493);
and U13035 (N_13035,N_12782,N_12533);
nand U13036 (N_13036,N_12719,N_12508);
nand U13037 (N_13037,N_12633,N_12468);
nor U13038 (N_13038,N_12568,N_12532);
or U13039 (N_13039,N_12433,N_12436);
and U13040 (N_13040,N_12752,N_12569);
or U13041 (N_13041,N_12648,N_12755);
and U13042 (N_13042,N_12788,N_12555);
nand U13043 (N_13043,N_12503,N_12495);
nand U13044 (N_13044,N_12736,N_12627);
or U13045 (N_13045,N_12653,N_12639);
and U13046 (N_13046,N_12579,N_12643);
nor U13047 (N_13047,N_12441,N_12466);
or U13048 (N_13048,N_12502,N_12706);
and U13049 (N_13049,N_12522,N_12435);
xor U13050 (N_13050,N_12422,N_12709);
nor U13051 (N_13051,N_12574,N_12542);
nand U13052 (N_13052,N_12495,N_12492);
or U13053 (N_13053,N_12571,N_12660);
or U13054 (N_13054,N_12527,N_12513);
and U13055 (N_13055,N_12622,N_12542);
or U13056 (N_13056,N_12495,N_12759);
and U13057 (N_13057,N_12506,N_12615);
nand U13058 (N_13058,N_12726,N_12534);
and U13059 (N_13059,N_12456,N_12573);
nand U13060 (N_13060,N_12656,N_12537);
nor U13061 (N_13061,N_12739,N_12531);
and U13062 (N_13062,N_12592,N_12770);
xor U13063 (N_13063,N_12550,N_12480);
nor U13064 (N_13064,N_12779,N_12446);
and U13065 (N_13065,N_12450,N_12416);
xor U13066 (N_13066,N_12500,N_12795);
nor U13067 (N_13067,N_12757,N_12660);
xnor U13068 (N_13068,N_12625,N_12505);
and U13069 (N_13069,N_12681,N_12447);
and U13070 (N_13070,N_12771,N_12716);
nor U13071 (N_13071,N_12651,N_12713);
nor U13072 (N_13072,N_12425,N_12417);
xor U13073 (N_13073,N_12469,N_12456);
and U13074 (N_13074,N_12674,N_12531);
xnor U13075 (N_13075,N_12771,N_12405);
or U13076 (N_13076,N_12441,N_12770);
or U13077 (N_13077,N_12468,N_12794);
nand U13078 (N_13078,N_12734,N_12436);
nor U13079 (N_13079,N_12649,N_12773);
xor U13080 (N_13080,N_12526,N_12600);
nor U13081 (N_13081,N_12421,N_12585);
nand U13082 (N_13082,N_12520,N_12442);
and U13083 (N_13083,N_12404,N_12546);
nand U13084 (N_13084,N_12622,N_12572);
and U13085 (N_13085,N_12591,N_12473);
or U13086 (N_13086,N_12499,N_12605);
and U13087 (N_13087,N_12544,N_12776);
xor U13088 (N_13088,N_12489,N_12691);
or U13089 (N_13089,N_12780,N_12590);
and U13090 (N_13090,N_12454,N_12556);
and U13091 (N_13091,N_12479,N_12708);
nor U13092 (N_13092,N_12556,N_12479);
and U13093 (N_13093,N_12489,N_12639);
nand U13094 (N_13094,N_12512,N_12537);
xnor U13095 (N_13095,N_12597,N_12616);
xor U13096 (N_13096,N_12723,N_12417);
xnor U13097 (N_13097,N_12741,N_12647);
or U13098 (N_13098,N_12508,N_12440);
and U13099 (N_13099,N_12503,N_12460);
and U13100 (N_13100,N_12700,N_12440);
nand U13101 (N_13101,N_12531,N_12470);
and U13102 (N_13102,N_12774,N_12436);
and U13103 (N_13103,N_12479,N_12725);
nor U13104 (N_13104,N_12556,N_12477);
xnor U13105 (N_13105,N_12685,N_12566);
nor U13106 (N_13106,N_12655,N_12626);
and U13107 (N_13107,N_12514,N_12461);
nor U13108 (N_13108,N_12722,N_12533);
xor U13109 (N_13109,N_12683,N_12795);
nor U13110 (N_13110,N_12622,N_12799);
or U13111 (N_13111,N_12524,N_12579);
and U13112 (N_13112,N_12731,N_12671);
or U13113 (N_13113,N_12527,N_12621);
and U13114 (N_13114,N_12630,N_12674);
nor U13115 (N_13115,N_12448,N_12402);
and U13116 (N_13116,N_12593,N_12576);
nor U13117 (N_13117,N_12571,N_12690);
nor U13118 (N_13118,N_12435,N_12739);
nor U13119 (N_13119,N_12688,N_12454);
nor U13120 (N_13120,N_12782,N_12685);
or U13121 (N_13121,N_12673,N_12783);
nor U13122 (N_13122,N_12590,N_12597);
nand U13123 (N_13123,N_12493,N_12764);
or U13124 (N_13124,N_12648,N_12534);
or U13125 (N_13125,N_12524,N_12438);
nor U13126 (N_13126,N_12513,N_12631);
or U13127 (N_13127,N_12415,N_12519);
nand U13128 (N_13128,N_12733,N_12521);
or U13129 (N_13129,N_12658,N_12723);
and U13130 (N_13130,N_12743,N_12799);
and U13131 (N_13131,N_12521,N_12424);
xor U13132 (N_13132,N_12642,N_12446);
nor U13133 (N_13133,N_12679,N_12475);
or U13134 (N_13134,N_12577,N_12783);
nor U13135 (N_13135,N_12788,N_12595);
xnor U13136 (N_13136,N_12580,N_12445);
and U13137 (N_13137,N_12681,N_12726);
nand U13138 (N_13138,N_12654,N_12750);
and U13139 (N_13139,N_12464,N_12422);
and U13140 (N_13140,N_12485,N_12568);
nor U13141 (N_13141,N_12709,N_12659);
nand U13142 (N_13142,N_12593,N_12409);
xnor U13143 (N_13143,N_12735,N_12415);
or U13144 (N_13144,N_12555,N_12423);
nor U13145 (N_13145,N_12513,N_12606);
xor U13146 (N_13146,N_12595,N_12707);
xnor U13147 (N_13147,N_12509,N_12419);
nor U13148 (N_13148,N_12726,N_12715);
xor U13149 (N_13149,N_12457,N_12447);
and U13150 (N_13150,N_12718,N_12524);
xnor U13151 (N_13151,N_12615,N_12473);
nor U13152 (N_13152,N_12756,N_12475);
and U13153 (N_13153,N_12426,N_12734);
or U13154 (N_13154,N_12773,N_12465);
or U13155 (N_13155,N_12691,N_12571);
xnor U13156 (N_13156,N_12760,N_12677);
or U13157 (N_13157,N_12786,N_12790);
nor U13158 (N_13158,N_12411,N_12438);
and U13159 (N_13159,N_12421,N_12580);
nor U13160 (N_13160,N_12763,N_12445);
nor U13161 (N_13161,N_12432,N_12722);
and U13162 (N_13162,N_12662,N_12549);
xnor U13163 (N_13163,N_12693,N_12611);
nand U13164 (N_13164,N_12415,N_12442);
nand U13165 (N_13165,N_12418,N_12564);
nor U13166 (N_13166,N_12611,N_12753);
nor U13167 (N_13167,N_12630,N_12742);
and U13168 (N_13168,N_12431,N_12520);
xor U13169 (N_13169,N_12429,N_12602);
and U13170 (N_13170,N_12488,N_12740);
nand U13171 (N_13171,N_12511,N_12723);
nand U13172 (N_13172,N_12428,N_12636);
nor U13173 (N_13173,N_12599,N_12616);
nor U13174 (N_13174,N_12522,N_12624);
and U13175 (N_13175,N_12400,N_12524);
nor U13176 (N_13176,N_12597,N_12516);
and U13177 (N_13177,N_12640,N_12449);
nand U13178 (N_13178,N_12795,N_12709);
and U13179 (N_13179,N_12614,N_12789);
nor U13180 (N_13180,N_12756,N_12635);
nand U13181 (N_13181,N_12743,N_12764);
and U13182 (N_13182,N_12682,N_12502);
xor U13183 (N_13183,N_12644,N_12684);
or U13184 (N_13184,N_12632,N_12606);
or U13185 (N_13185,N_12612,N_12778);
xor U13186 (N_13186,N_12718,N_12616);
xor U13187 (N_13187,N_12770,N_12520);
xnor U13188 (N_13188,N_12491,N_12745);
nand U13189 (N_13189,N_12696,N_12428);
or U13190 (N_13190,N_12445,N_12716);
xnor U13191 (N_13191,N_12503,N_12765);
xor U13192 (N_13192,N_12480,N_12458);
or U13193 (N_13193,N_12505,N_12523);
and U13194 (N_13194,N_12549,N_12604);
xor U13195 (N_13195,N_12791,N_12579);
xor U13196 (N_13196,N_12746,N_12634);
xor U13197 (N_13197,N_12587,N_12648);
nor U13198 (N_13198,N_12747,N_12794);
or U13199 (N_13199,N_12504,N_12413);
and U13200 (N_13200,N_13090,N_12992);
or U13201 (N_13201,N_13183,N_12845);
nor U13202 (N_13202,N_13058,N_13133);
xor U13203 (N_13203,N_13032,N_12838);
nor U13204 (N_13204,N_12927,N_13083);
or U13205 (N_13205,N_13068,N_13085);
or U13206 (N_13206,N_13117,N_12981);
nor U13207 (N_13207,N_13026,N_12949);
xor U13208 (N_13208,N_12819,N_12939);
or U13209 (N_13209,N_13097,N_12916);
nand U13210 (N_13210,N_13066,N_13126);
or U13211 (N_13211,N_13108,N_12945);
or U13212 (N_13212,N_13021,N_13060);
and U13213 (N_13213,N_12964,N_12911);
and U13214 (N_13214,N_12856,N_13182);
nand U13215 (N_13215,N_13132,N_12872);
nor U13216 (N_13216,N_13093,N_12835);
xnor U13217 (N_13217,N_12925,N_13120);
nand U13218 (N_13218,N_12898,N_12812);
and U13219 (N_13219,N_13158,N_12947);
and U13220 (N_13220,N_13003,N_13189);
nor U13221 (N_13221,N_12999,N_13038);
nand U13222 (N_13222,N_13107,N_12941);
xnor U13223 (N_13223,N_13101,N_13043);
and U13224 (N_13224,N_13130,N_13171);
or U13225 (N_13225,N_12952,N_12905);
nand U13226 (N_13226,N_13052,N_12912);
or U13227 (N_13227,N_12948,N_13063);
nor U13228 (N_13228,N_13013,N_13141);
and U13229 (N_13229,N_12896,N_13127);
nand U13230 (N_13230,N_13009,N_12890);
and U13231 (N_13231,N_12994,N_12814);
nand U13232 (N_13232,N_12832,N_12903);
nand U13233 (N_13233,N_12920,N_13007);
and U13234 (N_13234,N_12804,N_13184);
nor U13235 (N_13235,N_12961,N_13165);
or U13236 (N_13236,N_12970,N_12884);
or U13237 (N_13237,N_13096,N_13075);
nand U13238 (N_13238,N_12873,N_12885);
xnor U13239 (N_13239,N_13022,N_13062);
xnor U13240 (N_13240,N_12954,N_12892);
xnor U13241 (N_13241,N_12850,N_12882);
nand U13242 (N_13242,N_12955,N_13014);
or U13243 (N_13243,N_12816,N_13069);
or U13244 (N_13244,N_12888,N_12990);
and U13245 (N_13245,N_13175,N_12843);
or U13246 (N_13246,N_13124,N_12834);
nand U13247 (N_13247,N_12876,N_12844);
or U13248 (N_13248,N_13188,N_12889);
or U13249 (N_13249,N_12871,N_12914);
xnor U13250 (N_13250,N_12931,N_12946);
nand U13251 (N_13251,N_12960,N_12865);
nand U13252 (N_13252,N_12891,N_12822);
xor U13253 (N_13253,N_12842,N_13149);
or U13254 (N_13254,N_12906,N_12817);
and U13255 (N_13255,N_13027,N_13011);
nand U13256 (N_13256,N_13179,N_13154);
xnor U13257 (N_13257,N_13121,N_12953);
or U13258 (N_13258,N_13125,N_12900);
nor U13259 (N_13259,N_13150,N_12858);
nor U13260 (N_13260,N_13010,N_13109);
nor U13261 (N_13261,N_13181,N_12979);
and U13262 (N_13262,N_12963,N_13164);
or U13263 (N_13263,N_13018,N_13049);
nand U13264 (N_13264,N_13185,N_12830);
and U13265 (N_13265,N_12921,N_13077);
nor U13266 (N_13266,N_13145,N_12918);
nor U13267 (N_13267,N_12893,N_13102);
or U13268 (N_13268,N_13174,N_12870);
and U13269 (N_13269,N_13015,N_12840);
nor U13270 (N_13270,N_13129,N_13197);
nor U13271 (N_13271,N_12956,N_13196);
nand U13272 (N_13272,N_13106,N_13084);
or U13273 (N_13273,N_12922,N_12823);
and U13274 (N_13274,N_13000,N_13167);
or U13275 (N_13275,N_13023,N_13156);
nand U13276 (N_13276,N_13155,N_13157);
or U13277 (N_13277,N_12980,N_13016);
or U13278 (N_13278,N_12971,N_13180);
nand U13279 (N_13279,N_13142,N_12839);
xor U13280 (N_13280,N_12818,N_12908);
or U13281 (N_13281,N_13112,N_12877);
nand U13282 (N_13282,N_13136,N_13152);
xnor U13283 (N_13283,N_12988,N_13073);
and U13284 (N_13284,N_13033,N_12808);
or U13285 (N_13285,N_12909,N_12983);
nor U13286 (N_13286,N_13050,N_13059);
xnor U13287 (N_13287,N_13061,N_12824);
xor U13288 (N_13288,N_13161,N_13193);
nor U13289 (N_13289,N_13105,N_12861);
nand U13290 (N_13290,N_12875,N_12864);
and U13291 (N_13291,N_12984,N_13047);
xnor U13292 (N_13292,N_12851,N_12962);
xnor U13293 (N_13293,N_13095,N_12811);
xnor U13294 (N_13294,N_12902,N_12950);
and U13295 (N_13295,N_13192,N_12825);
nor U13296 (N_13296,N_13186,N_12951);
xor U13297 (N_13297,N_13148,N_12860);
nand U13298 (N_13298,N_12829,N_12894);
nor U13299 (N_13299,N_13048,N_13162);
or U13300 (N_13300,N_13113,N_13100);
and U13301 (N_13301,N_13036,N_12959);
and U13302 (N_13302,N_13025,N_13131);
nand U13303 (N_13303,N_12929,N_13122);
nor U13304 (N_13304,N_13064,N_13017);
or U13305 (N_13305,N_12915,N_13054);
and U13306 (N_13306,N_13081,N_12998);
xor U13307 (N_13307,N_12923,N_13044);
nor U13308 (N_13308,N_12813,N_12879);
nand U13309 (N_13309,N_12837,N_12828);
and U13310 (N_13310,N_13045,N_13187);
nor U13311 (N_13311,N_12801,N_12869);
xnor U13312 (N_13312,N_13039,N_13191);
xor U13313 (N_13313,N_13147,N_12978);
and U13314 (N_13314,N_13087,N_12836);
nor U13315 (N_13315,N_12933,N_12853);
nor U13316 (N_13316,N_12926,N_12886);
nand U13317 (N_13317,N_12967,N_13176);
xor U13318 (N_13318,N_13067,N_13159);
xor U13319 (N_13319,N_12874,N_13041);
nand U13320 (N_13320,N_13094,N_13128);
xor U13321 (N_13321,N_12975,N_13051);
and U13322 (N_13322,N_12965,N_12857);
nor U13323 (N_13323,N_13042,N_13029);
nor U13324 (N_13324,N_13040,N_13134);
xor U13325 (N_13325,N_13005,N_13056);
nand U13326 (N_13326,N_12901,N_12810);
and U13327 (N_13327,N_12815,N_13166);
nand U13328 (N_13328,N_12938,N_12820);
or U13329 (N_13329,N_12934,N_13012);
or U13330 (N_13330,N_13194,N_13089);
nor U13331 (N_13331,N_13076,N_12803);
nand U13332 (N_13332,N_13140,N_12826);
and U13333 (N_13333,N_13198,N_13070);
xnor U13334 (N_13334,N_12936,N_12800);
xnor U13335 (N_13335,N_12805,N_13037);
and U13336 (N_13336,N_13195,N_12942);
nor U13337 (N_13337,N_12995,N_13035);
and U13338 (N_13338,N_12932,N_12868);
xor U13339 (N_13339,N_12881,N_12957);
and U13340 (N_13340,N_13086,N_13151);
nor U13341 (N_13341,N_12993,N_13178);
or U13342 (N_13342,N_12969,N_12996);
nor U13343 (N_13343,N_12924,N_12928);
xor U13344 (N_13344,N_12880,N_12982);
xor U13345 (N_13345,N_13079,N_13053);
nor U13346 (N_13346,N_12987,N_12919);
or U13347 (N_13347,N_12913,N_13071);
xor U13348 (N_13348,N_12966,N_13034);
xnor U13349 (N_13349,N_13004,N_13190);
nand U13350 (N_13350,N_12827,N_12854);
xnor U13351 (N_13351,N_12943,N_12862);
xor U13352 (N_13352,N_13092,N_12833);
nor U13353 (N_13353,N_13104,N_13098);
nor U13354 (N_13354,N_13118,N_12989);
and U13355 (N_13355,N_13031,N_12930);
xnor U13356 (N_13356,N_13138,N_13088);
and U13357 (N_13357,N_13143,N_13024);
and U13358 (N_13358,N_12852,N_12849);
nand U13359 (N_13359,N_12866,N_13006);
or U13360 (N_13360,N_12991,N_13153);
xor U13361 (N_13361,N_12806,N_13074);
or U13362 (N_13362,N_13163,N_13080);
and U13363 (N_13363,N_13110,N_12940);
xnor U13364 (N_13364,N_12883,N_12841);
nand U13365 (N_13365,N_13082,N_12973);
nand U13366 (N_13366,N_13078,N_12904);
nand U13367 (N_13367,N_12972,N_13008);
nand U13368 (N_13368,N_12907,N_12986);
nor U13369 (N_13369,N_13114,N_13119);
nor U13370 (N_13370,N_13160,N_12867);
nand U13371 (N_13371,N_12944,N_12807);
nand U13372 (N_13372,N_12887,N_13137);
nor U13373 (N_13373,N_13135,N_13099);
and U13374 (N_13374,N_13057,N_13177);
and U13375 (N_13375,N_13144,N_13199);
or U13376 (N_13376,N_13055,N_13123);
xnor U13377 (N_13377,N_13030,N_12917);
xnor U13378 (N_13378,N_13001,N_13019);
xor U13379 (N_13379,N_12997,N_12878);
xnor U13380 (N_13380,N_12910,N_13002);
or U13381 (N_13381,N_12977,N_13170);
and U13382 (N_13382,N_13111,N_13065);
and U13383 (N_13383,N_12847,N_12831);
or U13384 (N_13384,N_13091,N_12899);
xor U13385 (N_13385,N_12968,N_13173);
nand U13386 (N_13386,N_12935,N_12976);
nand U13387 (N_13387,N_13103,N_12848);
xor U13388 (N_13388,N_12958,N_13169);
xor U13389 (N_13389,N_12863,N_13172);
nand U13390 (N_13390,N_13146,N_12897);
xor U13391 (N_13391,N_12895,N_13020);
xnor U13392 (N_13392,N_12974,N_13072);
nand U13393 (N_13393,N_12855,N_13046);
or U13394 (N_13394,N_12859,N_13168);
xor U13395 (N_13395,N_13115,N_12821);
xnor U13396 (N_13396,N_13028,N_13116);
or U13397 (N_13397,N_12846,N_12985);
nor U13398 (N_13398,N_12937,N_12809);
nor U13399 (N_13399,N_12802,N_13139);
nand U13400 (N_13400,N_13167,N_12935);
nor U13401 (N_13401,N_12945,N_12821);
xor U13402 (N_13402,N_13173,N_13031);
or U13403 (N_13403,N_12859,N_13094);
or U13404 (N_13404,N_12862,N_13124);
and U13405 (N_13405,N_12990,N_13100);
nor U13406 (N_13406,N_12874,N_12905);
nor U13407 (N_13407,N_13130,N_13005);
nor U13408 (N_13408,N_12889,N_12804);
nand U13409 (N_13409,N_12871,N_13136);
and U13410 (N_13410,N_13137,N_13106);
nor U13411 (N_13411,N_13161,N_12971);
and U13412 (N_13412,N_13074,N_13113);
nand U13413 (N_13413,N_13023,N_12866);
or U13414 (N_13414,N_13010,N_12833);
and U13415 (N_13415,N_13108,N_12827);
and U13416 (N_13416,N_13107,N_13024);
or U13417 (N_13417,N_13155,N_12968);
nor U13418 (N_13418,N_12923,N_12828);
and U13419 (N_13419,N_12961,N_12868);
nor U13420 (N_13420,N_13067,N_12947);
or U13421 (N_13421,N_12945,N_12971);
nand U13422 (N_13422,N_12932,N_12849);
nor U13423 (N_13423,N_13043,N_12901);
nand U13424 (N_13424,N_12975,N_13020);
nand U13425 (N_13425,N_13191,N_13117);
and U13426 (N_13426,N_13162,N_12869);
nand U13427 (N_13427,N_13047,N_12886);
nor U13428 (N_13428,N_13037,N_12974);
or U13429 (N_13429,N_13012,N_13122);
nand U13430 (N_13430,N_12865,N_12942);
and U13431 (N_13431,N_12897,N_12909);
and U13432 (N_13432,N_13179,N_12863);
nand U13433 (N_13433,N_12956,N_13131);
or U13434 (N_13434,N_13132,N_12908);
nor U13435 (N_13435,N_13161,N_12876);
nor U13436 (N_13436,N_12934,N_13074);
or U13437 (N_13437,N_12843,N_12972);
and U13438 (N_13438,N_12801,N_12910);
or U13439 (N_13439,N_13157,N_13124);
or U13440 (N_13440,N_12825,N_12835);
nor U13441 (N_13441,N_12991,N_13089);
and U13442 (N_13442,N_13037,N_12967);
nand U13443 (N_13443,N_13149,N_12958);
nand U13444 (N_13444,N_12905,N_12950);
nand U13445 (N_13445,N_12982,N_13060);
nor U13446 (N_13446,N_13029,N_13151);
nor U13447 (N_13447,N_12997,N_12981);
nand U13448 (N_13448,N_12930,N_12843);
xnor U13449 (N_13449,N_13143,N_12835);
or U13450 (N_13450,N_12831,N_13046);
or U13451 (N_13451,N_12947,N_13016);
nand U13452 (N_13452,N_12800,N_13187);
or U13453 (N_13453,N_13080,N_12917);
and U13454 (N_13454,N_12847,N_12917);
xor U13455 (N_13455,N_12833,N_13186);
nand U13456 (N_13456,N_13166,N_13070);
nand U13457 (N_13457,N_13094,N_13005);
and U13458 (N_13458,N_13191,N_13170);
and U13459 (N_13459,N_13081,N_12826);
xnor U13460 (N_13460,N_12927,N_13093);
nor U13461 (N_13461,N_13126,N_13039);
xnor U13462 (N_13462,N_13036,N_12805);
nor U13463 (N_13463,N_13171,N_12988);
and U13464 (N_13464,N_13176,N_13069);
nor U13465 (N_13465,N_12895,N_12872);
nor U13466 (N_13466,N_12851,N_12891);
and U13467 (N_13467,N_13068,N_12959);
nor U13468 (N_13468,N_13015,N_12946);
xor U13469 (N_13469,N_13126,N_12983);
nand U13470 (N_13470,N_12939,N_13198);
and U13471 (N_13471,N_13042,N_12954);
and U13472 (N_13472,N_13037,N_12802);
nor U13473 (N_13473,N_13087,N_13101);
nand U13474 (N_13474,N_13015,N_12882);
nand U13475 (N_13475,N_12827,N_12934);
and U13476 (N_13476,N_13189,N_12999);
nand U13477 (N_13477,N_13199,N_13121);
nor U13478 (N_13478,N_12911,N_12810);
xor U13479 (N_13479,N_13029,N_13123);
or U13480 (N_13480,N_12826,N_13051);
xor U13481 (N_13481,N_13058,N_13189);
nand U13482 (N_13482,N_12893,N_12804);
and U13483 (N_13483,N_12814,N_13164);
nand U13484 (N_13484,N_13011,N_13008);
nor U13485 (N_13485,N_12945,N_13064);
and U13486 (N_13486,N_13045,N_12876);
nor U13487 (N_13487,N_13079,N_13181);
and U13488 (N_13488,N_12924,N_12825);
nor U13489 (N_13489,N_12853,N_13099);
xnor U13490 (N_13490,N_12926,N_13141);
xor U13491 (N_13491,N_12906,N_13097);
nand U13492 (N_13492,N_12908,N_12932);
nand U13493 (N_13493,N_13060,N_12900);
xnor U13494 (N_13494,N_12822,N_13065);
nand U13495 (N_13495,N_12812,N_12938);
nor U13496 (N_13496,N_13058,N_13103);
nand U13497 (N_13497,N_12887,N_13065);
nor U13498 (N_13498,N_12926,N_12897);
nor U13499 (N_13499,N_13010,N_13182);
or U13500 (N_13500,N_12830,N_12938);
nor U13501 (N_13501,N_12899,N_12877);
and U13502 (N_13502,N_12819,N_13080);
xnor U13503 (N_13503,N_12938,N_13190);
or U13504 (N_13504,N_12826,N_13139);
nand U13505 (N_13505,N_13006,N_13010);
xnor U13506 (N_13506,N_12974,N_13074);
nor U13507 (N_13507,N_12977,N_13016);
or U13508 (N_13508,N_12912,N_12845);
nand U13509 (N_13509,N_12948,N_12938);
nand U13510 (N_13510,N_13171,N_13102);
nand U13511 (N_13511,N_12812,N_12996);
nand U13512 (N_13512,N_12869,N_13020);
or U13513 (N_13513,N_12886,N_13103);
nand U13514 (N_13514,N_12986,N_13188);
or U13515 (N_13515,N_12968,N_12885);
xor U13516 (N_13516,N_13172,N_12951);
xor U13517 (N_13517,N_13195,N_13036);
xnor U13518 (N_13518,N_13148,N_12800);
and U13519 (N_13519,N_12802,N_13130);
nor U13520 (N_13520,N_13122,N_12816);
or U13521 (N_13521,N_12820,N_13199);
and U13522 (N_13522,N_13070,N_13000);
nand U13523 (N_13523,N_13164,N_13098);
xnor U13524 (N_13524,N_13071,N_12834);
and U13525 (N_13525,N_12881,N_13076);
xor U13526 (N_13526,N_13064,N_13016);
nand U13527 (N_13527,N_13184,N_13185);
nand U13528 (N_13528,N_12908,N_13005);
nand U13529 (N_13529,N_13099,N_12946);
nor U13530 (N_13530,N_12893,N_13038);
nor U13531 (N_13531,N_13032,N_12942);
or U13532 (N_13532,N_13053,N_12824);
and U13533 (N_13533,N_12902,N_12995);
nand U13534 (N_13534,N_12978,N_13038);
nor U13535 (N_13535,N_13006,N_13144);
nor U13536 (N_13536,N_12853,N_12810);
nor U13537 (N_13537,N_12960,N_13016);
nor U13538 (N_13538,N_12967,N_12971);
nor U13539 (N_13539,N_12828,N_12882);
nand U13540 (N_13540,N_13066,N_13053);
nand U13541 (N_13541,N_13114,N_13130);
and U13542 (N_13542,N_13118,N_13072);
and U13543 (N_13543,N_13118,N_12863);
or U13544 (N_13544,N_13040,N_13017);
and U13545 (N_13545,N_12878,N_12950);
nand U13546 (N_13546,N_13019,N_12962);
or U13547 (N_13547,N_13084,N_13141);
nor U13548 (N_13548,N_12890,N_12801);
nand U13549 (N_13549,N_12804,N_13000);
and U13550 (N_13550,N_12907,N_12824);
xnor U13551 (N_13551,N_13169,N_12863);
and U13552 (N_13552,N_12809,N_13163);
nor U13553 (N_13553,N_12915,N_13137);
and U13554 (N_13554,N_13069,N_12840);
nand U13555 (N_13555,N_13096,N_13118);
xnor U13556 (N_13556,N_12958,N_13166);
and U13557 (N_13557,N_12901,N_12916);
nand U13558 (N_13558,N_13000,N_13061);
and U13559 (N_13559,N_12985,N_13130);
or U13560 (N_13560,N_13031,N_13097);
and U13561 (N_13561,N_12875,N_13017);
xnor U13562 (N_13562,N_13046,N_12994);
and U13563 (N_13563,N_13115,N_13101);
nand U13564 (N_13564,N_13137,N_12817);
nor U13565 (N_13565,N_12902,N_13056);
nor U13566 (N_13566,N_13016,N_13080);
or U13567 (N_13567,N_12967,N_13029);
and U13568 (N_13568,N_13194,N_12975);
nand U13569 (N_13569,N_12823,N_12808);
or U13570 (N_13570,N_12848,N_13188);
nor U13571 (N_13571,N_13098,N_12837);
nor U13572 (N_13572,N_12801,N_13009);
and U13573 (N_13573,N_13055,N_12885);
and U13574 (N_13574,N_12855,N_13165);
nor U13575 (N_13575,N_12836,N_12893);
nor U13576 (N_13576,N_13182,N_13135);
nand U13577 (N_13577,N_13154,N_12816);
nor U13578 (N_13578,N_13102,N_13168);
and U13579 (N_13579,N_12969,N_13129);
or U13580 (N_13580,N_12969,N_12829);
and U13581 (N_13581,N_13091,N_12916);
nor U13582 (N_13582,N_12888,N_13141);
nand U13583 (N_13583,N_12861,N_12954);
xor U13584 (N_13584,N_13087,N_12916);
or U13585 (N_13585,N_12822,N_13070);
or U13586 (N_13586,N_12850,N_12910);
or U13587 (N_13587,N_13098,N_13038);
or U13588 (N_13588,N_13055,N_12865);
nor U13589 (N_13589,N_12907,N_12897);
nand U13590 (N_13590,N_12949,N_13139);
nand U13591 (N_13591,N_12942,N_13010);
or U13592 (N_13592,N_13193,N_13074);
and U13593 (N_13593,N_12861,N_13162);
or U13594 (N_13594,N_13156,N_13185);
or U13595 (N_13595,N_13056,N_13142);
nor U13596 (N_13596,N_12963,N_12961);
xnor U13597 (N_13597,N_12887,N_12941);
nor U13598 (N_13598,N_12936,N_12850);
and U13599 (N_13599,N_12810,N_12959);
xnor U13600 (N_13600,N_13318,N_13564);
nand U13601 (N_13601,N_13543,N_13528);
nor U13602 (N_13602,N_13407,N_13297);
xor U13603 (N_13603,N_13413,N_13282);
nor U13604 (N_13604,N_13250,N_13520);
or U13605 (N_13605,N_13497,N_13551);
nand U13606 (N_13606,N_13510,N_13245);
nor U13607 (N_13607,N_13498,N_13306);
nand U13608 (N_13608,N_13236,N_13458);
xnor U13609 (N_13609,N_13415,N_13276);
nor U13610 (N_13610,N_13238,N_13588);
and U13611 (N_13611,N_13372,N_13295);
nand U13612 (N_13612,N_13358,N_13486);
xnor U13613 (N_13613,N_13204,N_13547);
nor U13614 (N_13614,N_13262,N_13400);
nand U13615 (N_13615,N_13232,N_13465);
or U13616 (N_13616,N_13502,N_13369);
nand U13617 (N_13617,N_13554,N_13428);
nand U13618 (N_13618,N_13353,N_13409);
or U13619 (N_13619,N_13557,N_13251);
xor U13620 (N_13620,N_13442,N_13203);
or U13621 (N_13621,N_13359,N_13539);
or U13622 (N_13622,N_13269,N_13258);
xnor U13623 (N_13623,N_13509,N_13341);
and U13624 (N_13624,N_13380,N_13491);
nand U13625 (N_13625,N_13538,N_13200);
nand U13626 (N_13626,N_13562,N_13367);
xnor U13627 (N_13627,N_13578,N_13416);
nor U13628 (N_13628,N_13566,N_13345);
or U13629 (N_13629,N_13508,N_13474);
nand U13630 (N_13630,N_13317,N_13363);
nor U13631 (N_13631,N_13266,N_13417);
xor U13632 (N_13632,N_13541,N_13558);
xnor U13633 (N_13633,N_13356,N_13255);
xnor U13634 (N_13634,N_13519,N_13506);
and U13635 (N_13635,N_13252,N_13215);
xnor U13636 (N_13636,N_13343,N_13433);
nor U13637 (N_13637,N_13309,N_13296);
nand U13638 (N_13638,N_13496,N_13438);
or U13639 (N_13639,N_13223,N_13585);
nor U13640 (N_13640,N_13454,N_13597);
nand U13641 (N_13641,N_13555,N_13436);
and U13642 (N_13642,N_13529,N_13336);
nand U13643 (N_13643,N_13459,N_13233);
xor U13644 (N_13644,N_13536,N_13228);
nor U13645 (N_13645,N_13259,N_13319);
nor U13646 (N_13646,N_13587,N_13207);
and U13647 (N_13647,N_13404,N_13337);
xor U13648 (N_13648,N_13396,N_13480);
or U13649 (N_13649,N_13390,N_13584);
and U13650 (N_13650,N_13248,N_13225);
or U13651 (N_13651,N_13446,N_13479);
xnor U13652 (N_13652,N_13441,N_13288);
nor U13653 (N_13653,N_13516,N_13494);
xnor U13654 (N_13654,N_13267,N_13290);
or U13655 (N_13655,N_13527,N_13472);
nor U13656 (N_13656,N_13371,N_13575);
and U13657 (N_13657,N_13549,N_13294);
xor U13658 (N_13658,N_13249,N_13265);
nand U13659 (N_13659,N_13402,N_13305);
nand U13660 (N_13660,N_13565,N_13270);
nor U13661 (N_13661,N_13213,N_13292);
or U13662 (N_13662,N_13456,N_13526);
nor U13663 (N_13663,N_13423,N_13299);
nor U13664 (N_13664,N_13385,N_13210);
nor U13665 (N_13665,N_13420,N_13389);
nor U13666 (N_13666,N_13214,N_13579);
and U13667 (N_13667,N_13589,N_13511);
or U13668 (N_13668,N_13518,N_13339);
or U13669 (N_13669,N_13287,N_13570);
nand U13670 (N_13670,N_13473,N_13544);
xor U13671 (N_13671,N_13531,N_13352);
xnor U13672 (N_13672,N_13350,N_13525);
xor U13673 (N_13673,N_13521,N_13361);
nor U13674 (N_13674,N_13328,N_13462);
nand U13675 (N_13675,N_13332,N_13524);
xnor U13676 (N_13676,N_13362,N_13260);
nand U13677 (N_13677,N_13576,N_13243);
nor U13678 (N_13678,N_13310,N_13383);
nor U13679 (N_13679,N_13439,N_13448);
xor U13680 (N_13680,N_13533,N_13279);
xnor U13681 (N_13681,N_13571,N_13398);
or U13682 (N_13682,N_13340,N_13284);
nor U13683 (N_13683,N_13393,N_13331);
or U13684 (N_13684,N_13573,N_13475);
nor U13685 (N_13685,N_13443,N_13552);
xnor U13686 (N_13686,N_13550,N_13447);
xnor U13687 (N_13687,N_13476,N_13487);
and U13688 (N_13688,N_13230,N_13360);
or U13689 (N_13689,N_13298,N_13212);
or U13690 (N_13690,N_13435,N_13410);
nand U13691 (N_13691,N_13217,N_13501);
or U13692 (N_13692,N_13308,N_13582);
nand U13693 (N_13693,N_13512,N_13285);
xor U13694 (N_13694,N_13515,N_13344);
or U13695 (N_13695,N_13419,N_13395);
nand U13696 (N_13696,N_13507,N_13467);
nor U13697 (N_13697,N_13586,N_13523);
and U13698 (N_13698,N_13239,N_13471);
and U13699 (N_13699,N_13355,N_13444);
xnor U13700 (N_13700,N_13221,N_13424);
nor U13701 (N_13701,N_13503,N_13261);
or U13702 (N_13702,N_13572,N_13440);
xor U13703 (N_13703,N_13202,N_13278);
xnor U13704 (N_13704,N_13324,N_13425);
or U13705 (N_13705,N_13422,N_13253);
nor U13706 (N_13706,N_13263,N_13411);
or U13707 (N_13707,N_13354,N_13379);
and U13708 (N_13708,N_13452,N_13593);
and U13709 (N_13709,N_13325,N_13437);
nor U13710 (N_13710,N_13408,N_13241);
nor U13711 (N_13711,N_13302,N_13590);
nor U13712 (N_13712,N_13545,N_13591);
and U13713 (N_13713,N_13569,N_13322);
nand U13714 (N_13714,N_13553,N_13495);
xnor U13715 (N_13715,N_13374,N_13463);
nor U13716 (N_13716,N_13488,N_13451);
nand U13717 (N_13717,N_13493,N_13429);
xor U13718 (N_13718,N_13468,N_13268);
nand U13719 (N_13719,N_13313,N_13351);
or U13720 (N_13720,N_13530,N_13574);
and U13721 (N_13721,N_13517,N_13235);
xnor U13722 (N_13722,N_13505,N_13485);
nor U13723 (N_13723,N_13542,N_13386);
nand U13724 (N_13724,N_13300,N_13492);
nor U13725 (N_13725,N_13535,N_13321);
or U13726 (N_13726,N_13218,N_13373);
nand U13727 (N_13727,N_13391,N_13381);
or U13728 (N_13728,N_13330,N_13427);
nand U13729 (N_13729,N_13231,N_13466);
xor U13730 (N_13730,N_13375,N_13477);
nor U13731 (N_13731,N_13399,N_13397);
xor U13732 (N_13732,N_13548,N_13418);
or U13733 (N_13733,N_13453,N_13388);
xor U13734 (N_13734,N_13430,N_13303);
nor U13735 (N_13735,N_13532,N_13208);
and U13736 (N_13736,N_13567,N_13273);
and U13737 (N_13737,N_13342,N_13434);
and U13738 (N_13738,N_13594,N_13432);
nor U13739 (N_13739,N_13333,N_13568);
or U13740 (N_13740,N_13504,N_13561);
xnor U13741 (N_13741,N_13312,N_13365);
nand U13742 (N_13742,N_13311,N_13271);
or U13743 (N_13743,N_13334,N_13481);
nand U13744 (N_13744,N_13599,N_13368);
and U13745 (N_13745,N_13357,N_13556);
and U13746 (N_13746,N_13499,N_13450);
or U13747 (N_13747,N_13220,N_13449);
or U13748 (N_13748,N_13254,N_13246);
nand U13749 (N_13749,N_13222,N_13370);
or U13750 (N_13750,N_13274,N_13483);
or U13751 (N_13751,N_13406,N_13490);
or U13752 (N_13752,N_13464,N_13247);
nor U13753 (N_13753,N_13540,N_13460);
nor U13754 (N_13754,N_13242,N_13546);
nor U13755 (N_13755,N_13392,N_13563);
nor U13756 (N_13756,N_13280,N_13275);
or U13757 (N_13757,N_13209,N_13478);
xor U13758 (N_13758,N_13583,N_13283);
and U13759 (N_13759,N_13240,N_13596);
nand U13760 (N_13760,N_13307,N_13377);
nor U13761 (N_13761,N_13216,N_13349);
or U13762 (N_13762,N_13277,N_13329);
nand U13763 (N_13763,N_13286,N_13500);
or U13764 (N_13764,N_13229,N_13226);
nor U13765 (N_13765,N_13513,N_13470);
nor U13766 (N_13766,N_13580,N_13384);
nor U13767 (N_13767,N_13378,N_13234);
nand U13768 (N_13768,N_13421,N_13522);
and U13769 (N_13769,N_13281,N_13205);
and U13770 (N_13770,N_13581,N_13316);
nor U13771 (N_13771,N_13346,N_13401);
xor U13772 (N_13772,N_13514,N_13264);
and U13773 (N_13773,N_13445,N_13394);
nor U13774 (N_13774,N_13387,N_13256);
nor U13775 (N_13775,N_13469,N_13537);
nand U13776 (N_13776,N_13326,N_13257);
and U13777 (N_13777,N_13577,N_13289);
nor U13778 (N_13778,N_13291,N_13482);
nor U13779 (N_13779,N_13457,N_13414);
nor U13780 (N_13780,N_13412,N_13272);
xnor U13781 (N_13781,N_13489,N_13201);
nor U13782 (N_13782,N_13376,N_13206);
and U13783 (N_13783,N_13227,N_13534);
or U13784 (N_13784,N_13382,N_13560);
xnor U13785 (N_13785,N_13364,N_13314);
xor U13786 (N_13786,N_13219,N_13347);
nand U13787 (N_13787,N_13592,N_13304);
nand U13788 (N_13788,N_13403,N_13335);
or U13789 (N_13789,N_13598,N_13405);
nand U13790 (N_13790,N_13315,N_13211);
or U13791 (N_13791,N_13338,N_13595);
or U13792 (N_13792,N_13426,N_13431);
nor U13793 (N_13793,N_13348,N_13559);
xor U13794 (N_13794,N_13237,N_13224);
nor U13795 (N_13795,N_13301,N_13244);
or U13796 (N_13796,N_13327,N_13484);
nor U13797 (N_13797,N_13320,N_13293);
or U13798 (N_13798,N_13461,N_13323);
nor U13799 (N_13799,N_13455,N_13366);
xnor U13800 (N_13800,N_13389,N_13490);
xnor U13801 (N_13801,N_13444,N_13336);
nand U13802 (N_13802,N_13559,N_13316);
nor U13803 (N_13803,N_13432,N_13378);
or U13804 (N_13804,N_13456,N_13384);
nor U13805 (N_13805,N_13493,N_13252);
or U13806 (N_13806,N_13211,N_13303);
nor U13807 (N_13807,N_13225,N_13323);
nor U13808 (N_13808,N_13480,N_13254);
or U13809 (N_13809,N_13472,N_13234);
xor U13810 (N_13810,N_13342,N_13220);
nor U13811 (N_13811,N_13514,N_13289);
and U13812 (N_13812,N_13213,N_13285);
xor U13813 (N_13813,N_13546,N_13477);
xnor U13814 (N_13814,N_13537,N_13545);
nand U13815 (N_13815,N_13581,N_13240);
xor U13816 (N_13816,N_13246,N_13523);
xor U13817 (N_13817,N_13350,N_13470);
nand U13818 (N_13818,N_13490,N_13529);
nand U13819 (N_13819,N_13424,N_13390);
nor U13820 (N_13820,N_13225,N_13439);
nor U13821 (N_13821,N_13307,N_13469);
and U13822 (N_13822,N_13445,N_13503);
nand U13823 (N_13823,N_13372,N_13343);
and U13824 (N_13824,N_13364,N_13329);
xnor U13825 (N_13825,N_13573,N_13547);
nor U13826 (N_13826,N_13583,N_13308);
nand U13827 (N_13827,N_13371,N_13478);
and U13828 (N_13828,N_13401,N_13579);
xnor U13829 (N_13829,N_13513,N_13474);
or U13830 (N_13830,N_13506,N_13511);
xnor U13831 (N_13831,N_13524,N_13225);
or U13832 (N_13832,N_13535,N_13294);
and U13833 (N_13833,N_13248,N_13243);
nand U13834 (N_13834,N_13314,N_13301);
and U13835 (N_13835,N_13589,N_13277);
and U13836 (N_13836,N_13222,N_13407);
nor U13837 (N_13837,N_13543,N_13213);
or U13838 (N_13838,N_13382,N_13232);
xnor U13839 (N_13839,N_13349,N_13334);
or U13840 (N_13840,N_13253,N_13244);
or U13841 (N_13841,N_13353,N_13382);
or U13842 (N_13842,N_13540,N_13519);
nand U13843 (N_13843,N_13435,N_13451);
or U13844 (N_13844,N_13453,N_13596);
xor U13845 (N_13845,N_13324,N_13421);
xnor U13846 (N_13846,N_13264,N_13467);
nor U13847 (N_13847,N_13386,N_13432);
and U13848 (N_13848,N_13590,N_13290);
nand U13849 (N_13849,N_13356,N_13206);
or U13850 (N_13850,N_13420,N_13290);
or U13851 (N_13851,N_13412,N_13203);
and U13852 (N_13852,N_13455,N_13364);
nand U13853 (N_13853,N_13578,N_13415);
or U13854 (N_13854,N_13522,N_13578);
nor U13855 (N_13855,N_13232,N_13373);
xnor U13856 (N_13856,N_13588,N_13342);
nand U13857 (N_13857,N_13468,N_13276);
nor U13858 (N_13858,N_13496,N_13231);
or U13859 (N_13859,N_13224,N_13242);
xnor U13860 (N_13860,N_13456,N_13217);
nand U13861 (N_13861,N_13350,N_13225);
nand U13862 (N_13862,N_13547,N_13398);
xnor U13863 (N_13863,N_13412,N_13540);
xnor U13864 (N_13864,N_13566,N_13347);
and U13865 (N_13865,N_13382,N_13447);
or U13866 (N_13866,N_13522,N_13228);
xor U13867 (N_13867,N_13423,N_13437);
or U13868 (N_13868,N_13277,N_13322);
nor U13869 (N_13869,N_13415,N_13503);
or U13870 (N_13870,N_13419,N_13374);
xor U13871 (N_13871,N_13224,N_13348);
xor U13872 (N_13872,N_13388,N_13454);
nor U13873 (N_13873,N_13370,N_13207);
nor U13874 (N_13874,N_13541,N_13445);
or U13875 (N_13875,N_13380,N_13475);
and U13876 (N_13876,N_13413,N_13474);
xnor U13877 (N_13877,N_13236,N_13334);
xor U13878 (N_13878,N_13382,N_13407);
and U13879 (N_13879,N_13449,N_13223);
nand U13880 (N_13880,N_13419,N_13577);
xnor U13881 (N_13881,N_13371,N_13583);
or U13882 (N_13882,N_13415,N_13510);
nand U13883 (N_13883,N_13502,N_13558);
and U13884 (N_13884,N_13296,N_13364);
xnor U13885 (N_13885,N_13344,N_13350);
xnor U13886 (N_13886,N_13207,N_13231);
and U13887 (N_13887,N_13287,N_13328);
nor U13888 (N_13888,N_13434,N_13580);
xnor U13889 (N_13889,N_13437,N_13390);
nor U13890 (N_13890,N_13584,N_13228);
nor U13891 (N_13891,N_13530,N_13411);
nor U13892 (N_13892,N_13326,N_13221);
or U13893 (N_13893,N_13319,N_13547);
nor U13894 (N_13894,N_13493,N_13516);
nand U13895 (N_13895,N_13489,N_13321);
and U13896 (N_13896,N_13278,N_13481);
and U13897 (N_13897,N_13551,N_13540);
and U13898 (N_13898,N_13410,N_13511);
nand U13899 (N_13899,N_13492,N_13537);
nand U13900 (N_13900,N_13260,N_13553);
nand U13901 (N_13901,N_13248,N_13391);
or U13902 (N_13902,N_13509,N_13257);
nand U13903 (N_13903,N_13438,N_13267);
nand U13904 (N_13904,N_13424,N_13211);
xor U13905 (N_13905,N_13305,N_13211);
nor U13906 (N_13906,N_13576,N_13494);
and U13907 (N_13907,N_13551,N_13322);
or U13908 (N_13908,N_13524,N_13309);
nand U13909 (N_13909,N_13226,N_13306);
or U13910 (N_13910,N_13399,N_13339);
or U13911 (N_13911,N_13508,N_13287);
and U13912 (N_13912,N_13262,N_13426);
nor U13913 (N_13913,N_13464,N_13306);
and U13914 (N_13914,N_13437,N_13590);
xnor U13915 (N_13915,N_13231,N_13378);
nor U13916 (N_13916,N_13270,N_13298);
xnor U13917 (N_13917,N_13419,N_13495);
xor U13918 (N_13918,N_13261,N_13454);
nor U13919 (N_13919,N_13467,N_13469);
and U13920 (N_13920,N_13380,N_13256);
or U13921 (N_13921,N_13414,N_13251);
and U13922 (N_13922,N_13313,N_13566);
and U13923 (N_13923,N_13520,N_13345);
and U13924 (N_13924,N_13369,N_13218);
or U13925 (N_13925,N_13267,N_13338);
xnor U13926 (N_13926,N_13377,N_13581);
xnor U13927 (N_13927,N_13252,N_13507);
xnor U13928 (N_13928,N_13275,N_13231);
nor U13929 (N_13929,N_13222,N_13596);
nand U13930 (N_13930,N_13488,N_13541);
nand U13931 (N_13931,N_13428,N_13340);
xor U13932 (N_13932,N_13495,N_13221);
or U13933 (N_13933,N_13307,N_13252);
nand U13934 (N_13934,N_13431,N_13536);
and U13935 (N_13935,N_13318,N_13426);
xor U13936 (N_13936,N_13569,N_13446);
and U13937 (N_13937,N_13222,N_13237);
nand U13938 (N_13938,N_13507,N_13582);
xnor U13939 (N_13939,N_13479,N_13464);
and U13940 (N_13940,N_13421,N_13349);
nor U13941 (N_13941,N_13532,N_13488);
and U13942 (N_13942,N_13540,N_13585);
nor U13943 (N_13943,N_13233,N_13529);
or U13944 (N_13944,N_13205,N_13527);
nand U13945 (N_13945,N_13381,N_13501);
xnor U13946 (N_13946,N_13222,N_13442);
and U13947 (N_13947,N_13593,N_13350);
and U13948 (N_13948,N_13448,N_13383);
or U13949 (N_13949,N_13595,N_13268);
nor U13950 (N_13950,N_13331,N_13221);
or U13951 (N_13951,N_13519,N_13504);
or U13952 (N_13952,N_13390,N_13409);
nand U13953 (N_13953,N_13211,N_13346);
or U13954 (N_13954,N_13288,N_13338);
nor U13955 (N_13955,N_13573,N_13533);
nand U13956 (N_13956,N_13589,N_13340);
or U13957 (N_13957,N_13299,N_13360);
or U13958 (N_13958,N_13309,N_13519);
nor U13959 (N_13959,N_13519,N_13478);
and U13960 (N_13960,N_13279,N_13506);
nor U13961 (N_13961,N_13321,N_13442);
or U13962 (N_13962,N_13560,N_13310);
or U13963 (N_13963,N_13256,N_13368);
nor U13964 (N_13964,N_13266,N_13253);
xnor U13965 (N_13965,N_13311,N_13437);
nor U13966 (N_13966,N_13350,N_13571);
nor U13967 (N_13967,N_13566,N_13222);
xor U13968 (N_13968,N_13491,N_13564);
and U13969 (N_13969,N_13486,N_13351);
nor U13970 (N_13970,N_13207,N_13529);
nor U13971 (N_13971,N_13579,N_13371);
and U13972 (N_13972,N_13328,N_13429);
nor U13973 (N_13973,N_13339,N_13578);
and U13974 (N_13974,N_13283,N_13416);
xnor U13975 (N_13975,N_13305,N_13511);
nand U13976 (N_13976,N_13519,N_13537);
or U13977 (N_13977,N_13343,N_13316);
nand U13978 (N_13978,N_13229,N_13438);
nand U13979 (N_13979,N_13445,N_13348);
xor U13980 (N_13980,N_13564,N_13539);
and U13981 (N_13981,N_13408,N_13470);
nand U13982 (N_13982,N_13250,N_13452);
or U13983 (N_13983,N_13588,N_13252);
xor U13984 (N_13984,N_13410,N_13588);
or U13985 (N_13985,N_13245,N_13539);
or U13986 (N_13986,N_13573,N_13512);
xnor U13987 (N_13987,N_13205,N_13320);
or U13988 (N_13988,N_13281,N_13399);
nor U13989 (N_13989,N_13279,N_13337);
nor U13990 (N_13990,N_13597,N_13258);
nor U13991 (N_13991,N_13559,N_13498);
and U13992 (N_13992,N_13239,N_13376);
nor U13993 (N_13993,N_13218,N_13375);
and U13994 (N_13994,N_13517,N_13367);
and U13995 (N_13995,N_13274,N_13530);
xnor U13996 (N_13996,N_13521,N_13208);
or U13997 (N_13997,N_13267,N_13476);
or U13998 (N_13998,N_13555,N_13250);
nor U13999 (N_13999,N_13275,N_13247);
nand U14000 (N_14000,N_13705,N_13856);
nand U14001 (N_14001,N_13918,N_13946);
nor U14002 (N_14002,N_13684,N_13879);
or U14003 (N_14003,N_13955,N_13672);
nand U14004 (N_14004,N_13942,N_13891);
nand U14005 (N_14005,N_13709,N_13881);
nor U14006 (N_14006,N_13952,N_13887);
xor U14007 (N_14007,N_13602,N_13744);
nand U14008 (N_14008,N_13653,N_13851);
nand U14009 (N_14009,N_13944,N_13817);
and U14010 (N_14010,N_13808,N_13896);
nand U14011 (N_14011,N_13658,N_13953);
nor U14012 (N_14012,N_13876,N_13917);
nor U14013 (N_14013,N_13991,N_13604);
or U14014 (N_14014,N_13877,N_13642);
nand U14015 (N_14015,N_13872,N_13628);
nor U14016 (N_14016,N_13692,N_13833);
or U14017 (N_14017,N_13816,N_13957);
and U14018 (N_14018,N_13906,N_13893);
xor U14019 (N_14019,N_13689,N_13998);
nor U14020 (N_14020,N_13741,N_13683);
or U14021 (N_14021,N_13976,N_13737);
and U14022 (N_14022,N_13646,N_13791);
xnor U14023 (N_14023,N_13787,N_13871);
and U14024 (N_14024,N_13948,N_13974);
xor U14025 (N_14025,N_13987,N_13822);
nand U14026 (N_14026,N_13753,N_13912);
and U14027 (N_14027,N_13936,N_13751);
and U14028 (N_14028,N_13983,N_13885);
xnor U14029 (N_14029,N_13864,N_13660);
and U14030 (N_14030,N_13767,N_13812);
and U14031 (N_14031,N_13947,N_13854);
and U14032 (N_14032,N_13675,N_13824);
or U14033 (N_14033,N_13670,N_13711);
nor U14034 (N_14034,N_13650,N_13779);
nor U14035 (N_14035,N_13723,N_13913);
xnor U14036 (N_14036,N_13997,N_13632);
nand U14037 (N_14037,N_13874,N_13752);
nand U14038 (N_14038,N_13810,N_13908);
nor U14039 (N_14039,N_13710,N_13659);
or U14040 (N_14040,N_13849,N_13673);
and U14041 (N_14041,N_13732,N_13820);
nor U14042 (N_14042,N_13743,N_13621);
nand U14043 (N_14043,N_13803,N_13749);
and U14044 (N_14044,N_13636,N_13964);
nand U14045 (N_14045,N_13631,N_13927);
nand U14046 (N_14046,N_13719,N_13839);
nor U14047 (N_14047,N_13725,N_13759);
or U14048 (N_14048,N_13645,N_13622);
nor U14049 (N_14049,N_13933,N_13866);
xnor U14050 (N_14050,N_13882,N_13657);
nand U14051 (N_14051,N_13625,N_13905);
or U14052 (N_14052,N_13945,N_13786);
nand U14053 (N_14053,N_13935,N_13720);
and U14054 (N_14054,N_13995,N_13931);
nor U14055 (N_14055,N_13682,N_13959);
nand U14056 (N_14056,N_13788,N_13669);
and U14057 (N_14057,N_13618,N_13686);
nor U14058 (N_14058,N_13716,N_13921);
nand U14059 (N_14059,N_13643,N_13920);
and U14060 (N_14060,N_13766,N_13815);
and U14061 (N_14061,N_13823,N_13674);
xor U14062 (N_14062,N_13700,N_13761);
xor U14063 (N_14063,N_13956,N_13966);
nor U14064 (N_14064,N_13789,N_13601);
xnor U14065 (N_14065,N_13718,N_13870);
nor U14066 (N_14066,N_13855,N_13688);
or U14067 (N_14067,N_13765,N_13802);
and U14068 (N_14068,N_13755,N_13850);
and U14069 (N_14069,N_13985,N_13950);
nor U14070 (N_14070,N_13840,N_13616);
xnor U14071 (N_14071,N_13804,N_13704);
xor U14072 (N_14072,N_13728,N_13968);
nand U14073 (N_14073,N_13671,N_13600);
and U14074 (N_14074,N_13706,N_13825);
or U14075 (N_14075,N_13880,N_13760);
or U14076 (N_14076,N_13687,N_13769);
nand U14077 (N_14077,N_13649,N_13970);
xor U14078 (N_14078,N_13862,N_13681);
and U14079 (N_14079,N_13852,N_13980);
and U14080 (N_14080,N_13608,N_13969);
xnor U14081 (N_14081,N_13842,N_13781);
nand U14082 (N_14082,N_13731,N_13832);
nand U14083 (N_14083,N_13619,N_13774);
nor U14084 (N_14084,N_13735,N_13609);
nor U14085 (N_14085,N_13702,N_13606);
nand U14086 (N_14086,N_13984,N_13777);
xor U14087 (N_14087,N_13928,N_13610);
nor U14088 (N_14088,N_13975,N_13757);
xnor U14089 (N_14089,N_13865,N_13793);
nor U14090 (N_14090,N_13979,N_13932);
xor U14091 (N_14091,N_13798,N_13794);
nor U14092 (N_14092,N_13992,N_13834);
or U14093 (N_14093,N_13801,N_13693);
or U14094 (N_14094,N_13890,N_13626);
xor U14095 (N_14095,N_13750,N_13962);
nor U14096 (N_14096,N_13652,N_13916);
and U14097 (N_14097,N_13911,N_13973);
or U14098 (N_14098,N_13617,N_13667);
nand U14099 (N_14099,N_13897,N_13915);
xor U14100 (N_14100,N_13624,N_13678);
nand U14101 (N_14101,N_13635,N_13662);
or U14102 (N_14102,N_13857,N_13770);
nand U14103 (N_14103,N_13988,N_13961);
nand U14104 (N_14104,N_13640,N_13685);
nor U14105 (N_14105,N_13827,N_13758);
nand U14106 (N_14106,N_13813,N_13922);
and U14107 (N_14107,N_13986,N_13907);
nand U14108 (N_14108,N_13861,N_13811);
nand U14109 (N_14109,N_13892,N_13754);
nand U14110 (N_14110,N_13698,N_13809);
and U14111 (N_14111,N_13796,N_13795);
nor U14112 (N_14112,N_13745,N_13613);
and U14113 (N_14113,N_13846,N_13886);
and U14114 (N_14114,N_13696,N_13638);
nand U14115 (N_14115,N_13665,N_13994);
or U14116 (N_14116,N_13859,N_13763);
or U14117 (N_14117,N_13776,N_13848);
nor U14118 (N_14118,N_13806,N_13620);
and U14119 (N_14119,N_13903,N_13900);
nand U14120 (N_14120,N_13972,N_13836);
or U14121 (N_14121,N_13703,N_13895);
or U14122 (N_14122,N_13629,N_13694);
nor U14123 (N_14123,N_13762,N_13925);
xor U14124 (N_14124,N_13778,N_13785);
and U14125 (N_14125,N_13965,N_13889);
nand U14126 (N_14126,N_13847,N_13989);
xor U14127 (N_14127,N_13899,N_13826);
or U14128 (N_14128,N_13722,N_13829);
nand U14129 (N_14129,N_13612,N_13873);
nand U14130 (N_14130,N_13938,N_13614);
xor U14131 (N_14131,N_13734,N_13999);
or U14132 (N_14132,N_13884,N_13726);
and U14133 (N_14133,N_13783,N_13981);
xor U14134 (N_14134,N_13923,N_13990);
nor U14135 (N_14135,N_13963,N_13715);
and U14136 (N_14136,N_13843,N_13739);
xor U14137 (N_14137,N_13663,N_13902);
and U14138 (N_14138,N_13771,N_13792);
nor U14139 (N_14139,N_13875,N_13883);
xor U14140 (N_14140,N_13831,N_13853);
nor U14141 (N_14141,N_13863,N_13647);
or U14142 (N_14142,N_13742,N_13951);
nand U14143 (N_14143,N_13637,N_13747);
nor U14144 (N_14144,N_13943,N_13828);
xnor U14145 (N_14145,N_13666,N_13627);
or U14146 (N_14146,N_13756,N_13837);
and U14147 (N_14147,N_13708,N_13634);
nor U14148 (N_14148,N_13651,N_13699);
or U14149 (N_14149,N_13707,N_13830);
and U14150 (N_14150,N_13654,N_13838);
nand U14151 (N_14151,N_13679,N_13910);
and U14152 (N_14152,N_13867,N_13639);
nand U14153 (N_14153,N_13814,N_13717);
xor U14154 (N_14154,N_13971,N_13784);
and U14155 (N_14155,N_13958,N_13929);
nor U14156 (N_14156,N_13605,N_13901);
xor U14157 (N_14157,N_13691,N_13697);
or U14158 (N_14158,N_13941,N_13695);
xnor U14159 (N_14159,N_13648,N_13615);
and U14160 (N_14160,N_13819,N_13655);
or U14161 (N_14161,N_13775,N_13919);
nor U14162 (N_14162,N_13712,N_13714);
xor U14163 (N_14163,N_13939,N_13926);
or U14164 (N_14164,N_13841,N_13729);
or U14165 (N_14165,N_13733,N_13730);
and U14166 (N_14166,N_13677,N_13644);
nand U14167 (N_14167,N_13940,N_13821);
nand U14168 (N_14168,N_13878,N_13797);
or U14169 (N_14169,N_13680,N_13860);
nand U14170 (N_14170,N_13954,N_13930);
nand U14171 (N_14171,N_13676,N_13937);
or U14172 (N_14172,N_13713,N_13967);
xnor U14173 (N_14173,N_13835,N_13934);
xnor U14174 (N_14174,N_13924,N_13607);
or U14175 (N_14175,N_13982,N_13978);
or U14176 (N_14176,N_13630,N_13768);
or U14177 (N_14177,N_13960,N_13800);
or U14178 (N_14178,N_13888,N_13603);
and U14179 (N_14179,N_13799,N_13904);
nand U14180 (N_14180,N_13805,N_13738);
nand U14181 (N_14181,N_13664,N_13868);
nor U14182 (N_14182,N_13845,N_13949);
or U14183 (N_14183,N_13909,N_13656);
and U14184 (N_14184,N_13858,N_13724);
and U14185 (N_14185,N_13818,N_13764);
xnor U14186 (N_14186,N_13844,N_13746);
nor U14187 (N_14187,N_13772,N_13898);
or U14188 (N_14188,N_13914,N_13668);
and U14189 (N_14189,N_13727,N_13690);
and U14190 (N_14190,N_13623,N_13993);
or U14191 (N_14191,N_13894,N_13641);
nand U14192 (N_14192,N_13748,N_13611);
xnor U14193 (N_14193,N_13807,N_13790);
xor U14194 (N_14194,N_13661,N_13721);
nor U14195 (N_14195,N_13740,N_13701);
and U14196 (N_14196,N_13782,N_13736);
and U14197 (N_14197,N_13996,N_13977);
nand U14198 (N_14198,N_13633,N_13780);
and U14199 (N_14199,N_13869,N_13773);
or U14200 (N_14200,N_13812,N_13721);
or U14201 (N_14201,N_13633,N_13727);
nor U14202 (N_14202,N_13697,N_13674);
nor U14203 (N_14203,N_13804,N_13758);
xnor U14204 (N_14204,N_13948,N_13793);
nor U14205 (N_14205,N_13752,N_13628);
nor U14206 (N_14206,N_13901,N_13916);
nor U14207 (N_14207,N_13987,N_13755);
xor U14208 (N_14208,N_13955,N_13764);
and U14209 (N_14209,N_13852,N_13630);
nand U14210 (N_14210,N_13993,N_13921);
and U14211 (N_14211,N_13945,N_13984);
and U14212 (N_14212,N_13880,N_13865);
or U14213 (N_14213,N_13742,N_13852);
and U14214 (N_14214,N_13875,N_13612);
xnor U14215 (N_14215,N_13998,N_13996);
xnor U14216 (N_14216,N_13865,N_13841);
and U14217 (N_14217,N_13753,N_13614);
xnor U14218 (N_14218,N_13944,N_13784);
nand U14219 (N_14219,N_13885,N_13938);
nand U14220 (N_14220,N_13654,N_13751);
or U14221 (N_14221,N_13813,N_13619);
xnor U14222 (N_14222,N_13929,N_13750);
and U14223 (N_14223,N_13737,N_13906);
nor U14224 (N_14224,N_13748,N_13947);
xor U14225 (N_14225,N_13778,N_13998);
nand U14226 (N_14226,N_13874,N_13668);
nor U14227 (N_14227,N_13709,N_13775);
xnor U14228 (N_14228,N_13693,N_13696);
nor U14229 (N_14229,N_13799,N_13778);
or U14230 (N_14230,N_13820,N_13681);
and U14231 (N_14231,N_13935,N_13924);
and U14232 (N_14232,N_13614,N_13744);
xor U14233 (N_14233,N_13918,N_13834);
nand U14234 (N_14234,N_13902,N_13724);
and U14235 (N_14235,N_13970,N_13884);
xnor U14236 (N_14236,N_13965,N_13857);
or U14237 (N_14237,N_13878,N_13766);
and U14238 (N_14238,N_13891,N_13844);
and U14239 (N_14239,N_13999,N_13909);
nor U14240 (N_14240,N_13740,N_13954);
xor U14241 (N_14241,N_13983,N_13795);
or U14242 (N_14242,N_13883,N_13700);
nand U14243 (N_14243,N_13964,N_13806);
nor U14244 (N_14244,N_13927,N_13820);
nand U14245 (N_14245,N_13717,N_13970);
nand U14246 (N_14246,N_13925,N_13606);
nand U14247 (N_14247,N_13742,N_13672);
or U14248 (N_14248,N_13970,N_13810);
or U14249 (N_14249,N_13812,N_13820);
nor U14250 (N_14250,N_13903,N_13673);
or U14251 (N_14251,N_13722,N_13901);
nand U14252 (N_14252,N_13978,N_13772);
or U14253 (N_14253,N_13652,N_13882);
nor U14254 (N_14254,N_13733,N_13681);
or U14255 (N_14255,N_13839,N_13985);
nand U14256 (N_14256,N_13618,N_13726);
or U14257 (N_14257,N_13881,N_13851);
xor U14258 (N_14258,N_13930,N_13992);
or U14259 (N_14259,N_13829,N_13669);
nor U14260 (N_14260,N_13659,N_13862);
or U14261 (N_14261,N_13822,N_13883);
xor U14262 (N_14262,N_13936,N_13729);
and U14263 (N_14263,N_13742,N_13945);
nor U14264 (N_14264,N_13937,N_13822);
nand U14265 (N_14265,N_13656,N_13862);
xor U14266 (N_14266,N_13720,N_13840);
or U14267 (N_14267,N_13831,N_13747);
nand U14268 (N_14268,N_13646,N_13872);
or U14269 (N_14269,N_13905,N_13603);
or U14270 (N_14270,N_13836,N_13621);
nor U14271 (N_14271,N_13720,N_13905);
and U14272 (N_14272,N_13753,N_13716);
nand U14273 (N_14273,N_13847,N_13802);
or U14274 (N_14274,N_13631,N_13612);
nand U14275 (N_14275,N_13956,N_13671);
or U14276 (N_14276,N_13936,N_13602);
or U14277 (N_14277,N_13762,N_13618);
nand U14278 (N_14278,N_13905,N_13750);
xnor U14279 (N_14279,N_13909,N_13762);
xor U14280 (N_14280,N_13864,N_13633);
and U14281 (N_14281,N_13880,N_13972);
xor U14282 (N_14282,N_13885,N_13770);
nand U14283 (N_14283,N_13857,N_13980);
and U14284 (N_14284,N_13867,N_13910);
nand U14285 (N_14285,N_13808,N_13608);
xor U14286 (N_14286,N_13659,N_13831);
nand U14287 (N_14287,N_13997,N_13746);
nand U14288 (N_14288,N_13789,N_13987);
and U14289 (N_14289,N_13798,N_13967);
or U14290 (N_14290,N_13869,N_13812);
nor U14291 (N_14291,N_13668,N_13719);
and U14292 (N_14292,N_13806,N_13791);
and U14293 (N_14293,N_13694,N_13627);
and U14294 (N_14294,N_13843,N_13889);
and U14295 (N_14295,N_13833,N_13785);
xnor U14296 (N_14296,N_13720,N_13873);
and U14297 (N_14297,N_13938,N_13631);
nor U14298 (N_14298,N_13748,N_13811);
nand U14299 (N_14299,N_13600,N_13952);
and U14300 (N_14300,N_13845,N_13884);
or U14301 (N_14301,N_13756,N_13997);
and U14302 (N_14302,N_13735,N_13705);
or U14303 (N_14303,N_13977,N_13757);
nor U14304 (N_14304,N_13878,N_13992);
or U14305 (N_14305,N_13773,N_13871);
nand U14306 (N_14306,N_13870,N_13656);
nor U14307 (N_14307,N_13882,N_13791);
or U14308 (N_14308,N_13990,N_13985);
nand U14309 (N_14309,N_13683,N_13994);
or U14310 (N_14310,N_13910,N_13896);
and U14311 (N_14311,N_13778,N_13777);
nand U14312 (N_14312,N_13915,N_13934);
and U14313 (N_14313,N_13679,N_13927);
xnor U14314 (N_14314,N_13771,N_13661);
and U14315 (N_14315,N_13894,N_13710);
xnor U14316 (N_14316,N_13872,N_13790);
and U14317 (N_14317,N_13801,N_13996);
nand U14318 (N_14318,N_13823,N_13653);
and U14319 (N_14319,N_13868,N_13754);
xnor U14320 (N_14320,N_13708,N_13619);
or U14321 (N_14321,N_13609,N_13726);
nor U14322 (N_14322,N_13639,N_13726);
nor U14323 (N_14323,N_13654,N_13948);
or U14324 (N_14324,N_13640,N_13686);
nor U14325 (N_14325,N_13678,N_13888);
or U14326 (N_14326,N_13717,N_13710);
nor U14327 (N_14327,N_13812,N_13705);
xor U14328 (N_14328,N_13891,N_13693);
nand U14329 (N_14329,N_13651,N_13721);
xor U14330 (N_14330,N_13850,N_13905);
and U14331 (N_14331,N_13808,N_13926);
xnor U14332 (N_14332,N_13816,N_13702);
or U14333 (N_14333,N_13659,N_13935);
nand U14334 (N_14334,N_13989,N_13676);
nor U14335 (N_14335,N_13985,N_13862);
and U14336 (N_14336,N_13670,N_13741);
nor U14337 (N_14337,N_13963,N_13810);
xor U14338 (N_14338,N_13996,N_13822);
xor U14339 (N_14339,N_13966,N_13918);
and U14340 (N_14340,N_13738,N_13679);
xor U14341 (N_14341,N_13656,N_13707);
and U14342 (N_14342,N_13703,N_13956);
nand U14343 (N_14343,N_13932,N_13854);
xnor U14344 (N_14344,N_13713,N_13925);
and U14345 (N_14345,N_13817,N_13913);
nor U14346 (N_14346,N_13821,N_13666);
nand U14347 (N_14347,N_13944,N_13899);
nor U14348 (N_14348,N_13805,N_13690);
nand U14349 (N_14349,N_13687,N_13689);
or U14350 (N_14350,N_13606,N_13891);
and U14351 (N_14351,N_13998,N_13846);
and U14352 (N_14352,N_13824,N_13935);
or U14353 (N_14353,N_13900,N_13656);
or U14354 (N_14354,N_13800,N_13974);
nor U14355 (N_14355,N_13785,N_13652);
and U14356 (N_14356,N_13715,N_13832);
or U14357 (N_14357,N_13792,N_13640);
xor U14358 (N_14358,N_13923,N_13784);
nor U14359 (N_14359,N_13919,N_13912);
nor U14360 (N_14360,N_13608,N_13904);
and U14361 (N_14361,N_13647,N_13815);
xnor U14362 (N_14362,N_13861,N_13756);
or U14363 (N_14363,N_13678,N_13683);
xnor U14364 (N_14364,N_13668,N_13747);
nand U14365 (N_14365,N_13920,N_13993);
nor U14366 (N_14366,N_13930,N_13890);
or U14367 (N_14367,N_13811,N_13818);
and U14368 (N_14368,N_13633,N_13717);
xnor U14369 (N_14369,N_13744,N_13955);
and U14370 (N_14370,N_13647,N_13931);
or U14371 (N_14371,N_13989,N_13877);
nand U14372 (N_14372,N_13877,N_13651);
nor U14373 (N_14373,N_13790,N_13841);
or U14374 (N_14374,N_13900,N_13890);
nand U14375 (N_14375,N_13769,N_13886);
and U14376 (N_14376,N_13752,N_13814);
nor U14377 (N_14377,N_13932,N_13831);
nor U14378 (N_14378,N_13665,N_13902);
xnor U14379 (N_14379,N_13837,N_13672);
xnor U14380 (N_14380,N_13623,N_13881);
xnor U14381 (N_14381,N_13964,N_13776);
nand U14382 (N_14382,N_13652,N_13670);
nand U14383 (N_14383,N_13909,N_13625);
nand U14384 (N_14384,N_13626,N_13609);
or U14385 (N_14385,N_13654,N_13866);
nand U14386 (N_14386,N_13969,N_13834);
xor U14387 (N_14387,N_13790,N_13779);
and U14388 (N_14388,N_13706,N_13639);
nand U14389 (N_14389,N_13697,N_13741);
and U14390 (N_14390,N_13677,N_13911);
xnor U14391 (N_14391,N_13810,N_13603);
or U14392 (N_14392,N_13601,N_13783);
or U14393 (N_14393,N_13646,N_13744);
nor U14394 (N_14394,N_13764,N_13911);
or U14395 (N_14395,N_13676,N_13875);
or U14396 (N_14396,N_13960,N_13645);
xnor U14397 (N_14397,N_13653,N_13854);
xnor U14398 (N_14398,N_13703,N_13745);
and U14399 (N_14399,N_13693,N_13812);
xor U14400 (N_14400,N_14236,N_14316);
nand U14401 (N_14401,N_14284,N_14078);
nand U14402 (N_14402,N_14358,N_14266);
or U14403 (N_14403,N_14228,N_14354);
or U14404 (N_14404,N_14116,N_14250);
or U14405 (N_14405,N_14083,N_14291);
or U14406 (N_14406,N_14375,N_14085);
xor U14407 (N_14407,N_14052,N_14339);
xnor U14408 (N_14408,N_14158,N_14245);
nand U14409 (N_14409,N_14209,N_14023);
xor U14410 (N_14410,N_14148,N_14094);
or U14411 (N_14411,N_14025,N_14383);
nand U14412 (N_14412,N_14002,N_14252);
nand U14413 (N_14413,N_14041,N_14362);
xor U14414 (N_14414,N_14243,N_14292);
nor U14415 (N_14415,N_14013,N_14214);
xor U14416 (N_14416,N_14318,N_14264);
nor U14417 (N_14417,N_14399,N_14283);
nor U14418 (N_14418,N_14035,N_14242);
and U14419 (N_14419,N_14056,N_14086);
nand U14420 (N_14420,N_14332,N_14281);
or U14421 (N_14421,N_14377,N_14040);
or U14422 (N_14422,N_14247,N_14215);
or U14423 (N_14423,N_14396,N_14326);
nand U14424 (N_14424,N_14033,N_14238);
or U14425 (N_14425,N_14046,N_14182);
and U14426 (N_14426,N_14343,N_14066);
or U14427 (N_14427,N_14299,N_14100);
nor U14428 (N_14428,N_14196,N_14153);
or U14429 (N_14429,N_14384,N_14123);
nand U14430 (N_14430,N_14061,N_14268);
and U14431 (N_14431,N_14072,N_14122);
and U14432 (N_14432,N_14135,N_14230);
and U14433 (N_14433,N_14051,N_14007);
or U14434 (N_14434,N_14234,N_14350);
nand U14435 (N_14435,N_14109,N_14068);
or U14436 (N_14436,N_14212,N_14095);
nand U14437 (N_14437,N_14315,N_14322);
nand U14438 (N_14438,N_14165,N_14314);
xnor U14439 (N_14439,N_14357,N_14003);
nor U14440 (N_14440,N_14352,N_14075);
nand U14441 (N_14441,N_14019,N_14138);
xnor U14442 (N_14442,N_14269,N_14192);
and U14443 (N_14443,N_14210,N_14296);
or U14444 (N_14444,N_14270,N_14047);
xnor U14445 (N_14445,N_14126,N_14156);
xor U14446 (N_14446,N_14336,N_14239);
and U14447 (N_14447,N_14166,N_14379);
and U14448 (N_14448,N_14278,N_14128);
nand U14449 (N_14449,N_14330,N_14275);
nand U14450 (N_14450,N_14170,N_14004);
xnor U14451 (N_14451,N_14331,N_14162);
nor U14452 (N_14452,N_14053,N_14241);
or U14453 (N_14453,N_14325,N_14254);
and U14454 (N_14454,N_14172,N_14089);
nor U14455 (N_14455,N_14273,N_14258);
or U14456 (N_14456,N_14308,N_14074);
xor U14457 (N_14457,N_14137,N_14108);
nor U14458 (N_14458,N_14136,N_14261);
xnor U14459 (N_14459,N_14161,N_14342);
nor U14460 (N_14460,N_14092,N_14351);
or U14461 (N_14461,N_14240,N_14310);
nor U14462 (N_14462,N_14029,N_14297);
nand U14463 (N_14463,N_14371,N_14050);
nand U14464 (N_14464,N_14285,N_14082);
or U14465 (N_14465,N_14012,N_14253);
and U14466 (N_14466,N_14014,N_14098);
nand U14467 (N_14467,N_14319,N_14144);
and U14468 (N_14468,N_14227,N_14361);
xor U14469 (N_14469,N_14114,N_14356);
xor U14470 (N_14470,N_14388,N_14080);
nand U14471 (N_14471,N_14305,N_14302);
xor U14472 (N_14472,N_14125,N_14101);
and U14473 (N_14473,N_14313,N_14244);
nand U14474 (N_14474,N_14341,N_14188);
and U14475 (N_14475,N_14304,N_14027);
nor U14476 (N_14476,N_14118,N_14367);
or U14477 (N_14477,N_14017,N_14380);
and U14478 (N_14478,N_14203,N_14088);
nand U14479 (N_14479,N_14191,N_14324);
and U14480 (N_14480,N_14286,N_14024);
nand U14481 (N_14481,N_14054,N_14199);
or U14482 (N_14482,N_14084,N_14360);
and U14483 (N_14483,N_14279,N_14001);
nand U14484 (N_14484,N_14186,N_14026);
and U14485 (N_14485,N_14171,N_14246);
nand U14486 (N_14486,N_14184,N_14366);
nand U14487 (N_14487,N_14251,N_14337);
nand U14488 (N_14488,N_14232,N_14364);
nor U14489 (N_14489,N_14201,N_14154);
nor U14490 (N_14490,N_14045,N_14229);
and U14491 (N_14491,N_14200,N_14179);
and U14492 (N_14492,N_14265,N_14398);
or U14493 (N_14493,N_14133,N_14376);
xor U14494 (N_14494,N_14290,N_14006);
nand U14495 (N_14495,N_14115,N_14222);
xnor U14496 (N_14496,N_14104,N_14204);
and U14497 (N_14497,N_14145,N_14022);
xnor U14498 (N_14498,N_14090,N_14120);
and U14499 (N_14499,N_14233,N_14225);
xnor U14500 (N_14500,N_14235,N_14231);
nor U14501 (N_14501,N_14363,N_14287);
or U14502 (N_14502,N_14187,N_14335);
and U14503 (N_14503,N_14217,N_14063);
nand U14504 (N_14504,N_14382,N_14065);
nand U14505 (N_14505,N_14119,N_14031);
xor U14506 (N_14506,N_14317,N_14130);
and U14507 (N_14507,N_14034,N_14106);
or U14508 (N_14508,N_14277,N_14077);
nor U14509 (N_14509,N_14000,N_14193);
or U14510 (N_14510,N_14005,N_14303);
nand U14511 (N_14511,N_14093,N_14271);
or U14512 (N_14512,N_14151,N_14345);
xnor U14513 (N_14513,N_14018,N_14211);
or U14514 (N_14514,N_14327,N_14195);
nand U14515 (N_14515,N_14394,N_14142);
and U14516 (N_14516,N_14346,N_14129);
and U14517 (N_14517,N_14015,N_14102);
xnor U14518 (N_14518,N_14389,N_14113);
or U14519 (N_14519,N_14349,N_14272);
nand U14520 (N_14520,N_14091,N_14174);
nand U14521 (N_14521,N_14307,N_14208);
nor U14522 (N_14522,N_14257,N_14152);
nor U14523 (N_14523,N_14057,N_14311);
and U14524 (N_14524,N_14218,N_14067);
xor U14525 (N_14525,N_14355,N_14062);
nor U14526 (N_14526,N_14016,N_14365);
nand U14527 (N_14527,N_14300,N_14373);
xor U14528 (N_14528,N_14219,N_14173);
nand U14529 (N_14529,N_14149,N_14030);
or U14530 (N_14530,N_14127,N_14096);
xnor U14531 (N_14531,N_14321,N_14385);
nand U14532 (N_14532,N_14185,N_14197);
or U14533 (N_14533,N_14180,N_14295);
xor U14534 (N_14534,N_14042,N_14160);
or U14535 (N_14535,N_14008,N_14392);
and U14536 (N_14536,N_14132,N_14039);
nor U14537 (N_14537,N_14028,N_14323);
or U14538 (N_14538,N_14395,N_14248);
xnor U14539 (N_14539,N_14255,N_14267);
xnor U14540 (N_14540,N_14155,N_14032);
and U14541 (N_14541,N_14070,N_14334);
nand U14542 (N_14542,N_14177,N_14205);
nand U14543 (N_14543,N_14181,N_14076);
xnor U14544 (N_14544,N_14221,N_14348);
nor U14545 (N_14545,N_14369,N_14058);
and U14546 (N_14546,N_14333,N_14393);
nand U14547 (N_14547,N_14298,N_14338);
nor U14548 (N_14548,N_14263,N_14198);
nand U14549 (N_14549,N_14274,N_14294);
and U14550 (N_14550,N_14011,N_14048);
nor U14551 (N_14551,N_14043,N_14381);
nand U14552 (N_14552,N_14293,N_14150);
or U14553 (N_14553,N_14167,N_14309);
nand U14554 (N_14554,N_14289,N_14260);
and U14555 (N_14555,N_14226,N_14259);
nand U14556 (N_14556,N_14194,N_14110);
nand U14557 (N_14557,N_14312,N_14157);
and U14558 (N_14558,N_14190,N_14347);
and U14559 (N_14559,N_14256,N_14372);
xor U14560 (N_14560,N_14140,N_14060);
nand U14561 (N_14561,N_14124,N_14071);
or U14562 (N_14562,N_14288,N_14036);
and U14563 (N_14563,N_14044,N_14378);
and U14564 (N_14564,N_14038,N_14390);
xnor U14565 (N_14565,N_14206,N_14069);
or U14566 (N_14566,N_14280,N_14134);
nor U14567 (N_14567,N_14021,N_14097);
nand U14568 (N_14568,N_14224,N_14131);
nand U14569 (N_14569,N_14175,N_14055);
xor U14570 (N_14570,N_14301,N_14163);
xnor U14571 (N_14571,N_14159,N_14237);
nand U14572 (N_14572,N_14249,N_14189);
or U14573 (N_14573,N_14282,N_14147);
xor U14574 (N_14574,N_14009,N_14387);
xnor U14575 (N_14575,N_14169,N_14183);
nand U14576 (N_14576,N_14168,N_14107);
nor U14577 (N_14577,N_14391,N_14202);
nand U14578 (N_14578,N_14099,N_14359);
or U14579 (N_14579,N_14105,N_14220);
and U14580 (N_14580,N_14353,N_14397);
or U14581 (N_14581,N_14117,N_14344);
nor U14582 (N_14582,N_14059,N_14176);
nor U14583 (N_14583,N_14146,N_14049);
xnor U14584 (N_14584,N_14073,N_14370);
and U14585 (N_14585,N_14037,N_14064);
nand U14586 (N_14586,N_14178,N_14139);
nor U14587 (N_14587,N_14328,N_14374);
or U14588 (N_14588,N_14213,N_14386);
nor U14589 (N_14589,N_14276,N_14103);
and U14590 (N_14590,N_14320,N_14010);
or U14591 (N_14591,N_14223,N_14121);
and U14592 (N_14592,N_14081,N_14329);
nor U14593 (N_14593,N_14020,N_14087);
or U14594 (N_14594,N_14141,N_14143);
nor U14595 (N_14595,N_14207,N_14340);
and U14596 (N_14596,N_14216,N_14368);
and U14597 (N_14597,N_14111,N_14306);
xnor U14598 (N_14598,N_14262,N_14164);
nand U14599 (N_14599,N_14112,N_14079);
and U14600 (N_14600,N_14376,N_14086);
or U14601 (N_14601,N_14060,N_14309);
nor U14602 (N_14602,N_14142,N_14386);
or U14603 (N_14603,N_14164,N_14026);
or U14604 (N_14604,N_14048,N_14352);
or U14605 (N_14605,N_14084,N_14087);
nor U14606 (N_14606,N_14235,N_14365);
nand U14607 (N_14607,N_14154,N_14149);
and U14608 (N_14608,N_14246,N_14008);
nand U14609 (N_14609,N_14071,N_14130);
and U14610 (N_14610,N_14057,N_14282);
nand U14611 (N_14611,N_14162,N_14157);
nor U14612 (N_14612,N_14231,N_14196);
and U14613 (N_14613,N_14199,N_14023);
xor U14614 (N_14614,N_14272,N_14228);
or U14615 (N_14615,N_14328,N_14155);
nor U14616 (N_14616,N_14128,N_14259);
and U14617 (N_14617,N_14318,N_14361);
xor U14618 (N_14618,N_14176,N_14386);
nor U14619 (N_14619,N_14112,N_14067);
or U14620 (N_14620,N_14227,N_14193);
nor U14621 (N_14621,N_14266,N_14311);
or U14622 (N_14622,N_14100,N_14297);
or U14623 (N_14623,N_14141,N_14064);
nand U14624 (N_14624,N_14204,N_14083);
nor U14625 (N_14625,N_14084,N_14191);
nor U14626 (N_14626,N_14316,N_14005);
or U14627 (N_14627,N_14087,N_14219);
xor U14628 (N_14628,N_14348,N_14090);
nand U14629 (N_14629,N_14258,N_14176);
or U14630 (N_14630,N_14257,N_14137);
nand U14631 (N_14631,N_14355,N_14284);
nand U14632 (N_14632,N_14247,N_14171);
nand U14633 (N_14633,N_14115,N_14084);
xnor U14634 (N_14634,N_14396,N_14220);
nor U14635 (N_14635,N_14293,N_14380);
xor U14636 (N_14636,N_14127,N_14062);
nand U14637 (N_14637,N_14301,N_14123);
nand U14638 (N_14638,N_14258,N_14195);
nand U14639 (N_14639,N_14085,N_14244);
and U14640 (N_14640,N_14349,N_14128);
and U14641 (N_14641,N_14160,N_14399);
nor U14642 (N_14642,N_14252,N_14137);
nand U14643 (N_14643,N_14383,N_14361);
nand U14644 (N_14644,N_14049,N_14150);
or U14645 (N_14645,N_14376,N_14347);
nand U14646 (N_14646,N_14030,N_14055);
xnor U14647 (N_14647,N_14031,N_14375);
xor U14648 (N_14648,N_14001,N_14321);
nor U14649 (N_14649,N_14124,N_14099);
xor U14650 (N_14650,N_14065,N_14342);
and U14651 (N_14651,N_14034,N_14327);
nand U14652 (N_14652,N_14220,N_14231);
nand U14653 (N_14653,N_14183,N_14020);
nor U14654 (N_14654,N_14014,N_14230);
nor U14655 (N_14655,N_14216,N_14086);
nand U14656 (N_14656,N_14046,N_14194);
or U14657 (N_14657,N_14341,N_14010);
xor U14658 (N_14658,N_14182,N_14131);
and U14659 (N_14659,N_14179,N_14056);
or U14660 (N_14660,N_14078,N_14109);
nand U14661 (N_14661,N_14360,N_14006);
nor U14662 (N_14662,N_14053,N_14344);
xor U14663 (N_14663,N_14372,N_14255);
or U14664 (N_14664,N_14398,N_14354);
xor U14665 (N_14665,N_14350,N_14274);
and U14666 (N_14666,N_14295,N_14320);
or U14667 (N_14667,N_14218,N_14235);
nand U14668 (N_14668,N_14380,N_14206);
nor U14669 (N_14669,N_14132,N_14287);
nor U14670 (N_14670,N_14298,N_14031);
nand U14671 (N_14671,N_14319,N_14147);
nand U14672 (N_14672,N_14264,N_14150);
nor U14673 (N_14673,N_14276,N_14137);
or U14674 (N_14674,N_14211,N_14241);
and U14675 (N_14675,N_14171,N_14305);
xnor U14676 (N_14676,N_14209,N_14304);
xnor U14677 (N_14677,N_14157,N_14217);
xor U14678 (N_14678,N_14122,N_14268);
xnor U14679 (N_14679,N_14157,N_14289);
or U14680 (N_14680,N_14251,N_14203);
xor U14681 (N_14681,N_14077,N_14286);
or U14682 (N_14682,N_14259,N_14047);
or U14683 (N_14683,N_14372,N_14079);
nand U14684 (N_14684,N_14349,N_14039);
nand U14685 (N_14685,N_14346,N_14298);
and U14686 (N_14686,N_14183,N_14121);
or U14687 (N_14687,N_14290,N_14337);
and U14688 (N_14688,N_14348,N_14182);
or U14689 (N_14689,N_14001,N_14138);
and U14690 (N_14690,N_14206,N_14008);
and U14691 (N_14691,N_14060,N_14067);
xor U14692 (N_14692,N_14101,N_14114);
nor U14693 (N_14693,N_14269,N_14164);
nor U14694 (N_14694,N_14140,N_14346);
nand U14695 (N_14695,N_14173,N_14145);
nor U14696 (N_14696,N_14301,N_14006);
xnor U14697 (N_14697,N_14185,N_14097);
nor U14698 (N_14698,N_14008,N_14193);
and U14699 (N_14699,N_14338,N_14139);
or U14700 (N_14700,N_14360,N_14340);
xor U14701 (N_14701,N_14151,N_14115);
and U14702 (N_14702,N_14074,N_14198);
xor U14703 (N_14703,N_14232,N_14354);
or U14704 (N_14704,N_14138,N_14305);
or U14705 (N_14705,N_14107,N_14334);
xor U14706 (N_14706,N_14181,N_14313);
xor U14707 (N_14707,N_14034,N_14095);
or U14708 (N_14708,N_14126,N_14085);
and U14709 (N_14709,N_14111,N_14319);
xnor U14710 (N_14710,N_14225,N_14381);
or U14711 (N_14711,N_14327,N_14387);
nor U14712 (N_14712,N_14129,N_14140);
nor U14713 (N_14713,N_14386,N_14049);
nand U14714 (N_14714,N_14280,N_14079);
and U14715 (N_14715,N_14277,N_14002);
xnor U14716 (N_14716,N_14211,N_14336);
nand U14717 (N_14717,N_14233,N_14165);
xor U14718 (N_14718,N_14104,N_14107);
or U14719 (N_14719,N_14237,N_14323);
nand U14720 (N_14720,N_14141,N_14358);
xor U14721 (N_14721,N_14107,N_14039);
nand U14722 (N_14722,N_14132,N_14256);
or U14723 (N_14723,N_14257,N_14080);
or U14724 (N_14724,N_14305,N_14367);
or U14725 (N_14725,N_14329,N_14109);
nand U14726 (N_14726,N_14078,N_14040);
nor U14727 (N_14727,N_14139,N_14094);
nand U14728 (N_14728,N_14378,N_14235);
or U14729 (N_14729,N_14399,N_14168);
xor U14730 (N_14730,N_14044,N_14144);
nor U14731 (N_14731,N_14145,N_14147);
and U14732 (N_14732,N_14220,N_14159);
nand U14733 (N_14733,N_14007,N_14175);
xor U14734 (N_14734,N_14391,N_14211);
and U14735 (N_14735,N_14327,N_14112);
and U14736 (N_14736,N_14196,N_14295);
xnor U14737 (N_14737,N_14014,N_14058);
nor U14738 (N_14738,N_14023,N_14251);
or U14739 (N_14739,N_14077,N_14326);
or U14740 (N_14740,N_14056,N_14381);
and U14741 (N_14741,N_14187,N_14157);
or U14742 (N_14742,N_14177,N_14133);
xnor U14743 (N_14743,N_14124,N_14103);
nor U14744 (N_14744,N_14051,N_14338);
nor U14745 (N_14745,N_14141,N_14359);
nand U14746 (N_14746,N_14053,N_14001);
and U14747 (N_14747,N_14183,N_14091);
xnor U14748 (N_14748,N_14368,N_14323);
or U14749 (N_14749,N_14059,N_14152);
nand U14750 (N_14750,N_14276,N_14050);
or U14751 (N_14751,N_14363,N_14006);
xor U14752 (N_14752,N_14194,N_14398);
or U14753 (N_14753,N_14308,N_14075);
xor U14754 (N_14754,N_14170,N_14237);
nand U14755 (N_14755,N_14219,N_14233);
and U14756 (N_14756,N_14079,N_14141);
and U14757 (N_14757,N_14181,N_14159);
nand U14758 (N_14758,N_14233,N_14034);
or U14759 (N_14759,N_14050,N_14261);
nand U14760 (N_14760,N_14341,N_14098);
nand U14761 (N_14761,N_14205,N_14022);
or U14762 (N_14762,N_14101,N_14159);
xnor U14763 (N_14763,N_14060,N_14225);
and U14764 (N_14764,N_14204,N_14388);
or U14765 (N_14765,N_14355,N_14353);
nand U14766 (N_14766,N_14153,N_14337);
and U14767 (N_14767,N_14367,N_14373);
and U14768 (N_14768,N_14319,N_14223);
or U14769 (N_14769,N_14092,N_14347);
nand U14770 (N_14770,N_14056,N_14336);
nand U14771 (N_14771,N_14123,N_14304);
and U14772 (N_14772,N_14338,N_14125);
nor U14773 (N_14773,N_14379,N_14009);
nor U14774 (N_14774,N_14397,N_14258);
xnor U14775 (N_14775,N_14255,N_14344);
nor U14776 (N_14776,N_14366,N_14213);
and U14777 (N_14777,N_14379,N_14294);
nand U14778 (N_14778,N_14067,N_14361);
xor U14779 (N_14779,N_14252,N_14237);
nor U14780 (N_14780,N_14350,N_14203);
nor U14781 (N_14781,N_14386,N_14190);
and U14782 (N_14782,N_14174,N_14089);
xor U14783 (N_14783,N_14272,N_14241);
xnor U14784 (N_14784,N_14097,N_14251);
or U14785 (N_14785,N_14052,N_14359);
xor U14786 (N_14786,N_14228,N_14151);
and U14787 (N_14787,N_14114,N_14058);
or U14788 (N_14788,N_14349,N_14155);
and U14789 (N_14789,N_14070,N_14302);
nor U14790 (N_14790,N_14327,N_14048);
nand U14791 (N_14791,N_14033,N_14064);
nor U14792 (N_14792,N_14016,N_14240);
nor U14793 (N_14793,N_14193,N_14265);
or U14794 (N_14794,N_14319,N_14031);
nor U14795 (N_14795,N_14235,N_14069);
xnor U14796 (N_14796,N_14215,N_14240);
and U14797 (N_14797,N_14226,N_14285);
nand U14798 (N_14798,N_14315,N_14161);
xnor U14799 (N_14799,N_14212,N_14307);
xnor U14800 (N_14800,N_14431,N_14596);
or U14801 (N_14801,N_14436,N_14734);
xnor U14802 (N_14802,N_14665,N_14643);
nor U14803 (N_14803,N_14788,N_14748);
nand U14804 (N_14804,N_14571,N_14453);
or U14805 (N_14805,N_14722,N_14441);
xor U14806 (N_14806,N_14486,N_14529);
and U14807 (N_14807,N_14750,N_14493);
xor U14808 (N_14808,N_14459,N_14662);
xor U14809 (N_14809,N_14651,N_14633);
nor U14810 (N_14810,N_14606,N_14515);
nand U14811 (N_14811,N_14597,N_14672);
nand U14812 (N_14812,N_14409,N_14553);
nor U14813 (N_14813,N_14548,N_14569);
nand U14814 (N_14814,N_14666,N_14730);
nand U14815 (N_14815,N_14659,N_14446);
and U14816 (N_14816,N_14520,N_14504);
or U14817 (N_14817,N_14638,N_14619);
and U14818 (N_14818,N_14702,N_14546);
xnor U14819 (N_14819,N_14600,N_14657);
xor U14820 (N_14820,N_14759,N_14528);
nand U14821 (N_14821,N_14521,N_14550);
or U14822 (N_14822,N_14468,N_14542);
nor U14823 (N_14823,N_14593,N_14795);
or U14824 (N_14824,N_14721,N_14719);
xnor U14825 (N_14825,N_14499,N_14654);
nor U14826 (N_14826,N_14667,N_14652);
or U14827 (N_14827,N_14456,N_14501);
xor U14828 (N_14828,N_14416,N_14492);
and U14829 (N_14829,N_14410,N_14647);
or U14830 (N_14830,N_14437,N_14790);
nor U14831 (N_14831,N_14602,N_14799);
xnor U14832 (N_14832,N_14494,N_14704);
nor U14833 (N_14833,N_14781,N_14589);
nand U14834 (N_14834,N_14474,N_14567);
nor U14835 (N_14835,N_14470,N_14525);
and U14836 (N_14836,N_14412,N_14469);
and U14837 (N_14837,N_14784,N_14541);
and U14838 (N_14838,N_14723,N_14505);
xor U14839 (N_14839,N_14603,N_14562);
nor U14840 (N_14840,N_14590,N_14682);
and U14841 (N_14841,N_14401,N_14439);
and U14842 (N_14842,N_14765,N_14406);
nand U14843 (N_14843,N_14736,N_14689);
or U14844 (N_14844,N_14570,N_14524);
and U14845 (N_14845,N_14735,N_14766);
and U14846 (N_14846,N_14645,N_14423);
nor U14847 (N_14847,N_14457,N_14710);
and U14848 (N_14848,N_14615,N_14552);
nand U14849 (N_14849,N_14400,N_14671);
xnor U14850 (N_14850,N_14407,N_14585);
or U14851 (N_14851,N_14714,N_14644);
nand U14852 (N_14852,N_14577,N_14678);
nand U14853 (N_14853,N_14697,N_14440);
and U14854 (N_14854,N_14793,N_14669);
nor U14855 (N_14855,N_14473,N_14578);
nand U14856 (N_14856,N_14425,N_14729);
or U14857 (N_14857,N_14777,N_14774);
nand U14858 (N_14858,N_14516,N_14428);
and U14859 (N_14859,N_14711,N_14498);
xnor U14860 (N_14860,N_14679,N_14614);
xor U14861 (N_14861,N_14502,N_14771);
or U14862 (N_14862,N_14471,N_14616);
and U14863 (N_14863,N_14716,N_14746);
and U14864 (N_14864,N_14485,N_14594);
nand U14865 (N_14865,N_14772,N_14677);
nand U14866 (N_14866,N_14674,N_14418);
nand U14867 (N_14867,N_14761,N_14581);
nor U14868 (N_14868,N_14426,N_14598);
or U14869 (N_14869,N_14435,N_14449);
or U14870 (N_14870,N_14693,N_14668);
xor U14871 (N_14871,N_14419,N_14708);
nand U14872 (N_14872,N_14465,N_14535);
nor U14873 (N_14873,N_14703,N_14442);
nand U14874 (N_14874,N_14495,N_14731);
xor U14875 (N_14875,N_14797,N_14534);
nand U14876 (N_14876,N_14692,N_14461);
and U14877 (N_14877,N_14532,N_14749);
nor U14878 (N_14878,N_14455,N_14753);
and U14879 (N_14879,N_14497,N_14745);
nand U14880 (N_14880,N_14610,N_14432);
xnor U14881 (N_14881,N_14740,N_14526);
nor U14882 (N_14882,N_14458,N_14760);
nor U14883 (N_14883,N_14509,N_14592);
nand U14884 (N_14884,N_14728,N_14792);
and U14885 (N_14885,N_14663,N_14743);
and U14886 (N_14886,N_14780,N_14568);
or U14887 (N_14887,N_14591,N_14582);
nand U14888 (N_14888,N_14786,N_14434);
nor U14889 (N_14889,N_14725,N_14653);
and U14890 (N_14890,N_14466,N_14408);
or U14891 (N_14891,N_14686,N_14768);
and U14892 (N_14892,N_14483,N_14413);
and U14893 (N_14893,N_14712,N_14506);
or U14894 (N_14894,N_14452,N_14450);
and U14895 (N_14895,N_14429,N_14403);
nand U14896 (N_14896,N_14696,N_14559);
and U14897 (N_14897,N_14579,N_14583);
or U14898 (N_14898,N_14531,N_14460);
nand U14899 (N_14899,N_14462,N_14608);
xor U14900 (N_14900,N_14464,N_14627);
and U14901 (N_14901,N_14572,N_14626);
xnor U14902 (N_14902,N_14764,N_14681);
nor U14903 (N_14903,N_14624,N_14635);
xnor U14904 (N_14904,N_14683,N_14620);
nand U14905 (N_14905,N_14404,N_14554);
xnor U14906 (N_14906,N_14560,N_14574);
nor U14907 (N_14907,N_14604,N_14763);
nand U14908 (N_14908,N_14726,N_14637);
and U14909 (N_14909,N_14747,N_14533);
or U14910 (N_14910,N_14670,N_14451);
xnor U14911 (N_14911,N_14754,N_14630);
and U14912 (N_14912,N_14642,N_14707);
nor U14913 (N_14913,N_14675,N_14555);
or U14914 (N_14914,N_14640,N_14755);
xor U14915 (N_14915,N_14539,N_14540);
and U14916 (N_14916,N_14751,N_14544);
or U14917 (N_14917,N_14724,N_14475);
or U14918 (N_14918,N_14656,N_14618);
xor U14919 (N_14919,N_14566,N_14463);
nand U14920 (N_14920,N_14776,N_14717);
nor U14921 (N_14921,N_14617,N_14639);
nand U14922 (N_14922,N_14530,N_14757);
and U14923 (N_14923,N_14732,N_14573);
or U14924 (N_14924,N_14580,N_14547);
nor U14925 (N_14925,N_14699,N_14785);
xor U14926 (N_14926,N_14587,N_14557);
nor U14927 (N_14927,N_14538,N_14690);
nand U14928 (N_14928,N_14479,N_14609);
xor U14929 (N_14929,N_14796,N_14705);
xnor U14930 (N_14930,N_14537,N_14742);
and U14931 (N_14931,N_14599,N_14477);
nand U14932 (N_14932,N_14522,N_14629);
xor U14933 (N_14933,N_14556,N_14673);
nand U14934 (N_14934,N_14762,N_14482);
nor U14935 (N_14935,N_14733,N_14769);
xnor U14936 (N_14936,N_14625,N_14698);
nor U14937 (N_14937,N_14517,N_14549);
or U14938 (N_14938,N_14467,N_14595);
or U14939 (N_14939,N_14767,N_14632);
nand U14940 (N_14940,N_14576,N_14503);
and U14941 (N_14941,N_14684,N_14448);
nor U14942 (N_14942,N_14514,N_14613);
xnor U14943 (N_14943,N_14621,N_14720);
or U14944 (N_14944,N_14789,N_14676);
and U14945 (N_14945,N_14489,N_14695);
and U14946 (N_14946,N_14472,N_14420);
and U14947 (N_14947,N_14564,N_14634);
nand U14948 (N_14948,N_14508,N_14565);
xnor U14949 (N_14949,N_14427,N_14688);
xor U14950 (N_14950,N_14770,N_14478);
nor U14951 (N_14951,N_14422,N_14445);
nand U14952 (N_14952,N_14417,N_14664);
or U14953 (N_14953,N_14631,N_14636);
or U14954 (N_14954,N_14438,N_14523);
xnor U14955 (N_14955,N_14611,N_14628);
and U14956 (N_14956,N_14490,N_14496);
and U14957 (N_14957,N_14443,N_14519);
and U14958 (N_14958,N_14424,N_14660);
xor U14959 (N_14959,N_14744,N_14480);
nor U14960 (N_14960,N_14447,N_14444);
nand U14961 (N_14961,N_14487,N_14787);
or U14962 (N_14962,N_14563,N_14791);
xnor U14963 (N_14963,N_14700,N_14738);
xor U14964 (N_14964,N_14601,N_14752);
nand U14965 (N_14965,N_14783,N_14649);
nand U14966 (N_14966,N_14561,N_14715);
and U14967 (N_14967,N_14623,N_14512);
nand U14968 (N_14968,N_14476,N_14709);
nor U14969 (N_14969,N_14402,N_14488);
nor U14970 (N_14970,N_14500,N_14646);
or U14971 (N_14971,N_14481,N_14607);
and U14972 (N_14972,N_14491,N_14415);
and U14973 (N_14973,N_14691,N_14513);
nand U14974 (N_14974,N_14782,N_14510);
nand U14975 (N_14975,N_14586,N_14430);
and U14976 (N_14976,N_14718,N_14588);
nand U14977 (N_14977,N_14551,N_14584);
nor U14978 (N_14978,N_14661,N_14741);
nor U14979 (N_14979,N_14641,N_14558);
nor U14980 (N_14980,N_14454,N_14758);
and U14981 (N_14981,N_14687,N_14411);
xor U14982 (N_14982,N_14701,N_14779);
or U14983 (N_14983,N_14605,N_14713);
xnor U14984 (N_14984,N_14706,N_14612);
nand U14985 (N_14985,N_14484,N_14575);
and U14986 (N_14986,N_14518,N_14405);
and U14987 (N_14987,N_14655,N_14737);
and U14988 (N_14988,N_14511,N_14650);
xnor U14989 (N_14989,N_14527,N_14756);
and U14990 (N_14990,N_14798,N_14775);
and U14991 (N_14991,N_14739,N_14658);
xor U14992 (N_14992,N_14545,N_14773);
and U14993 (N_14993,N_14414,N_14433);
or U14994 (N_14994,N_14543,N_14536);
nor U14995 (N_14995,N_14421,N_14622);
nor U14996 (N_14996,N_14794,N_14694);
xnor U14997 (N_14997,N_14685,N_14727);
xor U14998 (N_14998,N_14507,N_14648);
and U14999 (N_14999,N_14680,N_14778);
nor U15000 (N_15000,N_14712,N_14429);
nand U15001 (N_15001,N_14589,N_14736);
nand U15002 (N_15002,N_14736,N_14433);
or U15003 (N_15003,N_14698,N_14679);
and U15004 (N_15004,N_14552,N_14649);
xor U15005 (N_15005,N_14554,N_14753);
or U15006 (N_15006,N_14517,N_14624);
xnor U15007 (N_15007,N_14700,N_14694);
nand U15008 (N_15008,N_14514,N_14667);
or U15009 (N_15009,N_14575,N_14753);
nor U15010 (N_15010,N_14519,N_14701);
nor U15011 (N_15011,N_14557,N_14779);
or U15012 (N_15012,N_14461,N_14608);
nand U15013 (N_15013,N_14718,N_14665);
xnor U15014 (N_15014,N_14516,N_14661);
or U15015 (N_15015,N_14480,N_14607);
nor U15016 (N_15016,N_14778,N_14612);
nand U15017 (N_15017,N_14677,N_14555);
or U15018 (N_15018,N_14489,N_14712);
nor U15019 (N_15019,N_14491,N_14761);
xnor U15020 (N_15020,N_14561,N_14703);
nand U15021 (N_15021,N_14663,N_14446);
or U15022 (N_15022,N_14537,N_14572);
and U15023 (N_15023,N_14511,N_14465);
xnor U15024 (N_15024,N_14664,N_14515);
nor U15025 (N_15025,N_14706,N_14711);
nand U15026 (N_15026,N_14739,N_14556);
or U15027 (N_15027,N_14671,N_14724);
nor U15028 (N_15028,N_14419,N_14771);
or U15029 (N_15029,N_14768,N_14774);
or U15030 (N_15030,N_14527,N_14532);
and U15031 (N_15031,N_14699,N_14761);
nand U15032 (N_15032,N_14536,N_14731);
or U15033 (N_15033,N_14724,N_14613);
or U15034 (N_15034,N_14512,N_14433);
xor U15035 (N_15035,N_14470,N_14403);
and U15036 (N_15036,N_14459,N_14794);
xnor U15037 (N_15037,N_14663,N_14401);
xor U15038 (N_15038,N_14746,N_14500);
xnor U15039 (N_15039,N_14509,N_14588);
xnor U15040 (N_15040,N_14603,N_14400);
xnor U15041 (N_15041,N_14517,N_14557);
xnor U15042 (N_15042,N_14761,N_14653);
and U15043 (N_15043,N_14579,N_14687);
nand U15044 (N_15044,N_14400,N_14415);
nor U15045 (N_15045,N_14597,N_14756);
xor U15046 (N_15046,N_14703,N_14513);
nand U15047 (N_15047,N_14654,N_14453);
xor U15048 (N_15048,N_14783,N_14730);
or U15049 (N_15049,N_14558,N_14672);
and U15050 (N_15050,N_14793,N_14454);
or U15051 (N_15051,N_14567,N_14408);
nor U15052 (N_15052,N_14758,N_14716);
nor U15053 (N_15053,N_14517,N_14459);
nand U15054 (N_15054,N_14476,N_14494);
or U15055 (N_15055,N_14408,N_14750);
xnor U15056 (N_15056,N_14600,N_14636);
xnor U15057 (N_15057,N_14777,N_14444);
and U15058 (N_15058,N_14409,N_14588);
nand U15059 (N_15059,N_14766,N_14403);
xnor U15060 (N_15060,N_14452,N_14456);
nor U15061 (N_15061,N_14456,N_14457);
and U15062 (N_15062,N_14415,N_14734);
or U15063 (N_15063,N_14659,N_14758);
nand U15064 (N_15064,N_14453,N_14710);
nor U15065 (N_15065,N_14654,N_14745);
and U15066 (N_15066,N_14643,N_14605);
nand U15067 (N_15067,N_14412,N_14566);
or U15068 (N_15068,N_14528,N_14739);
and U15069 (N_15069,N_14576,N_14788);
nand U15070 (N_15070,N_14672,N_14418);
nor U15071 (N_15071,N_14690,N_14733);
xnor U15072 (N_15072,N_14571,N_14662);
nor U15073 (N_15073,N_14470,N_14780);
xnor U15074 (N_15074,N_14640,N_14544);
or U15075 (N_15075,N_14405,N_14413);
or U15076 (N_15076,N_14515,N_14653);
xnor U15077 (N_15077,N_14711,N_14620);
nor U15078 (N_15078,N_14407,N_14538);
nand U15079 (N_15079,N_14766,N_14657);
xnor U15080 (N_15080,N_14541,N_14629);
or U15081 (N_15081,N_14703,N_14691);
nor U15082 (N_15082,N_14770,N_14502);
and U15083 (N_15083,N_14447,N_14524);
nor U15084 (N_15084,N_14583,N_14481);
and U15085 (N_15085,N_14687,N_14765);
nor U15086 (N_15086,N_14775,N_14753);
or U15087 (N_15087,N_14699,N_14541);
and U15088 (N_15088,N_14783,N_14765);
and U15089 (N_15089,N_14539,N_14613);
nor U15090 (N_15090,N_14666,N_14437);
nor U15091 (N_15091,N_14681,N_14401);
or U15092 (N_15092,N_14558,N_14415);
nand U15093 (N_15093,N_14797,N_14619);
or U15094 (N_15094,N_14442,N_14663);
or U15095 (N_15095,N_14775,N_14493);
nand U15096 (N_15096,N_14530,N_14456);
or U15097 (N_15097,N_14450,N_14730);
or U15098 (N_15098,N_14769,N_14622);
nand U15099 (N_15099,N_14688,N_14546);
nand U15100 (N_15100,N_14467,N_14783);
and U15101 (N_15101,N_14421,N_14596);
or U15102 (N_15102,N_14557,N_14427);
xnor U15103 (N_15103,N_14789,N_14601);
nand U15104 (N_15104,N_14582,N_14617);
and U15105 (N_15105,N_14726,N_14779);
or U15106 (N_15106,N_14470,N_14420);
nand U15107 (N_15107,N_14592,N_14628);
and U15108 (N_15108,N_14419,N_14558);
nand U15109 (N_15109,N_14421,N_14684);
nor U15110 (N_15110,N_14710,N_14617);
or U15111 (N_15111,N_14498,N_14647);
and U15112 (N_15112,N_14463,N_14644);
xor U15113 (N_15113,N_14414,N_14486);
xnor U15114 (N_15114,N_14783,N_14541);
nand U15115 (N_15115,N_14565,N_14439);
xnor U15116 (N_15116,N_14412,N_14579);
xor U15117 (N_15117,N_14682,N_14418);
and U15118 (N_15118,N_14460,N_14710);
and U15119 (N_15119,N_14513,N_14504);
xor U15120 (N_15120,N_14789,N_14657);
xor U15121 (N_15121,N_14432,N_14408);
xor U15122 (N_15122,N_14447,N_14452);
xor U15123 (N_15123,N_14585,N_14618);
nor U15124 (N_15124,N_14486,N_14767);
nand U15125 (N_15125,N_14554,N_14522);
or U15126 (N_15126,N_14710,N_14745);
and U15127 (N_15127,N_14708,N_14590);
or U15128 (N_15128,N_14650,N_14424);
and U15129 (N_15129,N_14594,N_14691);
and U15130 (N_15130,N_14668,N_14698);
xor U15131 (N_15131,N_14792,N_14466);
nand U15132 (N_15132,N_14788,N_14405);
xor U15133 (N_15133,N_14551,N_14407);
and U15134 (N_15134,N_14699,N_14461);
or U15135 (N_15135,N_14661,N_14447);
or U15136 (N_15136,N_14491,N_14563);
or U15137 (N_15137,N_14646,N_14545);
or U15138 (N_15138,N_14414,N_14496);
xor U15139 (N_15139,N_14439,N_14612);
and U15140 (N_15140,N_14748,N_14601);
or U15141 (N_15141,N_14638,N_14400);
or U15142 (N_15142,N_14553,N_14533);
and U15143 (N_15143,N_14448,N_14788);
xnor U15144 (N_15144,N_14485,N_14592);
or U15145 (N_15145,N_14661,N_14546);
or U15146 (N_15146,N_14694,N_14796);
or U15147 (N_15147,N_14641,N_14595);
and U15148 (N_15148,N_14618,N_14731);
nor U15149 (N_15149,N_14789,N_14474);
xnor U15150 (N_15150,N_14722,N_14600);
nor U15151 (N_15151,N_14587,N_14472);
or U15152 (N_15152,N_14669,N_14584);
and U15153 (N_15153,N_14639,N_14756);
and U15154 (N_15154,N_14615,N_14746);
and U15155 (N_15155,N_14570,N_14527);
or U15156 (N_15156,N_14410,N_14574);
and U15157 (N_15157,N_14458,N_14511);
xor U15158 (N_15158,N_14658,N_14754);
xnor U15159 (N_15159,N_14530,N_14679);
xor U15160 (N_15160,N_14753,N_14494);
and U15161 (N_15161,N_14796,N_14568);
and U15162 (N_15162,N_14681,N_14665);
and U15163 (N_15163,N_14562,N_14758);
and U15164 (N_15164,N_14745,N_14486);
nor U15165 (N_15165,N_14421,N_14489);
and U15166 (N_15166,N_14756,N_14552);
and U15167 (N_15167,N_14403,N_14631);
nand U15168 (N_15168,N_14553,N_14494);
or U15169 (N_15169,N_14737,N_14785);
and U15170 (N_15170,N_14522,N_14483);
and U15171 (N_15171,N_14499,N_14556);
and U15172 (N_15172,N_14757,N_14551);
nand U15173 (N_15173,N_14701,N_14790);
and U15174 (N_15174,N_14542,N_14622);
or U15175 (N_15175,N_14592,N_14519);
nand U15176 (N_15176,N_14769,N_14737);
xnor U15177 (N_15177,N_14406,N_14554);
nor U15178 (N_15178,N_14778,N_14571);
xor U15179 (N_15179,N_14737,N_14746);
nor U15180 (N_15180,N_14413,N_14739);
nor U15181 (N_15181,N_14629,N_14455);
and U15182 (N_15182,N_14687,N_14750);
xor U15183 (N_15183,N_14641,N_14715);
xnor U15184 (N_15184,N_14440,N_14675);
nor U15185 (N_15185,N_14689,N_14682);
nor U15186 (N_15186,N_14776,N_14738);
nor U15187 (N_15187,N_14495,N_14440);
and U15188 (N_15188,N_14555,N_14711);
and U15189 (N_15189,N_14591,N_14605);
nand U15190 (N_15190,N_14437,N_14550);
nor U15191 (N_15191,N_14666,N_14722);
or U15192 (N_15192,N_14434,N_14754);
or U15193 (N_15193,N_14687,N_14563);
and U15194 (N_15194,N_14702,N_14637);
or U15195 (N_15195,N_14622,N_14593);
xnor U15196 (N_15196,N_14445,N_14672);
nand U15197 (N_15197,N_14792,N_14615);
or U15198 (N_15198,N_14614,N_14756);
or U15199 (N_15199,N_14457,N_14601);
and U15200 (N_15200,N_14930,N_14880);
nor U15201 (N_15201,N_15150,N_15080);
nand U15202 (N_15202,N_15087,N_15088);
nor U15203 (N_15203,N_14941,N_15132);
nand U15204 (N_15204,N_15149,N_15076);
and U15205 (N_15205,N_14905,N_14900);
or U15206 (N_15206,N_14846,N_15026);
xor U15207 (N_15207,N_15061,N_15131);
nor U15208 (N_15208,N_15106,N_14994);
nand U15209 (N_15209,N_15077,N_15012);
or U15210 (N_15210,N_14927,N_15144);
or U15211 (N_15211,N_14936,N_14970);
or U15212 (N_15212,N_14887,N_14862);
xnor U15213 (N_15213,N_15184,N_15005);
nand U15214 (N_15214,N_15045,N_14861);
xnor U15215 (N_15215,N_15146,N_15115);
or U15216 (N_15216,N_15127,N_15024);
and U15217 (N_15217,N_15017,N_15032);
nor U15218 (N_15218,N_15122,N_14844);
nand U15219 (N_15219,N_14950,N_14897);
nor U15220 (N_15220,N_15029,N_14892);
and U15221 (N_15221,N_14843,N_15015);
nand U15222 (N_15222,N_14866,N_15105);
nand U15223 (N_15223,N_14976,N_14997);
nor U15224 (N_15224,N_14934,N_15034);
or U15225 (N_15225,N_15137,N_14806);
xnor U15226 (N_15226,N_14845,N_15173);
xor U15227 (N_15227,N_14808,N_15160);
xor U15228 (N_15228,N_15193,N_14912);
or U15229 (N_15229,N_14807,N_15062);
xnor U15230 (N_15230,N_15103,N_14903);
or U15231 (N_15231,N_15179,N_14971);
nor U15232 (N_15232,N_14842,N_15096);
nor U15233 (N_15233,N_14876,N_14972);
and U15234 (N_15234,N_15022,N_14867);
xnor U15235 (N_15235,N_15086,N_14835);
or U15236 (N_15236,N_15028,N_14815);
nand U15237 (N_15237,N_15100,N_14926);
xnor U15238 (N_15238,N_14962,N_15041);
xor U15239 (N_15239,N_14904,N_15143);
nor U15240 (N_15240,N_15008,N_14804);
nor U15241 (N_15241,N_14938,N_14933);
and U15242 (N_15242,N_14919,N_15168);
nand U15243 (N_15243,N_15155,N_15071);
or U15244 (N_15244,N_14918,N_14984);
and U15245 (N_15245,N_15159,N_15133);
or U15246 (N_15246,N_14822,N_15064);
nor U15247 (N_15247,N_15037,N_14947);
or U15248 (N_15248,N_15134,N_15082);
and U15249 (N_15249,N_15060,N_14928);
or U15250 (N_15250,N_14975,N_14886);
xor U15251 (N_15251,N_15136,N_15188);
and U15252 (N_15252,N_15123,N_15180);
nand U15253 (N_15253,N_14883,N_15018);
nand U15254 (N_15254,N_14963,N_15092);
or U15255 (N_15255,N_15172,N_14853);
or U15256 (N_15256,N_15191,N_14959);
nand U15257 (N_15257,N_15070,N_15130);
or U15258 (N_15258,N_15046,N_15072);
and U15259 (N_15259,N_14939,N_15053);
xor U15260 (N_15260,N_15059,N_14952);
nand U15261 (N_15261,N_14906,N_15140);
xor U15262 (N_15262,N_14873,N_15175);
and U15263 (N_15263,N_15181,N_14893);
or U15264 (N_15264,N_15020,N_14878);
and U15265 (N_15265,N_14812,N_15010);
and U15266 (N_15266,N_14908,N_15176);
and U15267 (N_15267,N_14869,N_15167);
xor U15268 (N_15268,N_14855,N_14969);
nor U15269 (N_15269,N_14852,N_15013);
nand U15270 (N_15270,N_14973,N_14982);
and U15271 (N_15271,N_14872,N_15067);
or U15272 (N_15272,N_14818,N_15197);
and U15273 (N_15273,N_15192,N_14850);
nand U15274 (N_15274,N_15027,N_14868);
and U15275 (N_15275,N_15186,N_15019);
or U15276 (N_15276,N_14901,N_15090);
nand U15277 (N_15277,N_15178,N_15110);
or U15278 (N_15278,N_15025,N_15112);
nand U15279 (N_15279,N_14917,N_15114);
and U15280 (N_15280,N_14829,N_15058);
nor U15281 (N_15281,N_14924,N_14837);
or U15282 (N_15282,N_14813,N_14875);
nand U15283 (N_15283,N_15151,N_14942);
nand U15284 (N_15284,N_15121,N_14858);
and U15285 (N_15285,N_14921,N_15126);
nor U15286 (N_15286,N_15003,N_15109);
xor U15287 (N_15287,N_14820,N_15085);
nand U15288 (N_15288,N_14896,N_14957);
nor U15289 (N_15289,N_14965,N_14863);
nor U15290 (N_15290,N_14859,N_15091);
or U15291 (N_15291,N_15057,N_14977);
nand U15292 (N_15292,N_15171,N_15009);
or U15293 (N_15293,N_14956,N_15165);
or U15294 (N_15294,N_14838,N_14978);
or U15295 (N_15295,N_15016,N_15166);
nand U15296 (N_15296,N_14946,N_14967);
xnor U15297 (N_15297,N_15156,N_14920);
xor U15298 (N_15298,N_14981,N_14898);
or U15299 (N_15299,N_14840,N_15000);
xnor U15300 (N_15300,N_15040,N_15030);
and U15301 (N_15301,N_15147,N_15083);
nor U15302 (N_15302,N_15098,N_15031);
xor U15303 (N_15303,N_15095,N_14888);
nor U15304 (N_15304,N_15054,N_15107);
nor U15305 (N_15305,N_14864,N_15039);
or U15306 (N_15306,N_14895,N_15148);
xnor U15307 (N_15307,N_15089,N_14885);
xnor U15308 (N_15308,N_15050,N_15099);
nor U15309 (N_15309,N_14996,N_14841);
nand U15310 (N_15310,N_15048,N_14989);
nor U15311 (N_15311,N_14944,N_15125);
xnor U15312 (N_15312,N_14964,N_15035);
nand U15313 (N_15313,N_14834,N_14800);
nor U15314 (N_15314,N_15093,N_15073);
nand U15315 (N_15315,N_14902,N_15116);
xnor U15316 (N_15316,N_15014,N_15128);
and U15317 (N_15317,N_14839,N_14987);
xnor U15318 (N_15318,N_15047,N_15011);
nor U15319 (N_15319,N_15094,N_14986);
nand U15320 (N_15320,N_14909,N_14980);
and U15321 (N_15321,N_14865,N_15069);
xor U15322 (N_15322,N_14935,N_15141);
nand U15323 (N_15323,N_15036,N_15104);
and U15324 (N_15324,N_15164,N_14802);
xor U15325 (N_15325,N_14954,N_14915);
or U15326 (N_15326,N_14916,N_14999);
and U15327 (N_15327,N_14979,N_14890);
and U15328 (N_15328,N_14810,N_15157);
or U15329 (N_15329,N_15111,N_15033);
and U15330 (N_15330,N_15066,N_14856);
nand U15331 (N_15331,N_14960,N_14826);
nand U15332 (N_15332,N_15161,N_14940);
nand U15333 (N_15333,N_15101,N_14817);
xor U15334 (N_15334,N_15198,N_14913);
nor U15335 (N_15335,N_15084,N_14988);
or U15336 (N_15336,N_14910,N_15145);
xnor U15337 (N_15337,N_15129,N_14948);
or U15338 (N_15338,N_14851,N_14805);
nand U15339 (N_15339,N_15065,N_15118);
nand U15340 (N_15340,N_14823,N_15023);
nor U15341 (N_15341,N_14871,N_15163);
nand U15342 (N_15342,N_15075,N_14955);
and U15343 (N_15343,N_15001,N_14925);
and U15344 (N_15344,N_14811,N_14958);
nor U15345 (N_15345,N_14847,N_14816);
xnor U15346 (N_15346,N_14848,N_14992);
nor U15347 (N_15347,N_14966,N_14821);
or U15348 (N_15348,N_14891,N_14879);
and U15349 (N_15349,N_15056,N_14877);
nand U15350 (N_15350,N_15119,N_15169);
nor U15351 (N_15351,N_15185,N_15042);
xnor U15352 (N_15352,N_14881,N_15044);
or U15353 (N_15353,N_14884,N_15006);
or U15354 (N_15354,N_15097,N_15194);
nand U15355 (N_15355,N_14911,N_14833);
xor U15356 (N_15356,N_14907,N_14828);
xor U15357 (N_15357,N_14899,N_15138);
or U15358 (N_15358,N_15021,N_14801);
nor U15359 (N_15359,N_15182,N_15007);
nand U15360 (N_15360,N_15199,N_14990);
nor U15361 (N_15361,N_14968,N_15051);
and U15362 (N_15362,N_15120,N_14953);
or U15363 (N_15363,N_15142,N_14985);
or U15364 (N_15364,N_14993,N_15124);
nor U15365 (N_15365,N_15195,N_15063);
or U15366 (N_15366,N_15135,N_14974);
nand U15367 (N_15367,N_15049,N_14929);
xor U15368 (N_15368,N_14943,N_15002);
nand U15369 (N_15369,N_14870,N_15079);
xnor U15370 (N_15370,N_15081,N_14857);
xor U15371 (N_15371,N_14937,N_14932);
and U15372 (N_15372,N_14831,N_14827);
nand U15373 (N_15373,N_14951,N_15187);
xnor U15374 (N_15374,N_14991,N_14889);
nor U15375 (N_15375,N_14914,N_15158);
nor U15376 (N_15376,N_14860,N_14832);
nor U15377 (N_15377,N_14849,N_15190);
and U15378 (N_15378,N_15174,N_14882);
nand U15379 (N_15379,N_14949,N_14836);
nor U15380 (N_15380,N_15139,N_15102);
and U15381 (N_15381,N_14961,N_14945);
nor U15382 (N_15382,N_15177,N_15074);
xor U15383 (N_15383,N_14931,N_15043);
nand U15384 (N_15384,N_15153,N_14894);
nand U15385 (N_15385,N_14814,N_14874);
and U15386 (N_15386,N_14809,N_15052);
xnor U15387 (N_15387,N_14983,N_15078);
or U15388 (N_15388,N_15108,N_14923);
and U15389 (N_15389,N_14830,N_15068);
and U15390 (N_15390,N_14825,N_14854);
nand U15391 (N_15391,N_15196,N_15189);
nand U15392 (N_15392,N_14824,N_15113);
xor U15393 (N_15393,N_15038,N_15154);
and U15394 (N_15394,N_15152,N_15170);
or U15395 (N_15395,N_15183,N_14803);
nor U15396 (N_15396,N_14995,N_15055);
nor U15397 (N_15397,N_14819,N_15117);
xor U15398 (N_15398,N_15004,N_14922);
xor U15399 (N_15399,N_14998,N_15162);
or U15400 (N_15400,N_14833,N_14935);
nor U15401 (N_15401,N_15010,N_14985);
nand U15402 (N_15402,N_15009,N_15061);
nor U15403 (N_15403,N_14849,N_14875);
or U15404 (N_15404,N_15154,N_14810);
nand U15405 (N_15405,N_14951,N_14895);
and U15406 (N_15406,N_14991,N_14841);
xor U15407 (N_15407,N_15172,N_14857);
nor U15408 (N_15408,N_15095,N_15071);
xnor U15409 (N_15409,N_14956,N_15027);
xor U15410 (N_15410,N_14988,N_15060);
nand U15411 (N_15411,N_14881,N_14890);
xor U15412 (N_15412,N_14965,N_14981);
and U15413 (N_15413,N_14898,N_15108);
or U15414 (N_15414,N_15047,N_15040);
nor U15415 (N_15415,N_14965,N_15103);
nand U15416 (N_15416,N_15057,N_14883);
nand U15417 (N_15417,N_15026,N_14874);
or U15418 (N_15418,N_15097,N_15136);
or U15419 (N_15419,N_15180,N_15129);
or U15420 (N_15420,N_14946,N_14834);
xnor U15421 (N_15421,N_14819,N_14934);
xnor U15422 (N_15422,N_15067,N_14834);
xor U15423 (N_15423,N_14848,N_14850);
or U15424 (N_15424,N_14871,N_14950);
xnor U15425 (N_15425,N_14931,N_15179);
xnor U15426 (N_15426,N_15089,N_14847);
xor U15427 (N_15427,N_15173,N_15076);
nor U15428 (N_15428,N_15161,N_14812);
xor U15429 (N_15429,N_15169,N_14849);
nand U15430 (N_15430,N_14904,N_15124);
and U15431 (N_15431,N_14899,N_14818);
nand U15432 (N_15432,N_14949,N_15052);
xnor U15433 (N_15433,N_15007,N_15176);
nand U15434 (N_15434,N_14938,N_15029);
xnor U15435 (N_15435,N_15036,N_15086);
nand U15436 (N_15436,N_14882,N_14879);
xor U15437 (N_15437,N_15123,N_15067);
or U15438 (N_15438,N_15042,N_15132);
and U15439 (N_15439,N_15128,N_15074);
nor U15440 (N_15440,N_14920,N_15170);
nand U15441 (N_15441,N_14907,N_14889);
xnor U15442 (N_15442,N_14884,N_15002);
xor U15443 (N_15443,N_15135,N_15157);
nand U15444 (N_15444,N_15057,N_14986);
nor U15445 (N_15445,N_15007,N_15030);
xnor U15446 (N_15446,N_15156,N_14879);
or U15447 (N_15447,N_14945,N_15197);
nor U15448 (N_15448,N_14932,N_15034);
xnor U15449 (N_15449,N_15053,N_15101);
and U15450 (N_15450,N_14897,N_15139);
nor U15451 (N_15451,N_15014,N_15168);
nor U15452 (N_15452,N_15073,N_14976);
nor U15453 (N_15453,N_14829,N_14918);
or U15454 (N_15454,N_14877,N_14834);
and U15455 (N_15455,N_15068,N_15043);
or U15456 (N_15456,N_15126,N_15030);
nand U15457 (N_15457,N_14814,N_15119);
and U15458 (N_15458,N_14911,N_15103);
and U15459 (N_15459,N_15061,N_14909);
or U15460 (N_15460,N_15197,N_15146);
and U15461 (N_15461,N_14879,N_14843);
xnor U15462 (N_15462,N_15036,N_15164);
or U15463 (N_15463,N_15102,N_14985);
and U15464 (N_15464,N_14944,N_14820);
nor U15465 (N_15465,N_14823,N_14870);
xor U15466 (N_15466,N_15095,N_14880);
or U15467 (N_15467,N_15195,N_15078);
or U15468 (N_15468,N_15060,N_14941);
nor U15469 (N_15469,N_15180,N_15116);
nor U15470 (N_15470,N_14800,N_15005);
and U15471 (N_15471,N_14863,N_15189);
nor U15472 (N_15472,N_14902,N_14852);
xor U15473 (N_15473,N_15088,N_14806);
and U15474 (N_15474,N_14998,N_14910);
or U15475 (N_15475,N_14906,N_14826);
xnor U15476 (N_15476,N_14973,N_14881);
or U15477 (N_15477,N_15036,N_15184);
nand U15478 (N_15478,N_14873,N_15035);
nor U15479 (N_15479,N_15062,N_14897);
nand U15480 (N_15480,N_14895,N_14905);
and U15481 (N_15481,N_14954,N_15045);
nor U15482 (N_15482,N_14950,N_15177);
nor U15483 (N_15483,N_14877,N_15168);
or U15484 (N_15484,N_15117,N_14950);
xnor U15485 (N_15485,N_15144,N_14827);
nor U15486 (N_15486,N_14801,N_15020);
or U15487 (N_15487,N_14961,N_15004);
or U15488 (N_15488,N_15076,N_15192);
xor U15489 (N_15489,N_15114,N_14895);
and U15490 (N_15490,N_14806,N_15112);
or U15491 (N_15491,N_14950,N_14936);
xor U15492 (N_15492,N_15079,N_15069);
or U15493 (N_15493,N_15017,N_14908);
and U15494 (N_15494,N_15190,N_14811);
nand U15495 (N_15495,N_14917,N_15064);
nor U15496 (N_15496,N_14807,N_14909);
xnor U15497 (N_15497,N_14916,N_15026);
xnor U15498 (N_15498,N_14968,N_14918);
or U15499 (N_15499,N_15134,N_14822);
xnor U15500 (N_15500,N_14958,N_14852);
nor U15501 (N_15501,N_14941,N_15169);
nand U15502 (N_15502,N_15151,N_14929);
nor U15503 (N_15503,N_15196,N_14807);
nor U15504 (N_15504,N_14803,N_15035);
and U15505 (N_15505,N_14874,N_15039);
or U15506 (N_15506,N_14956,N_15191);
nor U15507 (N_15507,N_15110,N_14941);
xor U15508 (N_15508,N_14933,N_15046);
nor U15509 (N_15509,N_14825,N_14819);
or U15510 (N_15510,N_14805,N_14842);
nor U15511 (N_15511,N_14885,N_15076);
nor U15512 (N_15512,N_15183,N_15163);
nor U15513 (N_15513,N_15106,N_15180);
or U15514 (N_15514,N_14952,N_15138);
nand U15515 (N_15515,N_14993,N_15159);
or U15516 (N_15516,N_14872,N_15129);
and U15517 (N_15517,N_14919,N_14939);
or U15518 (N_15518,N_15103,N_15094);
or U15519 (N_15519,N_15035,N_15137);
and U15520 (N_15520,N_14888,N_15109);
or U15521 (N_15521,N_15159,N_15104);
and U15522 (N_15522,N_14872,N_14855);
nor U15523 (N_15523,N_15130,N_15185);
and U15524 (N_15524,N_14856,N_15164);
nand U15525 (N_15525,N_14978,N_15156);
xnor U15526 (N_15526,N_14932,N_14941);
nand U15527 (N_15527,N_14977,N_15022);
xnor U15528 (N_15528,N_14866,N_15147);
nand U15529 (N_15529,N_14860,N_14949);
nand U15530 (N_15530,N_15193,N_14810);
and U15531 (N_15531,N_14813,N_14848);
nand U15532 (N_15532,N_15038,N_15114);
nand U15533 (N_15533,N_14983,N_15047);
and U15534 (N_15534,N_15129,N_14808);
nor U15535 (N_15535,N_14894,N_14813);
and U15536 (N_15536,N_14970,N_15111);
nand U15537 (N_15537,N_14906,N_15189);
nor U15538 (N_15538,N_15110,N_14943);
and U15539 (N_15539,N_14823,N_14898);
or U15540 (N_15540,N_14809,N_14956);
xnor U15541 (N_15541,N_14956,N_14862);
nor U15542 (N_15542,N_15000,N_15087);
nand U15543 (N_15543,N_15056,N_14932);
or U15544 (N_15544,N_15080,N_15021);
xor U15545 (N_15545,N_14810,N_14832);
or U15546 (N_15546,N_14900,N_15095);
and U15547 (N_15547,N_14821,N_14844);
or U15548 (N_15548,N_15061,N_15097);
xor U15549 (N_15549,N_14965,N_15012);
nor U15550 (N_15550,N_15037,N_14809);
and U15551 (N_15551,N_15021,N_14830);
or U15552 (N_15552,N_14900,N_15159);
xnor U15553 (N_15553,N_14822,N_14823);
and U15554 (N_15554,N_15114,N_15185);
or U15555 (N_15555,N_15071,N_14923);
nand U15556 (N_15556,N_15023,N_14819);
xor U15557 (N_15557,N_15152,N_15038);
and U15558 (N_15558,N_15034,N_15113);
or U15559 (N_15559,N_14970,N_14848);
xnor U15560 (N_15560,N_15145,N_15089);
or U15561 (N_15561,N_14961,N_14983);
and U15562 (N_15562,N_15097,N_15003);
or U15563 (N_15563,N_15094,N_14819);
nand U15564 (N_15564,N_14943,N_15158);
and U15565 (N_15565,N_14866,N_14822);
or U15566 (N_15566,N_14952,N_15117);
and U15567 (N_15567,N_14840,N_14967);
and U15568 (N_15568,N_14883,N_15077);
and U15569 (N_15569,N_14909,N_15179);
xor U15570 (N_15570,N_15036,N_15072);
nand U15571 (N_15571,N_15106,N_15132);
nor U15572 (N_15572,N_14923,N_15174);
nand U15573 (N_15573,N_14869,N_15069);
and U15574 (N_15574,N_14816,N_14830);
and U15575 (N_15575,N_15143,N_14852);
nor U15576 (N_15576,N_14974,N_14805);
xnor U15577 (N_15577,N_15143,N_14850);
and U15578 (N_15578,N_15017,N_15149);
nand U15579 (N_15579,N_14872,N_14819);
and U15580 (N_15580,N_14922,N_14853);
and U15581 (N_15581,N_15140,N_15037);
nor U15582 (N_15582,N_14834,N_15124);
and U15583 (N_15583,N_15149,N_14826);
nand U15584 (N_15584,N_14912,N_14895);
nor U15585 (N_15585,N_14931,N_14805);
nand U15586 (N_15586,N_14864,N_15084);
or U15587 (N_15587,N_14995,N_15091);
or U15588 (N_15588,N_15096,N_14814);
nor U15589 (N_15589,N_15025,N_15129);
or U15590 (N_15590,N_14970,N_15126);
nor U15591 (N_15591,N_14856,N_14948);
nand U15592 (N_15592,N_15129,N_14949);
nor U15593 (N_15593,N_14812,N_14871);
nor U15594 (N_15594,N_15083,N_14833);
and U15595 (N_15595,N_15169,N_15137);
nand U15596 (N_15596,N_15184,N_15046);
xnor U15597 (N_15597,N_14837,N_14969);
or U15598 (N_15598,N_15043,N_15118);
nor U15599 (N_15599,N_14915,N_15195);
nand U15600 (N_15600,N_15496,N_15539);
xnor U15601 (N_15601,N_15305,N_15255);
nor U15602 (N_15602,N_15589,N_15592);
xor U15603 (N_15603,N_15298,N_15245);
nand U15604 (N_15604,N_15431,N_15316);
nand U15605 (N_15605,N_15246,N_15443);
nor U15606 (N_15606,N_15326,N_15216);
and U15607 (N_15607,N_15336,N_15438);
and U15608 (N_15608,N_15429,N_15304);
and U15609 (N_15609,N_15282,N_15537);
xor U15610 (N_15610,N_15457,N_15482);
nand U15611 (N_15611,N_15499,N_15385);
nand U15612 (N_15612,N_15310,N_15467);
nor U15613 (N_15613,N_15296,N_15534);
or U15614 (N_15614,N_15272,N_15535);
and U15615 (N_15615,N_15225,N_15346);
nor U15616 (N_15616,N_15521,N_15553);
nand U15617 (N_15617,N_15538,N_15583);
nor U15618 (N_15618,N_15408,N_15527);
or U15619 (N_15619,N_15354,N_15395);
and U15620 (N_15620,N_15484,N_15261);
nor U15621 (N_15621,N_15280,N_15444);
xor U15622 (N_15622,N_15409,N_15302);
nand U15623 (N_15623,N_15287,N_15450);
xnor U15624 (N_15624,N_15567,N_15413);
and U15625 (N_15625,N_15324,N_15436);
xnor U15626 (N_15626,N_15369,N_15559);
nor U15627 (N_15627,N_15506,N_15543);
xor U15628 (N_15628,N_15295,N_15585);
or U15629 (N_15629,N_15275,N_15208);
nand U15630 (N_15630,N_15425,N_15345);
and U15631 (N_15631,N_15503,N_15265);
or U15632 (N_15632,N_15259,N_15332);
nand U15633 (N_15633,N_15226,N_15476);
xor U15634 (N_15634,N_15516,N_15407);
nand U15635 (N_15635,N_15541,N_15262);
or U15636 (N_15636,N_15487,N_15230);
nor U15637 (N_15637,N_15209,N_15447);
nor U15638 (N_15638,N_15221,N_15594);
nor U15639 (N_15639,N_15264,N_15378);
nor U15640 (N_15640,N_15325,N_15581);
or U15641 (N_15641,N_15480,N_15333);
nor U15642 (N_15642,N_15513,N_15576);
and U15643 (N_15643,N_15432,N_15586);
nand U15644 (N_15644,N_15212,N_15515);
xor U15645 (N_15645,N_15213,N_15475);
nor U15646 (N_15646,N_15353,N_15376);
nor U15647 (N_15647,N_15200,N_15281);
xor U15648 (N_15648,N_15396,N_15462);
nand U15649 (N_15649,N_15224,N_15554);
or U15650 (N_15650,N_15379,N_15218);
and U15651 (N_15651,N_15366,N_15433);
xor U15652 (N_15652,N_15248,N_15341);
nand U15653 (N_15653,N_15373,N_15207);
and U15654 (N_15654,N_15290,N_15397);
or U15655 (N_15655,N_15337,N_15575);
nor U15656 (N_15656,N_15338,N_15365);
nand U15657 (N_15657,N_15321,N_15455);
nand U15658 (N_15658,N_15495,N_15456);
nor U15659 (N_15659,N_15377,N_15240);
nor U15660 (N_15660,N_15524,N_15550);
xnor U15661 (N_15661,N_15520,N_15466);
nor U15662 (N_15662,N_15247,N_15276);
xnor U15663 (N_15663,N_15367,N_15368);
xor U15664 (N_15664,N_15201,N_15279);
and U15665 (N_15665,N_15599,N_15232);
nor U15666 (N_15666,N_15303,N_15266);
nand U15667 (N_15667,N_15215,N_15315);
and U15668 (N_15668,N_15536,N_15414);
nand U15669 (N_15669,N_15299,N_15578);
nor U15670 (N_15670,N_15228,N_15351);
xor U15671 (N_15671,N_15381,N_15465);
xnor U15672 (N_15672,N_15330,N_15239);
and U15673 (N_15673,N_15364,N_15598);
or U15674 (N_15674,N_15517,N_15400);
nor U15675 (N_15675,N_15478,N_15460);
nand U15676 (N_15676,N_15360,N_15229);
or U15677 (N_15677,N_15204,N_15569);
nand U15678 (N_15678,N_15380,N_15522);
and U15679 (N_15679,N_15461,N_15300);
and U15680 (N_15680,N_15568,N_15549);
nand U15681 (N_15681,N_15510,N_15453);
and U15682 (N_15682,N_15406,N_15561);
or U15683 (N_15683,N_15440,N_15439);
and U15684 (N_15684,N_15533,N_15283);
nor U15685 (N_15685,N_15492,N_15386);
nand U15686 (N_15686,N_15356,N_15529);
nand U15687 (N_15687,N_15269,N_15579);
nand U15688 (N_15688,N_15595,N_15422);
xnor U15689 (N_15689,N_15390,N_15254);
or U15690 (N_15690,N_15394,N_15508);
xnor U15691 (N_15691,N_15344,N_15469);
nand U15692 (N_15692,N_15419,N_15382);
and U15693 (N_15693,N_15562,N_15320);
xnor U15694 (N_15694,N_15250,N_15301);
nor U15695 (N_15695,N_15222,N_15235);
nor U15696 (N_15696,N_15306,N_15424);
and U15697 (N_15697,N_15509,N_15588);
nand U15698 (N_15698,N_15311,N_15350);
or U15699 (N_15699,N_15493,N_15464);
and U15700 (N_15700,N_15448,N_15270);
and U15701 (N_15701,N_15342,N_15435);
xnor U15702 (N_15702,N_15548,N_15427);
nor U15703 (N_15703,N_15523,N_15442);
or U15704 (N_15704,N_15375,N_15319);
or U15705 (N_15705,N_15308,N_15387);
and U15706 (N_15706,N_15231,N_15584);
or U15707 (N_15707,N_15219,N_15434);
nor U15708 (N_15708,N_15256,N_15334);
xor U15709 (N_15709,N_15551,N_15577);
nand U15710 (N_15710,N_15339,N_15236);
nor U15711 (N_15711,N_15331,N_15343);
nor U15712 (N_15712,N_15416,N_15347);
or U15713 (N_15713,N_15532,N_15401);
xnor U15714 (N_15714,N_15542,N_15398);
nand U15715 (N_15715,N_15244,N_15260);
and U15716 (N_15716,N_15485,N_15405);
xnor U15717 (N_15717,N_15268,N_15211);
nand U15718 (N_15718,N_15445,N_15558);
nor U15719 (N_15719,N_15285,N_15288);
and U15720 (N_15720,N_15472,N_15504);
xnor U15721 (N_15721,N_15251,N_15459);
and U15722 (N_15722,N_15389,N_15363);
nand U15723 (N_15723,N_15312,N_15267);
or U15724 (N_15724,N_15210,N_15403);
nand U15725 (N_15725,N_15392,N_15596);
and U15726 (N_15726,N_15514,N_15545);
and U15727 (N_15727,N_15289,N_15202);
or U15728 (N_15728,N_15582,N_15307);
nand U15729 (N_15729,N_15399,N_15494);
nor U15730 (N_15730,N_15227,N_15490);
nor U15731 (N_15731,N_15544,N_15286);
or U15732 (N_15732,N_15446,N_15556);
and U15733 (N_15733,N_15359,N_15497);
nor U15734 (N_15734,N_15572,N_15323);
nand U15735 (N_15735,N_15470,N_15355);
nor U15736 (N_15736,N_15217,N_15234);
nand U15737 (N_15737,N_15252,N_15491);
nand U15738 (N_15738,N_15597,N_15546);
or U15739 (N_15739,N_15420,N_15393);
nand U15740 (N_15740,N_15340,N_15486);
or U15741 (N_15741,N_15371,N_15591);
nor U15742 (N_15742,N_15463,N_15291);
nand U15743 (N_15743,N_15511,N_15241);
or U15744 (N_15744,N_15253,N_15277);
xnor U15745 (N_15745,N_15540,N_15348);
nand U15746 (N_15746,N_15278,N_15512);
nor U15747 (N_15747,N_15415,N_15488);
or U15748 (N_15748,N_15417,N_15570);
and U15749 (N_15749,N_15214,N_15498);
or U15750 (N_15750,N_15441,N_15238);
nand U15751 (N_15751,N_15273,N_15587);
xnor U15752 (N_15752,N_15361,N_15526);
xnor U15753 (N_15753,N_15468,N_15309);
and U15754 (N_15754,N_15293,N_15418);
xor U15755 (N_15755,N_15421,N_15284);
xor U15756 (N_15756,N_15458,N_15451);
nor U15757 (N_15757,N_15519,N_15297);
xor U15758 (N_15758,N_15571,N_15370);
or U15759 (N_15759,N_15317,N_15507);
nor U15760 (N_15760,N_15530,N_15328);
or U15761 (N_15761,N_15391,N_15404);
nor U15762 (N_15762,N_15223,N_15590);
or U15763 (N_15763,N_15573,N_15565);
and U15764 (N_15764,N_15489,N_15372);
or U15765 (N_15765,N_15525,N_15258);
nor U15766 (N_15766,N_15313,N_15531);
nor U15767 (N_15767,N_15410,N_15502);
and U15768 (N_15768,N_15203,N_15564);
or U15769 (N_15769,N_15560,N_15449);
xnor U15770 (N_15770,N_15233,N_15552);
or U15771 (N_15771,N_15454,N_15473);
and U15772 (N_15772,N_15477,N_15437);
xor U15773 (N_15773,N_15383,N_15257);
xnor U15774 (N_15774,N_15237,N_15249);
nand U15775 (N_15775,N_15483,N_15481);
or U15776 (N_15776,N_15411,N_15566);
nand U15777 (N_15777,N_15349,N_15555);
and U15778 (N_15778,N_15501,N_15430);
nor U15779 (N_15779,N_15474,N_15593);
nor U15780 (N_15780,N_15352,N_15402);
nor U15781 (N_15781,N_15423,N_15205);
xor U15782 (N_15782,N_15242,N_15358);
xor U15783 (N_15783,N_15518,N_15271);
and U15784 (N_15784,N_15335,N_15505);
nand U15785 (N_15785,N_15479,N_15563);
or U15786 (N_15786,N_15357,N_15318);
xor U15787 (N_15787,N_15452,N_15426);
or U15788 (N_15788,N_15384,N_15206);
nand U15789 (N_15789,N_15322,N_15574);
or U15790 (N_15790,N_15362,N_15388);
or U15791 (N_15791,N_15580,N_15374);
or U15792 (N_15792,N_15428,N_15243);
and U15793 (N_15793,N_15528,N_15327);
nand U15794 (N_15794,N_15220,N_15274);
nand U15795 (N_15795,N_15500,N_15314);
and U15796 (N_15796,N_15471,N_15329);
or U15797 (N_15797,N_15294,N_15263);
nor U15798 (N_15798,N_15292,N_15412);
or U15799 (N_15799,N_15547,N_15557);
and U15800 (N_15800,N_15578,N_15455);
nor U15801 (N_15801,N_15465,N_15338);
or U15802 (N_15802,N_15578,N_15568);
nor U15803 (N_15803,N_15556,N_15304);
nor U15804 (N_15804,N_15387,N_15273);
xor U15805 (N_15805,N_15569,N_15305);
xor U15806 (N_15806,N_15400,N_15301);
or U15807 (N_15807,N_15596,N_15274);
xnor U15808 (N_15808,N_15540,N_15487);
nand U15809 (N_15809,N_15514,N_15230);
nor U15810 (N_15810,N_15242,N_15375);
and U15811 (N_15811,N_15204,N_15510);
nor U15812 (N_15812,N_15380,N_15354);
nand U15813 (N_15813,N_15257,N_15441);
nand U15814 (N_15814,N_15386,N_15502);
nand U15815 (N_15815,N_15538,N_15430);
or U15816 (N_15816,N_15382,N_15242);
xor U15817 (N_15817,N_15428,N_15531);
xnor U15818 (N_15818,N_15341,N_15278);
and U15819 (N_15819,N_15439,N_15323);
or U15820 (N_15820,N_15379,N_15280);
nor U15821 (N_15821,N_15386,N_15451);
nand U15822 (N_15822,N_15583,N_15273);
nor U15823 (N_15823,N_15215,N_15399);
and U15824 (N_15824,N_15269,N_15585);
or U15825 (N_15825,N_15483,N_15549);
and U15826 (N_15826,N_15370,N_15556);
xor U15827 (N_15827,N_15495,N_15293);
or U15828 (N_15828,N_15491,N_15333);
nor U15829 (N_15829,N_15507,N_15347);
or U15830 (N_15830,N_15221,N_15286);
nand U15831 (N_15831,N_15252,N_15463);
xnor U15832 (N_15832,N_15312,N_15392);
nand U15833 (N_15833,N_15204,N_15276);
xor U15834 (N_15834,N_15427,N_15420);
or U15835 (N_15835,N_15307,N_15436);
xnor U15836 (N_15836,N_15351,N_15275);
nor U15837 (N_15837,N_15298,N_15259);
xnor U15838 (N_15838,N_15490,N_15527);
nand U15839 (N_15839,N_15427,N_15514);
xor U15840 (N_15840,N_15431,N_15468);
xor U15841 (N_15841,N_15308,N_15409);
and U15842 (N_15842,N_15225,N_15246);
and U15843 (N_15843,N_15279,N_15342);
and U15844 (N_15844,N_15294,N_15341);
xnor U15845 (N_15845,N_15369,N_15204);
nand U15846 (N_15846,N_15360,N_15472);
nor U15847 (N_15847,N_15282,N_15404);
nand U15848 (N_15848,N_15456,N_15327);
nand U15849 (N_15849,N_15347,N_15571);
or U15850 (N_15850,N_15330,N_15309);
nand U15851 (N_15851,N_15431,N_15599);
nand U15852 (N_15852,N_15573,N_15320);
and U15853 (N_15853,N_15467,N_15270);
nor U15854 (N_15854,N_15294,N_15483);
nor U15855 (N_15855,N_15348,N_15320);
nor U15856 (N_15856,N_15522,N_15535);
nand U15857 (N_15857,N_15408,N_15290);
nor U15858 (N_15858,N_15350,N_15234);
and U15859 (N_15859,N_15373,N_15272);
and U15860 (N_15860,N_15501,N_15462);
and U15861 (N_15861,N_15448,N_15281);
xor U15862 (N_15862,N_15543,N_15314);
xor U15863 (N_15863,N_15294,N_15381);
or U15864 (N_15864,N_15509,N_15515);
nand U15865 (N_15865,N_15586,N_15572);
and U15866 (N_15866,N_15274,N_15387);
nand U15867 (N_15867,N_15238,N_15402);
and U15868 (N_15868,N_15397,N_15482);
nand U15869 (N_15869,N_15494,N_15478);
nor U15870 (N_15870,N_15441,N_15239);
xor U15871 (N_15871,N_15407,N_15356);
xnor U15872 (N_15872,N_15589,N_15445);
and U15873 (N_15873,N_15590,N_15369);
and U15874 (N_15874,N_15327,N_15245);
nand U15875 (N_15875,N_15425,N_15510);
or U15876 (N_15876,N_15294,N_15367);
or U15877 (N_15877,N_15369,N_15261);
or U15878 (N_15878,N_15330,N_15492);
xor U15879 (N_15879,N_15549,N_15206);
xor U15880 (N_15880,N_15332,N_15461);
nand U15881 (N_15881,N_15243,N_15535);
and U15882 (N_15882,N_15494,N_15332);
and U15883 (N_15883,N_15298,N_15466);
or U15884 (N_15884,N_15472,N_15381);
or U15885 (N_15885,N_15240,N_15223);
nand U15886 (N_15886,N_15568,N_15393);
or U15887 (N_15887,N_15392,N_15311);
nor U15888 (N_15888,N_15378,N_15442);
or U15889 (N_15889,N_15469,N_15287);
nor U15890 (N_15890,N_15276,N_15205);
or U15891 (N_15891,N_15534,N_15368);
and U15892 (N_15892,N_15515,N_15379);
nor U15893 (N_15893,N_15503,N_15510);
nand U15894 (N_15894,N_15490,N_15512);
or U15895 (N_15895,N_15253,N_15393);
and U15896 (N_15896,N_15245,N_15346);
or U15897 (N_15897,N_15320,N_15218);
nor U15898 (N_15898,N_15465,N_15440);
xor U15899 (N_15899,N_15292,N_15526);
nand U15900 (N_15900,N_15458,N_15267);
or U15901 (N_15901,N_15594,N_15422);
or U15902 (N_15902,N_15259,N_15283);
or U15903 (N_15903,N_15368,N_15431);
nand U15904 (N_15904,N_15485,N_15372);
nand U15905 (N_15905,N_15395,N_15430);
nor U15906 (N_15906,N_15541,N_15362);
xnor U15907 (N_15907,N_15515,N_15353);
xor U15908 (N_15908,N_15542,N_15501);
xor U15909 (N_15909,N_15578,N_15221);
nor U15910 (N_15910,N_15448,N_15235);
or U15911 (N_15911,N_15537,N_15545);
nand U15912 (N_15912,N_15479,N_15294);
xnor U15913 (N_15913,N_15546,N_15232);
or U15914 (N_15914,N_15526,N_15580);
nand U15915 (N_15915,N_15542,N_15354);
nor U15916 (N_15916,N_15341,N_15363);
and U15917 (N_15917,N_15246,N_15556);
nand U15918 (N_15918,N_15566,N_15569);
nand U15919 (N_15919,N_15432,N_15421);
or U15920 (N_15920,N_15278,N_15413);
or U15921 (N_15921,N_15409,N_15378);
nor U15922 (N_15922,N_15598,N_15539);
nand U15923 (N_15923,N_15274,N_15286);
or U15924 (N_15924,N_15496,N_15422);
and U15925 (N_15925,N_15324,N_15582);
and U15926 (N_15926,N_15573,N_15486);
nand U15927 (N_15927,N_15545,N_15507);
or U15928 (N_15928,N_15478,N_15289);
xnor U15929 (N_15929,N_15300,N_15396);
and U15930 (N_15930,N_15499,N_15512);
or U15931 (N_15931,N_15233,N_15200);
nand U15932 (N_15932,N_15413,N_15541);
nand U15933 (N_15933,N_15248,N_15277);
and U15934 (N_15934,N_15423,N_15502);
nor U15935 (N_15935,N_15309,N_15324);
and U15936 (N_15936,N_15249,N_15325);
or U15937 (N_15937,N_15510,N_15356);
and U15938 (N_15938,N_15256,N_15584);
or U15939 (N_15939,N_15574,N_15212);
nand U15940 (N_15940,N_15322,N_15386);
or U15941 (N_15941,N_15290,N_15379);
and U15942 (N_15942,N_15336,N_15331);
and U15943 (N_15943,N_15598,N_15286);
xnor U15944 (N_15944,N_15570,N_15210);
nor U15945 (N_15945,N_15343,N_15384);
xnor U15946 (N_15946,N_15221,N_15279);
nand U15947 (N_15947,N_15261,N_15343);
or U15948 (N_15948,N_15380,N_15564);
xnor U15949 (N_15949,N_15428,N_15212);
nand U15950 (N_15950,N_15347,N_15220);
nor U15951 (N_15951,N_15392,N_15232);
xor U15952 (N_15952,N_15446,N_15403);
nor U15953 (N_15953,N_15487,N_15427);
nand U15954 (N_15954,N_15455,N_15584);
or U15955 (N_15955,N_15367,N_15520);
nor U15956 (N_15956,N_15438,N_15409);
or U15957 (N_15957,N_15557,N_15591);
nand U15958 (N_15958,N_15580,N_15299);
and U15959 (N_15959,N_15451,N_15519);
and U15960 (N_15960,N_15225,N_15302);
nand U15961 (N_15961,N_15578,N_15465);
xnor U15962 (N_15962,N_15403,N_15348);
and U15963 (N_15963,N_15240,N_15560);
nand U15964 (N_15964,N_15266,N_15319);
nor U15965 (N_15965,N_15293,N_15566);
nand U15966 (N_15966,N_15221,N_15244);
and U15967 (N_15967,N_15518,N_15406);
nor U15968 (N_15968,N_15441,N_15247);
or U15969 (N_15969,N_15423,N_15362);
nand U15970 (N_15970,N_15450,N_15260);
and U15971 (N_15971,N_15504,N_15386);
and U15972 (N_15972,N_15438,N_15461);
nand U15973 (N_15973,N_15243,N_15446);
nor U15974 (N_15974,N_15423,N_15355);
nand U15975 (N_15975,N_15226,N_15251);
and U15976 (N_15976,N_15562,N_15499);
or U15977 (N_15977,N_15552,N_15463);
nand U15978 (N_15978,N_15226,N_15373);
xnor U15979 (N_15979,N_15238,N_15555);
xnor U15980 (N_15980,N_15484,N_15385);
or U15981 (N_15981,N_15273,N_15506);
nand U15982 (N_15982,N_15274,N_15507);
or U15983 (N_15983,N_15318,N_15334);
nand U15984 (N_15984,N_15330,N_15414);
and U15985 (N_15985,N_15246,N_15410);
and U15986 (N_15986,N_15517,N_15330);
nand U15987 (N_15987,N_15445,N_15317);
nand U15988 (N_15988,N_15534,N_15458);
nand U15989 (N_15989,N_15300,N_15230);
and U15990 (N_15990,N_15304,N_15328);
nor U15991 (N_15991,N_15510,N_15490);
nor U15992 (N_15992,N_15256,N_15479);
and U15993 (N_15993,N_15254,N_15231);
nand U15994 (N_15994,N_15586,N_15457);
xor U15995 (N_15995,N_15374,N_15262);
and U15996 (N_15996,N_15366,N_15397);
and U15997 (N_15997,N_15548,N_15206);
and U15998 (N_15998,N_15462,N_15407);
and U15999 (N_15999,N_15204,N_15378);
nor U16000 (N_16000,N_15641,N_15742);
xor U16001 (N_16001,N_15835,N_15834);
or U16002 (N_16002,N_15612,N_15951);
and U16003 (N_16003,N_15729,N_15795);
nand U16004 (N_16004,N_15746,N_15622);
or U16005 (N_16005,N_15791,N_15775);
nand U16006 (N_16006,N_15845,N_15985);
nand U16007 (N_16007,N_15721,N_15956);
nor U16008 (N_16008,N_15656,N_15643);
xor U16009 (N_16009,N_15943,N_15824);
nor U16010 (N_16010,N_15696,N_15973);
and U16011 (N_16011,N_15779,N_15843);
nand U16012 (N_16012,N_15889,N_15933);
nor U16013 (N_16013,N_15821,N_15735);
or U16014 (N_16014,N_15836,N_15832);
or U16015 (N_16015,N_15777,N_15819);
nand U16016 (N_16016,N_15904,N_15755);
and U16017 (N_16017,N_15784,N_15658);
or U16018 (N_16018,N_15668,N_15928);
xor U16019 (N_16019,N_15661,N_15686);
xnor U16020 (N_16020,N_15961,N_15914);
nand U16021 (N_16021,N_15740,N_15760);
nor U16022 (N_16022,N_15960,N_15603);
xor U16023 (N_16023,N_15601,N_15998);
or U16024 (N_16024,N_15693,N_15888);
nand U16025 (N_16025,N_15639,N_15844);
nand U16026 (N_16026,N_15886,N_15830);
or U16027 (N_16027,N_15919,N_15977);
nand U16028 (N_16028,N_15979,N_15811);
nor U16029 (N_16029,N_15850,N_15852);
and U16030 (N_16030,N_15682,N_15714);
and U16031 (N_16031,N_15997,N_15699);
xor U16032 (N_16032,N_15861,N_15781);
and U16033 (N_16033,N_15631,N_15774);
nor U16034 (N_16034,N_15865,N_15866);
nand U16035 (N_16035,N_15780,N_15778);
and U16036 (N_16036,N_15924,N_15932);
nor U16037 (N_16037,N_15651,N_15680);
and U16038 (N_16038,N_15801,N_15992);
and U16039 (N_16039,N_15627,N_15691);
nor U16040 (N_16040,N_15654,N_15615);
and U16041 (N_16041,N_15754,N_15891);
or U16042 (N_16042,N_15665,N_15946);
or U16043 (N_16043,N_15982,N_15797);
xor U16044 (N_16044,N_15640,N_15911);
xnor U16045 (N_16045,N_15805,N_15766);
and U16046 (N_16046,N_15787,N_15848);
and U16047 (N_16047,N_15873,N_15625);
nand U16048 (N_16048,N_15934,N_15923);
xor U16049 (N_16049,N_15783,N_15959);
and U16050 (N_16050,N_15609,N_15829);
nand U16051 (N_16051,N_15744,N_15604);
or U16052 (N_16052,N_15710,N_15814);
or U16053 (N_16053,N_15606,N_15907);
or U16054 (N_16054,N_15720,N_15823);
and U16055 (N_16055,N_15969,N_15681);
nor U16056 (N_16056,N_15994,N_15800);
and U16057 (N_16057,N_15828,N_15980);
xor U16058 (N_16058,N_15990,N_15678);
and U16059 (N_16059,N_15812,N_15872);
nand U16060 (N_16060,N_15770,N_15894);
and U16061 (N_16061,N_15944,N_15790);
xnor U16062 (N_16062,N_15895,N_15776);
nor U16063 (N_16063,N_15751,N_15723);
nor U16064 (N_16064,N_15942,N_15987);
xor U16065 (N_16065,N_15764,N_15859);
or U16066 (N_16066,N_15831,N_15816);
nor U16067 (N_16067,N_15900,N_15773);
xnor U16068 (N_16068,N_15981,N_15975);
xnor U16069 (N_16069,N_15624,N_15820);
nor U16070 (N_16070,N_15673,N_15822);
or U16071 (N_16071,N_15739,N_15728);
and U16072 (N_16072,N_15763,N_15663);
and U16073 (N_16073,N_15683,N_15854);
or U16074 (N_16074,N_15709,N_15613);
or U16075 (N_16075,N_15793,N_15733);
nor U16076 (N_16076,N_15737,N_15918);
and U16077 (N_16077,N_15748,N_15753);
nor U16078 (N_16078,N_15995,N_15926);
or U16079 (N_16079,N_15711,N_15638);
xor U16080 (N_16080,N_15752,N_15750);
or U16081 (N_16081,N_15620,N_15885);
or U16082 (N_16082,N_15772,N_15947);
or U16083 (N_16083,N_15929,N_15853);
nand U16084 (N_16084,N_15867,N_15930);
xnor U16085 (N_16085,N_15749,N_15978);
nand U16086 (N_16086,N_15660,N_15608);
nand U16087 (N_16087,N_15610,N_15782);
or U16088 (N_16088,N_15789,N_15698);
and U16089 (N_16089,N_15803,N_15667);
or U16090 (N_16090,N_15666,N_15771);
xnor U16091 (N_16091,N_15734,N_15689);
or U16092 (N_16092,N_15652,N_15917);
or U16093 (N_16093,N_15840,N_15882);
or U16094 (N_16094,N_15684,N_15838);
nand U16095 (N_16095,N_15738,N_15993);
and U16096 (N_16096,N_15972,N_15692);
nor U16097 (N_16097,N_15921,N_15762);
nor U16098 (N_16098,N_15810,N_15989);
or U16099 (N_16099,N_15675,N_15605);
and U16100 (N_16100,N_15851,N_15788);
nor U16101 (N_16101,N_15644,N_15881);
or U16102 (N_16102,N_15826,N_15635);
or U16103 (N_16103,N_15860,N_15768);
and U16104 (N_16104,N_15717,N_15976);
nor U16105 (N_16105,N_15815,N_15818);
or U16106 (N_16106,N_15621,N_15700);
xnor U16107 (N_16107,N_15949,N_15945);
and U16108 (N_16108,N_15708,N_15971);
and U16109 (N_16109,N_15948,N_15716);
nor U16110 (N_16110,N_15846,N_15707);
or U16111 (N_16111,N_15954,N_15952);
or U16112 (N_16112,N_15988,N_15690);
and U16113 (N_16113,N_15685,N_15999);
xnor U16114 (N_16114,N_15827,N_15722);
nand U16115 (N_16115,N_15653,N_15679);
nor U16116 (N_16116,N_15937,N_15983);
and U16117 (N_16117,N_15953,N_15931);
xor U16118 (N_16118,N_15796,N_15847);
xnor U16119 (N_16119,N_15808,N_15662);
xor U16120 (N_16120,N_15649,N_15804);
and U16121 (N_16121,N_15633,N_15842);
xnor U16122 (N_16122,N_15671,N_15628);
xnor U16123 (N_16123,N_15607,N_15713);
nor U16124 (N_16124,N_15802,N_15758);
or U16125 (N_16125,N_15743,N_15887);
nor U16126 (N_16126,N_15925,N_15871);
or U16127 (N_16127,N_15634,N_15965);
or U16128 (N_16128,N_15912,N_15893);
nand U16129 (N_16129,N_15941,N_15636);
nor U16130 (N_16130,N_15664,N_15726);
nand U16131 (N_16131,N_15984,N_15897);
nor U16132 (N_16132,N_15697,N_15825);
and U16133 (N_16133,N_15786,N_15922);
nor U16134 (N_16134,N_15880,N_15909);
nand U16135 (N_16135,N_15630,N_15940);
nand U16136 (N_16136,N_15855,N_15884);
nor U16137 (N_16137,N_15646,N_15869);
nand U16138 (N_16138,N_15875,N_15837);
xnor U16139 (N_16139,N_15715,N_15807);
or U16140 (N_16140,N_15876,N_15968);
nand U16141 (N_16141,N_15647,N_15903);
nor U16142 (N_16142,N_15955,N_15614);
or U16143 (N_16143,N_15669,N_15920);
nor U16144 (N_16144,N_15712,N_15676);
nand U16145 (N_16145,N_15718,N_15899);
and U16146 (N_16146,N_15727,N_15898);
and U16147 (N_16147,N_15747,N_15618);
or U16148 (N_16148,N_15833,N_15868);
and U16149 (N_16149,N_15839,N_15938);
xor U16150 (N_16150,N_15759,N_15902);
or U16151 (N_16151,N_15706,N_15677);
xor U16152 (N_16152,N_15642,N_15694);
nor U16153 (N_16153,N_15632,N_15874);
xnor U16154 (N_16154,N_15864,N_15725);
nor U16155 (N_16155,N_15986,N_15916);
nor U16156 (N_16156,N_15896,N_15890);
xor U16157 (N_16157,N_15849,N_15927);
and U16158 (N_16158,N_15765,N_15719);
nor U16159 (N_16159,N_15906,N_15957);
or U16160 (N_16160,N_15910,N_15806);
nor U16161 (N_16161,N_15616,N_15602);
nor U16162 (N_16162,N_15936,N_15650);
and U16163 (N_16163,N_15745,N_15674);
nand U16164 (N_16164,N_15905,N_15761);
nand U16165 (N_16165,N_15817,N_15672);
or U16166 (N_16166,N_15915,N_15670);
nand U16167 (N_16167,N_15883,N_15939);
nor U16168 (N_16168,N_15862,N_15648);
nand U16169 (N_16169,N_15870,N_15769);
nor U16170 (N_16170,N_15756,N_15702);
xor U16171 (N_16171,N_15687,N_15974);
xnor U16172 (N_16172,N_15623,N_15813);
nor U16173 (N_16173,N_15705,N_15879);
or U16174 (N_16174,N_15858,N_15703);
xor U16175 (N_16175,N_15863,N_15701);
or U16176 (N_16176,N_15794,N_15963);
xnor U16177 (N_16177,N_15695,N_15856);
and U16178 (N_16178,N_15619,N_15617);
xnor U16179 (N_16179,N_15966,N_15657);
and U16180 (N_16180,N_15913,N_15841);
xnor U16181 (N_16181,N_15799,N_15724);
and U16182 (N_16182,N_15731,N_15600);
nor U16183 (N_16183,N_15704,N_15736);
xnor U16184 (N_16184,N_15785,N_15767);
xnor U16185 (N_16185,N_15991,N_15908);
xor U16186 (N_16186,N_15757,N_15798);
nor U16187 (N_16187,N_15958,N_15892);
nand U16188 (N_16188,N_15996,N_15857);
nand U16189 (N_16189,N_15688,N_15970);
nor U16190 (N_16190,N_15950,N_15935);
xnor U16191 (N_16191,N_15792,N_15637);
nand U16192 (N_16192,N_15901,N_15659);
and U16193 (N_16193,N_15741,N_15877);
nor U16194 (N_16194,N_15629,N_15809);
nand U16195 (N_16195,N_15655,N_15962);
and U16196 (N_16196,N_15964,N_15967);
nand U16197 (N_16197,N_15878,N_15611);
xor U16198 (N_16198,N_15626,N_15732);
and U16199 (N_16199,N_15645,N_15730);
nor U16200 (N_16200,N_15651,N_15656);
and U16201 (N_16201,N_15883,N_15808);
nand U16202 (N_16202,N_15621,N_15615);
or U16203 (N_16203,N_15982,N_15949);
xor U16204 (N_16204,N_15802,N_15881);
and U16205 (N_16205,N_15796,N_15628);
nand U16206 (N_16206,N_15862,N_15604);
or U16207 (N_16207,N_15875,N_15872);
nand U16208 (N_16208,N_15702,N_15620);
xnor U16209 (N_16209,N_15855,N_15828);
or U16210 (N_16210,N_15699,N_15710);
xor U16211 (N_16211,N_15689,N_15783);
nand U16212 (N_16212,N_15816,N_15858);
or U16213 (N_16213,N_15846,N_15762);
nor U16214 (N_16214,N_15630,N_15938);
nand U16215 (N_16215,N_15965,N_15715);
xor U16216 (N_16216,N_15759,N_15864);
nor U16217 (N_16217,N_15781,N_15896);
nand U16218 (N_16218,N_15614,N_15869);
nand U16219 (N_16219,N_15682,N_15787);
nor U16220 (N_16220,N_15720,N_15629);
xnor U16221 (N_16221,N_15913,N_15929);
xnor U16222 (N_16222,N_15710,N_15707);
nand U16223 (N_16223,N_15915,N_15721);
xor U16224 (N_16224,N_15647,N_15892);
and U16225 (N_16225,N_15732,N_15728);
nor U16226 (N_16226,N_15960,N_15901);
and U16227 (N_16227,N_15802,N_15793);
nand U16228 (N_16228,N_15925,N_15870);
or U16229 (N_16229,N_15887,N_15674);
nand U16230 (N_16230,N_15637,N_15936);
and U16231 (N_16231,N_15974,N_15874);
xnor U16232 (N_16232,N_15914,N_15863);
or U16233 (N_16233,N_15946,N_15880);
nand U16234 (N_16234,N_15830,N_15957);
xnor U16235 (N_16235,N_15845,N_15635);
xnor U16236 (N_16236,N_15775,N_15774);
xnor U16237 (N_16237,N_15904,N_15742);
and U16238 (N_16238,N_15679,N_15661);
xor U16239 (N_16239,N_15775,N_15800);
nand U16240 (N_16240,N_15667,N_15908);
xor U16241 (N_16241,N_15819,N_15604);
nand U16242 (N_16242,N_15785,N_15783);
nand U16243 (N_16243,N_15906,N_15900);
nand U16244 (N_16244,N_15754,N_15823);
nor U16245 (N_16245,N_15750,N_15782);
xor U16246 (N_16246,N_15903,N_15608);
and U16247 (N_16247,N_15733,N_15803);
or U16248 (N_16248,N_15719,N_15944);
xnor U16249 (N_16249,N_15888,N_15993);
xor U16250 (N_16250,N_15933,N_15834);
xnor U16251 (N_16251,N_15910,N_15970);
or U16252 (N_16252,N_15838,N_15914);
nor U16253 (N_16253,N_15864,N_15742);
nand U16254 (N_16254,N_15620,N_15978);
xor U16255 (N_16255,N_15637,N_15913);
nor U16256 (N_16256,N_15956,N_15920);
and U16257 (N_16257,N_15722,N_15681);
or U16258 (N_16258,N_15735,N_15672);
and U16259 (N_16259,N_15763,N_15671);
xnor U16260 (N_16260,N_15926,N_15909);
nor U16261 (N_16261,N_15822,N_15856);
and U16262 (N_16262,N_15709,N_15733);
and U16263 (N_16263,N_15975,N_15758);
xor U16264 (N_16264,N_15640,N_15620);
xor U16265 (N_16265,N_15991,N_15791);
and U16266 (N_16266,N_15943,N_15896);
nand U16267 (N_16267,N_15737,N_15619);
and U16268 (N_16268,N_15914,N_15619);
and U16269 (N_16269,N_15850,N_15800);
nand U16270 (N_16270,N_15994,N_15822);
and U16271 (N_16271,N_15816,N_15811);
and U16272 (N_16272,N_15666,N_15854);
nand U16273 (N_16273,N_15990,N_15728);
and U16274 (N_16274,N_15973,N_15975);
nor U16275 (N_16275,N_15772,N_15939);
and U16276 (N_16276,N_15866,N_15975);
nor U16277 (N_16277,N_15899,N_15846);
and U16278 (N_16278,N_15639,N_15735);
nor U16279 (N_16279,N_15925,N_15740);
nor U16280 (N_16280,N_15830,N_15811);
nand U16281 (N_16281,N_15921,N_15806);
nand U16282 (N_16282,N_15873,N_15699);
nand U16283 (N_16283,N_15605,N_15878);
or U16284 (N_16284,N_15829,N_15775);
or U16285 (N_16285,N_15811,N_15841);
nand U16286 (N_16286,N_15937,N_15767);
or U16287 (N_16287,N_15909,N_15933);
or U16288 (N_16288,N_15614,N_15668);
or U16289 (N_16289,N_15767,N_15932);
and U16290 (N_16290,N_15761,N_15857);
and U16291 (N_16291,N_15677,N_15827);
or U16292 (N_16292,N_15943,N_15630);
or U16293 (N_16293,N_15831,N_15829);
nor U16294 (N_16294,N_15880,N_15860);
or U16295 (N_16295,N_15884,N_15838);
or U16296 (N_16296,N_15885,N_15986);
or U16297 (N_16297,N_15600,N_15818);
nand U16298 (N_16298,N_15988,N_15919);
or U16299 (N_16299,N_15916,N_15774);
nor U16300 (N_16300,N_15773,N_15610);
nor U16301 (N_16301,N_15974,N_15745);
nor U16302 (N_16302,N_15947,N_15997);
and U16303 (N_16303,N_15783,N_15843);
and U16304 (N_16304,N_15621,N_15772);
or U16305 (N_16305,N_15992,N_15908);
or U16306 (N_16306,N_15902,N_15610);
xor U16307 (N_16307,N_15787,N_15856);
nor U16308 (N_16308,N_15968,N_15996);
xor U16309 (N_16309,N_15908,N_15661);
nor U16310 (N_16310,N_15875,N_15600);
nand U16311 (N_16311,N_15632,N_15762);
or U16312 (N_16312,N_15743,N_15937);
or U16313 (N_16313,N_15652,N_15859);
nor U16314 (N_16314,N_15937,N_15608);
and U16315 (N_16315,N_15906,N_15620);
or U16316 (N_16316,N_15919,N_15889);
nand U16317 (N_16317,N_15759,N_15919);
nand U16318 (N_16318,N_15927,N_15772);
and U16319 (N_16319,N_15913,N_15704);
nor U16320 (N_16320,N_15899,N_15978);
nand U16321 (N_16321,N_15847,N_15818);
or U16322 (N_16322,N_15723,N_15754);
nor U16323 (N_16323,N_15934,N_15869);
nand U16324 (N_16324,N_15737,N_15889);
or U16325 (N_16325,N_15896,N_15937);
nor U16326 (N_16326,N_15867,N_15616);
nor U16327 (N_16327,N_15741,N_15672);
nor U16328 (N_16328,N_15970,N_15994);
or U16329 (N_16329,N_15814,N_15877);
xor U16330 (N_16330,N_15641,N_15686);
nand U16331 (N_16331,N_15907,N_15654);
and U16332 (N_16332,N_15969,N_15837);
nand U16333 (N_16333,N_15918,N_15683);
or U16334 (N_16334,N_15892,N_15751);
xor U16335 (N_16335,N_15913,N_15769);
xnor U16336 (N_16336,N_15626,N_15980);
or U16337 (N_16337,N_15841,N_15654);
nand U16338 (N_16338,N_15895,N_15976);
nand U16339 (N_16339,N_15917,N_15927);
or U16340 (N_16340,N_15631,N_15862);
nor U16341 (N_16341,N_15785,N_15831);
or U16342 (N_16342,N_15897,N_15963);
and U16343 (N_16343,N_15763,N_15810);
nand U16344 (N_16344,N_15733,N_15906);
or U16345 (N_16345,N_15839,N_15741);
nor U16346 (N_16346,N_15940,N_15625);
or U16347 (N_16347,N_15923,N_15957);
and U16348 (N_16348,N_15635,N_15792);
and U16349 (N_16349,N_15618,N_15679);
or U16350 (N_16350,N_15835,N_15803);
or U16351 (N_16351,N_15676,N_15892);
and U16352 (N_16352,N_15921,N_15891);
xnor U16353 (N_16353,N_15985,N_15667);
or U16354 (N_16354,N_15835,N_15762);
and U16355 (N_16355,N_15796,N_15977);
xor U16356 (N_16356,N_15798,N_15895);
nand U16357 (N_16357,N_15757,N_15638);
nand U16358 (N_16358,N_15900,N_15676);
nand U16359 (N_16359,N_15968,N_15808);
nand U16360 (N_16360,N_15703,N_15693);
nand U16361 (N_16361,N_15683,N_15649);
or U16362 (N_16362,N_15712,N_15904);
xor U16363 (N_16363,N_15802,N_15725);
or U16364 (N_16364,N_15980,N_15814);
nor U16365 (N_16365,N_15762,N_15987);
or U16366 (N_16366,N_15923,N_15940);
nor U16367 (N_16367,N_15695,N_15696);
nand U16368 (N_16368,N_15935,N_15979);
xor U16369 (N_16369,N_15901,N_15955);
or U16370 (N_16370,N_15943,N_15737);
nor U16371 (N_16371,N_15703,N_15733);
xor U16372 (N_16372,N_15715,N_15907);
nor U16373 (N_16373,N_15880,N_15763);
nor U16374 (N_16374,N_15643,N_15979);
nand U16375 (N_16375,N_15677,N_15912);
xor U16376 (N_16376,N_15890,N_15786);
nand U16377 (N_16377,N_15821,N_15859);
nor U16378 (N_16378,N_15980,N_15886);
nor U16379 (N_16379,N_15798,N_15802);
and U16380 (N_16380,N_15728,N_15889);
or U16381 (N_16381,N_15675,N_15869);
or U16382 (N_16382,N_15788,N_15767);
nand U16383 (N_16383,N_15622,N_15621);
nor U16384 (N_16384,N_15777,N_15642);
nand U16385 (N_16385,N_15855,N_15995);
xor U16386 (N_16386,N_15765,N_15953);
xor U16387 (N_16387,N_15607,N_15743);
xor U16388 (N_16388,N_15688,N_15620);
nand U16389 (N_16389,N_15632,N_15610);
nand U16390 (N_16390,N_15841,N_15744);
xnor U16391 (N_16391,N_15861,N_15770);
and U16392 (N_16392,N_15821,N_15709);
nor U16393 (N_16393,N_15656,N_15833);
or U16394 (N_16394,N_15938,N_15767);
nor U16395 (N_16395,N_15676,N_15894);
nor U16396 (N_16396,N_15677,N_15721);
nand U16397 (N_16397,N_15699,N_15787);
xor U16398 (N_16398,N_15993,N_15938);
and U16399 (N_16399,N_15840,N_15635);
and U16400 (N_16400,N_16275,N_16379);
and U16401 (N_16401,N_16328,N_16239);
xnor U16402 (N_16402,N_16125,N_16087);
or U16403 (N_16403,N_16250,N_16258);
nand U16404 (N_16404,N_16214,N_16143);
or U16405 (N_16405,N_16383,N_16118);
nor U16406 (N_16406,N_16339,N_16005);
xor U16407 (N_16407,N_16131,N_16164);
or U16408 (N_16408,N_16015,N_16206);
xor U16409 (N_16409,N_16191,N_16303);
xnor U16410 (N_16410,N_16331,N_16014);
nand U16411 (N_16411,N_16182,N_16170);
nor U16412 (N_16412,N_16376,N_16268);
and U16413 (N_16413,N_16196,N_16247);
or U16414 (N_16414,N_16262,N_16381);
nor U16415 (N_16415,N_16129,N_16309);
or U16416 (N_16416,N_16066,N_16204);
xnor U16417 (N_16417,N_16366,N_16117);
or U16418 (N_16418,N_16220,N_16388);
nor U16419 (N_16419,N_16148,N_16045);
nand U16420 (N_16420,N_16107,N_16340);
and U16421 (N_16421,N_16279,N_16332);
nand U16422 (N_16422,N_16166,N_16302);
nand U16423 (N_16423,N_16189,N_16396);
or U16424 (N_16424,N_16380,N_16197);
xor U16425 (N_16425,N_16307,N_16075);
xor U16426 (N_16426,N_16171,N_16245);
nor U16427 (N_16427,N_16174,N_16217);
and U16428 (N_16428,N_16119,N_16313);
nand U16429 (N_16429,N_16329,N_16176);
and U16430 (N_16430,N_16116,N_16321);
nand U16431 (N_16431,N_16318,N_16024);
xor U16432 (N_16432,N_16076,N_16081);
xnor U16433 (N_16433,N_16195,N_16147);
and U16434 (N_16434,N_16157,N_16311);
nand U16435 (N_16435,N_16265,N_16298);
nand U16436 (N_16436,N_16221,N_16351);
xor U16437 (N_16437,N_16084,N_16008);
xor U16438 (N_16438,N_16280,N_16226);
xnor U16439 (N_16439,N_16062,N_16139);
and U16440 (N_16440,N_16378,N_16273);
nor U16441 (N_16441,N_16326,N_16151);
nor U16442 (N_16442,N_16223,N_16295);
nand U16443 (N_16443,N_16061,N_16229);
or U16444 (N_16444,N_16057,N_16193);
and U16445 (N_16445,N_16306,N_16278);
nor U16446 (N_16446,N_16259,N_16106);
nand U16447 (N_16447,N_16361,N_16249);
nand U16448 (N_16448,N_16054,N_16232);
nand U16449 (N_16449,N_16113,N_16070);
nor U16450 (N_16450,N_16104,N_16183);
nor U16451 (N_16451,N_16260,N_16333);
and U16452 (N_16452,N_16053,N_16165);
or U16453 (N_16453,N_16101,N_16392);
or U16454 (N_16454,N_16093,N_16293);
nor U16455 (N_16455,N_16023,N_16068);
nand U16456 (N_16456,N_16094,N_16072);
or U16457 (N_16457,N_16325,N_16327);
or U16458 (N_16458,N_16255,N_16112);
and U16459 (N_16459,N_16345,N_16224);
nand U16460 (N_16460,N_16297,N_16025);
or U16461 (N_16461,N_16200,N_16288);
xor U16462 (N_16462,N_16059,N_16031);
nand U16463 (N_16463,N_16092,N_16021);
or U16464 (N_16464,N_16338,N_16291);
xor U16465 (N_16465,N_16294,N_16287);
nor U16466 (N_16466,N_16160,N_16363);
nand U16467 (N_16467,N_16150,N_16362);
nand U16468 (N_16468,N_16185,N_16141);
and U16469 (N_16469,N_16169,N_16199);
or U16470 (N_16470,N_16190,N_16036);
and U16471 (N_16471,N_16099,N_16124);
nor U16472 (N_16472,N_16144,N_16091);
nand U16473 (N_16473,N_16198,N_16349);
and U16474 (N_16474,N_16315,N_16242);
xnor U16475 (N_16475,N_16034,N_16310);
xor U16476 (N_16476,N_16370,N_16252);
nor U16477 (N_16477,N_16052,N_16347);
or U16478 (N_16478,N_16060,N_16234);
or U16479 (N_16479,N_16020,N_16108);
xor U16480 (N_16480,N_16028,N_16277);
xor U16481 (N_16481,N_16312,N_16127);
and U16482 (N_16482,N_16161,N_16138);
nor U16483 (N_16483,N_16359,N_16071);
nor U16484 (N_16484,N_16386,N_16030);
xor U16485 (N_16485,N_16213,N_16394);
and U16486 (N_16486,N_16358,N_16056);
and U16487 (N_16487,N_16123,N_16022);
nand U16488 (N_16488,N_16369,N_16033);
xnor U16489 (N_16489,N_16097,N_16238);
xor U16490 (N_16490,N_16391,N_16159);
xor U16491 (N_16491,N_16050,N_16371);
xor U16492 (N_16492,N_16355,N_16142);
or U16493 (N_16493,N_16122,N_16109);
xnor U16494 (N_16494,N_16393,N_16373);
and U16495 (N_16495,N_16317,N_16181);
and U16496 (N_16496,N_16257,N_16114);
and U16497 (N_16497,N_16001,N_16336);
and U16498 (N_16498,N_16248,N_16105);
xor U16499 (N_16499,N_16365,N_16137);
and U16500 (N_16500,N_16067,N_16018);
or U16501 (N_16501,N_16368,N_16322);
nor U16502 (N_16502,N_16314,N_16051);
nor U16503 (N_16503,N_16046,N_16212);
or U16504 (N_16504,N_16389,N_16134);
nand U16505 (N_16505,N_16003,N_16284);
nand U16506 (N_16506,N_16384,N_16342);
nand U16507 (N_16507,N_16017,N_16374);
nor U16508 (N_16508,N_16341,N_16039);
nand U16509 (N_16509,N_16065,N_16089);
or U16510 (N_16510,N_16375,N_16283);
or U16511 (N_16511,N_16103,N_16296);
nor U16512 (N_16512,N_16304,N_16230);
and U16513 (N_16513,N_16344,N_16095);
or U16514 (N_16514,N_16064,N_16222);
xnor U16515 (N_16515,N_16156,N_16299);
and U16516 (N_16516,N_16082,N_16290);
xor U16517 (N_16517,N_16135,N_16043);
nor U16518 (N_16518,N_16038,N_16184);
nor U16519 (N_16519,N_16074,N_16251);
nand U16520 (N_16520,N_16019,N_16289);
or U16521 (N_16521,N_16350,N_16180);
or U16522 (N_16522,N_16011,N_16240);
or U16523 (N_16523,N_16016,N_16348);
nor U16524 (N_16524,N_16382,N_16080);
nand U16525 (N_16525,N_16264,N_16208);
or U16526 (N_16526,N_16175,N_16167);
xor U16527 (N_16527,N_16237,N_16177);
or U16528 (N_16528,N_16246,N_16115);
nand U16529 (N_16529,N_16120,N_16187);
nand U16530 (N_16530,N_16155,N_16002);
nor U16531 (N_16531,N_16110,N_16292);
xnor U16532 (N_16532,N_16352,N_16320);
or U16533 (N_16533,N_16211,N_16272);
and U16534 (N_16534,N_16395,N_16337);
nand U16535 (N_16535,N_16281,N_16090);
nand U16536 (N_16536,N_16048,N_16269);
and U16537 (N_16537,N_16244,N_16286);
and U16538 (N_16538,N_16098,N_16077);
or U16539 (N_16539,N_16044,N_16276);
xor U16540 (N_16540,N_16004,N_16227);
and U16541 (N_16541,N_16192,N_16356);
nand U16542 (N_16542,N_16367,N_16063);
xor U16543 (N_16543,N_16319,N_16168);
and U16544 (N_16544,N_16387,N_16083);
and U16545 (N_16545,N_16216,N_16377);
nor U16546 (N_16546,N_16146,N_16069);
and U16547 (N_16547,N_16241,N_16390);
or U16548 (N_16548,N_16163,N_16149);
nor U16549 (N_16549,N_16305,N_16042);
xnor U16550 (N_16550,N_16007,N_16398);
and U16551 (N_16551,N_16308,N_16145);
nor U16552 (N_16552,N_16256,N_16372);
xor U16553 (N_16553,N_16225,N_16055);
nand U16554 (N_16554,N_16158,N_16133);
xor U16555 (N_16555,N_16330,N_16153);
and U16556 (N_16556,N_16049,N_16334);
or U16557 (N_16557,N_16209,N_16357);
and U16558 (N_16558,N_16041,N_16354);
and U16559 (N_16559,N_16270,N_16009);
or U16560 (N_16560,N_16316,N_16086);
xnor U16561 (N_16561,N_16032,N_16010);
and U16562 (N_16562,N_16035,N_16397);
and U16563 (N_16563,N_16207,N_16254);
nor U16564 (N_16564,N_16323,N_16186);
and U16565 (N_16565,N_16324,N_16100);
xor U16566 (N_16566,N_16088,N_16364);
nor U16567 (N_16567,N_16228,N_16140);
nand U16568 (N_16568,N_16274,N_16037);
nor U16569 (N_16569,N_16029,N_16013);
nand U16570 (N_16570,N_16271,N_16136);
nor U16571 (N_16571,N_16231,N_16203);
nor U16572 (N_16572,N_16235,N_16202);
xor U16573 (N_16573,N_16210,N_16128);
nand U16574 (N_16574,N_16027,N_16085);
and U16575 (N_16575,N_16194,N_16126);
xor U16576 (N_16576,N_16353,N_16243);
nand U16577 (N_16577,N_16219,N_16006);
or U16578 (N_16578,N_16178,N_16179);
nor U16579 (N_16579,N_16253,N_16040);
xor U16580 (N_16580,N_16152,N_16012);
xor U16581 (N_16581,N_16058,N_16385);
or U16582 (N_16582,N_16162,N_16267);
xnor U16583 (N_16583,N_16188,N_16399);
xnor U16584 (N_16584,N_16173,N_16073);
nand U16585 (N_16585,N_16079,N_16102);
or U16586 (N_16586,N_16201,N_16026);
or U16587 (N_16587,N_16111,N_16078);
xor U16588 (N_16588,N_16282,N_16000);
xor U16589 (N_16589,N_16121,N_16130);
nor U16590 (N_16590,N_16263,N_16132);
and U16591 (N_16591,N_16346,N_16300);
xnor U16592 (N_16592,N_16285,N_16233);
nand U16593 (N_16593,N_16205,N_16301);
xor U16594 (N_16594,N_16172,N_16266);
nand U16595 (N_16595,N_16343,N_16215);
or U16596 (N_16596,N_16154,N_16047);
nor U16597 (N_16597,N_16360,N_16218);
xor U16598 (N_16598,N_16236,N_16261);
or U16599 (N_16599,N_16096,N_16335);
and U16600 (N_16600,N_16233,N_16248);
and U16601 (N_16601,N_16395,N_16130);
xor U16602 (N_16602,N_16097,N_16117);
nor U16603 (N_16603,N_16350,N_16140);
or U16604 (N_16604,N_16286,N_16298);
nor U16605 (N_16605,N_16274,N_16322);
xnor U16606 (N_16606,N_16162,N_16080);
nor U16607 (N_16607,N_16250,N_16127);
xor U16608 (N_16608,N_16271,N_16097);
and U16609 (N_16609,N_16182,N_16343);
xnor U16610 (N_16610,N_16233,N_16219);
or U16611 (N_16611,N_16080,N_16282);
xnor U16612 (N_16612,N_16317,N_16143);
nand U16613 (N_16613,N_16075,N_16110);
xnor U16614 (N_16614,N_16243,N_16010);
or U16615 (N_16615,N_16109,N_16040);
and U16616 (N_16616,N_16210,N_16200);
nor U16617 (N_16617,N_16180,N_16211);
or U16618 (N_16618,N_16329,N_16261);
and U16619 (N_16619,N_16264,N_16029);
or U16620 (N_16620,N_16095,N_16148);
and U16621 (N_16621,N_16097,N_16308);
and U16622 (N_16622,N_16295,N_16010);
and U16623 (N_16623,N_16193,N_16048);
xor U16624 (N_16624,N_16073,N_16293);
xnor U16625 (N_16625,N_16014,N_16023);
and U16626 (N_16626,N_16087,N_16226);
nand U16627 (N_16627,N_16392,N_16179);
nor U16628 (N_16628,N_16063,N_16345);
or U16629 (N_16629,N_16231,N_16020);
xnor U16630 (N_16630,N_16119,N_16263);
and U16631 (N_16631,N_16191,N_16026);
xnor U16632 (N_16632,N_16297,N_16305);
and U16633 (N_16633,N_16179,N_16089);
and U16634 (N_16634,N_16034,N_16050);
and U16635 (N_16635,N_16134,N_16210);
nor U16636 (N_16636,N_16049,N_16389);
and U16637 (N_16637,N_16224,N_16367);
nor U16638 (N_16638,N_16303,N_16112);
and U16639 (N_16639,N_16182,N_16269);
and U16640 (N_16640,N_16219,N_16159);
xor U16641 (N_16641,N_16233,N_16003);
and U16642 (N_16642,N_16367,N_16061);
or U16643 (N_16643,N_16150,N_16221);
nor U16644 (N_16644,N_16014,N_16361);
nand U16645 (N_16645,N_16170,N_16338);
xnor U16646 (N_16646,N_16342,N_16306);
and U16647 (N_16647,N_16229,N_16068);
and U16648 (N_16648,N_16165,N_16303);
and U16649 (N_16649,N_16149,N_16304);
nor U16650 (N_16650,N_16129,N_16059);
xnor U16651 (N_16651,N_16075,N_16271);
xor U16652 (N_16652,N_16183,N_16145);
nor U16653 (N_16653,N_16186,N_16170);
xor U16654 (N_16654,N_16392,N_16095);
nand U16655 (N_16655,N_16329,N_16205);
xor U16656 (N_16656,N_16389,N_16088);
nand U16657 (N_16657,N_16126,N_16376);
nor U16658 (N_16658,N_16081,N_16064);
nor U16659 (N_16659,N_16282,N_16068);
xor U16660 (N_16660,N_16368,N_16389);
nand U16661 (N_16661,N_16196,N_16076);
nand U16662 (N_16662,N_16210,N_16354);
and U16663 (N_16663,N_16175,N_16363);
or U16664 (N_16664,N_16251,N_16158);
and U16665 (N_16665,N_16066,N_16237);
xnor U16666 (N_16666,N_16160,N_16070);
and U16667 (N_16667,N_16298,N_16091);
and U16668 (N_16668,N_16257,N_16134);
or U16669 (N_16669,N_16125,N_16024);
nand U16670 (N_16670,N_16360,N_16073);
nor U16671 (N_16671,N_16064,N_16385);
xnor U16672 (N_16672,N_16154,N_16057);
nand U16673 (N_16673,N_16134,N_16159);
nor U16674 (N_16674,N_16105,N_16389);
nand U16675 (N_16675,N_16371,N_16299);
or U16676 (N_16676,N_16264,N_16117);
and U16677 (N_16677,N_16163,N_16198);
xnor U16678 (N_16678,N_16240,N_16257);
and U16679 (N_16679,N_16320,N_16161);
nand U16680 (N_16680,N_16380,N_16134);
xnor U16681 (N_16681,N_16374,N_16224);
xnor U16682 (N_16682,N_16017,N_16128);
nand U16683 (N_16683,N_16070,N_16049);
or U16684 (N_16684,N_16278,N_16105);
nor U16685 (N_16685,N_16219,N_16347);
nand U16686 (N_16686,N_16121,N_16261);
nor U16687 (N_16687,N_16187,N_16314);
nand U16688 (N_16688,N_16059,N_16212);
and U16689 (N_16689,N_16155,N_16337);
or U16690 (N_16690,N_16365,N_16394);
and U16691 (N_16691,N_16139,N_16164);
and U16692 (N_16692,N_16387,N_16010);
nand U16693 (N_16693,N_16066,N_16063);
nand U16694 (N_16694,N_16219,N_16077);
nor U16695 (N_16695,N_16060,N_16151);
and U16696 (N_16696,N_16200,N_16053);
or U16697 (N_16697,N_16209,N_16036);
and U16698 (N_16698,N_16163,N_16154);
and U16699 (N_16699,N_16155,N_16275);
or U16700 (N_16700,N_16166,N_16153);
xor U16701 (N_16701,N_16203,N_16124);
xor U16702 (N_16702,N_16111,N_16346);
or U16703 (N_16703,N_16320,N_16315);
nand U16704 (N_16704,N_16267,N_16251);
xor U16705 (N_16705,N_16352,N_16147);
nand U16706 (N_16706,N_16222,N_16066);
nand U16707 (N_16707,N_16138,N_16103);
xor U16708 (N_16708,N_16395,N_16128);
nor U16709 (N_16709,N_16384,N_16307);
or U16710 (N_16710,N_16110,N_16230);
and U16711 (N_16711,N_16193,N_16066);
xor U16712 (N_16712,N_16313,N_16352);
or U16713 (N_16713,N_16005,N_16368);
xor U16714 (N_16714,N_16118,N_16041);
and U16715 (N_16715,N_16297,N_16291);
and U16716 (N_16716,N_16183,N_16146);
nand U16717 (N_16717,N_16298,N_16231);
nand U16718 (N_16718,N_16351,N_16313);
or U16719 (N_16719,N_16125,N_16382);
and U16720 (N_16720,N_16277,N_16303);
nand U16721 (N_16721,N_16051,N_16383);
xor U16722 (N_16722,N_16250,N_16337);
or U16723 (N_16723,N_16379,N_16396);
or U16724 (N_16724,N_16324,N_16302);
or U16725 (N_16725,N_16083,N_16332);
or U16726 (N_16726,N_16006,N_16393);
nand U16727 (N_16727,N_16387,N_16373);
or U16728 (N_16728,N_16117,N_16188);
nor U16729 (N_16729,N_16173,N_16124);
or U16730 (N_16730,N_16011,N_16342);
and U16731 (N_16731,N_16263,N_16204);
and U16732 (N_16732,N_16097,N_16346);
xnor U16733 (N_16733,N_16055,N_16296);
nor U16734 (N_16734,N_16355,N_16001);
or U16735 (N_16735,N_16020,N_16211);
or U16736 (N_16736,N_16277,N_16077);
nand U16737 (N_16737,N_16293,N_16113);
or U16738 (N_16738,N_16124,N_16382);
nor U16739 (N_16739,N_16277,N_16049);
or U16740 (N_16740,N_16367,N_16054);
xnor U16741 (N_16741,N_16396,N_16039);
and U16742 (N_16742,N_16272,N_16138);
xnor U16743 (N_16743,N_16120,N_16102);
xnor U16744 (N_16744,N_16053,N_16034);
xor U16745 (N_16745,N_16025,N_16039);
nand U16746 (N_16746,N_16280,N_16248);
or U16747 (N_16747,N_16329,N_16376);
and U16748 (N_16748,N_16396,N_16027);
xnor U16749 (N_16749,N_16289,N_16122);
nand U16750 (N_16750,N_16306,N_16254);
nand U16751 (N_16751,N_16052,N_16026);
and U16752 (N_16752,N_16312,N_16281);
nand U16753 (N_16753,N_16200,N_16250);
nor U16754 (N_16754,N_16172,N_16014);
xor U16755 (N_16755,N_16002,N_16371);
nor U16756 (N_16756,N_16297,N_16347);
xnor U16757 (N_16757,N_16112,N_16249);
nor U16758 (N_16758,N_16365,N_16115);
and U16759 (N_16759,N_16016,N_16225);
xnor U16760 (N_16760,N_16366,N_16230);
or U16761 (N_16761,N_16034,N_16147);
nand U16762 (N_16762,N_16016,N_16182);
xnor U16763 (N_16763,N_16328,N_16306);
xor U16764 (N_16764,N_16383,N_16251);
nand U16765 (N_16765,N_16386,N_16103);
or U16766 (N_16766,N_16076,N_16209);
nor U16767 (N_16767,N_16023,N_16197);
or U16768 (N_16768,N_16301,N_16254);
nor U16769 (N_16769,N_16093,N_16274);
and U16770 (N_16770,N_16096,N_16020);
nand U16771 (N_16771,N_16104,N_16207);
or U16772 (N_16772,N_16227,N_16373);
or U16773 (N_16773,N_16269,N_16119);
or U16774 (N_16774,N_16072,N_16053);
and U16775 (N_16775,N_16013,N_16078);
and U16776 (N_16776,N_16074,N_16281);
xnor U16777 (N_16777,N_16163,N_16247);
xnor U16778 (N_16778,N_16014,N_16314);
nor U16779 (N_16779,N_16083,N_16134);
or U16780 (N_16780,N_16389,N_16226);
xnor U16781 (N_16781,N_16147,N_16190);
nor U16782 (N_16782,N_16210,N_16086);
nor U16783 (N_16783,N_16279,N_16114);
nand U16784 (N_16784,N_16185,N_16304);
nor U16785 (N_16785,N_16313,N_16058);
or U16786 (N_16786,N_16037,N_16031);
nand U16787 (N_16787,N_16197,N_16314);
and U16788 (N_16788,N_16357,N_16025);
or U16789 (N_16789,N_16127,N_16159);
nor U16790 (N_16790,N_16019,N_16147);
nor U16791 (N_16791,N_16270,N_16127);
xor U16792 (N_16792,N_16198,N_16111);
and U16793 (N_16793,N_16318,N_16361);
or U16794 (N_16794,N_16021,N_16089);
and U16795 (N_16795,N_16158,N_16043);
xnor U16796 (N_16796,N_16324,N_16222);
or U16797 (N_16797,N_16002,N_16085);
nand U16798 (N_16798,N_16281,N_16393);
nand U16799 (N_16799,N_16042,N_16111);
or U16800 (N_16800,N_16655,N_16621);
nand U16801 (N_16801,N_16403,N_16753);
nor U16802 (N_16802,N_16523,N_16515);
and U16803 (N_16803,N_16718,N_16686);
xnor U16804 (N_16804,N_16464,N_16486);
or U16805 (N_16805,N_16483,N_16541);
or U16806 (N_16806,N_16462,N_16591);
or U16807 (N_16807,N_16592,N_16522);
and U16808 (N_16808,N_16411,N_16578);
nor U16809 (N_16809,N_16780,N_16642);
and U16810 (N_16810,N_16645,N_16704);
nand U16811 (N_16811,N_16683,N_16404);
nand U16812 (N_16812,N_16558,N_16764);
and U16813 (N_16813,N_16465,N_16456);
xnor U16814 (N_16814,N_16530,N_16689);
nor U16815 (N_16815,N_16536,N_16401);
nor U16816 (N_16816,N_16739,N_16710);
nand U16817 (N_16817,N_16428,N_16663);
nor U16818 (N_16818,N_16490,N_16613);
and U16819 (N_16819,N_16502,N_16409);
or U16820 (N_16820,N_16793,N_16791);
nor U16821 (N_16821,N_16737,N_16677);
and U16822 (N_16822,N_16609,N_16550);
and U16823 (N_16823,N_16773,N_16416);
and U16824 (N_16824,N_16487,N_16499);
and U16825 (N_16825,N_16583,N_16664);
xor U16826 (N_16826,N_16461,N_16412);
xnor U16827 (N_16827,N_16444,N_16797);
or U16828 (N_16828,N_16784,N_16746);
nand U16829 (N_16829,N_16770,N_16496);
or U16830 (N_16830,N_16440,N_16652);
nand U16831 (N_16831,N_16457,N_16567);
nor U16832 (N_16832,N_16501,N_16633);
nor U16833 (N_16833,N_16666,N_16426);
xnor U16834 (N_16834,N_16561,N_16738);
xor U16835 (N_16835,N_16529,N_16714);
nor U16836 (N_16836,N_16629,N_16580);
and U16837 (N_16837,N_16625,N_16607);
nor U16838 (N_16838,N_16482,N_16604);
or U16839 (N_16839,N_16754,N_16507);
or U16840 (N_16840,N_16598,N_16495);
and U16841 (N_16841,N_16460,N_16623);
or U16842 (N_16842,N_16468,N_16463);
nor U16843 (N_16843,N_16469,N_16509);
nand U16844 (N_16844,N_16493,N_16698);
xor U16845 (N_16845,N_16672,N_16762);
nand U16846 (N_16846,N_16640,N_16631);
or U16847 (N_16847,N_16721,N_16521);
nor U16848 (N_16848,N_16707,N_16685);
xor U16849 (N_16849,N_16741,N_16505);
nor U16850 (N_16850,N_16615,N_16566);
or U16851 (N_16851,N_16436,N_16681);
xor U16852 (N_16852,N_16451,N_16545);
xor U16853 (N_16853,N_16750,N_16555);
xor U16854 (N_16854,N_16573,N_16595);
and U16855 (N_16855,N_16790,N_16571);
xor U16856 (N_16856,N_16405,N_16605);
nand U16857 (N_16857,N_16705,N_16455);
or U16858 (N_16858,N_16572,N_16442);
nor U16859 (N_16859,N_16799,N_16568);
xnor U16860 (N_16860,N_16745,N_16727);
and U16861 (N_16861,N_16528,N_16674);
and U16862 (N_16862,N_16726,N_16648);
nor U16863 (N_16863,N_16516,N_16679);
nor U16864 (N_16864,N_16637,N_16650);
or U16865 (N_16865,N_16636,N_16749);
xor U16866 (N_16866,N_16448,N_16435);
xor U16867 (N_16867,N_16671,N_16611);
or U16868 (N_16868,N_16701,N_16743);
and U16869 (N_16869,N_16688,N_16508);
xor U16870 (N_16870,N_16434,N_16747);
or U16871 (N_16871,N_16706,N_16406);
nor U16872 (N_16872,N_16540,N_16447);
or U16873 (N_16873,N_16775,N_16470);
and U16874 (N_16874,N_16531,N_16582);
nand U16875 (N_16875,N_16788,N_16560);
nor U16876 (N_16876,N_16777,N_16699);
nor U16877 (N_16877,N_16789,N_16513);
nand U16878 (N_16878,N_16692,N_16641);
and U16879 (N_16879,N_16662,N_16657);
or U16880 (N_16880,N_16602,N_16771);
nand U16881 (N_16881,N_16562,N_16458);
and U16882 (N_16882,N_16415,N_16511);
xor U16883 (N_16883,N_16712,N_16731);
nor U16884 (N_16884,N_16723,N_16450);
and U16885 (N_16885,N_16472,N_16553);
nor U16886 (N_16886,N_16425,N_16594);
and U16887 (N_16887,N_16787,N_16722);
nor U16888 (N_16888,N_16433,N_16713);
nand U16889 (N_16889,N_16684,N_16599);
xor U16890 (N_16890,N_16510,N_16763);
nor U16891 (N_16891,N_16579,N_16556);
nand U16892 (N_16892,N_16772,N_16413);
nor U16893 (N_16893,N_16638,N_16612);
nor U16894 (N_16894,N_16708,N_16497);
xor U16895 (N_16895,N_16660,N_16766);
or U16896 (N_16896,N_16441,N_16622);
and U16897 (N_16897,N_16628,N_16418);
or U16898 (N_16898,N_16479,N_16608);
xor U16899 (N_16899,N_16740,N_16673);
and U16900 (N_16900,N_16539,N_16634);
xnor U16901 (N_16901,N_16627,N_16700);
xor U16902 (N_16902,N_16644,N_16734);
and U16903 (N_16903,N_16702,N_16659);
and U16904 (N_16904,N_16500,N_16724);
or U16905 (N_16905,N_16581,N_16577);
or U16906 (N_16906,N_16669,N_16676);
or U16907 (N_16907,N_16732,N_16410);
or U16908 (N_16908,N_16619,N_16761);
nand U16909 (N_16909,N_16620,N_16488);
xor U16910 (N_16910,N_16554,N_16533);
and U16911 (N_16911,N_16653,N_16446);
xnor U16912 (N_16912,N_16779,N_16400);
nand U16913 (N_16913,N_16768,N_16757);
nor U16914 (N_16914,N_16570,N_16736);
xnor U16915 (N_16915,N_16711,N_16494);
xor U16916 (N_16916,N_16574,N_16796);
and U16917 (N_16917,N_16564,N_16670);
xor U16918 (N_16918,N_16559,N_16667);
or U16919 (N_16919,N_16693,N_16774);
xnor U16920 (N_16920,N_16569,N_16597);
xnor U16921 (N_16921,N_16534,N_16514);
nor U16922 (N_16922,N_16475,N_16551);
nor U16923 (N_16923,N_16719,N_16614);
nand U16924 (N_16924,N_16481,N_16618);
xnor U16925 (N_16925,N_16437,N_16624);
nand U16926 (N_16926,N_16525,N_16626);
xor U16927 (N_16927,N_16651,N_16695);
xnor U16928 (N_16928,N_16744,N_16675);
nor U16929 (N_16929,N_16584,N_16431);
and U16930 (N_16930,N_16476,N_16492);
xnor U16931 (N_16931,N_16538,N_16765);
nand U16932 (N_16932,N_16544,N_16548);
and U16933 (N_16933,N_16678,N_16785);
or U16934 (N_16934,N_16647,N_16422);
nor U16935 (N_16935,N_16680,N_16429);
or U16936 (N_16936,N_16546,N_16643);
nand U16937 (N_16937,N_16424,N_16616);
nand U16938 (N_16938,N_16658,N_16438);
nand U16939 (N_16939,N_16601,N_16782);
nor U16940 (N_16940,N_16617,N_16795);
xnor U16941 (N_16941,N_16519,N_16503);
and U16942 (N_16942,N_16439,N_16535);
xnor U16943 (N_16943,N_16668,N_16557);
nor U16944 (N_16944,N_16407,N_16474);
or U16945 (N_16945,N_16600,N_16547);
or U16946 (N_16946,N_16419,N_16445);
nand U16947 (N_16947,N_16512,N_16691);
nand U16948 (N_16948,N_16414,N_16717);
or U16949 (N_16949,N_16697,N_16466);
nand U16950 (N_16950,N_16593,N_16646);
xor U16951 (N_16951,N_16752,N_16665);
nor U16952 (N_16952,N_16575,N_16526);
nor U16953 (N_16953,N_16524,N_16781);
nor U16954 (N_16954,N_16729,N_16755);
and U16955 (N_16955,N_16798,N_16506);
nor U16956 (N_16956,N_16527,N_16402);
nand U16957 (N_16957,N_16543,N_16480);
nand U16958 (N_16958,N_16532,N_16491);
or U16959 (N_16959,N_16730,N_16751);
or U16960 (N_16960,N_16408,N_16517);
and U16961 (N_16961,N_16709,N_16537);
nand U16962 (N_16962,N_16715,N_16759);
and U16963 (N_16963,N_16735,N_16610);
xnor U16964 (N_16964,N_16587,N_16453);
xnor U16965 (N_16965,N_16760,N_16661);
or U16966 (N_16966,N_16767,N_16725);
nand U16967 (N_16967,N_16748,N_16682);
nor U16968 (N_16968,N_16769,N_16504);
xnor U16969 (N_16969,N_16432,N_16518);
nand U16970 (N_16970,N_16485,N_16471);
or U16971 (N_16971,N_16452,N_16417);
nor U16972 (N_16972,N_16489,N_16783);
xor U16973 (N_16973,N_16549,N_16716);
and U16974 (N_16974,N_16454,N_16459);
nor U16975 (N_16975,N_16588,N_16478);
xor U16976 (N_16976,N_16443,N_16477);
nor U16977 (N_16977,N_16728,N_16654);
and U16978 (N_16978,N_16687,N_16576);
and U16979 (N_16979,N_16484,N_16656);
and U16980 (N_16980,N_16585,N_16703);
and U16981 (N_16981,N_16590,N_16520);
nor U16982 (N_16982,N_16786,N_16649);
or U16983 (N_16983,N_16498,N_16603);
xnor U16984 (N_16984,N_16776,N_16635);
or U16985 (N_16985,N_16589,N_16420);
nand U16986 (N_16986,N_16720,N_16421);
nand U16987 (N_16987,N_16794,N_16696);
or U16988 (N_16988,N_16733,N_16563);
or U16989 (N_16989,N_16427,N_16742);
and U16990 (N_16990,N_16586,N_16552);
and U16991 (N_16991,N_16756,N_16690);
nand U16992 (N_16992,N_16792,N_16596);
xor U16993 (N_16993,N_16758,N_16430);
nand U16994 (N_16994,N_16542,N_16694);
nor U16995 (N_16995,N_16473,N_16778);
nor U16996 (N_16996,N_16449,N_16606);
or U16997 (N_16997,N_16630,N_16639);
xnor U16998 (N_16998,N_16565,N_16632);
or U16999 (N_16999,N_16467,N_16423);
nor U17000 (N_17000,N_16636,N_16656);
xnor U17001 (N_17001,N_16702,N_16705);
nand U17002 (N_17002,N_16664,N_16416);
xnor U17003 (N_17003,N_16687,N_16561);
nor U17004 (N_17004,N_16737,N_16435);
and U17005 (N_17005,N_16604,N_16446);
nor U17006 (N_17006,N_16405,N_16642);
and U17007 (N_17007,N_16562,N_16599);
nand U17008 (N_17008,N_16463,N_16597);
nor U17009 (N_17009,N_16473,N_16599);
or U17010 (N_17010,N_16753,N_16659);
and U17011 (N_17011,N_16680,N_16442);
and U17012 (N_17012,N_16781,N_16439);
nand U17013 (N_17013,N_16553,N_16639);
or U17014 (N_17014,N_16574,N_16572);
or U17015 (N_17015,N_16759,N_16518);
or U17016 (N_17016,N_16479,N_16448);
xnor U17017 (N_17017,N_16689,N_16475);
xor U17018 (N_17018,N_16607,N_16437);
or U17019 (N_17019,N_16452,N_16610);
nor U17020 (N_17020,N_16660,N_16728);
or U17021 (N_17021,N_16537,N_16470);
or U17022 (N_17022,N_16674,N_16641);
nor U17023 (N_17023,N_16684,N_16607);
and U17024 (N_17024,N_16514,N_16574);
xnor U17025 (N_17025,N_16563,N_16656);
and U17026 (N_17026,N_16423,N_16553);
nand U17027 (N_17027,N_16442,N_16752);
xor U17028 (N_17028,N_16742,N_16468);
nand U17029 (N_17029,N_16468,N_16734);
nand U17030 (N_17030,N_16405,N_16789);
and U17031 (N_17031,N_16776,N_16563);
xor U17032 (N_17032,N_16760,N_16683);
xor U17033 (N_17033,N_16528,N_16468);
and U17034 (N_17034,N_16718,N_16501);
xor U17035 (N_17035,N_16470,N_16651);
nor U17036 (N_17036,N_16465,N_16541);
nor U17037 (N_17037,N_16469,N_16576);
nand U17038 (N_17038,N_16501,N_16620);
nand U17039 (N_17039,N_16485,N_16715);
nand U17040 (N_17040,N_16713,N_16464);
and U17041 (N_17041,N_16426,N_16429);
nor U17042 (N_17042,N_16554,N_16537);
or U17043 (N_17043,N_16607,N_16468);
or U17044 (N_17044,N_16419,N_16469);
or U17045 (N_17045,N_16788,N_16411);
nand U17046 (N_17046,N_16779,N_16759);
or U17047 (N_17047,N_16779,N_16587);
or U17048 (N_17048,N_16631,N_16454);
or U17049 (N_17049,N_16787,N_16784);
nor U17050 (N_17050,N_16525,N_16630);
nor U17051 (N_17051,N_16678,N_16733);
or U17052 (N_17052,N_16527,N_16492);
nand U17053 (N_17053,N_16645,N_16695);
or U17054 (N_17054,N_16617,N_16522);
nor U17055 (N_17055,N_16665,N_16722);
or U17056 (N_17056,N_16763,N_16408);
and U17057 (N_17057,N_16770,N_16447);
nand U17058 (N_17058,N_16681,N_16618);
nor U17059 (N_17059,N_16430,N_16629);
nand U17060 (N_17060,N_16628,N_16588);
or U17061 (N_17061,N_16441,N_16598);
nor U17062 (N_17062,N_16561,N_16679);
and U17063 (N_17063,N_16578,N_16463);
nor U17064 (N_17064,N_16564,N_16774);
nand U17065 (N_17065,N_16656,N_16439);
nor U17066 (N_17066,N_16418,N_16493);
nand U17067 (N_17067,N_16537,N_16762);
and U17068 (N_17068,N_16655,N_16521);
and U17069 (N_17069,N_16675,N_16571);
nor U17070 (N_17070,N_16644,N_16795);
xor U17071 (N_17071,N_16770,N_16578);
nand U17072 (N_17072,N_16424,N_16618);
nand U17073 (N_17073,N_16759,N_16490);
xnor U17074 (N_17074,N_16487,N_16414);
nand U17075 (N_17075,N_16740,N_16543);
and U17076 (N_17076,N_16581,N_16724);
xor U17077 (N_17077,N_16780,N_16647);
nand U17078 (N_17078,N_16551,N_16732);
nor U17079 (N_17079,N_16618,N_16666);
and U17080 (N_17080,N_16795,N_16775);
nor U17081 (N_17081,N_16625,N_16470);
nor U17082 (N_17082,N_16530,N_16601);
nand U17083 (N_17083,N_16605,N_16569);
xnor U17084 (N_17084,N_16534,N_16783);
nor U17085 (N_17085,N_16606,N_16754);
or U17086 (N_17086,N_16605,N_16591);
nor U17087 (N_17087,N_16602,N_16556);
or U17088 (N_17088,N_16748,N_16619);
xor U17089 (N_17089,N_16582,N_16469);
nor U17090 (N_17090,N_16431,N_16461);
and U17091 (N_17091,N_16580,N_16583);
and U17092 (N_17092,N_16741,N_16409);
nor U17093 (N_17093,N_16615,N_16599);
nand U17094 (N_17094,N_16454,N_16614);
nor U17095 (N_17095,N_16478,N_16492);
and U17096 (N_17096,N_16416,N_16452);
or U17097 (N_17097,N_16747,N_16706);
nor U17098 (N_17098,N_16748,N_16405);
nor U17099 (N_17099,N_16509,N_16492);
or U17100 (N_17100,N_16592,N_16723);
xnor U17101 (N_17101,N_16777,N_16731);
and U17102 (N_17102,N_16446,N_16640);
and U17103 (N_17103,N_16719,N_16641);
xnor U17104 (N_17104,N_16469,N_16568);
or U17105 (N_17105,N_16694,N_16494);
xor U17106 (N_17106,N_16572,N_16509);
or U17107 (N_17107,N_16523,N_16665);
xnor U17108 (N_17108,N_16670,N_16459);
or U17109 (N_17109,N_16753,N_16638);
and U17110 (N_17110,N_16751,N_16475);
nand U17111 (N_17111,N_16767,N_16667);
xnor U17112 (N_17112,N_16742,N_16690);
or U17113 (N_17113,N_16545,N_16655);
and U17114 (N_17114,N_16702,N_16430);
nand U17115 (N_17115,N_16705,N_16487);
and U17116 (N_17116,N_16605,N_16604);
or U17117 (N_17117,N_16756,N_16559);
nor U17118 (N_17118,N_16780,N_16722);
nand U17119 (N_17119,N_16784,N_16619);
or U17120 (N_17120,N_16484,N_16716);
and U17121 (N_17121,N_16490,N_16637);
nor U17122 (N_17122,N_16557,N_16762);
and U17123 (N_17123,N_16613,N_16716);
xnor U17124 (N_17124,N_16487,N_16583);
or U17125 (N_17125,N_16650,N_16706);
nand U17126 (N_17126,N_16550,N_16736);
nand U17127 (N_17127,N_16487,N_16452);
and U17128 (N_17128,N_16782,N_16420);
nand U17129 (N_17129,N_16560,N_16786);
xor U17130 (N_17130,N_16536,N_16676);
xnor U17131 (N_17131,N_16730,N_16472);
xor U17132 (N_17132,N_16759,N_16559);
or U17133 (N_17133,N_16588,N_16415);
nor U17134 (N_17134,N_16794,N_16507);
or U17135 (N_17135,N_16557,N_16409);
or U17136 (N_17136,N_16439,N_16583);
xnor U17137 (N_17137,N_16770,N_16592);
or U17138 (N_17138,N_16640,N_16441);
and U17139 (N_17139,N_16471,N_16620);
and U17140 (N_17140,N_16644,N_16613);
xor U17141 (N_17141,N_16764,N_16659);
nor U17142 (N_17142,N_16527,N_16534);
nand U17143 (N_17143,N_16404,N_16694);
xor U17144 (N_17144,N_16586,N_16786);
nand U17145 (N_17145,N_16730,N_16480);
and U17146 (N_17146,N_16652,N_16678);
nand U17147 (N_17147,N_16487,N_16453);
nor U17148 (N_17148,N_16754,N_16716);
and U17149 (N_17149,N_16474,N_16452);
and U17150 (N_17150,N_16400,N_16754);
and U17151 (N_17151,N_16605,N_16685);
nand U17152 (N_17152,N_16700,N_16438);
or U17153 (N_17153,N_16682,N_16594);
nor U17154 (N_17154,N_16596,N_16675);
or U17155 (N_17155,N_16761,N_16763);
xor U17156 (N_17156,N_16774,N_16730);
nor U17157 (N_17157,N_16488,N_16646);
or U17158 (N_17158,N_16440,N_16579);
nand U17159 (N_17159,N_16423,N_16759);
nand U17160 (N_17160,N_16773,N_16503);
xnor U17161 (N_17161,N_16715,N_16654);
or U17162 (N_17162,N_16456,N_16742);
or U17163 (N_17163,N_16631,N_16628);
xor U17164 (N_17164,N_16429,N_16419);
and U17165 (N_17165,N_16768,N_16543);
and U17166 (N_17166,N_16594,N_16655);
xor U17167 (N_17167,N_16651,N_16639);
nor U17168 (N_17168,N_16437,N_16522);
nand U17169 (N_17169,N_16530,N_16425);
nor U17170 (N_17170,N_16640,N_16737);
nor U17171 (N_17171,N_16537,N_16552);
and U17172 (N_17172,N_16662,N_16723);
and U17173 (N_17173,N_16649,N_16622);
nand U17174 (N_17174,N_16463,N_16581);
nand U17175 (N_17175,N_16625,N_16567);
and U17176 (N_17176,N_16589,N_16422);
nand U17177 (N_17177,N_16605,N_16466);
nor U17178 (N_17178,N_16741,N_16576);
or U17179 (N_17179,N_16663,N_16729);
and U17180 (N_17180,N_16436,N_16753);
nor U17181 (N_17181,N_16798,N_16699);
and U17182 (N_17182,N_16734,N_16472);
nor U17183 (N_17183,N_16413,N_16737);
nor U17184 (N_17184,N_16654,N_16641);
xnor U17185 (N_17185,N_16583,N_16653);
or U17186 (N_17186,N_16627,N_16579);
and U17187 (N_17187,N_16688,N_16591);
and U17188 (N_17188,N_16481,N_16635);
xnor U17189 (N_17189,N_16721,N_16481);
or U17190 (N_17190,N_16576,N_16483);
nand U17191 (N_17191,N_16748,N_16518);
and U17192 (N_17192,N_16748,N_16674);
nor U17193 (N_17193,N_16555,N_16507);
and U17194 (N_17194,N_16521,N_16679);
nand U17195 (N_17195,N_16778,N_16658);
and U17196 (N_17196,N_16708,N_16498);
and U17197 (N_17197,N_16490,N_16768);
xor U17198 (N_17198,N_16438,N_16408);
and U17199 (N_17199,N_16766,N_16662);
nor U17200 (N_17200,N_17035,N_16862);
xnor U17201 (N_17201,N_17127,N_17114);
and U17202 (N_17202,N_16938,N_16936);
nor U17203 (N_17203,N_17084,N_16836);
xor U17204 (N_17204,N_16863,N_17030);
xor U17205 (N_17205,N_16985,N_17181);
nor U17206 (N_17206,N_17109,N_16963);
xnor U17207 (N_17207,N_16926,N_17031);
nor U17208 (N_17208,N_17088,N_16902);
nor U17209 (N_17209,N_16982,N_17089);
or U17210 (N_17210,N_17072,N_16945);
nor U17211 (N_17211,N_16823,N_17070);
nand U17212 (N_17212,N_17166,N_17029);
xnor U17213 (N_17213,N_17157,N_16852);
nand U17214 (N_17214,N_17062,N_17074);
xor U17215 (N_17215,N_17125,N_16988);
and U17216 (N_17216,N_16879,N_16978);
or U17217 (N_17217,N_17052,N_16972);
or U17218 (N_17218,N_16832,N_17008);
nor U17219 (N_17219,N_16840,N_17093);
xnor U17220 (N_17220,N_17133,N_16843);
nor U17221 (N_17221,N_16890,N_17020);
and U17222 (N_17222,N_16921,N_16818);
and U17223 (N_17223,N_17021,N_16971);
xnor U17224 (N_17224,N_17078,N_16829);
and U17225 (N_17225,N_16857,N_17150);
xor U17226 (N_17226,N_16946,N_16990);
nor U17227 (N_17227,N_16906,N_17138);
nand U17228 (N_17228,N_17082,N_16922);
or U17229 (N_17229,N_17137,N_17081);
xor U17230 (N_17230,N_16868,N_17152);
and U17231 (N_17231,N_17180,N_16838);
nor U17232 (N_17232,N_16809,N_17048);
or U17233 (N_17233,N_17095,N_16846);
nor U17234 (N_17234,N_17184,N_17186);
nor U17235 (N_17235,N_17174,N_17019);
and U17236 (N_17236,N_16820,N_17053);
and U17237 (N_17237,N_17050,N_16804);
and U17238 (N_17238,N_16911,N_16958);
nand U17239 (N_17239,N_16813,N_16930);
nand U17240 (N_17240,N_17059,N_16835);
nor U17241 (N_17241,N_17124,N_17042);
nor U17242 (N_17242,N_16855,N_17037);
and U17243 (N_17243,N_17135,N_16924);
or U17244 (N_17244,N_16912,N_17141);
xnor U17245 (N_17245,N_17147,N_17188);
or U17246 (N_17246,N_17120,N_17002);
nor U17247 (N_17247,N_16901,N_16967);
or U17248 (N_17248,N_16872,N_16827);
nand U17249 (N_17249,N_16894,N_16933);
and U17250 (N_17250,N_17017,N_17055);
and U17251 (N_17251,N_17000,N_16875);
xnor U17252 (N_17252,N_17061,N_16960);
and U17253 (N_17253,N_17197,N_16842);
and U17254 (N_17254,N_16854,N_16889);
xor U17255 (N_17255,N_16919,N_16821);
or U17256 (N_17256,N_17145,N_17027);
nand U17257 (N_17257,N_16943,N_17163);
nor U17258 (N_17258,N_16801,N_17116);
and U17259 (N_17259,N_17032,N_17190);
and U17260 (N_17260,N_17057,N_16909);
nand U17261 (N_17261,N_16815,N_17126);
nand U17262 (N_17262,N_16989,N_17170);
nand U17263 (N_17263,N_16810,N_16914);
nor U17264 (N_17264,N_17199,N_17117);
nand U17265 (N_17265,N_16830,N_17155);
or U17266 (N_17266,N_16940,N_16987);
and U17267 (N_17267,N_17187,N_17183);
nand U17268 (N_17268,N_16848,N_16931);
or U17269 (N_17269,N_17179,N_16891);
and U17270 (N_17270,N_16952,N_17142);
or U17271 (N_17271,N_16976,N_17130);
or U17272 (N_17272,N_16867,N_16900);
nand U17273 (N_17273,N_16893,N_17169);
nor U17274 (N_17274,N_17079,N_16844);
or U17275 (N_17275,N_17185,N_16925);
or U17276 (N_17276,N_17077,N_17009);
or U17277 (N_17277,N_16850,N_17086);
and U17278 (N_17278,N_17143,N_17098);
xnor U17279 (N_17279,N_16883,N_16929);
nand U17280 (N_17280,N_17006,N_16884);
or U17281 (N_17281,N_16950,N_16897);
nor U17282 (N_17282,N_16845,N_17063);
xor U17283 (N_17283,N_16856,N_16837);
and U17284 (N_17284,N_17051,N_17039);
nor U17285 (N_17285,N_17054,N_16917);
xor U17286 (N_17286,N_17043,N_16920);
nand U17287 (N_17287,N_16955,N_16876);
nor U17288 (N_17288,N_17195,N_17038);
nor U17289 (N_17289,N_17164,N_16977);
xnor U17290 (N_17290,N_17097,N_16904);
xor U17291 (N_17291,N_17122,N_17131);
or U17292 (N_17292,N_17171,N_16824);
xnor U17293 (N_17293,N_17129,N_16953);
nor U17294 (N_17294,N_17191,N_17162);
or U17295 (N_17295,N_17026,N_16887);
nor U17296 (N_17296,N_16803,N_16928);
or U17297 (N_17297,N_17119,N_17041);
and U17298 (N_17298,N_16905,N_17121);
and U17299 (N_17299,N_16993,N_16834);
nand U17300 (N_17300,N_16881,N_17044);
and U17301 (N_17301,N_17069,N_16828);
or U17302 (N_17302,N_16907,N_17115);
nand U17303 (N_17303,N_17146,N_17189);
or U17304 (N_17304,N_17011,N_17148);
or U17305 (N_17305,N_16878,N_16973);
nor U17306 (N_17306,N_16870,N_17075);
or U17307 (N_17307,N_16877,N_16849);
nand U17308 (N_17308,N_17104,N_16961);
nor U17309 (N_17309,N_17046,N_17112);
or U17310 (N_17310,N_17005,N_17024);
nand U17311 (N_17311,N_16941,N_16861);
nand U17312 (N_17312,N_16954,N_17103);
nor U17313 (N_17313,N_17108,N_17192);
nand U17314 (N_17314,N_16984,N_17036);
or U17315 (N_17315,N_17058,N_16979);
or U17316 (N_17316,N_16981,N_17165);
nor U17317 (N_17317,N_16825,N_17014);
nand U17318 (N_17318,N_16847,N_17105);
and U17319 (N_17319,N_16970,N_17159);
xnor U17320 (N_17320,N_16858,N_16948);
nand U17321 (N_17321,N_16860,N_16975);
nor U17322 (N_17322,N_16910,N_17100);
nor U17323 (N_17323,N_16811,N_17068);
nor U17324 (N_17324,N_16956,N_17139);
nor U17325 (N_17325,N_17160,N_16916);
nor U17326 (N_17326,N_17004,N_17007);
nor U17327 (N_17327,N_16962,N_16998);
nand U17328 (N_17328,N_16944,N_17132);
or U17329 (N_17329,N_16964,N_17060);
and U17330 (N_17330,N_16807,N_17151);
nor U17331 (N_17331,N_17056,N_16898);
xnor U17332 (N_17332,N_16888,N_16817);
or U17333 (N_17333,N_16934,N_16822);
and U17334 (N_17334,N_16974,N_17111);
or U17335 (N_17335,N_17182,N_16996);
nor U17336 (N_17336,N_17194,N_17136);
and U17337 (N_17337,N_17092,N_16992);
nor U17338 (N_17338,N_16800,N_17045);
or U17339 (N_17339,N_16874,N_16947);
or U17340 (N_17340,N_17025,N_17010);
or U17341 (N_17341,N_16957,N_17012);
nand U17342 (N_17342,N_16969,N_16923);
and U17343 (N_17343,N_17066,N_16932);
xnor U17344 (N_17344,N_17175,N_16995);
xnor U17345 (N_17345,N_17144,N_17101);
xnor U17346 (N_17346,N_16968,N_17177);
nand U17347 (N_17347,N_16997,N_16939);
or U17348 (N_17348,N_17167,N_16983);
nand U17349 (N_17349,N_17064,N_16986);
and U17350 (N_17350,N_17033,N_16859);
nor U17351 (N_17351,N_17003,N_17196);
or U17352 (N_17352,N_16880,N_16873);
nand U17353 (N_17353,N_16966,N_16895);
or U17354 (N_17354,N_17083,N_17065);
nand U17355 (N_17355,N_17015,N_17173);
and U17356 (N_17356,N_16814,N_16866);
nor U17357 (N_17357,N_17113,N_17154);
nor U17358 (N_17358,N_16913,N_16965);
nand U17359 (N_17359,N_17016,N_17134);
and U17360 (N_17360,N_16853,N_17128);
xnor U17361 (N_17361,N_17087,N_16885);
xnor U17362 (N_17362,N_16808,N_17073);
nand U17363 (N_17363,N_16882,N_17023);
xor U17364 (N_17364,N_16994,N_17153);
xnor U17365 (N_17365,N_16959,N_16927);
and U17366 (N_17366,N_17156,N_17047);
xnor U17367 (N_17367,N_17071,N_17176);
xor U17368 (N_17368,N_16871,N_17091);
and U17369 (N_17369,N_16851,N_17040);
or U17370 (N_17370,N_17034,N_17080);
nor U17371 (N_17371,N_17161,N_16865);
nand U17372 (N_17372,N_17090,N_17076);
xnor U17373 (N_17373,N_16831,N_16951);
and U17374 (N_17374,N_17158,N_17028);
and U17375 (N_17375,N_17118,N_17123);
xnor U17376 (N_17376,N_16918,N_16806);
nor U17377 (N_17377,N_16816,N_17193);
xor U17378 (N_17378,N_17049,N_17168);
nor U17379 (N_17379,N_16991,N_16826);
nand U17380 (N_17380,N_17178,N_16805);
and U17381 (N_17381,N_17018,N_16819);
or U17382 (N_17382,N_17198,N_17001);
xnor U17383 (N_17383,N_17149,N_17013);
or U17384 (N_17384,N_16903,N_17085);
or U17385 (N_17385,N_16942,N_16999);
and U17386 (N_17386,N_17094,N_16841);
nor U17387 (N_17387,N_16896,N_16908);
and U17388 (N_17388,N_16892,N_17022);
xor U17389 (N_17389,N_16937,N_16949);
or U17390 (N_17390,N_16886,N_16812);
or U17391 (N_17391,N_16980,N_16802);
and U17392 (N_17392,N_17102,N_17067);
or U17393 (N_17393,N_16839,N_16864);
or U17394 (N_17394,N_16915,N_17172);
nand U17395 (N_17395,N_17107,N_16899);
and U17396 (N_17396,N_16869,N_16935);
nand U17397 (N_17397,N_17099,N_17140);
or U17398 (N_17398,N_17106,N_17110);
xor U17399 (N_17399,N_17096,N_16833);
or U17400 (N_17400,N_17118,N_17111);
or U17401 (N_17401,N_17126,N_16859);
nand U17402 (N_17402,N_16950,N_17146);
nand U17403 (N_17403,N_16887,N_16832);
nor U17404 (N_17404,N_16960,N_17195);
and U17405 (N_17405,N_16961,N_16818);
or U17406 (N_17406,N_16999,N_16923);
nor U17407 (N_17407,N_17195,N_16813);
nor U17408 (N_17408,N_16971,N_16801);
and U17409 (N_17409,N_17097,N_17120);
xnor U17410 (N_17410,N_17122,N_16841);
nor U17411 (N_17411,N_16841,N_17090);
xor U17412 (N_17412,N_17149,N_16818);
or U17413 (N_17413,N_16948,N_16949);
nor U17414 (N_17414,N_16826,N_16884);
nor U17415 (N_17415,N_16990,N_16913);
and U17416 (N_17416,N_16857,N_16836);
nand U17417 (N_17417,N_17011,N_16940);
nor U17418 (N_17418,N_17153,N_16863);
nor U17419 (N_17419,N_16928,N_17189);
and U17420 (N_17420,N_16898,N_16845);
nor U17421 (N_17421,N_17100,N_17099);
and U17422 (N_17422,N_16876,N_16963);
or U17423 (N_17423,N_16961,N_16840);
and U17424 (N_17424,N_16963,N_16837);
and U17425 (N_17425,N_16947,N_17025);
or U17426 (N_17426,N_17122,N_16957);
and U17427 (N_17427,N_17140,N_16919);
nor U17428 (N_17428,N_16839,N_17123);
and U17429 (N_17429,N_16810,N_16983);
xnor U17430 (N_17430,N_17020,N_17002);
xor U17431 (N_17431,N_17172,N_17020);
or U17432 (N_17432,N_16853,N_17070);
or U17433 (N_17433,N_17071,N_17001);
xor U17434 (N_17434,N_17030,N_16862);
nor U17435 (N_17435,N_17193,N_17082);
nand U17436 (N_17436,N_17165,N_17040);
xnor U17437 (N_17437,N_16958,N_17118);
nor U17438 (N_17438,N_17001,N_16816);
nor U17439 (N_17439,N_17005,N_16982);
or U17440 (N_17440,N_17151,N_17085);
nand U17441 (N_17441,N_17079,N_16931);
xor U17442 (N_17442,N_17005,N_17085);
or U17443 (N_17443,N_17157,N_16916);
xor U17444 (N_17444,N_17110,N_17148);
nor U17445 (N_17445,N_17101,N_16913);
and U17446 (N_17446,N_17193,N_16888);
xnor U17447 (N_17447,N_17080,N_16972);
or U17448 (N_17448,N_17052,N_16900);
and U17449 (N_17449,N_16964,N_17066);
and U17450 (N_17450,N_16885,N_17002);
and U17451 (N_17451,N_16800,N_17189);
or U17452 (N_17452,N_16912,N_16985);
and U17453 (N_17453,N_17111,N_17122);
nor U17454 (N_17454,N_17152,N_16851);
nand U17455 (N_17455,N_16938,N_17096);
or U17456 (N_17456,N_16807,N_16985);
and U17457 (N_17457,N_17090,N_17035);
and U17458 (N_17458,N_16933,N_16868);
or U17459 (N_17459,N_17007,N_16960);
and U17460 (N_17460,N_16988,N_17173);
xnor U17461 (N_17461,N_17132,N_17100);
xor U17462 (N_17462,N_17044,N_17137);
and U17463 (N_17463,N_16824,N_16889);
and U17464 (N_17464,N_17174,N_17118);
or U17465 (N_17465,N_17001,N_16921);
xnor U17466 (N_17466,N_17104,N_16985);
or U17467 (N_17467,N_17096,N_17053);
or U17468 (N_17468,N_17123,N_17198);
or U17469 (N_17469,N_17149,N_17027);
or U17470 (N_17470,N_16960,N_16841);
or U17471 (N_17471,N_16861,N_16802);
nor U17472 (N_17472,N_17158,N_16914);
or U17473 (N_17473,N_16930,N_17101);
or U17474 (N_17474,N_17092,N_16995);
nand U17475 (N_17475,N_17150,N_16866);
xor U17476 (N_17476,N_16957,N_17133);
nor U17477 (N_17477,N_16893,N_17135);
or U17478 (N_17478,N_17074,N_16835);
and U17479 (N_17479,N_17172,N_16955);
and U17480 (N_17480,N_16836,N_16848);
or U17481 (N_17481,N_16906,N_16987);
nor U17482 (N_17482,N_16836,N_16850);
nor U17483 (N_17483,N_17119,N_17018);
nand U17484 (N_17484,N_17000,N_17060);
nor U17485 (N_17485,N_17076,N_16925);
and U17486 (N_17486,N_16968,N_16870);
and U17487 (N_17487,N_17118,N_16891);
nor U17488 (N_17488,N_17119,N_17089);
nand U17489 (N_17489,N_16960,N_16950);
or U17490 (N_17490,N_16938,N_17015);
xor U17491 (N_17491,N_16993,N_17022);
nand U17492 (N_17492,N_17184,N_16958);
nand U17493 (N_17493,N_17185,N_16841);
or U17494 (N_17494,N_16813,N_16833);
or U17495 (N_17495,N_16947,N_16970);
nand U17496 (N_17496,N_17197,N_16908);
and U17497 (N_17497,N_16875,N_16824);
or U17498 (N_17498,N_17053,N_17150);
or U17499 (N_17499,N_17110,N_17009);
nor U17500 (N_17500,N_16826,N_16934);
nand U17501 (N_17501,N_17026,N_16961);
or U17502 (N_17502,N_17181,N_17003);
nand U17503 (N_17503,N_17166,N_16814);
nor U17504 (N_17504,N_16814,N_16815);
and U17505 (N_17505,N_16860,N_17023);
nand U17506 (N_17506,N_17040,N_17153);
xnor U17507 (N_17507,N_16851,N_16905);
nand U17508 (N_17508,N_16852,N_17021);
nor U17509 (N_17509,N_16973,N_17115);
nor U17510 (N_17510,N_17171,N_17034);
or U17511 (N_17511,N_16826,N_17191);
xnor U17512 (N_17512,N_17168,N_16923);
nor U17513 (N_17513,N_16817,N_16824);
nor U17514 (N_17514,N_16939,N_16812);
nand U17515 (N_17515,N_16813,N_17191);
nand U17516 (N_17516,N_16887,N_16823);
nand U17517 (N_17517,N_16905,N_16935);
or U17518 (N_17518,N_16885,N_17086);
or U17519 (N_17519,N_16854,N_16869);
or U17520 (N_17520,N_17189,N_16990);
nor U17521 (N_17521,N_17114,N_16955);
or U17522 (N_17522,N_16852,N_17117);
nand U17523 (N_17523,N_17031,N_17009);
nand U17524 (N_17524,N_17102,N_17153);
nor U17525 (N_17525,N_16816,N_17002);
and U17526 (N_17526,N_16860,N_16847);
or U17527 (N_17527,N_16873,N_16854);
or U17528 (N_17528,N_17133,N_17175);
nand U17529 (N_17529,N_17182,N_17125);
nor U17530 (N_17530,N_16872,N_17189);
nand U17531 (N_17531,N_16834,N_17007);
and U17532 (N_17532,N_16889,N_16815);
and U17533 (N_17533,N_17085,N_17001);
nand U17534 (N_17534,N_16800,N_16905);
nand U17535 (N_17535,N_17078,N_17062);
xor U17536 (N_17536,N_16943,N_17008);
xnor U17537 (N_17537,N_16922,N_16806);
xor U17538 (N_17538,N_16996,N_16891);
and U17539 (N_17539,N_16854,N_17128);
and U17540 (N_17540,N_16920,N_17104);
and U17541 (N_17541,N_17122,N_16971);
nand U17542 (N_17542,N_16871,N_16952);
nor U17543 (N_17543,N_16809,N_17014);
or U17544 (N_17544,N_17181,N_17034);
nor U17545 (N_17545,N_17196,N_16981);
xnor U17546 (N_17546,N_16959,N_16964);
xor U17547 (N_17547,N_17124,N_17012);
and U17548 (N_17548,N_17063,N_16891);
or U17549 (N_17549,N_17198,N_17082);
xor U17550 (N_17550,N_17105,N_16841);
nand U17551 (N_17551,N_16865,N_17010);
or U17552 (N_17552,N_16856,N_16893);
or U17553 (N_17553,N_17084,N_16881);
nor U17554 (N_17554,N_17134,N_16826);
xor U17555 (N_17555,N_17196,N_16959);
xnor U17556 (N_17556,N_17199,N_17044);
nand U17557 (N_17557,N_16874,N_16854);
xor U17558 (N_17558,N_17162,N_17192);
or U17559 (N_17559,N_16809,N_17077);
nand U17560 (N_17560,N_17182,N_17068);
or U17561 (N_17561,N_16888,N_16911);
nand U17562 (N_17562,N_17130,N_16960);
xor U17563 (N_17563,N_17101,N_17047);
nor U17564 (N_17564,N_16907,N_17050);
nand U17565 (N_17565,N_17153,N_16989);
nor U17566 (N_17566,N_16801,N_16979);
and U17567 (N_17567,N_17194,N_16883);
xnor U17568 (N_17568,N_16971,N_17178);
nor U17569 (N_17569,N_16810,N_16943);
nand U17570 (N_17570,N_16814,N_16937);
nor U17571 (N_17571,N_17148,N_16846);
nand U17572 (N_17572,N_17000,N_17135);
nor U17573 (N_17573,N_16923,N_17141);
nand U17574 (N_17574,N_17148,N_17166);
or U17575 (N_17575,N_17003,N_16866);
nand U17576 (N_17576,N_17106,N_17084);
or U17577 (N_17577,N_17107,N_17140);
nand U17578 (N_17578,N_16991,N_16844);
nor U17579 (N_17579,N_16856,N_17117);
nand U17580 (N_17580,N_17167,N_16949);
xnor U17581 (N_17581,N_16901,N_17157);
and U17582 (N_17582,N_16952,N_16929);
xnor U17583 (N_17583,N_17120,N_16807);
or U17584 (N_17584,N_17050,N_16861);
and U17585 (N_17585,N_17171,N_17114);
or U17586 (N_17586,N_17093,N_16863);
or U17587 (N_17587,N_17008,N_16970);
nand U17588 (N_17588,N_17182,N_17060);
xnor U17589 (N_17589,N_16809,N_17130);
or U17590 (N_17590,N_16920,N_17090);
and U17591 (N_17591,N_17086,N_16844);
and U17592 (N_17592,N_16937,N_16942);
xnor U17593 (N_17593,N_17186,N_16802);
nand U17594 (N_17594,N_17016,N_16940);
xnor U17595 (N_17595,N_16822,N_17169);
nand U17596 (N_17596,N_16896,N_16882);
xor U17597 (N_17597,N_17155,N_17142);
nand U17598 (N_17598,N_16972,N_16954);
or U17599 (N_17599,N_16957,N_16984);
and U17600 (N_17600,N_17391,N_17570);
xnor U17601 (N_17601,N_17498,N_17386);
or U17602 (N_17602,N_17238,N_17257);
nand U17603 (N_17603,N_17338,N_17354);
or U17604 (N_17604,N_17266,N_17526);
or U17605 (N_17605,N_17418,N_17421);
nand U17606 (N_17606,N_17561,N_17237);
nand U17607 (N_17607,N_17568,N_17360);
xnor U17608 (N_17608,N_17283,N_17542);
and U17609 (N_17609,N_17582,N_17328);
xnor U17610 (N_17610,N_17554,N_17477);
nor U17611 (N_17611,N_17289,N_17510);
nand U17612 (N_17612,N_17430,N_17446);
nand U17613 (N_17613,N_17547,N_17507);
xnor U17614 (N_17614,N_17303,N_17520);
nor U17615 (N_17615,N_17545,N_17374);
xor U17616 (N_17616,N_17341,N_17455);
or U17617 (N_17617,N_17308,N_17415);
xor U17618 (N_17618,N_17471,N_17594);
nor U17619 (N_17619,N_17497,N_17527);
and U17620 (N_17620,N_17433,N_17427);
xnor U17621 (N_17621,N_17440,N_17249);
and U17622 (N_17622,N_17394,N_17295);
and U17623 (N_17623,N_17371,N_17368);
nand U17624 (N_17624,N_17343,N_17284);
and U17625 (N_17625,N_17550,N_17382);
xor U17626 (N_17626,N_17327,N_17480);
nor U17627 (N_17627,N_17560,N_17558);
xor U17628 (N_17628,N_17207,N_17276);
xor U17629 (N_17629,N_17468,N_17378);
xor U17630 (N_17630,N_17204,N_17512);
xor U17631 (N_17631,N_17333,N_17346);
or U17632 (N_17632,N_17272,N_17592);
nor U17633 (N_17633,N_17541,N_17205);
xor U17634 (N_17634,N_17364,N_17254);
and U17635 (N_17635,N_17400,N_17267);
or U17636 (N_17636,N_17574,N_17564);
or U17637 (N_17637,N_17598,N_17302);
and U17638 (N_17638,N_17451,N_17465);
xnor U17639 (N_17639,N_17460,N_17385);
or U17640 (N_17640,N_17401,N_17549);
and U17641 (N_17641,N_17369,N_17273);
nand U17642 (N_17642,N_17201,N_17226);
nor U17643 (N_17643,N_17423,N_17563);
and U17644 (N_17644,N_17467,N_17488);
or U17645 (N_17645,N_17531,N_17405);
and U17646 (N_17646,N_17297,N_17265);
or U17647 (N_17647,N_17412,N_17450);
xnor U17648 (N_17648,N_17219,N_17492);
or U17649 (N_17649,N_17387,N_17370);
and U17650 (N_17650,N_17355,N_17458);
or U17651 (N_17651,N_17392,N_17281);
and U17652 (N_17652,N_17350,N_17268);
xnor U17653 (N_17653,N_17389,N_17588);
and U17654 (N_17654,N_17390,N_17539);
and U17655 (N_17655,N_17524,N_17571);
or U17656 (N_17656,N_17383,N_17584);
xor U17657 (N_17657,N_17351,N_17483);
or U17658 (N_17658,N_17376,N_17280);
nand U17659 (N_17659,N_17326,N_17323);
nor U17660 (N_17660,N_17573,N_17208);
nor U17661 (N_17661,N_17453,N_17525);
xor U17662 (N_17662,N_17230,N_17292);
nor U17663 (N_17663,N_17528,N_17210);
or U17664 (N_17664,N_17569,N_17589);
nor U17665 (N_17665,N_17250,N_17288);
nand U17666 (N_17666,N_17585,N_17414);
nand U17667 (N_17667,N_17435,N_17486);
nor U17668 (N_17668,N_17479,N_17363);
and U17669 (N_17669,N_17517,N_17220);
nor U17670 (N_17670,N_17321,N_17565);
nor U17671 (N_17671,N_17474,N_17529);
and U17672 (N_17672,N_17264,N_17461);
nor U17673 (N_17673,N_17431,N_17499);
and U17674 (N_17674,N_17519,N_17214);
nand U17675 (N_17675,N_17339,N_17318);
nor U17676 (N_17676,N_17501,N_17227);
nand U17677 (N_17677,N_17434,N_17365);
nand U17678 (N_17678,N_17506,N_17239);
nand U17679 (N_17679,N_17409,N_17322);
nand U17680 (N_17680,N_17299,N_17375);
xnor U17681 (N_17681,N_17305,N_17263);
xor U17682 (N_17682,N_17411,N_17271);
and U17683 (N_17683,N_17353,N_17223);
nand U17684 (N_17684,N_17330,N_17590);
or U17685 (N_17685,N_17438,N_17398);
nor U17686 (N_17686,N_17535,N_17315);
nor U17687 (N_17687,N_17285,N_17314);
nand U17688 (N_17688,N_17290,N_17359);
xnor U17689 (N_17689,N_17576,N_17247);
and U17690 (N_17690,N_17566,N_17206);
xnor U17691 (N_17691,N_17599,N_17437);
xnor U17692 (N_17692,N_17511,N_17296);
and U17693 (N_17693,N_17429,N_17252);
and U17694 (N_17694,N_17476,N_17522);
or U17695 (N_17695,N_17259,N_17540);
nand U17696 (N_17696,N_17551,N_17472);
or U17697 (N_17697,N_17457,N_17523);
xor U17698 (N_17698,N_17513,N_17335);
xor U17699 (N_17699,N_17396,N_17262);
xor U17700 (N_17700,N_17203,N_17586);
xnor U17701 (N_17701,N_17393,N_17298);
or U17702 (N_17702,N_17381,N_17340);
xnor U17703 (N_17703,N_17441,N_17362);
nand U17704 (N_17704,N_17543,N_17337);
xor U17705 (N_17705,N_17482,N_17417);
nor U17706 (N_17706,N_17278,N_17304);
and U17707 (N_17707,N_17242,N_17319);
and U17708 (N_17708,N_17478,N_17253);
nor U17709 (N_17709,N_17518,N_17231);
and U17710 (N_17710,N_17222,N_17361);
nand U17711 (N_17711,N_17596,N_17533);
xor U17712 (N_17712,N_17348,N_17494);
nand U17713 (N_17713,N_17384,N_17552);
and U17714 (N_17714,N_17424,N_17491);
nand U17715 (N_17715,N_17502,N_17516);
or U17716 (N_17716,N_17397,N_17442);
xor U17717 (N_17717,N_17228,N_17279);
xor U17718 (N_17718,N_17293,N_17349);
nand U17719 (N_17719,N_17420,N_17216);
and U17720 (N_17720,N_17294,N_17320);
nor U17721 (N_17721,N_17422,N_17342);
nand U17722 (N_17722,N_17403,N_17557);
and U17723 (N_17723,N_17372,N_17311);
nand U17724 (N_17724,N_17240,N_17331);
xnor U17725 (N_17725,N_17277,N_17466);
nand U17726 (N_17726,N_17530,N_17505);
nand U17727 (N_17727,N_17515,N_17291);
and U17728 (N_17728,N_17444,N_17470);
nand U17729 (N_17729,N_17258,N_17274);
or U17730 (N_17730,N_17555,N_17218);
nor U17731 (N_17731,N_17200,N_17357);
nand U17732 (N_17732,N_17581,N_17336);
or U17733 (N_17733,N_17225,N_17232);
or U17734 (N_17734,N_17439,N_17413);
nor U17735 (N_17735,N_17324,N_17312);
or U17736 (N_17736,N_17309,N_17593);
and U17737 (N_17737,N_17202,N_17416);
and U17738 (N_17738,N_17495,N_17493);
xor U17739 (N_17739,N_17452,N_17241);
or U17740 (N_17740,N_17356,N_17432);
or U17741 (N_17741,N_17487,N_17306);
nor U17742 (N_17742,N_17402,N_17211);
xnor U17743 (N_17743,N_17251,N_17475);
or U17744 (N_17744,N_17233,N_17408);
xor U17745 (N_17745,N_17246,N_17462);
nor U17746 (N_17746,N_17484,N_17256);
or U17747 (N_17747,N_17469,N_17436);
xnor U17748 (N_17748,N_17559,N_17504);
nor U17749 (N_17749,N_17485,N_17538);
xor U17750 (N_17750,N_17345,N_17366);
xnor U17751 (N_17751,N_17591,N_17443);
or U17752 (N_17752,N_17229,N_17380);
xor U17753 (N_17753,N_17329,N_17500);
or U17754 (N_17754,N_17217,N_17358);
nor U17755 (N_17755,N_17379,N_17532);
nor U17756 (N_17756,N_17367,N_17514);
and U17757 (N_17757,N_17334,N_17445);
nand U17758 (N_17758,N_17377,N_17473);
nor U17759 (N_17759,N_17419,N_17399);
xor U17760 (N_17760,N_17406,N_17286);
xor U17761 (N_17761,N_17496,N_17572);
and U17762 (N_17762,N_17261,N_17587);
or U17763 (N_17763,N_17248,N_17508);
or U17764 (N_17764,N_17553,N_17235);
nor U17765 (N_17765,N_17301,N_17300);
nor U17766 (N_17766,N_17234,N_17347);
and U17767 (N_17767,N_17307,N_17395);
nor U17768 (N_17768,N_17580,N_17410);
nor U17769 (N_17769,N_17454,N_17224);
nor U17770 (N_17770,N_17464,N_17583);
nor U17771 (N_17771,N_17260,N_17577);
and U17772 (N_17772,N_17352,N_17428);
xor U17773 (N_17773,N_17310,N_17578);
and U17774 (N_17774,N_17490,N_17509);
nor U17775 (N_17775,N_17536,N_17562);
and U17776 (N_17776,N_17544,N_17317);
nand U17777 (N_17777,N_17534,N_17537);
and U17778 (N_17778,N_17597,N_17344);
nand U17779 (N_17779,N_17213,N_17316);
nor U17780 (N_17780,N_17244,N_17325);
nor U17781 (N_17781,N_17255,N_17425);
xor U17782 (N_17782,N_17521,N_17243);
nand U17783 (N_17783,N_17459,N_17209);
xnor U17784 (N_17784,N_17503,N_17481);
and U17785 (N_17785,N_17332,N_17489);
nor U17786 (N_17786,N_17595,N_17426);
and U17787 (N_17787,N_17546,N_17236);
and U17788 (N_17788,N_17407,N_17548);
and U17789 (N_17789,N_17388,N_17463);
nor U17790 (N_17790,N_17269,N_17221);
xnor U17791 (N_17791,N_17287,N_17579);
nor U17792 (N_17792,N_17282,N_17373);
xnor U17793 (N_17793,N_17456,N_17245);
and U17794 (N_17794,N_17567,N_17313);
nand U17795 (N_17795,N_17448,N_17556);
nand U17796 (N_17796,N_17575,N_17404);
nor U17797 (N_17797,N_17215,N_17212);
nand U17798 (N_17798,N_17447,N_17270);
and U17799 (N_17799,N_17449,N_17275);
xor U17800 (N_17800,N_17300,N_17548);
nor U17801 (N_17801,N_17486,N_17573);
or U17802 (N_17802,N_17490,N_17267);
and U17803 (N_17803,N_17232,N_17458);
and U17804 (N_17804,N_17307,N_17309);
nand U17805 (N_17805,N_17235,N_17598);
or U17806 (N_17806,N_17297,N_17459);
xor U17807 (N_17807,N_17467,N_17566);
and U17808 (N_17808,N_17593,N_17223);
nor U17809 (N_17809,N_17405,N_17331);
and U17810 (N_17810,N_17484,N_17460);
or U17811 (N_17811,N_17269,N_17566);
nand U17812 (N_17812,N_17327,N_17227);
and U17813 (N_17813,N_17224,N_17563);
nand U17814 (N_17814,N_17522,N_17293);
or U17815 (N_17815,N_17259,N_17320);
nor U17816 (N_17816,N_17222,N_17254);
nand U17817 (N_17817,N_17251,N_17449);
nand U17818 (N_17818,N_17267,N_17246);
or U17819 (N_17819,N_17385,N_17338);
and U17820 (N_17820,N_17409,N_17382);
or U17821 (N_17821,N_17382,N_17255);
xnor U17822 (N_17822,N_17381,N_17254);
and U17823 (N_17823,N_17583,N_17580);
nand U17824 (N_17824,N_17410,N_17243);
nand U17825 (N_17825,N_17506,N_17308);
nor U17826 (N_17826,N_17281,N_17371);
nor U17827 (N_17827,N_17599,N_17207);
nand U17828 (N_17828,N_17370,N_17331);
or U17829 (N_17829,N_17228,N_17545);
nand U17830 (N_17830,N_17539,N_17362);
and U17831 (N_17831,N_17473,N_17503);
or U17832 (N_17832,N_17367,N_17414);
nand U17833 (N_17833,N_17358,N_17575);
and U17834 (N_17834,N_17537,N_17309);
or U17835 (N_17835,N_17434,N_17519);
nand U17836 (N_17836,N_17492,N_17234);
and U17837 (N_17837,N_17507,N_17369);
nor U17838 (N_17838,N_17430,N_17359);
nor U17839 (N_17839,N_17246,N_17508);
and U17840 (N_17840,N_17578,N_17260);
or U17841 (N_17841,N_17354,N_17445);
xor U17842 (N_17842,N_17465,N_17410);
or U17843 (N_17843,N_17563,N_17363);
nor U17844 (N_17844,N_17222,N_17252);
nand U17845 (N_17845,N_17204,N_17377);
xor U17846 (N_17846,N_17486,N_17468);
nor U17847 (N_17847,N_17423,N_17532);
nand U17848 (N_17848,N_17412,N_17553);
nor U17849 (N_17849,N_17342,N_17488);
xor U17850 (N_17850,N_17311,N_17237);
and U17851 (N_17851,N_17588,N_17305);
nand U17852 (N_17852,N_17442,N_17290);
xnor U17853 (N_17853,N_17436,N_17322);
and U17854 (N_17854,N_17553,N_17520);
nor U17855 (N_17855,N_17438,N_17268);
or U17856 (N_17856,N_17485,N_17469);
nor U17857 (N_17857,N_17465,N_17430);
nor U17858 (N_17858,N_17433,N_17226);
nor U17859 (N_17859,N_17244,N_17540);
or U17860 (N_17860,N_17251,N_17369);
nand U17861 (N_17861,N_17216,N_17534);
nand U17862 (N_17862,N_17309,N_17202);
nand U17863 (N_17863,N_17472,N_17530);
or U17864 (N_17864,N_17325,N_17202);
nor U17865 (N_17865,N_17511,N_17200);
nor U17866 (N_17866,N_17555,N_17413);
or U17867 (N_17867,N_17445,N_17513);
nor U17868 (N_17868,N_17454,N_17461);
xnor U17869 (N_17869,N_17206,N_17496);
or U17870 (N_17870,N_17287,N_17585);
xnor U17871 (N_17871,N_17281,N_17437);
and U17872 (N_17872,N_17241,N_17373);
or U17873 (N_17873,N_17480,N_17404);
xor U17874 (N_17874,N_17440,N_17332);
and U17875 (N_17875,N_17440,N_17513);
or U17876 (N_17876,N_17237,N_17256);
or U17877 (N_17877,N_17332,N_17266);
or U17878 (N_17878,N_17431,N_17340);
nand U17879 (N_17879,N_17534,N_17473);
nand U17880 (N_17880,N_17232,N_17265);
nand U17881 (N_17881,N_17382,N_17517);
or U17882 (N_17882,N_17396,N_17542);
nand U17883 (N_17883,N_17408,N_17503);
or U17884 (N_17884,N_17531,N_17384);
or U17885 (N_17885,N_17332,N_17338);
xor U17886 (N_17886,N_17385,N_17262);
xor U17887 (N_17887,N_17505,N_17422);
nor U17888 (N_17888,N_17453,N_17318);
or U17889 (N_17889,N_17399,N_17450);
and U17890 (N_17890,N_17593,N_17225);
xnor U17891 (N_17891,N_17376,N_17215);
nor U17892 (N_17892,N_17477,N_17568);
xnor U17893 (N_17893,N_17251,N_17317);
nor U17894 (N_17894,N_17241,N_17532);
or U17895 (N_17895,N_17309,N_17352);
or U17896 (N_17896,N_17472,N_17410);
and U17897 (N_17897,N_17577,N_17254);
nand U17898 (N_17898,N_17233,N_17348);
xor U17899 (N_17899,N_17560,N_17517);
and U17900 (N_17900,N_17538,N_17384);
nand U17901 (N_17901,N_17518,N_17292);
nand U17902 (N_17902,N_17358,N_17449);
nor U17903 (N_17903,N_17297,N_17492);
nand U17904 (N_17904,N_17226,N_17365);
nor U17905 (N_17905,N_17380,N_17320);
nor U17906 (N_17906,N_17530,N_17502);
nand U17907 (N_17907,N_17460,N_17383);
or U17908 (N_17908,N_17335,N_17545);
xor U17909 (N_17909,N_17552,N_17468);
and U17910 (N_17910,N_17301,N_17594);
xor U17911 (N_17911,N_17415,N_17284);
nor U17912 (N_17912,N_17509,N_17477);
and U17913 (N_17913,N_17272,N_17366);
xor U17914 (N_17914,N_17333,N_17241);
nor U17915 (N_17915,N_17281,N_17417);
nor U17916 (N_17916,N_17340,N_17539);
and U17917 (N_17917,N_17447,N_17358);
nor U17918 (N_17918,N_17489,N_17201);
and U17919 (N_17919,N_17260,N_17483);
xor U17920 (N_17920,N_17420,N_17576);
or U17921 (N_17921,N_17390,N_17446);
or U17922 (N_17922,N_17502,N_17238);
or U17923 (N_17923,N_17598,N_17241);
nor U17924 (N_17924,N_17224,N_17429);
nand U17925 (N_17925,N_17324,N_17282);
nand U17926 (N_17926,N_17420,N_17353);
nand U17927 (N_17927,N_17368,N_17590);
xor U17928 (N_17928,N_17397,N_17291);
nand U17929 (N_17929,N_17325,N_17531);
xor U17930 (N_17930,N_17537,N_17513);
and U17931 (N_17931,N_17532,N_17436);
nor U17932 (N_17932,N_17528,N_17492);
or U17933 (N_17933,N_17310,N_17284);
and U17934 (N_17934,N_17574,N_17314);
nor U17935 (N_17935,N_17338,N_17347);
and U17936 (N_17936,N_17262,N_17366);
xor U17937 (N_17937,N_17458,N_17512);
nand U17938 (N_17938,N_17420,N_17375);
and U17939 (N_17939,N_17421,N_17295);
or U17940 (N_17940,N_17344,N_17459);
or U17941 (N_17941,N_17561,N_17349);
nand U17942 (N_17942,N_17494,N_17378);
or U17943 (N_17943,N_17351,N_17519);
and U17944 (N_17944,N_17311,N_17479);
nor U17945 (N_17945,N_17371,N_17459);
and U17946 (N_17946,N_17503,N_17499);
or U17947 (N_17947,N_17212,N_17409);
and U17948 (N_17948,N_17487,N_17253);
and U17949 (N_17949,N_17333,N_17321);
or U17950 (N_17950,N_17361,N_17535);
and U17951 (N_17951,N_17334,N_17447);
and U17952 (N_17952,N_17339,N_17430);
nand U17953 (N_17953,N_17475,N_17436);
and U17954 (N_17954,N_17258,N_17430);
xnor U17955 (N_17955,N_17254,N_17501);
nor U17956 (N_17956,N_17237,N_17585);
or U17957 (N_17957,N_17212,N_17565);
nand U17958 (N_17958,N_17451,N_17589);
nand U17959 (N_17959,N_17389,N_17550);
or U17960 (N_17960,N_17473,N_17284);
or U17961 (N_17961,N_17244,N_17446);
and U17962 (N_17962,N_17380,N_17565);
nand U17963 (N_17963,N_17251,N_17456);
nor U17964 (N_17964,N_17352,N_17353);
nand U17965 (N_17965,N_17281,N_17431);
nand U17966 (N_17966,N_17468,N_17434);
xor U17967 (N_17967,N_17425,N_17487);
nor U17968 (N_17968,N_17490,N_17575);
or U17969 (N_17969,N_17418,N_17490);
xor U17970 (N_17970,N_17444,N_17262);
and U17971 (N_17971,N_17215,N_17585);
xnor U17972 (N_17972,N_17589,N_17564);
nor U17973 (N_17973,N_17271,N_17518);
nand U17974 (N_17974,N_17286,N_17573);
nor U17975 (N_17975,N_17406,N_17334);
nand U17976 (N_17976,N_17323,N_17381);
and U17977 (N_17977,N_17249,N_17484);
nand U17978 (N_17978,N_17496,N_17217);
xnor U17979 (N_17979,N_17452,N_17407);
nand U17980 (N_17980,N_17583,N_17591);
or U17981 (N_17981,N_17347,N_17441);
xnor U17982 (N_17982,N_17545,N_17331);
and U17983 (N_17983,N_17363,N_17213);
and U17984 (N_17984,N_17317,N_17501);
nor U17985 (N_17985,N_17397,N_17334);
xnor U17986 (N_17986,N_17297,N_17248);
and U17987 (N_17987,N_17504,N_17541);
nor U17988 (N_17988,N_17520,N_17513);
nand U17989 (N_17989,N_17223,N_17432);
or U17990 (N_17990,N_17261,N_17414);
nor U17991 (N_17991,N_17436,N_17356);
xnor U17992 (N_17992,N_17343,N_17356);
xor U17993 (N_17993,N_17335,N_17221);
and U17994 (N_17994,N_17340,N_17344);
nand U17995 (N_17995,N_17398,N_17385);
or U17996 (N_17996,N_17566,N_17502);
and U17997 (N_17997,N_17263,N_17409);
xnor U17998 (N_17998,N_17458,N_17548);
or U17999 (N_17999,N_17226,N_17545);
or U18000 (N_18000,N_17643,N_17785);
or U18001 (N_18001,N_17759,N_17720);
xor U18002 (N_18002,N_17986,N_17747);
and U18003 (N_18003,N_17983,N_17931);
nand U18004 (N_18004,N_17802,N_17792);
nor U18005 (N_18005,N_17945,N_17949);
nor U18006 (N_18006,N_17903,N_17880);
nand U18007 (N_18007,N_17970,N_17781);
nor U18008 (N_18008,N_17887,N_17667);
xnor U18009 (N_18009,N_17700,N_17602);
and U18010 (N_18010,N_17961,N_17758);
nand U18011 (N_18011,N_17614,N_17803);
nand U18012 (N_18012,N_17672,N_17982);
xnor U18013 (N_18013,N_17648,N_17862);
or U18014 (N_18014,N_17975,N_17812);
nand U18015 (N_18015,N_17858,N_17901);
and U18016 (N_18016,N_17883,N_17628);
and U18017 (N_18017,N_17640,N_17838);
or U18018 (N_18018,N_17791,N_17991);
nand U18019 (N_18019,N_17874,N_17859);
xnor U18020 (N_18020,N_17852,N_17879);
and U18021 (N_18021,N_17656,N_17809);
xnor U18022 (N_18022,N_17936,N_17717);
xor U18023 (N_18023,N_17711,N_17616);
nor U18024 (N_18024,N_17670,N_17855);
xor U18025 (N_18025,N_17894,N_17610);
and U18026 (N_18026,N_17882,N_17703);
nor U18027 (N_18027,N_17822,N_17772);
nor U18028 (N_18028,N_17891,N_17689);
nor U18029 (N_18029,N_17981,N_17682);
xor U18030 (N_18030,N_17836,N_17861);
nand U18031 (N_18031,N_17749,N_17946);
xnor U18032 (N_18032,N_17736,N_17729);
nand U18033 (N_18033,N_17770,N_17743);
or U18034 (N_18034,N_17893,N_17666);
and U18035 (N_18035,N_17683,N_17625);
nand U18036 (N_18036,N_17696,N_17846);
nor U18037 (N_18037,N_17713,N_17827);
or U18038 (N_18038,N_17789,N_17715);
nor U18039 (N_18039,N_17635,N_17878);
nor U18040 (N_18040,N_17826,N_17871);
and U18041 (N_18041,N_17613,N_17662);
nand U18042 (N_18042,N_17764,N_17686);
or U18043 (N_18043,N_17940,N_17828);
xnor U18044 (N_18044,N_17820,N_17606);
or U18045 (N_18045,N_17771,N_17853);
or U18046 (N_18046,N_17765,N_17877);
nand U18047 (N_18047,N_17793,N_17751);
and U18048 (N_18048,N_17886,N_17950);
and U18049 (N_18049,N_17608,N_17676);
and U18050 (N_18050,N_17997,N_17933);
nand U18051 (N_18051,N_17671,N_17884);
nor U18052 (N_18052,N_17953,N_17787);
nand U18053 (N_18053,N_17994,N_17724);
and U18054 (N_18054,N_17889,N_17782);
nor U18055 (N_18055,N_17954,N_17956);
xor U18056 (N_18056,N_17609,N_17757);
and U18057 (N_18057,N_17753,N_17847);
nand U18058 (N_18058,N_17731,N_17929);
xnor U18059 (N_18059,N_17661,N_17763);
or U18060 (N_18060,N_17928,N_17664);
nand U18061 (N_18061,N_17626,N_17863);
nand U18062 (N_18062,N_17816,N_17677);
or U18063 (N_18063,N_17817,N_17815);
or U18064 (N_18064,N_17857,N_17864);
or U18065 (N_18065,N_17627,N_17721);
or U18066 (N_18066,N_17850,N_17669);
xor U18067 (N_18067,N_17649,N_17996);
and U18068 (N_18068,N_17779,N_17607);
nor U18069 (N_18069,N_17760,N_17632);
xor U18070 (N_18070,N_17800,N_17653);
nand U18071 (N_18071,N_17837,N_17995);
xor U18072 (N_18072,N_17819,N_17911);
and U18073 (N_18073,N_17848,N_17698);
nor U18074 (N_18074,N_17795,N_17748);
xnor U18075 (N_18075,N_17824,N_17835);
xnor U18076 (N_18076,N_17909,N_17900);
and U18077 (N_18077,N_17681,N_17907);
or U18078 (N_18078,N_17947,N_17993);
xor U18079 (N_18079,N_17639,N_17725);
and U18080 (N_18080,N_17774,N_17968);
nor U18081 (N_18081,N_17942,N_17839);
nand U18082 (N_18082,N_17741,N_17637);
or U18083 (N_18083,N_17896,N_17904);
or U18084 (N_18084,N_17926,N_17615);
and U18085 (N_18085,N_17892,N_17979);
nand U18086 (N_18086,N_17605,N_17801);
or U18087 (N_18087,N_17638,N_17612);
nor U18088 (N_18088,N_17844,N_17723);
xor U18089 (N_18089,N_17799,N_17823);
nand U18090 (N_18090,N_17733,N_17849);
nor U18091 (N_18091,N_17796,N_17964);
xor U18092 (N_18092,N_17930,N_17663);
nand U18093 (N_18093,N_17697,N_17987);
nand U18094 (N_18094,N_17642,N_17754);
or U18095 (N_18095,N_17808,N_17906);
nor U18096 (N_18096,N_17927,N_17619);
nor U18097 (N_18097,N_17657,N_17768);
nor U18098 (N_18098,N_17620,N_17644);
nand U18099 (N_18099,N_17756,N_17727);
xnor U18100 (N_18100,N_17914,N_17865);
or U18101 (N_18101,N_17888,N_17641);
xor U18102 (N_18102,N_17722,N_17962);
nand U18103 (N_18103,N_17692,N_17684);
or U18104 (N_18104,N_17941,N_17966);
xor U18105 (N_18105,N_17814,N_17634);
nand U18106 (N_18106,N_17650,N_17805);
xnor U18107 (N_18107,N_17984,N_17960);
nor U18108 (N_18108,N_17674,N_17840);
xor U18109 (N_18109,N_17989,N_17813);
or U18110 (N_18110,N_17750,N_17690);
nand U18111 (N_18111,N_17876,N_17999);
xnor U18112 (N_18112,N_17773,N_17948);
or U18113 (N_18113,N_17680,N_17745);
and U18114 (N_18114,N_17739,N_17617);
and U18115 (N_18115,N_17985,N_17973);
xor U18116 (N_18116,N_17631,N_17794);
nor U18117 (N_18117,N_17622,N_17709);
nand U18118 (N_18118,N_17937,N_17744);
nand U18119 (N_18119,N_17707,N_17730);
nand U18120 (N_18120,N_17710,N_17735);
nor U18121 (N_18121,N_17963,N_17691);
nand U18122 (N_18122,N_17762,N_17869);
nor U18123 (N_18123,N_17830,N_17959);
nand U18124 (N_18124,N_17766,N_17734);
nand U18125 (N_18125,N_17678,N_17786);
xnor U18126 (N_18126,N_17624,N_17842);
nor U18127 (N_18127,N_17923,N_17687);
nor U18128 (N_18128,N_17623,N_17921);
and U18129 (N_18129,N_17712,N_17977);
or U18130 (N_18130,N_17755,N_17732);
nand U18131 (N_18131,N_17647,N_17841);
and U18132 (N_18132,N_17737,N_17831);
or U18133 (N_18133,N_17988,N_17980);
or U18134 (N_18134,N_17645,N_17807);
nand U18135 (N_18135,N_17908,N_17881);
xor U18136 (N_18136,N_17851,N_17821);
and U18137 (N_18137,N_17829,N_17742);
nor U18138 (N_18138,N_17905,N_17897);
xnor U18139 (N_18139,N_17899,N_17965);
nor U18140 (N_18140,N_17600,N_17752);
and U18141 (N_18141,N_17912,N_17767);
nor U18142 (N_18142,N_17990,N_17798);
and U18143 (N_18143,N_17646,N_17957);
xnor U18144 (N_18144,N_17902,N_17740);
nor U18145 (N_18145,N_17706,N_17971);
xnor U18146 (N_18146,N_17958,N_17716);
and U18147 (N_18147,N_17969,N_17668);
nor U18148 (N_18148,N_17719,N_17636);
nor U18149 (N_18149,N_17685,N_17704);
xor U18150 (N_18150,N_17952,N_17976);
nor U18151 (N_18151,N_17967,N_17992);
and U18152 (N_18152,N_17804,N_17944);
or U18153 (N_18153,N_17665,N_17833);
or U18154 (N_18154,N_17784,N_17695);
xor U18155 (N_18155,N_17898,N_17699);
nor U18156 (N_18156,N_17955,N_17916);
nand U18157 (N_18157,N_17834,N_17769);
and U18158 (N_18158,N_17675,N_17630);
nand U18159 (N_18159,N_17780,N_17705);
and U18160 (N_18160,N_17806,N_17843);
and U18161 (N_18161,N_17660,N_17920);
xor U18162 (N_18162,N_17790,N_17845);
nand U18163 (N_18163,N_17726,N_17694);
nand U18164 (N_18164,N_17693,N_17974);
nor U18165 (N_18165,N_17797,N_17673);
xor U18166 (N_18166,N_17978,N_17810);
and U18167 (N_18167,N_17618,N_17924);
or U18168 (N_18168,N_17603,N_17688);
or U18169 (N_18169,N_17856,N_17832);
nor U18170 (N_18170,N_17621,N_17708);
and U18171 (N_18171,N_17890,N_17825);
or U18172 (N_18172,N_17761,N_17658);
xnor U18173 (N_18173,N_17746,N_17652);
xnor U18174 (N_18174,N_17917,N_17918);
nor U18175 (N_18175,N_17860,N_17866);
and U18176 (N_18176,N_17932,N_17910);
xor U18177 (N_18177,N_17788,N_17951);
nor U18178 (N_18178,N_17601,N_17728);
nand U18179 (N_18179,N_17654,N_17783);
or U18180 (N_18180,N_17611,N_17629);
and U18181 (N_18181,N_17872,N_17939);
and U18182 (N_18182,N_17913,N_17811);
or U18183 (N_18183,N_17778,N_17738);
and U18184 (N_18184,N_17818,N_17873);
and U18185 (N_18185,N_17633,N_17870);
and U18186 (N_18186,N_17885,N_17925);
and U18187 (N_18187,N_17679,N_17659);
and U18188 (N_18188,N_17922,N_17972);
nor U18189 (N_18189,N_17775,N_17868);
nand U18190 (N_18190,N_17998,N_17714);
and U18191 (N_18191,N_17604,N_17938);
or U18192 (N_18192,N_17702,N_17895);
or U18193 (N_18193,N_17934,N_17777);
or U18194 (N_18194,N_17943,N_17854);
and U18195 (N_18195,N_17867,N_17655);
and U18196 (N_18196,N_17776,N_17935);
nor U18197 (N_18197,N_17718,N_17701);
and U18198 (N_18198,N_17651,N_17915);
and U18199 (N_18199,N_17875,N_17919);
or U18200 (N_18200,N_17752,N_17868);
or U18201 (N_18201,N_17657,N_17807);
and U18202 (N_18202,N_17789,N_17666);
or U18203 (N_18203,N_17750,N_17730);
and U18204 (N_18204,N_17922,N_17964);
and U18205 (N_18205,N_17881,N_17809);
nand U18206 (N_18206,N_17762,N_17806);
nand U18207 (N_18207,N_17637,N_17859);
nand U18208 (N_18208,N_17979,N_17941);
and U18209 (N_18209,N_17816,N_17809);
xnor U18210 (N_18210,N_17690,N_17840);
or U18211 (N_18211,N_17734,N_17791);
or U18212 (N_18212,N_17672,N_17622);
xnor U18213 (N_18213,N_17985,N_17626);
and U18214 (N_18214,N_17648,N_17971);
or U18215 (N_18215,N_17672,N_17704);
nand U18216 (N_18216,N_17971,N_17877);
nand U18217 (N_18217,N_17750,N_17885);
or U18218 (N_18218,N_17850,N_17801);
nor U18219 (N_18219,N_17701,N_17625);
nand U18220 (N_18220,N_17817,N_17869);
xnor U18221 (N_18221,N_17745,N_17751);
nor U18222 (N_18222,N_17935,N_17726);
xor U18223 (N_18223,N_17758,N_17765);
and U18224 (N_18224,N_17932,N_17934);
nand U18225 (N_18225,N_17654,N_17623);
nand U18226 (N_18226,N_17691,N_17836);
nor U18227 (N_18227,N_17985,N_17646);
or U18228 (N_18228,N_17908,N_17804);
or U18229 (N_18229,N_17894,N_17674);
xor U18230 (N_18230,N_17779,N_17863);
or U18231 (N_18231,N_17607,N_17894);
or U18232 (N_18232,N_17947,N_17909);
and U18233 (N_18233,N_17901,N_17926);
and U18234 (N_18234,N_17708,N_17918);
xor U18235 (N_18235,N_17650,N_17637);
or U18236 (N_18236,N_17755,N_17939);
xor U18237 (N_18237,N_17782,N_17894);
or U18238 (N_18238,N_17661,N_17932);
xor U18239 (N_18239,N_17622,N_17798);
nand U18240 (N_18240,N_17782,N_17999);
nor U18241 (N_18241,N_17630,N_17609);
nand U18242 (N_18242,N_17988,N_17642);
and U18243 (N_18243,N_17651,N_17831);
nor U18244 (N_18244,N_17693,N_17935);
xnor U18245 (N_18245,N_17721,N_17942);
and U18246 (N_18246,N_17831,N_17720);
nand U18247 (N_18247,N_17666,N_17754);
nor U18248 (N_18248,N_17698,N_17808);
nand U18249 (N_18249,N_17743,N_17687);
xor U18250 (N_18250,N_17744,N_17707);
nand U18251 (N_18251,N_17699,N_17892);
or U18252 (N_18252,N_17667,N_17673);
xor U18253 (N_18253,N_17778,N_17623);
nand U18254 (N_18254,N_17942,N_17736);
and U18255 (N_18255,N_17743,N_17846);
nor U18256 (N_18256,N_17610,N_17993);
nor U18257 (N_18257,N_17781,N_17946);
or U18258 (N_18258,N_17800,N_17903);
nand U18259 (N_18259,N_17852,N_17933);
xor U18260 (N_18260,N_17859,N_17987);
and U18261 (N_18261,N_17751,N_17825);
and U18262 (N_18262,N_17973,N_17939);
nand U18263 (N_18263,N_17985,N_17950);
or U18264 (N_18264,N_17683,N_17639);
nand U18265 (N_18265,N_17786,N_17620);
or U18266 (N_18266,N_17874,N_17601);
nand U18267 (N_18267,N_17991,N_17674);
xnor U18268 (N_18268,N_17761,N_17893);
or U18269 (N_18269,N_17773,N_17626);
nor U18270 (N_18270,N_17647,N_17919);
nand U18271 (N_18271,N_17959,N_17847);
xor U18272 (N_18272,N_17796,N_17770);
xor U18273 (N_18273,N_17617,N_17870);
nor U18274 (N_18274,N_17749,N_17861);
and U18275 (N_18275,N_17938,N_17804);
and U18276 (N_18276,N_17871,N_17944);
nor U18277 (N_18277,N_17959,N_17624);
and U18278 (N_18278,N_17992,N_17610);
and U18279 (N_18279,N_17976,N_17914);
nand U18280 (N_18280,N_17896,N_17825);
nand U18281 (N_18281,N_17653,N_17737);
nand U18282 (N_18282,N_17647,N_17847);
nand U18283 (N_18283,N_17937,N_17815);
or U18284 (N_18284,N_17645,N_17986);
xnor U18285 (N_18285,N_17873,N_17682);
nor U18286 (N_18286,N_17894,N_17955);
and U18287 (N_18287,N_17637,N_17988);
nand U18288 (N_18288,N_17894,N_17864);
nor U18289 (N_18289,N_17902,N_17666);
and U18290 (N_18290,N_17961,N_17764);
nand U18291 (N_18291,N_17622,N_17602);
or U18292 (N_18292,N_17868,N_17642);
nor U18293 (N_18293,N_17644,N_17782);
xnor U18294 (N_18294,N_17682,N_17658);
nand U18295 (N_18295,N_17816,N_17985);
nor U18296 (N_18296,N_17616,N_17871);
or U18297 (N_18297,N_17669,N_17648);
nand U18298 (N_18298,N_17697,N_17994);
nand U18299 (N_18299,N_17754,N_17942);
and U18300 (N_18300,N_17787,N_17776);
nand U18301 (N_18301,N_17646,N_17927);
and U18302 (N_18302,N_17748,N_17733);
nor U18303 (N_18303,N_17771,N_17641);
nand U18304 (N_18304,N_17795,N_17777);
nand U18305 (N_18305,N_17821,N_17966);
xnor U18306 (N_18306,N_17685,N_17673);
xor U18307 (N_18307,N_17990,N_17962);
xor U18308 (N_18308,N_17776,N_17959);
or U18309 (N_18309,N_17632,N_17693);
xor U18310 (N_18310,N_17634,N_17978);
nor U18311 (N_18311,N_17857,N_17674);
or U18312 (N_18312,N_17715,N_17779);
xnor U18313 (N_18313,N_17922,N_17898);
nand U18314 (N_18314,N_17731,N_17756);
xnor U18315 (N_18315,N_17871,N_17639);
nand U18316 (N_18316,N_17647,N_17958);
or U18317 (N_18317,N_17726,N_17665);
and U18318 (N_18318,N_17800,N_17723);
nor U18319 (N_18319,N_17824,N_17879);
nand U18320 (N_18320,N_17668,N_17646);
and U18321 (N_18321,N_17996,N_17953);
nor U18322 (N_18322,N_17919,N_17796);
xor U18323 (N_18323,N_17634,N_17604);
nor U18324 (N_18324,N_17983,N_17875);
xnor U18325 (N_18325,N_17873,N_17974);
nand U18326 (N_18326,N_17981,N_17675);
nor U18327 (N_18327,N_17920,N_17670);
xnor U18328 (N_18328,N_17886,N_17708);
or U18329 (N_18329,N_17936,N_17697);
nand U18330 (N_18330,N_17876,N_17913);
or U18331 (N_18331,N_17711,N_17995);
nand U18332 (N_18332,N_17913,N_17726);
and U18333 (N_18333,N_17862,N_17979);
and U18334 (N_18334,N_17897,N_17606);
xor U18335 (N_18335,N_17923,N_17646);
and U18336 (N_18336,N_17834,N_17611);
and U18337 (N_18337,N_17874,N_17706);
nor U18338 (N_18338,N_17865,N_17786);
and U18339 (N_18339,N_17708,N_17815);
nand U18340 (N_18340,N_17650,N_17737);
xnor U18341 (N_18341,N_17614,N_17753);
nand U18342 (N_18342,N_17743,N_17933);
or U18343 (N_18343,N_17746,N_17872);
and U18344 (N_18344,N_17961,N_17815);
or U18345 (N_18345,N_17614,N_17711);
nor U18346 (N_18346,N_17893,N_17738);
xor U18347 (N_18347,N_17888,N_17798);
or U18348 (N_18348,N_17836,N_17965);
xor U18349 (N_18349,N_17610,N_17927);
or U18350 (N_18350,N_17744,N_17963);
xnor U18351 (N_18351,N_17707,N_17883);
xor U18352 (N_18352,N_17741,N_17849);
or U18353 (N_18353,N_17990,N_17790);
nor U18354 (N_18354,N_17628,N_17697);
nor U18355 (N_18355,N_17917,N_17672);
nor U18356 (N_18356,N_17965,N_17873);
and U18357 (N_18357,N_17629,N_17637);
xor U18358 (N_18358,N_17985,N_17994);
nor U18359 (N_18359,N_17931,N_17922);
nor U18360 (N_18360,N_17902,N_17865);
and U18361 (N_18361,N_17729,N_17889);
and U18362 (N_18362,N_17805,N_17678);
and U18363 (N_18363,N_17819,N_17756);
nor U18364 (N_18364,N_17980,N_17973);
xnor U18365 (N_18365,N_17959,N_17867);
xnor U18366 (N_18366,N_17682,N_17753);
nand U18367 (N_18367,N_17624,N_17712);
nor U18368 (N_18368,N_17725,N_17856);
or U18369 (N_18369,N_17901,N_17827);
and U18370 (N_18370,N_17700,N_17905);
or U18371 (N_18371,N_17847,N_17744);
and U18372 (N_18372,N_17840,N_17647);
and U18373 (N_18373,N_17999,N_17922);
nor U18374 (N_18374,N_17879,N_17665);
and U18375 (N_18375,N_17740,N_17862);
xnor U18376 (N_18376,N_17651,N_17813);
xor U18377 (N_18377,N_17965,N_17855);
or U18378 (N_18378,N_17872,N_17695);
nor U18379 (N_18379,N_17689,N_17962);
xnor U18380 (N_18380,N_17751,N_17934);
and U18381 (N_18381,N_17897,N_17972);
nor U18382 (N_18382,N_17850,N_17963);
nor U18383 (N_18383,N_17783,N_17924);
nor U18384 (N_18384,N_17655,N_17988);
or U18385 (N_18385,N_17623,N_17773);
nand U18386 (N_18386,N_17877,N_17974);
xnor U18387 (N_18387,N_17777,N_17979);
xor U18388 (N_18388,N_17771,N_17718);
nor U18389 (N_18389,N_17670,N_17863);
nor U18390 (N_18390,N_17896,N_17782);
or U18391 (N_18391,N_17710,N_17929);
or U18392 (N_18392,N_17657,N_17843);
or U18393 (N_18393,N_17966,N_17731);
or U18394 (N_18394,N_17810,N_17854);
nand U18395 (N_18395,N_17606,N_17732);
nor U18396 (N_18396,N_17873,N_17868);
nor U18397 (N_18397,N_17736,N_17969);
and U18398 (N_18398,N_17782,N_17852);
nand U18399 (N_18399,N_17850,N_17712);
nor U18400 (N_18400,N_18218,N_18225);
xor U18401 (N_18401,N_18228,N_18231);
nor U18402 (N_18402,N_18142,N_18196);
nor U18403 (N_18403,N_18131,N_18141);
or U18404 (N_18404,N_18011,N_18184);
or U18405 (N_18405,N_18329,N_18073);
nand U18406 (N_18406,N_18034,N_18028);
xnor U18407 (N_18407,N_18064,N_18311);
xnor U18408 (N_18408,N_18236,N_18113);
xor U18409 (N_18409,N_18327,N_18058);
or U18410 (N_18410,N_18166,N_18177);
or U18411 (N_18411,N_18182,N_18092);
nor U18412 (N_18412,N_18180,N_18193);
xnor U18413 (N_18413,N_18385,N_18285);
or U18414 (N_18414,N_18122,N_18148);
and U18415 (N_18415,N_18264,N_18276);
nand U18416 (N_18416,N_18227,N_18202);
nor U18417 (N_18417,N_18192,N_18077);
or U18418 (N_18418,N_18002,N_18300);
nor U18419 (N_18419,N_18232,N_18140);
and U18420 (N_18420,N_18353,N_18293);
nor U18421 (N_18421,N_18207,N_18395);
nor U18422 (N_18422,N_18208,N_18079);
xor U18423 (N_18423,N_18169,N_18033);
or U18424 (N_18424,N_18319,N_18025);
xnor U18425 (N_18425,N_18154,N_18265);
nand U18426 (N_18426,N_18351,N_18151);
and U18427 (N_18427,N_18239,N_18200);
nand U18428 (N_18428,N_18054,N_18022);
xnor U18429 (N_18429,N_18100,N_18050);
nor U18430 (N_18430,N_18240,N_18349);
nand U18431 (N_18431,N_18355,N_18290);
nand U18432 (N_18432,N_18284,N_18063);
nand U18433 (N_18433,N_18283,N_18376);
or U18434 (N_18434,N_18205,N_18174);
and U18435 (N_18435,N_18134,N_18031);
nor U18436 (N_18436,N_18155,N_18282);
xnor U18437 (N_18437,N_18065,N_18335);
and U18438 (N_18438,N_18137,N_18060);
nand U18439 (N_18439,N_18072,N_18186);
and U18440 (N_18440,N_18374,N_18326);
or U18441 (N_18441,N_18315,N_18248);
or U18442 (N_18442,N_18256,N_18222);
or U18443 (N_18443,N_18348,N_18216);
nand U18444 (N_18444,N_18171,N_18107);
or U18445 (N_18445,N_18294,N_18263);
nand U18446 (N_18446,N_18378,N_18023);
and U18447 (N_18447,N_18246,N_18001);
nor U18448 (N_18448,N_18295,N_18244);
nand U18449 (N_18449,N_18118,N_18210);
and U18450 (N_18450,N_18270,N_18241);
xnor U18451 (N_18451,N_18388,N_18088);
xor U18452 (N_18452,N_18046,N_18379);
xor U18453 (N_18453,N_18078,N_18350);
or U18454 (N_18454,N_18359,N_18255);
nor U18455 (N_18455,N_18303,N_18217);
nor U18456 (N_18456,N_18391,N_18150);
and U18457 (N_18457,N_18167,N_18066);
xnor U18458 (N_18458,N_18213,N_18048);
nor U18459 (N_18459,N_18106,N_18039);
and U18460 (N_18460,N_18322,N_18009);
or U18461 (N_18461,N_18111,N_18070);
xor U18462 (N_18462,N_18115,N_18384);
and U18463 (N_18463,N_18051,N_18252);
xor U18464 (N_18464,N_18361,N_18334);
xnor U18465 (N_18465,N_18056,N_18108);
nand U18466 (N_18466,N_18116,N_18143);
nand U18467 (N_18467,N_18021,N_18105);
and U18468 (N_18468,N_18268,N_18067);
nor U18469 (N_18469,N_18027,N_18052);
or U18470 (N_18470,N_18185,N_18080);
xnor U18471 (N_18471,N_18187,N_18242);
nor U18472 (N_18472,N_18237,N_18250);
xor U18473 (N_18473,N_18132,N_18269);
and U18474 (N_18474,N_18018,N_18392);
nor U18475 (N_18475,N_18110,N_18147);
nand U18476 (N_18476,N_18189,N_18203);
nand U18477 (N_18477,N_18215,N_18238);
nand U18478 (N_18478,N_18342,N_18325);
nand U18479 (N_18479,N_18211,N_18386);
xor U18480 (N_18480,N_18099,N_18121);
xnor U18481 (N_18481,N_18119,N_18197);
nor U18482 (N_18482,N_18053,N_18380);
nand U18483 (N_18483,N_18226,N_18090);
and U18484 (N_18484,N_18133,N_18006);
nand U18485 (N_18485,N_18059,N_18398);
xnor U18486 (N_18486,N_18362,N_18040);
or U18487 (N_18487,N_18013,N_18096);
and U18488 (N_18488,N_18135,N_18313);
nand U18489 (N_18489,N_18199,N_18370);
and U18490 (N_18490,N_18375,N_18396);
and U18491 (N_18491,N_18043,N_18206);
and U18492 (N_18492,N_18162,N_18343);
nor U18493 (N_18493,N_18347,N_18082);
nor U18494 (N_18494,N_18083,N_18038);
xnor U18495 (N_18495,N_18383,N_18145);
nand U18496 (N_18496,N_18047,N_18259);
nand U18497 (N_18497,N_18320,N_18209);
nor U18498 (N_18498,N_18340,N_18288);
and U18499 (N_18499,N_18287,N_18175);
and U18500 (N_18500,N_18117,N_18165);
xor U18501 (N_18501,N_18109,N_18057);
or U18502 (N_18502,N_18258,N_18041);
or U18503 (N_18503,N_18330,N_18298);
and U18504 (N_18504,N_18366,N_18097);
nor U18505 (N_18505,N_18306,N_18005);
nor U18506 (N_18506,N_18178,N_18221);
xnor U18507 (N_18507,N_18345,N_18045);
and U18508 (N_18508,N_18091,N_18032);
nor U18509 (N_18509,N_18084,N_18317);
nand U18510 (N_18510,N_18243,N_18318);
nor U18511 (N_18511,N_18170,N_18289);
nand U18512 (N_18512,N_18249,N_18247);
and U18513 (N_18513,N_18003,N_18044);
xor U18514 (N_18514,N_18389,N_18332);
and U18515 (N_18515,N_18219,N_18007);
xor U18516 (N_18516,N_18161,N_18069);
and U18517 (N_18517,N_18149,N_18278);
nand U18518 (N_18518,N_18194,N_18297);
nor U18519 (N_18519,N_18030,N_18382);
nand U18520 (N_18520,N_18312,N_18234);
or U18521 (N_18521,N_18172,N_18017);
xnor U18522 (N_18522,N_18144,N_18314);
xnor U18523 (N_18523,N_18214,N_18124);
xor U18524 (N_18524,N_18333,N_18302);
nand U18525 (N_18525,N_18015,N_18020);
xor U18526 (N_18526,N_18128,N_18114);
nand U18527 (N_18527,N_18341,N_18160);
and U18528 (N_18528,N_18338,N_18014);
or U18529 (N_18529,N_18371,N_18062);
xnor U18530 (N_18530,N_18230,N_18266);
or U18531 (N_18531,N_18000,N_18394);
xnor U18532 (N_18532,N_18273,N_18008);
xnor U18533 (N_18533,N_18168,N_18220);
nand U18534 (N_18534,N_18120,N_18377);
or U18535 (N_18535,N_18254,N_18195);
and U18536 (N_18536,N_18201,N_18123);
nand U18537 (N_18537,N_18095,N_18304);
nor U18538 (N_18538,N_18159,N_18127);
and U18539 (N_18539,N_18235,N_18309);
nor U18540 (N_18540,N_18024,N_18233);
nand U18541 (N_18541,N_18271,N_18071);
or U18542 (N_18542,N_18272,N_18036);
or U18543 (N_18543,N_18364,N_18204);
or U18544 (N_18544,N_18397,N_18093);
and U18545 (N_18545,N_18344,N_18373);
or U18546 (N_18546,N_18112,N_18365);
xnor U18547 (N_18547,N_18081,N_18004);
nor U18548 (N_18548,N_18223,N_18352);
xnor U18549 (N_18549,N_18367,N_18104);
or U18550 (N_18550,N_18354,N_18358);
nor U18551 (N_18551,N_18224,N_18068);
or U18552 (N_18552,N_18360,N_18176);
and U18553 (N_18553,N_18191,N_18245);
and U18554 (N_18554,N_18183,N_18163);
nand U18555 (N_18555,N_18010,N_18262);
nand U18556 (N_18556,N_18087,N_18156);
xor U18557 (N_18557,N_18356,N_18103);
and U18558 (N_18558,N_18037,N_18153);
xnor U18559 (N_18559,N_18049,N_18130);
and U18560 (N_18560,N_18181,N_18126);
nor U18561 (N_18561,N_18055,N_18381);
or U18562 (N_18562,N_18261,N_18173);
nand U18563 (N_18563,N_18212,N_18363);
nor U18564 (N_18564,N_18146,N_18296);
nor U18565 (N_18565,N_18399,N_18152);
nand U18566 (N_18566,N_18337,N_18089);
or U18567 (N_18567,N_18321,N_18035);
or U18568 (N_18568,N_18251,N_18308);
xnor U18569 (N_18569,N_18257,N_18129);
nor U18570 (N_18570,N_18102,N_18042);
and U18571 (N_18571,N_18291,N_18292);
and U18572 (N_18572,N_18286,N_18339);
or U18573 (N_18573,N_18281,N_18346);
nor U18574 (N_18574,N_18336,N_18164);
and U18575 (N_18575,N_18260,N_18158);
or U18576 (N_18576,N_18368,N_18138);
or U18577 (N_18577,N_18012,N_18026);
or U18578 (N_18578,N_18075,N_18393);
and U18579 (N_18579,N_18074,N_18016);
nor U18580 (N_18580,N_18307,N_18328);
nor U18581 (N_18581,N_18274,N_18253);
nand U18582 (N_18582,N_18190,N_18029);
xor U18583 (N_18583,N_18198,N_18101);
or U18584 (N_18584,N_18019,N_18188);
or U18585 (N_18585,N_18267,N_18136);
or U18586 (N_18586,N_18301,N_18316);
or U18587 (N_18587,N_18061,N_18157);
and U18588 (N_18588,N_18139,N_18085);
xnor U18589 (N_18589,N_18390,N_18275);
and U18590 (N_18590,N_18279,N_18098);
or U18591 (N_18591,N_18387,N_18086);
nand U18592 (N_18592,N_18125,N_18094);
or U18593 (N_18593,N_18299,N_18076);
nor U18594 (N_18594,N_18229,N_18323);
nand U18595 (N_18595,N_18372,N_18280);
xor U18596 (N_18596,N_18324,N_18179);
nand U18597 (N_18597,N_18369,N_18331);
nor U18598 (N_18598,N_18277,N_18357);
or U18599 (N_18599,N_18310,N_18305);
nand U18600 (N_18600,N_18021,N_18318);
nor U18601 (N_18601,N_18097,N_18137);
and U18602 (N_18602,N_18225,N_18114);
nand U18603 (N_18603,N_18364,N_18231);
nor U18604 (N_18604,N_18195,N_18001);
or U18605 (N_18605,N_18109,N_18105);
and U18606 (N_18606,N_18332,N_18307);
xnor U18607 (N_18607,N_18298,N_18189);
xor U18608 (N_18608,N_18375,N_18057);
and U18609 (N_18609,N_18228,N_18201);
or U18610 (N_18610,N_18097,N_18131);
xor U18611 (N_18611,N_18096,N_18360);
nand U18612 (N_18612,N_18214,N_18051);
nor U18613 (N_18613,N_18090,N_18373);
or U18614 (N_18614,N_18316,N_18079);
or U18615 (N_18615,N_18164,N_18123);
xnor U18616 (N_18616,N_18276,N_18243);
and U18617 (N_18617,N_18289,N_18250);
or U18618 (N_18618,N_18074,N_18172);
and U18619 (N_18619,N_18321,N_18164);
nand U18620 (N_18620,N_18291,N_18344);
xnor U18621 (N_18621,N_18339,N_18328);
or U18622 (N_18622,N_18335,N_18022);
nand U18623 (N_18623,N_18107,N_18143);
xor U18624 (N_18624,N_18068,N_18175);
xnor U18625 (N_18625,N_18130,N_18199);
nand U18626 (N_18626,N_18315,N_18137);
or U18627 (N_18627,N_18071,N_18202);
nor U18628 (N_18628,N_18119,N_18329);
nor U18629 (N_18629,N_18106,N_18159);
nand U18630 (N_18630,N_18148,N_18357);
and U18631 (N_18631,N_18320,N_18356);
xor U18632 (N_18632,N_18192,N_18175);
nor U18633 (N_18633,N_18025,N_18348);
or U18634 (N_18634,N_18269,N_18172);
or U18635 (N_18635,N_18182,N_18141);
or U18636 (N_18636,N_18001,N_18292);
xor U18637 (N_18637,N_18232,N_18359);
and U18638 (N_18638,N_18032,N_18126);
or U18639 (N_18639,N_18197,N_18250);
nor U18640 (N_18640,N_18261,N_18262);
nand U18641 (N_18641,N_18034,N_18096);
nand U18642 (N_18642,N_18244,N_18261);
and U18643 (N_18643,N_18025,N_18041);
xnor U18644 (N_18644,N_18096,N_18113);
nor U18645 (N_18645,N_18302,N_18298);
nand U18646 (N_18646,N_18189,N_18113);
xor U18647 (N_18647,N_18105,N_18281);
xor U18648 (N_18648,N_18105,N_18108);
xnor U18649 (N_18649,N_18104,N_18332);
and U18650 (N_18650,N_18007,N_18033);
xor U18651 (N_18651,N_18048,N_18275);
or U18652 (N_18652,N_18126,N_18104);
nor U18653 (N_18653,N_18201,N_18136);
nor U18654 (N_18654,N_18231,N_18361);
and U18655 (N_18655,N_18126,N_18220);
nand U18656 (N_18656,N_18356,N_18285);
and U18657 (N_18657,N_18343,N_18381);
nor U18658 (N_18658,N_18367,N_18264);
or U18659 (N_18659,N_18107,N_18220);
or U18660 (N_18660,N_18023,N_18066);
nor U18661 (N_18661,N_18017,N_18344);
xnor U18662 (N_18662,N_18206,N_18030);
xor U18663 (N_18663,N_18153,N_18157);
xnor U18664 (N_18664,N_18264,N_18013);
nor U18665 (N_18665,N_18348,N_18341);
nor U18666 (N_18666,N_18188,N_18161);
nor U18667 (N_18667,N_18337,N_18059);
or U18668 (N_18668,N_18153,N_18349);
nand U18669 (N_18669,N_18369,N_18384);
nor U18670 (N_18670,N_18297,N_18267);
or U18671 (N_18671,N_18183,N_18016);
nor U18672 (N_18672,N_18211,N_18354);
and U18673 (N_18673,N_18241,N_18348);
or U18674 (N_18674,N_18109,N_18382);
and U18675 (N_18675,N_18181,N_18262);
and U18676 (N_18676,N_18380,N_18209);
nand U18677 (N_18677,N_18317,N_18174);
xnor U18678 (N_18678,N_18372,N_18317);
nand U18679 (N_18679,N_18188,N_18202);
nand U18680 (N_18680,N_18158,N_18095);
nand U18681 (N_18681,N_18064,N_18270);
or U18682 (N_18682,N_18089,N_18141);
and U18683 (N_18683,N_18329,N_18010);
xnor U18684 (N_18684,N_18046,N_18361);
or U18685 (N_18685,N_18056,N_18054);
or U18686 (N_18686,N_18312,N_18119);
xor U18687 (N_18687,N_18276,N_18037);
and U18688 (N_18688,N_18009,N_18347);
or U18689 (N_18689,N_18231,N_18305);
and U18690 (N_18690,N_18247,N_18098);
or U18691 (N_18691,N_18079,N_18108);
xnor U18692 (N_18692,N_18146,N_18224);
xnor U18693 (N_18693,N_18318,N_18291);
xnor U18694 (N_18694,N_18195,N_18143);
nor U18695 (N_18695,N_18138,N_18396);
nand U18696 (N_18696,N_18310,N_18136);
and U18697 (N_18697,N_18155,N_18059);
xnor U18698 (N_18698,N_18110,N_18254);
and U18699 (N_18699,N_18052,N_18197);
nor U18700 (N_18700,N_18073,N_18296);
xnor U18701 (N_18701,N_18094,N_18234);
nand U18702 (N_18702,N_18080,N_18161);
nand U18703 (N_18703,N_18312,N_18340);
or U18704 (N_18704,N_18210,N_18169);
or U18705 (N_18705,N_18240,N_18041);
xor U18706 (N_18706,N_18034,N_18245);
nand U18707 (N_18707,N_18397,N_18228);
xor U18708 (N_18708,N_18069,N_18016);
nor U18709 (N_18709,N_18189,N_18146);
nand U18710 (N_18710,N_18039,N_18251);
xor U18711 (N_18711,N_18340,N_18201);
xor U18712 (N_18712,N_18113,N_18074);
and U18713 (N_18713,N_18341,N_18136);
nor U18714 (N_18714,N_18067,N_18076);
and U18715 (N_18715,N_18190,N_18257);
and U18716 (N_18716,N_18217,N_18368);
or U18717 (N_18717,N_18056,N_18088);
nand U18718 (N_18718,N_18058,N_18362);
and U18719 (N_18719,N_18036,N_18055);
and U18720 (N_18720,N_18271,N_18011);
nor U18721 (N_18721,N_18267,N_18380);
nor U18722 (N_18722,N_18390,N_18213);
xor U18723 (N_18723,N_18234,N_18113);
nand U18724 (N_18724,N_18309,N_18374);
and U18725 (N_18725,N_18268,N_18189);
or U18726 (N_18726,N_18055,N_18122);
or U18727 (N_18727,N_18212,N_18273);
nand U18728 (N_18728,N_18218,N_18033);
and U18729 (N_18729,N_18188,N_18268);
nand U18730 (N_18730,N_18291,N_18398);
and U18731 (N_18731,N_18208,N_18230);
nor U18732 (N_18732,N_18330,N_18135);
and U18733 (N_18733,N_18190,N_18201);
nor U18734 (N_18734,N_18260,N_18263);
and U18735 (N_18735,N_18186,N_18178);
or U18736 (N_18736,N_18152,N_18245);
or U18737 (N_18737,N_18221,N_18369);
xor U18738 (N_18738,N_18062,N_18119);
or U18739 (N_18739,N_18258,N_18392);
nor U18740 (N_18740,N_18116,N_18075);
nand U18741 (N_18741,N_18043,N_18331);
nor U18742 (N_18742,N_18311,N_18206);
or U18743 (N_18743,N_18244,N_18070);
nor U18744 (N_18744,N_18399,N_18053);
or U18745 (N_18745,N_18360,N_18194);
nor U18746 (N_18746,N_18166,N_18209);
and U18747 (N_18747,N_18143,N_18086);
and U18748 (N_18748,N_18336,N_18346);
nand U18749 (N_18749,N_18160,N_18095);
or U18750 (N_18750,N_18335,N_18371);
or U18751 (N_18751,N_18167,N_18044);
nand U18752 (N_18752,N_18307,N_18116);
xor U18753 (N_18753,N_18269,N_18115);
and U18754 (N_18754,N_18023,N_18256);
nand U18755 (N_18755,N_18243,N_18135);
xor U18756 (N_18756,N_18288,N_18337);
or U18757 (N_18757,N_18019,N_18392);
or U18758 (N_18758,N_18060,N_18366);
xnor U18759 (N_18759,N_18168,N_18315);
and U18760 (N_18760,N_18078,N_18386);
or U18761 (N_18761,N_18031,N_18317);
xor U18762 (N_18762,N_18214,N_18022);
or U18763 (N_18763,N_18264,N_18244);
and U18764 (N_18764,N_18113,N_18393);
xnor U18765 (N_18765,N_18096,N_18078);
or U18766 (N_18766,N_18324,N_18112);
and U18767 (N_18767,N_18250,N_18297);
nand U18768 (N_18768,N_18019,N_18359);
nand U18769 (N_18769,N_18291,N_18116);
nand U18770 (N_18770,N_18242,N_18118);
or U18771 (N_18771,N_18396,N_18149);
nand U18772 (N_18772,N_18271,N_18046);
and U18773 (N_18773,N_18144,N_18152);
or U18774 (N_18774,N_18037,N_18118);
nor U18775 (N_18775,N_18197,N_18303);
or U18776 (N_18776,N_18380,N_18365);
xnor U18777 (N_18777,N_18032,N_18339);
xnor U18778 (N_18778,N_18261,N_18366);
or U18779 (N_18779,N_18048,N_18247);
or U18780 (N_18780,N_18299,N_18310);
or U18781 (N_18781,N_18115,N_18381);
nor U18782 (N_18782,N_18218,N_18238);
and U18783 (N_18783,N_18230,N_18180);
nor U18784 (N_18784,N_18155,N_18392);
nand U18785 (N_18785,N_18196,N_18270);
nand U18786 (N_18786,N_18006,N_18321);
and U18787 (N_18787,N_18037,N_18232);
and U18788 (N_18788,N_18234,N_18011);
xor U18789 (N_18789,N_18055,N_18148);
nor U18790 (N_18790,N_18169,N_18146);
nor U18791 (N_18791,N_18059,N_18007);
nor U18792 (N_18792,N_18194,N_18142);
nor U18793 (N_18793,N_18018,N_18219);
and U18794 (N_18794,N_18279,N_18276);
nor U18795 (N_18795,N_18232,N_18223);
nand U18796 (N_18796,N_18231,N_18130);
xor U18797 (N_18797,N_18079,N_18137);
or U18798 (N_18798,N_18015,N_18191);
and U18799 (N_18799,N_18136,N_18142);
nand U18800 (N_18800,N_18447,N_18763);
or U18801 (N_18801,N_18726,N_18436);
nor U18802 (N_18802,N_18737,N_18516);
nor U18803 (N_18803,N_18733,N_18739);
xor U18804 (N_18804,N_18607,N_18478);
xnor U18805 (N_18805,N_18654,N_18753);
nor U18806 (N_18806,N_18774,N_18765);
xor U18807 (N_18807,N_18466,N_18522);
or U18808 (N_18808,N_18464,N_18661);
and U18809 (N_18809,N_18676,N_18598);
nand U18810 (N_18810,N_18677,N_18584);
xnor U18811 (N_18811,N_18787,N_18727);
nand U18812 (N_18812,N_18651,N_18603);
xor U18813 (N_18813,N_18762,N_18565);
xor U18814 (N_18814,N_18553,N_18628);
nand U18815 (N_18815,N_18793,N_18622);
nand U18816 (N_18816,N_18587,N_18784);
or U18817 (N_18817,N_18498,N_18467);
xor U18818 (N_18818,N_18644,N_18557);
nor U18819 (N_18819,N_18564,N_18673);
or U18820 (N_18820,N_18761,N_18766);
nand U18821 (N_18821,N_18519,N_18650);
and U18822 (N_18822,N_18764,N_18488);
nand U18823 (N_18823,N_18655,N_18600);
xor U18824 (N_18824,N_18544,N_18614);
nand U18825 (N_18825,N_18441,N_18653);
and U18826 (N_18826,N_18593,N_18668);
xnor U18827 (N_18827,N_18537,N_18575);
or U18828 (N_18828,N_18546,N_18558);
and U18829 (N_18829,N_18683,N_18635);
nor U18830 (N_18830,N_18620,N_18752);
nor U18831 (N_18831,N_18716,N_18405);
nor U18832 (N_18832,N_18714,N_18696);
nor U18833 (N_18833,N_18798,N_18486);
or U18834 (N_18834,N_18626,N_18461);
nand U18835 (N_18835,N_18539,N_18406);
and U18836 (N_18836,N_18453,N_18559);
or U18837 (N_18837,N_18450,N_18408);
nand U18838 (N_18838,N_18786,N_18538);
and U18839 (N_18839,N_18484,N_18670);
nor U18840 (N_18840,N_18616,N_18757);
xnor U18841 (N_18841,N_18728,N_18790);
xor U18842 (N_18842,N_18497,N_18609);
and U18843 (N_18843,N_18551,N_18529);
nand U18844 (N_18844,N_18432,N_18597);
xor U18845 (N_18845,N_18578,N_18638);
nor U18846 (N_18846,N_18783,N_18604);
and U18847 (N_18847,N_18476,N_18610);
nand U18848 (N_18848,N_18583,N_18427);
and U18849 (N_18849,N_18772,N_18706);
and U18850 (N_18850,N_18404,N_18634);
nand U18851 (N_18851,N_18499,N_18732);
nand U18852 (N_18852,N_18526,N_18411);
nor U18853 (N_18853,N_18779,N_18745);
and U18854 (N_18854,N_18658,N_18445);
nor U18855 (N_18855,N_18645,N_18724);
xor U18856 (N_18856,N_18505,N_18504);
nand U18857 (N_18857,N_18701,N_18680);
xor U18858 (N_18858,N_18443,N_18707);
or U18859 (N_18859,N_18734,N_18589);
and U18860 (N_18860,N_18400,N_18605);
nor U18861 (N_18861,N_18490,N_18588);
nand U18862 (N_18862,N_18699,N_18794);
or U18863 (N_18863,N_18652,N_18448);
nor U18864 (N_18864,N_18555,N_18754);
nand U18865 (N_18865,N_18465,N_18751);
nor U18866 (N_18866,N_18425,N_18694);
xor U18867 (N_18867,N_18483,N_18615);
nand U18868 (N_18868,N_18449,N_18534);
and U18869 (N_18869,N_18416,N_18639);
nor U18870 (N_18870,N_18574,N_18722);
and U18871 (N_18871,N_18741,N_18462);
and U18872 (N_18872,N_18672,N_18426);
xor U18873 (N_18873,N_18552,N_18735);
nand U18874 (N_18874,N_18641,N_18550);
xor U18875 (N_18875,N_18586,N_18682);
nand U18876 (N_18876,N_18776,N_18479);
nand U18877 (N_18877,N_18494,N_18617);
or U18878 (N_18878,N_18629,N_18520);
nand U18879 (N_18879,N_18729,N_18460);
nor U18880 (N_18880,N_18401,N_18591);
xor U18881 (N_18881,N_18611,N_18503);
and U18882 (N_18882,N_18511,N_18723);
xor U18883 (N_18883,N_18768,N_18797);
or U18884 (N_18884,N_18648,N_18523);
xnor U18885 (N_18885,N_18657,N_18469);
nand U18886 (N_18886,N_18767,N_18744);
nor U18887 (N_18887,N_18590,N_18627);
nor U18888 (N_18888,N_18545,N_18533);
nand U18889 (N_18889,N_18688,N_18665);
nor U18890 (N_18890,N_18632,N_18775);
or U18891 (N_18891,N_18571,N_18777);
nand U18892 (N_18892,N_18536,N_18746);
xnor U18893 (N_18893,N_18690,N_18618);
nor U18894 (N_18894,N_18518,N_18513);
nor U18895 (N_18895,N_18624,N_18780);
and U18896 (N_18896,N_18561,N_18759);
or U18897 (N_18897,N_18528,N_18407);
nand U18898 (N_18898,N_18472,N_18541);
and U18899 (N_18899,N_18771,N_18412);
nand U18900 (N_18900,N_18686,N_18548);
nand U18901 (N_18901,N_18585,N_18477);
nor U18902 (N_18902,N_18413,N_18693);
and U18903 (N_18903,N_18691,N_18451);
xor U18904 (N_18904,N_18760,N_18474);
xnor U18905 (N_18905,N_18778,N_18507);
nor U18906 (N_18906,N_18681,N_18791);
and U18907 (N_18907,N_18481,N_18749);
or U18908 (N_18908,N_18560,N_18619);
or U18909 (N_18909,N_18580,N_18656);
or U18910 (N_18910,N_18500,N_18799);
and U18911 (N_18911,N_18532,N_18527);
or U18912 (N_18912,N_18687,N_18444);
nor U18913 (N_18913,N_18418,N_18457);
xnor U18914 (N_18914,N_18662,N_18501);
nor U18915 (N_18915,N_18485,N_18421);
nand U18916 (N_18916,N_18514,N_18581);
xnor U18917 (N_18917,N_18623,N_18667);
or U18918 (N_18918,N_18702,N_18409);
xor U18919 (N_18919,N_18633,N_18703);
and U18920 (N_18920,N_18755,N_18606);
nand U18921 (N_18921,N_18473,N_18637);
nor U18922 (N_18922,N_18625,N_18640);
and U18923 (N_18923,N_18417,N_18795);
nand U18924 (N_18924,N_18666,N_18709);
and U18925 (N_18925,N_18758,N_18684);
or U18926 (N_18926,N_18705,N_18521);
nor U18927 (N_18927,N_18738,N_18423);
nor U18928 (N_18928,N_18643,N_18402);
and U18929 (N_18929,N_18595,N_18569);
and U18930 (N_18930,N_18750,N_18489);
and U18931 (N_18931,N_18612,N_18496);
and U18932 (N_18932,N_18543,N_18547);
xor U18933 (N_18933,N_18506,N_18740);
and U18934 (N_18934,N_18422,N_18711);
nor U18935 (N_18935,N_18608,N_18660);
xnor U18936 (N_18936,N_18446,N_18736);
xnor U18937 (N_18937,N_18669,N_18592);
or U18938 (N_18938,N_18649,N_18785);
xor U18939 (N_18939,N_18782,N_18512);
nand U18940 (N_18940,N_18563,N_18540);
nand U18941 (N_18941,N_18456,N_18430);
or U18942 (N_18942,N_18685,N_18470);
or U18943 (N_18943,N_18602,N_18577);
and U18944 (N_18944,N_18594,N_18742);
or U18945 (N_18945,N_18630,N_18573);
nor U18946 (N_18946,N_18475,N_18549);
nor U18947 (N_18947,N_18433,N_18434);
or U18948 (N_18948,N_18773,N_18769);
and U18949 (N_18949,N_18420,N_18596);
nand U18950 (N_18950,N_18419,N_18468);
and U18951 (N_18951,N_18502,N_18459);
or U18952 (N_18952,N_18509,N_18487);
xnor U18953 (N_18953,N_18613,N_18492);
and U18954 (N_18954,N_18570,N_18730);
or U18955 (N_18955,N_18671,N_18679);
or U18956 (N_18956,N_18458,N_18743);
xor U18957 (N_18957,N_18471,N_18788);
nor U18958 (N_18958,N_18566,N_18715);
or U18959 (N_18959,N_18663,N_18525);
or U18960 (N_18960,N_18770,N_18695);
nor U18961 (N_18961,N_18455,N_18576);
and U18962 (N_18962,N_18718,N_18535);
xnor U18963 (N_18963,N_18431,N_18495);
nand U18964 (N_18964,N_18524,N_18572);
xnor U18965 (N_18965,N_18725,N_18438);
or U18966 (N_18966,N_18428,N_18435);
xor U18967 (N_18967,N_18747,N_18717);
xnor U18968 (N_18968,N_18437,N_18756);
and U18969 (N_18969,N_18567,N_18631);
xor U18970 (N_18970,N_18636,N_18720);
or U18971 (N_18971,N_18582,N_18517);
nand U18972 (N_18972,N_18674,N_18599);
xnor U18973 (N_18973,N_18710,N_18698);
nor U18974 (N_18974,N_18414,N_18424);
xor U18975 (N_18975,N_18439,N_18579);
xnor U18976 (N_18976,N_18748,N_18659);
and U18977 (N_18977,N_18482,N_18664);
nand U18978 (N_18978,N_18689,N_18480);
xnor U18979 (N_18979,N_18556,N_18719);
or U18980 (N_18980,N_18692,N_18554);
or U18981 (N_18981,N_18704,N_18646);
or U18982 (N_18982,N_18642,N_18621);
and U18983 (N_18983,N_18647,N_18452);
nand U18984 (N_18984,N_18491,N_18601);
or U18985 (N_18985,N_18568,N_18493);
xnor U18986 (N_18986,N_18796,N_18697);
nor U18987 (N_18987,N_18508,N_18515);
nor U18988 (N_18988,N_18792,N_18562);
nand U18989 (N_18989,N_18700,N_18721);
xnor U18990 (N_18990,N_18789,N_18708);
xnor U18991 (N_18991,N_18429,N_18410);
nand U18992 (N_18992,N_18542,N_18530);
nor U18993 (N_18993,N_18403,N_18440);
xor U18994 (N_18994,N_18712,N_18454);
xnor U18995 (N_18995,N_18678,N_18713);
nor U18996 (N_18996,N_18781,N_18731);
or U18997 (N_18997,N_18463,N_18675);
nor U18998 (N_18998,N_18415,N_18531);
nand U18999 (N_18999,N_18442,N_18510);
and U19000 (N_19000,N_18645,N_18682);
xnor U19001 (N_19001,N_18595,N_18498);
or U19002 (N_19002,N_18710,N_18620);
xnor U19003 (N_19003,N_18636,N_18675);
or U19004 (N_19004,N_18596,N_18728);
xnor U19005 (N_19005,N_18718,N_18795);
and U19006 (N_19006,N_18461,N_18568);
and U19007 (N_19007,N_18493,N_18776);
and U19008 (N_19008,N_18613,N_18533);
xor U19009 (N_19009,N_18710,N_18676);
xnor U19010 (N_19010,N_18790,N_18592);
and U19011 (N_19011,N_18464,N_18524);
xor U19012 (N_19012,N_18604,N_18711);
xnor U19013 (N_19013,N_18486,N_18608);
nor U19014 (N_19014,N_18680,N_18656);
and U19015 (N_19015,N_18590,N_18549);
or U19016 (N_19016,N_18496,N_18501);
and U19017 (N_19017,N_18503,N_18566);
nand U19018 (N_19018,N_18543,N_18600);
xor U19019 (N_19019,N_18716,N_18781);
xnor U19020 (N_19020,N_18765,N_18544);
xor U19021 (N_19021,N_18607,N_18599);
or U19022 (N_19022,N_18622,N_18657);
nand U19023 (N_19023,N_18447,N_18591);
nand U19024 (N_19024,N_18635,N_18728);
or U19025 (N_19025,N_18518,N_18686);
nor U19026 (N_19026,N_18517,N_18512);
nor U19027 (N_19027,N_18699,N_18560);
or U19028 (N_19028,N_18508,N_18414);
nand U19029 (N_19029,N_18412,N_18501);
nor U19030 (N_19030,N_18489,N_18524);
nand U19031 (N_19031,N_18563,N_18766);
nor U19032 (N_19032,N_18720,N_18443);
and U19033 (N_19033,N_18760,N_18614);
nand U19034 (N_19034,N_18625,N_18430);
nor U19035 (N_19035,N_18574,N_18501);
and U19036 (N_19036,N_18411,N_18436);
xnor U19037 (N_19037,N_18508,N_18550);
and U19038 (N_19038,N_18488,N_18598);
or U19039 (N_19039,N_18607,N_18724);
xnor U19040 (N_19040,N_18752,N_18734);
nand U19041 (N_19041,N_18635,N_18490);
nand U19042 (N_19042,N_18676,N_18733);
and U19043 (N_19043,N_18611,N_18492);
and U19044 (N_19044,N_18661,N_18509);
and U19045 (N_19045,N_18639,N_18746);
nand U19046 (N_19046,N_18658,N_18715);
and U19047 (N_19047,N_18691,N_18455);
xor U19048 (N_19048,N_18590,N_18566);
and U19049 (N_19049,N_18593,N_18664);
or U19050 (N_19050,N_18581,N_18421);
xor U19051 (N_19051,N_18559,N_18482);
xor U19052 (N_19052,N_18646,N_18781);
and U19053 (N_19053,N_18451,N_18530);
and U19054 (N_19054,N_18681,N_18658);
nand U19055 (N_19055,N_18617,N_18484);
nor U19056 (N_19056,N_18479,N_18692);
or U19057 (N_19057,N_18411,N_18564);
or U19058 (N_19058,N_18569,N_18610);
xor U19059 (N_19059,N_18551,N_18603);
or U19060 (N_19060,N_18536,N_18682);
or U19061 (N_19061,N_18735,N_18614);
or U19062 (N_19062,N_18548,N_18735);
xor U19063 (N_19063,N_18738,N_18461);
xnor U19064 (N_19064,N_18439,N_18493);
nor U19065 (N_19065,N_18722,N_18582);
nor U19066 (N_19066,N_18573,N_18422);
xor U19067 (N_19067,N_18560,N_18443);
or U19068 (N_19068,N_18761,N_18515);
nor U19069 (N_19069,N_18662,N_18742);
or U19070 (N_19070,N_18560,N_18766);
or U19071 (N_19071,N_18730,N_18554);
and U19072 (N_19072,N_18757,N_18726);
nor U19073 (N_19073,N_18623,N_18764);
or U19074 (N_19074,N_18637,N_18442);
nand U19075 (N_19075,N_18708,N_18673);
nand U19076 (N_19076,N_18481,N_18516);
and U19077 (N_19077,N_18442,N_18646);
nor U19078 (N_19078,N_18699,N_18484);
and U19079 (N_19079,N_18444,N_18555);
or U19080 (N_19080,N_18484,N_18691);
and U19081 (N_19081,N_18561,N_18425);
nor U19082 (N_19082,N_18501,N_18709);
nand U19083 (N_19083,N_18662,N_18751);
or U19084 (N_19084,N_18569,N_18631);
nor U19085 (N_19085,N_18437,N_18653);
or U19086 (N_19086,N_18460,N_18578);
nor U19087 (N_19087,N_18486,N_18620);
nand U19088 (N_19088,N_18429,N_18493);
and U19089 (N_19089,N_18569,N_18760);
nand U19090 (N_19090,N_18404,N_18540);
xnor U19091 (N_19091,N_18443,N_18420);
xnor U19092 (N_19092,N_18490,N_18628);
and U19093 (N_19093,N_18762,N_18487);
or U19094 (N_19094,N_18745,N_18403);
or U19095 (N_19095,N_18512,N_18626);
and U19096 (N_19096,N_18798,N_18619);
and U19097 (N_19097,N_18547,N_18669);
and U19098 (N_19098,N_18669,N_18716);
xnor U19099 (N_19099,N_18618,N_18578);
xnor U19100 (N_19100,N_18573,N_18605);
and U19101 (N_19101,N_18774,N_18619);
xor U19102 (N_19102,N_18584,N_18582);
or U19103 (N_19103,N_18513,N_18579);
nand U19104 (N_19104,N_18725,N_18466);
xor U19105 (N_19105,N_18739,N_18488);
xnor U19106 (N_19106,N_18588,N_18766);
and U19107 (N_19107,N_18689,N_18743);
or U19108 (N_19108,N_18530,N_18434);
and U19109 (N_19109,N_18682,N_18515);
nand U19110 (N_19110,N_18403,N_18775);
or U19111 (N_19111,N_18527,N_18781);
nand U19112 (N_19112,N_18551,N_18554);
nor U19113 (N_19113,N_18637,N_18406);
nor U19114 (N_19114,N_18710,N_18424);
or U19115 (N_19115,N_18769,N_18482);
nand U19116 (N_19116,N_18731,N_18565);
or U19117 (N_19117,N_18657,N_18617);
xor U19118 (N_19118,N_18761,N_18623);
nor U19119 (N_19119,N_18726,N_18630);
and U19120 (N_19120,N_18552,N_18535);
nand U19121 (N_19121,N_18514,N_18714);
xnor U19122 (N_19122,N_18584,N_18697);
and U19123 (N_19123,N_18794,N_18509);
or U19124 (N_19124,N_18677,N_18420);
xnor U19125 (N_19125,N_18538,N_18771);
or U19126 (N_19126,N_18468,N_18571);
nor U19127 (N_19127,N_18692,N_18495);
xnor U19128 (N_19128,N_18640,N_18791);
nand U19129 (N_19129,N_18583,N_18561);
or U19130 (N_19130,N_18766,N_18593);
nand U19131 (N_19131,N_18772,N_18579);
nor U19132 (N_19132,N_18706,N_18731);
nand U19133 (N_19133,N_18537,N_18670);
xor U19134 (N_19134,N_18541,N_18455);
nand U19135 (N_19135,N_18772,N_18751);
and U19136 (N_19136,N_18751,N_18565);
and U19137 (N_19137,N_18785,N_18528);
nand U19138 (N_19138,N_18624,N_18761);
or U19139 (N_19139,N_18646,N_18491);
or U19140 (N_19140,N_18402,N_18549);
xor U19141 (N_19141,N_18771,N_18456);
nand U19142 (N_19142,N_18525,N_18680);
nand U19143 (N_19143,N_18472,N_18486);
and U19144 (N_19144,N_18711,N_18463);
nand U19145 (N_19145,N_18720,N_18623);
nand U19146 (N_19146,N_18650,N_18679);
nor U19147 (N_19147,N_18694,N_18570);
nor U19148 (N_19148,N_18621,N_18541);
nor U19149 (N_19149,N_18468,N_18709);
xor U19150 (N_19150,N_18705,N_18416);
or U19151 (N_19151,N_18408,N_18718);
and U19152 (N_19152,N_18733,N_18404);
nor U19153 (N_19153,N_18536,N_18718);
and U19154 (N_19154,N_18613,N_18758);
or U19155 (N_19155,N_18656,N_18473);
and U19156 (N_19156,N_18628,N_18520);
and U19157 (N_19157,N_18624,N_18593);
or U19158 (N_19158,N_18493,N_18704);
nor U19159 (N_19159,N_18403,N_18638);
nand U19160 (N_19160,N_18458,N_18742);
and U19161 (N_19161,N_18601,N_18773);
and U19162 (N_19162,N_18476,N_18759);
and U19163 (N_19163,N_18686,N_18723);
and U19164 (N_19164,N_18790,N_18428);
and U19165 (N_19165,N_18615,N_18717);
xnor U19166 (N_19166,N_18596,N_18519);
and U19167 (N_19167,N_18756,N_18608);
or U19168 (N_19168,N_18561,N_18414);
xor U19169 (N_19169,N_18669,N_18520);
nand U19170 (N_19170,N_18744,N_18755);
xor U19171 (N_19171,N_18404,N_18487);
xor U19172 (N_19172,N_18547,N_18584);
nand U19173 (N_19173,N_18508,N_18421);
or U19174 (N_19174,N_18641,N_18441);
nor U19175 (N_19175,N_18602,N_18461);
and U19176 (N_19176,N_18608,N_18421);
xnor U19177 (N_19177,N_18603,N_18660);
or U19178 (N_19178,N_18618,N_18581);
nor U19179 (N_19179,N_18700,N_18628);
and U19180 (N_19180,N_18496,N_18431);
nand U19181 (N_19181,N_18787,N_18669);
nor U19182 (N_19182,N_18468,N_18404);
nor U19183 (N_19183,N_18584,N_18544);
and U19184 (N_19184,N_18675,N_18771);
and U19185 (N_19185,N_18651,N_18788);
xor U19186 (N_19186,N_18512,N_18587);
nand U19187 (N_19187,N_18644,N_18454);
and U19188 (N_19188,N_18548,N_18695);
or U19189 (N_19189,N_18636,N_18461);
and U19190 (N_19190,N_18598,N_18502);
xor U19191 (N_19191,N_18695,N_18458);
nor U19192 (N_19192,N_18686,N_18409);
xor U19193 (N_19193,N_18647,N_18665);
nor U19194 (N_19194,N_18538,N_18548);
or U19195 (N_19195,N_18558,N_18548);
xnor U19196 (N_19196,N_18637,N_18403);
or U19197 (N_19197,N_18498,N_18557);
nand U19198 (N_19198,N_18455,N_18414);
or U19199 (N_19199,N_18603,N_18522);
or U19200 (N_19200,N_18898,N_19161);
nor U19201 (N_19201,N_19124,N_19115);
xor U19202 (N_19202,N_19151,N_18873);
or U19203 (N_19203,N_18809,N_18992);
xor U19204 (N_19204,N_19006,N_19178);
xnor U19205 (N_19205,N_19080,N_19194);
xor U19206 (N_19206,N_19136,N_19010);
nand U19207 (N_19207,N_19116,N_18911);
nor U19208 (N_19208,N_19030,N_18814);
or U19209 (N_19209,N_19065,N_19135);
or U19210 (N_19210,N_18946,N_18906);
nor U19211 (N_19211,N_19113,N_18917);
nand U19212 (N_19212,N_18940,N_18936);
or U19213 (N_19213,N_19049,N_19199);
xnor U19214 (N_19214,N_18895,N_19078);
nand U19215 (N_19215,N_19003,N_18942);
nand U19216 (N_19216,N_19037,N_18830);
or U19217 (N_19217,N_19104,N_18851);
nor U19218 (N_19218,N_18881,N_19072);
nor U19219 (N_19219,N_18897,N_18944);
nor U19220 (N_19220,N_18833,N_18891);
nand U19221 (N_19221,N_19012,N_18935);
or U19222 (N_19222,N_18822,N_19097);
or U19223 (N_19223,N_19190,N_19160);
xnor U19224 (N_19224,N_19034,N_19064);
nor U19225 (N_19225,N_19150,N_18888);
nor U19226 (N_19226,N_19172,N_19058);
and U19227 (N_19227,N_18913,N_18981);
nor U19228 (N_19228,N_19120,N_18959);
xor U19229 (N_19229,N_18912,N_18988);
and U19230 (N_19230,N_18815,N_18871);
xnor U19231 (N_19231,N_19093,N_18952);
nand U19232 (N_19232,N_19070,N_19192);
xnor U19233 (N_19233,N_19167,N_19028);
and U19234 (N_19234,N_19019,N_18941);
and U19235 (N_19235,N_18987,N_19016);
and U19236 (N_19236,N_19011,N_18982);
or U19237 (N_19237,N_18965,N_19189);
nand U19238 (N_19238,N_19043,N_19153);
or U19239 (N_19239,N_19023,N_19108);
nor U19240 (N_19240,N_19089,N_18824);
xnor U19241 (N_19241,N_18933,N_19057);
and U19242 (N_19242,N_18893,N_18882);
nand U19243 (N_19243,N_19038,N_19056);
and U19244 (N_19244,N_18819,N_19148);
nand U19245 (N_19245,N_18909,N_18872);
nand U19246 (N_19246,N_19159,N_19177);
nand U19247 (N_19247,N_18949,N_19143);
xnor U19248 (N_19248,N_18900,N_19081);
nor U19249 (N_19249,N_18957,N_19195);
xnor U19250 (N_19250,N_18969,N_19087);
and U19251 (N_19251,N_19067,N_18995);
and U19252 (N_19252,N_19032,N_19026);
xnor U19253 (N_19253,N_18915,N_19005);
nor U19254 (N_19254,N_18876,N_18825);
and U19255 (N_19255,N_19013,N_18805);
and U19256 (N_19256,N_18828,N_18963);
and U19257 (N_19257,N_19186,N_18863);
and U19258 (N_19258,N_19083,N_18804);
or U19259 (N_19259,N_19193,N_19074);
nor U19260 (N_19260,N_18829,N_18993);
or U19261 (N_19261,N_19176,N_18928);
xnor U19262 (N_19262,N_18803,N_18978);
or U19263 (N_19263,N_18996,N_18999);
nand U19264 (N_19264,N_18997,N_18938);
xor U19265 (N_19265,N_18954,N_19145);
and U19266 (N_19266,N_19060,N_19029);
or U19267 (N_19267,N_19059,N_18813);
xnor U19268 (N_19268,N_19147,N_18967);
or U19269 (N_19269,N_18958,N_18847);
xor U19270 (N_19270,N_18855,N_18848);
nor U19271 (N_19271,N_18979,N_18905);
nand U19272 (N_19272,N_19095,N_18924);
nor U19273 (N_19273,N_18904,N_19133);
and U19274 (N_19274,N_19175,N_18826);
nand U19275 (N_19275,N_19140,N_19007);
nor U19276 (N_19276,N_19126,N_18930);
xnor U19277 (N_19277,N_19179,N_19073);
or U19278 (N_19278,N_18887,N_18885);
xnor U19279 (N_19279,N_18820,N_19017);
and U19280 (N_19280,N_19048,N_19168);
nand U19281 (N_19281,N_19085,N_19122);
xor U19282 (N_19282,N_19014,N_18810);
or U19283 (N_19283,N_19198,N_19157);
xnor U19284 (N_19284,N_18970,N_18836);
nor U19285 (N_19285,N_19053,N_19101);
nand U19286 (N_19286,N_18947,N_19075);
nand U19287 (N_19287,N_18832,N_18914);
nand U19288 (N_19288,N_19050,N_19027);
nand U19289 (N_19289,N_18844,N_19106);
and U19290 (N_19290,N_19098,N_18899);
xor U19291 (N_19291,N_18922,N_18870);
and U19292 (N_19292,N_18837,N_18983);
and U19293 (N_19293,N_18955,N_19197);
or U19294 (N_19294,N_19054,N_19045);
xor U19295 (N_19295,N_18934,N_18960);
xor U19296 (N_19296,N_18968,N_18869);
and U19297 (N_19297,N_18961,N_18849);
and U19298 (N_19298,N_18834,N_19127);
nand U19299 (N_19299,N_18910,N_19099);
nor U19300 (N_19300,N_19139,N_18854);
xor U19301 (N_19301,N_18916,N_18994);
or U19302 (N_19302,N_18927,N_18861);
or U19303 (N_19303,N_19042,N_18807);
nand U19304 (N_19304,N_18806,N_18908);
nand U19305 (N_19305,N_18894,N_18956);
xor U19306 (N_19306,N_18835,N_19103);
and U19307 (N_19307,N_18989,N_19020);
nand U19308 (N_19308,N_18827,N_19066);
or U19309 (N_19309,N_19171,N_18932);
nand U19310 (N_19310,N_18831,N_18976);
nand U19311 (N_19311,N_19021,N_18842);
xor U19312 (N_19312,N_19094,N_19111);
xor U19313 (N_19313,N_18853,N_19117);
or U19314 (N_19314,N_19142,N_19022);
xnor U19315 (N_19315,N_18817,N_18858);
or U19316 (N_19316,N_18953,N_19096);
nand U19317 (N_19317,N_19182,N_18864);
nand U19318 (N_19318,N_18821,N_18943);
nor U19319 (N_19319,N_18883,N_18902);
or U19320 (N_19320,N_19044,N_18921);
nand U19321 (N_19321,N_19138,N_19123);
nor U19322 (N_19322,N_18856,N_18901);
xnor U19323 (N_19323,N_19162,N_19137);
and U19324 (N_19324,N_19125,N_19033);
nor U19325 (N_19325,N_19181,N_19082);
and U19326 (N_19326,N_18991,N_18950);
nor U19327 (N_19327,N_18865,N_19128);
xor U19328 (N_19328,N_18962,N_18931);
and U19329 (N_19329,N_19114,N_18878);
or U19330 (N_19330,N_18801,N_19149);
xnor U19331 (N_19331,N_19134,N_19121);
or U19332 (N_19332,N_18918,N_18811);
nor U19333 (N_19333,N_18966,N_18859);
nor U19334 (N_19334,N_19119,N_19000);
and U19335 (N_19335,N_19112,N_19154);
xor U19336 (N_19336,N_18802,N_18846);
xnor U19337 (N_19337,N_19166,N_18937);
or U19338 (N_19338,N_19184,N_19001);
xnor U19339 (N_19339,N_18977,N_18860);
xnor U19340 (N_19340,N_18926,N_19025);
nor U19341 (N_19341,N_18880,N_18852);
xnor U19342 (N_19342,N_18986,N_18980);
nor U19343 (N_19343,N_19035,N_19055);
nand U19344 (N_19344,N_19163,N_18998);
nand U19345 (N_19345,N_19152,N_19187);
nand U19346 (N_19346,N_19110,N_18886);
and U19347 (N_19347,N_19024,N_19141);
xor U19348 (N_19348,N_19046,N_18973);
or U19349 (N_19349,N_19041,N_19077);
or U19350 (N_19350,N_19183,N_19156);
nor U19351 (N_19351,N_18866,N_19088);
nand U19352 (N_19352,N_19170,N_19144);
nor U19353 (N_19353,N_18875,N_19052);
and U19354 (N_19354,N_18948,N_18919);
and U19355 (N_19355,N_19174,N_18816);
nand U19356 (N_19356,N_19062,N_18951);
and U19357 (N_19357,N_18975,N_19102);
and U19358 (N_19358,N_19031,N_18964);
nand U19359 (N_19359,N_19018,N_19090);
or U19360 (N_19360,N_18974,N_19109);
and U19361 (N_19361,N_19196,N_19146);
or U19362 (N_19362,N_19188,N_19084);
nand U19363 (N_19363,N_18923,N_19185);
and U19364 (N_19364,N_19076,N_18939);
or U19365 (N_19365,N_19173,N_18985);
nand U19366 (N_19366,N_18800,N_19061);
xnor U19367 (N_19367,N_19036,N_19107);
nor U19368 (N_19368,N_19165,N_19129);
xor U19369 (N_19369,N_19004,N_19180);
nor U19370 (N_19370,N_19009,N_19051);
xor U19371 (N_19371,N_19039,N_18903);
and U19372 (N_19372,N_19132,N_19047);
xnor U19373 (N_19373,N_18838,N_18843);
nor U19374 (N_19374,N_19040,N_18818);
xnor U19375 (N_19375,N_19091,N_19068);
nand U19376 (N_19376,N_19015,N_19169);
and U19377 (N_19377,N_18839,N_18857);
and U19378 (N_19378,N_18862,N_18907);
nor U19379 (N_19379,N_18868,N_19008);
xnor U19380 (N_19380,N_19105,N_18971);
xnor U19381 (N_19381,N_19164,N_19071);
nor U19382 (N_19382,N_18925,N_19155);
and U19383 (N_19383,N_18892,N_18845);
xor U19384 (N_19384,N_19063,N_18984);
nor U19385 (N_19385,N_18884,N_19191);
xnor U19386 (N_19386,N_18972,N_18877);
xor U19387 (N_19387,N_18945,N_18840);
xor U19388 (N_19388,N_18879,N_18889);
nand U19389 (N_19389,N_19130,N_18929);
nand U19390 (N_19390,N_19086,N_18850);
and U19391 (N_19391,N_18812,N_19131);
nand U19392 (N_19392,N_18920,N_18808);
nor U19393 (N_19393,N_18874,N_19002);
nor U19394 (N_19394,N_18867,N_19158);
or U19395 (N_19395,N_19079,N_19118);
and U19396 (N_19396,N_19100,N_19092);
nor U19397 (N_19397,N_18896,N_18823);
or U19398 (N_19398,N_18990,N_18890);
nor U19399 (N_19399,N_18841,N_19069);
nand U19400 (N_19400,N_18898,N_18837);
nand U19401 (N_19401,N_18956,N_19076);
nand U19402 (N_19402,N_19084,N_18830);
nand U19403 (N_19403,N_18956,N_19195);
nand U19404 (N_19404,N_18974,N_18868);
nor U19405 (N_19405,N_19033,N_18991);
or U19406 (N_19406,N_18934,N_18969);
and U19407 (N_19407,N_19098,N_19021);
and U19408 (N_19408,N_18865,N_19033);
xnor U19409 (N_19409,N_18848,N_19097);
or U19410 (N_19410,N_18910,N_18889);
nand U19411 (N_19411,N_19028,N_19018);
nor U19412 (N_19412,N_18966,N_19053);
nand U19413 (N_19413,N_18854,N_19173);
or U19414 (N_19414,N_19157,N_19188);
and U19415 (N_19415,N_18801,N_18985);
nor U19416 (N_19416,N_18881,N_18873);
and U19417 (N_19417,N_18817,N_19048);
or U19418 (N_19418,N_19074,N_18991);
xnor U19419 (N_19419,N_19162,N_19181);
nor U19420 (N_19420,N_18901,N_19079);
nor U19421 (N_19421,N_18841,N_19013);
and U19422 (N_19422,N_19133,N_18803);
and U19423 (N_19423,N_18812,N_19004);
nor U19424 (N_19424,N_19129,N_19147);
nor U19425 (N_19425,N_19185,N_18971);
or U19426 (N_19426,N_19085,N_18823);
nand U19427 (N_19427,N_19013,N_19145);
or U19428 (N_19428,N_18976,N_19061);
xor U19429 (N_19429,N_19093,N_19164);
and U19430 (N_19430,N_19025,N_19191);
or U19431 (N_19431,N_19030,N_19097);
or U19432 (N_19432,N_19109,N_18998);
xnor U19433 (N_19433,N_19151,N_18853);
or U19434 (N_19434,N_18803,N_18843);
and U19435 (N_19435,N_19108,N_18978);
and U19436 (N_19436,N_19131,N_18837);
and U19437 (N_19437,N_18820,N_18815);
nand U19438 (N_19438,N_18890,N_19080);
or U19439 (N_19439,N_19197,N_18825);
xor U19440 (N_19440,N_18994,N_19187);
nor U19441 (N_19441,N_18964,N_19124);
or U19442 (N_19442,N_19047,N_18970);
and U19443 (N_19443,N_18884,N_19133);
or U19444 (N_19444,N_18939,N_19095);
nand U19445 (N_19445,N_19072,N_19062);
nand U19446 (N_19446,N_18890,N_19123);
xnor U19447 (N_19447,N_19125,N_18984);
or U19448 (N_19448,N_19059,N_18850);
xor U19449 (N_19449,N_19038,N_18937);
nor U19450 (N_19450,N_18814,N_18809);
nand U19451 (N_19451,N_18853,N_18941);
or U19452 (N_19452,N_19082,N_18839);
nand U19453 (N_19453,N_19077,N_19107);
nor U19454 (N_19454,N_18882,N_19035);
xnor U19455 (N_19455,N_18930,N_19058);
xnor U19456 (N_19456,N_18945,N_18803);
or U19457 (N_19457,N_19171,N_19121);
and U19458 (N_19458,N_18804,N_18976);
or U19459 (N_19459,N_18865,N_18979);
nor U19460 (N_19460,N_18971,N_19003);
or U19461 (N_19461,N_19109,N_18801);
nor U19462 (N_19462,N_19077,N_19002);
nor U19463 (N_19463,N_19058,N_19046);
xnor U19464 (N_19464,N_19176,N_19095);
xor U19465 (N_19465,N_19048,N_18871);
or U19466 (N_19466,N_19066,N_19032);
nand U19467 (N_19467,N_19125,N_18869);
or U19468 (N_19468,N_19050,N_18881);
and U19469 (N_19469,N_19035,N_19010);
nand U19470 (N_19470,N_19075,N_18857);
xor U19471 (N_19471,N_19020,N_18897);
or U19472 (N_19472,N_19160,N_18875);
nand U19473 (N_19473,N_19020,N_19025);
xor U19474 (N_19474,N_18892,N_19125);
and U19475 (N_19475,N_18939,N_19156);
nor U19476 (N_19476,N_19188,N_19062);
and U19477 (N_19477,N_19005,N_18941);
and U19478 (N_19478,N_18895,N_18912);
nand U19479 (N_19479,N_19189,N_19161);
or U19480 (N_19480,N_19177,N_18933);
xor U19481 (N_19481,N_19170,N_18986);
and U19482 (N_19482,N_18902,N_19187);
or U19483 (N_19483,N_19044,N_18864);
and U19484 (N_19484,N_18953,N_19163);
or U19485 (N_19485,N_19136,N_19158);
nor U19486 (N_19486,N_19005,N_19195);
nand U19487 (N_19487,N_18921,N_19154);
and U19488 (N_19488,N_19109,N_18973);
nor U19489 (N_19489,N_19003,N_19199);
nand U19490 (N_19490,N_19133,N_19110);
xor U19491 (N_19491,N_18868,N_18982);
nand U19492 (N_19492,N_18961,N_18837);
nand U19493 (N_19493,N_18946,N_19178);
and U19494 (N_19494,N_19172,N_19060);
xnor U19495 (N_19495,N_19062,N_18806);
and U19496 (N_19496,N_19147,N_19197);
nor U19497 (N_19497,N_18824,N_19009);
or U19498 (N_19498,N_18860,N_19156);
and U19499 (N_19499,N_19064,N_19178);
nand U19500 (N_19500,N_19051,N_18981);
nand U19501 (N_19501,N_19056,N_18864);
and U19502 (N_19502,N_19061,N_19101);
xnor U19503 (N_19503,N_19170,N_18968);
or U19504 (N_19504,N_18851,N_19158);
and U19505 (N_19505,N_19037,N_19174);
and U19506 (N_19506,N_19142,N_18835);
and U19507 (N_19507,N_19015,N_18952);
nor U19508 (N_19508,N_19025,N_19019);
xor U19509 (N_19509,N_18865,N_18998);
nand U19510 (N_19510,N_18986,N_18984);
and U19511 (N_19511,N_18932,N_18996);
and U19512 (N_19512,N_19152,N_19061);
or U19513 (N_19513,N_19027,N_19092);
and U19514 (N_19514,N_18826,N_18952);
xnor U19515 (N_19515,N_18800,N_19003);
or U19516 (N_19516,N_18923,N_19057);
and U19517 (N_19517,N_18940,N_19145);
nand U19518 (N_19518,N_18939,N_19084);
or U19519 (N_19519,N_19036,N_18901);
or U19520 (N_19520,N_19042,N_19090);
nor U19521 (N_19521,N_19066,N_19115);
xnor U19522 (N_19522,N_18916,N_19089);
nor U19523 (N_19523,N_19019,N_18814);
nor U19524 (N_19524,N_19182,N_18867);
or U19525 (N_19525,N_19078,N_18830);
or U19526 (N_19526,N_18862,N_19185);
xnor U19527 (N_19527,N_19127,N_18825);
xnor U19528 (N_19528,N_18906,N_19013);
nor U19529 (N_19529,N_18895,N_19159);
nor U19530 (N_19530,N_19051,N_19163);
nand U19531 (N_19531,N_19047,N_18849);
or U19532 (N_19532,N_18956,N_18821);
xnor U19533 (N_19533,N_18930,N_19161);
and U19534 (N_19534,N_19060,N_18873);
and U19535 (N_19535,N_18931,N_18861);
and U19536 (N_19536,N_18839,N_19052);
or U19537 (N_19537,N_18958,N_19056);
nand U19538 (N_19538,N_18801,N_18831);
nand U19539 (N_19539,N_18812,N_18939);
and U19540 (N_19540,N_19111,N_19080);
nor U19541 (N_19541,N_18804,N_18809);
nand U19542 (N_19542,N_19126,N_19088);
or U19543 (N_19543,N_19112,N_18982);
or U19544 (N_19544,N_18800,N_19104);
or U19545 (N_19545,N_19154,N_18990);
nor U19546 (N_19546,N_19081,N_19171);
and U19547 (N_19547,N_18901,N_18950);
nand U19548 (N_19548,N_18965,N_18911);
and U19549 (N_19549,N_19007,N_18932);
and U19550 (N_19550,N_18973,N_19027);
nand U19551 (N_19551,N_19171,N_18971);
xnor U19552 (N_19552,N_18812,N_19198);
nor U19553 (N_19553,N_19046,N_18991);
and U19554 (N_19554,N_18897,N_19080);
nor U19555 (N_19555,N_19047,N_18841);
nor U19556 (N_19556,N_19187,N_19133);
nand U19557 (N_19557,N_19022,N_18865);
or U19558 (N_19558,N_19093,N_18871);
or U19559 (N_19559,N_19032,N_19096);
or U19560 (N_19560,N_19092,N_18836);
or U19561 (N_19561,N_18932,N_18843);
xor U19562 (N_19562,N_18994,N_18854);
xnor U19563 (N_19563,N_19003,N_19027);
nor U19564 (N_19564,N_19078,N_18892);
nor U19565 (N_19565,N_18814,N_18829);
nor U19566 (N_19566,N_18862,N_18950);
nand U19567 (N_19567,N_18882,N_19128);
xnor U19568 (N_19568,N_19050,N_18960);
nor U19569 (N_19569,N_19000,N_18863);
and U19570 (N_19570,N_19072,N_18862);
nor U19571 (N_19571,N_19058,N_19181);
and U19572 (N_19572,N_18933,N_18981);
xnor U19573 (N_19573,N_19139,N_19147);
and U19574 (N_19574,N_18908,N_18814);
nand U19575 (N_19575,N_19012,N_19188);
or U19576 (N_19576,N_19038,N_18981);
xnor U19577 (N_19577,N_19102,N_18880);
xnor U19578 (N_19578,N_19078,N_18826);
xnor U19579 (N_19579,N_19004,N_19081);
and U19580 (N_19580,N_19049,N_18835);
and U19581 (N_19581,N_18944,N_18863);
or U19582 (N_19582,N_19160,N_18873);
or U19583 (N_19583,N_19069,N_18830);
nor U19584 (N_19584,N_19000,N_18813);
xnor U19585 (N_19585,N_19130,N_18918);
or U19586 (N_19586,N_18985,N_19170);
or U19587 (N_19587,N_18966,N_18811);
nand U19588 (N_19588,N_18897,N_19097);
nor U19589 (N_19589,N_19101,N_18995);
xor U19590 (N_19590,N_19061,N_18809);
and U19591 (N_19591,N_19129,N_18998);
nand U19592 (N_19592,N_18896,N_19086);
and U19593 (N_19593,N_18821,N_19034);
and U19594 (N_19594,N_18850,N_19020);
nor U19595 (N_19595,N_18878,N_19128);
nand U19596 (N_19596,N_18842,N_18873);
and U19597 (N_19597,N_18821,N_19138);
xnor U19598 (N_19598,N_19054,N_19167);
xnor U19599 (N_19599,N_18915,N_19046);
and U19600 (N_19600,N_19406,N_19306);
nor U19601 (N_19601,N_19481,N_19388);
nand U19602 (N_19602,N_19597,N_19462);
or U19603 (N_19603,N_19452,N_19568);
or U19604 (N_19604,N_19264,N_19276);
nor U19605 (N_19605,N_19522,N_19420);
and U19606 (N_19606,N_19407,N_19281);
and U19607 (N_19607,N_19556,N_19582);
xnor U19608 (N_19608,N_19552,N_19313);
or U19609 (N_19609,N_19256,N_19223);
xor U19610 (N_19610,N_19561,N_19501);
nand U19611 (N_19611,N_19360,N_19373);
or U19612 (N_19612,N_19327,N_19247);
xnor U19613 (N_19613,N_19357,N_19206);
and U19614 (N_19614,N_19564,N_19227);
xor U19615 (N_19615,N_19450,N_19216);
and U19616 (N_19616,N_19362,N_19576);
xor U19617 (N_19617,N_19364,N_19479);
or U19618 (N_19618,N_19555,N_19574);
nand U19619 (N_19619,N_19330,N_19415);
or U19620 (N_19620,N_19288,N_19549);
xnor U19621 (N_19621,N_19525,N_19397);
xnor U19622 (N_19622,N_19521,N_19465);
nand U19623 (N_19623,N_19245,N_19225);
nand U19624 (N_19624,N_19200,N_19296);
xor U19625 (N_19625,N_19535,N_19548);
nand U19626 (N_19626,N_19207,N_19229);
nand U19627 (N_19627,N_19546,N_19346);
nand U19628 (N_19628,N_19591,N_19380);
and U19629 (N_19629,N_19491,N_19512);
or U19630 (N_19630,N_19459,N_19429);
xnor U19631 (N_19631,N_19280,N_19454);
or U19632 (N_19632,N_19218,N_19285);
and U19633 (N_19633,N_19414,N_19493);
and U19634 (N_19634,N_19349,N_19248);
nand U19635 (N_19635,N_19261,N_19215);
xor U19636 (N_19636,N_19560,N_19352);
xnor U19637 (N_19637,N_19550,N_19500);
nand U19638 (N_19638,N_19508,N_19209);
xor U19639 (N_19639,N_19490,N_19234);
or U19640 (N_19640,N_19316,N_19343);
xnor U19641 (N_19641,N_19580,N_19401);
and U19642 (N_19642,N_19290,N_19437);
nand U19643 (N_19643,N_19328,N_19539);
nand U19644 (N_19644,N_19531,N_19260);
xnor U19645 (N_19645,N_19404,N_19381);
xor U19646 (N_19646,N_19503,N_19312);
and U19647 (N_19647,N_19228,N_19272);
xnor U19648 (N_19648,N_19338,N_19433);
nand U19649 (N_19649,N_19239,N_19505);
and U19650 (N_19650,N_19213,N_19271);
xor U19651 (N_19651,N_19219,N_19377);
xnor U19652 (N_19652,N_19417,N_19473);
nand U19653 (N_19653,N_19208,N_19257);
nand U19654 (N_19654,N_19575,N_19412);
nand U19655 (N_19655,N_19446,N_19483);
nand U19656 (N_19656,N_19291,N_19400);
nor U19657 (N_19657,N_19474,N_19476);
nor U19658 (N_19658,N_19551,N_19587);
or U19659 (N_19659,N_19590,N_19589);
and U19660 (N_19660,N_19513,N_19457);
xor U19661 (N_19661,N_19463,N_19598);
xnor U19662 (N_19662,N_19409,N_19244);
xor U19663 (N_19663,N_19263,N_19329);
nor U19664 (N_19664,N_19382,N_19235);
xnor U19665 (N_19665,N_19466,N_19249);
nand U19666 (N_19666,N_19595,N_19325);
or U19667 (N_19667,N_19449,N_19231);
or U19668 (N_19668,N_19480,N_19443);
xnor U19669 (N_19669,N_19277,N_19341);
and U19670 (N_19670,N_19565,N_19251);
and U19671 (N_19671,N_19342,N_19335);
xor U19672 (N_19672,N_19396,N_19445);
or U19673 (N_19673,N_19541,N_19435);
nor U19674 (N_19674,N_19308,N_19258);
xor U19675 (N_19675,N_19403,N_19562);
nand U19676 (N_19676,N_19210,N_19532);
nand U19677 (N_19677,N_19475,N_19353);
and U19678 (N_19678,N_19497,N_19485);
nor U19679 (N_19679,N_19460,N_19310);
or U19680 (N_19680,N_19202,N_19242);
and U19681 (N_19681,N_19205,N_19274);
or U19682 (N_19682,N_19366,N_19509);
xor U19683 (N_19683,N_19356,N_19348);
nor U19684 (N_19684,N_19599,N_19461);
nor U19685 (N_19685,N_19370,N_19594);
and U19686 (N_19686,N_19393,N_19447);
or U19687 (N_19687,N_19593,N_19442);
or U19688 (N_19688,N_19266,N_19596);
and U19689 (N_19689,N_19292,N_19336);
xor U19690 (N_19690,N_19468,N_19286);
and U19691 (N_19691,N_19577,N_19214);
xnor U19692 (N_19692,N_19499,N_19334);
and U19693 (N_19693,N_19471,N_19279);
and U19694 (N_19694,N_19217,N_19554);
nand U19695 (N_19695,N_19518,N_19472);
xor U19696 (N_19696,N_19451,N_19585);
xnor U19697 (N_19697,N_19455,N_19318);
xor U19698 (N_19698,N_19424,N_19211);
and U19699 (N_19699,N_19507,N_19302);
or U19700 (N_19700,N_19421,N_19265);
and U19701 (N_19701,N_19317,N_19324);
or U19702 (N_19702,N_19416,N_19394);
xnor U19703 (N_19703,N_19492,N_19367);
or U19704 (N_19704,N_19395,N_19220);
nor U19705 (N_19705,N_19536,N_19289);
or U19706 (N_19706,N_19444,N_19544);
xnor U19707 (N_19707,N_19203,N_19303);
and U19708 (N_19708,N_19458,N_19384);
nor U19709 (N_19709,N_19246,N_19307);
xnor U19710 (N_19710,N_19523,N_19224);
or U19711 (N_19711,N_19326,N_19273);
xnor U19712 (N_19712,N_19305,N_19557);
nor U19713 (N_19713,N_19520,N_19230);
nor U19714 (N_19714,N_19448,N_19301);
nor U19715 (N_19715,N_19254,N_19262);
or U19716 (N_19716,N_19269,N_19365);
nor U19717 (N_19717,N_19579,N_19383);
or U19718 (N_19718,N_19375,N_19354);
and U19719 (N_19719,N_19243,N_19559);
and U19720 (N_19720,N_19470,N_19592);
nor U19721 (N_19721,N_19250,N_19320);
or U19722 (N_19722,N_19293,N_19322);
nand U19723 (N_19723,N_19515,N_19432);
xor U19724 (N_19724,N_19545,N_19331);
nor U19725 (N_19725,N_19478,N_19363);
nand U19726 (N_19726,N_19498,N_19268);
xor U19727 (N_19727,N_19410,N_19398);
and U19728 (N_19728,N_19411,N_19201);
nand U19729 (N_19729,N_19389,N_19232);
nand U19730 (N_19730,N_19438,N_19297);
or U19731 (N_19731,N_19440,N_19391);
xor U19732 (N_19732,N_19436,N_19319);
xnor U19733 (N_19733,N_19212,N_19300);
or U19734 (N_19734,N_19309,N_19372);
nor U19735 (N_19735,N_19588,N_19431);
and U19736 (N_19736,N_19495,N_19540);
or U19737 (N_19737,N_19529,N_19204);
nand U19738 (N_19738,N_19526,N_19236);
nor U19739 (N_19739,N_19369,N_19314);
and U19740 (N_19740,N_19486,N_19405);
xor U19741 (N_19741,N_19477,N_19517);
nor U19742 (N_19742,N_19238,N_19527);
nor U19743 (N_19743,N_19299,N_19355);
xor U19744 (N_19744,N_19347,N_19259);
or U19745 (N_19745,N_19487,N_19456);
or U19746 (N_19746,N_19441,N_19226);
xor U19747 (N_19747,N_19344,N_19506);
nor U19748 (N_19748,N_19385,N_19543);
or U19749 (N_19749,N_19376,N_19553);
xnor U19750 (N_19750,N_19566,N_19578);
and U19751 (N_19751,N_19534,N_19586);
nand U19752 (N_19752,N_19418,N_19430);
and U19753 (N_19753,N_19399,N_19408);
xnor U19754 (N_19754,N_19287,N_19533);
xor U19755 (N_19755,N_19359,N_19295);
nor U19756 (N_19756,N_19240,N_19221);
and U19757 (N_19757,N_19275,N_19402);
nor U19758 (N_19758,N_19439,N_19558);
nor U19759 (N_19759,N_19390,N_19547);
nor U19760 (N_19760,N_19374,N_19222);
nor U19761 (N_19761,N_19237,N_19282);
or U19762 (N_19762,N_19488,N_19583);
xnor U19763 (N_19763,N_19584,N_19422);
xor U19764 (N_19764,N_19252,N_19581);
nor U19765 (N_19765,N_19255,N_19528);
xor U19766 (N_19766,N_19361,N_19502);
xor U19767 (N_19767,N_19484,N_19464);
nor U19768 (N_19768,N_19453,N_19351);
nand U19769 (N_19769,N_19315,N_19340);
or U19770 (N_19770,N_19514,N_19428);
nor U19771 (N_19771,N_19538,N_19570);
and U19772 (N_19772,N_19304,N_19426);
nand U19773 (N_19773,N_19358,N_19567);
xor U19774 (N_19774,N_19278,N_19524);
nor U19775 (N_19775,N_19427,N_19425);
and U19776 (N_19776,N_19387,N_19511);
or U19777 (N_19777,N_19494,N_19392);
nor U19778 (N_19778,N_19339,N_19298);
xnor U19779 (N_19779,N_19542,N_19284);
xor U19780 (N_19780,N_19504,N_19510);
nor U19781 (N_19781,N_19337,N_19332);
nor U19782 (N_19782,N_19378,N_19573);
nand U19783 (N_19783,N_19333,N_19233);
nor U19784 (N_19784,N_19323,N_19419);
nand U19785 (N_19785,N_19379,N_19572);
and U19786 (N_19786,N_19371,N_19469);
and U19787 (N_19787,N_19423,N_19413);
or U19788 (N_19788,N_19563,N_19350);
nand U19789 (N_19789,N_19253,N_19267);
or U19790 (N_19790,N_19516,N_19496);
or U19791 (N_19791,N_19482,N_19467);
nor U19792 (N_19792,N_19321,N_19283);
nand U19793 (N_19793,N_19270,N_19294);
nor U19794 (N_19794,N_19368,N_19569);
xnor U19795 (N_19795,N_19241,N_19345);
and U19796 (N_19796,N_19311,N_19530);
xnor U19797 (N_19797,N_19537,N_19519);
nand U19798 (N_19798,N_19434,N_19386);
and U19799 (N_19799,N_19489,N_19571);
and U19800 (N_19800,N_19580,N_19543);
or U19801 (N_19801,N_19245,N_19268);
and U19802 (N_19802,N_19501,N_19535);
or U19803 (N_19803,N_19459,N_19268);
xnor U19804 (N_19804,N_19523,N_19381);
and U19805 (N_19805,N_19273,N_19354);
nand U19806 (N_19806,N_19585,N_19345);
or U19807 (N_19807,N_19462,N_19585);
nor U19808 (N_19808,N_19296,N_19363);
and U19809 (N_19809,N_19233,N_19578);
nand U19810 (N_19810,N_19397,N_19592);
or U19811 (N_19811,N_19343,N_19275);
nand U19812 (N_19812,N_19595,N_19319);
nand U19813 (N_19813,N_19471,N_19343);
or U19814 (N_19814,N_19411,N_19382);
or U19815 (N_19815,N_19475,N_19238);
xor U19816 (N_19816,N_19369,N_19502);
and U19817 (N_19817,N_19322,N_19383);
or U19818 (N_19818,N_19563,N_19528);
and U19819 (N_19819,N_19404,N_19502);
nand U19820 (N_19820,N_19478,N_19243);
and U19821 (N_19821,N_19405,N_19503);
xnor U19822 (N_19822,N_19470,N_19430);
nand U19823 (N_19823,N_19505,N_19475);
nor U19824 (N_19824,N_19422,N_19454);
nor U19825 (N_19825,N_19377,N_19239);
nand U19826 (N_19826,N_19509,N_19270);
nand U19827 (N_19827,N_19382,N_19259);
or U19828 (N_19828,N_19237,N_19580);
nand U19829 (N_19829,N_19291,N_19526);
nand U19830 (N_19830,N_19264,N_19320);
nor U19831 (N_19831,N_19530,N_19211);
xor U19832 (N_19832,N_19406,N_19557);
xor U19833 (N_19833,N_19566,N_19426);
and U19834 (N_19834,N_19335,N_19451);
or U19835 (N_19835,N_19432,N_19484);
nor U19836 (N_19836,N_19563,N_19426);
nor U19837 (N_19837,N_19234,N_19350);
or U19838 (N_19838,N_19593,N_19359);
nand U19839 (N_19839,N_19315,N_19532);
nand U19840 (N_19840,N_19399,N_19357);
xnor U19841 (N_19841,N_19419,N_19224);
or U19842 (N_19842,N_19395,N_19504);
and U19843 (N_19843,N_19362,N_19536);
xor U19844 (N_19844,N_19475,N_19498);
xor U19845 (N_19845,N_19318,N_19434);
or U19846 (N_19846,N_19428,N_19227);
xor U19847 (N_19847,N_19467,N_19280);
or U19848 (N_19848,N_19200,N_19337);
nand U19849 (N_19849,N_19274,N_19466);
xor U19850 (N_19850,N_19365,N_19278);
and U19851 (N_19851,N_19239,N_19533);
nand U19852 (N_19852,N_19307,N_19430);
or U19853 (N_19853,N_19345,N_19253);
xor U19854 (N_19854,N_19357,N_19213);
and U19855 (N_19855,N_19427,N_19376);
nor U19856 (N_19856,N_19547,N_19326);
xnor U19857 (N_19857,N_19438,N_19291);
nand U19858 (N_19858,N_19488,N_19572);
and U19859 (N_19859,N_19354,N_19551);
or U19860 (N_19860,N_19475,N_19347);
and U19861 (N_19861,N_19521,N_19432);
nor U19862 (N_19862,N_19513,N_19406);
xnor U19863 (N_19863,N_19311,N_19422);
xor U19864 (N_19864,N_19244,N_19230);
or U19865 (N_19865,N_19488,N_19304);
nand U19866 (N_19866,N_19308,N_19572);
xor U19867 (N_19867,N_19467,N_19236);
nor U19868 (N_19868,N_19333,N_19501);
xnor U19869 (N_19869,N_19435,N_19342);
and U19870 (N_19870,N_19313,N_19318);
xnor U19871 (N_19871,N_19503,N_19378);
nand U19872 (N_19872,N_19317,N_19499);
xnor U19873 (N_19873,N_19460,N_19554);
and U19874 (N_19874,N_19391,N_19414);
nor U19875 (N_19875,N_19498,N_19335);
xor U19876 (N_19876,N_19238,N_19331);
and U19877 (N_19877,N_19568,N_19496);
and U19878 (N_19878,N_19483,N_19207);
xnor U19879 (N_19879,N_19508,N_19576);
xnor U19880 (N_19880,N_19421,N_19290);
nor U19881 (N_19881,N_19382,N_19229);
nor U19882 (N_19882,N_19420,N_19393);
xor U19883 (N_19883,N_19530,N_19231);
and U19884 (N_19884,N_19553,N_19463);
nand U19885 (N_19885,N_19409,N_19591);
or U19886 (N_19886,N_19536,N_19434);
and U19887 (N_19887,N_19592,N_19529);
nand U19888 (N_19888,N_19222,N_19204);
and U19889 (N_19889,N_19506,N_19372);
xnor U19890 (N_19890,N_19463,N_19239);
and U19891 (N_19891,N_19571,N_19419);
and U19892 (N_19892,N_19233,N_19398);
nand U19893 (N_19893,N_19267,N_19314);
nand U19894 (N_19894,N_19528,N_19217);
and U19895 (N_19895,N_19265,N_19441);
or U19896 (N_19896,N_19561,N_19297);
xnor U19897 (N_19897,N_19421,N_19255);
xnor U19898 (N_19898,N_19419,N_19424);
xnor U19899 (N_19899,N_19487,N_19256);
xnor U19900 (N_19900,N_19410,N_19241);
nand U19901 (N_19901,N_19510,N_19397);
nor U19902 (N_19902,N_19533,N_19549);
nor U19903 (N_19903,N_19477,N_19430);
nand U19904 (N_19904,N_19267,N_19537);
and U19905 (N_19905,N_19321,N_19270);
nor U19906 (N_19906,N_19317,N_19503);
or U19907 (N_19907,N_19455,N_19590);
or U19908 (N_19908,N_19351,N_19554);
xor U19909 (N_19909,N_19338,N_19275);
nor U19910 (N_19910,N_19308,N_19335);
and U19911 (N_19911,N_19584,N_19341);
nor U19912 (N_19912,N_19399,N_19229);
and U19913 (N_19913,N_19229,N_19266);
xor U19914 (N_19914,N_19458,N_19354);
and U19915 (N_19915,N_19355,N_19360);
nor U19916 (N_19916,N_19491,N_19315);
and U19917 (N_19917,N_19570,N_19467);
xnor U19918 (N_19918,N_19492,N_19414);
and U19919 (N_19919,N_19269,N_19296);
nor U19920 (N_19920,N_19339,N_19567);
or U19921 (N_19921,N_19214,N_19280);
nand U19922 (N_19922,N_19417,N_19423);
and U19923 (N_19923,N_19441,N_19525);
nand U19924 (N_19924,N_19472,N_19560);
and U19925 (N_19925,N_19317,N_19286);
or U19926 (N_19926,N_19262,N_19386);
nor U19927 (N_19927,N_19482,N_19201);
or U19928 (N_19928,N_19513,N_19242);
nor U19929 (N_19929,N_19223,N_19222);
xor U19930 (N_19930,N_19560,N_19274);
nand U19931 (N_19931,N_19427,N_19358);
nand U19932 (N_19932,N_19324,N_19238);
nor U19933 (N_19933,N_19278,N_19570);
or U19934 (N_19934,N_19288,N_19306);
or U19935 (N_19935,N_19429,N_19445);
nor U19936 (N_19936,N_19421,N_19526);
or U19937 (N_19937,N_19391,N_19516);
and U19938 (N_19938,N_19457,N_19431);
or U19939 (N_19939,N_19587,N_19360);
or U19940 (N_19940,N_19531,N_19468);
xnor U19941 (N_19941,N_19428,N_19581);
or U19942 (N_19942,N_19340,N_19382);
nand U19943 (N_19943,N_19344,N_19364);
xnor U19944 (N_19944,N_19458,N_19213);
and U19945 (N_19945,N_19510,N_19477);
and U19946 (N_19946,N_19344,N_19443);
xnor U19947 (N_19947,N_19516,N_19299);
xor U19948 (N_19948,N_19377,N_19388);
xnor U19949 (N_19949,N_19420,N_19286);
and U19950 (N_19950,N_19564,N_19203);
and U19951 (N_19951,N_19406,N_19389);
nor U19952 (N_19952,N_19432,N_19542);
nor U19953 (N_19953,N_19552,N_19447);
nor U19954 (N_19954,N_19505,N_19340);
or U19955 (N_19955,N_19570,N_19230);
nand U19956 (N_19956,N_19417,N_19318);
xnor U19957 (N_19957,N_19319,N_19520);
or U19958 (N_19958,N_19312,N_19585);
xnor U19959 (N_19959,N_19284,N_19340);
or U19960 (N_19960,N_19438,N_19203);
or U19961 (N_19961,N_19205,N_19285);
and U19962 (N_19962,N_19253,N_19255);
nor U19963 (N_19963,N_19218,N_19296);
or U19964 (N_19964,N_19447,N_19389);
and U19965 (N_19965,N_19497,N_19472);
xnor U19966 (N_19966,N_19388,N_19518);
and U19967 (N_19967,N_19426,N_19447);
nand U19968 (N_19968,N_19451,N_19565);
and U19969 (N_19969,N_19425,N_19588);
nand U19970 (N_19970,N_19244,N_19463);
nand U19971 (N_19971,N_19507,N_19295);
nor U19972 (N_19972,N_19595,N_19280);
and U19973 (N_19973,N_19358,N_19554);
nand U19974 (N_19974,N_19308,N_19295);
xnor U19975 (N_19975,N_19430,N_19473);
or U19976 (N_19976,N_19300,N_19220);
nand U19977 (N_19977,N_19334,N_19435);
nor U19978 (N_19978,N_19387,N_19479);
xor U19979 (N_19979,N_19296,N_19476);
or U19980 (N_19980,N_19445,N_19484);
and U19981 (N_19981,N_19375,N_19542);
and U19982 (N_19982,N_19287,N_19488);
nand U19983 (N_19983,N_19310,N_19211);
or U19984 (N_19984,N_19216,N_19545);
nor U19985 (N_19985,N_19248,N_19333);
nor U19986 (N_19986,N_19391,N_19275);
or U19987 (N_19987,N_19226,N_19208);
nand U19988 (N_19988,N_19342,N_19457);
and U19989 (N_19989,N_19562,N_19550);
or U19990 (N_19990,N_19257,N_19534);
and U19991 (N_19991,N_19360,N_19474);
or U19992 (N_19992,N_19577,N_19303);
nand U19993 (N_19993,N_19211,N_19359);
nor U19994 (N_19994,N_19531,N_19447);
nand U19995 (N_19995,N_19483,N_19448);
nand U19996 (N_19996,N_19569,N_19532);
and U19997 (N_19997,N_19455,N_19258);
and U19998 (N_19998,N_19592,N_19580);
and U19999 (N_19999,N_19465,N_19220);
nor UO_0 (O_0,N_19943,N_19703);
xor UO_1 (O_1,N_19882,N_19929);
nand UO_2 (O_2,N_19822,N_19836);
xor UO_3 (O_3,N_19958,N_19709);
or UO_4 (O_4,N_19831,N_19696);
or UO_5 (O_5,N_19897,N_19750);
xnor UO_6 (O_6,N_19772,N_19987);
nand UO_7 (O_7,N_19942,N_19994);
xor UO_8 (O_8,N_19634,N_19902);
xor UO_9 (O_9,N_19936,N_19900);
xnor UO_10 (O_10,N_19632,N_19635);
xnor UO_11 (O_11,N_19778,N_19601);
nor UO_12 (O_12,N_19931,N_19712);
nor UO_13 (O_13,N_19705,N_19957);
nor UO_14 (O_14,N_19913,N_19926);
and UO_15 (O_15,N_19797,N_19764);
or UO_16 (O_16,N_19690,N_19891);
nand UO_17 (O_17,N_19667,N_19768);
nor UO_18 (O_18,N_19780,N_19654);
and UO_19 (O_19,N_19606,N_19854);
nor UO_20 (O_20,N_19646,N_19684);
xor UO_21 (O_21,N_19815,N_19642);
or UO_22 (O_22,N_19748,N_19969);
or UO_23 (O_23,N_19842,N_19857);
and UO_24 (O_24,N_19906,N_19701);
or UO_25 (O_25,N_19614,N_19692);
nand UO_26 (O_26,N_19636,N_19977);
and UO_27 (O_27,N_19718,N_19885);
and UO_28 (O_28,N_19872,N_19860);
or UO_29 (O_29,N_19875,N_19964);
and UO_30 (O_30,N_19825,N_19617);
and UO_31 (O_31,N_19769,N_19742);
nand UO_32 (O_32,N_19674,N_19631);
and UO_33 (O_33,N_19826,N_19856);
xnor UO_34 (O_34,N_19736,N_19681);
or UO_35 (O_35,N_19791,N_19770);
nand UO_36 (O_36,N_19911,N_19615);
or UO_37 (O_37,N_19795,N_19814);
nand UO_38 (O_38,N_19616,N_19877);
nand UO_39 (O_39,N_19820,N_19671);
and UO_40 (O_40,N_19702,N_19980);
nand UO_41 (O_41,N_19811,N_19847);
nand UO_42 (O_42,N_19816,N_19727);
and UO_43 (O_43,N_19890,N_19801);
nor UO_44 (O_44,N_19894,N_19608);
and UO_45 (O_45,N_19868,N_19986);
or UO_46 (O_46,N_19630,N_19650);
and UO_47 (O_47,N_19638,N_19664);
xnor UO_48 (O_48,N_19939,N_19832);
nor UO_49 (O_49,N_19851,N_19922);
nor UO_50 (O_50,N_19715,N_19721);
nand UO_51 (O_51,N_19876,N_19659);
xor UO_52 (O_52,N_19898,N_19782);
and UO_53 (O_53,N_19951,N_19932);
and UO_54 (O_54,N_19962,N_19880);
xnor UO_55 (O_55,N_19907,N_19938);
nand UO_56 (O_56,N_19730,N_19657);
xor UO_57 (O_57,N_19903,N_19947);
xor UO_58 (O_58,N_19666,N_19817);
or UO_59 (O_59,N_19804,N_19949);
and UO_60 (O_60,N_19910,N_19798);
nand UO_61 (O_61,N_19746,N_19837);
xor UO_62 (O_62,N_19848,N_19744);
xnor UO_63 (O_63,N_19706,N_19724);
nor UO_64 (O_64,N_19774,N_19863);
nor UO_65 (O_65,N_19756,N_19800);
nor UO_66 (O_66,N_19629,N_19827);
xnor UO_67 (O_67,N_19895,N_19745);
nand UO_68 (O_68,N_19694,N_19934);
and UO_69 (O_69,N_19751,N_19766);
xnor UO_70 (O_70,N_19993,N_19807);
xor UO_71 (O_71,N_19669,N_19991);
or UO_72 (O_72,N_19940,N_19733);
xor UO_73 (O_73,N_19792,N_19767);
xnor UO_74 (O_74,N_19946,N_19653);
and UO_75 (O_75,N_19812,N_19786);
or UO_76 (O_76,N_19883,N_19641);
and UO_77 (O_77,N_19834,N_19651);
xor UO_78 (O_78,N_19693,N_19610);
xnor UO_79 (O_79,N_19723,N_19862);
and UO_80 (O_80,N_19983,N_19874);
nand UO_81 (O_81,N_19648,N_19725);
or UO_82 (O_82,N_19948,N_19968);
nor UO_83 (O_83,N_19867,N_19633);
nand UO_84 (O_84,N_19915,N_19870);
nand UO_85 (O_85,N_19680,N_19966);
nand UO_86 (O_86,N_19660,N_19916);
nand UO_87 (O_87,N_19652,N_19924);
nor UO_88 (O_88,N_19626,N_19810);
nand UO_89 (O_89,N_19708,N_19695);
and UO_90 (O_90,N_19805,N_19729);
or UO_91 (O_91,N_19689,N_19697);
and UO_92 (O_92,N_19789,N_19656);
xnor UO_93 (O_93,N_19661,N_19973);
or UO_94 (O_94,N_19989,N_19955);
nor UO_95 (O_95,N_19886,N_19873);
nand UO_96 (O_96,N_19981,N_19763);
nor UO_97 (O_97,N_19861,N_19784);
nor UO_98 (O_98,N_19719,N_19828);
nor UO_99 (O_99,N_19758,N_19979);
and UO_100 (O_100,N_19662,N_19893);
or UO_101 (O_101,N_19691,N_19665);
nand UO_102 (O_102,N_19609,N_19639);
and UO_103 (O_103,N_19707,N_19982);
xor UO_104 (O_104,N_19960,N_19686);
nor UO_105 (O_105,N_19749,N_19643);
and UO_106 (O_106,N_19622,N_19941);
or UO_107 (O_107,N_19850,N_19710);
or UO_108 (O_108,N_19761,N_19625);
or UO_109 (O_109,N_19704,N_19790);
or UO_110 (O_110,N_19624,N_19735);
nand UO_111 (O_111,N_19920,N_19794);
xnor UO_112 (O_112,N_19658,N_19732);
nand UO_113 (O_113,N_19846,N_19679);
xnor UO_114 (O_114,N_19602,N_19663);
nand UO_115 (O_115,N_19841,N_19688);
nand UO_116 (O_116,N_19967,N_19655);
nor UO_117 (O_117,N_19923,N_19714);
or UO_118 (O_118,N_19904,N_19912);
nand UO_119 (O_119,N_19621,N_19809);
and UO_120 (O_120,N_19963,N_19953);
nor UO_121 (O_121,N_19921,N_19728);
xor UO_122 (O_122,N_19781,N_19919);
nor UO_123 (O_123,N_19835,N_19859);
or UO_124 (O_124,N_19775,N_19858);
nor UO_125 (O_125,N_19866,N_19845);
and UO_126 (O_126,N_19914,N_19984);
nor UO_127 (O_127,N_19687,N_19881);
and UO_128 (O_128,N_19855,N_19699);
or UO_129 (O_129,N_19970,N_19788);
or UO_130 (O_130,N_19640,N_19716);
nand UO_131 (O_131,N_19765,N_19743);
nor UO_132 (O_132,N_19961,N_19773);
nand UO_133 (O_133,N_19779,N_19618);
xor UO_134 (O_134,N_19783,N_19647);
nor UO_135 (O_135,N_19829,N_19917);
or UO_136 (O_136,N_19678,N_19739);
nor UO_137 (O_137,N_19755,N_19600);
nand UO_138 (O_138,N_19677,N_19752);
nor UO_139 (O_139,N_19999,N_19711);
nor UO_140 (O_140,N_19759,N_19802);
and UO_141 (O_141,N_19933,N_19909);
or UO_142 (O_142,N_19889,N_19787);
or UO_143 (O_143,N_19685,N_19864);
nor UO_144 (O_144,N_19905,N_19908);
and UO_145 (O_145,N_19771,N_19888);
and UO_146 (O_146,N_19808,N_19734);
xnor UO_147 (O_147,N_19945,N_19887);
or UO_148 (O_148,N_19871,N_19760);
nand UO_149 (O_149,N_19720,N_19682);
nand UO_150 (O_150,N_19819,N_19777);
nand UO_151 (O_151,N_19965,N_19944);
nand UO_152 (O_152,N_19676,N_19813);
xnor UO_153 (O_153,N_19627,N_19731);
or UO_154 (O_154,N_19988,N_19896);
and UO_155 (O_155,N_19928,N_19853);
and UO_156 (O_156,N_19985,N_19918);
nor UO_157 (O_157,N_19603,N_19978);
nor UO_158 (O_158,N_19605,N_19722);
nor UO_159 (O_159,N_19952,N_19673);
or UO_160 (O_160,N_19806,N_19956);
and UO_161 (O_161,N_19762,N_19757);
xor UO_162 (O_162,N_19899,N_19972);
and UO_163 (O_163,N_19954,N_19830);
nand UO_164 (O_164,N_19878,N_19844);
nor UO_165 (O_165,N_19698,N_19869);
xor UO_166 (O_166,N_19628,N_19776);
and UO_167 (O_167,N_19753,N_19821);
xnor UO_168 (O_168,N_19996,N_19927);
and UO_169 (O_169,N_19607,N_19741);
or UO_170 (O_170,N_19747,N_19796);
xnor UO_171 (O_171,N_19738,N_19930);
nand UO_172 (O_172,N_19799,N_19726);
xor UO_173 (O_173,N_19740,N_19824);
nand UO_174 (O_174,N_19976,N_19839);
and UO_175 (O_175,N_19683,N_19700);
nand UO_176 (O_176,N_19713,N_19992);
xor UO_177 (O_177,N_19604,N_19884);
and UO_178 (O_178,N_19818,N_19998);
nand UO_179 (O_179,N_19612,N_19668);
nor UO_180 (O_180,N_19935,N_19754);
and UO_181 (O_181,N_19737,N_19974);
xor UO_182 (O_182,N_19971,N_19645);
nor UO_183 (O_183,N_19975,N_19623);
or UO_184 (O_184,N_19843,N_19959);
and UO_185 (O_185,N_19619,N_19879);
xnor UO_186 (O_186,N_19901,N_19644);
nand UO_187 (O_187,N_19995,N_19892);
nand UO_188 (O_188,N_19950,N_19675);
nor UO_189 (O_189,N_19840,N_19937);
nand UO_190 (O_190,N_19649,N_19613);
and UO_191 (O_191,N_19611,N_19865);
and UO_192 (O_192,N_19620,N_19852);
and UO_193 (O_193,N_19823,N_19833);
nand UO_194 (O_194,N_19717,N_19925);
nand UO_195 (O_195,N_19990,N_19670);
and UO_196 (O_196,N_19672,N_19785);
or UO_197 (O_197,N_19997,N_19793);
and UO_198 (O_198,N_19637,N_19838);
nor UO_199 (O_199,N_19803,N_19849);
nand UO_200 (O_200,N_19847,N_19788);
nand UO_201 (O_201,N_19640,N_19809);
nand UO_202 (O_202,N_19940,N_19620);
xnor UO_203 (O_203,N_19986,N_19880);
nand UO_204 (O_204,N_19877,N_19961);
and UO_205 (O_205,N_19622,N_19759);
nand UO_206 (O_206,N_19622,N_19724);
and UO_207 (O_207,N_19743,N_19721);
nand UO_208 (O_208,N_19731,N_19773);
nor UO_209 (O_209,N_19910,N_19894);
nor UO_210 (O_210,N_19616,N_19615);
xor UO_211 (O_211,N_19970,N_19627);
or UO_212 (O_212,N_19721,N_19629);
nand UO_213 (O_213,N_19712,N_19772);
or UO_214 (O_214,N_19887,N_19979);
and UO_215 (O_215,N_19828,N_19658);
nand UO_216 (O_216,N_19824,N_19988);
nand UO_217 (O_217,N_19718,N_19803);
and UO_218 (O_218,N_19683,N_19602);
nor UO_219 (O_219,N_19744,N_19926);
and UO_220 (O_220,N_19968,N_19986);
nor UO_221 (O_221,N_19964,N_19654);
nor UO_222 (O_222,N_19855,N_19771);
nand UO_223 (O_223,N_19885,N_19735);
xnor UO_224 (O_224,N_19813,N_19723);
xor UO_225 (O_225,N_19604,N_19754);
xnor UO_226 (O_226,N_19641,N_19832);
and UO_227 (O_227,N_19894,N_19700);
or UO_228 (O_228,N_19766,N_19907);
or UO_229 (O_229,N_19940,N_19821);
xnor UO_230 (O_230,N_19795,N_19825);
nand UO_231 (O_231,N_19856,N_19762);
or UO_232 (O_232,N_19677,N_19969);
and UO_233 (O_233,N_19798,N_19706);
or UO_234 (O_234,N_19759,N_19909);
and UO_235 (O_235,N_19661,N_19716);
xnor UO_236 (O_236,N_19967,N_19830);
nand UO_237 (O_237,N_19703,N_19701);
and UO_238 (O_238,N_19635,N_19946);
or UO_239 (O_239,N_19826,N_19635);
nor UO_240 (O_240,N_19751,N_19972);
nand UO_241 (O_241,N_19927,N_19651);
or UO_242 (O_242,N_19632,N_19659);
and UO_243 (O_243,N_19921,N_19672);
and UO_244 (O_244,N_19850,N_19936);
or UO_245 (O_245,N_19973,N_19948);
nor UO_246 (O_246,N_19802,N_19897);
nand UO_247 (O_247,N_19854,N_19963);
nor UO_248 (O_248,N_19945,N_19735);
or UO_249 (O_249,N_19739,N_19801);
or UO_250 (O_250,N_19936,N_19956);
or UO_251 (O_251,N_19648,N_19763);
xor UO_252 (O_252,N_19718,N_19678);
nand UO_253 (O_253,N_19850,N_19810);
and UO_254 (O_254,N_19926,N_19845);
nand UO_255 (O_255,N_19861,N_19652);
and UO_256 (O_256,N_19830,N_19626);
xnor UO_257 (O_257,N_19992,N_19683);
xnor UO_258 (O_258,N_19723,N_19729);
or UO_259 (O_259,N_19857,N_19872);
nand UO_260 (O_260,N_19791,N_19859);
or UO_261 (O_261,N_19620,N_19986);
xor UO_262 (O_262,N_19656,N_19611);
and UO_263 (O_263,N_19930,N_19974);
nor UO_264 (O_264,N_19633,N_19681);
xnor UO_265 (O_265,N_19906,N_19870);
or UO_266 (O_266,N_19682,N_19725);
xor UO_267 (O_267,N_19674,N_19898);
or UO_268 (O_268,N_19908,N_19812);
xnor UO_269 (O_269,N_19963,N_19603);
nor UO_270 (O_270,N_19741,N_19805);
or UO_271 (O_271,N_19911,N_19870);
and UO_272 (O_272,N_19882,N_19751);
xor UO_273 (O_273,N_19863,N_19745);
xor UO_274 (O_274,N_19607,N_19617);
and UO_275 (O_275,N_19720,N_19702);
nand UO_276 (O_276,N_19982,N_19895);
or UO_277 (O_277,N_19690,N_19799);
or UO_278 (O_278,N_19634,N_19853);
nand UO_279 (O_279,N_19642,N_19773);
or UO_280 (O_280,N_19956,N_19837);
xnor UO_281 (O_281,N_19830,N_19997);
nand UO_282 (O_282,N_19781,N_19984);
nand UO_283 (O_283,N_19983,N_19924);
xor UO_284 (O_284,N_19907,N_19651);
or UO_285 (O_285,N_19634,N_19956);
nand UO_286 (O_286,N_19869,N_19736);
or UO_287 (O_287,N_19970,N_19734);
xor UO_288 (O_288,N_19942,N_19765);
xor UO_289 (O_289,N_19812,N_19792);
and UO_290 (O_290,N_19677,N_19726);
or UO_291 (O_291,N_19880,N_19864);
and UO_292 (O_292,N_19617,N_19742);
nand UO_293 (O_293,N_19826,N_19622);
nor UO_294 (O_294,N_19688,N_19652);
nand UO_295 (O_295,N_19992,N_19759);
or UO_296 (O_296,N_19890,N_19932);
nand UO_297 (O_297,N_19635,N_19894);
nor UO_298 (O_298,N_19858,N_19887);
nand UO_299 (O_299,N_19991,N_19606);
nand UO_300 (O_300,N_19940,N_19866);
or UO_301 (O_301,N_19673,N_19662);
xnor UO_302 (O_302,N_19817,N_19975);
nand UO_303 (O_303,N_19697,N_19641);
xor UO_304 (O_304,N_19707,N_19862);
and UO_305 (O_305,N_19712,N_19647);
xnor UO_306 (O_306,N_19753,N_19948);
and UO_307 (O_307,N_19650,N_19826);
and UO_308 (O_308,N_19864,N_19993);
nor UO_309 (O_309,N_19997,N_19876);
and UO_310 (O_310,N_19980,N_19808);
and UO_311 (O_311,N_19873,N_19769);
nand UO_312 (O_312,N_19799,N_19745);
or UO_313 (O_313,N_19922,N_19752);
and UO_314 (O_314,N_19943,N_19826);
or UO_315 (O_315,N_19687,N_19777);
and UO_316 (O_316,N_19956,N_19942);
or UO_317 (O_317,N_19874,N_19662);
nor UO_318 (O_318,N_19649,N_19699);
or UO_319 (O_319,N_19960,N_19725);
and UO_320 (O_320,N_19862,N_19950);
xnor UO_321 (O_321,N_19678,N_19860);
nor UO_322 (O_322,N_19608,N_19789);
or UO_323 (O_323,N_19913,N_19677);
and UO_324 (O_324,N_19855,N_19656);
xnor UO_325 (O_325,N_19986,N_19812);
nand UO_326 (O_326,N_19712,N_19859);
nor UO_327 (O_327,N_19748,N_19956);
nor UO_328 (O_328,N_19847,N_19754);
or UO_329 (O_329,N_19879,N_19951);
and UO_330 (O_330,N_19782,N_19690);
and UO_331 (O_331,N_19991,N_19747);
nand UO_332 (O_332,N_19789,N_19745);
or UO_333 (O_333,N_19887,N_19913);
and UO_334 (O_334,N_19914,N_19838);
or UO_335 (O_335,N_19744,N_19804);
nor UO_336 (O_336,N_19948,N_19877);
or UO_337 (O_337,N_19987,N_19767);
xor UO_338 (O_338,N_19882,N_19910);
nand UO_339 (O_339,N_19724,N_19950);
or UO_340 (O_340,N_19717,N_19961);
nor UO_341 (O_341,N_19968,N_19913);
nor UO_342 (O_342,N_19985,N_19700);
nor UO_343 (O_343,N_19802,N_19622);
or UO_344 (O_344,N_19697,N_19979);
xnor UO_345 (O_345,N_19645,N_19740);
xnor UO_346 (O_346,N_19642,N_19703);
or UO_347 (O_347,N_19830,N_19853);
and UO_348 (O_348,N_19933,N_19736);
nand UO_349 (O_349,N_19783,N_19635);
nand UO_350 (O_350,N_19905,N_19727);
xnor UO_351 (O_351,N_19673,N_19760);
and UO_352 (O_352,N_19771,N_19978);
xor UO_353 (O_353,N_19696,N_19822);
xnor UO_354 (O_354,N_19860,N_19788);
xnor UO_355 (O_355,N_19979,N_19878);
and UO_356 (O_356,N_19949,N_19945);
and UO_357 (O_357,N_19852,N_19899);
xor UO_358 (O_358,N_19850,N_19932);
or UO_359 (O_359,N_19899,N_19978);
nand UO_360 (O_360,N_19635,N_19623);
xnor UO_361 (O_361,N_19994,N_19812);
xnor UO_362 (O_362,N_19808,N_19923);
and UO_363 (O_363,N_19875,N_19739);
xnor UO_364 (O_364,N_19834,N_19650);
or UO_365 (O_365,N_19887,N_19695);
xor UO_366 (O_366,N_19884,N_19711);
and UO_367 (O_367,N_19793,N_19794);
nor UO_368 (O_368,N_19612,N_19840);
and UO_369 (O_369,N_19688,N_19638);
and UO_370 (O_370,N_19670,N_19836);
and UO_371 (O_371,N_19859,N_19932);
xor UO_372 (O_372,N_19998,N_19903);
or UO_373 (O_373,N_19723,N_19710);
and UO_374 (O_374,N_19666,N_19988);
and UO_375 (O_375,N_19977,N_19728);
and UO_376 (O_376,N_19792,N_19834);
nor UO_377 (O_377,N_19604,N_19779);
xor UO_378 (O_378,N_19921,N_19851);
xor UO_379 (O_379,N_19971,N_19707);
or UO_380 (O_380,N_19638,N_19883);
xnor UO_381 (O_381,N_19795,N_19848);
xnor UO_382 (O_382,N_19697,N_19790);
nand UO_383 (O_383,N_19869,N_19849);
nand UO_384 (O_384,N_19740,N_19901);
nand UO_385 (O_385,N_19849,N_19816);
and UO_386 (O_386,N_19688,N_19777);
or UO_387 (O_387,N_19716,N_19852);
or UO_388 (O_388,N_19847,N_19692);
xnor UO_389 (O_389,N_19905,N_19873);
or UO_390 (O_390,N_19956,N_19702);
nor UO_391 (O_391,N_19883,N_19973);
or UO_392 (O_392,N_19844,N_19944);
nor UO_393 (O_393,N_19721,N_19930);
or UO_394 (O_394,N_19759,N_19692);
and UO_395 (O_395,N_19678,N_19909);
nor UO_396 (O_396,N_19852,N_19611);
and UO_397 (O_397,N_19883,N_19834);
xnor UO_398 (O_398,N_19794,N_19632);
xor UO_399 (O_399,N_19754,N_19902);
nand UO_400 (O_400,N_19881,N_19605);
nand UO_401 (O_401,N_19736,N_19804);
nor UO_402 (O_402,N_19731,N_19640);
nor UO_403 (O_403,N_19923,N_19869);
and UO_404 (O_404,N_19882,N_19729);
and UO_405 (O_405,N_19633,N_19774);
nor UO_406 (O_406,N_19985,N_19685);
xor UO_407 (O_407,N_19626,N_19639);
nor UO_408 (O_408,N_19633,N_19750);
nor UO_409 (O_409,N_19928,N_19953);
nor UO_410 (O_410,N_19657,N_19637);
and UO_411 (O_411,N_19777,N_19743);
xor UO_412 (O_412,N_19603,N_19739);
xor UO_413 (O_413,N_19966,N_19733);
xnor UO_414 (O_414,N_19753,N_19931);
nor UO_415 (O_415,N_19904,N_19899);
and UO_416 (O_416,N_19867,N_19855);
xor UO_417 (O_417,N_19693,N_19791);
nor UO_418 (O_418,N_19625,N_19791);
nor UO_419 (O_419,N_19833,N_19683);
nor UO_420 (O_420,N_19826,N_19831);
or UO_421 (O_421,N_19621,N_19872);
xor UO_422 (O_422,N_19906,N_19856);
nand UO_423 (O_423,N_19981,N_19642);
and UO_424 (O_424,N_19794,N_19986);
and UO_425 (O_425,N_19618,N_19657);
or UO_426 (O_426,N_19731,N_19861);
or UO_427 (O_427,N_19891,N_19978);
nand UO_428 (O_428,N_19718,N_19816);
and UO_429 (O_429,N_19668,N_19952);
nor UO_430 (O_430,N_19710,N_19640);
xor UO_431 (O_431,N_19604,N_19944);
xnor UO_432 (O_432,N_19646,N_19839);
or UO_433 (O_433,N_19789,N_19901);
nor UO_434 (O_434,N_19793,N_19618);
or UO_435 (O_435,N_19659,N_19893);
xnor UO_436 (O_436,N_19838,N_19605);
nor UO_437 (O_437,N_19893,N_19646);
or UO_438 (O_438,N_19750,N_19802);
xor UO_439 (O_439,N_19667,N_19785);
nor UO_440 (O_440,N_19958,N_19634);
and UO_441 (O_441,N_19886,N_19806);
xor UO_442 (O_442,N_19658,N_19601);
nand UO_443 (O_443,N_19716,N_19873);
xor UO_444 (O_444,N_19662,N_19771);
nand UO_445 (O_445,N_19642,N_19963);
and UO_446 (O_446,N_19796,N_19693);
xor UO_447 (O_447,N_19962,N_19602);
and UO_448 (O_448,N_19787,N_19645);
nand UO_449 (O_449,N_19912,N_19922);
nand UO_450 (O_450,N_19619,N_19851);
xnor UO_451 (O_451,N_19924,N_19846);
xor UO_452 (O_452,N_19971,N_19860);
nand UO_453 (O_453,N_19960,N_19997);
nor UO_454 (O_454,N_19960,N_19878);
nor UO_455 (O_455,N_19880,N_19875);
or UO_456 (O_456,N_19920,N_19786);
xnor UO_457 (O_457,N_19836,N_19782);
nand UO_458 (O_458,N_19845,N_19912);
nor UO_459 (O_459,N_19844,N_19635);
and UO_460 (O_460,N_19999,N_19935);
and UO_461 (O_461,N_19697,N_19638);
xnor UO_462 (O_462,N_19771,N_19689);
nand UO_463 (O_463,N_19997,N_19777);
nand UO_464 (O_464,N_19787,N_19679);
xnor UO_465 (O_465,N_19711,N_19785);
or UO_466 (O_466,N_19900,N_19933);
xnor UO_467 (O_467,N_19728,N_19825);
nand UO_468 (O_468,N_19630,N_19938);
or UO_469 (O_469,N_19724,N_19816);
nand UO_470 (O_470,N_19609,N_19999);
xor UO_471 (O_471,N_19942,N_19880);
xor UO_472 (O_472,N_19786,N_19823);
nor UO_473 (O_473,N_19915,N_19649);
nand UO_474 (O_474,N_19915,N_19799);
and UO_475 (O_475,N_19919,N_19642);
nand UO_476 (O_476,N_19634,N_19730);
nand UO_477 (O_477,N_19939,N_19796);
xnor UO_478 (O_478,N_19631,N_19996);
nor UO_479 (O_479,N_19608,N_19936);
and UO_480 (O_480,N_19999,N_19922);
or UO_481 (O_481,N_19919,N_19818);
xnor UO_482 (O_482,N_19919,N_19856);
or UO_483 (O_483,N_19660,N_19649);
nand UO_484 (O_484,N_19927,N_19776);
and UO_485 (O_485,N_19991,N_19814);
nor UO_486 (O_486,N_19951,N_19608);
xor UO_487 (O_487,N_19763,N_19859);
nor UO_488 (O_488,N_19823,N_19728);
xnor UO_489 (O_489,N_19912,N_19658);
and UO_490 (O_490,N_19991,N_19804);
nand UO_491 (O_491,N_19975,N_19774);
nand UO_492 (O_492,N_19807,N_19963);
nand UO_493 (O_493,N_19672,N_19977);
xor UO_494 (O_494,N_19857,N_19897);
xnor UO_495 (O_495,N_19800,N_19896);
nand UO_496 (O_496,N_19753,N_19732);
and UO_497 (O_497,N_19615,N_19767);
nand UO_498 (O_498,N_19805,N_19899);
xnor UO_499 (O_499,N_19722,N_19695);
nor UO_500 (O_500,N_19807,N_19658);
or UO_501 (O_501,N_19678,N_19904);
xor UO_502 (O_502,N_19600,N_19737);
or UO_503 (O_503,N_19787,N_19750);
nand UO_504 (O_504,N_19684,N_19894);
nand UO_505 (O_505,N_19606,N_19696);
xnor UO_506 (O_506,N_19840,N_19644);
or UO_507 (O_507,N_19866,N_19776);
nand UO_508 (O_508,N_19691,N_19633);
nand UO_509 (O_509,N_19601,N_19685);
xnor UO_510 (O_510,N_19671,N_19799);
nor UO_511 (O_511,N_19646,N_19808);
and UO_512 (O_512,N_19861,N_19664);
xnor UO_513 (O_513,N_19743,N_19864);
xnor UO_514 (O_514,N_19864,N_19884);
and UO_515 (O_515,N_19992,N_19879);
nand UO_516 (O_516,N_19632,N_19997);
and UO_517 (O_517,N_19639,N_19620);
and UO_518 (O_518,N_19934,N_19841);
and UO_519 (O_519,N_19724,N_19964);
nand UO_520 (O_520,N_19816,N_19801);
xnor UO_521 (O_521,N_19602,N_19753);
nor UO_522 (O_522,N_19609,N_19992);
nand UO_523 (O_523,N_19884,N_19837);
nor UO_524 (O_524,N_19650,N_19718);
and UO_525 (O_525,N_19842,N_19880);
xor UO_526 (O_526,N_19979,N_19814);
and UO_527 (O_527,N_19860,N_19911);
xnor UO_528 (O_528,N_19769,N_19825);
nand UO_529 (O_529,N_19973,N_19674);
or UO_530 (O_530,N_19924,N_19765);
or UO_531 (O_531,N_19968,N_19833);
or UO_532 (O_532,N_19688,N_19966);
nor UO_533 (O_533,N_19967,N_19721);
xnor UO_534 (O_534,N_19695,N_19638);
nand UO_535 (O_535,N_19660,N_19668);
and UO_536 (O_536,N_19743,N_19719);
or UO_537 (O_537,N_19887,N_19867);
and UO_538 (O_538,N_19926,N_19742);
or UO_539 (O_539,N_19717,N_19795);
xor UO_540 (O_540,N_19720,N_19621);
and UO_541 (O_541,N_19880,N_19798);
nor UO_542 (O_542,N_19718,N_19826);
nand UO_543 (O_543,N_19798,N_19753);
nor UO_544 (O_544,N_19983,N_19940);
xor UO_545 (O_545,N_19775,N_19973);
nand UO_546 (O_546,N_19922,N_19834);
nand UO_547 (O_547,N_19976,N_19861);
or UO_548 (O_548,N_19672,N_19787);
nand UO_549 (O_549,N_19908,N_19791);
nand UO_550 (O_550,N_19877,N_19934);
nor UO_551 (O_551,N_19704,N_19908);
xor UO_552 (O_552,N_19905,N_19715);
and UO_553 (O_553,N_19811,N_19605);
or UO_554 (O_554,N_19635,N_19871);
or UO_555 (O_555,N_19788,N_19686);
nand UO_556 (O_556,N_19780,N_19981);
nand UO_557 (O_557,N_19714,N_19734);
and UO_558 (O_558,N_19807,N_19964);
and UO_559 (O_559,N_19625,N_19897);
nand UO_560 (O_560,N_19858,N_19894);
xnor UO_561 (O_561,N_19887,N_19707);
nor UO_562 (O_562,N_19976,N_19666);
or UO_563 (O_563,N_19934,N_19800);
nand UO_564 (O_564,N_19748,N_19699);
nor UO_565 (O_565,N_19816,N_19827);
and UO_566 (O_566,N_19772,N_19823);
and UO_567 (O_567,N_19871,N_19817);
nand UO_568 (O_568,N_19994,N_19947);
xor UO_569 (O_569,N_19827,N_19835);
and UO_570 (O_570,N_19611,N_19784);
and UO_571 (O_571,N_19798,N_19773);
or UO_572 (O_572,N_19915,N_19611);
nor UO_573 (O_573,N_19887,N_19619);
nand UO_574 (O_574,N_19731,N_19968);
xnor UO_575 (O_575,N_19658,N_19729);
xnor UO_576 (O_576,N_19707,N_19777);
and UO_577 (O_577,N_19600,N_19605);
nor UO_578 (O_578,N_19730,N_19971);
nand UO_579 (O_579,N_19704,N_19946);
nand UO_580 (O_580,N_19764,N_19798);
nand UO_581 (O_581,N_19982,N_19983);
nor UO_582 (O_582,N_19899,N_19686);
and UO_583 (O_583,N_19741,N_19957);
or UO_584 (O_584,N_19797,N_19721);
nor UO_585 (O_585,N_19782,N_19674);
nor UO_586 (O_586,N_19839,N_19698);
or UO_587 (O_587,N_19758,N_19775);
xor UO_588 (O_588,N_19747,N_19732);
nand UO_589 (O_589,N_19610,N_19711);
xnor UO_590 (O_590,N_19961,N_19930);
nor UO_591 (O_591,N_19841,N_19741);
xor UO_592 (O_592,N_19806,N_19951);
xnor UO_593 (O_593,N_19793,N_19839);
nand UO_594 (O_594,N_19984,N_19610);
xnor UO_595 (O_595,N_19896,N_19672);
nor UO_596 (O_596,N_19947,N_19852);
nor UO_597 (O_597,N_19979,N_19825);
and UO_598 (O_598,N_19706,N_19868);
xnor UO_599 (O_599,N_19718,N_19752);
or UO_600 (O_600,N_19957,N_19696);
or UO_601 (O_601,N_19684,N_19713);
nand UO_602 (O_602,N_19868,N_19850);
and UO_603 (O_603,N_19677,N_19672);
xor UO_604 (O_604,N_19996,N_19628);
nor UO_605 (O_605,N_19978,N_19929);
nor UO_606 (O_606,N_19615,N_19802);
xnor UO_607 (O_607,N_19881,N_19811);
nand UO_608 (O_608,N_19981,N_19618);
xor UO_609 (O_609,N_19838,N_19888);
nor UO_610 (O_610,N_19956,N_19692);
or UO_611 (O_611,N_19677,N_19681);
or UO_612 (O_612,N_19740,N_19910);
xnor UO_613 (O_613,N_19732,N_19620);
or UO_614 (O_614,N_19833,N_19631);
or UO_615 (O_615,N_19670,N_19610);
nor UO_616 (O_616,N_19608,N_19645);
nor UO_617 (O_617,N_19619,N_19630);
xor UO_618 (O_618,N_19756,N_19703);
and UO_619 (O_619,N_19801,N_19609);
and UO_620 (O_620,N_19950,N_19996);
nand UO_621 (O_621,N_19701,N_19870);
nor UO_622 (O_622,N_19666,N_19634);
or UO_623 (O_623,N_19823,N_19656);
nand UO_624 (O_624,N_19932,N_19991);
and UO_625 (O_625,N_19660,N_19707);
and UO_626 (O_626,N_19817,N_19797);
and UO_627 (O_627,N_19961,N_19952);
or UO_628 (O_628,N_19705,N_19952);
xor UO_629 (O_629,N_19735,N_19939);
xnor UO_630 (O_630,N_19851,N_19961);
nor UO_631 (O_631,N_19897,N_19986);
nor UO_632 (O_632,N_19995,N_19847);
nand UO_633 (O_633,N_19711,N_19871);
or UO_634 (O_634,N_19947,N_19735);
and UO_635 (O_635,N_19827,N_19730);
or UO_636 (O_636,N_19652,N_19610);
or UO_637 (O_637,N_19858,N_19829);
nand UO_638 (O_638,N_19610,N_19836);
xor UO_639 (O_639,N_19776,N_19609);
or UO_640 (O_640,N_19820,N_19773);
xor UO_641 (O_641,N_19942,N_19890);
and UO_642 (O_642,N_19940,N_19868);
and UO_643 (O_643,N_19908,N_19967);
and UO_644 (O_644,N_19885,N_19715);
and UO_645 (O_645,N_19803,N_19955);
nor UO_646 (O_646,N_19929,N_19851);
nor UO_647 (O_647,N_19840,N_19676);
or UO_648 (O_648,N_19744,N_19688);
and UO_649 (O_649,N_19885,N_19936);
and UO_650 (O_650,N_19923,N_19997);
or UO_651 (O_651,N_19910,N_19917);
nand UO_652 (O_652,N_19611,N_19646);
or UO_653 (O_653,N_19657,N_19773);
and UO_654 (O_654,N_19650,N_19913);
and UO_655 (O_655,N_19709,N_19861);
nor UO_656 (O_656,N_19698,N_19783);
xnor UO_657 (O_657,N_19957,N_19970);
nor UO_658 (O_658,N_19640,N_19842);
nor UO_659 (O_659,N_19971,N_19979);
nand UO_660 (O_660,N_19763,N_19934);
nor UO_661 (O_661,N_19771,N_19646);
xnor UO_662 (O_662,N_19601,N_19924);
and UO_663 (O_663,N_19817,N_19901);
and UO_664 (O_664,N_19694,N_19856);
nand UO_665 (O_665,N_19725,N_19639);
xor UO_666 (O_666,N_19741,N_19792);
or UO_667 (O_667,N_19857,N_19657);
and UO_668 (O_668,N_19829,N_19777);
nand UO_669 (O_669,N_19741,N_19995);
nand UO_670 (O_670,N_19767,N_19878);
or UO_671 (O_671,N_19713,N_19709);
or UO_672 (O_672,N_19661,N_19669);
nand UO_673 (O_673,N_19625,N_19623);
and UO_674 (O_674,N_19802,N_19839);
or UO_675 (O_675,N_19879,N_19774);
nor UO_676 (O_676,N_19937,N_19891);
and UO_677 (O_677,N_19638,N_19992);
or UO_678 (O_678,N_19882,N_19968);
or UO_679 (O_679,N_19657,N_19959);
or UO_680 (O_680,N_19727,N_19808);
nand UO_681 (O_681,N_19691,N_19853);
nand UO_682 (O_682,N_19888,N_19783);
nor UO_683 (O_683,N_19950,N_19755);
and UO_684 (O_684,N_19962,N_19621);
or UO_685 (O_685,N_19618,N_19787);
xnor UO_686 (O_686,N_19991,N_19777);
or UO_687 (O_687,N_19970,N_19887);
nor UO_688 (O_688,N_19913,N_19875);
nand UO_689 (O_689,N_19607,N_19764);
nand UO_690 (O_690,N_19679,N_19788);
xor UO_691 (O_691,N_19654,N_19913);
nand UO_692 (O_692,N_19770,N_19746);
xor UO_693 (O_693,N_19630,N_19848);
or UO_694 (O_694,N_19981,N_19807);
nor UO_695 (O_695,N_19678,N_19720);
xnor UO_696 (O_696,N_19972,N_19789);
and UO_697 (O_697,N_19825,N_19743);
nand UO_698 (O_698,N_19897,N_19883);
or UO_699 (O_699,N_19756,N_19768);
and UO_700 (O_700,N_19648,N_19957);
or UO_701 (O_701,N_19724,N_19828);
xor UO_702 (O_702,N_19697,N_19840);
xor UO_703 (O_703,N_19807,N_19707);
nor UO_704 (O_704,N_19888,N_19884);
and UO_705 (O_705,N_19683,N_19919);
or UO_706 (O_706,N_19754,N_19738);
and UO_707 (O_707,N_19732,N_19774);
nand UO_708 (O_708,N_19695,N_19700);
and UO_709 (O_709,N_19606,N_19951);
xor UO_710 (O_710,N_19873,N_19707);
or UO_711 (O_711,N_19634,N_19901);
nand UO_712 (O_712,N_19636,N_19924);
nor UO_713 (O_713,N_19801,N_19842);
and UO_714 (O_714,N_19652,N_19639);
nand UO_715 (O_715,N_19749,N_19863);
nor UO_716 (O_716,N_19948,N_19934);
xor UO_717 (O_717,N_19612,N_19766);
xnor UO_718 (O_718,N_19840,N_19917);
and UO_719 (O_719,N_19741,N_19608);
nor UO_720 (O_720,N_19791,N_19613);
xnor UO_721 (O_721,N_19775,N_19997);
or UO_722 (O_722,N_19688,N_19771);
and UO_723 (O_723,N_19653,N_19839);
nand UO_724 (O_724,N_19659,N_19859);
nand UO_725 (O_725,N_19756,N_19864);
and UO_726 (O_726,N_19806,N_19675);
and UO_727 (O_727,N_19617,N_19814);
nand UO_728 (O_728,N_19823,N_19775);
and UO_729 (O_729,N_19733,N_19863);
nor UO_730 (O_730,N_19989,N_19685);
xnor UO_731 (O_731,N_19946,N_19668);
xor UO_732 (O_732,N_19713,N_19741);
or UO_733 (O_733,N_19894,N_19919);
nor UO_734 (O_734,N_19937,N_19907);
xnor UO_735 (O_735,N_19656,N_19913);
and UO_736 (O_736,N_19980,N_19930);
xnor UO_737 (O_737,N_19730,N_19650);
xor UO_738 (O_738,N_19817,N_19939);
nor UO_739 (O_739,N_19802,N_19992);
nor UO_740 (O_740,N_19735,N_19907);
and UO_741 (O_741,N_19672,N_19850);
and UO_742 (O_742,N_19939,N_19744);
or UO_743 (O_743,N_19625,N_19633);
nand UO_744 (O_744,N_19796,N_19854);
and UO_745 (O_745,N_19654,N_19704);
xor UO_746 (O_746,N_19685,N_19971);
or UO_747 (O_747,N_19768,N_19998);
xor UO_748 (O_748,N_19679,N_19606);
xor UO_749 (O_749,N_19777,N_19686);
xor UO_750 (O_750,N_19740,N_19770);
nor UO_751 (O_751,N_19973,N_19632);
and UO_752 (O_752,N_19950,N_19788);
and UO_753 (O_753,N_19899,N_19856);
nand UO_754 (O_754,N_19812,N_19839);
nand UO_755 (O_755,N_19625,N_19823);
nor UO_756 (O_756,N_19961,N_19968);
nor UO_757 (O_757,N_19958,N_19887);
xor UO_758 (O_758,N_19801,N_19724);
nand UO_759 (O_759,N_19659,N_19886);
xor UO_760 (O_760,N_19600,N_19850);
nor UO_761 (O_761,N_19705,N_19936);
xor UO_762 (O_762,N_19636,N_19821);
nor UO_763 (O_763,N_19607,N_19919);
or UO_764 (O_764,N_19896,N_19667);
and UO_765 (O_765,N_19985,N_19832);
or UO_766 (O_766,N_19737,N_19657);
nand UO_767 (O_767,N_19854,N_19802);
xnor UO_768 (O_768,N_19750,N_19801);
xnor UO_769 (O_769,N_19679,N_19651);
nand UO_770 (O_770,N_19755,N_19736);
or UO_771 (O_771,N_19684,N_19647);
nor UO_772 (O_772,N_19956,N_19861);
nand UO_773 (O_773,N_19929,N_19853);
or UO_774 (O_774,N_19927,N_19680);
nor UO_775 (O_775,N_19777,N_19932);
or UO_776 (O_776,N_19650,N_19726);
nand UO_777 (O_777,N_19691,N_19680);
or UO_778 (O_778,N_19633,N_19646);
nor UO_779 (O_779,N_19611,N_19760);
nand UO_780 (O_780,N_19963,N_19819);
nand UO_781 (O_781,N_19602,N_19775);
nand UO_782 (O_782,N_19870,N_19842);
nand UO_783 (O_783,N_19643,N_19786);
nor UO_784 (O_784,N_19720,N_19614);
or UO_785 (O_785,N_19613,N_19605);
or UO_786 (O_786,N_19903,N_19804);
nand UO_787 (O_787,N_19714,N_19944);
nor UO_788 (O_788,N_19847,N_19612);
nand UO_789 (O_789,N_19986,N_19982);
or UO_790 (O_790,N_19824,N_19878);
xor UO_791 (O_791,N_19876,N_19877);
and UO_792 (O_792,N_19672,N_19649);
and UO_793 (O_793,N_19795,N_19702);
or UO_794 (O_794,N_19943,N_19940);
xnor UO_795 (O_795,N_19734,N_19759);
xor UO_796 (O_796,N_19966,N_19804);
nor UO_797 (O_797,N_19654,N_19870);
nand UO_798 (O_798,N_19626,N_19651);
nor UO_799 (O_799,N_19895,N_19806);
xor UO_800 (O_800,N_19782,N_19607);
or UO_801 (O_801,N_19792,N_19619);
and UO_802 (O_802,N_19883,N_19857);
xor UO_803 (O_803,N_19991,N_19818);
or UO_804 (O_804,N_19632,N_19917);
nand UO_805 (O_805,N_19766,N_19666);
nand UO_806 (O_806,N_19617,N_19783);
and UO_807 (O_807,N_19695,N_19967);
xor UO_808 (O_808,N_19766,N_19937);
and UO_809 (O_809,N_19750,N_19828);
nor UO_810 (O_810,N_19684,N_19748);
xor UO_811 (O_811,N_19632,N_19937);
nor UO_812 (O_812,N_19971,N_19937);
or UO_813 (O_813,N_19691,N_19621);
xnor UO_814 (O_814,N_19981,N_19632);
and UO_815 (O_815,N_19930,N_19784);
or UO_816 (O_816,N_19943,N_19678);
or UO_817 (O_817,N_19708,N_19808);
and UO_818 (O_818,N_19809,N_19931);
or UO_819 (O_819,N_19893,N_19699);
nor UO_820 (O_820,N_19858,N_19697);
nor UO_821 (O_821,N_19901,N_19724);
nor UO_822 (O_822,N_19971,N_19772);
or UO_823 (O_823,N_19974,N_19727);
xor UO_824 (O_824,N_19902,N_19859);
or UO_825 (O_825,N_19777,N_19994);
or UO_826 (O_826,N_19623,N_19712);
nor UO_827 (O_827,N_19673,N_19924);
and UO_828 (O_828,N_19804,N_19615);
xor UO_829 (O_829,N_19857,N_19922);
nand UO_830 (O_830,N_19952,N_19793);
and UO_831 (O_831,N_19746,N_19931);
xor UO_832 (O_832,N_19990,N_19723);
xnor UO_833 (O_833,N_19658,N_19821);
nand UO_834 (O_834,N_19749,N_19993);
or UO_835 (O_835,N_19870,N_19967);
nand UO_836 (O_836,N_19766,N_19755);
and UO_837 (O_837,N_19785,N_19728);
or UO_838 (O_838,N_19741,N_19824);
and UO_839 (O_839,N_19983,N_19643);
xnor UO_840 (O_840,N_19810,N_19635);
xor UO_841 (O_841,N_19715,N_19882);
or UO_842 (O_842,N_19881,N_19979);
or UO_843 (O_843,N_19900,N_19643);
xnor UO_844 (O_844,N_19899,N_19983);
nand UO_845 (O_845,N_19724,N_19838);
nand UO_846 (O_846,N_19628,N_19650);
xor UO_847 (O_847,N_19626,N_19657);
nand UO_848 (O_848,N_19749,N_19702);
nor UO_849 (O_849,N_19900,N_19767);
and UO_850 (O_850,N_19648,N_19828);
nor UO_851 (O_851,N_19685,N_19953);
xnor UO_852 (O_852,N_19624,N_19649);
or UO_853 (O_853,N_19950,N_19930);
xor UO_854 (O_854,N_19860,N_19655);
or UO_855 (O_855,N_19773,N_19682);
nand UO_856 (O_856,N_19969,N_19627);
nor UO_857 (O_857,N_19638,N_19851);
or UO_858 (O_858,N_19926,N_19871);
nand UO_859 (O_859,N_19659,N_19948);
xor UO_860 (O_860,N_19884,N_19708);
nor UO_861 (O_861,N_19978,N_19751);
and UO_862 (O_862,N_19755,N_19687);
xnor UO_863 (O_863,N_19815,N_19998);
xor UO_864 (O_864,N_19731,N_19734);
nand UO_865 (O_865,N_19802,N_19650);
nand UO_866 (O_866,N_19967,N_19928);
xnor UO_867 (O_867,N_19863,N_19841);
nor UO_868 (O_868,N_19740,N_19943);
or UO_869 (O_869,N_19757,N_19780);
nor UO_870 (O_870,N_19805,N_19896);
and UO_871 (O_871,N_19744,N_19665);
nand UO_872 (O_872,N_19935,N_19873);
or UO_873 (O_873,N_19745,N_19991);
nor UO_874 (O_874,N_19926,N_19814);
nor UO_875 (O_875,N_19951,N_19861);
nand UO_876 (O_876,N_19888,N_19668);
or UO_877 (O_877,N_19837,N_19809);
xnor UO_878 (O_878,N_19689,N_19655);
xnor UO_879 (O_879,N_19797,N_19742);
and UO_880 (O_880,N_19729,N_19903);
nand UO_881 (O_881,N_19636,N_19960);
nor UO_882 (O_882,N_19643,N_19641);
xor UO_883 (O_883,N_19710,N_19965);
nor UO_884 (O_884,N_19642,N_19970);
nor UO_885 (O_885,N_19829,N_19790);
and UO_886 (O_886,N_19899,N_19703);
nor UO_887 (O_887,N_19906,N_19712);
or UO_888 (O_888,N_19957,N_19672);
nor UO_889 (O_889,N_19692,N_19712);
xnor UO_890 (O_890,N_19976,N_19943);
or UO_891 (O_891,N_19960,N_19632);
or UO_892 (O_892,N_19904,N_19718);
nor UO_893 (O_893,N_19722,N_19816);
or UO_894 (O_894,N_19698,N_19697);
nor UO_895 (O_895,N_19690,N_19931);
xnor UO_896 (O_896,N_19864,N_19840);
xor UO_897 (O_897,N_19778,N_19625);
nand UO_898 (O_898,N_19790,N_19777);
nor UO_899 (O_899,N_19945,N_19833);
and UO_900 (O_900,N_19686,N_19700);
or UO_901 (O_901,N_19945,N_19741);
nor UO_902 (O_902,N_19744,N_19783);
nand UO_903 (O_903,N_19692,N_19804);
and UO_904 (O_904,N_19714,N_19620);
xnor UO_905 (O_905,N_19962,N_19950);
nand UO_906 (O_906,N_19670,N_19804);
nand UO_907 (O_907,N_19761,N_19716);
and UO_908 (O_908,N_19712,N_19860);
nand UO_909 (O_909,N_19965,N_19963);
nor UO_910 (O_910,N_19944,N_19945);
nand UO_911 (O_911,N_19778,N_19793);
nand UO_912 (O_912,N_19889,N_19776);
and UO_913 (O_913,N_19614,N_19601);
xor UO_914 (O_914,N_19688,N_19976);
nand UO_915 (O_915,N_19615,N_19746);
or UO_916 (O_916,N_19671,N_19878);
nand UO_917 (O_917,N_19855,N_19643);
nor UO_918 (O_918,N_19789,N_19860);
nand UO_919 (O_919,N_19683,N_19934);
and UO_920 (O_920,N_19774,N_19631);
nor UO_921 (O_921,N_19630,N_19614);
and UO_922 (O_922,N_19655,N_19641);
nand UO_923 (O_923,N_19963,N_19772);
nor UO_924 (O_924,N_19891,N_19668);
nand UO_925 (O_925,N_19870,N_19934);
nand UO_926 (O_926,N_19930,N_19603);
or UO_927 (O_927,N_19813,N_19604);
nor UO_928 (O_928,N_19939,N_19903);
nand UO_929 (O_929,N_19778,N_19685);
and UO_930 (O_930,N_19900,N_19795);
and UO_931 (O_931,N_19630,N_19942);
and UO_932 (O_932,N_19874,N_19764);
nand UO_933 (O_933,N_19728,N_19886);
and UO_934 (O_934,N_19608,N_19643);
xnor UO_935 (O_935,N_19951,N_19771);
or UO_936 (O_936,N_19660,N_19918);
and UO_937 (O_937,N_19714,N_19658);
and UO_938 (O_938,N_19907,N_19883);
or UO_939 (O_939,N_19848,N_19867);
xnor UO_940 (O_940,N_19795,N_19913);
nand UO_941 (O_941,N_19657,N_19798);
and UO_942 (O_942,N_19848,N_19972);
or UO_943 (O_943,N_19669,N_19647);
nor UO_944 (O_944,N_19798,N_19830);
nand UO_945 (O_945,N_19928,N_19800);
and UO_946 (O_946,N_19979,N_19959);
xnor UO_947 (O_947,N_19718,N_19980);
nor UO_948 (O_948,N_19980,N_19664);
nor UO_949 (O_949,N_19955,N_19802);
nand UO_950 (O_950,N_19956,N_19973);
and UO_951 (O_951,N_19933,N_19906);
or UO_952 (O_952,N_19658,N_19809);
xor UO_953 (O_953,N_19783,N_19631);
nand UO_954 (O_954,N_19845,N_19857);
nand UO_955 (O_955,N_19990,N_19721);
nor UO_956 (O_956,N_19789,N_19856);
nand UO_957 (O_957,N_19765,N_19715);
and UO_958 (O_958,N_19739,N_19830);
nor UO_959 (O_959,N_19873,N_19693);
or UO_960 (O_960,N_19899,N_19661);
nor UO_961 (O_961,N_19708,N_19872);
or UO_962 (O_962,N_19688,N_19832);
nand UO_963 (O_963,N_19908,N_19876);
and UO_964 (O_964,N_19936,N_19988);
nand UO_965 (O_965,N_19842,N_19602);
or UO_966 (O_966,N_19649,N_19603);
nor UO_967 (O_967,N_19676,N_19939);
nor UO_968 (O_968,N_19715,N_19819);
or UO_969 (O_969,N_19875,N_19753);
xnor UO_970 (O_970,N_19876,N_19751);
nor UO_971 (O_971,N_19839,N_19875);
nor UO_972 (O_972,N_19764,N_19996);
xor UO_973 (O_973,N_19735,N_19799);
or UO_974 (O_974,N_19867,N_19922);
nand UO_975 (O_975,N_19766,N_19616);
nand UO_976 (O_976,N_19781,N_19887);
or UO_977 (O_977,N_19750,N_19954);
and UO_978 (O_978,N_19852,N_19767);
xor UO_979 (O_979,N_19639,N_19985);
xor UO_980 (O_980,N_19865,N_19879);
and UO_981 (O_981,N_19883,N_19809);
nor UO_982 (O_982,N_19807,N_19897);
and UO_983 (O_983,N_19782,N_19855);
or UO_984 (O_984,N_19673,N_19865);
or UO_985 (O_985,N_19715,N_19997);
nand UO_986 (O_986,N_19808,N_19699);
nor UO_987 (O_987,N_19825,N_19845);
and UO_988 (O_988,N_19946,N_19684);
nor UO_989 (O_989,N_19861,N_19857);
nand UO_990 (O_990,N_19877,N_19798);
xor UO_991 (O_991,N_19913,N_19836);
and UO_992 (O_992,N_19869,N_19872);
xnor UO_993 (O_993,N_19784,N_19723);
and UO_994 (O_994,N_19691,N_19953);
nand UO_995 (O_995,N_19682,N_19797);
nand UO_996 (O_996,N_19767,N_19962);
nor UO_997 (O_997,N_19917,N_19725);
and UO_998 (O_998,N_19842,N_19646);
and UO_999 (O_999,N_19696,N_19804);
nor UO_1000 (O_1000,N_19984,N_19863);
nor UO_1001 (O_1001,N_19759,N_19961);
and UO_1002 (O_1002,N_19601,N_19739);
nor UO_1003 (O_1003,N_19858,N_19734);
or UO_1004 (O_1004,N_19818,N_19959);
or UO_1005 (O_1005,N_19894,N_19870);
and UO_1006 (O_1006,N_19979,N_19696);
nor UO_1007 (O_1007,N_19698,N_19695);
and UO_1008 (O_1008,N_19945,N_19935);
nand UO_1009 (O_1009,N_19917,N_19967);
and UO_1010 (O_1010,N_19669,N_19876);
and UO_1011 (O_1011,N_19624,N_19858);
nand UO_1012 (O_1012,N_19963,N_19771);
and UO_1013 (O_1013,N_19959,N_19819);
nor UO_1014 (O_1014,N_19934,N_19909);
nor UO_1015 (O_1015,N_19772,N_19993);
and UO_1016 (O_1016,N_19744,N_19791);
nor UO_1017 (O_1017,N_19841,N_19759);
or UO_1018 (O_1018,N_19931,N_19631);
and UO_1019 (O_1019,N_19889,N_19742);
xor UO_1020 (O_1020,N_19856,N_19729);
nand UO_1021 (O_1021,N_19941,N_19714);
and UO_1022 (O_1022,N_19659,N_19683);
or UO_1023 (O_1023,N_19920,N_19965);
or UO_1024 (O_1024,N_19917,N_19669);
nand UO_1025 (O_1025,N_19829,N_19675);
nand UO_1026 (O_1026,N_19876,N_19921);
or UO_1027 (O_1027,N_19716,N_19692);
and UO_1028 (O_1028,N_19979,N_19822);
nor UO_1029 (O_1029,N_19600,N_19747);
nor UO_1030 (O_1030,N_19960,N_19875);
or UO_1031 (O_1031,N_19968,N_19969);
xnor UO_1032 (O_1032,N_19990,N_19766);
or UO_1033 (O_1033,N_19945,N_19897);
xnor UO_1034 (O_1034,N_19963,N_19793);
xnor UO_1035 (O_1035,N_19675,N_19947);
nor UO_1036 (O_1036,N_19934,N_19911);
nor UO_1037 (O_1037,N_19831,N_19844);
nor UO_1038 (O_1038,N_19621,N_19712);
or UO_1039 (O_1039,N_19757,N_19898);
or UO_1040 (O_1040,N_19993,N_19641);
or UO_1041 (O_1041,N_19789,N_19653);
nor UO_1042 (O_1042,N_19940,N_19784);
xnor UO_1043 (O_1043,N_19983,N_19813);
nor UO_1044 (O_1044,N_19721,N_19679);
xor UO_1045 (O_1045,N_19647,N_19985);
or UO_1046 (O_1046,N_19988,N_19831);
and UO_1047 (O_1047,N_19995,N_19766);
or UO_1048 (O_1048,N_19640,N_19826);
xnor UO_1049 (O_1049,N_19891,N_19783);
nor UO_1050 (O_1050,N_19854,N_19769);
or UO_1051 (O_1051,N_19742,N_19627);
xor UO_1052 (O_1052,N_19689,N_19610);
and UO_1053 (O_1053,N_19868,N_19774);
nand UO_1054 (O_1054,N_19884,N_19961);
nand UO_1055 (O_1055,N_19664,N_19961);
nand UO_1056 (O_1056,N_19879,N_19850);
and UO_1057 (O_1057,N_19722,N_19831);
xnor UO_1058 (O_1058,N_19748,N_19743);
nor UO_1059 (O_1059,N_19678,N_19777);
nor UO_1060 (O_1060,N_19681,N_19948);
xnor UO_1061 (O_1061,N_19642,N_19986);
xnor UO_1062 (O_1062,N_19787,N_19839);
xnor UO_1063 (O_1063,N_19881,N_19678);
nor UO_1064 (O_1064,N_19978,N_19956);
nand UO_1065 (O_1065,N_19776,N_19647);
xnor UO_1066 (O_1066,N_19932,N_19724);
nand UO_1067 (O_1067,N_19762,N_19837);
nand UO_1068 (O_1068,N_19833,N_19906);
nor UO_1069 (O_1069,N_19895,N_19738);
and UO_1070 (O_1070,N_19801,N_19644);
nor UO_1071 (O_1071,N_19680,N_19945);
nor UO_1072 (O_1072,N_19923,N_19959);
xor UO_1073 (O_1073,N_19943,N_19748);
xnor UO_1074 (O_1074,N_19838,N_19945);
and UO_1075 (O_1075,N_19839,N_19674);
and UO_1076 (O_1076,N_19762,N_19696);
xor UO_1077 (O_1077,N_19902,N_19673);
and UO_1078 (O_1078,N_19857,N_19948);
xor UO_1079 (O_1079,N_19914,N_19902);
nor UO_1080 (O_1080,N_19684,N_19988);
or UO_1081 (O_1081,N_19807,N_19823);
nand UO_1082 (O_1082,N_19705,N_19648);
xor UO_1083 (O_1083,N_19995,N_19695);
nand UO_1084 (O_1084,N_19855,N_19973);
nor UO_1085 (O_1085,N_19937,N_19719);
or UO_1086 (O_1086,N_19872,N_19881);
or UO_1087 (O_1087,N_19677,N_19731);
and UO_1088 (O_1088,N_19789,N_19774);
xor UO_1089 (O_1089,N_19891,N_19855);
and UO_1090 (O_1090,N_19985,N_19716);
and UO_1091 (O_1091,N_19968,N_19664);
or UO_1092 (O_1092,N_19777,N_19870);
or UO_1093 (O_1093,N_19891,N_19970);
nor UO_1094 (O_1094,N_19835,N_19760);
nor UO_1095 (O_1095,N_19756,N_19952);
and UO_1096 (O_1096,N_19897,N_19837);
or UO_1097 (O_1097,N_19736,N_19829);
xnor UO_1098 (O_1098,N_19825,N_19631);
nor UO_1099 (O_1099,N_19920,N_19789);
or UO_1100 (O_1100,N_19743,N_19664);
nand UO_1101 (O_1101,N_19692,N_19740);
nor UO_1102 (O_1102,N_19761,N_19754);
xnor UO_1103 (O_1103,N_19824,N_19853);
and UO_1104 (O_1104,N_19921,N_19954);
nand UO_1105 (O_1105,N_19818,N_19835);
or UO_1106 (O_1106,N_19831,N_19787);
nor UO_1107 (O_1107,N_19721,N_19793);
and UO_1108 (O_1108,N_19989,N_19678);
or UO_1109 (O_1109,N_19717,N_19865);
xnor UO_1110 (O_1110,N_19951,N_19691);
or UO_1111 (O_1111,N_19835,N_19783);
xnor UO_1112 (O_1112,N_19742,N_19998);
nor UO_1113 (O_1113,N_19657,N_19979);
nand UO_1114 (O_1114,N_19967,N_19907);
or UO_1115 (O_1115,N_19848,N_19691);
or UO_1116 (O_1116,N_19855,N_19691);
and UO_1117 (O_1117,N_19981,N_19932);
xnor UO_1118 (O_1118,N_19915,N_19694);
xnor UO_1119 (O_1119,N_19938,N_19767);
xnor UO_1120 (O_1120,N_19651,N_19719);
nand UO_1121 (O_1121,N_19624,N_19846);
and UO_1122 (O_1122,N_19790,N_19826);
nand UO_1123 (O_1123,N_19784,N_19988);
nand UO_1124 (O_1124,N_19905,N_19746);
and UO_1125 (O_1125,N_19923,N_19965);
nand UO_1126 (O_1126,N_19611,N_19790);
and UO_1127 (O_1127,N_19670,N_19664);
or UO_1128 (O_1128,N_19940,N_19679);
nand UO_1129 (O_1129,N_19772,N_19859);
nand UO_1130 (O_1130,N_19824,N_19629);
nand UO_1131 (O_1131,N_19995,N_19976);
and UO_1132 (O_1132,N_19819,N_19989);
and UO_1133 (O_1133,N_19686,N_19901);
and UO_1134 (O_1134,N_19703,N_19741);
and UO_1135 (O_1135,N_19994,N_19938);
and UO_1136 (O_1136,N_19955,N_19894);
and UO_1137 (O_1137,N_19695,N_19811);
and UO_1138 (O_1138,N_19780,N_19735);
and UO_1139 (O_1139,N_19725,N_19830);
nor UO_1140 (O_1140,N_19983,N_19969);
nand UO_1141 (O_1141,N_19907,N_19692);
nor UO_1142 (O_1142,N_19858,N_19946);
nor UO_1143 (O_1143,N_19881,N_19922);
or UO_1144 (O_1144,N_19879,N_19837);
xor UO_1145 (O_1145,N_19888,N_19687);
nor UO_1146 (O_1146,N_19673,N_19797);
nor UO_1147 (O_1147,N_19730,N_19669);
and UO_1148 (O_1148,N_19777,N_19861);
nor UO_1149 (O_1149,N_19760,N_19894);
nor UO_1150 (O_1150,N_19869,N_19784);
and UO_1151 (O_1151,N_19763,N_19809);
or UO_1152 (O_1152,N_19927,N_19691);
nand UO_1153 (O_1153,N_19757,N_19638);
xnor UO_1154 (O_1154,N_19834,N_19866);
or UO_1155 (O_1155,N_19907,N_19993);
or UO_1156 (O_1156,N_19656,N_19963);
nand UO_1157 (O_1157,N_19876,N_19736);
nor UO_1158 (O_1158,N_19974,N_19934);
xor UO_1159 (O_1159,N_19976,N_19733);
and UO_1160 (O_1160,N_19987,N_19736);
xnor UO_1161 (O_1161,N_19927,N_19797);
nor UO_1162 (O_1162,N_19667,N_19817);
or UO_1163 (O_1163,N_19928,N_19923);
nor UO_1164 (O_1164,N_19762,N_19606);
and UO_1165 (O_1165,N_19747,N_19969);
or UO_1166 (O_1166,N_19839,N_19835);
nand UO_1167 (O_1167,N_19953,N_19997);
nor UO_1168 (O_1168,N_19761,N_19628);
xor UO_1169 (O_1169,N_19693,N_19624);
nand UO_1170 (O_1170,N_19879,N_19648);
nor UO_1171 (O_1171,N_19678,N_19976);
nand UO_1172 (O_1172,N_19764,N_19613);
xnor UO_1173 (O_1173,N_19644,N_19643);
nor UO_1174 (O_1174,N_19753,N_19825);
nor UO_1175 (O_1175,N_19810,N_19676);
nor UO_1176 (O_1176,N_19654,N_19644);
nor UO_1177 (O_1177,N_19684,N_19678);
xnor UO_1178 (O_1178,N_19618,N_19799);
nor UO_1179 (O_1179,N_19777,N_19781);
xnor UO_1180 (O_1180,N_19968,N_19632);
and UO_1181 (O_1181,N_19683,N_19898);
nor UO_1182 (O_1182,N_19729,N_19864);
nand UO_1183 (O_1183,N_19876,N_19992);
nand UO_1184 (O_1184,N_19934,N_19805);
nand UO_1185 (O_1185,N_19629,N_19939);
xor UO_1186 (O_1186,N_19776,N_19741);
or UO_1187 (O_1187,N_19803,N_19712);
xnor UO_1188 (O_1188,N_19850,N_19984);
xor UO_1189 (O_1189,N_19607,N_19843);
xor UO_1190 (O_1190,N_19932,N_19999);
or UO_1191 (O_1191,N_19929,N_19969);
nor UO_1192 (O_1192,N_19794,N_19826);
and UO_1193 (O_1193,N_19923,N_19613);
nor UO_1194 (O_1194,N_19832,N_19798);
nand UO_1195 (O_1195,N_19914,N_19621);
nand UO_1196 (O_1196,N_19873,N_19676);
or UO_1197 (O_1197,N_19864,N_19690);
and UO_1198 (O_1198,N_19908,N_19958);
or UO_1199 (O_1199,N_19923,N_19849);
and UO_1200 (O_1200,N_19994,N_19646);
or UO_1201 (O_1201,N_19935,N_19748);
nor UO_1202 (O_1202,N_19732,N_19919);
and UO_1203 (O_1203,N_19760,N_19771);
nand UO_1204 (O_1204,N_19693,N_19652);
xor UO_1205 (O_1205,N_19798,N_19950);
nor UO_1206 (O_1206,N_19997,N_19739);
and UO_1207 (O_1207,N_19655,N_19885);
and UO_1208 (O_1208,N_19835,N_19697);
or UO_1209 (O_1209,N_19669,N_19955);
nand UO_1210 (O_1210,N_19974,N_19917);
nand UO_1211 (O_1211,N_19818,N_19852);
or UO_1212 (O_1212,N_19902,N_19644);
or UO_1213 (O_1213,N_19716,N_19648);
xor UO_1214 (O_1214,N_19926,N_19779);
nand UO_1215 (O_1215,N_19950,N_19985);
nand UO_1216 (O_1216,N_19889,N_19986);
or UO_1217 (O_1217,N_19972,N_19764);
nor UO_1218 (O_1218,N_19697,N_19735);
xnor UO_1219 (O_1219,N_19729,N_19737);
xnor UO_1220 (O_1220,N_19754,N_19711);
xor UO_1221 (O_1221,N_19982,N_19831);
and UO_1222 (O_1222,N_19855,N_19642);
xor UO_1223 (O_1223,N_19741,N_19668);
nor UO_1224 (O_1224,N_19802,N_19720);
xor UO_1225 (O_1225,N_19829,N_19661);
nand UO_1226 (O_1226,N_19856,N_19699);
and UO_1227 (O_1227,N_19632,N_19623);
or UO_1228 (O_1228,N_19747,N_19840);
and UO_1229 (O_1229,N_19849,N_19793);
xnor UO_1230 (O_1230,N_19662,N_19750);
or UO_1231 (O_1231,N_19956,N_19632);
xor UO_1232 (O_1232,N_19900,N_19781);
xnor UO_1233 (O_1233,N_19776,N_19904);
or UO_1234 (O_1234,N_19774,N_19982);
and UO_1235 (O_1235,N_19939,N_19979);
or UO_1236 (O_1236,N_19611,N_19742);
xnor UO_1237 (O_1237,N_19731,N_19770);
xnor UO_1238 (O_1238,N_19662,N_19866);
nor UO_1239 (O_1239,N_19686,N_19851);
and UO_1240 (O_1240,N_19997,N_19602);
and UO_1241 (O_1241,N_19733,N_19885);
xor UO_1242 (O_1242,N_19908,N_19971);
xnor UO_1243 (O_1243,N_19921,N_19931);
or UO_1244 (O_1244,N_19978,N_19998);
xor UO_1245 (O_1245,N_19699,N_19976);
and UO_1246 (O_1246,N_19740,N_19698);
nor UO_1247 (O_1247,N_19945,N_19628);
or UO_1248 (O_1248,N_19799,N_19922);
and UO_1249 (O_1249,N_19672,N_19842);
xnor UO_1250 (O_1250,N_19976,N_19608);
and UO_1251 (O_1251,N_19743,N_19639);
and UO_1252 (O_1252,N_19739,N_19676);
xnor UO_1253 (O_1253,N_19785,N_19678);
or UO_1254 (O_1254,N_19643,N_19738);
or UO_1255 (O_1255,N_19901,N_19826);
and UO_1256 (O_1256,N_19744,N_19609);
and UO_1257 (O_1257,N_19852,N_19925);
xor UO_1258 (O_1258,N_19825,N_19720);
xor UO_1259 (O_1259,N_19863,N_19928);
or UO_1260 (O_1260,N_19960,N_19964);
xnor UO_1261 (O_1261,N_19790,N_19955);
and UO_1262 (O_1262,N_19665,N_19896);
or UO_1263 (O_1263,N_19774,N_19916);
nor UO_1264 (O_1264,N_19613,N_19921);
nand UO_1265 (O_1265,N_19732,N_19812);
nand UO_1266 (O_1266,N_19943,N_19997);
nand UO_1267 (O_1267,N_19765,N_19644);
nor UO_1268 (O_1268,N_19614,N_19904);
xor UO_1269 (O_1269,N_19749,N_19819);
or UO_1270 (O_1270,N_19929,N_19819);
nand UO_1271 (O_1271,N_19944,N_19739);
nand UO_1272 (O_1272,N_19997,N_19745);
and UO_1273 (O_1273,N_19708,N_19811);
and UO_1274 (O_1274,N_19811,N_19719);
nor UO_1275 (O_1275,N_19610,N_19625);
xnor UO_1276 (O_1276,N_19680,N_19899);
nor UO_1277 (O_1277,N_19671,N_19998);
nand UO_1278 (O_1278,N_19850,N_19744);
and UO_1279 (O_1279,N_19739,N_19631);
and UO_1280 (O_1280,N_19790,N_19726);
nand UO_1281 (O_1281,N_19802,N_19716);
nor UO_1282 (O_1282,N_19787,N_19811);
xor UO_1283 (O_1283,N_19822,N_19648);
or UO_1284 (O_1284,N_19671,N_19725);
and UO_1285 (O_1285,N_19816,N_19790);
or UO_1286 (O_1286,N_19616,N_19935);
xor UO_1287 (O_1287,N_19665,N_19871);
nor UO_1288 (O_1288,N_19815,N_19868);
nand UO_1289 (O_1289,N_19954,N_19908);
nand UO_1290 (O_1290,N_19676,N_19653);
xnor UO_1291 (O_1291,N_19700,N_19606);
and UO_1292 (O_1292,N_19942,N_19747);
or UO_1293 (O_1293,N_19735,N_19971);
xnor UO_1294 (O_1294,N_19726,N_19975);
or UO_1295 (O_1295,N_19662,N_19770);
nor UO_1296 (O_1296,N_19602,N_19737);
and UO_1297 (O_1297,N_19623,N_19618);
nor UO_1298 (O_1298,N_19716,N_19636);
nand UO_1299 (O_1299,N_19881,N_19919);
nand UO_1300 (O_1300,N_19952,N_19986);
nor UO_1301 (O_1301,N_19642,N_19716);
and UO_1302 (O_1302,N_19766,N_19844);
xor UO_1303 (O_1303,N_19827,N_19602);
nand UO_1304 (O_1304,N_19693,N_19822);
or UO_1305 (O_1305,N_19639,N_19836);
xnor UO_1306 (O_1306,N_19785,N_19610);
nor UO_1307 (O_1307,N_19790,N_19636);
and UO_1308 (O_1308,N_19855,N_19827);
nor UO_1309 (O_1309,N_19977,N_19804);
and UO_1310 (O_1310,N_19704,N_19609);
nor UO_1311 (O_1311,N_19882,N_19948);
nand UO_1312 (O_1312,N_19970,N_19853);
and UO_1313 (O_1313,N_19685,N_19698);
nor UO_1314 (O_1314,N_19779,N_19624);
or UO_1315 (O_1315,N_19612,N_19974);
or UO_1316 (O_1316,N_19737,N_19787);
xor UO_1317 (O_1317,N_19811,N_19983);
nand UO_1318 (O_1318,N_19867,N_19782);
nor UO_1319 (O_1319,N_19835,N_19792);
nand UO_1320 (O_1320,N_19788,N_19905);
xnor UO_1321 (O_1321,N_19785,N_19965);
and UO_1322 (O_1322,N_19823,N_19606);
and UO_1323 (O_1323,N_19957,N_19647);
nor UO_1324 (O_1324,N_19955,N_19742);
and UO_1325 (O_1325,N_19996,N_19779);
and UO_1326 (O_1326,N_19943,N_19705);
xnor UO_1327 (O_1327,N_19714,N_19708);
or UO_1328 (O_1328,N_19639,N_19619);
and UO_1329 (O_1329,N_19894,N_19845);
and UO_1330 (O_1330,N_19625,N_19875);
and UO_1331 (O_1331,N_19675,N_19754);
nor UO_1332 (O_1332,N_19882,N_19676);
and UO_1333 (O_1333,N_19934,N_19789);
xnor UO_1334 (O_1334,N_19764,N_19846);
xor UO_1335 (O_1335,N_19878,N_19905);
nor UO_1336 (O_1336,N_19966,N_19633);
or UO_1337 (O_1337,N_19666,N_19917);
and UO_1338 (O_1338,N_19661,N_19625);
xnor UO_1339 (O_1339,N_19602,N_19977);
nand UO_1340 (O_1340,N_19840,N_19874);
or UO_1341 (O_1341,N_19870,N_19863);
nand UO_1342 (O_1342,N_19794,N_19768);
nor UO_1343 (O_1343,N_19814,N_19891);
and UO_1344 (O_1344,N_19806,N_19818);
and UO_1345 (O_1345,N_19939,N_19624);
xor UO_1346 (O_1346,N_19801,N_19676);
xor UO_1347 (O_1347,N_19654,N_19914);
and UO_1348 (O_1348,N_19739,N_19868);
and UO_1349 (O_1349,N_19903,N_19749);
nand UO_1350 (O_1350,N_19960,N_19950);
or UO_1351 (O_1351,N_19823,N_19791);
and UO_1352 (O_1352,N_19967,N_19944);
nand UO_1353 (O_1353,N_19874,N_19817);
or UO_1354 (O_1354,N_19789,N_19728);
nor UO_1355 (O_1355,N_19924,N_19768);
and UO_1356 (O_1356,N_19690,N_19770);
or UO_1357 (O_1357,N_19923,N_19701);
nor UO_1358 (O_1358,N_19656,N_19793);
nand UO_1359 (O_1359,N_19728,N_19956);
nor UO_1360 (O_1360,N_19760,N_19774);
and UO_1361 (O_1361,N_19914,N_19794);
or UO_1362 (O_1362,N_19745,N_19825);
xor UO_1363 (O_1363,N_19790,N_19998);
and UO_1364 (O_1364,N_19881,N_19897);
and UO_1365 (O_1365,N_19766,N_19809);
nand UO_1366 (O_1366,N_19673,N_19722);
nor UO_1367 (O_1367,N_19628,N_19801);
nand UO_1368 (O_1368,N_19820,N_19791);
and UO_1369 (O_1369,N_19859,N_19801);
or UO_1370 (O_1370,N_19940,N_19842);
xnor UO_1371 (O_1371,N_19831,N_19610);
nand UO_1372 (O_1372,N_19727,N_19923);
nor UO_1373 (O_1373,N_19697,N_19907);
or UO_1374 (O_1374,N_19999,N_19861);
and UO_1375 (O_1375,N_19883,N_19870);
and UO_1376 (O_1376,N_19699,N_19936);
and UO_1377 (O_1377,N_19611,N_19608);
nor UO_1378 (O_1378,N_19901,N_19637);
and UO_1379 (O_1379,N_19665,N_19934);
or UO_1380 (O_1380,N_19854,N_19731);
and UO_1381 (O_1381,N_19777,N_19809);
nand UO_1382 (O_1382,N_19964,N_19727);
or UO_1383 (O_1383,N_19784,N_19809);
nand UO_1384 (O_1384,N_19784,N_19635);
xnor UO_1385 (O_1385,N_19900,N_19687);
nand UO_1386 (O_1386,N_19800,N_19688);
or UO_1387 (O_1387,N_19833,N_19908);
nand UO_1388 (O_1388,N_19788,N_19661);
nand UO_1389 (O_1389,N_19924,N_19896);
or UO_1390 (O_1390,N_19901,N_19864);
xnor UO_1391 (O_1391,N_19662,N_19861);
xor UO_1392 (O_1392,N_19842,N_19818);
nor UO_1393 (O_1393,N_19674,N_19981);
or UO_1394 (O_1394,N_19733,N_19859);
xor UO_1395 (O_1395,N_19865,N_19939);
and UO_1396 (O_1396,N_19987,N_19607);
or UO_1397 (O_1397,N_19954,N_19879);
nor UO_1398 (O_1398,N_19635,N_19607);
or UO_1399 (O_1399,N_19912,N_19929);
nand UO_1400 (O_1400,N_19811,N_19643);
nand UO_1401 (O_1401,N_19814,N_19725);
or UO_1402 (O_1402,N_19656,N_19868);
or UO_1403 (O_1403,N_19837,N_19700);
nand UO_1404 (O_1404,N_19926,N_19993);
xnor UO_1405 (O_1405,N_19634,N_19839);
and UO_1406 (O_1406,N_19622,N_19615);
and UO_1407 (O_1407,N_19848,N_19807);
nand UO_1408 (O_1408,N_19652,N_19748);
and UO_1409 (O_1409,N_19686,N_19896);
nor UO_1410 (O_1410,N_19623,N_19719);
xnor UO_1411 (O_1411,N_19670,N_19736);
nor UO_1412 (O_1412,N_19978,N_19967);
nand UO_1413 (O_1413,N_19969,N_19609);
nor UO_1414 (O_1414,N_19796,N_19672);
and UO_1415 (O_1415,N_19610,N_19633);
xor UO_1416 (O_1416,N_19828,N_19900);
nand UO_1417 (O_1417,N_19950,N_19841);
or UO_1418 (O_1418,N_19778,N_19964);
xor UO_1419 (O_1419,N_19785,N_19914);
nor UO_1420 (O_1420,N_19866,N_19927);
nand UO_1421 (O_1421,N_19915,N_19804);
nor UO_1422 (O_1422,N_19884,N_19738);
or UO_1423 (O_1423,N_19710,N_19976);
xor UO_1424 (O_1424,N_19656,N_19888);
or UO_1425 (O_1425,N_19798,N_19758);
nand UO_1426 (O_1426,N_19716,N_19856);
xor UO_1427 (O_1427,N_19636,N_19958);
xnor UO_1428 (O_1428,N_19614,N_19728);
nand UO_1429 (O_1429,N_19772,N_19817);
and UO_1430 (O_1430,N_19670,N_19710);
nor UO_1431 (O_1431,N_19764,N_19943);
nand UO_1432 (O_1432,N_19793,N_19907);
nand UO_1433 (O_1433,N_19981,N_19879);
xor UO_1434 (O_1434,N_19806,N_19793);
and UO_1435 (O_1435,N_19759,N_19697);
or UO_1436 (O_1436,N_19606,N_19707);
xnor UO_1437 (O_1437,N_19948,N_19601);
and UO_1438 (O_1438,N_19931,N_19831);
and UO_1439 (O_1439,N_19742,N_19643);
or UO_1440 (O_1440,N_19959,N_19956);
or UO_1441 (O_1441,N_19913,N_19765);
nand UO_1442 (O_1442,N_19648,N_19960);
and UO_1443 (O_1443,N_19994,N_19815);
xor UO_1444 (O_1444,N_19827,N_19885);
nor UO_1445 (O_1445,N_19944,N_19973);
nor UO_1446 (O_1446,N_19983,N_19808);
or UO_1447 (O_1447,N_19909,N_19961);
nand UO_1448 (O_1448,N_19765,N_19982);
and UO_1449 (O_1449,N_19771,N_19694);
and UO_1450 (O_1450,N_19632,N_19795);
or UO_1451 (O_1451,N_19800,N_19883);
nand UO_1452 (O_1452,N_19909,N_19778);
nand UO_1453 (O_1453,N_19995,N_19800);
and UO_1454 (O_1454,N_19872,N_19766);
nor UO_1455 (O_1455,N_19653,N_19821);
nor UO_1456 (O_1456,N_19975,N_19955);
and UO_1457 (O_1457,N_19820,N_19609);
nor UO_1458 (O_1458,N_19881,N_19698);
nand UO_1459 (O_1459,N_19757,N_19994);
nor UO_1460 (O_1460,N_19799,N_19683);
or UO_1461 (O_1461,N_19686,N_19907);
nor UO_1462 (O_1462,N_19807,N_19660);
and UO_1463 (O_1463,N_19882,N_19946);
and UO_1464 (O_1464,N_19692,N_19757);
and UO_1465 (O_1465,N_19779,N_19895);
xor UO_1466 (O_1466,N_19986,N_19919);
nor UO_1467 (O_1467,N_19908,N_19719);
nor UO_1468 (O_1468,N_19997,N_19753);
and UO_1469 (O_1469,N_19688,N_19839);
nand UO_1470 (O_1470,N_19691,N_19655);
and UO_1471 (O_1471,N_19691,N_19776);
xor UO_1472 (O_1472,N_19783,N_19837);
xor UO_1473 (O_1473,N_19837,N_19706);
nor UO_1474 (O_1474,N_19770,N_19640);
nor UO_1475 (O_1475,N_19946,N_19821);
nor UO_1476 (O_1476,N_19652,N_19873);
xnor UO_1477 (O_1477,N_19685,N_19890);
or UO_1478 (O_1478,N_19777,N_19723);
nand UO_1479 (O_1479,N_19610,N_19720);
xor UO_1480 (O_1480,N_19607,N_19907);
or UO_1481 (O_1481,N_19752,N_19611);
nor UO_1482 (O_1482,N_19792,N_19889);
xor UO_1483 (O_1483,N_19976,N_19789);
nand UO_1484 (O_1484,N_19785,N_19810);
or UO_1485 (O_1485,N_19848,N_19815);
nor UO_1486 (O_1486,N_19784,N_19724);
or UO_1487 (O_1487,N_19776,N_19917);
nand UO_1488 (O_1488,N_19687,N_19761);
nand UO_1489 (O_1489,N_19991,N_19857);
and UO_1490 (O_1490,N_19883,N_19893);
or UO_1491 (O_1491,N_19997,N_19940);
xor UO_1492 (O_1492,N_19867,N_19754);
nor UO_1493 (O_1493,N_19837,N_19684);
nand UO_1494 (O_1494,N_19615,N_19782);
xnor UO_1495 (O_1495,N_19684,N_19935);
nor UO_1496 (O_1496,N_19618,N_19924);
nor UO_1497 (O_1497,N_19919,N_19912);
and UO_1498 (O_1498,N_19921,N_19731);
or UO_1499 (O_1499,N_19849,N_19942);
nor UO_1500 (O_1500,N_19754,N_19610);
nand UO_1501 (O_1501,N_19913,N_19758);
nand UO_1502 (O_1502,N_19969,N_19871);
xnor UO_1503 (O_1503,N_19765,N_19901);
or UO_1504 (O_1504,N_19957,N_19732);
nor UO_1505 (O_1505,N_19821,N_19797);
or UO_1506 (O_1506,N_19706,N_19695);
nor UO_1507 (O_1507,N_19992,N_19770);
nand UO_1508 (O_1508,N_19878,N_19760);
or UO_1509 (O_1509,N_19787,N_19978);
or UO_1510 (O_1510,N_19855,N_19879);
and UO_1511 (O_1511,N_19605,N_19960);
nand UO_1512 (O_1512,N_19682,N_19924);
and UO_1513 (O_1513,N_19895,N_19601);
and UO_1514 (O_1514,N_19793,N_19931);
xnor UO_1515 (O_1515,N_19815,N_19988);
nor UO_1516 (O_1516,N_19881,N_19666);
nor UO_1517 (O_1517,N_19697,N_19758);
nor UO_1518 (O_1518,N_19963,N_19930);
nor UO_1519 (O_1519,N_19773,N_19951);
or UO_1520 (O_1520,N_19919,N_19832);
nand UO_1521 (O_1521,N_19861,N_19728);
nor UO_1522 (O_1522,N_19899,N_19801);
nand UO_1523 (O_1523,N_19823,N_19981);
xnor UO_1524 (O_1524,N_19845,N_19773);
xor UO_1525 (O_1525,N_19988,N_19703);
nand UO_1526 (O_1526,N_19852,N_19997);
and UO_1527 (O_1527,N_19689,N_19953);
or UO_1528 (O_1528,N_19614,N_19797);
and UO_1529 (O_1529,N_19940,N_19751);
or UO_1530 (O_1530,N_19679,N_19681);
or UO_1531 (O_1531,N_19985,N_19699);
nor UO_1532 (O_1532,N_19938,N_19895);
nor UO_1533 (O_1533,N_19665,N_19865);
nor UO_1534 (O_1534,N_19790,N_19945);
or UO_1535 (O_1535,N_19812,N_19953);
or UO_1536 (O_1536,N_19810,N_19971);
nand UO_1537 (O_1537,N_19679,N_19693);
xor UO_1538 (O_1538,N_19744,N_19674);
nand UO_1539 (O_1539,N_19641,N_19725);
nor UO_1540 (O_1540,N_19843,N_19700);
and UO_1541 (O_1541,N_19668,N_19961);
or UO_1542 (O_1542,N_19666,N_19848);
and UO_1543 (O_1543,N_19751,N_19928);
and UO_1544 (O_1544,N_19806,N_19838);
nor UO_1545 (O_1545,N_19624,N_19790);
nor UO_1546 (O_1546,N_19982,N_19814);
nor UO_1547 (O_1547,N_19985,N_19884);
and UO_1548 (O_1548,N_19969,N_19770);
and UO_1549 (O_1549,N_19741,N_19947);
and UO_1550 (O_1550,N_19842,N_19784);
nor UO_1551 (O_1551,N_19805,N_19879);
nand UO_1552 (O_1552,N_19944,N_19898);
nor UO_1553 (O_1553,N_19738,N_19914);
nand UO_1554 (O_1554,N_19727,N_19649);
or UO_1555 (O_1555,N_19793,N_19775);
xnor UO_1556 (O_1556,N_19725,N_19899);
xor UO_1557 (O_1557,N_19667,N_19732);
xnor UO_1558 (O_1558,N_19642,N_19872);
nand UO_1559 (O_1559,N_19694,N_19952);
nand UO_1560 (O_1560,N_19697,N_19642);
or UO_1561 (O_1561,N_19741,N_19630);
nor UO_1562 (O_1562,N_19644,N_19805);
xnor UO_1563 (O_1563,N_19867,N_19702);
nand UO_1564 (O_1564,N_19779,N_19776);
nand UO_1565 (O_1565,N_19769,N_19764);
and UO_1566 (O_1566,N_19609,N_19939);
nor UO_1567 (O_1567,N_19677,N_19917);
and UO_1568 (O_1568,N_19875,N_19714);
or UO_1569 (O_1569,N_19889,N_19871);
or UO_1570 (O_1570,N_19900,N_19607);
or UO_1571 (O_1571,N_19921,N_19882);
and UO_1572 (O_1572,N_19681,N_19722);
xor UO_1573 (O_1573,N_19805,N_19969);
and UO_1574 (O_1574,N_19892,N_19811);
xor UO_1575 (O_1575,N_19610,N_19761);
and UO_1576 (O_1576,N_19895,N_19671);
xor UO_1577 (O_1577,N_19857,N_19994);
and UO_1578 (O_1578,N_19738,N_19618);
and UO_1579 (O_1579,N_19730,N_19910);
nor UO_1580 (O_1580,N_19759,N_19611);
xor UO_1581 (O_1581,N_19788,N_19606);
and UO_1582 (O_1582,N_19764,N_19670);
nor UO_1583 (O_1583,N_19912,N_19744);
and UO_1584 (O_1584,N_19821,N_19889);
or UO_1585 (O_1585,N_19870,N_19680);
nor UO_1586 (O_1586,N_19644,N_19918);
or UO_1587 (O_1587,N_19874,N_19992);
nand UO_1588 (O_1588,N_19969,N_19671);
nor UO_1589 (O_1589,N_19685,N_19625);
nand UO_1590 (O_1590,N_19781,N_19948);
xor UO_1591 (O_1591,N_19712,N_19952);
or UO_1592 (O_1592,N_19603,N_19947);
or UO_1593 (O_1593,N_19998,N_19653);
or UO_1594 (O_1594,N_19681,N_19892);
nor UO_1595 (O_1595,N_19617,N_19686);
or UO_1596 (O_1596,N_19741,N_19938);
nor UO_1597 (O_1597,N_19812,N_19626);
xor UO_1598 (O_1598,N_19616,N_19638);
xor UO_1599 (O_1599,N_19977,N_19637);
or UO_1600 (O_1600,N_19805,N_19617);
xnor UO_1601 (O_1601,N_19669,N_19626);
or UO_1602 (O_1602,N_19821,N_19853);
xor UO_1603 (O_1603,N_19826,N_19938);
and UO_1604 (O_1604,N_19872,N_19905);
nor UO_1605 (O_1605,N_19679,N_19797);
nor UO_1606 (O_1606,N_19824,N_19790);
nand UO_1607 (O_1607,N_19765,N_19602);
nand UO_1608 (O_1608,N_19795,N_19643);
nand UO_1609 (O_1609,N_19933,N_19945);
xor UO_1610 (O_1610,N_19849,N_19733);
xor UO_1611 (O_1611,N_19638,N_19749);
nor UO_1612 (O_1612,N_19694,N_19673);
nor UO_1613 (O_1613,N_19621,N_19749);
xor UO_1614 (O_1614,N_19969,N_19670);
xnor UO_1615 (O_1615,N_19694,N_19641);
and UO_1616 (O_1616,N_19835,N_19833);
or UO_1617 (O_1617,N_19680,N_19888);
nor UO_1618 (O_1618,N_19699,N_19707);
xor UO_1619 (O_1619,N_19634,N_19757);
nand UO_1620 (O_1620,N_19608,N_19762);
and UO_1621 (O_1621,N_19999,N_19997);
xnor UO_1622 (O_1622,N_19774,N_19831);
or UO_1623 (O_1623,N_19623,N_19760);
xor UO_1624 (O_1624,N_19780,N_19696);
and UO_1625 (O_1625,N_19852,N_19672);
xor UO_1626 (O_1626,N_19753,N_19616);
nor UO_1627 (O_1627,N_19717,N_19732);
or UO_1628 (O_1628,N_19954,N_19681);
and UO_1629 (O_1629,N_19760,N_19847);
nor UO_1630 (O_1630,N_19850,N_19685);
or UO_1631 (O_1631,N_19840,N_19926);
xnor UO_1632 (O_1632,N_19710,N_19907);
and UO_1633 (O_1633,N_19640,N_19670);
and UO_1634 (O_1634,N_19653,N_19757);
and UO_1635 (O_1635,N_19703,N_19717);
nand UO_1636 (O_1636,N_19780,N_19647);
nand UO_1637 (O_1637,N_19666,N_19631);
or UO_1638 (O_1638,N_19850,N_19921);
and UO_1639 (O_1639,N_19811,N_19939);
xor UO_1640 (O_1640,N_19899,N_19727);
nor UO_1641 (O_1641,N_19941,N_19814);
xnor UO_1642 (O_1642,N_19785,N_19982);
and UO_1643 (O_1643,N_19860,N_19898);
xor UO_1644 (O_1644,N_19892,N_19610);
nand UO_1645 (O_1645,N_19826,N_19908);
nor UO_1646 (O_1646,N_19890,N_19818);
and UO_1647 (O_1647,N_19660,N_19686);
or UO_1648 (O_1648,N_19839,N_19726);
or UO_1649 (O_1649,N_19685,N_19796);
and UO_1650 (O_1650,N_19793,N_19948);
nand UO_1651 (O_1651,N_19925,N_19800);
and UO_1652 (O_1652,N_19977,N_19661);
or UO_1653 (O_1653,N_19774,N_19924);
or UO_1654 (O_1654,N_19711,N_19608);
xor UO_1655 (O_1655,N_19899,N_19626);
and UO_1656 (O_1656,N_19931,N_19885);
xnor UO_1657 (O_1657,N_19918,N_19621);
xnor UO_1658 (O_1658,N_19971,N_19946);
nand UO_1659 (O_1659,N_19715,N_19786);
and UO_1660 (O_1660,N_19641,N_19669);
nor UO_1661 (O_1661,N_19842,N_19918);
xor UO_1662 (O_1662,N_19791,N_19978);
and UO_1663 (O_1663,N_19892,N_19766);
or UO_1664 (O_1664,N_19673,N_19616);
xnor UO_1665 (O_1665,N_19792,N_19705);
nor UO_1666 (O_1666,N_19604,N_19906);
nand UO_1667 (O_1667,N_19872,N_19693);
nor UO_1668 (O_1668,N_19844,N_19993);
nand UO_1669 (O_1669,N_19660,N_19881);
nand UO_1670 (O_1670,N_19711,N_19652);
nor UO_1671 (O_1671,N_19772,N_19705);
or UO_1672 (O_1672,N_19904,N_19950);
xor UO_1673 (O_1673,N_19669,N_19613);
or UO_1674 (O_1674,N_19670,N_19654);
or UO_1675 (O_1675,N_19656,N_19601);
xor UO_1676 (O_1676,N_19831,N_19624);
or UO_1677 (O_1677,N_19942,N_19759);
xor UO_1678 (O_1678,N_19647,N_19633);
nand UO_1679 (O_1679,N_19733,N_19945);
nor UO_1680 (O_1680,N_19847,N_19795);
or UO_1681 (O_1681,N_19935,N_19963);
xor UO_1682 (O_1682,N_19707,N_19886);
nor UO_1683 (O_1683,N_19923,N_19649);
and UO_1684 (O_1684,N_19864,N_19984);
nor UO_1685 (O_1685,N_19753,N_19722);
nand UO_1686 (O_1686,N_19758,N_19956);
nor UO_1687 (O_1687,N_19880,N_19820);
or UO_1688 (O_1688,N_19781,N_19636);
nand UO_1689 (O_1689,N_19921,N_19991);
and UO_1690 (O_1690,N_19733,N_19899);
or UO_1691 (O_1691,N_19935,N_19721);
and UO_1692 (O_1692,N_19769,N_19639);
nand UO_1693 (O_1693,N_19819,N_19810);
nand UO_1694 (O_1694,N_19931,N_19988);
nand UO_1695 (O_1695,N_19953,N_19601);
or UO_1696 (O_1696,N_19925,N_19835);
nor UO_1697 (O_1697,N_19756,N_19617);
nor UO_1698 (O_1698,N_19800,N_19805);
xnor UO_1699 (O_1699,N_19697,N_19734);
or UO_1700 (O_1700,N_19667,N_19834);
nor UO_1701 (O_1701,N_19625,N_19963);
nand UO_1702 (O_1702,N_19877,N_19834);
or UO_1703 (O_1703,N_19929,N_19833);
xnor UO_1704 (O_1704,N_19943,N_19687);
nand UO_1705 (O_1705,N_19633,N_19866);
and UO_1706 (O_1706,N_19619,N_19911);
and UO_1707 (O_1707,N_19694,N_19794);
xnor UO_1708 (O_1708,N_19698,N_19943);
nand UO_1709 (O_1709,N_19738,N_19906);
nand UO_1710 (O_1710,N_19875,N_19923);
nand UO_1711 (O_1711,N_19622,N_19662);
or UO_1712 (O_1712,N_19880,N_19668);
nor UO_1713 (O_1713,N_19801,N_19769);
nand UO_1714 (O_1714,N_19746,N_19910);
or UO_1715 (O_1715,N_19626,N_19643);
and UO_1716 (O_1716,N_19813,N_19792);
or UO_1717 (O_1717,N_19744,N_19766);
and UO_1718 (O_1718,N_19990,N_19604);
and UO_1719 (O_1719,N_19998,N_19851);
xnor UO_1720 (O_1720,N_19836,N_19858);
or UO_1721 (O_1721,N_19968,N_19674);
and UO_1722 (O_1722,N_19795,N_19765);
nor UO_1723 (O_1723,N_19752,N_19732);
and UO_1724 (O_1724,N_19920,N_19697);
nor UO_1725 (O_1725,N_19777,N_19864);
xor UO_1726 (O_1726,N_19820,N_19945);
or UO_1727 (O_1727,N_19640,N_19892);
nand UO_1728 (O_1728,N_19751,N_19799);
xnor UO_1729 (O_1729,N_19845,N_19766);
nand UO_1730 (O_1730,N_19851,N_19685);
and UO_1731 (O_1731,N_19870,N_19865);
nand UO_1732 (O_1732,N_19697,N_19768);
nand UO_1733 (O_1733,N_19615,N_19786);
nor UO_1734 (O_1734,N_19925,N_19766);
nand UO_1735 (O_1735,N_19730,N_19980);
nand UO_1736 (O_1736,N_19925,N_19940);
nand UO_1737 (O_1737,N_19971,N_19713);
and UO_1738 (O_1738,N_19786,N_19918);
nand UO_1739 (O_1739,N_19767,N_19668);
xor UO_1740 (O_1740,N_19630,N_19704);
nor UO_1741 (O_1741,N_19600,N_19904);
and UO_1742 (O_1742,N_19772,N_19985);
and UO_1743 (O_1743,N_19846,N_19784);
or UO_1744 (O_1744,N_19737,N_19840);
or UO_1745 (O_1745,N_19732,N_19639);
xnor UO_1746 (O_1746,N_19964,N_19906);
nand UO_1747 (O_1747,N_19940,N_19760);
nor UO_1748 (O_1748,N_19922,N_19747);
xor UO_1749 (O_1749,N_19877,N_19996);
nand UO_1750 (O_1750,N_19814,N_19616);
or UO_1751 (O_1751,N_19637,N_19879);
nand UO_1752 (O_1752,N_19978,N_19742);
or UO_1753 (O_1753,N_19841,N_19682);
and UO_1754 (O_1754,N_19830,N_19646);
nor UO_1755 (O_1755,N_19732,N_19885);
and UO_1756 (O_1756,N_19984,N_19824);
nand UO_1757 (O_1757,N_19887,N_19814);
xor UO_1758 (O_1758,N_19687,N_19998);
nand UO_1759 (O_1759,N_19928,N_19895);
and UO_1760 (O_1760,N_19633,N_19741);
nand UO_1761 (O_1761,N_19600,N_19687);
and UO_1762 (O_1762,N_19611,N_19822);
and UO_1763 (O_1763,N_19910,N_19697);
and UO_1764 (O_1764,N_19824,N_19653);
xor UO_1765 (O_1765,N_19623,N_19669);
nand UO_1766 (O_1766,N_19603,N_19831);
nor UO_1767 (O_1767,N_19939,N_19787);
or UO_1768 (O_1768,N_19624,N_19869);
xor UO_1769 (O_1769,N_19816,N_19882);
xnor UO_1770 (O_1770,N_19602,N_19987);
and UO_1771 (O_1771,N_19954,N_19772);
xor UO_1772 (O_1772,N_19796,N_19929);
and UO_1773 (O_1773,N_19690,N_19689);
xnor UO_1774 (O_1774,N_19926,N_19882);
xnor UO_1775 (O_1775,N_19767,N_19713);
xnor UO_1776 (O_1776,N_19957,N_19801);
nand UO_1777 (O_1777,N_19849,N_19804);
nand UO_1778 (O_1778,N_19867,N_19931);
and UO_1779 (O_1779,N_19744,N_19790);
nand UO_1780 (O_1780,N_19639,N_19734);
and UO_1781 (O_1781,N_19848,N_19977);
or UO_1782 (O_1782,N_19642,N_19820);
or UO_1783 (O_1783,N_19805,N_19771);
nand UO_1784 (O_1784,N_19883,N_19617);
nor UO_1785 (O_1785,N_19812,N_19917);
nand UO_1786 (O_1786,N_19862,N_19989);
nand UO_1787 (O_1787,N_19818,N_19762);
and UO_1788 (O_1788,N_19834,N_19982);
and UO_1789 (O_1789,N_19781,N_19863);
and UO_1790 (O_1790,N_19952,N_19963);
nor UO_1791 (O_1791,N_19895,N_19621);
and UO_1792 (O_1792,N_19793,N_19769);
and UO_1793 (O_1793,N_19818,N_19923);
nand UO_1794 (O_1794,N_19868,N_19700);
and UO_1795 (O_1795,N_19625,N_19659);
or UO_1796 (O_1796,N_19723,N_19847);
nand UO_1797 (O_1797,N_19775,N_19818);
nand UO_1798 (O_1798,N_19934,N_19883);
and UO_1799 (O_1799,N_19872,N_19954);
or UO_1800 (O_1800,N_19879,N_19801);
nor UO_1801 (O_1801,N_19792,N_19902);
or UO_1802 (O_1802,N_19622,N_19786);
nand UO_1803 (O_1803,N_19990,N_19747);
xnor UO_1804 (O_1804,N_19818,N_19619);
nor UO_1805 (O_1805,N_19836,N_19602);
nand UO_1806 (O_1806,N_19735,N_19604);
xor UO_1807 (O_1807,N_19605,N_19614);
or UO_1808 (O_1808,N_19918,N_19616);
nor UO_1809 (O_1809,N_19948,N_19924);
or UO_1810 (O_1810,N_19917,N_19799);
nor UO_1811 (O_1811,N_19865,N_19735);
xor UO_1812 (O_1812,N_19848,N_19739);
nand UO_1813 (O_1813,N_19681,N_19907);
and UO_1814 (O_1814,N_19744,N_19774);
xor UO_1815 (O_1815,N_19786,N_19859);
nor UO_1816 (O_1816,N_19743,N_19873);
xor UO_1817 (O_1817,N_19807,N_19664);
or UO_1818 (O_1818,N_19828,N_19925);
nand UO_1819 (O_1819,N_19937,N_19717);
xnor UO_1820 (O_1820,N_19946,N_19879);
xnor UO_1821 (O_1821,N_19812,N_19863);
xor UO_1822 (O_1822,N_19748,N_19755);
nand UO_1823 (O_1823,N_19808,N_19778);
and UO_1824 (O_1824,N_19733,N_19980);
and UO_1825 (O_1825,N_19658,N_19835);
nor UO_1826 (O_1826,N_19949,N_19788);
or UO_1827 (O_1827,N_19879,N_19859);
nor UO_1828 (O_1828,N_19908,N_19767);
and UO_1829 (O_1829,N_19966,N_19989);
and UO_1830 (O_1830,N_19621,N_19920);
and UO_1831 (O_1831,N_19892,N_19904);
nor UO_1832 (O_1832,N_19904,N_19734);
and UO_1833 (O_1833,N_19995,N_19634);
xnor UO_1834 (O_1834,N_19645,N_19763);
and UO_1835 (O_1835,N_19872,N_19991);
and UO_1836 (O_1836,N_19937,N_19897);
or UO_1837 (O_1837,N_19674,N_19859);
xor UO_1838 (O_1838,N_19954,N_19983);
xnor UO_1839 (O_1839,N_19646,N_19873);
and UO_1840 (O_1840,N_19736,N_19925);
xor UO_1841 (O_1841,N_19717,N_19958);
xor UO_1842 (O_1842,N_19646,N_19984);
or UO_1843 (O_1843,N_19722,N_19706);
xnor UO_1844 (O_1844,N_19665,N_19900);
nor UO_1845 (O_1845,N_19611,N_19699);
and UO_1846 (O_1846,N_19988,N_19848);
or UO_1847 (O_1847,N_19855,N_19950);
and UO_1848 (O_1848,N_19731,N_19826);
xor UO_1849 (O_1849,N_19722,N_19853);
and UO_1850 (O_1850,N_19696,N_19645);
nor UO_1851 (O_1851,N_19974,N_19761);
and UO_1852 (O_1852,N_19989,N_19760);
or UO_1853 (O_1853,N_19905,N_19898);
and UO_1854 (O_1854,N_19743,N_19847);
nand UO_1855 (O_1855,N_19831,N_19606);
nand UO_1856 (O_1856,N_19774,N_19680);
and UO_1857 (O_1857,N_19928,N_19894);
or UO_1858 (O_1858,N_19759,N_19844);
nand UO_1859 (O_1859,N_19924,N_19790);
and UO_1860 (O_1860,N_19626,N_19824);
nand UO_1861 (O_1861,N_19820,N_19704);
or UO_1862 (O_1862,N_19938,N_19784);
xnor UO_1863 (O_1863,N_19723,N_19965);
xnor UO_1864 (O_1864,N_19967,N_19930);
nand UO_1865 (O_1865,N_19984,N_19670);
and UO_1866 (O_1866,N_19642,N_19991);
nand UO_1867 (O_1867,N_19695,N_19804);
and UO_1868 (O_1868,N_19912,N_19678);
xor UO_1869 (O_1869,N_19665,N_19651);
nand UO_1870 (O_1870,N_19973,N_19620);
nand UO_1871 (O_1871,N_19903,N_19610);
or UO_1872 (O_1872,N_19822,N_19906);
and UO_1873 (O_1873,N_19844,N_19656);
nor UO_1874 (O_1874,N_19846,N_19794);
xor UO_1875 (O_1875,N_19914,N_19675);
nand UO_1876 (O_1876,N_19657,N_19649);
and UO_1877 (O_1877,N_19630,N_19988);
nand UO_1878 (O_1878,N_19762,N_19746);
and UO_1879 (O_1879,N_19777,N_19910);
nand UO_1880 (O_1880,N_19761,N_19888);
xor UO_1881 (O_1881,N_19632,N_19769);
or UO_1882 (O_1882,N_19621,N_19862);
or UO_1883 (O_1883,N_19976,N_19849);
nand UO_1884 (O_1884,N_19673,N_19626);
nor UO_1885 (O_1885,N_19850,N_19819);
nor UO_1886 (O_1886,N_19709,N_19960);
nor UO_1887 (O_1887,N_19688,N_19639);
or UO_1888 (O_1888,N_19769,N_19808);
or UO_1889 (O_1889,N_19761,N_19703);
and UO_1890 (O_1890,N_19787,N_19627);
xor UO_1891 (O_1891,N_19967,N_19787);
xnor UO_1892 (O_1892,N_19790,N_19634);
and UO_1893 (O_1893,N_19739,N_19916);
nor UO_1894 (O_1894,N_19909,N_19868);
xor UO_1895 (O_1895,N_19604,N_19915);
or UO_1896 (O_1896,N_19640,N_19750);
or UO_1897 (O_1897,N_19863,N_19929);
nor UO_1898 (O_1898,N_19761,N_19727);
or UO_1899 (O_1899,N_19634,N_19786);
xnor UO_1900 (O_1900,N_19802,N_19725);
nand UO_1901 (O_1901,N_19689,N_19656);
and UO_1902 (O_1902,N_19712,N_19613);
xor UO_1903 (O_1903,N_19615,N_19822);
nor UO_1904 (O_1904,N_19977,N_19879);
and UO_1905 (O_1905,N_19897,N_19935);
and UO_1906 (O_1906,N_19922,N_19954);
xnor UO_1907 (O_1907,N_19892,N_19613);
xnor UO_1908 (O_1908,N_19796,N_19769);
nor UO_1909 (O_1909,N_19757,N_19985);
nor UO_1910 (O_1910,N_19786,N_19982);
xor UO_1911 (O_1911,N_19771,N_19897);
and UO_1912 (O_1912,N_19962,N_19684);
and UO_1913 (O_1913,N_19611,N_19635);
and UO_1914 (O_1914,N_19760,N_19959);
or UO_1915 (O_1915,N_19765,N_19831);
nand UO_1916 (O_1916,N_19734,N_19603);
nor UO_1917 (O_1917,N_19824,N_19887);
or UO_1918 (O_1918,N_19870,N_19843);
or UO_1919 (O_1919,N_19779,N_19614);
and UO_1920 (O_1920,N_19850,N_19664);
nor UO_1921 (O_1921,N_19650,N_19957);
nor UO_1922 (O_1922,N_19744,N_19695);
nand UO_1923 (O_1923,N_19728,N_19834);
or UO_1924 (O_1924,N_19708,N_19825);
nor UO_1925 (O_1925,N_19752,N_19817);
and UO_1926 (O_1926,N_19748,N_19877);
and UO_1927 (O_1927,N_19910,N_19605);
and UO_1928 (O_1928,N_19971,N_19992);
and UO_1929 (O_1929,N_19834,N_19997);
and UO_1930 (O_1930,N_19831,N_19976);
nor UO_1931 (O_1931,N_19817,N_19927);
nand UO_1932 (O_1932,N_19957,N_19934);
nand UO_1933 (O_1933,N_19629,N_19781);
or UO_1934 (O_1934,N_19696,N_19882);
nand UO_1935 (O_1935,N_19616,N_19757);
nor UO_1936 (O_1936,N_19615,N_19703);
nand UO_1937 (O_1937,N_19606,N_19805);
nand UO_1938 (O_1938,N_19892,N_19710);
nand UO_1939 (O_1939,N_19727,N_19882);
and UO_1940 (O_1940,N_19817,N_19919);
and UO_1941 (O_1941,N_19963,N_19699);
nand UO_1942 (O_1942,N_19878,N_19630);
or UO_1943 (O_1943,N_19892,N_19997);
or UO_1944 (O_1944,N_19709,N_19776);
nand UO_1945 (O_1945,N_19917,N_19854);
or UO_1946 (O_1946,N_19865,N_19857);
or UO_1947 (O_1947,N_19941,N_19620);
nor UO_1948 (O_1948,N_19731,N_19696);
xnor UO_1949 (O_1949,N_19953,N_19757);
and UO_1950 (O_1950,N_19957,N_19744);
xnor UO_1951 (O_1951,N_19989,N_19829);
nand UO_1952 (O_1952,N_19668,N_19927);
nand UO_1953 (O_1953,N_19986,N_19646);
nor UO_1954 (O_1954,N_19902,N_19705);
or UO_1955 (O_1955,N_19850,N_19607);
or UO_1956 (O_1956,N_19785,N_19978);
nor UO_1957 (O_1957,N_19601,N_19684);
nor UO_1958 (O_1958,N_19694,N_19942);
nand UO_1959 (O_1959,N_19955,N_19650);
and UO_1960 (O_1960,N_19887,N_19786);
or UO_1961 (O_1961,N_19612,N_19888);
nor UO_1962 (O_1962,N_19988,N_19891);
xnor UO_1963 (O_1963,N_19770,N_19833);
nand UO_1964 (O_1964,N_19631,N_19664);
nor UO_1965 (O_1965,N_19702,N_19846);
and UO_1966 (O_1966,N_19961,N_19613);
and UO_1967 (O_1967,N_19871,N_19802);
nand UO_1968 (O_1968,N_19704,N_19750);
xnor UO_1969 (O_1969,N_19763,N_19863);
nand UO_1970 (O_1970,N_19880,N_19804);
or UO_1971 (O_1971,N_19706,N_19866);
and UO_1972 (O_1972,N_19677,N_19646);
nand UO_1973 (O_1973,N_19986,N_19869);
or UO_1974 (O_1974,N_19760,N_19809);
nand UO_1975 (O_1975,N_19900,N_19747);
or UO_1976 (O_1976,N_19853,N_19919);
nor UO_1977 (O_1977,N_19998,N_19990);
and UO_1978 (O_1978,N_19868,N_19610);
nand UO_1979 (O_1979,N_19774,N_19794);
and UO_1980 (O_1980,N_19866,N_19705);
and UO_1981 (O_1981,N_19631,N_19882);
nand UO_1982 (O_1982,N_19757,N_19983);
and UO_1983 (O_1983,N_19793,N_19646);
or UO_1984 (O_1984,N_19765,N_19890);
and UO_1985 (O_1985,N_19912,N_19826);
or UO_1986 (O_1986,N_19610,N_19907);
nand UO_1987 (O_1987,N_19629,N_19624);
xnor UO_1988 (O_1988,N_19868,N_19870);
xnor UO_1989 (O_1989,N_19982,N_19950);
nor UO_1990 (O_1990,N_19763,N_19668);
xnor UO_1991 (O_1991,N_19686,N_19793);
nor UO_1992 (O_1992,N_19625,N_19773);
and UO_1993 (O_1993,N_19604,N_19984);
xnor UO_1994 (O_1994,N_19786,N_19635);
nand UO_1995 (O_1995,N_19735,N_19658);
or UO_1996 (O_1996,N_19801,N_19692);
nand UO_1997 (O_1997,N_19671,N_19786);
xnor UO_1998 (O_1998,N_19862,N_19669);
nand UO_1999 (O_1999,N_19831,N_19861);
xnor UO_2000 (O_2000,N_19719,N_19708);
nor UO_2001 (O_2001,N_19824,N_19934);
xor UO_2002 (O_2002,N_19749,N_19947);
or UO_2003 (O_2003,N_19890,N_19655);
or UO_2004 (O_2004,N_19625,N_19746);
xnor UO_2005 (O_2005,N_19929,N_19986);
xor UO_2006 (O_2006,N_19730,N_19694);
xor UO_2007 (O_2007,N_19974,N_19673);
nand UO_2008 (O_2008,N_19605,N_19903);
nand UO_2009 (O_2009,N_19927,N_19934);
nor UO_2010 (O_2010,N_19761,N_19790);
xnor UO_2011 (O_2011,N_19619,N_19940);
nand UO_2012 (O_2012,N_19941,N_19868);
xnor UO_2013 (O_2013,N_19646,N_19613);
or UO_2014 (O_2014,N_19821,N_19798);
xnor UO_2015 (O_2015,N_19966,N_19946);
xnor UO_2016 (O_2016,N_19905,N_19600);
xnor UO_2017 (O_2017,N_19790,N_19690);
or UO_2018 (O_2018,N_19717,N_19970);
or UO_2019 (O_2019,N_19967,N_19863);
nor UO_2020 (O_2020,N_19836,N_19864);
or UO_2021 (O_2021,N_19940,N_19688);
or UO_2022 (O_2022,N_19696,N_19883);
xor UO_2023 (O_2023,N_19888,N_19749);
and UO_2024 (O_2024,N_19985,N_19741);
and UO_2025 (O_2025,N_19710,N_19804);
nor UO_2026 (O_2026,N_19845,N_19708);
nor UO_2027 (O_2027,N_19925,N_19778);
xor UO_2028 (O_2028,N_19996,N_19769);
and UO_2029 (O_2029,N_19998,N_19727);
xor UO_2030 (O_2030,N_19602,N_19614);
xor UO_2031 (O_2031,N_19962,N_19731);
xnor UO_2032 (O_2032,N_19974,N_19823);
or UO_2033 (O_2033,N_19840,N_19843);
nand UO_2034 (O_2034,N_19753,N_19809);
xor UO_2035 (O_2035,N_19757,N_19699);
xnor UO_2036 (O_2036,N_19773,N_19933);
nor UO_2037 (O_2037,N_19846,N_19688);
xnor UO_2038 (O_2038,N_19831,N_19758);
nor UO_2039 (O_2039,N_19904,N_19985);
xnor UO_2040 (O_2040,N_19870,N_19889);
xnor UO_2041 (O_2041,N_19927,N_19830);
or UO_2042 (O_2042,N_19979,N_19771);
or UO_2043 (O_2043,N_19734,N_19893);
or UO_2044 (O_2044,N_19858,N_19841);
or UO_2045 (O_2045,N_19721,N_19827);
nor UO_2046 (O_2046,N_19867,N_19792);
and UO_2047 (O_2047,N_19800,N_19815);
nor UO_2048 (O_2048,N_19787,N_19751);
nor UO_2049 (O_2049,N_19638,N_19751);
nor UO_2050 (O_2050,N_19777,N_19894);
xnor UO_2051 (O_2051,N_19818,N_19913);
or UO_2052 (O_2052,N_19914,N_19917);
nor UO_2053 (O_2053,N_19872,N_19666);
and UO_2054 (O_2054,N_19703,N_19612);
and UO_2055 (O_2055,N_19882,N_19888);
and UO_2056 (O_2056,N_19797,N_19666);
nand UO_2057 (O_2057,N_19841,N_19969);
xnor UO_2058 (O_2058,N_19838,N_19994);
nor UO_2059 (O_2059,N_19761,N_19600);
xor UO_2060 (O_2060,N_19904,N_19983);
nand UO_2061 (O_2061,N_19958,N_19610);
or UO_2062 (O_2062,N_19758,N_19753);
or UO_2063 (O_2063,N_19926,N_19670);
or UO_2064 (O_2064,N_19917,N_19768);
and UO_2065 (O_2065,N_19936,N_19786);
and UO_2066 (O_2066,N_19600,N_19625);
and UO_2067 (O_2067,N_19757,N_19900);
or UO_2068 (O_2068,N_19888,N_19625);
xnor UO_2069 (O_2069,N_19673,N_19842);
nand UO_2070 (O_2070,N_19984,N_19913);
and UO_2071 (O_2071,N_19978,N_19866);
and UO_2072 (O_2072,N_19740,N_19649);
nand UO_2073 (O_2073,N_19675,N_19652);
and UO_2074 (O_2074,N_19836,N_19863);
or UO_2075 (O_2075,N_19855,N_19668);
or UO_2076 (O_2076,N_19697,N_19909);
or UO_2077 (O_2077,N_19922,N_19963);
or UO_2078 (O_2078,N_19827,N_19833);
nor UO_2079 (O_2079,N_19870,N_19986);
nand UO_2080 (O_2080,N_19653,N_19747);
xnor UO_2081 (O_2081,N_19985,N_19976);
nor UO_2082 (O_2082,N_19748,N_19955);
xor UO_2083 (O_2083,N_19898,N_19655);
and UO_2084 (O_2084,N_19636,N_19997);
nand UO_2085 (O_2085,N_19854,N_19835);
nand UO_2086 (O_2086,N_19889,N_19925);
or UO_2087 (O_2087,N_19641,N_19983);
or UO_2088 (O_2088,N_19690,N_19622);
nand UO_2089 (O_2089,N_19918,N_19661);
xnor UO_2090 (O_2090,N_19739,N_19887);
or UO_2091 (O_2091,N_19869,N_19851);
nand UO_2092 (O_2092,N_19931,N_19898);
nor UO_2093 (O_2093,N_19823,N_19886);
xnor UO_2094 (O_2094,N_19927,N_19800);
nand UO_2095 (O_2095,N_19692,N_19912);
and UO_2096 (O_2096,N_19829,N_19804);
or UO_2097 (O_2097,N_19927,N_19877);
xnor UO_2098 (O_2098,N_19800,N_19900);
and UO_2099 (O_2099,N_19978,N_19621);
nand UO_2100 (O_2100,N_19892,N_19864);
xnor UO_2101 (O_2101,N_19801,N_19686);
nor UO_2102 (O_2102,N_19646,N_19829);
and UO_2103 (O_2103,N_19713,N_19989);
xor UO_2104 (O_2104,N_19741,N_19944);
nand UO_2105 (O_2105,N_19754,N_19965);
or UO_2106 (O_2106,N_19791,N_19897);
xor UO_2107 (O_2107,N_19773,N_19828);
nand UO_2108 (O_2108,N_19919,N_19829);
nand UO_2109 (O_2109,N_19666,N_19836);
or UO_2110 (O_2110,N_19891,N_19647);
or UO_2111 (O_2111,N_19845,N_19836);
xor UO_2112 (O_2112,N_19867,N_19935);
nand UO_2113 (O_2113,N_19760,N_19646);
nand UO_2114 (O_2114,N_19847,N_19751);
nor UO_2115 (O_2115,N_19835,N_19682);
xor UO_2116 (O_2116,N_19974,N_19966);
xnor UO_2117 (O_2117,N_19851,N_19902);
and UO_2118 (O_2118,N_19747,N_19968);
nor UO_2119 (O_2119,N_19658,N_19615);
xnor UO_2120 (O_2120,N_19840,N_19684);
nor UO_2121 (O_2121,N_19832,N_19846);
and UO_2122 (O_2122,N_19651,N_19702);
nand UO_2123 (O_2123,N_19738,N_19853);
or UO_2124 (O_2124,N_19722,N_19762);
xor UO_2125 (O_2125,N_19777,N_19815);
xor UO_2126 (O_2126,N_19609,N_19648);
xor UO_2127 (O_2127,N_19757,N_19840);
and UO_2128 (O_2128,N_19962,N_19669);
nor UO_2129 (O_2129,N_19648,N_19849);
or UO_2130 (O_2130,N_19896,N_19704);
nand UO_2131 (O_2131,N_19985,N_19944);
nand UO_2132 (O_2132,N_19712,N_19620);
or UO_2133 (O_2133,N_19645,N_19758);
and UO_2134 (O_2134,N_19831,N_19986);
and UO_2135 (O_2135,N_19969,N_19700);
and UO_2136 (O_2136,N_19693,N_19815);
nor UO_2137 (O_2137,N_19816,N_19976);
or UO_2138 (O_2138,N_19961,N_19886);
or UO_2139 (O_2139,N_19670,N_19902);
nor UO_2140 (O_2140,N_19985,N_19833);
xnor UO_2141 (O_2141,N_19866,N_19660);
or UO_2142 (O_2142,N_19621,N_19658);
nand UO_2143 (O_2143,N_19999,N_19741);
nor UO_2144 (O_2144,N_19828,N_19747);
xor UO_2145 (O_2145,N_19840,N_19865);
nor UO_2146 (O_2146,N_19754,N_19653);
or UO_2147 (O_2147,N_19890,N_19783);
nand UO_2148 (O_2148,N_19873,N_19799);
or UO_2149 (O_2149,N_19933,N_19701);
nand UO_2150 (O_2150,N_19959,N_19895);
or UO_2151 (O_2151,N_19900,N_19863);
xor UO_2152 (O_2152,N_19895,N_19756);
nor UO_2153 (O_2153,N_19969,N_19629);
and UO_2154 (O_2154,N_19984,N_19807);
nor UO_2155 (O_2155,N_19687,N_19608);
and UO_2156 (O_2156,N_19723,N_19939);
and UO_2157 (O_2157,N_19604,N_19958);
or UO_2158 (O_2158,N_19659,N_19919);
nand UO_2159 (O_2159,N_19829,N_19639);
and UO_2160 (O_2160,N_19643,N_19704);
and UO_2161 (O_2161,N_19820,N_19778);
or UO_2162 (O_2162,N_19764,N_19951);
or UO_2163 (O_2163,N_19815,N_19801);
nor UO_2164 (O_2164,N_19870,N_19965);
nand UO_2165 (O_2165,N_19631,N_19612);
nand UO_2166 (O_2166,N_19708,N_19877);
nand UO_2167 (O_2167,N_19734,N_19692);
xnor UO_2168 (O_2168,N_19823,N_19704);
xnor UO_2169 (O_2169,N_19954,N_19782);
nand UO_2170 (O_2170,N_19810,N_19912);
nor UO_2171 (O_2171,N_19694,N_19832);
or UO_2172 (O_2172,N_19775,N_19643);
nand UO_2173 (O_2173,N_19902,N_19932);
xnor UO_2174 (O_2174,N_19611,N_19697);
or UO_2175 (O_2175,N_19966,N_19641);
and UO_2176 (O_2176,N_19774,N_19914);
xor UO_2177 (O_2177,N_19710,N_19604);
nand UO_2178 (O_2178,N_19811,N_19679);
xnor UO_2179 (O_2179,N_19747,N_19658);
nor UO_2180 (O_2180,N_19633,N_19764);
xor UO_2181 (O_2181,N_19820,N_19874);
or UO_2182 (O_2182,N_19616,N_19678);
nor UO_2183 (O_2183,N_19759,N_19986);
nand UO_2184 (O_2184,N_19877,N_19838);
and UO_2185 (O_2185,N_19991,N_19697);
and UO_2186 (O_2186,N_19997,N_19984);
nor UO_2187 (O_2187,N_19618,N_19926);
nand UO_2188 (O_2188,N_19612,N_19729);
nor UO_2189 (O_2189,N_19744,N_19807);
nand UO_2190 (O_2190,N_19933,N_19768);
nor UO_2191 (O_2191,N_19800,N_19889);
nor UO_2192 (O_2192,N_19842,N_19942);
and UO_2193 (O_2193,N_19708,N_19985);
nor UO_2194 (O_2194,N_19694,N_19721);
xnor UO_2195 (O_2195,N_19702,N_19602);
nand UO_2196 (O_2196,N_19802,N_19943);
nand UO_2197 (O_2197,N_19910,N_19630);
or UO_2198 (O_2198,N_19864,N_19679);
xnor UO_2199 (O_2199,N_19959,N_19719);
or UO_2200 (O_2200,N_19841,N_19630);
or UO_2201 (O_2201,N_19771,N_19901);
or UO_2202 (O_2202,N_19887,N_19653);
or UO_2203 (O_2203,N_19817,N_19839);
or UO_2204 (O_2204,N_19979,N_19734);
nand UO_2205 (O_2205,N_19709,N_19801);
or UO_2206 (O_2206,N_19715,N_19667);
xor UO_2207 (O_2207,N_19816,N_19992);
or UO_2208 (O_2208,N_19896,N_19933);
or UO_2209 (O_2209,N_19713,N_19972);
nor UO_2210 (O_2210,N_19667,N_19824);
and UO_2211 (O_2211,N_19921,N_19663);
nand UO_2212 (O_2212,N_19842,N_19606);
or UO_2213 (O_2213,N_19897,N_19605);
xnor UO_2214 (O_2214,N_19870,N_19737);
and UO_2215 (O_2215,N_19825,N_19794);
or UO_2216 (O_2216,N_19831,N_19670);
xor UO_2217 (O_2217,N_19831,N_19622);
or UO_2218 (O_2218,N_19615,N_19798);
nand UO_2219 (O_2219,N_19861,N_19729);
nand UO_2220 (O_2220,N_19964,N_19677);
and UO_2221 (O_2221,N_19968,N_19787);
and UO_2222 (O_2222,N_19879,N_19638);
nand UO_2223 (O_2223,N_19772,N_19633);
and UO_2224 (O_2224,N_19914,N_19846);
nand UO_2225 (O_2225,N_19940,N_19965);
or UO_2226 (O_2226,N_19649,N_19736);
nand UO_2227 (O_2227,N_19771,N_19704);
nor UO_2228 (O_2228,N_19670,N_19632);
xor UO_2229 (O_2229,N_19970,N_19762);
nor UO_2230 (O_2230,N_19912,N_19605);
xnor UO_2231 (O_2231,N_19870,N_19970);
nor UO_2232 (O_2232,N_19666,N_19843);
nor UO_2233 (O_2233,N_19882,N_19901);
nor UO_2234 (O_2234,N_19647,N_19932);
and UO_2235 (O_2235,N_19783,N_19655);
nor UO_2236 (O_2236,N_19865,N_19686);
xor UO_2237 (O_2237,N_19927,N_19883);
xor UO_2238 (O_2238,N_19999,N_19615);
nand UO_2239 (O_2239,N_19833,N_19703);
xor UO_2240 (O_2240,N_19977,N_19761);
and UO_2241 (O_2241,N_19616,N_19931);
and UO_2242 (O_2242,N_19935,N_19834);
and UO_2243 (O_2243,N_19782,N_19906);
and UO_2244 (O_2244,N_19986,N_19964);
nor UO_2245 (O_2245,N_19874,N_19628);
nor UO_2246 (O_2246,N_19985,N_19655);
nor UO_2247 (O_2247,N_19666,N_19740);
nor UO_2248 (O_2248,N_19749,N_19905);
nand UO_2249 (O_2249,N_19651,N_19610);
or UO_2250 (O_2250,N_19976,N_19882);
nor UO_2251 (O_2251,N_19982,N_19897);
nand UO_2252 (O_2252,N_19954,N_19741);
nand UO_2253 (O_2253,N_19672,N_19790);
xor UO_2254 (O_2254,N_19994,N_19719);
or UO_2255 (O_2255,N_19712,N_19854);
nor UO_2256 (O_2256,N_19977,N_19934);
and UO_2257 (O_2257,N_19887,N_19807);
or UO_2258 (O_2258,N_19956,N_19920);
nor UO_2259 (O_2259,N_19818,N_19785);
nor UO_2260 (O_2260,N_19738,N_19916);
or UO_2261 (O_2261,N_19778,N_19932);
nor UO_2262 (O_2262,N_19762,N_19735);
and UO_2263 (O_2263,N_19611,N_19605);
xor UO_2264 (O_2264,N_19711,N_19813);
xor UO_2265 (O_2265,N_19797,N_19759);
xor UO_2266 (O_2266,N_19932,N_19723);
and UO_2267 (O_2267,N_19621,N_19662);
xor UO_2268 (O_2268,N_19674,N_19896);
and UO_2269 (O_2269,N_19958,N_19791);
nand UO_2270 (O_2270,N_19985,N_19829);
xor UO_2271 (O_2271,N_19886,N_19632);
nand UO_2272 (O_2272,N_19860,N_19835);
nand UO_2273 (O_2273,N_19802,N_19812);
or UO_2274 (O_2274,N_19652,N_19757);
nand UO_2275 (O_2275,N_19914,N_19798);
or UO_2276 (O_2276,N_19665,N_19846);
nand UO_2277 (O_2277,N_19736,N_19746);
and UO_2278 (O_2278,N_19655,N_19735);
xnor UO_2279 (O_2279,N_19825,N_19813);
xor UO_2280 (O_2280,N_19929,N_19937);
and UO_2281 (O_2281,N_19870,N_19797);
xnor UO_2282 (O_2282,N_19607,N_19747);
nand UO_2283 (O_2283,N_19901,N_19955);
nand UO_2284 (O_2284,N_19735,N_19934);
xor UO_2285 (O_2285,N_19682,N_19878);
and UO_2286 (O_2286,N_19810,N_19662);
xor UO_2287 (O_2287,N_19721,N_19988);
nand UO_2288 (O_2288,N_19937,N_19676);
or UO_2289 (O_2289,N_19652,N_19966);
or UO_2290 (O_2290,N_19668,N_19743);
or UO_2291 (O_2291,N_19996,N_19790);
or UO_2292 (O_2292,N_19922,N_19728);
nand UO_2293 (O_2293,N_19739,N_19664);
xnor UO_2294 (O_2294,N_19985,N_19828);
nand UO_2295 (O_2295,N_19837,N_19616);
nor UO_2296 (O_2296,N_19821,N_19627);
xnor UO_2297 (O_2297,N_19613,N_19662);
or UO_2298 (O_2298,N_19987,N_19799);
nor UO_2299 (O_2299,N_19814,N_19701);
or UO_2300 (O_2300,N_19865,N_19951);
and UO_2301 (O_2301,N_19812,N_19680);
xor UO_2302 (O_2302,N_19836,N_19770);
or UO_2303 (O_2303,N_19683,N_19791);
nor UO_2304 (O_2304,N_19741,N_19683);
or UO_2305 (O_2305,N_19610,N_19719);
or UO_2306 (O_2306,N_19923,N_19722);
or UO_2307 (O_2307,N_19611,N_19983);
nor UO_2308 (O_2308,N_19840,N_19812);
nand UO_2309 (O_2309,N_19698,N_19759);
or UO_2310 (O_2310,N_19833,N_19829);
and UO_2311 (O_2311,N_19634,N_19617);
nor UO_2312 (O_2312,N_19669,N_19620);
xor UO_2313 (O_2313,N_19806,N_19904);
nor UO_2314 (O_2314,N_19973,N_19653);
nand UO_2315 (O_2315,N_19694,N_19643);
or UO_2316 (O_2316,N_19993,N_19791);
xor UO_2317 (O_2317,N_19866,N_19844);
and UO_2318 (O_2318,N_19652,N_19667);
nor UO_2319 (O_2319,N_19812,N_19914);
nand UO_2320 (O_2320,N_19660,N_19635);
xnor UO_2321 (O_2321,N_19932,N_19961);
and UO_2322 (O_2322,N_19924,N_19911);
or UO_2323 (O_2323,N_19857,N_19802);
nor UO_2324 (O_2324,N_19821,N_19837);
or UO_2325 (O_2325,N_19815,N_19646);
nor UO_2326 (O_2326,N_19695,N_19983);
nor UO_2327 (O_2327,N_19759,N_19749);
nand UO_2328 (O_2328,N_19966,N_19832);
and UO_2329 (O_2329,N_19925,N_19957);
nor UO_2330 (O_2330,N_19912,N_19935);
and UO_2331 (O_2331,N_19648,N_19871);
or UO_2332 (O_2332,N_19870,N_19978);
nand UO_2333 (O_2333,N_19926,N_19881);
nor UO_2334 (O_2334,N_19627,N_19963);
nand UO_2335 (O_2335,N_19805,N_19922);
xnor UO_2336 (O_2336,N_19997,N_19701);
xnor UO_2337 (O_2337,N_19823,N_19679);
nand UO_2338 (O_2338,N_19924,N_19755);
nand UO_2339 (O_2339,N_19845,N_19692);
and UO_2340 (O_2340,N_19873,N_19986);
or UO_2341 (O_2341,N_19960,N_19627);
nand UO_2342 (O_2342,N_19951,N_19779);
and UO_2343 (O_2343,N_19928,N_19875);
nor UO_2344 (O_2344,N_19718,N_19884);
nor UO_2345 (O_2345,N_19674,N_19955);
xor UO_2346 (O_2346,N_19721,N_19953);
and UO_2347 (O_2347,N_19913,N_19826);
nand UO_2348 (O_2348,N_19718,N_19932);
nand UO_2349 (O_2349,N_19707,N_19780);
and UO_2350 (O_2350,N_19620,N_19892);
or UO_2351 (O_2351,N_19670,N_19874);
nor UO_2352 (O_2352,N_19770,N_19999);
xnor UO_2353 (O_2353,N_19728,N_19975);
xor UO_2354 (O_2354,N_19961,N_19813);
or UO_2355 (O_2355,N_19710,N_19642);
xnor UO_2356 (O_2356,N_19950,N_19662);
nor UO_2357 (O_2357,N_19721,N_19658);
nor UO_2358 (O_2358,N_19799,N_19935);
or UO_2359 (O_2359,N_19848,N_19859);
xor UO_2360 (O_2360,N_19809,N_19779);
or UO_2361 (O_2361,N_19761,N_19718);
nand UO_2362 (O_2362,N_19603,N_19976);
nor UO_2363 (O_2363,N_19809,N_19769);
or UO_2364 (O_2364,N_19999,N_19816);
xnor UO_2365 (O_2365,N_19665,N_19841);
nand UO_2366 (O_2366,N_19656,N_19923);
xnor UO_2367 (O_2367,N_19737,N_19955);
or UO_2368 (O_2368,N_19692,N_19764);
or UO_2369 (O_2369,N_19654,N_19803);
xnor UO_2370 (O_2370,N_19741,N_19882);
nor UO_2371 (O_2371,N_19947,N_19799);
xor UO_2372 (O_2372,N_19975,N_19772);
xor UO_2373 (O_2373,N_19984,N_19692);
nand UO_2374 (O_2374,N_19693,N_19916);
and UO_2375 (O_2375,N_19890,N_19841);
and UO_2376 (O_2376,N_19787,N_19929);
or UO_2377 (O_2377,N_19776,N_19999);
and UO_2378 (O_2378,N_19958,N_19767);
and UO_2379 (O_2379,N_19692,N_19613);
xnor UO_2380 (O_2380,N_19868,N_19691);
or UO_2381 (O_2381,N_19905,N_19612);
or UO_2382 (O_2382,N_19652,N_19784);
nor UO_2383 (O_2383,N_19972,N_19662);
or UO_2384 (O_2384,N_19675,N_19674);
or UO_2385 (O_2385,N_19802,N_19778);
and UO_2386 (O_2386,N_19704,N_19669);
xnor UO_2387 (O_2387,N_19665,N_19772);
and UO_2388 (O_2388,N_19995,N_19937);
or UO_2389 (O_2389,N_19956,N_19968);
nand UO_2390 (O_2390,N_19965,N_19978);
nor UO_2391 (O_2391,N_19949,N_19825);
nand UO_2392 (O_2392,N_19998,N_19822);
xnor UO_2393 (O_2393,N_19894,N_19633);
nand UO_2394 (O_2394,N_19789,N_19948);
nor UO_2395 (O_2395,N_19622,N_19773);
and UO_2396 (O_2396,N_19998,N_19946);
xor UO_2397 (O_2397,N_19933,N_19800);
xor UO_2398 (O_2398,N_19644,N_19703);
nand UO_2399 (O_2399,N_19755,N_19851);
xor UO_2400 (O_2400,N_19609,N_19954);
and UO_2401 (O_2401,N_19732,N_19980);
nand UO_2402 (O_2402,N_19903,N_19643);
or UO_2403 (O_2403,N_19820,N_19810);
xor UO_2404 (O_2404,N_19665,N_19703);
or UO_2405 (O_2405,N_19852,N_19645);
xor UO_2406 (O_2406,N_19824,N_19812);
or UO_2407 (O_2407,N_19780,N_19790);
nor UO_2408 (O_2408,N_19633,N_19690);
nand UO_2409 (O_2409,N_19810,N_19802);
xor UO_2410 (O_2410,N_19864,N_19667);
or UO_2411 (O_2411,N_19845,N_19731);
xor UO_2412 (O_2412,N_19730,N_19767);
or UO_2413 (O_2413,N_19962,N_19892);
or UO_2414 (O_2414,N_19742,N_19969);
nor UO_2415 (O_2415,N_19979,N_19693);
nor UO_2416 (O_2416,N_19764,N_19617);
nand UO_2417 (O_2417,N_19785,N_19907);
or UO_2418 (O_2418,N_19907,N_19846);
and UO_2419 (O_2419,N_19847,N_19894);
xnor UO_2420 (O_2420,N_19768,N_19749);
nor UO_2421 (O_2421,N_19686,N_19986);
or UO_2422 (O_2422,N_19865,N_19881);
xor UO_2423 (O_2423,N_19870,N_19728);
nor UO_2424 (O_2424,N_19990,N_19922);
and UO_2425 (O_2425,N_19808,N_19962);
nand UO_2426 (O_2426,N_19775,N_19746);
nor UO_2427 (O_2427,N_19772,N_19807);
and UO_2428 (O_2428,N_19943,N_19640);
nor UO_2429 (O_2429,N_19916,N_19869);
and UO_2430 (O_2430,N_19602,N_19871);
xnor UO_2431 (O_2431,N_19845,N_19710);
nand UO_2432 (O_2432,N_19832,N_19961);
nand UO_2433 (O_2433,N_19809,N_19714);
xnor UO_2434 (O_2434,N_19645,N_19693);
or UO_2435 (O_2435,N_19924,N_19873);
nor UO_2436 (O_2436,N_19615,N_19973);
xor UO_2437 (O_2437,N_19998,N_19912);
and UO_2438 (O_2438,N_19776,N_19985);
nand UO_2439 (O_2439,N_19824,N_19656);
and UO_2440 (O_2440,N_19911,N_19690);
nor UO_2441 (O_2441,N_19600,N_19829);
nand UO_2442 (O_2442,N_19792,N_19811);
nor UO_2443 (O_2443,N_19807,N_19638);
xor UO_2444 (O_2444,N_19923,N_19853);
xnor UO_2445 (O_2445,N_19816,N_19959);
nand UO_2446 (O_2446,N_19863,N_19804);
or UO_2447 (O_2447,N_19829,N_19830);
or UO_2448 (O_2448,N_19653,N_19680);
and UO_2449 (O_2449,N_19658,N_19881);
nor UO_2450 (O_2450,N_19759,N_19746);
xnor UO_2451 (O_2451,N_19651,N_19751);
nor UO_2452 (O_2452,N_19840,N_19727);
and UO_2453 (O_2453,N_19720,N_19626);
nand UO_2454 (O_2454,N_19785,N_19650);
xnor UO_2455 (O_2455,N_19805,N_19806);
or UO_2456 (O_2456,N_19658,N_19843);
or UO_2457 (O_2457,N_19919,N_19964);
and UO_2458 (O_2458,N_19973,N_19868);
or UO_2459 (O_2459,N_19651,N_19676);
nor UO_2460 (O_2460,N_19781,N_19724);
and UO_2461 (O_2461,N_19624,N_19719);
xnor UO_2462 (O_2462,N_19791,N_19710);
nand UO_2463 (O_2463,N_19742,N_19941);
xnor UO_2464 (O_2464,N_19656,N_19871);
nor UO_2465 (O_2465,N_19801,N_19785);
xor UO_2466 (O_2466,N_19612,N_19711);
or UO_2467 (O_2467,N_19784,N_19623);
nand UO_2468 (O_2468,N_19719,N_19815);
nor UO_2469 (O_2469,N_19908,N_19627);
and UO_2470 (O_2470,N_19980,N_19715);
and UO_2471 (O_2471,N_19879,N_19717);
xnor UO_2472 (O_2472,N_19718,N_19625);
or UO_2473 (O_2473,N_19745,N_19860);
nor UO_2474 (O_2474,N_19661,N_19856);
nand UO_2475 (O_2475,N_19866,N_19806);
and UO_2476 (O_2476,N_19607,N_19830);
or UO_2477 (O_2477,N_19991,N_19853);
nor UO_2478 (O_2478,N_19845,N_19775);
nand UO_2479 (O_2479,N_19659,N_19960);
or UO_2480 (O_2480,N_19903,N_19877);
xor UO_2481 (O_2481,N_19934,N_19672);
xor UO_2482 (O_2482,N_19870,N_19897);
and UO_2483 (O_2483,N_19805,N_19701);
nor UO_2484 (O_2484,N_19933,N_19846);
xnor UO_2485 (O_2485,N_19655,N_19714);
nand UO_2486 (O_2486,N_19976,N_19767);
and UO_2487 (O_2487,N_19752,N_19706);
xor UO_2488 (O_2488,N_19999,N_19668);
or UO_2489 (O_2489,N_19825,N_19817);
xor UO_2490 (O_2490,N_19723,N_19703);
or UO_2491 (O_2491,N_19839,N_19625);
xor UO_2492 (O_2492,N_19913,N_19992);
nor UO_2493 (O_2493,N_19772,N_19783);
nand UO_2494 (O_2494,N_19677,N_19869);
nor UO_2495 (O_2495,N_19644,N_19775);
xnor UO_2496 (O_2496,N_19900,N_19803);
or UO_2497 (O_2497,N_19834,N_19912);
xnor UO_2498 (O_2498,N_19879,N_19800);
xor UO_2499 (O_2499,N_19635,N_19684);
endmodule