module basic_750_5000_1000_50_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_216,In_293);
and U1 (N_1,In_33,In_200);
nand U2 (N_2,In_8,In_307);
and U3 (N_3,In_591,In_692);
xnor U4 (N_4,In_31,In_537);
nand U5 (N_5,In_746,In_413);
nor U6 (N_6,In_109,In_674);
nand U7 (N_7,In_618,In_539);
nor U8 (N_8,In_503,In_191);
and U9 (N_9,In_96,In_261);
nand U10 (N_10,In_641,In_323);
xor U11 (N_11,In_246,In_226);
or U12 (N_12,In_207,In_110);
xnor U13 (N_13,In_352,In_172);
xor U14 (N_14,In_556,In_648);
and U15 (N_15,In_277,In_297);
xor U16 (N_16,In_138,In_568);
and U17 (N_17,In_533,In_37);
and U18 (N_18,In_462,In_131);
nor U19 (N_19,In_504,In_256);
xnor U20 (N_20,In_466,In_468);
nor U21 (N_21,In_624,In_174);
and U22 (N_22,In_565,In_40);
nand U23 (N_23,In_278,In_74);
xor U24 (N_24,In_600,In_638);
and U25 (N_25,In_558,In_672);
and U26 (N_26,In_235,In_108);
nor U27 (N_27,In_369,In_64);
nand U28 (N_28,In_727,In_419);
and U29 (N_29,In_385,In_481);
xnor U30 (N_30,In_378,In_421);
nand U31 (N_31,In_720,In_527);
xor U32 (N_32,In_711,In_264);
xor U33 (N_33,In_268,In_405);
nand U34 (N_34,In_670,In_717);
or U35 (N_35,In_185,In_382);
nand U36 (N_36,In_347,In_322);
xnor U37 (N_37,In_585,In_328);
xnor U38 (N_38,In_222,In_463);
nand U39 (N_39,In_669,In_286);
nor U40 (N_40,In_240,In_687);
or U41 (N_41,In_281,In_491);
or U42 (N_42,In_11,In_554);
xnor U43 (N_43,In_160,In_380);
or U44 (N_44,In_306,In_374);
and U45 (N_45,In_302,In_735);
and U46 (N_46,In_335,In_141);
nor U47 (N_47,In_195,In_742);
nand U48 (N_48,In_87,In_267);
xnor U49 (N_49,In_423,In_171);
nor U50 (N_50,In_162,In_528);
and U51 (N_51,In_694,In_697);
or U52 (N_52,In_215,In_633);
nand U53 (N_53,In_471,In_204);
and U54 (N_54,In_111,In_346);
and U55 (N_55,In_148,In_315);
or U56 (N_56,In_234,In_397);
nand U57 (N_57,In_353,In_379);
and U58 (N_58,In_80,In_209);
nand U59 (N_59,In_337,In_124);
nand U60 (N_60,In_258,In_310);
nor U61 (N_61,In_744,In_154);
nand U62 (N_62,In_57,In_407);
or U63 (N_63,In_688,In_545);
and U64 (N_64,In_390,In_26);
nand U65 (N_65,In_440,In_400);
xnor U66 (N_66,In_68,In_683);
and U67 (N_67,In_479,In_701);
nand U68 (N_68,In_476,In_112);
and U69 (N_69,In_381,In_88);
xor U70 (N_70,In_737,In_182);
nand U71 (N_71,In_354,In_709);
or U72 (N_72,In_581,In_675);
xor U73 (N_73,In_645,In_16);
or U74 (N_74,In_355,In_333);
or U75 (N_75,In_738,In_576);
and U76 (N_76,In_516,In_401);
nand U77 (N_77,In_309,In_329);
xnor U78 (N_78,In_43,In_34);
nor U79 (N_79,In_1,In_298);
nand U80 (N_80,In_480,In_599);
nor U81 (N_81,In_231,In_395);
or U82 (N_82,In_699,In_220);
nand U83 (N_83,In_497,In_289);
or U84 (N_84,In_540,In_54);
xor U85 (N_85,In_358,In_649);
xor U86 (N_86,In_56,In_529);
and U87 (N_87,In_534,In_320);
xor U88 (N_88,In_336,In_399);
or U89 (N_89,In_45,In_577);
nor U90 (N_90,In_630,In_501);
and U91 (N_91,In_150,In_729);
and U92 (N_92,In_582,In_520);
and U93 (N_93,In_588,In_144);
nor U94 (N_94,In_460,In_509);
xnor U95 (N_95,In_183,In_560);
nor U96 (N_96,In_485,In_607);
xnor U97 (N_97,In_636,In_189);
nor U98 (N_98,In_3,In_44);
or U99 (N_99,In_23,In_2);
nand U100 (N_100,In_728,In_69);
xnor U101 (N_101,In_304,In_133);
xor U102 (N_102,In_324,In_175);
or U103 (N_103,In_187,In_619);
or U104 (N_104,In_660,In_237);
nand U105 (N_105,N_73,In_656);
xor U106 (N_106,In_272,In_500);
nand U107 (N_107,N_58,N_25);
and U108 (N_108,In_538,In_444);
nand U109 (N_109,In_548,In_430);
nand U110 (N_110,In_224,N_3);
nor U111 (N_111,In_622,In_211);
nand U112 (N_112,In_251,In_357);
nor U113 (N_113,In_127,In_487);
nor U114 (N_114,In_27,N_72);
and U115 (N_115,In_655,In_680);
and U116 (N_116,In_135,N_24);
nand U117 (N_117,In_280,In_523);
nand U118 (N_118,In_55,In_242);
and U119 (N_119,In_79,In_257);
nor U120 (N_120,In_105,In_370);
and U121 (N_121,In_446,In_426);
nand U122 (N_122,In_208,In_349);
xnor U123 (N_123,In_488,In_412);
nand U124 (N_124,In_75,In_291);
or U125 (N_125,In_104,N_43);
or U126 (N_126,In_679,In_388);
nor U127 (N_127,In_731,In_61);
nor U128 (N_128,In_602,In_132);
or U129 (N_129,N_29,In_348);
nand U130 (N_130,In_586,In_326);
nor U131 (N_131,In_4,In_708);
or U132 (N_132,In_72,In_39);
xor U133 (N_133,In_563,In_723);
and U134 (N_134,In_252,N_53);
nand U135 (N_135,In_404,N_28);
or U136 (N_136,In_495,In_254);
xnor U137 (N_137,In_681,In_194);
nor U138 (N_138,N_98,In_572);
nor U139 (N_139,N_85,N_35);
and U140 (N_140,In_305,In_312);
nand U141 (N_141,In_682,N_4);
xnor U142 (N_142,N_56,In_89);
nor U143 (N_143,In_288,In_179);
and U144 (N_144,In_351,In_719);
or U145 (N_145,In_51,In_574);
and U146 (N_146,In_263,In_238);
and U147 (N_147,N_12,In_70);
xnor U148 (N_148,In_259,N_6);
xor U149 (N_149,In_580,In_695);
nand U150 (N_150,In_749,In_95);
nand U151 (N_151,In_654,In_244);
or U152 (N_152,In_592,In_9);
and U153 (N_153,In_543,In_700);
nor U154 (N_154,In_167,In_415);
nand U155 (N_155,N_5,In_196);
nand U156 (N_156,In_696,In_253);
nand U157 (N_157,In_340,In_170);
nand U158 (N_158,In_389,In_436);
nor U159 (N_159,In_546,N_38);
or U160 (N_160,In_76,N_71);
nor U161 (N_161,In_623,In_705);
nand U162 (N_162,N_69,In_443);
or U163 (N_163,In_726,N_95);
nand U164 (N_164,In_601,In_646);
xnor U165 (N_165,In_120,In_375);
xor U166 (N_166,N_60,In_512);
nor U167 (N_167,In_663,In_373);
nand U168 (N_168,In_589,In_279);
nor U169 (N_169,N_39,In_707);
and U170 (N_170,In_459,In_608);
xnor U171 (N_171,N_0,In_386);
or U172 (N_172,In_526,In_439);
nor U173 (N_173,N_1,In_557);
or U174 (N_174,In_248,In_221);
nor U175 (N_175,In_684,In_483);
nand U176 (N_176,In_327,In_217);
or U177 (N_177,In_308,N_82);
or U178 (N_178,In_603,In_106);
or U179 (N_179,In_46,N_7);
nand U180 (N_180,N_52,In_651);
and U181 (N_181,In_671,In_584);
nor U182 (N_182,N_14,In_712);
nor U183 (N_183,In_275,In_561);
or U184 (N_184,In_145,In_83);
xnor U185 (N_185,In_489,In_449);
nand U186 (N_186,In_102,In_676);
xor U187 (N_187,In_693,N_77);
or U188 (N_188,In_566,In_420);
nor U189 (N_189,N_89,In_361);
nor U190 (N_190,In_610,In_409);
xnor U191 (N_191,In_153,In_285);
nand U192 (N_192,In_721,N_94);
and U193 (N_193,In_35,In_318);
nor U194 (N_194,In_21,In_716);
nor U195 (N_195,In_428,In_225);
or U196 (N_196,In_303,In_559);
xor U197 (N_197,N_47,In_245);
and U198 (N_198,In_621,In_213);
and U199 (N_199,In_255,In_416);
and U200 (N_200,N_160,In_58);
and U201 (N_201,In_32,N_172);
nor U202 (N_202,In_311,N_62);
and U203 (N_203,In_658,In_178);
or U204 (N_204,In_435,In_198);
and U205 (N_205,N_142,N_26);
nor U206 (N_206,In_472,In_233);
xor U207 (N_207,In_274,In_223);
xnor U208 (N_208,In_722,In_437);
xnor U209 (N_209,In_117,N_10);
and U210 (N_210,In_90,In_343);
and U211 (N_211,N_9,N_108);
nor U212 (N_212,In_743,In_492);
or U213 (N_213,In_524,In_344);
nor U214 (N_214,In_19,In_486);
nand U215 (N_215,N_110,N_170);
xnor U216 (N_216,In_521,N_75);
nand U217 (N_217,In_301,N_151);
xor U218 (N_218,In_15,N_74);
nor U219 (N_219,In_550,In_113);
nand U220 (N_220,In_456,In_639);
nand U221 (N_221,N_162,N_45);
nand U222 (N_222,N_147,In_5);
xor U223 (N_223,In_575,In_640);
and U224 (N_224,N_104,In_249);
nor U225 (N_225,In_535,N_64);
nand U226 (N_226,N_42,N_78);
xnor U227 (N_227,N_46,In_186);
and U228 (N_228,In_232,In_66);
nand U229 (N_229,In_482,In_92);
or U230 (N_230,In_445,In_473);
xor U231 (N_231,N_156,In_202);
and U232 (N_232,N_116,In_690);
nand U233 (N_233,N_102,In_715);
nor U234 (N_234,N_113,In_101);
or U235 (N_235,In_734,N_59);
or U236 (N_236,N_57,N_158);
nand U237 (N_237,In_201,In_71);
nor U238 (N_238,In_632,N_67);
and U239 (N_239,N_61,In_625);
xor U240 (N_240,In_531,N_111);
nor U241 (N_241,In_241,N_84);
xor U242 (N_242,In_562,In_522);
and U243 (N_243,In_123,N_92);
and U244 (N_244,In_14,In_551);
xnor U245 (N_245,N_37,N_83);
xor U246 (N_246,In_530,In_93);
or U247 (N_247,In_611,In_316);
and U248 (N_248,In_338,N_198);
xnor U249 (N_249,In_166,In_447);
xnor U250 (N_250,In_136,In_142);
nor U251 (N_251,In_702,N_121);
nor U252 (N_252,In_13,In_129);
or U253 (N_253,In_490,N_161);
and U254 (N_254,N_36,N_32);
nand U255 (N_255,N_114,N_23);
nor U256 (N_256,In_156,N_140);
xnor U257 (N_257,In_161,In_685);
xnor U258 (N_258,In_432,In_270);
xor U259 (N_259,In_642,N_178);
or U260 (N_260,In_49,In_615);
or U261 (N_261,In_152,N_128);
or U262 (N_262,In_745,In_555);
nand U263 (N_263,N_131,In_260);
nor U264 (N_264,In_714,In_553);
or U265 (N_265,N_164,In_461);
nand U266 (N_266,N_11,In_100);
or U267 (N_267,N_120,N_189);
and U268 (N_268,In_544,N_154);
nor U269 (N_269,In_6,In_330);
or U270 (N_270,In_292,N_148);
xor U271 (N_271,In_396,In_192);
and U272 (N_272,In_24,In_125);
nor U273 (N_273,N_177,In_314);
nor U274 (N_274,In_299,In_514);
nor U275 (N_275,In_571,N_139);
and U276 (N_276,In_653,In_620);
nor U277 (N_277,N_144,In_143);
xor U278 (N_278,In_391,In_718);
nor U279 (N_279,In_659,In_36);
xor U280 (N_280,In_747,In_507);
nand U281 (N_281,In_18,In_469);
xnor U282 (N_282,In_63,In_350);
or U283 (N_283,In_210,N_48);
and U284 (N_284,In_730,In_371);
nor U285 (N_285,In_376,In_85);
and U286 (N_286,In_668,In_441);
nor U287 (N_287,In_450,N_93);
nor U288 (N_288,N_186,In_403);
nor U289 (N_289,In_10,In_107);
nor U290 (N_290,In_139,In_29);
nand U291 (N_291,In_243,N_133);
xnor U292 (N_292,N_41,In_661);
nor U293 (N_293,In_290,In_230);
nand U294 (N_294,N_149,N_19);
xnor U295 (N_295,In_703,In_205);
and U296 (N_296,N_192,In_184);
nor U297 (N_297,N_153,In_236);
nand U298 (N_298,In_146,N_124);
nand U299 (N_299,In_227,In_587);
or U300 (N_300,In_394,In_455);
and U301 (N_301,In_53,N_88);
and U302 (N_302,In_513,In_627);
nand U303 (N_303,In_98,N_49);
nand U304 (N_304,In_366,N_180);
xnor U305 (N_305,N_202,In_331);
and U306 (N_306,In_387,In_541);
or U307 (N_307,N_168,N_97);
or U308 (N_308,In_494,N_33);
or U309 (N_309,N_117,N_276);
or U310 (N_310,N_283,In_402);
or U311 (N_311,N_298,N_15);
or U312 (N_312,In_181,In_159);
xnor U313 (N_313,In_470,In_736);
xnor U314 (N_314,In_519,In_48);
or U315 (N_315,N_236,N_218);
xnor U316 (N_316,N_238,In_38);
nand U317 (N_317,N_253,N_209);
and U318 (N_318,In_282,In_363);
nand U319 (N_319,In_149,In_505);
nand U320 (N_320,N_115,In_22);
and U321 (N_321,N_268,N_227);
nor U322 (N_322,N_27,In_452);
nand U323 (N_323,In_686,N_291);
xor U324 (N_324,In_67,N_219);
or U325 (N_325,N_79,N_81);
and U326 (N_326,In_42,N_240);
nand U327 (N_327,In_62,In_239);
nand U328 (N_328,N_181,In_130);
xnor U329 (N_329,N_263,In_614);
nor U330 (N_330,In_262,N_234);
and U331 (N_331,In_451,In_665);
xor U332 (N_332,In_368,In_266);
xnor U333 (N_333,In_629,N_193);
xnor U334 (N_334,N_100,In_164);
xor U335 (N_335,N_196,In_657);
xor U336 (N_336,In_177,In_30);
and U337 (N_337,In_478,In_594);
nor U338 (N_338,N_86,In_163);
nand U339 (N_339,N_216,In_99);
nor U340 (N_340,In_570,In_276);
nand U341 (N_341,In_103,In_542);
and U342 (N_342,In_84,In_190);
nor U343 (N_343,N_281,N_212);
nand U344 (N_344,N_296,In_453);
nand U345 (N_345,In_28,In_739);
or U346 (N_346,N_91,N_267);
and U347 (N_347,In_97,In_25);
nand U348 (N_348,In_334,In_508);
and U349 (N_349,N_272,N_269);
nand U350 (N_350,In_283,In_713);
xor U351 (N_351,In_583,In_578);
nor U352 (N_352,In_20,N_87);
nor U353 (N_353,In_525,In_339);
or U354 (N_354,In_605,In_91);
and U355 (N_355,N_259,N_132);
nor U356 (N_356,In_496,In_609);
or U357 (N_357,In_532,N_260);
xor U358 (N_358,N_159,N_21);
nand U359 (N_359,N_138,N_54);
xnor U360 (N_360,In_424,In_82);
or U361 (N_361,N_190,N_230);
nor U362 (N_362,In_691,N_119);
or U363 (N_363,In_579,In_332);
or U364 (N_364,In_271,In_273);
nand U365 (N_365,In_60,In_457);
nand U366 (N_366,N_182,N_166);
xnor U367 (N_367,N_65,In_287);
and U368 (N_368,N_195,In_408);
nand U369 (N_369,N_251,N_90);
nand U370 (N_370,N_107,N_130);
and U371 (N_371,In_199,In_81);
xnor U372 (N_372,N_210,N_235);
nor U373 (N_373,N_217,In_362);
nor U374 (N_374,N_125,N_280);
xor U375 (N_375,In_590,N_290);
or U376 (N_376,In_269,In_536);
nor U377 (N_377,N_106,In_626);
nand U378 (N_378,In_429,N_279);
and U379 (N_379,In_73,N_208);
or U380 (N_380,N_292,N_213);
xor U381 (N_381,In_17,In_212);
and U382 (N_382,In_612,In_422);
xor U383 (N_383,In_484,In_733);
nand U384 (N_384,In_417,In_398);
or U385 (N_385,N_101,In_502);
nand U386 (N_386,N_297,In_511);
and U387 (N_387,In_549,N_220);
and U388 (N_388,In_128,In_662);
xor U389 (N_389,In_114,N_275);
nor U390 (N_390,In_342,In_477);
nor U391 (N_391,N_265,In_325);
and U392 (N_392,N_225,N_145);
nor U393 (N_393,N_243,In_115);
and U394 (N_394,N_40,In_664);
and U395 (N_395,In_377,N_22);
xnor U396 (N_396,In_433,In_673);
nor U397 (N_397,N_266,In_365);
nand U398 (N_398,In_510,In_203);
or U399 (N_399,N_55,In_265);
nand U400 (N_400,N_229,In_547);
or U401 (N_401,N_308,In_740);
xnor U402 (N_402,N_335,N_322);
nor U403 (N_403,In_157,N_163);
nand U404 (N_404,N_303,In_228);
nand U405 (N_405,In_442,N_381);
nand U406 (N_406,N_214,N_314);
and U407 (N_407,In_168,N_262);
and U408 (N_408,In_597,N_18);
and U409 (N_409,N_362,N_174);
nor U410 (N_410,N_364,In_41);
or U411 (N_411,N_379,In_515);
xor U412 (N_412,N_169,N_380);
or U413 (N_413,N_337,N_350);
nor U414 (N_414,N_359,N_301);
and U415 (N_415,N_248,N_317);
and U416 (N_416,N_109,In_474);
nand U417 (N_417,In_119,N_336);
nor U418 (N_418,N_320,N_30);
nor U419 (N_419,N_309,N_171);
nand U420 (N_420,N_331,In_188);
nand U421 (N_421,In_438,N_2);
xnor U422 (N_422,N_273,In_604);
nand U423 (N_423,N_261,N_304);
and U424 (N_424,In_313,In_180);
or U425 (N_425,In_724,N_370);
or U426 (N_426,In_725,N_173);
xor U427 (N_427,N_288,N_390);
xor U428 (N_428,In_598,N_256);
nor U429 (N_429,In_193,In_499);
or U430 (N_430,In_126,N_387);
nand U431 (N_431,In_411,N_398);
and U432 (N_432,In_666,N_211);
xor U433 (N_433,N_325,N_231);
and U434 (N_434,N_328,In_606);
nor U435 (N_435,N_306,In_0);
or U436 (N_436,In_569,In_635);
nand U437 (N_437,In_321,N_17);
xor U438 (N_438,N_254,In_165);
nor U439 (N_439,In_706,In_151);
nand U440 (N_440,N_315,N_237);
xnor U441 (N_441,N_185,N_63);
or U442 (N_442,In_383,In_140);
or U443 (N_443,N_318,N_126);
or U444 (N_444,N_374,N_361);
nand U445 (N_445,In_506,In_137);
nand U446 (N_446,In_704,N_76);
xor U447 (N_447,N_228,N_352);
or U448 (N_448,N_369,N_226);
and U449 (N_449,In_284,N_233);
or U450 (N_450,N_310,In_667);
xnor U451 (N_451,N_252,In_206);
or U452 (N_452,N_396,N_284);
nor U453 (N_453,N_242,In_341);
or U454 (N_454,N_287,In_631);
or U455 (N_455,N_199,In_467);
and U456 (N_456,N_112,N_395);
nand U457 (N_457,In_741,N_191);
or U458 (N_458,N_353,In_359);
and U459 (N_459,In_493,N_319);
xnor U460 (N_460,In_732,N_333);
and U461 (N_461,N_241,N_203);
or U462 (N_462,In_372,N_385);
and U463 (N_463,N_313,N_293);
and U464 (N_464,In_698,N_224);
and U465 (N_465,In_643,N_299);
and U466 (N_466,N_295,N_285);
xor U467 (N_467,N_244,In_122);
and U468 (N_468,In_613,N_80);
nand U469 (N_469,N_305,In_59);
xnor U470 (N_470,N_270,N_146);
or U471 (N_471,N_187,N_68);
xor U472 (N_472,In_596,N_70);
and U473 (N_473,N_339,In_295);
and U474 (N_474,In_47,N_340);
nor U475 (N_475,In_116,In_393);
and U476 (N_476,N_105,N_134);
xor U477 (N_477,In_434,N_363);
nand U478 (N_478,N_345,N_344);
nor U479 (N_479,N_136,N_311);
nand U480 (N_480,N_356,In_748);
or U481 (N_481,In_458,In_427);
nor U482 (N_482,In_517,N_391);
xnor U483 (N_483,In_317,N_143);
xnor U484 (N_484,In_431,N_367);
or U485 (N_485,In_78,In_425);
nor U486 (N_486,N_373,N_348);
nand U487 (N_487,N_223,N_330);
and U488 (N_488,N_232,In_637);
or U489 (N_489,N_13,N_397);
nor U490 (N_490,In_628,In_647);
or U491 (N_491,N_99,N_8);
nand U492 (N_492,N_388,In_518);
xnor U493 (N_493,N_264,N_316);
nor U494 (N_494,N_355,N_239);
nor U495 (N_495,N_179,In_319);
nor U496 (N_496,In_677,N_324);
or U497 (N_497,N_155,In_567);
xor U498 (N_498,N_271,In_7);
xor U499 (N_499,N_300,N_375);
nor U500 (N_500,N_433,In_710);
or U501 (N_501,N_389,N_496);
nand U502 (N_502,N_440,In_214);
nand U503 (N_503,N_127,N_383);
xor U504 (N_504,N_429,N_150);
and U505 (N_505,N_349,N_473);
xor U506 (N_506,N_122,N_466);
or U507 (N_507,N_201,N_460);
and U508 (N_508,In_410,N_194);
nand U509 (N_509,In_247,In_294);
and U510 (N_510,N_475,N_34);
nand U511 (N_511,N_498,N_463);
nand U512 (N_512,N_477,In_158);
nand U513 (N_513,N_312,N_386);
nor U514 (N_514,N_494,N_250);
xnor U515 (N_515,N_137,N_278);
nand U516 (N_516,N_222,N_499);
nand U517 (N_517,N_205,N_418);
and U518 (N_518,N_257,In_650);
and U519 (N_519,N_354,N_286);
xnor U520 (N_520,N_200,N_382);
and U521 (N_521,N_403,N_409);
nor U522 (N_522,N_394,N_425);
nand U523 (N_523,N_426,In_678);
xnor U524 (N_524,N_413,N_371);
nor U525 (N_525,N_393,N_338);
or U526 (N_526,N_417,N_407);
or U527 (N_527,N_488,N_470);
xnor U528 (N_528,N_135,N_31);
or U529 (N_529,N_44,N_326);
nand U530 (N_530,N_495,N_294);
xor U531 (N_531,N_368,N_416);
xor U532 (N_532,In_414,N_459);
nor U533 (N_533,N_411,In_384);
xor U534 (N_534,N_377,N_323);
and U535 (N_535,N_410,N_401);
nand U536 (N_536,In_176,In_644);
xnor U537 (N_537,N_432,N_351);
and U538 (N_538,In_77,N_96);
nand U539 (N_539,In_65,N_455);
and U540 (N_540,N_456,In_564);
or U541 (N_541,N_346,N_165);
xnor U542 (N_542,In_356,N_51);
and U543 (N_543,N_255,N_357);
xnor U544 (N_544,In_454,N_342);
nand U545 (N_545,N_497,N_402);
nand U546 (N_546,N_448,N_347);
xor U547 (N_547,N_422,In_418);
nand U548 (N_548,N_480,N_444);
xnor U549 (N_549,N_461,N_221);
xnor U550 (N_550,In_464,N_405);
or U551 (N_551,N_366,N_439);
nor U552 (N_552,N_484,N_157);
xnor U553 (N_553,In_406,N_452);
and U554 (N_554,N_20,N_334);
xor U555 (N_555,N_446,N_176);
nor U556 (N_556,N_436,N_204);
nand U557 (N_557,In_296,N_438);
nand U558 (N_558,N_412,N_454);
or U559 (N_559,N_184,N_360);
and U560 (N_560,N_329,N_490);
or U561 (N_561,N_427,N_453);
nor U562 (N_562,N_129,N_207);
xor U563 (N_563,N_443,N_483);
or U564 (N_564,N_246,N_197);
or U565 (N_565,N_450,N_365);
or U566 (N_566,N_445,In_250);
nand U567 (N_567,In_52,In_12);
and U568 (N_568,N_123,N_378);
and U569 (N_569,In_595,In_169);
nand U570 (N_570,In_367,In_498);
and U571 (N_571,N_341,N_141);
xnor U572 (N_572,N_249,N_167);
nor U573 (N_573,N_332,In_229);
and U574 (N_574,N_282,N_485);
and U575 (N_575,N_482,N_486);
nor U576 (N_576,In_552,N_399);
or U577 (N_577,N_487,N_321);
or U578 (N_578,N_478,N_245);
or U579 (N_579,N_247,In_94);
or U580 (N_580,In_616,N_175);
nor U581 (N_581,N_465,N_458);
and U582 (N_582,In_219,N_423);
or U583 (N_583,N_447,N_415);
nand U584 (N_584,N_188,N_307);
and U585 (N_585,N_472,N_474);
nand U586 (N_586,N_302,N_492);
or U587 (N_587,In_689,N_206);
and U588 (N_588,N_152,N_449);
nand U589 (N_589,N_430,In_345);
and U590 (N_590,In_465,N_215);
and U591 (N_591,N_50,N_421);
or U592 (N_592,N_493,In_118);
or U593 (N_593,N_343,N_431);
nand U594 (N_594,N_384,N_66);
nand U595 (N_595,N_376,N_462);
and U596 (N_596,N_183,N_103);
and U597 (N_597,In_197,In_218);
nor U598 (N_598,In_475,In_86);
or U599 (N_599,N_400,N_471);
and U600 (N_600,N_527,In_634);
nor U601 (N_601,N_550,N_467);
and U602 (N_602,N_569,N_579);
nand U603 (N_603,N_521,N_585);
nand U604 (N_604,N_544,N_500);
or U605 (N_605,N_501,N_506);
nor U606 (N_606,N_570,N_534);
or U607 (N_607,N_591,N_518);
nand U608 (N_608,N_580,N_532);
nor U609 (N_609,In_617,N_575);
and U610 (N_610,In_147,In_155);
xor U611 (N_611,In_652,N_408);
or U612 (N_612,N_520,N_592);
and U613 (N_613,In_448,N_504);
nor U614 (N_614,N_548,N_503);
or U615 (N_615,N_476,N_118);
and U616 (N_616,N_479,N_529);
and U617 (N_617,In_392,N_435);
and U618 (N_618,N_568,N_565);
nor U619 (N_619,In_360,N_593);
xnor U620 (N_620,N_553,N_590);
nor U621 (N_621,N_442,N_567);
nand U622 (N_622,N_538,N_551);
nand U623 (N_623,N_594,N_451);
and U624 (N_624,N_576,In_121);
and U625 (N_625,N_525,N_584);
nand U626 (N_626,N_489,In_300);
and U627 (N_627,N_531,N_556);
nor U628 (N_628,N_563,N_424);
or U629 (N_629,N_533,N_516);
xor U630 (N_630,N_457,N_586);
and U631 (N_631,In_134,N_513);
or U632 (N_632,N_514,N_577);
nand U633 (N_633,N_258,N_571);
xnor U634 (N_634,N_578,N_558);
xnor U635 (N_635,N_566,N_552);
xnor U636 (N_636,N_277,N_540);
nor U637 (N_637,N_528,N_539);
nand U638 (N_638,N_511,N_512);
nor U639 (N_639,N_464,N_559);
nor U640 (N_640,N_524,N_589);
and U641 (N_641,N_510,N_515);
xor U642 (N_642,In_573,N_508);
nor U643 (N_643,N_560,N_572);
and U644 (N_644,N_434,N_530);
nand U645 (N_645,N_505,N_428);
nor U646 (N_646,N_406,In_593);
or U647 (N_647,N_519,In_50);
xnor U648 (N_648,In_173,N_546);
nand U649 (N_649,N_542,N_481);
and U650 (N_650,N_583,N_507);
or U651 (N_651,N_555,N_588);
nand U652 (N_652,N_522,N_526);
xor U653 (N_653,N_595,N_597);
and U654 (N_654,N_392,N_420);
or U655 (N_655,N_372,N_469);
nor U656 (N_656,N_536,N_554);
and U657 (N_657,N_549,N_289);
nand U658 (N_658,N_419,N_414);
nor U659 (N_659,N_557,N_545);
and U660 (N_660,N_581,N_404);
and U661 (N_661,N_441,N_274);
or U662 (N_662,N_573,N_468);
nand U663 (N_663,N_574,N_547);
nor U664 (N_664,N_541,N_582);
or U665 (N_665,N_491,N_502);
and U666 (N_666,N_537,N_16);
nand U667 (N_667,N_437,In_364);
nor U668 (N_668,N_596,N_599);
or U669 (N_669,N_517,N_535);
and U670 (N_670,N_523,N_358);
nand U671 (N_671,N_543,N_327);
nor U672 (N_672,N_587,N_562);
and U673 (N_673,N_598,N_561);
xor U674 (N_674,N_509,N_564);
and U675 (N_675,N_589,N_510);
or U676 (N_676,N_527,N_574);
nand U677 (N_677,N_414,N_527);
or U678 (N_678,In_134,N_451);
nor U679 (N_679,N_522,N_570);
or U680 (N_680,N_502,N_580);
xor U681 (N_681,N_517,N_504);
xor U682 (N_682,N_544,N_590);
xor U683 (N_683,N_567,N_469);
or U684 (N_684,N_525,N_594);
or U685 (N_685,N_557,N_502);
or U686 (N_686,N_468,N_506);
nor U687 (N_687,N_289,N_548);
xor U688 (N_688,N_546,N_575);
or U689 (N_689,N_420,N_515);
nor U690 (N_690,N_481,N_392);
xor U691 (N_691,In_50,N_552);
nor U692 (N_692,N_504,N_520);
nor U693 (N_693,N_505,N_414);
nor U694 (N_694,In_652,N_582);
or U695 (N_695,N_587,N_514);
nand U696 (N_696,N_521,N_441);
nand U697 (N_697,N_555,N_596);
nor U698 (N_698,N_528,N_543);
or U699 (N_699,N_524,N_457);
or U700 (N_700,N_692,N_647);
nand U701 (N_701,N_681,N_651);
nand U702 (N_702,N_653,N_646);
or U703 (N_703,N_677,N_698);
nand U704 (N_704,N_691,N_617);
nand U705 (N_705,N_669,N_637);
nand U706 (N_706,N_609,N_674);
nor U707 (N_707,N_694,N_645);
nand U708 (N_708,N_606,N_630);
nor U709 (N_709,N_643,N_699);
nor U710 (N_710,N_619,N_659);
or U711 (N_711,N_664,N_623);
and U712 (N_712,N_649,N_628);
and U713 (N_713,N_658,N_661);
or U714 (N_714,N_603,N_654);
nor U715 (N_715,N_666,N_679);
or U716 (N_716,N_607,N_673);
nand U717 (N_717,N_693,N_625);
or U718 (N_718,N_686,N_601);
nor U719 (N_719,N_675,N_638);
nand U720 (N_720,N_652,N_634);
or U721 (N_721,N_618,N_621);
and U722 (N_722,N_676,N_672);
or U723 (N_723,N_627,N_690);
and U724 (N_724,N_635,N_656);
nor U725 (N_725,N_695,N_668);
xor U726 (N_726,N_662,N_612);
and U727 (N_727,N_622,N_639);
nand U728 (N_728,N_629,N_608);
nor U729 (N_729,N_650,N_620);
nor U730 (N_730,N_602,N_604);
and U731 (N_731,N_636,N_611);
nand U732 (N_732,N_667,N_688);
and U733 (N_733,N_626,N_697);
nand U734 (N_734,N_670,N_610);
nor U735 (N_735,N_642,N_689);
xor U736 (N_736,N_633,N_665);
nand U737 (N_737,N_678,N_680);
nand U738 (N_738,N_687,N_640);
nor U739 (N_739,N_641,N_663);
and U740 (N_740,N_682,N_615);
or U741 (N_741,N_683,N_684);
and U742 (N_742,N_657,N_671);
and U743 (N_743,N_624,N_632);
xnor U744 (N_744,N_600,N_605);
nor U745 (N_745,N_696,N_660);
xor U746 (N_746,N_616,N_613);
and U747 (N_747,N_631,N_685);
and U748 (N_748,N_655,N_644);
nor U749 (N_749,N_614,N_648);
and U750 (N_750,N_671,N_675);
xnor U751 (N_751,N_657,N_691);
and U752 (N_752,N_600,N_628);
nand U753 (N_753,N_625,N_659);
or U754 (N_754,N_656,N_609);
xor U755 (N_755,N_600,N_660);
and U756 (N_756,N_655,N_683);
nand U757 (N_757,N_677,N_670);
xor U758 (N_758,N_659,N_628);
and U759 (N_759,N_602,N_697);
or U760 (N_760,N_614,N_649);
xor U761 (N_761,N_679,N_604);
nand U762 (N_762,N_674,N_667);
or U763 (N_763,N_699,N_603);
nor U764 (N_764,N_684,N_694);
nor U765 (N_765,N_627,N_683);
nand U766 (N_766,N_683,N_698);
or U767 (N_767,N_639,N_614);
or U768 (N_768,N_684,N_602);
nand U769 (N_769,N_658,N_674);
xor U770 (N_770,N_617,N_696);
or U771 (N_771,N_603,N_658);
xnor U772 (N_772,N_632,N_609);
nor U773 (N_773,N_698,N_664);
xor U774 (N_774,N_682,N_658);
nand U775 (N_775,N_662,N_646);
or U776 (N_776,N_668,N_616);
and U777 (N_777,N_657,N_655);
and U778 (N_778,N_629,N_683);
and U779 (N_779,N_601,N_681);
nand U780 (N_780,N_600,N_651);
or U781 (N_781,N_660,N_619);
xor U782 (N_782,N_625,N_652);
and U783 (N_783,N_622,N_644);
nor U784 (N_784,N_662,N_613);
and U785 (N_785,N_633,N_660);
and U786 (N_786,N_699,N_681);
xor U787 (N_787,N_602,N_625);
xor U788 (N_788,N_639,N_660);
and U789 (N_789,N_644,N_629);
xnor U790 (N_790,N_639,N_682);
nand U791 (N_791,N_697,N_655);
and U792 (N_792,N_654,N_689);
or U793 (N_793,N_600,N_657);
nor U794 (N_794,N_611,N_612);
xnor U795 (N_795,N_636,N_610);
xnor U796 (N_796,N_689,N_695);
xnor U797 (N_797,N_669,N_684);
nor U798 (N_798,N_681,N_619);
xnor U799 (N_799,N_643,N_609);
nand U800 (N_800,N_746,N_721);
or U801 (N_801,N_750,N_710);
or U802 (N_802,N_732,N_772);
nor U803 (N_803,N_742,N_794);
and U804 (N_804,N_740,N_730);
or U805 (N_805,N_759,N_712);
and U806 (N_806,N_773,N_797);
nor U807 (N_807,N_793,N_719);
nand U808 (N_808,N_741,N_702);
nand U809 (N_809,N_766,N_723);
xnor U810 (N_810,N_769,N_782);
and U811 (N_811,N_718,N_745);
or U812 (N_812,N_715,N_765);
nand U813 (N_813,N_787,N_753);
or U814 (N_814,N_798,N_761);
or U815 (N_815,N_703,N_733);
or U816 (N_816,N_704,N_725);
and U817 (N_817,N_735,N_763);
and U818 (N_818,N_711,N_777);
and U819 (N_819,N_713,N_729);
xnor U820 (N_820,N_754,N_736);
or U821 (N_821,N_700,N_714);
nor U822 (N_822,N_778,N_705);
nand U823 (N_823,N_779,N_717);
or U824 (N_824,N_796,N_731);
nand U825 (N_825,N_738,N_774);
nand U826 (N_826,N_748,N_771);
and U827 (N_827,N_764,N_776);
and U828 (N_828,N_784,N_727);
or U829 (N_829,N_783,N_790);
nor U830 (N_830,N_770,N_728);
and U831 (N_831,N_706,N_762);
nand U832 (N_832,N_788,N_708);
nor U833 (N_833,N_707,N_743);
nor U834 (N_834,N_744,N_757);
nand U835 (N_835,N_789,N_758);
xor U836 (N_836,N_747,N_767);
and U837 (N_837,N_709,N_749);
nand U838 (N_838,N_768,N_775);
or U839 (N_839,N_791,N_781);
xor U840 (N_840,N_752,N_751);
and U841 (N_841,N_734,N_739);
nand U842 (N_842,N_756,N_760);
nand U843 (N_843,N_780,N_722);
nor U844 (N_844,N_785,N_724);
xnor U845 (N_845,N_737,N_716);
xor U846 (N_846,N_755,N_701);
and U847 (N_847,N_799,N_786);
or U848 (N_848,N_720,N_726);
xnor U849 (N_849,N_795,N_792);
xnor U850 (N_850,N_731,N_761);
and U851 (N_851,N_761,N_760);
nand U852 (N_852,N_765,N_741);
and U853 (N_853,N_780,N_797);
xor U854 (N_854,N_761,N_701);
and U855 (N_855,N_719,N_734);
and U856 (N_856,N_787,N_750);
xor U857 (N_857,N_747,N_784);
and U858 (N_858,N_746,N_704);
xor U859 (N_859,N_752,N_762);
nor U860 (N_860,N_791,N_797);
xor U861 (N_861,N_732,N_735);
and U862 (N_862,N_791,N_785);
xor U863 (N_863,N_798,N_732);
and U864 (N_864,N_744,N_761);
nor U865 (N_865,N_773,N_799);
nor U866 (N_866,N_737,N_712);
nor U867 (N_867,N_767,N_790);
xor U868 (N_868,N_705,N_716);
or U869 (N_869,N_748,N_774);
xnor U870 (N_870,N_735,N_725);
nor U871 (N_871,N_796,N_789);
or U872 (N_872,N_706,N_790);
and U873 (N_873,N_703,N_739);
nand U874 (N_874,N_760,N_794);
xnor U875 (N_875,N_788,N_721);
xor U876 (N_876,N_710,N_766);
or U877 (N_877,N_750,N_765);
nor U878 (N_878,N_744,N_781);
and U879 (N_879,N_763,N_741);
nor U880 (N_880,N_757,N_771);
nor U881 (N_881,N_764,N_734);
and U882 (N_882,N_718,N_764);
or U883 (N_883,N_733,N_737);
and U884 (N_884,N_759,N_700);
nor U885 (N_885,N_701,N_721);
and U886 (N_886,N_760,N_793);
nor U887 (N_887,N_745,N_706);
or U888 (N_888,N_768,N_702);
nor U889 (N_889,N_738,N_743);
xnor U890 (N_890,N_779,N_766);
or U891 (N_891,N_792,N_780);
or U892 (N_892,N_765,N_786);
and U893 (N_893,N_737,N_747);
xnor U894 (N_894,N_759,N_715);
or U895 (N_895,N_771,N_746);
nor U896 (N_896,N_738,N_740);
nand U897 (N_897,N_709,N_798);
or U898 (N_898,N_795,N_755);
or U899 (N_899,N_730,N_739);
nand U900 (N_900,N_843,N_831);
nand U901 (N_901,N_847,N_826);
or U902 (N_902,N_835,N_870);
xor U903 (N_903,N_882,N_880);
nor U904 (N_904,N_811,N_816);
nor U905 (N_905,N_853,N_829);
nor U906 (N_906,N_866,N_894);
and U907 (N_907,N_838,N_879);
or U908 (N_908,N_846,N_868);
nor U909 (N_909,N_814,N_832);
nand U910 (N_910,N_892,N_807);
nand U911 (N_911,N_839,N_808);
or U912 (N_912,N_803,N_889);
xor U913 (N_913,N_865,N_822);
nor U914 (N_914,N_899,N_810);
or U915 (N_915,N_836,N_898);
nand U916 (N_916,N_888,N_852);
nand U917 (N_917,N_802,N_812);
xor U918 (N_918,N_896,N_821);
and U919 (N_919,N_897,N_881);
or U920 (N_920,N_815,N_817);
xor U921 (N_921,N_884,N_857);
nand U922 (N_922,N_856,N_813);
or U923 (N_923,N_893,N_809);
nor U924 (N_924,N_827,N_873);
nor U925 (N_925,N_891,N_860);
or U926 (N_926,N_850,N_869);
nand U927 (N_927,N_848,N_878);
and U928 (N_928,N_883,N_859);
and U929 (N_929,N_820,N_804);
and U930 (N_930,N_874,N_877);
nand U931 (N_931,N_890,N_819);
xor U932 (N_932,N_841,N_834);
nor U933 (N_933,N_858,N_825);
xor U934 (N_934,N_855,N_872);
nor U935 (N_935,N_800,N_842);
nor U936 (N_936,N_837,N_887);
nor U937 (N_937,N_871,N_849);
nand U938 (N_938,N_885,N_861);
nor U939 (N_939,N_851,N_823);
and U940 (N_940,N_824,N_833);
nand U941 (N_941,N_830,N_801);
or U942 (N_942,N_844,N_854);
nand U943 (N_943,N_876,N_840);
and U944 (N_944,N_805,N_886);
nor U945 (N_945,N_818,N_867);
or U946 (N_946,N_875,N_863);
and U947 (N_947,N_806,N_845);
nor U948 (N_948,N_862,N_828);
or U949 (N_949,N_895,N_864);
and U950 (N_950,N_802,N_860);
xnor U951 (N_951,N_873,N_835);
and U952 (N_952,N_856,N_839);
nor U953 (N_953,N_850,N_875);
nor U954 (N_954,N_808,N_877);
xnor U955 (N_955,N_828,N_847);
xor U956 (N_956,N_815,N_831);
or U957 (N_957,N_855,N_892);
xor U958 (N_958,N_884,N_883);
nand U959 (N_959,N_857,N_807);
or U960 (N_960,N_837,N_843);
nand U961 (N_961,N_816,N_861);
xnor U962 (N_962,N_847,N_885);
nor U963 (N_963,N_866,N_825);
nor U964 (N_964,N_892,N_804);
nor U965 (N_965,N_845,N_820);
or U966 (N_966,N_802,N_845);
xnor U967 (N_967,N_850,N_845);
nand U968 (N_968,N_899,N_863);
nor U969 (N_969,N_854,N_813);
nand U970 (N_970,N_839,N_893);
and U971 (N_971,N_824,N_897);
xnor U972 (N_972,N_812,N_835);
nor U973 (N_973,N_898,N_848);
xnor U974 (N_974,N_859,N_890);
nor U975 (N_975,N_854,N_800);
nand U976 (N_976,N_893,N_888);
nand U977 (N_977,N_833,N_811);
nand U978 (N_978,N_828,N_835);
nand U979 (N_979,N_890,N_879);
or U980 (N_980,N_894,N_812);
nand U981 (N_981,N_891,N_880);
xnor U982 (N_982,N_868,N_855);
xor U983 (N_983,N_845,N_834);
nand U984 (N_984,N_853,N_823);
xnor U985 (N_985,N_826,N_899);
nor U986 (N_986,N_811,N_891);
nand U987 (N_987,N_804,N_874);
xnor U988 (N_988,N_862,N_836);
xor U989 (N_989,N_878,N_881);
xor U990 (N_990,N_810,N_850);
and U991 (N_991,N_828,N_804);
and U992 (N_992,N_851,N_898);
or U993 (N_993,N_878,N_855);
or U994 (N_994,N_853,N_869);
nor U995 (N_995,N_826,N_850);
nor U996 (N_996,N_898,N_825);
and U997 (N_997,N_896,N_863);
nand U998 (N_998,N_819,N_826);
xor U999 (N_999,N_834,N_814);
nand U1000 (N_1000,N_948,N_979);
nor U1001 (N_1001,N_992,N_969);
nor U1002 (N_1002,N_954,N_999);
xnor U1003 (N_1003,N_944,N_964);
nand U1004 (N_1004,N_917,N_961);
xor U1005 (N_1005,N_980,N_913);
nand U1006 (N_1006,N_963,N_972);
nand U1007 (N_1007,N_940,N_930);
nand U1008 (N_1008,N_973,N_978);
nand U1009 (N_1009,N_957,N_971);
nor U1010 (N_1010,N_905,N_931);
nand U1011 (N_1011,N_932,N_991);
nand U1012 (N_1012,N_924,N_958);
nand U1013 (N_1013,N_935,N_970);
nor U1014 (N_1014,N_928,N_995);
nand U1015 (N_1015,N_901,N_989);
nor U1016 (N_1016,N_923,N_916);
and U1017 (N_1017,N_962,N_939);
nand U1018 (N_1018,N_946,N_959);
xnor U1019 (N_1019,N_900,N_919);
or U1020 (N_1020,N_976,N_967);
nor U1021 (N_1021,N_938,N_996);
xor U1022 (N_1022,N_910,N_906);
or U1023 (N_1023,N_912,N_927);
xor U1024 (N_1024,N_987,N_903);
nand U1025 (N_1025,N_918,N_997);
nor U1026 (N_1026,N_926,N_994);
or U1027 (N_1027,N_922,N_952);
nand U1028 (N_1028,N_950,N_929);
xnor U1029 (N_1029,N_909,N_986);
xnor U1030 (N_1030,N_998,N_925);
nor U1031 (N_1031,N_949,N_984);
and U1032 (N_1032,N_947,N_933);
and U1033 (N_1033,N_968,N_902);
and U1034 (N_1034,N_953,N_911);
nor U1035 (N_1035,N_966,N_988);
nand U1036 (N_1036,N_914,N_981);
xnor U1037 (N_1037,N_942,N_907);
nand U1038 (N_1038,N_983,N_951);
nor U1039 (N_1039,N_936,N_965);
or U1040 (N_1040,N_943,N_915);
nand U1041 (N_1041,N_934,N_921);
and U1042 (N_1042,N_975,N_974);
nand U1043 (N_1043,N_920,N_993);
nor U1044 (N_1044,N_982,N_960);
nand U1045 (N_1045,N_977,N_945);
xnor U1046 (N_1046,N_955,N_990);
xor U1047 (N_1047,N_941,N_937);
and U1048 (N_1048,N_908,N_985);
nand U1049 (N_1049,N_904,N_956);
nand U1050 (N_1050,N_996,N_933);
nor U1051 (N_1051,N_974,N_923);
or U1052 (N_1052,N_974,N_987);
nor U1053 (N_1053,N_967,N_907);
or U1054 (N_1054,N_945,N_925);
nor U1055 (N_1055,N_933,N_927);
nor U1056 (N_1056,N_937,N_914);
xor U1057 (N_1057,N_910,N_931);
nand U1058 (N_1058,N_924,N_901);
nor U1059 (N_1059,N_986,N_930);
nor U1060 (N_1060,N_903,N_951);
nor U1061 (N_1061,N_996,N_918);
nand U1062 (N_1062,N_991,N_913);
and U1063 (N_1063,N_941,N_949);
and U1064 (N_1064,N_980,N_952);
and U1065 (N_1065,N_933,N_921);
or U1066 (N_1066,N_986,N_996);
or U1067 (N_1067,N_956,N_991);
and U1068 (N_1068,N_997,N_940);
xor U1069 (N_1069,N_928,N_931);
nor U1070 (N_1070,N_929,N_954);
and U1071 (N_1071,N_978,N_909);
xor U1072 (N_1072,N_991,N_974);
and U1073 (N_1073,N_936,N_951);
or U1074 (N_1074,N_966,N_928);
xnor U1075 (N_1075,N_920,N_964);
or U1076 (N_1076,N_950,N_959);
nand U1077 (N_1077,N_953,N_979);
xor U1078 (N_1078,N_967,N_987);
xnor U1079 (N_1079,N_988,N_918);
xor U1080 (N_1080,N_977,N_960);
nor U1081 (N_1081,N_982,N_909);
nor U1082 (N_1082,N_934,N_915);
xnor U1083 (N_1083,N_925,N_979);
nor U1084 (N_1084,N_907,N_973);
and U1085 (N_1085,N_931,N_912);
nor U1086 (N_1086,N_935,N_929);
and U1087 (N_1087,N_940,N_923);
nand U1088 (N_1088,N_924,N_990);
nor U1089 (N_1089,N_924,N_959);
and U1090 (N_1090,N_920,N_930);
nor U1091 (N_1091,N_934,N_991);
nor U1092 (N_1092,N_930,N_918);
nor U1093 (N_1093,N_998,N_991);
or U1094 (N_1094,N_950,N_934);
xor U1095 (N_1095,N_968,N_931);
or U1096 (N_1096,N_986,N_962);
and U1097 (N_1097,N_941,N_905);
or U1098 (N_1098,N_980,N_987);
xor U1099 (N_1099,N_971,N_970);
and U1100 (N_1100,N_1056,N_1062);
or U1101 (N_1101,N_1001,N_1058);
xor U1102 (N_1102,N_1043,N_1003);
xnor U1103 (N_1103,N_1094,N_1038);
and U1104 (N_1104,N_1080,N_1095);
nor U1105 (N_1105,N_1030,N_1034);
and U1106 (N_1106,N_1021,N_1037);
xor U1107 (N_1107,N_1004,N_1072);
and U1108 (N_1108,N_1020,N_1067);
or U1109 (N_1109,N_1079,N_1013);
nand U1110 (N_1110,N_1077,N_1090);
and U1111 (N_1111,N_1098,N_1089);
and U1112 (N_1112,N_1093,N_1005);
nand U1113 (N_1113,N_1002,N_1018);
xnor U1114 (N_1114,N_1084,N_1039);
nor U1115 (N_1115,N_1099,N_1085);
nor U1116 (N_1116,N_1053,N_1014);
nor U1117 (N_1117,N_1000,N_1012);
nor U1118 (N_1118,N_1009,N_1073);
or U1119 (N_1119,N_1048,N_1031);
nand U1120 (N_1120,N_1060,N_1059);
nor U1121 (N_1121,N_1087,N_1096);
or U1122 (N_1122,N_1025,N_1015);
nor U1123 (N_1123,N_1055,N_1028);
nand U1124 (N_1124,N_1024,N_1049);
nor U1125 (N_1125,N_1081,N_1086);
and U1126 (N_1126,N_1019,N_1076);
and U1127 (N_1127,N_1091,N_1075);
nand U1128 (N_1128,N_1088,N_1016);
nand U1129 (N_1129,N_1032,N_1041);
xnor U1130 (N_1130,N_1082,N_1023);
nor U1131 (N_1131,N_1054,N_1050);
nand U1132 (N_1132,N_1051,N_1042);
xnor U1133 (N_1133,N_1047,N_1070);
nand U1134 (N_1134,N_1045,N_1069);
nand U1135 (N_1135,N_1064,N_1036);
nand U1136 (N_1136,N_1097,N_1022);
nor U1137 (N_1137,N_1006,N_1052);
nor U1138 (N_1138,N_1029,N_1063);
xnor U1139 (N_1139,N_1061,N_1011);
xor U1140 (N_1140,N_1083,N_1017);
nand U1141 (N_1141,N_1057,N_1044);
or U1142 (N_1142,N_1071,N_1066);
nand U1143 (N_1143,N_1026,N_1007);
nand U1144 (N_1144,N_1074,N_1068);
or U1145 (N_1145,N_1092,N_1046);
xnor U1146 (N_1146,N_1008,N_1065);
xor U1147 (N_1147,N_1035,N_1027);
xor U1148 (N_1148,N_1010,N_1078);
and U1149 (N_1149,N_1040,N_1033);
nor U1150 (N_1150,N_1009,N_1024);
xor U1151 (N_1151,N_1033,N_1055);
and U1152 (N_1152,N_1054,N_1043);
nor U1153 (N_1153,N_1090,N_1082);
and U1154 (N_1154,N_1009,N_1010);
nand U1155 (N_1155,N_1029,N_1051);
xnor U1156 (N_1156,N_1062,N_1035);
or U1157 (N_1157,N_1074,N_1072);
nand U1158 (N_1158,N_1093,N_1089);
or U1159 (N_1159,N_1049,N_1099);
nor U1160 (N_1160,N_1023,N_1097);
nor U1161 (N_1161,N_1051,N_1000);
nor U1162 (N_1162,N_1038,N_1089);
nor U1163 (N_1163,N_1079,N_1095);
nand U1164 (N_1164,N_1055,N_1030);
xnor U1165 (N_1165,N_1050,N_1096);
nor U1166 (N_1166,N_1091,N_1067);
nand U1167 (N_1167,N_1067,N_1087);
and U1168 (N_1168,N_1076,N_1027);
nand U1169 (N_1169,N_1051,N_1040);
nand U1170 (N_1170,N_1085,N_1035);
xor U1171 (N_1171,N_1091,N_1016);
nor U1172 (N_1172,N_1084,N_1059);
nor U1173 (N_1173,N_1057,N_1024);
or U1174 (N_1174,N_1025,N_1026);
or U1175 (N_1175,N_1098,N_1002);
nand U1176 (N_1176,N_1030,N_1095);
nor U1177 (N_1177,N_1093,N_1007);
and U1178 (N_1178,N_1040,N_1078);
nor U1179 (N_1179,N_1081,N_1091);
nand U1180 (N_1180,N_1047,N_1064);
xnor U1181 (N_1181,N_1021,N_1000);
nor U1182 (N_1182,N_1030,N_1079);
xor U1183 (N_1183,N_1062,N_1022);
or U1184 (N_1184,N_1004,N_1046);
and U1185 (N_1185,N_1028,N_1042);
or U1186 (N_1186,N_1055,N_1063);
xor U1187 (N_1187,N_1076,N_1031);
or U1188 (N_1188,N_1056,N_1003);
nand U1189 (N_1189,N_1085,N_1078);
and U1190 (N_1190,N_1090,N_1093);
and U1191 (N_1191,N_1092,N_1002);
xor U1192 (N_1192,N_1060,N_1035);
xnor U1193 (N_1193,N_1010,N_1016);
nand U1194 (N_1194,N_1076,N_1036);
nor U1195 (N_1195,N_1029,N_1061);
or U1196 (N_1196,N_1006,N_1065);
xor U1197 (N_1197,N_1036,N_1014);
nor U1198 (N_1198,N_1018,N_1023);
xor U1199 (N_1199,N_1086,N_1082);
and U1200 (N_1200,N_1136,N_1100);
and U1201 (N_1201,N_1123,N_1199);
nand U1202 (N_1202,N_1172,N_1106);
and U1203 (N_1203,N_1135,N_1162);
xnor U1204 (N_1204,N_1117,N_1152);
and U1205 (N_1205,N_1157,N_1145);
nor U1206 (N_1206,N_1104,N_1134);
nand U1207 (N_1207,N_1137,N_1155);
or U1208 (N_1208,N_1146,N_1122);
nor U1209 (N_1209,N_1161,N_1133);
or U1210 (N_1210,N_1120,N_1138);
xor U1211 (N_1211,N_1114,N_1171);
nor U1212 (N_1212,N_1101,N_1175);
nand U1213 (N_1213,N_1143,N_1193);
xnor U1214 (N_1214,N_1197,N_1128);
xor U1215 (N_1215,N_1154,N_1151);
and U1216 (N_1216,N_1125,N_1156);
nand U1217 (N_1217,N_1194,N_1196);
nor U1218 (N_1218,N_1174,N_1164);
and U1219 (N_1219,N_1108,N_1183);
and U1220 (N_1220,N_1195,N_1102);
xor U1221 (N_1221,N_1176,N_1139);
xor U1222 (N_1222,N_1118,N_1181);
nor U1223 (N_1223,N_1112,N_1185);
nand U1224 (N_1224,N_1148,N_1142);
and U1225 (N_1225,N_1173,N_1159);
or U1226 (N_1226,N_1182,N_1153);
nand U1227 (N_1227,N_1187,N_1180);
nand U1228 (N_1228,N_1111,N_1124);
nand U1229 (N_1229,N_1144,N_1158);
or U1230 (N_1230,N_1163,N_1130);
or U1231 (N_1231,N_1177,N_1170);
and U1232 (N_1232,N_1150,N_1103);
xor U1233 (N_1233,N_1166,N_1191);
and U1234 (N_1234,N_1131,N_1160);
and U1235 (N_1235,N_1105,N_1132);
nand U1236 (N_1236,N_1188,N_1198);
nor U1237 (N_1237,N_1113,N_1107);
or U1238 (N_1238,N_1179,N_1110);
and U1239 (N_1239,N_1186,N_1127);
xnor U1240 (N_1240,N_1116,N_1184);
nor U1241 (N_1241,N_1129,N_1190);
or U1242 (N_1242,N_1121,N_1147);
or U1243 (N_1243,N_1168,N_1189);
and U1244 (N_1244,N_1126,N_1149);
nand U1245 (N_1245,N_1115,N_1192);
xnor U1246 (N_1246,N_1169,N_1178);
nand U1247 (N_1247,N_1119,N_1165);
or U1248 (N_1248,N_1109,N_1167);
and U1249 (N_1249,N_1141,N_1140);
xnor U1250 (N_1250,N_1178,N_1139);
xnor U1251 (N_1251,N_1186,N_1155);
nand U1252 (N_1252,N_1173,N_1141);
or U1253 (N_1253,N_1165,N_1145);
nor U1254 (N_1254,N_1148,N_1128);
and U1255 (N_1255,N_1191,N_1147);
and U1256 (N_1256,N_1162,N_1175);
or U1257 (N_1257,N_1101,N_1147);
nor U1258 (N_1258,N_1157,N_1195);
xor U1259 (N_1259,N_1180,N_1100);
nand U1260 (N_1260,N_1192,N_1142);
nor U1261 (N_1261,N_1158,N_1182);
or U1262 (N_1262,N_1197,N_1188);
and U1263 (N_1263,N_1140,N_1195);
xor U1264 (N_1264,N_1175,N_1109);
nor U1265 (N_1265,N_1181,N_1125);
xor U1266 (N_1266,N_1102,N_1146);
nor U1267 (N_1267,N_1170,N_1123);
nand U1268 (N_1268,N_1153,N_1171);
nand U1269 (N_1269,N_1118,N_1107);
or U1270 (N_1270,N_1190,N_1121);
and U1271 (N_1271,N_1151,N_1160);
nand U1272 (N_1272,N_1140,N_1129);
xnor U1273 (N_1273,N_1138,N_1181);
xnor U1274 (N_1274,N_1152,N_1145);
nor U1275 (N_1275,N_1107,N_1170);
xor U1276 (N_1276,N_1142,N_1183);
or U1277 (N_1277,N_1170,N_1110);
nand U1278 (N_1278,N_1154,N_1167);
nand U1279 (N_1279,N_1196,N_1162);
nand U1280 (N_1280,N_1104,N_1160);
or U1281 (N_1281,N_1126,N_1166);
and U1282 (N_1282,N_1168,N_1106);
nor U1283 (N_1283,N_1111,N_1173);
nand U1284 (N_1284,N_1141,N_1106);
and U1285 (N_1285,N_1125,N_1194);
nand U1286 (N_1286,N_1187,N_1129);
xor U1287 (N_1287,N_1173,N_1163);
and U1288 (N_1288,N_1157,N_1125);
xor U1289 (N_1289,N_1144,N_1123);
nand U1290 (N_1290,N_1170,N_1136);
nor U1291 (N_1291,N_1109,N_1140);
nand U1292 (N_1292,N_1181,N_1179);
nor U1293 (N_1293,N_1176,N_1133);
or U1294 (N_1294,N_1131,N_1159);
and U1295 (N_1295,N_1138,N_1147);
and U1296 (N_1296,N_1198,N_1118);
or U1297 (N_1297,N_1144,N_1126);
nor U1298 (N_1298,N_1113,N_1123);
nand U1299 (N_1299,N_1168,N_1112);
nand U1300 (N_1300,N_1286,N_1273);
nand U1301 (N_1301,N_1251,N_1237);
and U1302 (N_1302,N_1229,N_1239);
xnor U1303 (N_1303,N_1247,N_1228);
and U1304 (N_1304,N_1202,N_1253);
or U1305 (N_1305,N_1218,N_1275);
nand U1306 (N_1306,N_1200,N_1249);
xor U1307 (N_1307,N_1285,N_1242);
nand U1308 (N_1308,N_1277,N_1296);
nand U1309 (N_1309,N_1256,N_1283);
nand U1310 (N_1310,N_1222,N_1294);
or U1311 (N_1311,N_1205,N_1209);
nor U1312 (N_1312,N_1244,N_1262);
nand U1313 (N_1313,N_1252,N_1258);
or U1314 (N_1314,N_1264,N_1240);
xor U1315 (N_1315,N_1219,N_1238);
xor U1316 (N_1316,N_1223,N_1267);
nand U1317 (N_1317,N_1214,N_1213);
or U1318 (N_1318,N_1207,N_1203);
or U1319 (N_1319,N_1234,N_1260);
xor U1320 (N_1320,N_1255,N_1276);
and U1321 (N_1321,N_1254,N_1216);
nand U1322 (N_1322,N_1295,N_1243);
nand U1323 (N_1323,N_1280,N_1279);
xor U1324 (N_1324,N_1221,N_1248);
and U1325 (N_1325,N_1261,N_1263);
nor U1326 (N_1326,N_1259,N_1265);
xnor U1327 (N_1327,N_1271,N_1233);
nor U1328 (N_1328,N_1293,N_1212);
and U1329 (N_1329,N_1246,N_1230);
nand U1330 (N_1330,N_1274,N_1288);
or U1331 (N_1331,N_1245,N_1217);
xor U1332 (N_1332,N_1236,N_1266);
and U1333 (N_1333,N_1270,N_1292);
nand U1334 (N_1334,N_1287,N_1284);
and U1335 (N_1335,N_1235,N_1224);
nand U1336 (N_1336,N_1206,N_1298);
nand U1337 (N_1337,N_1268,N_1278);
and U1338 (N_1338,N_1290,N_1225);
nand U1339 (N_1339,N_1204,N_1250);
or U1340 (N_1340,N_1201,N_1232);
nand U1341 (N_1341,N_1210,N_1281);
or U1342 (N_1342,N_1289,N_1215);
or U1343 (N_1343,N_1231,N_1297);
and U1344 (N_1344,N_1299,N_1291);
and U1345 (N_1345,N_1272,N_1220);
and U1346 (N_1346,N_1208,N_1257);
and U1347 (N_1347,N_1211,N_1269);
nor U1348 (N_1348,N_1241,N_1226);
or U1349 (N_1349,N_1282,N_1227);
and U1350 (N_1350,N_1272,N_1295);
and U1351 (N_1351,N_1261,N_1280);
or U1352 (N_1352,N_1252,N_1291);
nand U1353 (N_1353,N_1213,N_1265);
nor U1354 (N_1354,N_1282,N_1262);
xor U1355 (N_1355,N_1263,N_1268);
nand U1356 (N_1356,N_1226,N_1228);
or U1357 (N_1357,N_1219,N_1217);
and U1358 (N_1358,N_1266,N_1271);
nand U1359 (N_1359,N_1270,N_1254);
xnor U1360 (N_1360,N_1207,N_1295);
or U1361 (N_1361,N_1258,N_1249);
and U1362 (N_1362,N_1255,N_1235);
or U1363 (N_1363,N_1275,N_1285);
or U1364 (N_1364,N_1230,N_1259);
and U1365 (N_1365,N_1298,N_1259);
nand U1366 (N_1366,N_1287,N_1242);
xnor U1367 (N_1367,N_1272,N_1286);
nand U1368 (N_1368,N_1261,N_1234);
nor U1369 (N_1369,N_1239,N_1225);
nor U1370 (N_1370,N_1207,N_1263);
nand U1371 (N_1371,N_1236,N_1232);
nor U1372 (N_1372,N_1230,N_1295);
nor U1373 (N_1373,N_1213,N_1293);
xor U1374 (N_1374,N_1216,N_1241);
xor U1375 (N_1375,N_1215,N_1266);
and U1376 (N_1376,N_1251,N_1244);
xnor U1377 (N_1377,N_1211,N_1213);
or U1378 (N_1378,N_1256,N_1232);
and U1379 (N_1379,N_1296,N_1213);
nor U1380 (N_1380,N_1241,N_1286);
nor U1381 (N_1381,N_1274,N_1205);
nand U1382 (N_1382,N_1259,N_1211);
or U1383 (N_1383,N_1272,N_1252);
nand U1384 (N_1384,N_1215,N_1217);
and U1385 (N_1385,N_1233,N_1274);
xor U1386 (N_1386,N_1201,N_1210);
nor U1387 (N_1387,N_1287,N_1228);
xnor U1388 (N_1388,N_1290,N_1269);
or U1389 (N_1389,N_1218,N_1274);
nor U1390 (N_1390,N_1262,N_1290);
nor U1391 (N_1391,N_1235,N_1201);
or U1392 (N_1392,N_1228,N_1204);
nor U1393 (N_1393,N_1289,N_1269);
and U1394 (N_1394,N_1232,N_1202);
xnor U1395 (N_1395,N_1271,N_1298);
nand U1396 (N_1396,N_1201,N_1215);
xnor U1397 (N_1397,N_1259,N_1251);
nor U1398 (N_1398,N_1248,N_1207);
and U1399 (N_1399,N_1221,N_1222);
nand U1400 (N_1400,N_1315,N_1349);
nor U1401 (N_1401,N_1312,N_1356);
and U1402 (N_1402,N_1351,N_1355);
xnor U1403 (N_1403,N_1347,N_1353);
or U1404 (N_1404,N_1332,N_1328);
xor U1405 (N_1405,N_1389,N_1333);
nand U1406 (N_1406,N_1304,N_1343);
nand U1407 (N_1407,N_1399,N_1361);
and U1408 (N_1408,N_1320,N_1324);
nor U1409 (N_1409,N_1314,N_1307);
or U1410 (N_1410,N_1310,N_1377);
nor U1411 (N_1411,N_1301,N_1398);
xnor U1412 (N_1412,N_1388,N_1311);
xnor U1413 (N_1413,N_1372,N_1363);
nand U1414 (N_1414,N_1346,N_1326);
nor U1415 (N_1415,N_1348,N_1316);
or U1416 (N_1416,N_1385,N_1395);
nand U1417 (N_1417,N_1306,N_1382);
nand U1418 (N_1418,N_1336,N_1394);
nand U1419 (N_1419,N_1367,N_1321);
nor U1420 (N_1420,N_1340,N_1325);
nand U1421 (N_1421,N_1327,N_1329);
and U1422 (N_1422,N_1342,N_1335);
xor U1423 (N_1423,N_1302,N_1319);
or U1424 (N_1424,N_1339,N_1368);
nand U1425 (N_1425,N_1397,N_1366);
xnor U1426 (N_1426,N_1323,N_1344);
nor U1427 (N_1427,N_1392,N_1300);
xor U1428 (N_1428,N_1341,N_1345);
and U1429 (N_1429,N_1359,N_1331);
or U1430 (N_1430,N_1358,N_1330);
xnor U1431 (N_1431,N_1373,N_1387);
and U1432 (N_1432,N_1374,N_1393);
nor U1433 (N_1433,N_1309,N_1338);
nand U1434 (N_1434,N_1365,N_1380);
and U1435 (N_1435,N_1390,N_1313);
or U1436 (N_1436,N_1360,N_1334);
xnor U1437 (N_1437,N_1371,N_1383);
nand U1438 (N_1438,N_1379,N_1376);
nand U1439 (N_1439,N_1322,N_1357);
or U1440 (N_1440,N_1317,N_1318);
or U1441 (N_1441,N_1370,N_1369);
and U1442 (N_1442,N_1305,N_1396);
xnor U1443 (N_1443,N_1354,N_1350);
xor U1444 (N_1444,N_1384,N_1303);
nor U1445 (N_1445,N_1391,N_1378);
and U1446 (N_1446,N_1352,N_1337);
nor U1447 (N_1447,N_1308,N_1364);
nor U1448 (N_1448,N_1386,N_1362);
nand U1449 (N_1449,N_1375,N_1381);
and U1450 (N_1450,N_1325,N_1365);
nand U1451 (N_1451,N_1331,N_1372);
nor U1452 (N_1452,N_1374,N_1366);
nor U1453 (N_1453,N_1354,N_1323);
or U1454 (N_1454,N_1320,N_1312);
xor U1455 (N_1455,N_1343,N_1306);
xor U1456 (N_1456,N_1396,N_1303);
xnor U1457 (N_1457,N_1305,N_1392);
xor U1458 (N_1458,N_1367,N_1397);
nor U1459 (N_1459,N_1350,N_1347);
xnor U1460 (N_1460,N_1393,N_1338);
nor U1461 (N_1461,N_1381,N_1342);
nand U1462 (N_1462,N_1329,N_1378);
nand U1463 (N_1463,N_1348,N_1366);
or U1464 (N_1464,N_1330,N_1305);
xor U1465 (N_1465,N_1325,N_1348);
or U1466 (N_1466,N_1316,N_1351);
or U1467 (N_1467,N_1363,N_1333);
nor U1468 (N_1468,N_1334,N_1324);
or U1469 (N_1469,N_1308,N_1386);
or U1470 (N_1470,N_1359,N_1317);
nor U1471 (N_1471,N_1389,N_1366);
xnor U1472 (N_1472,N_1335,N_1321);
and U1473 (N_1473,N_1301,N_1308);
or U1474 (N_1474,N_1335,N_1388);
nand U1475 (N_1475,N_1398,N_1387);
or U1476 (N_1476,N_1389,N_1391);
nand U1477 (N_1477,N_1367,N_1304);
xor U1478 (N_1478,N_1356,N_1350);
xnor U1479 (N_1479,N_1376,N_1398);
and U1480 (N_1480,N_1341,N_1310);
nand U1481 (N_1481,N_1352,N_1396);
xor U1482 (N_1482,N_1330,N_1374);
nand U1483 (N_1483,N_1389,N_1317);
or U1484 (N_1484,N_1349,N_1305);
nand U1485 (N_1485,N_1393,N_1369);
nand U1486 (N_1486,N_1342,N_1366);
xor U1487 (N_1487,N_1396,N_1350);
xor U1488 (N_1488,N_1322,N_1381);
and U1489 (N_1489,N_1378,N_1359);
or U1490 (N_1490,N_1337,N_1335);
nand U1491 (N_1491,N_1329,N_1347);
nand U1492 (N_1492,N_1398,N_1305);
xnor U1493 (N_1493,N_1349,N_1325);
or U1494 (N_1494,N_1317,N_1324);
xor U1495 (N_1495,N_1358,N_1373);
xor U1496 (N_1496,N_1329,N_1395);
nor U1497 (N_1497,N_1397,N_1331);
xor U1498 (N_1498,N_1352,N_1399);
and U1499 (N_1499,N_1394,N_1382);
xor U1500 (N_1500,N_1412,N_1495);
or U1501 (N_1501,N_1413,N_1457);
xor U1502 (N_1502,N_1449,N_1422);
nor U1503 (N_1503,N_1421,N_1453);
nand U1504 (N_1504,N_1487,N_1490);
xor U1505 (N_1505,N_1444,N_1423);
nand U1506 (N_1506,N_1472,N_1451);
or U1507 (N_1507,N_1499,N_1435);
or U1508 (N_1508,N_1401,N_1478);
or U1509 (N_1509,N_1493,N_1476);
and U1510 (N_1510,N_1479,N_1450);
nand U1511 (N_1511,N_1459,N_1481);
and U1512 (N_1512,N_1447,N_1410);
nand U1513 (N_1513,N_1416,N_1455);
xnor U1514 (N_1514,N_1466,N_1438);
nand U1515 (N_1515,N_1484,N_1477);
nand U1516 (N_1516,N_1441,N_1436);
nor U1517 (N_1517,N_1400,N_1419);
or U1518 (N_1518,N_1446,N_1492);
nor U1519 (N_1519,N_1431,N_1468);
or U1520 (N_1520,N_1483,N_1496);
or U1521 (N_1521,N_1461,N_1433);
or U1522 (N_1522,N_1420,N_1482);
xor U1523 (N_1523,N_1428,N_1475);
xor U1524 (N_1524,N_1440,N_1469);
or U1525 (N_1525,N_1488,N_1454);
and U1526 (N_1526,N_1424,N_1491);
nand U1527 (N_1527,N_1448,N_1427);
or U1528 (N_1528,N_1437,N_1439);
nand U1529 (N_1529,N_1458,N_1443);
xor U1530 (N_1530,N_1425,N_1467);
and U1531 (N_1531,N_1464,N_1471);
or U1532 (N_1532,N_1497,N_1411);
or U1533 (N_1533,N_1432,N_1473);
nor U1534 (N_1534,N_1445,N_1405);
nand U1535 (N_1535,N_1494,N_1426);
nor U1536 (N_1536,N_1460,N_1456);
and U1537 (N_1537,N_1409,N_1404);
nand U1538 (N_1538,N_1452,N_1498);
and U1539 (N_1539,N_1485,N_1402);
nand U1540 (N_1540,N_1462,N_1403);
nand U1541 (N_1541,N_1489,N_1430);
or U1542 (N_1542,N_1465,N_1474);
nand U1543 (N_1543,N_1408,N_1406);
and U1544 (N_1544,N_1470,N_1434);
or U1545 (N_1545,N_1463,N_1480);
and U1546 (N_1546,N_1442,N_1486);
and U1547 (N_1547,N_1407,N_1415);
nor U1548 (N_1548,N_1414,N_1429);
nand U1549 (N_1549,N_1417,N_1418);
nand U1550 (N_1550,N_1411,N_1419);
xnor U1551 (N_1551,N_1471,N_1492);
or U1552 (N_1552,N_1490,N_1450);
nand U1553 (N_1553,N_1403,N_1404);
or U1554 (N_1554,N_1412,N_1469);
xnor U1555 (N_1555,N_1492,N_1405);
xnor U1556 (N_1556,N_1487,N_1462);
nor U1557 (N_1557,N_1470,N_1432);
xor U1558 (N_1558,N_1438,N_1487);
and U1559 (N_1559,N_1491,N_1429);
or U1560 (N_1560,N_1434,N_1427);
nor U1561 (N_1561,N_1436,N_1477);
nand U1562 (N_1562,N_1484,N_1486);
or U1563 (N_1563,N_1475,N_1417);
xor U1564 (N_1564,N_1446,N_1404);
nand U1565 (N_1565,N_1487,N_1421);
nand U1566 (N_1566,N_1439,N_1495);
nand U1567 (N_1567,N_1407,N_1432);
and U1568 (N_1568,N_1446,N_1466);
xnor U1569 (N_1569,N_1455,N_1410);
nand U1570 (N_1570,N_1428,N_1450);
and U1571 (N_1571,N_1415,N_1461);
nor U1572 (N_1572,N_1422,N_1437);
xnor U1573 (N_1573,N_1409,N_1490);
or U1574 (N_1574,N_1454,N_1447);
nor U1575 (N_1575,N_1467,N_1423);
xnor U1576 (N_1576,N_1443,N_1446);
or U1577 (N_1577,N_1439,N_1456);
or U1578 (N_1578,N_1478,N_1459);
nor U1579 (N_1579,N_1435,N_1455);
and U1580 (N_1580,N_1489,N_1429);
nand U1581 (N_1581,N_1454,N_1420);
xnor U1582 (N_1582,N_1496,N_1473);
and U1583 (N_1583,N_1414,N_1483);
nand U1584 (N_1584,N_1455,N_1486);
xor U1585 (N_1585,N_1498,N_1455);
nor U1586 (N_1586,N_1484,N_1433);
or U1587 (N_1587,N_1406,N_1453);
or U1588 (N_1588,N_1447,N_1424);
xor U1589 (N_1589,N_1439,N_1485);
nand U1590 (N_1590,N_1486,N_1404);
xor U1591 (N_1591,N_1430,N_1465);
or U1592 (N_1592,N_1449,N_1494);
nor U1593 (N_1593,N_1494,N_1400);
or U1594 (N_1594,N_1496,N_1485);
nor U1595 (N_1595,N_1414,N_1442);
nor U1596 (N_1596,N_1422,N_1453);
and U1597 (N_1597,N_1430,N_1444);
and U1598 (N_1598,N_1403,N_1459);
xor U1599 (N_1599,N_1478,N_1432);
nand U1600 (N_1600,N_1500,N_1593);
nand U1601 (N_1601,N_1530,N_1557);
or U1602 (N_1602,N_1586,N_1572);
nor U1603 (N_1603,N_1529,N_1502);
xnor U1604 (N_1604,N_1516,N_1551);
nor U1605 (N_1605,N_1594,N_1576);
nand U1606 (N_1606,N_1562,N_1589);
nand U1607 (N_1607,N_1565,N_1536);
xor U1608 (N_1608,N_1584,N_1509);
and U1609 (N_1609,N_1553,N_1528);
or U1610 (N_1610,N_1579,N_1521);
nor U1611 (N_1611,N_1596,N_1559);
nand U1612 (N_1612,N_1585,N_1567);
nor U1613 (N_1613,N_1505,N_1545);
nand U1614 (N_1614,N_1501,N_1515);
nor U1615 (N_1615,N_1513,N_1549);
or U1616 (N_1616,N_1560,N_1543);
and U1617 (N_1617,N_1541,N_1510);
and U1618 (N_1618,N_1526,N_1566);
and U1619 (N_1619,N_1558,N_1522);
nand U1620 (N_1620,N_1574,N_1580);
nand U1621 (N_1621,N_1535,N_1544);
nor U1622 (N_1622,N_1547,N_1512);
xor U1623 (N_1623,N_1578,N_1518);
nand U1624 (N_1624,N_1592,N_1588);
xor U1625 (N_1625,N_1568,N_1590);
and U1626 (N_1626,N_1599,N_1561);
or U1627 (N_1627,N_1548,N_1507);
and U1628 (N_1628,N_1571,N_1597);
nor U1629 (N_1629,N_1514,N_1575);
nor U1630 (N_1630,N_1573,N_1524);
and U1631 (N_1631,N_1570,N_1581);
and U1632 (N_1632,N_1537,N_1546);
or U1633 (N_1633,N_1569,N_1503);
nand U1634 (N_1634,N_1583,N_1564);
or U1635 (N_1635,N_1539,N_1550);
or U1636 (N_1636,N_1540,N_1517);
and U1637 (N_1637,N_1533,N_1520);
and U1638 (N_1638,N_1506,N_1531);
and U1639 (N_1639,N_1582,N_1508);
or U1640 (N_1640,N_1587,N_1534);
nor U1641 (N_1641,N_1598,N_1595);
nand U1642 (N_1642,N_1563,N_1504);
nand U1643 (N_1643,N_1532,N_1555);
nand U1644 (N_1644,N_1591,N_1525);
nand U1645 (N_1645,N_1511,N_1523);
and U1646 (N_1646,N_1542,N_1519);
or U1647 (N_1647,N_1556,N_1527);
xnor U1648 (N_1648,N_1538,N_1554);
nor U1649 (N_1649,N_1552,N_1577);
nand U1650 (N_1650,N_1581,N_1539);
nand U1651 (N_1651,N_1551,N_1536);
nor U1652 (N_1652,N_1551,N_1556);
nand U1653 (N_1653,N_1596,N_1553);
and U1654 (N_1654,N_1526,N_1597);
and U1655 (N_1655,N_1547,N_1511);
nand U1656 (N_1656,N_1500,N_1514);
xor U1657 (N_1657,N_1540,N_1574);
and U1658 (N_1658,N_1546,N_1545);
nand U1659 (N_1659,N_1550,N_1532);
nor U1660 (N_1660,N_1509,N_1549);
xor U1661 (N_1661,N_1570,N_1508);
or U1662 (N_1662,N_1514,N_1597);
nor U1663 (N_1663,N_1504,N_1519);
or U1664 (N_1664,N_1561,N_1572);
or U1665 (N_1665,N_1563,N_1523);
xnor U1666 (N_1666,N_1570,N_1573);
nand U1667 (N_1667,N_1518,N_1561);
xor U1668 (N_1668,N_1578,N_1571);
and U1669 (N_1669,N_1599,N_1501);
nor U1670 (N_1670,N_1564,N_1592);
nor U1671 (N_1671,N_1500,N_1524);
and U1672 (N_1672,N_1527,N_1580);
and U1673 (N_1673,N_1543,N_1514);
xnor U1674 (N_1674,N_1547,N_1505);
nand U1675 (N_1675,N_1548,N_1503);
and U1676 (N_1676,N_1592,N_1590);
xor U1677 (N_1677,N_1576,N_1529);
or U1678 (N_1678,N_1569,N_1515);
or U1679 (N_1679,N_1559,N_1572);
and U1680 (N_1680,N_1573,N_1592);
and U1681 (N_1681,N_1560,N_1501);
or U1682 (N_1682,N_1519,N_1527);
nor U1683 (N_1683,N_1505,N_1500);
nand U1684 (N_1684,N_1554,N_1518);
nand U1685 (N_1685,N_1516,N_1565);
nor U1686 (N_1686,N_1512,N_1516);
nand U1687 (N_1687,N_1508,N_1513);
and U1688 (N_1688,N_1514,N_1593);
and U1689 (N_1689,N_1524,N_1577);
or U1690 (N_1690,N_1501,N_1586);
or U1691 (N_1691,N_1566,N_1588);
and U1692 (N_1692,N_1512,N_1567);
nor U1693 (N_1693,N_1569,N_1558);
nor U1694 (N_1694,N_1501,N_1539);
nand U1695 (N_1695,N_1597,N_1578);
nor U1696 (N_1696,N_1508,N_1568);
and U1697 (N_1697,N_1568,N_1515);
nand U1698 (N_1698,N_1570,N_1517);
xnor U1699 (N_1699,N_1528,N_1578);
and U1700 (N_1700,N_1619,N_1622);
nand U1701 (N_1701,N_1654,N_1610);
and U1702 (N_1702,N_1609,N_1682);
xnor U1703 (N_1703,N_1628,N_1644);
xor U1704 (N_1704,N_1631,N_1638);
or U1705 (N_1705,N_1647,N_1608);
xor U1706 (N_1706,N_1679,N_1681);
xor U1707 (N_1707,N_1666,N_1688);
xnor U1708 (N_1708,N_1613,N_1669);
xnor U1709 (N_1709,N_1648,N_1671);
nor U1710 (N_1710,N_1603,N_1637);
xor U1711 (N_1711,N_1615,N_1636);
and U1712 (N_1712,N_1658,N_1607);
or U1713 (N_1713,N_1686,N_1612);
nor U1714 (N_1714,N_1616,N_1640);
or U1715 (N_1715,N_1620,N_1651);
nand U1716 (N_1716,N_1618,N_1675);
nand U1717 (N_1717,N_1627,N_1602);
and U1718 (N_1718,N_1650,N_1659);
and U1719 (N_1719,N_1652,N_1625);
nand U1720 (N_1720,N_1655,N_1660);
and U1721 (N_1721,N_1614,N_1606);
xor U1722 (N_1722,N_1639,N_1698);
or U1723 (N_1723,N_1656,N_1653);
nor U1724 (N_1724,N_1633,N_1674);
nor U1725 (N_1725,N_1632,N_1667);
nor U1726 (N_1726,N_1626,N_1611);
xnor U1727 (N_1727,N_1617,N_1604);
or U1728 (N_1728,N_1663,N_1680);
xor U1729 (N_1729,N_1643,N_1642);
xor U1730 (N_1730,N_1694,N_1623);
nand U1731 (N_1731,N_1641,N_1629);
xor U1732 (N_1732,N_1621,N_1657);
nor U1733 (N_1733,N_1678,N_1600);
nor U1734 (N_1734,N_1691,N_1664);
xnor U1735 (N_1735,N_1699,N_1649);
nand U1736 (N_1736,N_1635,N_1605);
nand U1737 (N_1737,N_1670,N_1661);
xor U1738 (N_1738,N_1693,N_1646);
nor U1739 (N_1739,N_1687,N_1695);
nand U1740 (N_1740,N_1665,N_1673);
nor U1741 (N_1741,N_1634,N_1677);
nand U1742 (N_1742,N_1676,N_1692);
and U1743 (N_1743,N_1684,N_1672);
nor U1744 (N_1744,N_1689,N_1685);
nand U1745 (N_1745,N_1690,N_1624);
nand U1746 (N_1746,N_1696,N_1630);
xor U1747 (N_1747,N_1697,N_1662);
xnor U1748 (N_1748,N_1683,N_1601);
xor U1749 (N_1749,N_1645,N_1668);
xor U1750 (N_1750,N_1629,N_1655);
nor U1751 (N_1751,N_1625,N_1623);
nand U1752 (N_1752,N_1642,N_1639);
nor U1753 (N_1753,N_1651,N_1664);
xnor U1754 (N_1754,N_1611,N_1628);
nand U1755 (N_1755,N_1623,N_1624);
nor U1756 (N_1756,N_1652,N_1646);
and U1757 (N_1757,N_1695,N_1642);
xnor U1758 (N_1758,N_1692,N_1635);
nor U1759 (N_1759,N_1667,N_1699);
and U1760 (N_1760,N_1650,N_1643);
nand U1761 (N_1761,N_1617,N_1631);
or U1762 (N_1762,N_1665,N_1667);
or U1763 (N_1763,N_1616,N_1633);
xnor U1764 (N_1764,N_1691,N_1603);
or U1765 (N_1765,N_1693,N_1671);
xor U1766 (N_1766,N_1640,N_1635);
nand U1767 (N_1767,N_1699,N_1601);
and U1768 (N_1768,N_1615,N_1652);
nor U1769 (N_1769,N_1603,N_1607);
and U1770 (N_1770,N_1674,N_1621);
and U1771 (N_1771,N_1652,N_1626);
nand U1772 (N_1772,N_1695,N_1653);
xor U1773 (N_1773,N_1654,N_1630);
and U1774 (N_1774,N_1695,N_1663);
and U1775 (N_1775,N_1623,N_1660);
nor U1776 (N_1776,N_1655,N_1668);
and U1777 (N_1777,N_1628,N_1647);
or U1778 (N_1778,N_1682,N_1624);
nor U1779 (N_1779,N_1620,N_1630);
nand U1780 (N_1780,N_1648,N_1678);
nor U1781 (N_1781,N_1687,N_1605);
nand U1782 (N_1782,N_1644,N_1605);
or U1783 (N_1783,N_1605,N_1620);
nand U1784 (N_1784,N_1637,N_1664);
nor U1785 (N_1785,N_1605,N_1688);
nor U1786 (N_1786,N_1686,N_1624);
and U1787 (N_1787,N_1640,N_1634);
nand U1788 (N_1788,N_1630,N_1608);
xor U1789 (N_1789,N_1673,N_1659);
and U1790 (N_1790,N_1695,N_1640);
xor U1791 (N_1791,N_1653,N_1621);
nand U1792 (N_1792,N_1692,N_1685);
xor U1793 (N_1793,N_1686,N_1668);
nand U1794 (N_1794,N_1603,N_1682);
xnor U1795 (N_1795,N_1600,N_1652);
or U1796 (N_1796,N_1648,N_1699);
or U1797 (N_1797,N_1651,N_1606);
xnor U1798 (N_1798,N_1637,N_1696);
nor U1799 (N_1799,N_1668,N_1682);
xnor U1800 (N_1800,N_1733,N_1782);
nor U1801 (N_1801,N_1786,N_1788);
or U1802 (N_1802,N_1787,N_1735);
nand U1803 (N_1803,N_1719,N_1758);
nand U1804 (N_1804,N_1771,N_1752);
and U1805 (N_1805,N_1741,N_1784);
nor U1806 (N_1806,N_1764,N_1785);
nand U1807 (N_1807,N_1777,N_1701);
nand U1808 (N_1808,N_1770,N_1760);
and U1809 (N_1809,N_1772,N_1710);
or U1810 (N_1810,N_1713,N_1723);
and U1811 (N_1811,N_1793,N_1774);
nand U1812 (N_1812,N_1751,N_1778);
nor U1813 (N_1813,N_1729,N_1700);
nor U1814 (N_1814,N_1716,N_1766);
and U1815 (N_1815,N_1715,N_1757);
xor U1816 (N_1816,N_1756,N_1753);
and U1817 (N_1817,N_1794,N_1799);
nor U1818 (N_1818,N_1797,N_1755);
nor U1819 (N_1819,N_1724,N_1722);
xor U1820 (N_1820,N_1792,N_1769);
nand U1821 (N_1821,N_1725,N_1790);
and U1822 (N_1822,N_1732,N_1706);
nor U1823 (N_1823,N_1783,N_1718);
nand U1824 (N_1824,N_1773,N_1740);
nand U1825 (N_1825,N_1707,N_1759);
or U1826 (N_1826,N_1762,N_1711);
xnor U1827 (N_1827,N_1728,N_1795);
nor U1828 (N_1828,N_1763,N_1714);
xor U1829 (N_1829,N_1776,N_1743);
nor U1830 (N_1830,N_1798,N_1761);
and U1831 (N_1831,N_1791,N_1779);
nor U1832 (N_1832,N_1721,N_1730);
xnor U1833 (N_1833,N_1767,N_1739);
and U1834 (N_1834,N_1745,N_1748);
xor U1835 (N_1835,N_1775,N_1746);
nand U1836 (N_1836,N_1734,N_1720);
or U1837 (N_1837,N_1749,N_1709);
nor U1838 (N_1838,N_1731,N_1704);
nor U1839 (N_1839,N_1744,N_1727);
nand U1840 (N_1840,N_1702,N_1742);
nand U1841 (N_1841,N_1780,N_1747);
and U1842 (N_1842,N_1726,N_1712);
nor U1843 (N_1843,N_1796,N_1765);
nand U1844 (N_1844,N_1703,N_1738);
nand U1845 (N_1845,N_1717,N_1781);
and U1846 (N_1846,N_1754,N_1750);
nand U1847 (N_1847,N_1708,N_1705);
nand U1848 (N_1848,N_1768,N_1789);
nand U1849 (N_1849,N_1737,N_1736);
nand U1850 (N_1850,N_1756,N_1741);
and U1851 (N_1851,N_1752,N_1779);
and U1852 (N_1852,N_1758,N_1706);
nor U1853 (N_1853,N_1741,N_1746);
or U1854 (N_1854,N_1792,N_1738);
nor U1855 (N_1855,N_1774,N_1783);
and U1856 (N_1856,N_1709,N_1748);
xor U1857 (N_1857,N_1704,N_1707);
or U1858 (N_1858,N_1743,N_1748);
xnor U1859 (N_1859,N_1768,N_1729);
nand U1860 (N_1860,N_1720,N_1795);
xnor U1861 (N_1861,N_1737,N_1783);
and U1862 (N_1862,N_1719,N_1786);
xnor U1863 (N_1863,N_1720,N_1732);
xnor U1864 (N_1864,N_1763,N_1718);
nand U1865 (N_1865,N_1751,N_1745);
nand U1866 (N_1866,N_1744,N_1797);
and U1867 (N_1867,N_1752,N_1705);
or U1868 (N_1868,N_1786,N_1750);
and U1869 (N_1869,N_1778,N_1712);
or U1870 (N_1870,N_1728,N_1715);
nor U1871 (N_1871,N_1759,N_1789);
or U1872 (N_1872,N_1745,N_1736);
nand U1873 (N_1873,N_1702,N_1740);
nor U1874 (N_1874,N_1725,N_1722);
or U1875 (N_1875,N_1796,N_1716);
or U1876 (N_1876,N_1774,N_1794);
nor U1877 (N_1877,N_1749,N_1767);
xnor U1878 (N_1878,N_1772,N_1747);
or U1879 (N_1879,N_1786,N_1798);
nor U1880 (N_1880,N_1754,N_1701);
nand U1881 (N_1881,N_1753,N_1795);
or U1882 (N_1882,N_1714,N_1732);
nor U1883 (N_1883,N_1757,N_1777);
nor U1884 (N_1884,N_1731,N_1730);
nand U1885 (N_1885,N_1787,N_1729);
or U1886 (N_1886,N_1768,N_1749);
and U1887 (N_1887,N_1798,N_1726);
xnor U1888 (N_1888,N_1768,N_1765);
or U1889 (N_1889,N_1708,N_1717);
nand U1890 (N_1890,N_1713,N_1736);
xor U1891 (N_1891,N_1737,N_1755);
and U1892 (N_1892,N_1770,N_1780);
or U1893 (N_1893,N_1751,N_1785);
and U1894 (N_1894,N_1713,N_1756);
nor U1895 (N_1895,N_1792,N_1753);
or U1896 (N_1896,N_1793,N_1765);
and U1897 (N_1897,N_1765,N_1794);
or U1898 (N_1898,N_1707,N_1738);
xor U1899 (N_1899,N_1792,N_1798);
nand U1900 (N_1900,N_1880,N_1866);
or U1901 (N_1901,N_1845,N_1841);
or U1902 (N_1902,N_1897,N_1894);
and U1903 (N_1903,N_1870,N_1861);
nor U1904 (N_1904,N_1822,N_1832);
xor U1905 (N_1905,N_1884,N_1854);
nand U1906 (N_1906,N_1821,N_1848);
nand U1907 (N_1907,N_1833,N_1804);
nand U1908 (N_1908,N_1859,N_1840);
or U1909 (N_1909,N_1842,N_1802);
or U1910 (N_1910,N_1887,N_1851);
nor U1911 (N_1911,N_1839,N_1846);
and U1912 (N_1912,N_1850,N_1810);
and U1913 (N_1913,N_1883,N_1844);
or U1914 (N_1914,N_1814,N_1811);
nand U1915 (N_1915,N_1827,N_1834);
nand U1916 (N_1916,N_1888,N_1873);
nand U1917 (N_1917,N_1820,N_1815);
nand U1918 (N_1918,N_1891,N_1806);
and U1919 (N_1919,N_1863,N_1869);
or U1920 (N_1920,N_1860,N_1823);
nand U1921 (N_1921,N_1886,N_1862);
or U1922 (N_1922,N_1895,N_1843);
nand U1923 (N_1923,N_1865,N_1836);
nand U1924 (N_1924,N_1801,N_1856);
xnor U1925 (N_1925,N_1831,N_1812);
nor U1926 (N_1926,N_1878,N_1808);
or U1927 (N_1927,N_1825,N_1818);
nor U1928 (N_1928,N_1881,N_1809);
and U1929 (N_1929,N_1871,N_1858);
or U1930 (N_1930,N_1857,N_1893);
or U1931 (N_1931,N_1807,N_1849);
xnor U1932 (N_1932,N_1877,N_1838);
or U1933 (N_1933,N_1898,N_1835);
nor U1934 (N_1934,N_1816,N_1867);
nor U1935 (N_1935,N_1868,N_1803);
and U1936 (N_1936,N_1847,N_1837);
or U1937 (N_1937,N_1899,N_1896);
and U1938 (N_1938,N_1879,N_1890);
nor U1939 (N_1939,N_1852,N_1875);
and U1940 (N_1940,N_1826,N_1819);
xor U1941 (N_1941,N_1892,N_1872);
nand U1942 (N_1942,N_1824,N_1876);
and U1943 (N_1943,N_1829,N_1817);
or U1944 (N_1944,N_1882,N_1853);
or U1945 (N_1945,N_1813,N_1864);
nand U1946 (N_1946,N_1855,N_1805);
xnor U1947 (N_1947,N_1874,N_1885);
and U1948 (N_1948,N_1830,N_1889);
nand U1949 (N_1949,N_1800,N_1828);
nand U1950 (N_1950,N_1862,N_1868);
and U1951 (N_1951,N_1850,N_1883);
nand U1952 (N_1952,N_1890,N_1801);
nand U1953 (N_1953,N_1889,N_1814);
xor U1954 (N_1954,N_1857,N_1854);
and U1955 (N_1955,N_1872,N_1833);
and U1956 (N_1956,N_1830,N_1805);
and U1957 (N_1957,N_1838,N_1841);
xnor U1958 (N_1958,N_1862,N_1872);
xor U1959 (N_1959,N_1871,N_1855);
xnor U1960 (N_1960,N_1828,N_1814);
and U1961 (N_1961,N_1831,N_1832);
nand U1962 (N_1962,N_1800,N_1853);
or U1963 (N_1963,N_1827,N_1889);
and U1964 (N_1964,N_1883,N_1878);
or U1965 (N_1965,N_1865,N_1818);
nor U1966 (N_1966,N_1847,N_1809);
or U1967 (N_1967,N_1883,N_1826);
nand U1968 (N_1968,N_1801,N_1811);
and U1969 (N_1969,N_1848,N_1849);
and U1970 (N_1970,N_1803,N_1838);
or U1971 (N_1971,N_1897,N_1810);
xor U1972 (N_1972,N_1875,N_1857);
or U1973 (N_1973,N_1855,N_1856);
or U1974 (N_1974,N_1855,N_1866);
nor U1975 (N_1975,N_1852,N_1820);
xnor U1976 (N_1976,N_1865,N_1854);
or U1977 (N_1977,N_1810,N_1820);
and U1978 (N_1978,N_1802,N_1877);
or U1979 (N_1979,N_1832,N_1846);
nand U1980 (N_1980,N_1845,N_1874);
nor U1981 (N_1981,N_1854,N_1833);
and U1982 (N_1982,N_1808,N_1803);
or U1983 (N_1983,N_1863,N_1848);
and U1984 (N_1984,N_1866,N_1838);
nand U1985 (N_1985,N_1829,N_1890);
and U1986 (N_1986,N_1814,N_1855);
xor U1987 (N_1987,N_1894,N_1848);
xnor U1988 (N_1988,N_1877,N_1817);
xnor U1989 (N_1989,N_1884,N_1822);
or U1990 (N_1990,N_1845,N_1810);
xor U1991 (N_1991,N_1821,N_1809);
nor U1992 (N_1992,N_1825,N_1848);
nor U1993 (N_1993,N_1856,N_1899);
or U1994 (N_1994,N_1886,N_1816);
nand U1995 (N_1995,N_1830,N_1893);
nand U1996 (N_1996,N_1854,N_1826);
xnor U1997 (N_1997,N_1859,N_1838);
xor U1998 (N_1998,N_1843,N_1845);
xor U1999 (N_1999,N_1838,N_1893);
or U2000 (N_2000,N_1908,N_1909);
xnor U2001 (N_2001,N_1974,N_1956);
nor U2002 (N_2002,N_1971,N_1972);
or U2003 (N_2003,N_1912,N_1989);
nor U2004 (N_2004,N_1977,N_1910);
or U2005 (N_2005,N_1959,N_1934);
nor U2006 (N_2006,N_1995,N_1979);
nand U2007 (N_2007,N_1903,N_1946);
nand U2008 (N_2008,N_1975,N_1928);
and U2009 (N_2009,N_1930,N_1943);
and U2010 (N_2010,N_1944,N_1968);
nand U2011 (N_2011,N_1963,N_1998);
and U2012 (N_2012,N_1911,N_1970);
or U2013 (N_2013,N_1905,N_1980);
and U2014 (N_2014,N_1904,N_1957);
nor U2015 (N_2015,N_1951,N_1921);
and U2016 (N_2016,N_1954,N_1940);
nor U2017 (N_2017,N_1913,N_1932);
nand U2018 (N_2018,N_1960,N_1918);
nand U2019 (N_2019,N_1981,N_1991);
xnor U2020 (N_2020,N_1955,N_1952);
nor U2021 (N_2021,N_1987,N_1994);
nand U2022 (N_2022,N_1966,N_1922);
nor U2023 (N_2023,N_1917,N_1942);
nor U2024 (N_2024,N_1950,N_1993);
and U2025 (N_2025,N_1906,N_1953);
nor U2026 (N_2026,N_1958,N_1997);
nor U2027 (N_2027,N_1933,N_1964);
nand U2028 (N_2028,N_1916,N_1969);
or U2029 (N_2029,N_1945,N_1907);
or U2030 (N_2030,N_1948,N_1947);
or U2031 (N_2031,N_1962,N_1927);
or U2032 (N_2032,N_1965,N_1914);
nand U2033 (N_2033,N_1935,N_1926);
nor U2034 (N_2034,N_1902,N_1982);
nand U2035 (N_2035,N_1924,N_1985);
nand U2036 (N_2036,N_1938,N_1973);
or U2037 (N_2037,N_1984,N_1967);
xor U2038 (N_2038,N_1978,N_1936);
or U2039 (N_2039,N_1999,N_1990);
nand U2040 (N_2040,N_1992,N_1976);
nor U2041 (N_2041,N_1988,N_1939);
xnor U2042 (N_2042,N_1931,N_1920);
nand U2043 (N_2043,N_1919,N_1996);
nand U2044 (N_2044,N_1986,N_1949);
and U2045 (N_2045,N_1941,N_1925);
nor U2046 (N_2046,N_1937,N_1900);
nand U2047 (N_2047,N_1983,N_1923);
nand U2048 (N_2048,N_1961,N_1901);
and U2049 (N_2049,N_1915,N_1929);
nor U2050 (N_2050,N_1951,N_1985);
nand U2051 (N_2051,N_1942,N_1978);
nor U2052 (N_2052,N_1965,N_1939);
and U2053 (N_2053,N_1924,N_1926);
nand U2054 (N_2054,N_1960,N_1981);
xnor U2055 (N_2055,N_1959,N_1920);
xor U2056 (N_2056,N_1983,N_1949);
nand U2057 (N_2057,N_1981,N_1994);
nand U2058 (N_2058,N_1970,N_1992);
or U2059 (N_2059,N_1980,N_1948);
nor U2060 (N_2060,N_1955,N_1949);
or U2061 (N_2061,N_1990,N_1998);
nor U2062 (N_2062,N_1990,N_1908);
nor U2063 (N_2063,N_1900,N_1963);
or U2064 (N_2064,N_1928,N_1981);
nand U2065 (N_2065,N_1974,N_1910);
nor U2066 (N_2066,N_1927,N_1988);
xnor U2067 (N_2067,N_1990,N_1915);
and U2068 (N_2068,N_1955,N_1956);
xor U2069 (N_2069,N_1907,N_1991);
nor U2070 (N_2070,N_1958,N_1974);
and U2071 (N_2071,N_1911,N_1979);
xnor U2072 (N_2072,N_1914,N_1944);
or U2073 (N_2073,N_1960,N_1939);
nor U2074 (N_2074,N_1982,N_1961);
nand U2075 (N_2075,N_1915,N_1918);
nor U2076 (N_2076,N_1977,N_1917);
or U2077 (N_2077,N_1925,N_1900);
xor U2078 (N_2078,N_1907,N_1967);
xor U2079 (N_2079,N_1969,N_1999);
nor U2080 (N_2080,N_1986,N_1932);
or U2081 (N_2081,N_1973,N_1989);
and U2082 (N_2082,N_1996,N_1954);
nor U2083 (N_2083,N_1970,N_1967);
xnor U2084 (N_2084,N_1958,N_1906);
or U2085 (N_2085,N_1907,N_1994);
or U2086 (N_2086,N_1999,N_1913);
and U2087 (N_2087,N_1915,N_1983);
or U2088 (N_2088,N_1983,N_1963);
xor U2089 (N_2089,N_1924,N_1950);
xor U2090 (N_2090,N_1946,N_1962);
xor U2091 (N_2091,N_1973,N_1920);
nand U2092 (N_2092,N_1926,N_1925);
and U2093 (N_2093,N_1934,N_1923);
nand U2094 (N_2094,N_1930,N_1945);
nor U2095 (N_2095,N_1936,N_1915);
nand U2096 (N_2096,N_1976,N_1930);
or U2097 (N_2097,N_1954,N_1907);
nor U2098 (N_2098,N_1928,N_1965);
nand U2099 (N_2099,N_1963,N_1989);
and U2100 (N_2100,N_2010,N_2055);
or U2101 (N_2101,N_2093,N_2057);
nor U2102 (N_2102,N_2052,N_2086);
xor U2103 (N_2103,N_2061,N_2034);
and U2104 (N_2104,N_2036,N_2000);
or U2105 (N_2105,N_2085,N_2054);
or U2106 (N_2106,N_2026,N_2067);
nand U2107 (N_2107,N_2035,N_2043);
xnor U2108 (N_2108,N_2002,N_2009);
nor U2109 (N_2109,N_2063,N_2016);
nor U2110 (N_2110,N_2082,N_2006);
nor U2111 (N_2111,N_2097,N_2053);
or U2112 (N_2112,N_2089,N_2033);
or U2113 (N_2113,N_2094,N_2024);
nor U2114 (N_2114,N_2059,N_2015);
nand U2115 (N_2115,N_2066,N_2008);
nand U2116 (N_2116,N_2073,N_2001);
nor U2117 (N_2117,N_2072,N_2076);
nor U2118 (N_2118,N_2004,N_2079);
xor U2119 (N_2119,N_2062,N_2037);
nand U2120 (N_2120,N_2083,N_2003);
nor U2121 (N_2121,N_2013,N_2018);
and U2122 (N_2122,N_2092,N_2040);
or U2123 (N_2123,N_2050,N_2080);
xor U2124 (N_2124,N_2058,N_2095);
xor U2125 (N_2125,N_2084,N_2005);
and U2126 (N_2126,N_2099,N_2088);
nor U2127 (N_2127,N_2014,N_2064);
nor U2128 (N_2128,N_2046,N_2032);
nor U2129 (N_2129,N_2007,N_2074);
xor U2130 (N_2130,N_2012,N_2039);
or U2131 (N_2131,N_2056,N_2098);
nand U2132 (N_2132,N_2077,N_2027);
nor U2133 (N_2133,N_2069,N_2044);
xor U2134 (N_2134,N_2087,N_2045);
and U2135 (N_2135,N_2030,N_2081);
or U2136 (N_2136,N_2021,N_2051);
xnor U2137 (N_2137,N_2022,N_2020);
or U2138 (N_2138,N_2031,N_2017);
nand U2139 (N_2139,N_2038,N_2070);
or U2140 (N_2140,N_2041,N_2090);
nand U2141 (N_2141,N_2065,N_2049);
and U2142 (N_2142,N_2068,N_2071);
xor U2143 (N_2143,N_2028,N_2075);
or U2144 (N_2144,N_2091,N_2096);
and U2145 (N_2145,N_2060,N_2025);
xor U2146 (N_2146,N_2019,N_2042);
and U2147 (N_2147,N_2048,N_2078);
or U2148 (N_2148,N_2047,N_2029);
nor U2149 (N_2149,N_2011,N_2023);
or U2150 (N_2150,N_2050,N_2079);
xnor U2151 (N_2151,N_2023,N_2060);
nor U2152 (N_2152,N_2023,N_2058);
and U2153 (N_2153,N_2063,N_2061);
or U2154 (N_2154,N_2071,N_2040);
and U2155 (N_2155,N_2059,N_2027);
or U2156 (N_2156,N_2060,N_2066);
and U2157 (N_2157,N_2069,N_2065);
nor U2158 (N_2158,N_2032,N_2040);
xor U2159 (N_2159,N_2048,N_2021);
or U2160 (N_2160,N_2014,N_2045);
or U2161 (N_2161,N_2097,N_2036);
xnor U2162 (N_2162,N_2021,N_2047);
xor U2163 (N_2163,N_2008,N_2081);
xnor U2164 (N_2164,N_2066,N_2042);
and U2165 (N_2165,N_2033,N_2025);
or U2166 (N_2166,N_2000,N_2040);
nor U2167 (N_2167,N_2044,N_2043);
xnor U2168 (N_2168,N_2065,N_2040);
or U2169 (N_2169,N_2046,N_2041);
or U2170 (N_2170,N_2033,N_2021);
or U2171 (N_2171,N_2016,N_2074);
and U2172 (N_2172,N_2048,N_2014);
nor U2173 (N_2173,N_2000,N_2016);
or U2174 (N_2174,N_2050,N_2090);
nand U2175 (N_2175,N_2033,N_2018);
and U2176 (N_2176,N_2089,N_2080);
nand U2177 (N_2177,N_2020,N_2090);
or U2178 (N_2178,N_2075,N_2023);
or U2179 (N_2179,N_2062,N_2018);
and U2180 (N_2180,N_2005,N_2089);
or U2181 (N_2181,N_2059,N_2021);
or U2182 (N_2182,N_2034,N_2044);
and U2183 (N_2183,N_2047,N_2003);
and U2184 (N_2184,N_2084,N_2038);
or U2185 (N_2185,N_2009,N_2003);
nor U2186 (N_2186,N_2045,N_2039);
nand U2187 (N_2187,N_2020,N_2066);
nor U2188 (N_2188,N_2069,N_2058);
xnor U2189 (N_2189,N_2093,N_2037);
and U2190 (N_2190,N_2086,N_2061);
nor U2191 (N_2191,N_2090,N_2096);
and U2192 (N_2192,N_2061,N_2040);
and U2193 (N_2193,N_2083,N_2035);
nand U2194 (N_2194,N_2044,N_2054);
and U2195 (N_2195,N_2048,N_2074);
xor U2196 (N_2196,N_2084,N_2013);
nor U2197 (N_2197,N_2027,N_2003);
nand U2198 (N_2198,N_2090,N_2085);
nor U2199 (N_2199,N_2016,N_2061);
nor U2200 (N_2200,N_2169,N_2147);
and U2201 (N_2201,N_2192,N_2110);
or U2202 (N_2202,N_2149,N_2160);
nand U2203 (N_2203,N_2198,N_2115);
nand U2204 (N_2204,N_2148,N_2165);
or U2205 (N_2205,N_2154,N_2162);
and U2206 (N_2206,N_2190,N_2177);
xor U2207 (N_2207,N_2111,N_2157);
nand U2208 (N_2208,N_2193,N_2129);
xor U2209 (N_2209,N_2100,N_2144);
and U2210 (N_2210,N_2143,N_2194);
xnor U2211 (N_2211,N_2121,N_2142);
and U2212 (N_2212,N_2191,N_2120);
xor U2213 (N_2213,N_2178,N_2127);
xor U2214 (N_2214,N_2101,N_2186);
xnor U2215 (N_2215,N_2156,N_2153);
nor U2216 (N_2216,N_2114,N_2113);
and U2217 (N_2217,N_2109,N_2103);
nand U2218 (N_2218,N_2173,N_2105);
or U2219 (N_2219,N_2197,N_2189);
or U2220 (N_2220,N_2180,N_2168);
nand U2221 (N_2221,N_2184,N_2104);
nand U2222 (N_2222,N_2199,N_2146);
and U2223 (N_2223,N_2125,N_2135);
and U2224 (N_2224,N_2133,N_2108);
xor U2225 (N_2225,N_2136,N_2122);
nor U2226 (N_2226,N_2106,N_2195);
nor U2227 (N_2227,N_2107,N_2158);
xnor U2228 (N_2228,N_2155,N_2130);
nand U2229 (N_2229,N_2161,N_2188);
nor U2230 (N_2230,N_2112,N_2164);
nor U2231 (N_2231,N_2172,N_2138);
xnor U2232 (N_2232,N_2196,N_2159);
and U2233 (N_2233,N_2119,N_2117);
nand U2234 (N_2234,N_2102,N_2131);
and U2235 (N_2235,N_2124,N_2183);
nor U2236 (N_2236,N_2150,N_2166);
and U2237 (N_2237,N_2181,N_2179);
xor U2238 (N_2238,N_2176,N_2185);
and U2239 (N_2239,N_2171,N_2137);
nand U2240 (N_2240,N_2174,N_2141);
or U2241 (N_2241,N_2132,N_2175);
nand U2242 (N_2242,N_2118,N_2167);
and U2243 (N_2243,N_2123,N_2140);
xor U2244 (N_2244,N_2116,N_2170);
xor U2245 (N_2245,N_2151,N_2126);
or U2246 (N_2246,N_2152,N_2182);
xnor U2247 (N_2247,N_2145,N_2134);
nand U2248 (N_2248,N_2187,N_2163);
xor U2249 (N_2249,N_2128,N_2139);
and U2250 (N_2250,N_2175,N_2107);
nand U2251 (N_2251,N_2197,N_2161);
nor U2252 (N_2252,N_2183,N_2161);
and U2253 (N_2253,N_2178,N_2108);
nand U2254 (N_2254,N_2147,N_2179);
nor U2255 (N_2255,N_2126,N_2161);
nor U2256 (N_2256,N_2188,N_2138);
xnor U2257 (N_2257,N_2185,N_2114);
and U2258 (N_2258,N_2191,N_2125);
and U2259 (N_2259,N_2130,N_2198);
nand U2260 (N_2260,N_2196,N_2121);
or U2261 (N_2261,N_2180,N_2116);
xnor U2262 (N_2262,N_2119,N_2149);
nor U2263 (N_2263,N_2165,N_2105);
nor U2264 (N_2264,N_2178,N_2190);
nor U2265 (N_2265,N_2143,N_2183);
and U2266 (N_2266,N_2197,N_2134);
nor U2267 (N_2267,N_2124,N_2163);
xnor U2268 (N_2268,N_2174,N_2173);
or U2269 (N_2269,N_2125,N_2190);
nor U2270 (N_2270,N_2171,N_2139);
or U2271 (N_2271,N_2166,N_2199);
and U2272 (N_2272,N_2149,N_2128);
nand U2273 (N_2273,N_2107,N_2160);
nand U2274 (N_2274,N_2129,N_2180);
nor U2275 (N_2275,N_2113,N_2137);
and U2276 (N_2276,N_2131,N_2180);
nand U2277 (N_2277,N_2115,N_2167);
and U2278 (N_2278,N_2140,N_2120);
xnor U2279 (N_2279,N_2138,N_2114);
nand U2280 (N_2280,N_2145,N_2131);
or U2281 (N_2281,N_2188,N_2105);
and U2282 (N_2282,N_2196,N_2184);
and U2283 (N_2283,N_2167,N_2174);
nand U2284 (N_2284,N_2179,N_2156);
nand U2285 (N_2285,N_2143,N_2109);
nand U2286 (N_2286,N_2194,N_2166);
and U2287 (N_2287,N_2192,N_2138);
nand U2288 (N_2288,N_2129,N_2156);
nor U2289 (N_2289,N_2125,N_2104);
nor U2290 (N_2290,N_2122,N_2198);
or U2291 (N_2291,N_2135,N_2191);
xnor U2292 (N_2292,N_2136,N_2164);
nand U2293 (N_2293,N_2135,N_2161);
nor U2294 (N_2294,N_2142,N_2184);
and U2295 (N_2295,N_2180,N_2175);
or U2296 (N_2296,N_2190,N_2168);
nand U2297 (N_2297,N_2167,N_2124);
nor U2298 (N_2298,N_2175,N_2128);
or U2299 (N_2299,N_2173,N_2168);
nand U2300 (N_2300,N_2223,N_2281);
or U2301 (N_2301,N_2221,N_2225);
and U2302 (N_2302,N_2267,N_2282);
and U2303 (N_2303,N_2211,N_2251);
nand U2304 (N_2304,N_2250,N_2274);
nand U2305 (N_2305,N_2212,N_2208);
and U2306 (N_2306,N_2240,N_2292);
nor U2307 (N_2307,N_2255,N_2224);
nand U2308 (N_2308,N_2286,N_2265);
nor U2309 (N_2309,N_2295,N_2226);
xor U2310 (N_2310,N_2218,N_2247);
and U2311 (N_2311,N_2273,N_2233);
or U2312 (N_2312,N_2278,N_2257);
xor U2313 (N_2313,N_2220,N_2217);
or U2314 (N_2314,N_2239,N_2289);
or U2315 (N_2315,N_2203,N_2230);
or U2316 (N_2316,N_2280,N_2213);
or U2317 (N_2317,N_2238,N_2231);
xor U2318 (N_2318,N_2277,N_2261);
xor U2319 (N_2319,N_2236,N_2200);
nor U2320 (N_2320,N_2241,N_2264);
and U2321 (N_2321,N_2294,N_2210);
xnor U2322 (N_2322,N_2254,N_2287);
or U2323 (N_2323,N_2263,N_2272);
nand U2324 (N_2324,N_2204,N_2216);
or U2325 (N_2325,N_2243,N_2252);
nor U2326 (N_2326,N_2249,N_2209);
and U2327 (N_2327,N_2290,N_2288);
and U2328 (N_2328,N_2279,N_2299);
nand U2329 (N_2329,N_2283,N_2234);
or U2330 (N_2330,N_2262,N_2202);
and U2331 (N_2331,N_2206,N_2235);
and U2332 (N_2332,N_2296,N_2256);
or U2333 (N_2333,N_2270,N_2207);
or U2334 (N_2334,N_2229,N_2266);
or U2335 (N_2335,N_2275,N_2291);
xnor U2336 (N_2336,N_2260,N_2285);
xnor U2337 (N_2337,N_2237,N_2259);
and U2338 (N_2338,N_2214,N_2269);
nor U2339 (N_2339,N_2268,N_2228);
and U2340 (N_2340,N_2298,N_2242);
or U2341 (N_2341,N_2205,N_2246);
nand U2342 (N_2342,N_2258,N_2227);
and U2343 (N_2343,N_2232,N_2215);
or U2344 (N_2344,N_2271,N_2219);
nor U2345 (N_2345,N_2245,N_2201);
nor U2346 (N_2346,N_2244,N_2253);
nand U2347 (N_2347,N_2297,N_2293);
nand U2348 (N_2348,N_2284,N_2248);
or U2349 (N_2349,N_2276,N_2222);
xor U2350 (N_2350,N_2288,N_2201);
and U2351 (N_2351,N_2224,N_2287);
or U2352 (N_2352,N_2244,N_2296);
or U2353 (N_2353,N_2284,N_2291);
xor U2354 (N_2354,N_2286,N_2241);
nand U2355 (N_2355,N_2203,N_2211);
xnor U2356 (N_2356,N_2292,N_2277);
nor U2357 (N_2357,N_2242,N_2207);
xor U2358 (N_2358,N_2275,N_2221);
or U2359 (N_2359,N_2219,N_2265);
xor U2360 (N_2360,N_2267,N_2260);
and U2361 (N_2361,N_2241,N_2282);
nor U2362 (N_2362,N_2267,N_2240);
and U2363 (N_2363,N_2208,N_2288);
or U2364 (N_2364,N_2223,N_2263);
and U2365 (N_2365,N_2205,N_2294);
nor U2366 (N_2366,N_2204,N_2291);
xor U2367 (N_2367,N_2230,N_2298);
and U2368 (N_2368,N_2266,N_2295);
xor U2369 (N_2369,N_2200,N_2251);
or U2370 (N_2370,N_2281,N_2263);
and U2371 (N_2371,N_2267,N_2200);
xor U2372 (N_2372,N_2214,N_2290);
xnor U2373 (N_2373,N_2233,N_2264);
xnor U2374 (N_2374,N_2208,N_2295);
and U2375 (N_2375,N_2232,N_2254);
and U2376 (N_2376,N_2240,N_2207);
xor U2377 (N_2377,N_2214,N_2299);
or U2378 (N_2378,N_2229,N_2219);
and U2379 (N_2379,N_2297,N_2212);
nor U2380 (N_2380,N_2255,N_2285);
xor U2381 (N_2381,N_2223,N_2275);
nor U2382 (N_2382,N_2271,N_2255);
nor U2383 (N_2383,N_2236,N_2267);
and U2384 (N_2384,N_2254,N_2276);
or U2385 (N_2385,N_2220,N_2235);
or U2386 (N_2386,N_2206,N_2282);
or U2387 (N_2387,N_2227,N_2213);
and U2388 (N_2388,N_2287,N_2216);
xor U2389 (N_2389,N_2270,N_2208);
nor U2390 (N_2390,N_2298,N_2289);
nor U2391 (N_2391,N_2283,N_2244);
xor U2392 (N_2392,N_2213,N_2239);
nor U2393 (N_2393,N_2264,N_2203);
or U2394 (N_2394,N_2230,N_2244);
or U2395 (N_2395,N_2228,N_2223);
nor U2396 (N_2396,N_2285,N_2257);
or U2397 (N_2397,N_2235,N_2292);
nand U2398 (N_2398,N_2245,N_2251);
nand U2399 (N_2399,N_2238,N_2224);
xor U2400 (N_2400,N_2324,N_2352);
nor U2401 (N_2401,N_2312,N_2390);
and U2402 (N_2402,N_2389,N_2383);
xor U2403 (N_2403,N_2371,N_2356);
and U2404 (N_2404,N_2365,N_2349);
and U2405 (N_2405,N_2362,N_2376);
or U2406 (N_2406,N_2384,N_2310);
xor U2407 (N_2407,N_2363,N_2372);
xnor U2408 (N_2408,N_2344,N_2313);
xnor U2409 (N_2409,N_2330,N_2386);
nor U2410 (N_2410,N_2302,N_2333);
xor U2411 (N_2411,N_2327,N_2347);
and U2412 (N_2412,N_2311,N_2366);
nand U2413 (N_2413,N_2323,N_2331);
nand U2414 (N_2414,N_2326,N_2357);
or U2415 (N_2415,N_2343,N_2348);
or U2416 (N_2416,N_2317,N_2375);
nand U2417 (N_2417,N_2322,N_2301);
and U2418 (N_2418,N_2385,N_2318);
and U2419 (N_2419,N_2320,N_2307);
xnor U2420 (N_2420,N_2380,N_2339);
xor U2421 (N_2421,N_2304,N_2398);
and U2422 (N_2422,N_2300,N_2394);
and U2423 (N_2423,N_2373,N_2315);
or U2424 (N_2424,N_2345,N_2337);
nand U2425 (N_2425,N_2340,N_2350);
nand U2426 (N_2426,N_2370,N_2368);
and U2427 (N_2427,N_2391,N_2351);
or U2428 (N_2428,N_2364,N_2378);
nand U2429 (N_2429,N_2314,N_2338);
nor U2430 (N_2430,N_2377,N_2361);
xnor U2431 (N_2431,N_2325,N_2346);
nor U2432 (N_2432,N_2341,N_2342);
and U2433 (N_2433,N_2308,N_2382);
nand U2434 (N_2434,N_2360,N_2309);
or U2435 (N_2435,N_2396,N_2388);
nand U2436 (N_2436,N_2332,N_2306);
xnor U2437 (N_2437,N_2334,N_2393);
and U2438 (N_2438,N_2335,N_2316);
xnor U2439 (N_2439,N_2358,N_2397);
xnor U2440 (N_2440,N_2379,N_2305);
xor U2441 (N_2441,N_2321,N_2336);
or U2442 (N_2442,N_2392,N_2395);
xor U2443 (N_2443,N_2354,N_2328);
and U2444 (N_2444,N_2355,N_2374);
nor U2445 (N_2445,N_2367,N_2399);
or U2446 (N_2446,N_2329,N_2369);
nand U2447 (N_2447,N_2381,N_2387);
or U2448 (N_2448,N_2319,N_2359);
nor U2449 (N_2449,N_2303,N_2353);
nor U2450 (N_2450,N_2369,N_2359);
xor U2451 (N_2451,N_2392,N_2378);
nand U2452 (N_2452,N_2394,N_2372);
or U2453 (N_2453,N_2310,N_2368);
nor U2454 (N_2454,N_2345,N_2342);
and U2455 (N_2455,N_2338,N_2310);
xnor U2456 (N_2456,N_2379,N_2328);
and U2457 (N_2457,N_2369,N_2375);
nand U2458 (N_2458,N_2328,N_2344);
xor U2459 (N_2459,N_2312,N_2385);
xor U2460 (N_2460,N_2309,N_2374);
xor U2461 (N_2461,N_2352,N_2317);
nor U2462 (N_2462,N_2369,N_2345);
and U2463 (N_2463,N_2343,N_2327);
nor U2464 (N_2464,N_2360,N_2333);
nand U2465 (N_2465,N_2310,N_2341);
nor U2466 (N_2466,N_2339,N_2343);
nand U2467 (N_2467,N_2311,N_2388);
xnor U2468 (N_2468,N_2385,N_2342);
xor U2469 (N_2469,N_2371,N_2346);
nor U2470 (N_2470,N_2301,N_2313);
nand U2471 (N_2471,N_2398,N_2362);
nor U2472 (N_2472,N_2371,N_2347);
xnor U2473 (N_2473,N_2392,N_2361);
nand U2474 (N_2474,N_2380,N_2388);
and U2475 (N_2475,N_2367,N_2351);
and U2476 (N_2476,N_2346,N_2389);
nor U2477 (N_2477,N_2302,N_2329);
or U2478 (N_2478,N_2320,N_2323);
or U2479 (N_2479,N_2311,N_2382);
and U2480 (N_2480,N_2386,N_2380);
xor U2481 (N_2481,N_2376,N_2377);
or U2482 (N_2482,N_2371,N_2343);
nand U2483 (N_2483,N_2328,N_2366);
nor U2484 (N_2484,N_2373,N_2355);
xnor U2485 (N_2485,N_2374,N_2326);
xnor U2486 (N_2486,N_2361,N_2309);
or U2487 (N_2487,N_2364,N_2310);
and U2488 (N_2488,N_2392,N_2349);
nand U2489 (N_2489,N_2350,N_2396);
and U2490 (N_2490,N_2375,N_2328);
xnor U2491 (N_2491,N_2341,N_2328);
xnor U2492 (N_2492,N_2398,N_2308);
and U2493 (N_2493,N_2341,N_2307);
nor U2494 (N_2494,N_2392,N_2356);
nand U2495 (N_2495,N_2315,N_2362);
and U2496 (N_2496,N_2302,N_2385);
nor U2497 (N_2497,N_2326,N_2385);
or U2498 (N_2498,N_2352,N_2366);
or U2499 (N_2499,N_2324,N_2388);
nor U2500 (N_2500,N_2477,N_2489);
nor U2501 (N_2501,N_2443,N_2458);
nor U2502 (N_2502,N_2474,N_2488);
nand U2503 (N_2503,N_2462,N_2422);
and U2504 (N_2504,N_2417,N_2494);
nand U2505 (N_2505,N_2436,N_2448);
and U2506 (N_2506,N_2492,N_2466);
and U2507 (N_2507,N_2419,N_2447);
or U2508 (N_2508,N_2421,N_2408);
or U2509 (N_2509,N_2442,N_2434);
xor U2510 (N_2510,N_2476,N_2499);
nor U2511 (N_2511,N_2433,N_2493);
nor U2512 (N_2512,N_2485,N_2467);
or U2513 (N_2513,N_2473,N_2491);
and U2514 (N_2514,N_2445,N_2478);
nor U2515 (N_2515,N_2452,N_2404);
xnor U2516 (N_2516,N_2457,N_2429);
and U2517 (N_2517,N_2427,N_2463);
nand U2518 (N_2518,N_2498,N_2409);
nand U2519 (N_2519,N_2479,N_2451);
nand U2520 (N_2520,N_2495,N_2414);
nand U2521 (N_2521,N_2413,N_2430);
nand U2522 (N_2522,N_2403,N_2483);
nand U2523 (N_2523,N_2464,N_2486);
or U2524 (N_2524,N_2438,N_2496);
nand U2525 (N_2525,N_2431,N_2446);
or U2526 (N_2526,N_2454,N_2456);
nor U2527 (N_2527,N_2415,N_2461);
or U2528 (N_2528,N_2455,N_2484);
nor U2529 (N_2529,N_2481,N_2420);
or U2530 (N_2530,N_2424,N_2471);
xnor U2531 (N_2531,N_2450,N_2407);
or U2532 (N_2532,N_2490,N_2410);
nand U2533 (N_2533,N_2425,N_2406);
and U2534 (N_2534,N_2402,N_2459);
xor U2535 (N_2535,N_2475,N_2469);
xnor U2536 (N_2536,N_2439,N_2487);
nor U2537 (N_2537,N_2412,N_2437);
and U2538 (N_2538,N_2441,N_2418);
nand U2539 (N_2539,N_2405,N_2428);
or U2540 (N_2540,N_2482,N_2411);
and U2541 (N_2541,N_2432,N_2423);
nor U2542 (N_2542,N_2435,N_2453);
and U2543 (N_2543,N_2449,N_2426);
nand U2544 (N_2544,N_2468,N_2401);
xnor U2545 (N_2545,N_2444,N_2416);
nor U2546 (N_2546,N_2497,N_2470);
and U2547 (N_2547,N_2472,N_2465);
nor U2548 (N_2548,N_2440,N_2480);
nand U2549 (N_2549,N_2400,N_2460);
nor U2550 (N_2550,N_2417,N_2460);
and U2551 (N_2551,N_2413,N_2409);
nand U2552 (N_2552,N_2440,N_2412);
nor U2553 (N_2553,N_2491,N_2426);
xor U2554 (N_2554,N_2498,N_2443);
xnor U2555 (N_2555,N_2473,N_2425);
and U2556 (N_2556,N_2493,N_2463);
or U2557 (N_2557,N_2440,N_2493);
nand U2558 (N_2558,N_2441,N_2471);
xor U2559 (N_2559,N_2440,N_2401);
xor U2560 (N_2560,N_2406,N_2471);
nor U2561 (N_2561,N_2419,N_2410);
xor U2562 (N_2562,N_2446,N_2495);
nand U2563 (N_2563,N_2464,N_2487);
and U2564 (N_2564,N_2438,N_2482);
xnor U2565 (N_2565,N_2430,N_2417);
xor U2566 (N_2566,N_2483,N_2491);
nor U2567 (N_2567,N_2403,N_2423);
or U2568 (N_2568,N_2424,N_2445);
nand U2569 (N_2569,N_2480,N_2412);
or U2570 (N_2570,N_2480,N_2493);
nor U2571 (N_2571,N_2492,N_2477);
nor U2572 (N_2572,N_2407,N_2478);
nor U2573 (N_2573,N_2478,N_2485);
and U2574 (N_2574,N_2426,N_2464);
nor U2575 (N_2575,N_2419,N_2404);
nand U2576 (N_2576,N_2473,N_2445);
or U2577 (N_2577,N_2455,N_2426);
nand U2578 (N_2578,N_2487,N_2406);
nor U2579 (N_2579,N_2402,N_2438);
or U2580 (N_2580,N_2412,N_2401);
or U2581 (N_2581,N_2407,N_2467);
nor U2582 (N_2582,N_2459,N_2496);
nor U2583 (N_2583,N_2449,N_2423);
xor U2584 (N_2584,N_2467,N_2419);
or U2585 (N_2585,N_2418,N_2475);
or U2586 (N_2586,N_2406,N_2481);
and U2587 (N_2587,N_2427,N_2462);
xnor U2588 (N_2588,N_2498,N_2446);
nor U2589 (N_2589,N_2479,N_2411);
and U2590 (N_2590,N_2493,N_2405);
nand U2591 (N_2591,N_2491,N_2443);
or U2592 (N_2592,N_2461,N_2452);
or U2593 (N_2593,N_2474,N_2455);
and U2594 (N_2594,N_2483,N_2450);
nor U2595 (N_2595,N_2473,N_2442);
xnor U2596 (N_2596,N_2485,N_2449);
xnor U2597 (N_2597,N_2455,N_2459);
or U2598 (N_2598,N_2419,N_2429);
xnor U2599 (N_2599,N_2465,N_2476);
nor U2600 (N_2600,N_2501,N_2597);
and U2601 (N_2601,N_2592,N_2546);
nand U2602 (N_2602,N_2509,N_2500);
nand U2603 (N_2603,N_2510,N_2532);
xor U2604 (N_2604,N_2514,N_2511);
xor U2605 (N_2605,N_2572,N_2587);
nor U2606 (N_2606,N_2521,N_2503);
xor U2607 (N_2607,N_2551,N_2549);
and U2608 (N_2608,N_2505,N_2547);
and U2609 (N_2609,N_2550,N_2512);
nand U2610 (N_2610,N_2595,N_2538);
nor U2611 (N_2611,N_2557,N_2504);
and U2612 (N_2612,N_2562,N_2519);
nor U2613 (N_2613,N_2515,N_2524);
xor U2614 (N_2614,N_2580,N_2541);
xor U2615 (N_2615,N_2506,N_2586);
and U2616 (N_2616,N_2566,N_2553);
and U2617 (N_2617,N_2579,N_2517);
xnor U2618 (N_2618,N_2507,N_2548);
nor U2619 (N_2619,N_2574,N_2529);
nor U2620 (N_2620,N_2528,N_2530);
xor U2621 (N_2621,N_2570,N_2596);
nor U2622 (N_2622,N_2584,N_2560);
and U2623 (N_2623,N_2577,N_2569);
or U2624 (N_2624,N_2535,N_2564);
nand U2625 (N_2625,N_2590,N_2578);
and U2626 (N_2626,N_2525,N_2527);
and U2627 (N_2627,N_2522,N_2576);
nor U2628 (N_2628,N_2599,N_2591);
nand U2629 (N_2629,N_2556,N_2526);
nor U2630 (N_2630,N_2581,N_2508);
and U2631 (N_2631,N_2555,N_2565);
xnor U2632 (N_2632,N_2537,N_2520);
or U2633 (N_2633,N_2568,N_2573);
xor U2634 (N_2634,N_2523,N_2539);
or U2635 (N_2635,N_2516,N_2513);
nor U2636 (N_2636,N_2575,N_2543);
or U2637 (N_2637,N_2542,N_2588);
and U2638 (N_2638,N_2502,N_2544);
nand U2639 (N_2639,N_2582,N_2563);
nand U2640 (N_2640,N_2554,N_2531);
or U2641 (N_2641,N_2559,N_2593);
nand U2642 (N_2642,N_2594,N_2518);
xor U2643 (N_2643,N_2552,N_2534);
xnor U2644 (N_2644,N_2583,N_2585);
and U2645 (N_2645,N_2598,N_2589);
or U2646 (N_2646,N_2571,N_2533);
xor U2647 (N_2647,N_2540,N_2545);
xnor U2648 (N_2648,N_2567,N_2558);
and U2649 (N_2649,N_2561,N_2536);
nand U2650 (N_2650,N_2591,N_2571);
xor U2651 (N_2651,N_2566,N_2560);
nor U2652 (N_2652,N_2544,N_2572);
or U2653 (N_2653,N_2535,N_2587);
and U2654 (N_2654,N_2519,N_2550);
nand U2655 (N_2655,N_2588,N_2543);
and U2656 (N_2656,N_2584,N_2513);
nor U2657 (N_2657,N_2520,N_2534);
nand U2658 (N_2658,N_2521,N_2581);
nand U2659 (N_2659,N_2535,N_2505);
and U2660 (N_2660,N_2539,N_2594);
xnor U2661 (N_2661,N_2554,N_2530);
xor U2662 (N_2662,N_2518,N_2570);
nand U2663 (N_2663,N_2563,N_2597);
or U2664 (N_2664,N_2504,N_2573);
nor U2665 (N_2665,N_2574,N_2570);
nor U2666 (N_2666,N_2550,N_2565);
nand U2667 (N_2667,N_2543,N_2525);
and U2668 (N_2668,N_2589,N_2513);
xnor U2669 (N_2669,N_2524,N_2533);
xor U2670 (N_2670,N_2593,N_2572);
or U2671 (N_2671,N_2519,N_2561);
or U2672 (N_2672,N_2534,N_2547);
or U2673 (N_2673,N_2526,N_2594);
xor U2674 (N_2674,N_2567,N_2584);
nand U2675 (N_2675,N_2559,N_2587);
nor U2676 (N_2676,N_2533,N_2563);
xor U2677 (N_2677,N_2566,N_2555);
nand U2678 (N_2678,N_2587,N_2534);
nand U2679 (N_2679,N_2593,N_2514);
nor U2680 (N_2680,N_2508,N_2549);
nand U2681 (N_2681,N_2505,N_2593);
or U2682 (N_2682,N_2595,N_2545);
or U2683 (N_2683,N_2574,N_2526);
and U2684 (N_2684,N_2513,N_2568);
nand U2685 (N_2685,N_2506,N_2511);
nand U2686 (N_2686,N_2517,N_2573);
and U2687 (N_2687,N_2590,N_2519);
or U2688 (N_2688,N_2530,N_2512);
nor U2689 (N_2689,N_2582,N_2502);
or U2690 (N_2690,N_2583,N_2579);
xnor U2691 (N_2691,N_2511,N_2585);
and U2692 (N_2692,N_2598,N_2534);
nor U2693 (N_2693,N_2567,N_2554);
nor U2694 (N_2694,N_2528,N_2577);
nor U2695 (N_2695,N_2599,N_2525);
nor U2696 (N_2696,N_2576,N_2588);
nor U2697 (N_2697,N_2594,N_2516);
or U2698 (N_2698,N_2553,N_2555);
or U2699 (N_2699,N_2540,N_2559);
nor U2700 (N_2700,N_2687,N_2686);
nand U2701 (N_2701,N_2645,N_2615);
nand U2702 (N_2702,N_2636,N_2673);
and U2703 (N_2703,N_2627,N_2678);
nor U2704 (N_2704,N_2658,N_2642);
or U2705 (N_2705,N_2633,N_2612);
or U2706 (N_2706,N_2648,N_2614);
xor U2707 (N_2707,N_2634,N_2693);
nor U2708 (N_2708,N_2692,N_2616);
nor U2709 (N_2709,N_2676,N_2689);
and U2710 (N_2710,N_2646,N_2618);
nor U2711 (N_2711,N_2684,N_2630);
xor U2712 (N_2712,N_2639,N_2606);
nand U2713 (N_2713,N_2660,N_2603);
and U2714 (N_2714,N_2655,N_2652);
or U2715 (N_2715,N_2649,N_2610);
and U2716 (N_2716,N_2657,N_2637);
nand U2717 (N_2717,N_2665,N_2674);
nand U2718 (N_2718,N_2619,N_2623);
xor U2719 (N_2719,N_2654,N_2608);
xor U2720 (N_2720,N_2690,N_2675);
or U2721 (N_2721,N_2659,N_2656);
nor U2722 (N_2722,N_2653,N_2666);
xor U2723 (N_2723,N_2669,N_2601);
nor U2724 (N_2724,N_2600,N_2647);
nor U2725 (N_2725,N_2605,N_2695);
and U2726 (N_2726,N_2651,N_2698);
and U2727 (N_2727,N_2685,N_2650);
or U2728 (N_2728,N_2688,N_2668);
xor U2729 (N_2729,N_2670,N_2671);
nand U2730 (N_2730,N_2638,N_2622);
nor U2731 (N_2731,N_2629,N_2680);
nor U2732 (N_2732,N_2683,N_2677);
or U2733 (N_2733,N_2664,N_2602);
and U2734 (N_2734,N_2661,N_2644);
xnor U2735 (N_2735,N_2699,N_2640);
nor U2736 (N_2736,N_2694,N_2641);
or U2737 (N_2737,N_2672,N_2624);
and U2738 (N_2738,N_2617,N_2682);
and U2739 (N_2739,N_2628,N_2626);
nand U2740 (N_2740,N_2679,N_2697);
and U2741 (N_2741,N_2667,N_2643);
and U2742 (N_2742,N_2691,N_2662);
or U2743 (N_2743,N_2620,N_2609);
xnor U2744 (N_2744,N_2607,N_2635);
and U2745 (N_2745,N_2696,N_2611);
xnor U2746 (N_2746,N_2663,N_2621);
and U2747 (N_2747,N_2604,N_2632);
nor U2748 (N_2748,N_2613,N_2631);
xnor U2749 (N_2749,N_2681,N_2625);
xnor U2750 (N_2750,N_2671,N_2660);
nor U2751 (N_2751,N_2682,N_2687);
or U2752 (N_2752,N_2669,N_2630);
and U2753 (N_2753,N_2615,N_2624);
nand U2754 (N_2754,N_2670,N_2605);
and U2755 (N_2755,N_2664,N_2631);
and U2756 (N_2756,N_2651,N_2677);
or U2757 (N_2757,N_2685,N_2629);
nor U2758 (N_2758,N_2682,N_2661);
nor U2759 (N_2759,N_2656,N_2626);
and U2760 (N_2760,N_2639,N_2698);
and U2761 (N_2761,N_2645,N_2646);
or U2762 (N_2762,N_2620,N_2655);
and U2763 (N_2763,N_2617,N_2696);
nand U2764 (N_2764,N_2626,N_2635);
or U2765 (N_2765,N_2637,N_2659);
nor U2766 (N_2766,N_2621,N_2683);
or U2767 (N_2767,N_2620,N_2645);
or U2768 (N_2768,N_2653,N_2692);
xnor U2769 (N_2769,N_2634,N_2635);
nand U2770 (N_2770,N_2625,N_2651);
nand U2771 (N_2771,N_2654,N_2609);
nor U2772 (N_2772,N_2676,N_2659);
or U2773 (N_2773,N_2635,N_2601);
xor U2774 (N_2774,N_2621,N_2666);
and U2775 (N_2775,N_2627,N_2692);
and U2776 (N_2776,N_2615,N_2674);
nand U2777 (N_2777,N_2673,N_2697);
and U2778 (N_2778,N_2622,N_2616);
and U2779 (N_2779,N_2653,N_2612);
or U2780 (N_2780,N_2601,N_2692);
nor U2781 (N_2781,N_2699,N_2609);
or U2782 (N_2782,N_2672,N_2699);
nor U2783 (N_2783,N_2621,N_2665);
and U2784 (N_2784,N_2622,N_2679);
or U2785 (N_2785,N_2670,N_2604);
or U2786 (N_2786,N_2601,N_2614);
nand U2787 (N_2787,N_2611,N_2652);
xnor U2788 (N_2788,N_2633,N_2624);
or U2789 (N_2789,N_2613,N_2660);
xor U2790 (N_2790,N_2615,N_2669);
or U2791 (N_2791,N_2659,N_2619);
nor U2792 (N_2792,N_2655,N_2696);
and U2793 (N_2793,N_2635,N_2602);
nor U2794 (N_2794,N_2617,N_2699);
and U2795 (N_2795,N_2683,N_2671);
xor U2796 (N_2796,N_2602,N_2639);
or U2797 (N_2797,N_2624,N_2623);
nor U2798 (N_2798,N_2605,N_2603);
or U2799 (N_2799,N_2668,N_2654);
or U2800 (N_2800,N_2749,N_2715);
or U2801 (N_2801,N_2796,N_2777);
or U2802 (N_2802,N_2723,N_2767);
nor U2803 (N_2803,N_2727,N_2719);
nor U2804 (N_2804,N_2790,N_2769);
xnor U2805 (N_2805,N_2720,N_2761);
xor U2806 (N_2806,N_2718,N_2739);
xnor U2807 (N_2807,N_2702,N_2730);
xnor U2808 (N_2808,N_2717,N_2766);
nor U2809 (N_2809,N_2707,N_2782);
nand U2810 (N_2810,N_2771,N_2774);
xor U2811 (N_2811,N_2797,N_2731);
and U2812 (N_2812,N_2736,N_2716);
or U2813 (N_2813,N_2746,N_2764);
and U2814 (N_2814,N_2747,N_2745);
and U2815 (N_2815,N_2780,N_2784);
and U2816 (N_2816,N_2708,N_2711);
xor U2817 (N_2817,N_2783,N_2795);
or U2818 (N_2818,N_2703,N_2733);
nand U2819 (N_2819,N_2781,N_2757);
nand U2820 (N_2820,N_2701,N_2778);
or U2821 (N_2821,N_2789,N_2776);
nor U2822 (N_2822,N_2721,N_2787);
or U2823 (N_2823,N_2775,N_2700);
and U2824 (N_2824,N_2725,N_2714);
xor U2825 (N_2825,N_2779,N_2704);
nand U2826 (N_2826,N_2758,N_2750);
and U2827 (N_2827,N_2737,N_2742);
or U2828 (N_2828,N_2786,N_2740);
or U2829 (N_2829,N_2751,N_2793);
and U2830 (N_2830,N_2755,N_2712);
nor U2831 (N_2831,N_2753,N_2744);
and U2832 (N_2832,N_2710,N_2738);
nor U2833 (N_2833,N_2728,N_2770);
or U2834 (N_2834,N_2754,N_2741);
xnor U2835 (N_2835,N_2799,N_2763);
or U2836 (N_2836,N_2773,N_2743);
xnor U2837 (N_2837,N_2735,N_2772);
and U2838 (N_2838,N_2768,N_2785);
nor U2839 (N_2839,N_2734,N_2794);
xor U2840 (N_2840,N_2726,N_2732);
nand U2841 (N_2841,N_2706,N_2709);
nand U2842 (N_2842,N_2729,N_2713);
xor U2843 (N_2843,N_2798,N_2748);
nand U2844 (N_2844,N_2792,N_2762);
xnor U2845 (N_2845,N_2791,N_2705);
and U2846 (N_2846,N_2756,N_2788);
xor U2847 (N_2847,N_2760,N_2722);
xnor U2848 (N_2848,N_2724,N_2765);
xnor U2849 (N_2849,N_2759,N_2752);
nand U2850 (N_2850,N_2767,N_2751);
and U2851 (N_2851,N_2748,N_2717);
or U2852 (N_2852,N_2756,N_2702);
and U2853 (N_2853,N_2762,N_2751);
xnor U2854 (N_2854,N_2787,N_2760);
or U2855 (N_2855,N_2752,N_2704);
nor U2856 (N_2856,N_2799,N_2720);
nor U2857 (N_2857,N_2738,N_2728);
and U2858 (N_2858,N_2749,N_2796);
or U2859 (N_2859,N_2752,N_2706);
or U2860 (N_2860,N_2765,N_2776);
xnor U2861 (N_2861,N_2799,N_2762);
xor U2862 (N_2862,N_2705,N_2746);
or U2863 (N_2863,N_2774,N_2770);
and U2864 (N_2864,N_2751,N_2768);
nand U2865 (N_2865,N_2708,N_2782);
nand U2866 (N_2866,N_2783,N_2746);
and U2867 (N_2867,N_2716,N_2759);
nand U2868 (N_2868,N_2793,N_2726);
nor U2869 (N_2869,N_2778,N_2724);
xor U2870 (N_2870,N_2728,N_2722);
and U2871 (N_2871,N_2779,N_2727);
and U2872 (N_2872,N_2755,N_2701);
and U2873 (N_2873,N_2774,N_2700);
nand U2874 (N_2874,N_2702,N_2719);
nor U2875 (N_2875,N_2737,N_2755);
xnor U2876 (N_2876,N_2786,N_2788);
or U2877 (N_2877,N_2706,N_2729);
xnor U2878 (N_2878,N_2740,N_2799);
xnor U2879 (N_2879,N_2739,N_2711);
nand U2880 (N_2880,N_2776,N_2745);
xnor U2881 (N_2881,N_2759,N_2753);
xnor U2882 (N_2882,N_2718,N_2714);
xnor U2883 (N_2883,N_2773,N_2709);
nor U2884 (N_2884,N_2702,N_2792);
or U2885 (N_2885,N_2724,N_2740);
nor U2886 (N_2886,N_2718,N_2793);
or U2887 (N_2887,N_2702,N_2758);
or U2888 (N_2888,N_2797,N_2728);
and U2889 (N_2889,N_2794,N_2770);
or U2890 (N_2890,N_2703,N_2764);
nor U2891 (N_2891,N_2762,N_2765);
xor U2892 (N_2892,N_2756,N_2729);
or U2893 (N_2893,N_2736,N_2734);
nor U2894 (N_2894,N_2745,N_2732);
nand U2895 (N_2895,N_2753,N_2763);
and U2896 (N_2896,N_2733,N_2797);
xnor U2897 (N_2897,N_2791,N_2750);
nand U2898 (N_2898,N_2761,N_2780);
and U2899 (N_2899,N_2766,N_2734);
or U2900 (N_2900,N_2893,N_2872);
or U2901 (N_2901,N_2810,N_2858);
xnor U2902 (N_2902,N_2874,N_2851);
and U2903 (N_2903,N_2830,N_2867);
nand U2904 (N_2904,N_2875,N_2876);
or U2905 (N_2905,N_2892,N_2806);
or U2906 (N_2906,N_2843,N_2871);
nand U2907 (N_2907,N_2852,N_2888);
nand U2908 (N_2908,N_2838,N_2805);
and U2909 (N_2909,N_2850,N_2824);
nor U2910 (N_2910,N_2821,N_2880);
nor U2911 (N_2911,N_2881,N_2866);
and U2912 (N_2912,N_2864,N_2800);
and U2913 (N_2913,N_2845,N_2822);
or U2914 (N_2914,N_2846,N_2829);
nor U2915 (N_2915,N_2889,N_2884);
nand U2916 (N_2916,N_2882,N_2807);
nand U2917 (N_2917,N_2826,N_2808);
xor U2918 (N_2918,N_2842,N_2883);
nand U2919 (N_2919,N_2878,N_2862);
nand U2920 (N_2920,N_2896,N_2801);
and U2921 (N_2921,N_2819,N_2802);
xnor U2922 (N_2922,N_2898,N_2855);
and U2923 (N_2923,N_2856,N_2811);
and U2924 (N_2924,N_2837,N_2818);
xnor U2925 (N_2925,N_2890,N_2877);
or U2926 (N_2926,N_2840,N_2836);
xnor U2927 (N_2927,N_2865,N_2869);
or U2928 (N_2928,N_2857,N_2834);
or U2929 (N_2929,N_2859,N_2854);
and U2930 (N_2930,N_2861,N_2817);
and U2931 (N_2931,N_2886,N_2897);
and U2932 (N_2932,N_2891,N_2820);
nand U2933 (N_2933,N_2879,N_2814);
or U2934 (N_2934,N_2849,N_2863);
xnor U2935 (N_2935,N_2870,N_2804);
nand U2936 (N_2936,N_2899,N_2832);
nor U2937 (N_2937,N_2868,N_2831);
xor U2938 (N_2938,N_2847,N_2823);
xor U2939 (N_2939,N_2825,N_2844);
or U2940 (N_2940,N_2815,N_2841);
nand U2941 (N_2941,N_2828,N_2827);
xor U2942 (N_2942,N_2833,N_2895);
nor U2943 (N_2943,N_2812,N_2803);
or U2944 (N_2944,N_2816,N_2839);
or U2945 (N_2945,N_2894,N_2887);
nand U2946 (N_2946,N_2873,N_2813);
or U2947 (N_2947,N_2848,N_2860);
xor U2948 (N_2948,N_2885,N_2835);
nor U2949 (N_2949,N_2809,N_2853);
xnor U2950 (N_2950,N_2865,N_2832);
nor U2951 (N_2951,N_2820,N_2827);
xnor U2952 (N_2952,N_2819,N_2817);
nand U2953 (N_2953,N_2893,N_2883);
nor U2954 (N_2954,N_2855,N_2896);
and U2955 (N_2955,N_2855,N_2819);
xor U2956 (N_2956,N_2833,N_2808);
or U2957 (N_2957,N_2887,N_2892);
and U2958 (N_2958,N_2860,N_2877);
or U2959 (N_2959,N_2877,N_2813);
and U2960 (N_2960,N_2894,N_2854);
nor U2961 (N_2961,N_2870,N_2826);
and U2962 (N_2962,N_2862,N_2812);
xnor U2963 (N_2963,N_2825,N_2822);
or U2964 (N_2964,N_2888,N_2886);
and U2965 (N_2965,N_2803,N_2809);
nand U2966 (N_2966,N_2835,N_2847);
xnor U2967 (N_2967,N_2826,N_2860);
or U2968 (N_2968,N_2861,N_2825);
and U2969 (N_2969,N_2871,N_2865);
nand U2970 (N_2970,N_2812,N_2877);
nand U2971 (N_2971,N_2838,N_2881);
or U2972 (N_2972,N_2862,N_2829);
nand U2973 (N_2973,N_2873,N_2830);
xnor U2974 (N_2974,N_2820,N_2821);
and U2975 (N_2975,N_2840,N_2808);
xnor U2976 (N_2976,N_2862,N_2891);
nand U2977 (N_2977,N_2813,N_2896);
nor U2978 (N_2978,N_2866,N_2854);
or U2979 (N_2979,N_2898,N_2831);
nand U2980 (N_2980,N_2846,N_2876);
nor U2981 (N_2981,N_2822,N_2833);
nand U2982 (N_2982,N_2815,N_2829);
xnor U2983 (N_2983,N_2825,N_2862);
nor U2984 (N_2984,N_2881,N_2839);
and U2985 (N_2985,N_2802,N_2801);
and U2986 (N_2986,N_2818,N_2813);
nor U2987 (N_2987,N_2831,N_2864);
nand U2988 (N_2988,N_2843,N_2891);
or U2989 (N_2989,N_2841,N_2804);
nand U2990 (N_2990,N_2874,N_2894);
nor U2991 (N_2991,N_2842,N_2819);
or U2992 (N_2992,N_2805,N_2814);
or U2993 (N_2993,N_2884,N_2851);
xor U2994 (N_2994,N_2839,N_2863);
or U2995 (N_2995,N_2813,N_2879);
or U2996 (N_2996,N_2879,N_2869);
nand U2997 (N_2997,N_2849,N_2888);
xnor U2998 (N_2998,N_2883,N_2806);
or U2999 (N_2999,N_2885,N_2819);
xor U3000 (N_3000,N_2986,N_2920);
and U3001 (N_3001,N_2996,N_2944);
nand U3002 (N_3002,N_2963,N_2968);
or U3003 (N_3003,N_2919,N_2993);
xor U3004 (N_3004,N_2943,N_2924);
and U3005 (N_3005,N_2902,N_2957);
or U3006 (N_3006,N_2997,N_2935);
and U3007 (N_3007,N_2907,N_2980);
xor U3008 (N_3008,N_2925,N_2921);
xor U3009 (N_3009,N_2969,N_2936);
or U3010 (N_3010,N_2926,N_2931);
and U3011 (N_3011,N_2950,N_2976);
or U3012 (N_3012,N_2956,N_2918);
nor U3013 (N_3013,N_2914,N_2961);
xnor U3014 (N_3014,N_2965,N_2942);
or U3015 (N_3015,N_2909,N_2930);
nand U3016 (N_3016,N_2971,N_2946);
and U3017 (N_3017,N_2962,N_2989);
and U3018 (N_3018,N_2967,N_2940);
xor U3019 (N_3019,N_2977,N_2912);
or U3020 (N_3020,N_2973,N_2917);
nand U3021 (N_3021,N_2945,N_2911);
xnor U3022 (N_3022,N_2928,N_2903);
nand U3023 (N_3023,N_2939,N_2974);
and U3024 (N_3024,N_2983,N_2913);
or U3025 (N_3025,N_2915,N_2922);
or U3026 (N_3026,N_2992,N_2985);
nand U3027 (N_3027,N_2933,N_2927);
nand U3028 (N_3028,N_2954,N_2908);
nand U3029 (N_3029,N_2966,N_2994);
nor U3030 (N_3030,N_2934,N_2995);
nand U3031 (N_3031,N_2972,N_2959);
xor U3032 (N_3032,N_2904,N_2988);
nor U3033 (N_3033,N_2929,N_2916);
or U3034 (N_3034,N_2970,N_2998);
xor U3035 (N_3035,N_2948,N_2990);
nand U3036 (N_3036,N_2941,N_2910);
or U3037 (N_3037,N_2978,N_2947);
nand U3038 (N_3038,N_2932,N_2999);
and U3039 (N_3039,N_2937,N_2900);
nor U3040 (N_3040,N_2982,N_2975);
nand U3041 (N_3041,N_2923,N_2991);
xor U3042 (N_3042,N_2951,N_2960);
nor U3043 (N_3043,N_2905,N_2906);
nand U3044 (N_3044,N_2984,N_2953);
and U3045 (N_3045,N_2952,N_2901);
and U3046 (N_3046,N_2949,N_2964);
nor U3047 (N_3047,N_2938,N_2955);
xnor U3048 (N_3048,N_2979,N_2958);
nand U3049 (N_3049,N_2981,N_2987);
nand U3050 (N_3050,N_2983,N_2904);
or U3051 (N_3051,N_2950,N_2919);
or U3052 (N_3052,N_2908,N_2986);
or U3053 (N_3053,N_2967,N_2961);
nand U3054 (N_3054,N_2940,N_2939);
nor U3055 (N_3055,N_2903,N_2972);
xnor U3056 (N_3056,N_2990,N_2902);
xnor U3057 (N_3057,N_2948,N_2999);
nor U3058 (N_3058,N_2936,N_2911);
xor U3059 (N_3059,N_2914,N_2956);
and U3060 (N_3060,N_2994,N_2976);
and U3061 (N_3061,N_2955,N_2932);
xor U3062 (N_3062,N_2956,N_2943);
nand U3063 (N_3063,N_2964,N_2924);
xnor U3064 (N_3064,N_2950,N_2927);
nor U3065 (N_3065,N_2967,N_2994);
and U3066 (N_3066,N_2950,N_2974);
xnor U3067 (N_3067,N_2931,N_2913);
or U3068 (N_3068,N_2900,N_2962);
nor U3069 (N_3069,N_2979,N_2961);
nor U3070 (N_3070,N_2939,N_2991);
or U3071 (N_3071,N_2996,N_2933);
and U3072 (N_3072,N_2913,N_2919);
nand U3073 (N_3073,N_2940,N_2980);
and U3074 (N_3074,N_2901,N_2973);
and U3075 (N_3075,N_2947,N_2998);
nand U3076 (N_3076,N_2968,N_2909);
nand U3077 (N_3077,N_2976,N_2986);
nand U3078 (N_3078,N_2988,N_2965);
or U3079 (N_3079,N_2934,N_2931);
and U3080 (N_3080,N_2965,N_2990);
and U3081 (N_3081,N_2923,N_2995);
nor U3082 (N_3082,N_2912,N_2969);
xnor U3083 (N_3083,N_2911,N_2972);
nand U3084 (N_3084,N_2964,N_2982);
and U3085 (N_3085,N_2970,N_2901);
or U3086 (N_3086,N_2917,N_2968);
xnor U3087 (N_3087,N_2985,N_2963);
nand U3088 (N_3088,N_2978,N_2993);
xnor U3089 (N_3089,N_2945,N_2976);
xor U3090 (N_3090,N_2947,N_2961);
or U3091 (N_3091,N_2906,N_2973);
or U3092 (N_3092,N_2977,N_2924);
nor U3093 (N_3093,N_2979,N_2987);
or U3094 (N_3094,N_2924,N_2995);
nand U3095 (N_3095,N_2940,N_2998);
nand U3096 (N_3096,N_2960,N_2915);
xor U3097 (N_3097,N_2961,N_2972);
nor U3098 (N_3098,N_2951,N_2914);
and U3099 (N_3099,N_2906,N_2986);
xor U3100 (N_3100,N_3076,N_3072);
and U3101 (N_3101,N_3031,N_3097);
and U3102 (N_3102,N_3091,N_3053);
nor U3103 (N_3103,N_3093,N_3090);
nand U3104 (N_3104,N_3078,N_3004);
nand U3105 (N_3105,N_3028,N_3060);
xor U3106 (N_3106,N_3026,N_3003);
nor U3107 (N_3107,N_3000,N_3018);
nand U3108 (N_3108,N_3039,N_3041);
or U3109 (N_3109,N_3092,N_3042);
or U3110 (N_3110,N_3069,N_3047);
nand U3111 (N_3111,N_3051,N_3019);
and U3112 (N_3112,N_3085,N_3055);
nand U3113 (N_3113,N_3066,N_3073);
nor U3114 (N_3114,N_3065,N_3050);
or U3115 (N_3115,N_3086,N_3035);
nand U3116 (N_3116,N_3037,N_3079);
and U3117 (N_3117,N_3045,N_3088);
or U3118 (N_3118,N_3022,N_3087);
or U3119 (N_3119,N_3056,N_3054);
or U3120 (N_3120,N_3011,N_3084);
nor U3121 (N_3121,N_3013,N_3009);
nor U3122 (N_3122,N_3030,N_3007);
xor U3123 (N_3123,N_3052,N_3001);
or U3124 (N_3124,N_3094,N_3067);
nand U3125 (N_3125,N_3099,N_3059);
and U3126 (N_3126,N_3048,N_3015);
nand U3127 (N_3127,N_3098,N_3071);
and U3128 (N_3128,N_3020,N_3025);
nor U3129 (N_3129,N_3032,N_3016);
xor U3130 (N_3130,N_3089,N_3081);
xor U3131 (N_3131,N_3005,N_3024);
nand U3132 (N_3132,N_3057,N_3083);
nand U3133 (N_3133,N_3068,N_3063);
xor U3134 (N_3134,N_3062,N_3043);
nor U3135 (N_3135,N_3074,N_3012);
and U3136 (N_3136,N_3070,N_3017);
or U3137 (N_3137,N_3095,N_3040);
nand U3138 (N_3138,N_3034,N_3027);
and U3139 (N_3139,N_3058,N_3002);
nor U3140 (N_3140,N_3029,N_3036);
xor U3141 (N_3141,N_3049,N_3075);
or U3142 (N_3142,N_3033,N_3014);
nor U3143 (N_3143,N_3023,N_3077);
xor U3144 (N_3144,N_3010,N_3082);
nor U3145 (N_3145,N_3061,N_3064);
nor U3146 (N_3146,N_3021,N_3006);
nand U3147 (N_3147,N_3080,N_3046);
nand U3148 (N_3148,N_3096,N_3038);
nor U3149 (N_3149,N_3044,N_3008);
nor U3150 (N_3150,N_3059,N_3097);
and U3151 (N_3151,N_3043,N_3090);
and U3152 (N_3152,N_3049,N_3021);
and U3153 (N_3153,N_3070,N_3022);
nor U3154 (N_3154,N_3036,N_3081);
nor U3155 (N_3155,N_3008,N_3055);
xor U3156 (N_3156,N_3004,N_3036);
nand U3157 (N_3157,N_3036,N_3089);
nor U3158 (N_3158,N_3061,N_3092);
nand U3159 (N_3159,N_3006,N_3025);
and U3160 (N_3160,N_3031,N_3006);
nor U3161 (N_3161,N_3001,N_3000);
and U3162 (N_3162,N_3006,N_3017);
or U3163 (N_3163,N_3091,N_3047);
or U3164 (N_3164,N_3052,N_3039);
xor U3165 (N_3165,N_3047,N_3087);
nor U3166 (N_3166,N_3060,N_3000);
and U3167 (N_3167,N_3043,N_3022);
xor U3168 (N_3168,N_3055,N_3080);
nor U3169 (N_3169,N_3084,N_3006);
and U3170 (N_3170,N_3025,N_3035);
nor U3171 (N_3171,N_3086,N_3048);
and U3172 (N_3172,N_3083,N_3071);
or U3173 (N_3173,N_3008,N_3089);
nand U3174 (N_3174,N_3045,N_3000);
or U3175 (N_3175,N_3007,N_3047);
xnor U3176 (N_3176,N_3054,N_3087);
or U3177 (N_3177,N_3014,N_3022);
and U3178 (N_3178,N_3018,N_3075);
nand U3179 (N_3179,N_3014,N_3048);
xnor U3180 (N_3180,N_3071,N_3046);
or U3181 (N_3181,N_3036,N_3076);
nor U3182 (N_3182,N_3088,N_3032);
nand U3183 (N_3183,N_3083,N_3041);
or U3184 (N_3184,N_3009,N_3059);
nor U3185 (N_3185,N_3053,N_3088);
nand U3186 (N_3186,N_3051,N_3037);
xor U3187 (N_3187,N_3024,N_3031);
nor U3188 (N_3188,N_3068,N_3043);
nor U3189 (N_3189,N_3019,N_3008);
nor U3190 (N_3190,N_3030,N_3002);
xnor U3191 (N_3191,N_3098,N_3073);
xor U3192 (N_3192,N_3020,N_3043);
nand U3193 (N_3193,N_3071,N_3073);
xor U3194 (N_3194,N_3066,N_3059);
and U3195 (N_3195,N_3056,N_3082);
or U3196 (N_3196,N_3069,N_3034);
nor U3197 (N_3197,N_3083,N_3029);
nand U3198 (N_3198,N_3062,N_3052);
nand U3199 (N_3199,N_3035,N_3088);
and U3200 (N_3200,N_3174,N_3122);
xor U3201 (N_3201,N_3147,N_3182);
nor U3202 (N_3202,N_3113,N_3157);
nor U3203 (N_3203,N_3184,N_3178);
and U3204 (N_3204,N_3180,N_3172);
and U3205 (N_3205,N_3127,N_3192);
xnor U3206 (N_3206,N_3156,N_3168);
xnor U3207 (N_3207,N_3139,N_3163);
nor U3208 (N_3208,N_3176,N_3189);
nor U3209 (N_3209,N_3165,N_3120);
or U3210 (N_3210,N_3193,N_3121);
xnor U3211 (N_3211,N_3128,N_3146);
xor U3212 (N_3212,N_3132,N_3153);
and U3213 (N_3213,N_3135,N_3166);
and U3214 (N_3214,N_3133,N_3105);
and U3215 (N_3215,N_3124,N_3130);
nor U3216 (N_3216,N_3143,N_3195);
nand U3217 (N_3217,N_3179,N_3117);
xnor U3218 (N_3218,N_3118,N_3142);
or U3219 (N_3219,N_3114,N_3112);
xnor U3220 (N_3220,N_3162,N_3167);
or U3221 (N_3221,N_3136,N_3164);
xnor U3222 (N_3222,N_3197,N_3129);
and U3223 (N_3223,N_3110,N_3151);
xnor U3224 (N_3224,N_3196,N_3123);
nand U3225 (N_3225,N_3131,N_3108);
nand U3226 (N_3226,N_3169,N_3111);
xnor U3227 (N_3227,N_3140,N_3116);
nor U3228 (N_3228,N_3119,N_3155);
and U3229 (N_3229,N_3191,N_3183);
nor U3230 (N_3230,N_3190,N_3138);
nand U3231 (N_3231,N_3186,N_3106);
or U3232 (N_3232,N_3109,N_3194);
or U3233 (N_3233,N_3126,N_3198);
xor U3234 (N_3234,N_3175,N_3134);
nor U3235 (N_3235,N_3161,N_3141);
and U3236 (N_3236,N_3159,N_3137);
nor U3237 (N_3237,N_3160,N_3152);
nand U3238 (N_3238,N_3145,N_3148);
and U3239 (N_3239,N_3171,N_3185);
and U3240 (N_3240,N_3115,N_3158);
or U3241 (N_3241,N_3150,N_3177);
xor U3242 (N_3242,N_3103,N_3104);
xor U3243 (N_3243,N_3187,N_3149);
nand U3244 (N_3244,N_3173,N_3100);
nand U3245 (N_3245,N_3107,N_3199);
nand U3246 (N_3246,N_3188,N_3170);
nor U3247 (N_3247,N_3181,N_3144);
xnor U3248 (N_3248,N_3101,N_3125);
or U3249 (N_3249,N_3102,N_3154);
nand U3250 (N_3250,N_3124,N_3160);
or U3251 (N_3251,N_3112,N_3185);
nor U3252 (N_3252,N_3175,N_3186);
or U3253 (N_3253,N_3137,N_3104);
nor U3254 (N_3254,N_3115,N_3143);
xnor U3255 (N_3255,N_3104,N_3136);
nand U3256 (N_3256,N_3124,N_3151);
xnor U3257 (N_3257,N_3125,N_3197);
xnor U3258 (N_3258,N_3147,N_3162);
xor U3259 (N_3259,N_3125,N_3172);
and U3260 (N_3260,N_3183,N_3177);
nor U3261 (N_3261,N_3136,N_3130);
xnor U3262 (N_3262,N_3111,N_3127);
nand U3263 (N_3263,N_3122,N_3110);
or U3264 (N_3264,N_3188,N_3158);
or U3265 (N_3265,N_3105,N_3166);
xor U3266 (N_3266,N_3196,N_3145);
and U3267 (N_3267,N_3150,N_3144);
xor U3268 (N_3268,N_3185,N_3174);
and U3269 (N_3269,N_3132,N_3120);
and U3270 (N_3270,N_3131,N_3141);
xnor U3271 (N_3271,N_3107,N_3192);
or U3272 (N_3272,N_3126,N_3129);
xor U3273 (N_3273,N_3182,N_3150);
or U3274 (N_3274,N_3146,N_3112);
and U3275 (N_3275,N_3107,N_3119);
and U3276 (N_3276,N_3158,N_3122);
and U3277 (N_3277,N_3116,N_3122);
or U3278 (N_3278,N_3112,N_3157);
or U3279 (N_3279,N_3199,N_3151);
or U3280 (N_3280,N_3157,N_3160);
and U3281 (N_3281,N_3183,N_3161);
nand U3282 (N_3282,N_3103,N_3198);
nor U3283 (N_3283,N_3189,N_3140);
nor U3284 (N_3284,N_3181,N_3102);
and U3285 (N_3285,N_3180,N_3188);
xnor U3286 (N_3286,N_3144,N_3131);
or U3287 (N_3287,N_3155,N_3170);
xnor U3288 (N_3288,N_3172,N_3144);
nor U3289 (N_3289,N_3104,N_3197);
or U3290 (N_3290,N_3162,N_3163);
nor U3291 (N_3291,N_3118,N_3170);
nand U3292 (N_3292,N_3173,N_3147);
nand U3293 (N_3293,N_3186,N_3149);
nand U3294 (N_3294,N_3162,N_3176);
or U3295 (N_3295,N_3119,N_3149);
xor U3296 (N_3296,N_3113,N_3164);
xor U3297 (N_3297,N_3193,N_3145);
nand U3298 (N_3298,N_3158,N_3173);
and U3299 (N_3299,N_3160,N_3142);
nand U3300 (N_3300,N_3236,N_3252);
nand U3301 (N_3301,N_3222,N_3262);
xor U3302 (N_3302,N_3272,N_3221);
and U3303 (N_3303,N_3261,N_3244);
xor U3304 (N_3304,N_3277,N_3285);
or U3305 (N_3305,N_3240,N_3228);
nor U3306 (N_3306,N_3284,N_3219);
nand U3307 (N_3307,N_3263,N_3220);
or U3308 (N_3308,N_3283,N_3259);
or U3309 (N_3309,N_3208,N_3212);
nor U3310 (N_3310,N_3250,N_3274);
nor U3311 (N_3311,N_3280,N_3276);
or U3312 (N_3312,N_3264,N_3286);
and U3313 (N_3313,N_3265,N_3282);
or U3314 (N_3314,N_3267,N_3239);
nand U3315 (N_3315,N_3205,N_3203);
nor U3316 (N_3316,N_3278,N_3216);
nor U3317 (N_3317,N_3245,N_3213);
or U3318 (N_3318,N_3233,N_3232);
and U3319 (N_3319,N_3255,N_3229);
and U3320 (N_3320,N_3269,N_3260);
nor U3321 (N_3321,N_3248,N_3257);
or U3322 (N_3322,N_3209,N_3218);
or U3323 (N_3323,N_3210,N_3243);
nor U3324 (N_3324,N_3200,N_3247);
or U3325 (N_3325,N_3227,N_3225);
nor U3326 (N_3326,N_3242,N_3254);
xnor U3327 (N_3327,N_3281,N_3224);
and U3328 (N_3328,N_3256,N_3298);
and U3329 (N_3329,N_3253,N_3202);
nor U3330 (N_3330,N_3204,N_3295);
nor U3331 (N_3331,N_3294,N_3258);
and U3332 (N_3332,N_3249,N_3296);
nor U3333 (N_3333,N_3238,N_3235);
and U3334 (N_3334,N_3291,N_3207);
nor U3335 (N_3335,N_3237,N_3211);
nand U3336 (N_3336,N_3292,N_3273);
and U3337 (N_3337,N_3206,N_3217);
or U3338 (N_3338,N_3230,N_3251);
or U3339 (N_3339,N_3271,N_3293);
or U3340 (N_3340,N_3275,N_3226);
or U3341 (N_3341,N_3214,N_3297);
xnor U3342 (N_3342,N_3289,N_3223);
nor U3343 (N_3343,N_3246,N_3288);
nor U3344 (N_3344,N_3268,N_3299);
nand U3345 (N_3345,N_3287,N_3231);
nand U3346 (N_3346,N_3234,N_3215);
and U3347 (N_3347,N_3270,N_3266);
xnor U3348 (N_3348,N_3201,N_3290);
and U3349 (N_3349,N_3279,N_3241);
nor U3350 (N_3350,N_3222,N_3228);
nand U3351 (N_3351,N_3248,N_3289);
xor U3352 (N_3352,N_3246,N_3290);
or U3353 (N_3353,N_3260,N_3281);
nand U3354 (N_3354,N_3278,N_3280);
xnor U3355 (N_3355,N_3288,N_3253);
and U3356 (N_3356,N_3273,N_3255);
and U3357 (N_3357,N_3251,N_3281);
xnor U3358 (N_3358,N_3277,N_3202);
and U3359 (N_3359,N_3295,N_3271);
xnor U3360 (N_3360,N_3221,N_3227);
nand U3361 (N_3361,N_3253,N_3201);
nor U3362 (N_3362,N_3201,N_3218);
or U3363 (N_3363,N_3233,N_3214);
and U3364 (N_3364,N_3207,N_3288);
nand U3365 (N_3365,N_3212,N_3275);
xor U3366 (N_3366,N_3219,N_3275);
nor U3367 (N_3367,N_3208,N_3200);
nor U3368 (N_3368,N_3207,N_3270);
nor U3369 (N_3369,N_3266,N_3246);
or U3370 (N_3370,N_3267,N_3279);
and U3371 (N_3371,N_3203,N_3220);
or U3372 (N_3372,N_3226,N_3260);
xnor U3373 (N_3373,N_3278,N_3225);
nor U3374 (N_3374,N_3235,N_3285);
and U3375 (N_3375,N_3254,N_3255);
xnor U3376 (N_3376,N_3204,N_3262);
or U3377 (N_3377,N_3297,N_3206);
and U3378 (N_3378,N_3269,N_3266);
or U3379 (N_3379,N_3245,N_3277);
nor U3380 (N_3380,N_3213,N_3279);
nor U3381 (N_3381,N_3237,N_3297);
xor U3382 (N_3382,N_3264,N_3262);
or U3383 (N_3383,N_3229,N_3237);
nand U3384 (N_3384,N_3281,N_3241);
nor U3385 (N_3385,N_3270,N_3239);
or U3386 (N_3386,N_3285,N_3230);
nand U3387 (N_3387,N_3273,N_3241);
nand U3388 (N_3388,N_3226,N_3223);
and U3389 (N_3389,N_3252,N_3254);
and U3390 (N_3390,N_3265,N_3200);
and U3391 (N_3391,N_3243,N_3260);
nor U3392 (N_3392,N_3234,N_3210);
nor U3393 (N_3393,N_3234,N_3229);
and U3394 (N_3394,N_3234,N_3243);
nor U3395 (N_3395,N_3220,N_3282);
nor U3396 (N_3396,N_3248,N_3226);
or U3397 (N_3397,N_3204,N_3297);
or U3398 (N_3398,N_3287,N_3206);
nand U3399 (N_3399,N_3249,N_3225);
xnor U3400 (N_3400,N_3372,N_3324);
or U3401 (N_3401,N_3337,N_3358);
nor U3402 (N_3402,N_3377,N_3392);
and U3403 (N_3403,N_3332,N_3344);
xnor U3404 (N_3404,N_3389,N_3349);
and U3405 (N_3405,N_3338,N_3348);
xnor U3406 (N_3406,N_3374,N_3347);
and U3407 (N_3407,N_3306,N_3315);
nand U3408 (N_3408,N_3346,N_3399);
or U3409 (N_3409,N_3376,N_3303);
or U3410 (N_3410,N_3368,N_3331);
nand U3411 (N_3411,N_3386,N_3381);
nor U3412 (N_3412,N_3353,N_3341);
nand U3413 (N_3413,N_3305,N_3339);
nand U3414 (N_3414,N_3340,N_3307);
nor U3415 (N_3415,N_3330,N_3327);
xor U3416 (N_3416,N_3383,N_3370);
and U3417 (N_3417,N_3336,N_3388);
xnor U3418 (N_3418,N_3334,N_3363);
and U3419 (N_3419,N_3395,N_3397);
and U3420 (N_3420,N_3355,N_3316);
xor U3421 (N_3421,N_3352,N_3321);
and U3422 (N_3422,N_3328,N_3359);
nand U3423 (N_3423,N_3385,N_3343);
and U3424 (N_3424,N_3329,N_3354);
or U3425 (N_3425,N_3371,N_3373);
nand U3426 (N_3426,N_3393,N_3320);
and U3427 (N_3427,N_3322,N_3351);
or U3428 (N_3428,N_3364,N_3345);
and U3429 (N_3429,N_3301,N_3323);
xnor U3430 (N_3430,N_3317,N_3304);
xor U3431 (N_3431,N_3380,N_3379);
xnor U3432 (N_3432,N_3387,N_3394);
xnor U3433 (N_3433,N_3360,N_3333);
and U3434 (N_3434,N_3312,N_3398);
nor U3435 (N_3435,N_3361,N_3362);
nand U3436 (N_3436,N_3309,N_3308);
xor U3437 (N_3437,N_3325,N_3365);
xor U3438 (N_3438,N_3378,N_3318);
and U3439 (N_3439,N_3319,N_3367);
nand U3440 (N_3440,N_3391,N_3350);
and U3441 (N_3441,N_3369,N_3326);
xnor U3442 (N_3442,N_3375,N_3310);
xnor U3443 (N_3443,N_3384,N_3300);
or U3444 (N_3444,N_3342,N_3396);
and U3445 (N_3445,N_3313,N_3390);
and U3446 (N_3446,N_3382,N_3357);
xnor U3447 (N_3447,N_3311,N_3314);
and U3448 (N_3448,N_3356,N_3302);
xor U3449 (N_3449,N_3335,N_3366);
nand U3450 (N_3450,N_3321,N_3309);
xor U3451 (N_3451,N_3375,N_3395);
or U3452 (N_3452,N_3319,N_3342);
or U3453 (N_3453,N_3374,N_3346);
xor U3454 (N_3454,N_3374,N_3315);
and U3455 (N_3455,N_3334,N_3353);
xnor U3456 (N_3456,N_3327,N_3341);
nor U3457 (N_3457,N_3380,N_3358);
nor U3458 (N_3458,N_3373,N_3334);
nor U3459 (N_3459,N_3324,N_3394);
and U3460 (N_3460,N_3371,N_3313);
and U3461 (N_3461,N_3329,N_3364);
and U3462 (N_3462,N_3363,N_3384);
nand U3463 (N_3463,N_3366,N_3354);
or U3464 (N_3464,N_3396,N_3359);
and U3465 (N_3465,N_3355,N_3374);
nand U3466 (N_3466,N_3303,N_3391);
nor U3467 (N_3467,N_3378,N_3355);
or U3468 (N_3468,N_3327,N_3343);
or U3469 (N_3469,N_3307,N_3313);
nand U3470 (N_3470,N_3366,N_3369);
xnor U3471 (N_3471,N_3358,N_3300);
nand U3472 (N_3472,N_3372,N_3367);
nor U3473 (N_3473,N_3334,N_3340);
xor U3474 (N_3474,N_3386,N_3311);
and U3475 (N_3475,N_3330,N_3378);
and U3476 (N_3476,N_3375,N_3380);
or U3477 (N_3477,N_3382,N_3361);
and U3478 (N_3478,N_3398,N_3308);
nor U3479 (N_3479,N_3318,N_3390);
nor U3480 (N_3480,N_3321,N_3329);
and U3481 (N_3481,N_3344,N_3334);
nor U3482 (N_3482,N_3373,N_3387);
or U3483 (N_3483,N_3317,N_3351);
xnor U3484 (N_3484,N_3364,N_3306);
nor U3485 (N_3485,N_3304,N_3387);
or U3486 (N_3486,N_3324,N_3384);
xor U3487 (N_3487,N_3363,N_3342);
and U3488 (N_3488,N_3374,N_3359);
nand U3489 (N_3489,N_3372,N_3319);
nand U3490 (N_3490,N_3341,N_3388);
or U3491 (N_3491,N_3339,N_3301);
xnor U3492 (N_3492,N_3368,N_3312);
or U3493 (N_3493,N_3377,N_3396);
nor U3494 (N_3494,N_3336,N_3325);
or U3495 (N_3495,N_3349,N_3373);
nor U3496 (N_3496,N_3369,N_3398);
nand U3497 (N_3497,N_3337,N_3312);
or U3498 (N_3498,N_3305,N_3350);
or U3499 (N_3499,N_3385,N_3311);
xnor U3500 (N_3500,N_3418,N_3439);
and U3501 (N_3501,N_3477,N_3436);
and U3502 (N_3502,N_3416,N_3454);
nand U3503 (N_3503,N_3433,N_3429);
nand U3504 (N_3504,N_3458,N_3456);
nor U3505 (N_3505,N_3486,N_3470);
and U3506 (N_3506,N_3484,N_3450);
nand U3507 (N_3507,N_3401,N_3400);
or U3508 (N_3508,N_3423,N_3421);
nor U3509 (N_3509,N_3499,N_3471);
nand U3510 (N_3510,N_3452,N_3478);
xnor U3511 (N_3511,N_3409,N_3414);
nand U3512 (N_3512,N_3437,N_3406);
nor U3513 (N_3513,N_3435,N_3492);
xor U3514 (N_3514,N_3428,N_3467);
and U3515 (N_3515,N_3404,N_3495);
and U3516 (N_3516,N_3475,N_3473);
nor U3517 (N_3517,N_3408,N_3403);
xor U3518 (N_3518,N_3446,N_3424);
nand U3519 (N_3519,N_3407,N_3417);
or U3520 (N_3520,N_3430,N_3419);
or U3521 (N_3521,N_3405,N_3472);
or U3522 (N_3522,N_3447,N_3459);
nand U3523 (N_3523,N_3402,N_3426);
xnor U3524 (N_3524,N_3457,N_3415);
and U3525 (N_3525,N_3448,N_3462);
and U3526 (N_3526,N_3451,N_3411);
or U3527 (N_3527,N_3464,N_3413);
xor U3528 (N_3528,N_3420,N_3412);
nor U3529 (N_3529,N_3443,N_3483);
xnor U3530 (N_3530,N_3476,N_3491);
and U3531 (N_3531,N_3485,N_3449);
or U3532 (N_3532,N_3480,N_3494);
and U3533 (N_3533,N_3427,N_3432);
nor U3534 (N_3534,N_3482,N_3490);
and U3535 (N_3535,N_3489,N_3445);
and U3536 (N_3536,N_3487,N_3444);
nor U3537 (N_3537,N_3440,N_3425);
and U3538 (N_3538,N_3466,N_3422);
or U3539 (N_3539,N_3460,N_3468);
or U3540 (N_3540,N_3442,N_3463);
and U3541 (N_3541,N_3455,N_3461);
or U3542 (N_3542,N_3474,N_3453);
nand U3543 (N_3543,N_3434,N_3479);
nand U3544 (N_3544,N_3481,N_3410);
xor U3545 (N_3545,N_3488,N_3497);
xor U3546 (N_3546,N_3469,N_3438);
or U3547 (N_3547,N_3496,N_3431);
nand U3548 (N_3548,N_3498,N_3441);
nand U3549 (N_3549,N_3493,N_3465);
and U3550 (N_3550,N_3470,N_3489);
nand U3551 (N_3551,N_3456,N_3432);
xnor U3552 (N_3552,N_3451,N_3424);
xor U3553 (N_3553,N_3450,N_3478);
and U3554 (N_3554,N_3470,N_3444);
or U3555 (N_3555,N_3451,N_3425);
nand U3556 (N_3556,N_3444,N_3485);
nor U3557 (N_3557,N_3451,N_3423);
and U3558 (N_3558,N_3446,N_3485);
nor U3559 (N_3559,N_3446,N_3479);
xor U3560 (N_3560,N_3490,N_3436);
or U3561 (N_3561,N_3400,N_3450);
xor U3562 (N_3562,N_3485,N_3423);
or U3563 (N_3563,N_3447,N_3475);
or U3564 (N_3564,N_3457,N_3446);
or U3565 (N_3565,N_3442,N_3444);
nand U3566 (N_3566,N_3475,N_3471);
xnor U3567 (N_3567,N_3464,N_3441);
xnor U3568 (N_3568,N_3463,N_3494);
nor U3569 (N_3569,N_3450,N_3423);
or U3570 (N_3570,N_3429,N_3493);
nor U3571 (N_3571,N_3471,N_3445);
and U3572 (N_3572,N_3410,N_3404);
or U3573 (N_3573,N_3412,N_3461);
nor U3574 (N_3574,N_3411,N_3460);
nand U3575 (N_3575,N_3423,N_3430);
nand U3576 (N_3576,N_3496,N_3454);
nor U3577 (N_3577,N_3466,N_3436);
nand U3578 (N_3578,N_3446,N_3458);
or U3579 (N_3579,N_3424,N_3444);
xor U3580 (N_3580,N_3488,N_3425);
and U3581 (N_3581,N_3444,N_3432);
or U3582 (N_3582,N_3429,N_3430);
xor U3583 (N_3583,N_3435,N_3486);
or U3584 (N_3584,N_3472,N_3418);
nand U3585 (N_3585,N_3495,N_3433);
or U3586 (N_3586,N_3450,N_3446);
xnor U3587 (N_3587,N_3459,N_3418);
nor U3588 (N_3588,N_3475,N_3496);
nand U3589 (N_3589,N_3404,N_3454);
or U3590 (N_3590,N_3407,N_3490);
or U3591 (N_3591,N_3482,N_3401);
nand U3592 (N_3592,N_3484,N_3469);
nor U3593 (N_3593,N_3444,N_3468);
and U3594 (N_3594,N_3469,N_3463);
or U3595 (N_3595,N_3471,N_3437);
and U3596 (N_3596,N_3478,N_3430);
nor U3597 (N_3597,N_3406,N_3447);
nor U3598 (N_3598,N_3479,N_3492);
and U3599 (N_3599,N_3477,N_3462);
xor U3600 (N_3600,N_3584,N_3510);
nor U3601 (N_3601,N_3526,N_3541);
or U3602 (N_3602,N_3594,N_3557);
xnor U3603 (N_3603,N_3525,N_3578);
or U3604 (N_3604,N_3555,N_3560);
nand U3605 (N_3605,N_3536,N_3576);
or U3606 (N_3606,N_3595,N_3501);
xor U3607 (N_3607,N_3551,N_3565);
nor U3608 (N_3608,N_3500,N_3567);
nor U3609 (N_3609,N_3558,N_3549);
and U3610 (N_3610,N_3599,N_3531);
xnor U3611 (N_3611,N_3529,N_3527);
nor U3612 (N_3612,N_3568,N_3596);
xor U3613 (N_3613,N_3559,N_3538);
nand U3614 (N_3614,N_3515,N_3547);
and U3615 (N_3615,N_3561,N_3553);
and U3616 (N_3616,N_3519,N_3514);
and U3617 (N_3617,N_3574,N_3548);
nand U3618 (N_3618,N_3522,N_3581);
xor U3619 (N_3619,N_3542,N_3521);
nand U3620 (N_3620,N_3545,N_3552);
or U3621 (N_3621,N_3573,N_3512);
nand U3622 (N_3622,N_3563,N_3585);
nand U3623 (N_3623,N_3537,N_3506);
xor U3624 (N_3624,N_3566,N_3523);
nor U3625 (N_3625,N_3524,N_3546);
xor U3626 (N_3626,N_3588,N_3535);
nand U3627 (N_3627,N_3532,N_3569);
nand U3628 (N_3628,N_3580,N_3598);
nor U3629 (N_3629,N_3575,N_3539);
and U3630 (N_3630,N_3533,N_3520);
or U3631 (N_3631,N_3583,N_3562);
nor U3632 (N_3632,N_3564,N_3556);
xor U3633 (N_3633,N_3505,N_3592);
nand U3634 (N_3634,N_3597,N_3572);
and U3635 (N_3635,N_3586,N_3571);
nor U3636 (N_3636,N_3589,N_3579);
nand U3637 (N_3637,N_3570,N_3543);
nand U3638 (N_3638,N_3516,N_3577);
or U3639 (N_3639,N_3544,N_3587);
nor U3640 (N_3640,N_3591,N_3504);
xor U3641 (N_3641,N_3590,N_3503);
and U3642 (N_3642,N_3534,N_3550);
nor U3643 (N_3643,N_3518,N_3582);
or U3644 (N_3644,N_3502,N_3508);
nor U3645 (N_3645,N_3530,N_3507);
xnor U3646 (N_3646,N_3511,N_3593);
xnor U3647 (N_3647,N_3509,N_3517);
nand U3648 (N_3648,N_3540,N_3528);
nand U3649 (N_3649,N_3554,N_3513);
and U3650 (N_3650,N_3559,N_3579);
nand U3651 (N_3651,N_3597,N_3552);
and U3652 (N_3652,N_3546,N_3535);
and U3653 (N_3653,N_3592,N_3543);
or U3654 (N_3654,N_3581,N_3569);
nor U3655 (N_3655,N_3539,N_3533);
or U3656 (N_3656,N_3571,N_3527);
and U3657 (N_3657,N_3560,N_3588);
nor U3658 (N_3658,N_3587,N_3510);
or U3659 (N_3659,N_3577,N_3572);
xor U3660 (N_3660,N_3553,N_3576);
nor U3661 (N_3661,N_3532,N_3519);
nand U3662 (N_3662,N_3537,N_3573);
xnor U3663 (N_3663,N_3530,N_3570);
nand U3664 (N_3664,N_3580,N_3540);
and U3665 (N_3665,N_3575,N_3546);
or U3666 (N_3666,N_3582,N_3566);
and U3667 (N_3667,N_3546,N_3513);
nand U3668 (N_3668,N_3562,N_3535);
nor U3669 (N_3669,N_3593,N_3595);
nor U3670 (N_3670,N_3515,N_3525);
nand U3671 (N_3671,N_3562,N_3592);
and U3672 (N_3672,N_3524,N_3554);
nand U3673 (N_3673,N_3563,N_3534);
xnor U3674 (N_3674,N_3580,N_3582);
xor U3675 (N_3675,N_3598,N_3528);
nor U3676 (N_3676,N_3579,N_3532);
xor U3677 (N_3677,N_3555,N_3514);
xor U3678 (N_3678,N_3533,N_3507);
and U3679 (N_3679,N_3587,N_3579);
nand U3680 (N_3680,N_3566,N_3577);
nand U3681 (N_3681,N_3579,N_3562);
and U3682 (N_3682,N_3596,N_3586);
or U3683 (N_3683,N_3532,N_3553);
and U3684 (N_3684,N_3597,N_3530);
or U3685 (N_3685,N_3553,N_3591);
nand U3686 (N_3686,N_3502,N_3536);
nor U3687 (N_3687,N_3550,N_3553);
nand U3688 (N_3688,N_3506,N_3574);
or U3689 (N_3689,N_3567,N_3597);
or U3690 (N_3690,N_3584,N_3563);
xor U3691 (N_3691,N_3575,N_3547);
nand U3692 (N_3692,N_3507,N_3560);
nor U3693 (N_3693,N_3501,N_3545);
xnor U3694 (N_3694,N_3565,N_3577);
nand U3695 (N_3695,N_3523,N_3535);
or U3696 (N_3696,N_3535,N_3584);
or U3697 (N_3697,N_3546,N_3504);
nand U3698 (N_3698,N_3559,N_3585);
xor U3699 (N_3699,N_3550,N_3548);
nand U3700 (N_3700,N_3668,N_3677);
or U3701 (N_3701,N_3662,N_3690);
xor U3702 (N_3702,N_3656,N_3626);
nand U3703 (N_3703,N_3619,N_3658);
and U3704 (N_3704,N_3628,N_3676);
xor U3705 (N_3705,N_3608,N_3603);
nor U3706 (N_3706,N_3661,N_3694);
xnor U3707 (N_3707,N_3614,N_3645);
nor U3708 (N_3708,N_3646,N_3625);
or U3709 (N_3709,N_3674,N_3657);
and U3710 (N_3710,N_3652,N_3687);
nand U3711 (N_3711,N_3648,N_3680);
or U3712 (N_3712,N_3612,N_3621);
and U3713 (N_3713,N_3613,N_3692);
and U3714 (N_3714,N_3671,N_3649);
and U3715 (N_3715,N_3643,N_3655);
or U3716 (N_3716,N_3650,N_3631);
nor U3717 (N_3717,N_3600,N_3601);
nand U3718 (N_3718,N_3602,N_3605);
or U3719 (N_3719,N_3675,N_3624);
or U3720 (N_3720,N_3691,N_3618);
and U3721 (N_3721,N_3635,N_3667);
or U3722 (N_3722,N_3670,N_3653);
nor U3723 (N_3723,N_3654,N_3647);
nor U3724 (N_3724,N_3607,N_3660);
or U3725 (N_3725,N_3684,N_3610);
nor U3726 (N_3726,N_3609,N_3634);
nand U3727 (N_3727,N_3632,N_3615);
nor U3728 (N_3728,N_3686,N_3688);
xor U3729 (N_3729,N_3636,N_3616);
or U3730 (N_3730,N_3681,N_3640);
nand U3731 (N_3731,N_3642,N_3693);
nor U3732 (N_3732,N_3678,N_3604);
and U3733 (N_3733,N_3630,N_3659);
nand U3734 (N_3734,N_3689,N_3637);
or U3735 (N_3735,N_3673,N_3696);
nor U3736 (N_3736,N_3669,N_3695);
nand U3737 (N_3737,N_3641,N_3620);
and U3738 (N_3738,N_3663,N_3629);
nand U3739 (N_3739,N_3697,N_3679);
xor U3740 (N_3740,N_3623,N_3606);
nand U3741 (N_3741,N_3639,N_3651);
nand U3742 (N_3742,N_3682,N_3666);
or U3743 (N_3743,N_3683,N_3617);
or U3744 (N_3744,N_3672,N_3633);
xnor U3745 (N_3745,N_3611,N_3664);
nor U3746 (N_3746,N_3644,N_3698);
nor U3747 (N_3747,N_3638,N_3622);
and U3748 (N_3748,N_3627,N_3665);
nor U3749 (N_3749,N_3685,N_3699);
nand U3750 (N_3750,N_3672,N_3645);
nor U3751 (N_3751,N_3668,N_3667);
nand U3752 (N_3752,N_3670,N_3683);
and U3753 (N_3753,N_3604,N_3644);
and U3754 (N_3754,N_3621,N_3671);
nand U3755 (N_3755,N_3601,N_3624);
nand U3756 (N_3756,N_3628,N_3642);
or U3757 (N_3757,N_3661,N_3688);
xor U3758 (N_3758,N_3660,N_3681);
xor U3759 (N_3759,N_3696,N_3625);
and U3760 (N_3760,N_3628,N_3645);
xor U3761 (N_3761,N_3693,N_3682);
xnor U3762 (N_3762,N_3647,N_3622);
xnor U3763 (N_3763,N_3656,N_3657);
or U3764 (N_3764,N_3669,N_3674);
nor U3765 (N_3765,N_3629,N_3645);
nor U3766 (N_3766,N_3644,N_3680);
nor U3767 (N_3767,N_3605,N_3674);
and U3768 (N_3768,N_3653,N_3614);
nand U3769 (N_3769,N_3605,N_3625);
and U3770 (N_3770,N_3693,N_3641);
xnor U3771 (N_3771,N_3691,N_3649);
or U3772 (N_3772,N_3629,N_3606);
nor U3773 (N_3773,N_3697,N_3622);
and U3774 (N_3774,N_3655,N_3660);
nor U3775 (N_3775,N_3676,N_3607);
nand U3776 (N_3776,N_3681,N_3686);
or U3777 (N_3777,N_3683,N_3622);
and U3778 (N_3778,N_3626,N_3691);
and U3779 (N_3779,N_3617,N_3612);
or U3780 (N_3780,N_3676,N_3600);
nand U3781 (N_3781,N_3642,N_3665);
nand U3782 (N_3782,N_3687,N_3682);
and U3783 (N_3783,N_3640,N_3657);
nor U3784 (N_3784,N_3658,N_3661);
and U3785 (N_3785,N_3671,N_3650);
nand U3786 (N_3786,N_3696,N_3605);
and U3787 (N_3787,N_3606,N_3639);
or U3788 (N_3788,N_3630,N_3638);
nor U3789 (N_3789,N_3621,N_3663);
or U3790 (N_3790,N_3642,N_3616);
nand U3791 (N_3791,N_3644,N_3661);
and U3792 (N_3792,N_3678,N_3657);
or U3793 (N_3793,N_3608,N_3636);
or U3794 (N_3794,N_3665,N_3695);
or U3795 (N_3795,N_3697,N_3659);
xor U3796 (N_3796,N_3617,N_3606);
nand U3797 (N_3797,N_3695,N_3680);
nand U3798 (N_3798,N_3666,N_3632);
and U3799 (N_3799,N_3685,N_3696);
or U3800 (N_3800,N_3784,N_3799);
nor U3801 (N_3801,N_3701,N_3758);
or U3802 (N_3802,N_3772,N_3794);
nor U3803 (N_3803,N_3722,N_3743);
and U3804 (N_3804,N_3707,N_3714);
or U3805 (N_3805,N_3749,N_3785);
xnor U3806 (N_3806,N_3765,N_3764);
and U3807 (N_3807,N_3730,N_3709);
and U3808 (N_3808,N_3735,N_3766);
or U3809 (N_3809,N_3780,N_3754);
or U3810 (N_3810,N_3751,N_3711);
nand U3811 (N_3811,N_3737,N_3795);
and U3812 (N_3812,N_3742,N_3752);
xor U3813 (N_3813,N_3725,N_3706);
or U3814 (N_3814,N_3715,N_3762);
or U3815 (N_3815,N_3724,N_3729);
or U3816 (N_3816,N_3787,N_3727);
xor U3817 (N_3817,N_3763,N_3741);
nor U3818 (N_3818,N_3704,N_3733);
and U3819 (N_3819,N_3790,N_3759);
and U3820 (N_3820,N_3775,N_3700);
nor U3821 (N_3821,N_3728,N_3761);
xor U3822 (N_3822,N_3753,N_3757);
nor U3823 (N_3823,N_3779,N_3720);
nor U3824 (N_3824,N_3755,N_3767);
or U3825 (N_3825,N_3726,N_3716);
and U3826 (N_3826,N_3770,N_3731);
xnor U3827 (N_3827,N_3782,N_3708);
and U3828 (N_3828,N_3776,N_3793);
and U3829 (N_3829,N_3791,N_3781);
nor U3830 (N_3830,N_3718,N_3797);
or U3831 (N_3831,N_3712,N_3705);
xor U3832 (N_3832,N_3748,N_3798);
xnor U3833 (N_3833,N_3703,N_3710);
nand U3834 (N_3834,N_3783,N_3773);
or U3835 (N_3835,N_3744,N_3771);
nand U3836 (N_3836,N_3746,N_3732);
or U3837 (N_3837,N_3789,N_3777);
xnor U3838 (N_3838,N_3745,N_3756);
and U3839 (N_3839,N_3760,N_3702);
nor U3840 (N_3840,N_3738,N_3713);
or U3841 (N_3841,N_3778,N_3774);
and U3842 (N_3842,N_3736,N_3739);
nor U3843 (N_3843,N_3796,N_3719);
xnor U3844 (N_3844,N_3723,N_3768);
nor U3845 (N_3845,N_3788,N_3721);
xor U3846 (N_3846,N_3786,N_3769);
or U3847 (N_3847,N_3792,N_3747);
xor U3848 (N_3848,N_3750,N_3734);
xor U3849 (N_3849,N_3717,N_3740);
nor U3850 (N_3850,N_3786,N_3775);
xor U3851 (N_3851,N_3768,N_3798);
or U3852 (N_3852,N_3757,N_3734);
nand U3853 (N_3853,N_3724,N_3711);
nand U3854 (N_3854,N_3720,N_3735);
xor U3855 (N_3855,N_3715,N_3787);
nand U3856 (N_3856,N_3712,N_3734);
nand U3857 (N_3857,N_3759,N_3794);
nand U3858 (N_3858,N_3768,N_3715);
nand U3859 (N_3859,N_3736,N_3721);
and U3860 (N_3860,N_3741,N_3730);
xor U3861 (N_3861,N_3773,N_3700);
or U3862 (N_3862,N_3740,N_3742);
nor U3863 (N_3863,N_3752,N_3769);
nand U3864 (N_3864,N_3722,N_3791);
nor U3865 (N_3865,N_3722,N_3760);
nor U3866 (N_3866,N_3726,N_3776);
nand U3867 (N_3867,N_3761,N_3744);
nor U3868 (N_3868,N_3768,N_3766);
nor U3869 (N_3869,N_3769,N_3719);
or U3870 (N_3870,N_3788,N_3723);
and U3871 (N_3871,N_3777,N_3713);
or U3872 (N_3872,N_3765,N_3756);
or U3873 (N_3873,N_3738,N_3733);
nand U3874 (N_3874,N_3767,N_3742);
or U3875 (N_3875,N_3771,N_3702);
nand U3876 (N_3876,N_3797,N_3724);
nor U3877 (N_3877,N_3760,N_3781);
xor U3878 (N_3878,N_3779,N_3761);
or U3879 (N_3879,N_3772,N_3716);
and U3880 (N_3880,N_3711,N_3777);
xnor U3881 (N_3881,N_3779,N_3750);
or U3882 (N_3882,N_3758,N_3708);
nor U3883 (N_3883,N_3745,N_3731);
and U3884 (N_3884,N_3736,N_3725);
nor U3885 (N_3885,N_3748,N_3767);
and U3886 (N_3886,N_3772,N_3796);
and U3887 (N_3887,N_3746,N_3701);
or U3888 (N_3888,N_3742,N_3793);
and U3889 (N_3889,N_3705,N_3780);
or U3890 (N_3890,N_3797,N_3783);
and U3891 (N_3891,N_3703,N_3706);
nor U3892 (N_3892,N_3788,N_3730);
nand U3893 (N_3893,N_3774,N_3729);
or U3894 (N_3894,N_3796,N_3765);
xor U3895 (N_3895,N_3715,N_3749);
xnor U3896 (N_3896,N_3726,N_3739);
xnor U3897 (N_3897,N_3746,N_3753);
and U3898 (N_3898,N_3760,N_3791);
xor U3899 (N_3899,N_3722,N_3737);
or U3900 (N_3900,N_3848,N_3865);
nor U3901 (N_3901,N_3831,N_3815);
xnor U3902 (N_3902,N_3811,N_3827);
xor U3903 (N_3903,N_3859,N_3899);
nand U3904 (N_3904,N_3808,N_3858);
xnor U3905 (N_3905,N_3843,N_3846);
nand U3906 (N_3906,N_3874,N_3802);
xnor U3907 (N_3907,N_3847,N_3841);
nor U3908 (N_3908,N_3885,N_3886);
nor U3909 (N_3909,N_3836,N_3849);
xor U3910 (N_3910,N_3889,N_3868);
or U3911 (N_3911,N_3879,N_3881);
nor U3912 (N_3912,N_3838,N_3807);
and U3913 (N_3913,N_3898,N_3829);
or U3914 (N_3914,N_3862,N_3896);
nand U3915 (N_3915,N_3816,N_3870);
and U3916 (N_3916,N_3852,N_3863);
xnor U3917 (N_3917,N_3825,N_3883);
nand U3918 (N_3918,N_3822,N_3869);
xor U3919 (N_3919,N_3866,N_3845);
xnor U3920 (N_3920,N_3830,N_3837);
and U3921 (N_3921,N_3835,N_3850);
nand U3922 (N_3922,N_3806,N_3860);
xnor U3923 (N_3923,N_3803,N_3804);
or U3924 (N_3924,N_3876,N_3867);
and U3925 (N_3925,N_3895,N_3891);
xnor U3926 (N_3926,N_3817,N_3834);
nand U3927 (N_3927,N_3872,N_3813);
and U3928 (N_3928,N_3833,N_3856);
xor U3929 (N_3929,N_3853,N_3819);
or U3930 (N_3930,N_3823,N_3839);
nor U3931 (N_3931,N_3892,N_3840);
xnor U3932 (N_3932,N_3855,N_3857);
nor U3933 (N_3933,N_3864,N_3809);
nand U3934 (N_3934,N_3854,N_3882);
xor U3935 (N_3935,N_3875,N_3805);
and U3936 (N_3936,N_3810,N_3890);
or U3937 (N_3937,N_3887,N_3801);
or U3938 (N_3938,N_3832,N_3826);
nor U3939 (N_3939,N_3897,N_3851);
or U3940 (N_3940,N_3800,N_3861);
nor U3941 (N_3941,N_3842,N_3884);
and U3942 (N_3942,N_3820,N_3814);
nand U3943 (N_3943,N_3894,N_3844);
xor U3944 (N_3944,N_3821,N_3871);
nor U3945 (N_3945,N_3818,N_3880);
nor U3946 (N_3946,N_3873,N_3878);
or U3947 (N_3947,N_3877,N_3812);
xor U3948 (N_3948,N_3893,N_3824);
and U3949 (N_3949,N_3888,N_3828);
nor U3950 (N_3950,N_3816,N_3863);
nor U3951 (N_3951,N_3846,N_3881);
and U3952 (N_3952,N_3891,N_3884);
xnor U3953 (N_3953,N_3807,N_3836);
xor U3954 (N_3954,N_3866,N_3850);
xor U3955 (N_3955,N_3829,N_3807);
nor U3956 (N_3956,N_3857,N_3816);
xnor U3957 (N_3957,N_3825,N_3817);
or U3958 (N_3958,N_3848,N_3816);
or U3959 (N_3959,N_3881,N_3813);
nor U3960 (N_3960,N_3823,N_3860);
and U3961 (N_3961,N_3875,N_3844);
nand U3962 (N_3962,N_3848,N_3893);
xnor U3963 (N_3963,N_3876,N_3822);
nor U3964 (N_3964,N_3823,N_3808);
xor U3965 (N_3965,N_3884,N_3817);
xnor U3966 (N_3966,N_3800,N_3837);
xor U3967 (N_3967,N_3894,N_3848);
or U3968 (N_3968,N_3858,N_3821);
nand U3969 (N_3969,N_3856,N_3841);
nand U3970 (N_3970,N_3828,N_3806);
nor U3971 (N_3971,N_3804,N_3845);
or U3972 (N_3972,N_3808,N_3819);
nor U3973 (N_3973,N_3849,N_3839);
and U3974 (N_3974,N_3878,N_3802);
or U3975 (N_3975,N_3893,N_3834);
nand U3976 (N_3976,N_3814,N_3840);
and U3977 (N_3977,N_3855,N_3825);
and U3978 (N_3978,N_3866,N_3869);
nor U3979 (N_3979,N_3805,N_3893);
or U3980 (N_3980,N_3853,N_3884);
nand U3981 (N_3981,N_3871,N_3808);
or U3982 (N_3982,N_3841,N_3889);
and U3983 (N_3983,N_3839,N_3854);
xnor U3984 (N_3984,N_3868,N_3884);
or U3985 (N_3985,N_3814,N_3866);
and U3986 (N_3986,N_3811,N_3808);
nand U3987 (N_3987,N_3825,N_3818);
xor U3988 (N_3988,N_3867,N_3819);
xnor U3989 (N_3989,N_3835,N_3806);
nor U3990 (N_3990,N_3887,N_3853);
or U3991 (N_3991,N_3898,N_3855);
or U3992 (N_3992,N_3891,N_3864);
nor U3993 (N_3993,N_3839,N_3824);
nand U3994 (N_3994,N_3823,N_3853);
nor U3995 (N_3995,N_3878,N_3858);
nor U3996 (N_3996,N_3825,N_3804);
nor U3997 (N_3997,N_3856,N_3836);
nor U3998 (N_3998,N_3858,N_3897);
nor U3999 (N_3999,N_3891,N_3840);
and U4000 (N_4000,N_3954,N_3914);
xnor U4001 (N_4001,N_3996,N_3963);
or U4002 (N_4002,N_3993,N_3988);
nor U4003 (N_4003,N_3976,N_3925);
xnor U4004 (N_4004,N_3992,N_3969);
xor U4005 (N_4005,N_3935,N_3921);
nor U4006 (N_4006,N_3972,N_3962);
nand U4007 (N_4007,N_3958,N_3922);
or U4008 (N_4008,N_3940,N_3973);
or U4009 (N_4009,N_3957,N_3952);
xnor U4010 (N_4010,N_3974,N_3989);
nand U4011 (N_4011,N_3908,N_3999);
nand U4012 (N_4012,N_3910,N_3977);
and U4013 (N_4013,N_3942,N_3941);
or U4014 (N_4014,N_3915,N_3933);
and U4015 (N_4015,N_3948,N_3911);
or U4016 (N_4016,N_3924,N_3961);
or U4017 (N_4017,N_3904,N_3929);
nand U4018 (N_4018,N_3913,N_3955);
nor U4019 (N_4019,N_3995,N_3928);
or U4020 (N_4020,N_3971,N_3938);
nor U4021 (N_4021,N_3986,N_3970);
and U4022 (N_4022,N_3953,N_3998);
or U4023 (N_4023,N_3917,N_3979);
nand U4024 (N_4024,N_3965,N_3919);
nor U4025 (N_4025,N_3981,N_3926);
or U4026 (N_4026,N_3901,N_3930);
nand U4027 (N_4027,N_3960,N_3967);
nor U4028 (N_4028,N_3906,N_3903);
or U4029 (N_4029,N_3980,N_3959);
or U4030 (N_4030,N_3956,N_3934);
xor U4031 (N_4031,N_3947,N_3918);
or U4032 (N_4032,N_3927,N_3949);
nand U4033 (N_4033,N_3944,N_3950);
nor U4034 (N_4034,N_3984,N_3909);
xor U4035 (N_4035,N_3931,N_3966);
or U4036 (N_4036,N_3964,N_3997);
nor U4037 (N_4037,N_3907,N_3912);
nand U4038 (N_4038,N_3920,N_3905);
nand U4039 (N_4039,N_3932,N_3916);
or U4040 (N_4040,N_3936,N_3982);
nand U4041 (N_4041,N_3902,N_3978);
and U4042 (N_4042,N_3983,N_3968);
xor U4043 (N_4043,N_3991,N_3945);
nor U4044 (N_4044,N_3990,N_3985);
and U4045 (N_4045,N_3939,N_3994);
nor U4046 (N_4046,N_3923,N_3943);
or U4047 (N_4047,N_3987,N_3946);
xor U4048 (N_4048,N_3975,N_3900);
nor U4049 (N_4049,N_3951,N_3937);
or U4050 (N_4050,N_3960,N_3983);
xnor U4051 (N_4051,N_3903,N_3997);
nand U4052 (N_4052,N_3969,N_3994);
nor U4053 (N_4053,N_3935,N_3918);
and U4054 (N_4054,N_3929,N_3980);
nand U4055 (N_4055,N_3948,N_3904);
nand U4056 (N_4056,N_3967,N_3943);
nand U4057 (N_4057,N_3933,N_3973);
nand U4058 (N_4058,N_3942,N_3908);
and U4059 (N_4059,N_3979,N_3955);
and U4060 (N_4060,N_3964,N_3993);
xor U4061 (N_4061,N_3940,N_3956);
and U4062 (N_4062,N_3933,N_3934);
nor U4063 (N_4063,N_3993,N_3953);
xnor U4064 (N_4064,N_3903,N_3927);
and U4065 (N_4065,N_3956,N_3920);
nor U4066 (N_4066,N_3976,N_3966);
xor U4067 (N_4067,N_3930,N_3948);
or U4068 (N_4068,N_3940,N_3913);
and U4069 (N_4069,N_3959,N_3971);
xor U4070 (N_4070,N_3989,N_3907);
nor U4071 (N_4071,N_3995,N_3936);
nor U4072 (N_4072,N_3930,N_3955);
or U4073 (N_4073,N_3915,N_3943);
and U4074 (N_4074,N_3977,N_3984);
nor U4075 (N_4075,N_3995,N_3933);
nand U4076 (N_4076,N_3982,N_3983);
or U4077 (N_4077,N_3932,N_3985);
or U4078 (N_4078,N_3954,N_3959);
xor U4079 (N_4079,N_3953,N_3990);
xor U4080 (N_4080,N_3963,N_3952);
or U4081 (N_4081,N_3902,N_3960);
and U4082 (N_4082,N_3976,N_3979);
nand U4083 (N_4083,N_3947,N_3935);
nand U4084 (N_4084,N_3974,N_3930);
nor U4085 (N_4085,N_3985,N_3931);
nor U4086 (N_4086,N_3994,N_3943);
or U4087 (N_4087,N_3988,N_3960);
and U4088 (N_4088,N_3906,N_3900);
and U4089 (N_4089,N_3998,N_3985);
xor U4090 (N_4090,N_3980,N_3921);
and U4091 (N_4091,N_3950,N_3937);
nor U4092 (N_4092,N_3963,N_3916);
or U4093 (N_4093,N_3919,N_3936);
nand U4094 (N_4094,N_3923,N_3917);
or U4095 (N_4095,N_3952,N_3953);
nand U4096 (N_4096,N_3955,N_3982);
xor U4097 (N_4097,N_3987,N_3909);
and U4098 (N_4098,N_3910,N_3960);
nor U4099 (N_4099,N_3975,N_3991);
xnor U4100 (N_4100,N_4026,N_4023);
nand U4101 (N_4101,N_4039,N_4058);
xor U4102 (N_4102,N_4017,N_4067);
nand U4103 (N_4103,N_4056,N_4097);
xnor U4104 (N_4104,N_4002,N_4006);
nor U4105 (N_4105,N_4091,N_4099);
and U4106 (N_4106,N_4094,N_4028);
or U4107 (N_4107,N_4089,N_4030);
or U4108 (N_4108,N_4083,N_4096);
nor U4109 (N_4109,N_4072,N_4005);
nor U4110 (N_4110,N_4055,N_4064);
or U4111 (N_4111,N_4013,N_4098);
nor U4112 (N_4112,N_4012,N_4016);
and U4113 (N_4113,N_4036,N_4062);
xor U4114 (N_4114,N_4073,N_4061);
xor U4115 (N_4115,N_4007,N_4088);
or U4116 (N_4116,N_4093,N_4087);
xor U4117 (N_4117,N_4020,N_4092);
nand U4118 (N_4118,N_4034,N_4024);
nand U4119 (N_4119,N_4042,N_4004);
nor U4120 (N_4120,N_4049,N_4000);
xnor U4121 (N_4121,N_4069,N_4051);
xor U4122 (N_4122,N_4003,N_4015);
or U4123 (N_4123,N_4053,N_4033);
nand U4124 (N_4124,N_4071,N_4050);
and U4125 (N_4125,N_4037,N_4022);
xor U4126 (N_4126,N_4095,N_4009);
and U4127 (N_4127,N_4054,N_4059);
nand U4128 (N_4128,N_4079,N_4085);
or U4129 (N_4129,N_4041,N_4084);
xor U4130 (N_4130,N_4076,N_4066);
xnor U4131 (N_4131,N_4078,N_4011);
nor U4132 (N_4132,N_4068,N_4047);
and U4133 (N_4133,N_4001,N_4014);
xnor U4134 (N_4134,N_4045,N_4027);
or U4135 (N_4135,N_4052,N_4046);
nor U4136 (N_4136,N_4021,N_4082);
xor U4137 (N_4137,N_4019,N_4057);
xor U4138 (N_4138,N_4038,N_4060);
xnor U4139 (N_4139,N_4063,N_4075);
or U4140 (N_4140,N_4086,N_4008);
nand U4141 (N_4141,N_4074,N_4048);
nand U4142 (N_4142,N_4070,N_4031);
nand U4143 (N_4143,N_4090,N_4018);
or U4144 (N_4144,N_4029,N_4010);
nand U4145 (N_4145,N_4025,N_4032);
nor U4146 (N_4146,N_4077,N_4080);
or U4147 (N_4147,N_4043,N_4065);
and U4148 (N_4148,N_4035,N_4040);
nand U4149 (N_4149,N_4081,N_4044);
nor U4150 (N_4150,N_4019,N_4037);
or U4151 (N_4151,N_4091,N_4000);
or U4152 (N_4152,N_4016,N_4040);
nand U4153 (N_4153,N_4057,N_4000);
xnor U4154 (N_4154,N_4056,N_4000);
nor U4155 (N_4155,N_4033,N_4018);
and U4156 (N_4156,N_4036,N_4025);
xor U4157 (N_4157,N_4005,N_4076);
nand U4158 (N_4158,N_4069,N_4002);
nor U4159 (N_4159,N_4064,N_4069);
nor U4160 (N_4160,N_4069,N_4074);
nand U4161 (N_4161,N_4084,N_4025);
xor U4162 (N_4162,N_4098,N_4033);
nand U4163 (N_4163,N_4094,N_4088);
and U4164 (N_4164,N_4025,N_4089);
and U4165 (N_4165,N_4034,N_4014);
nor U4166 (N_4166,N_4071,N_4066);
and U4167 (N_4167,N_4054,N_4025);
or U4168 (N_4168,N_4076,N_4043);
nand U4169 (N_4169,N_4096,N_4027);
and U4170 (N_4170,N_4061,N_4086);
nand U4171 (N_4171,N_4002,N_4027);
xor U4172 (N_4172,N_4079,N_4013);
nor U4173 (N_4173,N_4061,N_4053);
or U4174 (N_4174,N_4085,N_4012);
xor U4175 (N_4175,N_4032,N_4021);
nand U4176 (N_4176,N_4075,N_4068);
and U4177 (N_4177,N_4087,N_4076);
and U4178 (N_4178,N_4099,N_4024);
nand U4179 (N_4179,N_4033,N_4090);
and U4180 (N_4180,N_4058,N_4088);
xnor U4181 (N_4181,N_4021,N_4003);
and U4182 (N_4182,N_4084,N_4061);
and U4183 (N_4183,N_4040,N_4086);
nor U4184 (N_4184,N_4025,N_4047);
nand U4185 (N_4185,N_4093,N_4070);
nor U4186 (N_4186,N_4004,N_4064);
nor U4187 (N_4187,N_4068,N_4050);
or U4188 (N_4188,N_4042,N_4071);
and U4189 (N_4189,N_4073,N_4014);
nand U4190 (N_4190,N_4026,N_4094);
and U4191 (N_4191,N_4042,N_4012);
xor U4192 (N_4192,N_4088,N_4084);
and U4193 (N_4193,N_4044,N_4006);
and U4194 (N_4194,N_4013,N_4099);
nor U4195 (N_4195,N_4033,N_4085);
and U4196 (N_4196,N_4081,N_4025);
xnor U4197 (N_4197,N_4055,N_4072);
nand U4198 (N_4198,N_4081,N_4065);
or U4199 (N_4199,N_4072,N_4061);
and U4200 (N_4200,N_4176,N_4170);
nor U4201 (N_4201,N_4197,N_4160);
xnor U4202 (N_4202,N_4161,N_4139);
nor U4203 (N_4203,N_4192,N_4133);
and U4204 (N_4204,N_4121,N_4168);
or U4205 (N_4205,N_4155,N_4148);
xnor U4206 (N_4206,N_4114,N_4103);
or U4207 (N_4207,N_4162,N_4134);
nand U4208 (N_4208,N_4107,N_4123);
or U4209 (N_4209,N_4138,N_4172);
or U4210 (N_4210,N_4135,N_4194);
and U4211 (N_4211,N_4100,N_4154);
or U4212 (N_4212,N_4145,N_4129);
and U4213 (N_4213,N_4164,N_4142);
or U4214 (N_4214,N_4186,N_4151);
nand U4215 (N_4215,N_4177,N_4105);
or U4216 (N_4216,N_4195,N_4110);
or U4217 (N_4217,N_4136,N_4193);
nor U4218 (N_4218,N_4116,N_4165);
xor U4219 (N_4219,N_4131,N_4117);
and U4220 (N_4220,N_4173,N_4174);
nand U4221 (N_4221,N_4109,N_4126);
or U4222 (N_4222,N_4167,N_4189);
nor U4223 (N_4223,N_4157,N_4180);
xnor U4224 (N_4224,N_4108,N_4185);
or U4225 (N_4225,N_4178,N_4184);
nand U4226 (N_4226,N_4159,N_4146);
or U4227 (N_4227,N_4147,N_4187);
and U4228 (N_4228,N_4188,N_4130);
xnor U4229 (N_4229,N_4115,N_4149);
nor U4230 (N_4230,N_4182,N_4112);
nor U4231 (N_4231,N_4156,N_4144);
nor U4232 (N_4232,N_4181,N_4140);
nor U4233 (N_4233,N_4141,N_4152);
or U4234 (N_4234,N_4190,N_4119);
nand U4235 (N_4235,N_4166,N_4183);
xnor U4236 (N_4236,N_4158,N_4113);
nor U4237 (N_4237,N_4120,N_4143);
nand U4238 (N_4238,N_4169,N_4122);
or U4239 (N_4239,N_4175,N_4153);
nand U4240 (N_4240,N_4127,N_4199);
or U4241 (N_4241,N_4150,N_4196);
or U4242 (N_4242,N_4198,N_4102);
or U4243 (N_4243,N_4106,N_4118);
nor U4244 (N_4244,N_4171,N_4179);
nor U4245 (N_4245,N_4124,N_4128);
xor U4246 (N_4246,N_4191,N_4111);
nor U4247 (N_4247,N_4104,N_4101);
nand U4248 (N_4248,N_4125,N_4163);
and U4249 (N_4249,N_4137,N_4132);
nor U4250 (N_4250,N_4125,N_4109);
nand U4251 (N_4251,N_4177,N_4163);
or U4252 (N_4252,N_4163,N_4119);
and U4253 (N_4253,N_4151,N_4172);
xnor U4254 (N_4254,N_4146,N_4178);
nand U4255 (N_4255,N_4117,N_4138);
nor U4256 (N_4256,N_4113,N_4103);
and U4257 (N_4257,N_4150,N_4130);
xnor U4258 (N_4258,N_4149,N_4172);
nor U4259 (N_4259,N_4130,N_4118);
xnor U4260 (N_4260,N_4178,N_4117);
or U4261 (N_4261,N_4150,N_4104);
xor U4262 (N_4262,N_4133,N_4171);
xnor U4263 (N_4263,N_4142,N_4126);
nor U4264 (N_4264,N_4194,N_4107);
xor U4265 (N_4265,N_4183,N_4111);
nor U4266 (N_4266,N_4175,N_4171);
nand U4267 (N_4267,N_4195,N_4149);
and U4268 (N_4268,N_4110,N_4117);
and U4269 (N_4269,N_4127,N_4143);
xnor U4270 (N_4270,N_4131,N_4174);
or U4271 (N_4271,N_4101,N_4189);
or U4272 (N_4272,N_4198,N_4157);
xnor U4273 (N_4273,N_4102,N_4105);
and U4274 (N_4274,N_4111,N_4161);
nor U4275 (N_4275,N_4134,N_4114);
xnor U4276 (N_4276,N_4158,N_4137);
xnor U4277 (N_4277,N_4178,N_4100);
xor U4278 (N_4278,N_4112,N_4151);
xnor U4279 (N_4279,N_4195,N_4199);
and U4280 (N_4280,N_4141,N_4147);
or U4281 (N_4281,N_4194,N_4141);
nand U4282 (N_4282,N_4178,N_4112);
or U4283 (N_4283,N_4197,N_4195);
nor U4284 (N_4284,N_4135,N_4153);
nor U4285 (N_4285,N_4189,N_4173);
xnor U4286 (N_4286,N_4172,N_4106);
nand U4287 (N_4287,N_4148,N_4126);
and U4288 (N_4288,N_4106,N_4168);
nand U4289 (N_4289,N_4116,N_4194);
xnor U4290 (N_4290,N_4122,N_4153);
xnor U4291 (N_4291,N_4188,N_4109);
and U4292 (N_4292,N_4162,N_4198);
xnor U4293 (N_4293,N_4190,N_4152);
nand U4294 (N_4294,N_4166,N_4170);
and U4295 (N_4295,N_4144,N_4147);
nand U4296 (N_4296,N_4189,N_4139);
nor U4297 (N_4297,N_4125,N_4191);
nor U4298 (N_4298,N_4120,N_4139);
xor U4299 (N_4299,N_4180,N_4146);
xnor U4300 (N_4300,N_4298,N_4247);
nor U4301 (N_4301,N_4256,N_4225);
nand U4302 (N_4302,N_4254,N_4296);
and U4303 (N_4303,N_4292,N_4294);
nor U4304 (N_4304,N_4235,N_4259);
and U4305 (N_4305,N_4211,N_4203);
or U4306 (N_4306,N_4228,N_4248);
xor U4307 (N_4307,N_4231,N_4282);
xor U4308 (N_4308,N_4205,N_4260);
or U4309 (N_4309,N_4265,N_4255);
nand U4310 (N_4310,N_4210,N_4213);
xnor U4311 (N_4311,N_4284,N_4241);
xnor U4312 (N_4312,N_4271,N_4237);
xor U4313 (N_4313,N_4251,N_4230);
or U4314 (N_4314,N_4246,N_4287);
xor U4315 (N_4315,N_4244,N_4233);
nor U4316 (N_4316,N_4278,N_4291);
nor U4317 (N_4317,N_4269,N_4249);
nor U4318 (N_4318,N_4268,N_4214);
or U4319 (N_4319,N_4238,N_4280);
or U4320 (N_4320,N_4200,N_4216);
nand U4321 (N_4321,N_4222,N_4275);
and U4322 (N_4322,N_4219,N_4234);
nand U4323 (N_4323,N_4283,N_4277);
and U4324 (N_4324,N_4242,N_4267);
or U4325 (N_4325,N_4295,N_4297);
xor U4326 (N_4326,N_4262,N_4286);
nand U4327 (N_4327,N_4202,N_4252);
and U4328 (N_4328,N_4243,N_4273);
nor U4329 (N_4329,N_4299,N_4204);
or U4330 (N_4330,N_4293,N_4274);
nor U4331 (N_4331,N_4288,N_4281);
xor U4332 (N_4332,N_4220,N_4272);
xor U4333 (N_4333,N_4253,N_4276);
xor U4334 (N_4334,N_4224,N_4245);
or U4335 (N_4335,N_4289,N_4217);
nor U4336 (N_4336,N_4290,N_4250);
xnor U4337 (N_4337,N_4212,N_4208);
and U4338 (N_4338,N_4264,N_4227);
nor U4339 (N_4339,N_4207,N_4206);
nand U4340 (N_4340,N_4215,N_4232);
nand U4341 (N_4341,N_4221,N_4236);
nand U4342 (N_4342,N_4240,N_4270);
or U4343 (N_4343,N_4258,N_4226);
xnor U4344 (N_4344,N_4285,N_4201);
nand U4345 (N_4345,N_4257,N_4279);
xnor U4346 (N_4346,N_4239,N_4261);
and U4347 (N_4347,N_4229,N_4218);
xor U4348 (N_4348,N_4209,N_4266);
or U4349 (N_4349,N_4223,N_4263);
or U4350 (N_4350,N_4258,N_4230);
nand U4351 (N_4351,N_4260,N_4290);
and U4352 (N_4352,N_4298,N_4204);
xnor U4353 (N_4353,N_4298,N_4279);
xor U4354 (N_4354,N_4283,N_4214);
nand U4355 (N_4355,N_4281,N_4230);
and U4356 (N_4356,N_4239,N_4228);
and U4357 (N_4357,N_4241,N_4270);
nor U4358 (N_4358,N_4276,N_4261);
xnor U4359 (N_4359,N_4227,N_4203);
or U4360 (N_4360,N_4268,N_4245);
nor U4361 (N_4361,N_4251,N_4272);
nor U4362 (N_4362,N_4213,N_4247);
and U4363 (N_4363,N_4272,N_4219);
or U4364 (N_4364,N_4253,N_4236);
and U4365 (N_4365,N_4214,N_4256);
nand U4366 (N_4366,N_4264,N_4217);
or U4367 (N_4367,N_4244,N_4203);
and U4368 (N_4368,N_4299,N_4268);
or U4369 (N_4369,N_4233,N_4299);
and U4370 (N_4370,N_4268,N_4201);
or U4371 (N_4371,N_4233,N_4295);
nand U4372 (N_4372,N_4273,N_4280);
nor U4373 (N_4373,N_4257,N_4242);
nand U4374 (N_4374,N_4208,N_4203);
nor U4375 (N_4375,N_4212,N_4214);
and U4376 (N_4376,N_4291,N_4223);
or U4377 (N_4377,N_4264,N_4288);
xnor U4378 (N_4378,N_4200,N_4240);
nor U4379 (N_4379,N_4227,N_4251);
nand U4380 (N_4380,N_4244,N_4222);
nand U4381 (N_4381,N_4299,N_4288);
nand U4382 (N_4382,N_4228,N_4299);
and U4383 (N_4383,N_4245,N_4216);
nor U4384 (N_4384,N_4257,N_4203);
and U4385 (N_4385,N_4289,N_4203);
nor U4386 (N_4386,N_4207,N_4278);
nand U4387 (N_4387,N_4241,N_4213);
or U4388 (N_4388,N_4289,N_4286);
or U4389 (N_4389,N_4249,N_4206);
nand U4390 (N_4390,N_4209,N_4202);
or U4391 (N_4391,N_4268,N_4266);
xnor U4392 (N_4392,N_4218,N_4230);
and U4393 (N_4393,N_4205,N_4214);
and U4394 (N_4394,N_4255,N_4205);
nand U4395 (N_4395,N_4248,N_4291);
and U4396 (N_4396,N_4264,N_4266);
and U4397 (N_4397,N_4215,N_4291);
or U4398 (N_4398,N_4212,N_4229);
and U4399 (N_4399,N_4227,N_4206);
nand U4400 (N_4400,N_4399,N_4382);
xnor U4401 (N_4401,N_4397,N_4392);
nand U4402 (N_4402,N_4334,N_4362);
nand U4403 (N_4403,N_4386,N_4394);
and U4404 (N_4404,N_4302,N_4389);
xnor U4405 (N_4405,N_4384,N_4304);
nor U4406 (N_4406,N_4328,N_4360);
and U4407 (N_4407,N_4314,N_4357);
nand U4408 (N_4408,N_4333,N_4310);
or U4409 (N_4409,N_4352,N_4371);
or U4410 (N_4410,N_4378,N_4396);
xor U4411 (N_4411,N_4367,N_4372);
nand U4412 (N_4412,N_4353,N_4376);
and U4413 (N_4413,N_4349,N_4391);
xnor U4414 (N_4414,N_4385,N_4377);
and U4415 (N_4415,N_4341,N_4317);
nand U4416 (N_4416,N_4373,N_4315);
nand U4417 (N_4417,N_4332,N_4346);
or U4418 (N_4418,N_4345,N_4356);
nand U4419 (N_4419,N_4313,N_4379);
or U4420 (N_4420,N_4324,N_4308);
or U4421 (N_4421,N_4330,N_4320);
xnor U4422 (N_4422,N_4388,N_4387);
xor U4423 (N_4423,N_4325,N_4369);
and U4424 (N_4424,N_4354,N_4300);
nand U4425 (N_4425,N_4351,N_4342);
xnor U4426 (N_4426,N_4339,N_4316);
nor U4427 (N_4427,N_4361,N_4327);
nand U4428 (N_4428,N_4395,N_4318);
nor U4429 (N_4429,N_4363,N_4309);
nor U4430 (N_4430,N_4337,N_4319);
xnor U4431 (N_4431,N_4303,N_4321);
xnor U4432 (N_4432,N_4383,N_4381);
nor U4433 (N_4433,N_4347,N_4390);
or U4434 (N_4434,N_4307,N_4370);
xnor U4435 (N_4435,N_4322,N_4323);
or U4436 (N_4436,N_4366,N_4358);
nor U4437 (N_4437,N_4368,N_4398);
and U4438 (N_4438,N_4301,N_4306);
and U4439 (N_4439,N_4338,N_4335);
or U4440 (N_4440,N_4329,N_4380);
nor U4441 (N_4441,N_4340,N_4331);
xnor U4442 (N_4442,N_4359,N_4393);
nor U4443 (N_4443,N_4326,N_4312);
or U4444 (N_4444,N_4365,N_4305);
nor U4445 (N_4445,N_4343,N_4311);
and U4446 (N_4446,N_4350,N_4355);
or U4447 (N_4447,N_4348,N_4364);
or U4448 (N_4448,N_4374,N_4344);
and U4449 (N_4449,N_4336,N_4375);
nor U4450 (N_4450,N_4365,N_4347);
and U4451 (N_4451,N_4325,N_4332);
xnor U4452 (N_4452,N_4344,N_4361);
or U4453 (N_4453,N_4368,N_4371);
or U4454 (N_4454,N_4344,N_4384);
or U4455 (N_4455,N_4398,N_4335);
or U4456 (N_4456,N_4323,N_4347);
nor U4457 (N_4457,N_4352,N_4384);
nand U4458 (N_4458,N_4384,N_4315);
or U4459 (N_4459,N_4337,N_4399);
nor U4460 (N_4460,N_4393,N_4352);
xor U4461 (N_4461,N_4372,N_4315);
or U4462 (N_4462,N_4330,N_4344);
and U4463 (N_4463,N_4302,N_4308);
nand U4464 (N_4464,N_4310,N_4354);
xnor U4465 (N_4465,N_4378,N_4343);
xor U4466 (N_4466,N_4302,N_4374);
nand U4467 (N_4467,N_4325,N_4311);
or U4468 (N_4468,N_4311,N_4381);
nor U4469 (N_4469,N_4333,N_4313);
or U4470 (N_4470,N_4388,N_4345);
nor U4471 (N_4471,N_4345,N_4332);
xnor U4472 (N_4472,N_4385,N_4371);
or U4473 (N_4473,N_4352,N_4323);
nand U4474 (N_4474,N_4387,N_4339);
xor U4475 (N_4475,N_4388,N_4303);
nor U4476 (N_4476,N_4394,N_4311);
and U4477 (N_4477,N_4368,N_4379);
or U4478 (N_4478,N_4363,N_4340);
nand U4479 (N_4479,N_4317,N_4343);
and U4480 (N_4480,N_4399,N_4371);
nor U4481 (N_4481,N_4382,N_4386);
nor U4482 (N_4482,N_4341,N_4392);
or U4483 (N_4483,N_4367,N_4321);
and U4484 (N_4484,N_4333,N_4365);
nor U4485 (N_4485,N_4392,N_4369);
nand U4486 (N_4486,N_4399,N_4340);
or U4487 (N_4487,N_4397,N_4372);
or U4488 (N_4488,N_4341,N_4352);
xnor U4489 (N_4489,N_4392,N_4344);
nor U4490 (N_4490,N_4369,N_4399);
and U4491 (N_4491,N_4327,N_4384);
or U4492 (N_4492,N_4353,N_4371);
and U4493 (N_4493,N_4373,N_4375);
and U4494 (N_4494,N_4364,N_4359);
and U4495 (N_4495,N_4327,N_4376);
or U4496 (N_4496,N_4354,N_4388);
nor U4497 (N_4497,N_4302,N_4358);
xnor U4498 (N_4498,N_4325,N_4309);
and U4499 (N_4499,N_4375,N_4364);
nor U4500 (N_4500,N_4421,N_4428);
nor U4501 (N_4501,N_4400,N_4426);
nand U4502 (N_4502,N_4496,N_4405);
nor U4503 (N_4503,N_4443,N_4475);
xor U4504 (N_4504,N_4422,N_4451);
or U4505 (N_4505,N_4457,N_4414);
nand U4506 (N_4506,N_4485,N_4476);
nand U4507 (N_4507,N_4441,N_4412);
nand U4508 (N_4508,N_4431,N_4455);
and U4509 (N_4509,N_4473,N_4493);
or U4510 (N_4510,N_4429,N_4470);
nand U4511 (N_4511,N_4456,N_4413);
and U4512 (N_4512,N_4445,N_4494);
or U4513 (N_4513,N_4497,N_4402);
nor U4514 (N_4514,N_4452,N_4425);
and U4515 (N_4515,N_4479,N_4480);
nor U4516 (N_4516,N_4407,N_4499);
xnor U4517 (N_4517,N_4465,N_4444);
and U4518 (N_4518,N_4477,N_4432);
nor U4519 (N_4519,N_4442,N_4435);
and U4520 (N_4520,N_4498,N_4427);
nor U4521 (N_4521,N_4446,N_4416);
and U4522 (N_4522,N_4478,N_4418);
nor U4523 (N_4523,N_4492,N_4491);
nand U4524 (N_4524,N_4450,N_4449);
nand U4525 (N_4525,N_4468,N_4462);
nand U4526 (N_4526,N_4409,N_4439);
nand U4527 (N_4527,N_4464,N_4423);
and U4528 (N_4528,N_4467,N_4460);
xnor U4529 (N_4529,N_4481,N_4483);
or U4530 (N_4530,N_4471,N_4434);
or U4531 (N_4531,N_4453,N_4472);
and U4532 (N_4532,N_4437,N_4404);
or U4533 (N_4533,N_4410,N_4474);
nor U4534 (N_4534,N_4401,N_4488);
and U4535 (N_4535,N_4461,N_4417);
or U4536 (N_4536,N_4411,N_4440);
nand U4537 (N_4537,N_4495,N_4424);
nand U4538 (N_4538,N_4419,N_4408);
or U4539 (N_4539,N_4436,N_4448);
and U4540 (N_4540,N_4466,N_4403);
and U4541 (N_4541,N_4447,N_4482);
nor U4542 (N_4542,N_4430,N_4454);
nand U4543 (N_4543,N_4438,N_4463);
nor U4544 (N_4544,N_4490,N_4458);
xnor U4545 (N_4545,N_4406,N_4486);
xnor U4546 (N_4546,N_4433,N_4487);
or U4547 (N_4547,N_4469,N_4489);
and U4548 (N_4548,N_4420,N_4459);
nor U4549 (N_4549,N_4415,N_4484);
and U4550 (N_4550,N_4426,N_4410);
nand U4551 (N_4551,N_4484,N_4475);
nor U4552 (N_4552,N_4471,N_4404);
and U4553 (N_4553,N_4400,N_4436);
or U4554 (N_4554,N_4495,N_4469);
xnor U4555 (N_4555,N_4446,N_4457);
nand U4556 (N_4556,N_4460,N_4483);
or U4557 (N_4557,N_4498,N_4478);
or U4558 (N_4558,N_4489,N_4463);
xor U4559 (N_4559,N_4426,N_4491);
nor U4560 (N_4560,N_4426,N_4424);
nand U4561 (N_4561,N_4452,N_4494);
nand U4562 (N_4562,N_4481,N_4453);
and U4563 (N_4563,N_4417,N_4469);
and U4564 (N_4564,N_4462,N_4446);
and U4565 (N_4565,N_4435,N_4463);
xor U4566 (N_4566,N_4424,N_4472);
nand U4567 (N_4567,N_4463,N_4421);
and U4568 (N_4568,N_4455,N_4405);
and U4569 (N_4569,N_4408,N_4455);
nand U4570 (N_4570,N_4401,N_4455);
nand U4571 (N_4571,N_4402,N_4484);
xnor U4572 (N_4572,N_4438,N_4402);
nor U4573 (N_4573,N_4492,N_4446);
nor U4574 (N_4574,N_4416,N_4431);
or U4575 (N_4575,N_4492,N_4439);
xor U4576 (N_4576,N_4401,N_4413);
xnor U4577 (N_4577,N_4460,N_4443);
nand U4578 (N_4578,N_4491,N_4460);
nand U4579 (N_4579,N_4460,N_4456);
nor U4580 (N_4580,N_4414,N_4441);
nand U4581 (N_4581,N_4437,N_4467);
nor U4582 (N_4582,N_4423,N_4438);
xor U4583 (N_4583,N_4426,N_4473);
or U4584 (N_4584,N_4464,N_4407);
xor U4585 (N_4585,N_4410,N_4446);
or U4586 (N_4586,N_4483,N_4480);
nor U4587 (N_4587,N_4437,N_4478);
and U4588 (N_4588,N_4469,N_4450);
nor U4589 (N_4589,N_4407,N_4403);
and U4590 (N_4590,N_4453,N_4443);
nor U4591 (N_4591,N_4479,N_4492);
xnor U4592 (N_4592,N_4478,N_4470);
nand U4593 (N_4593,N_4427,N_4475);
and U4594 (N_4594,N_4471,N_4450);
and U4595 (N_4595,N_4499,N_4447);
or U4596 (N_4596,N_4412,N_4431);
nand U4597 (N_4597,N_4444,N_4467);
nor U4598 (N_4598,N_4434,N_4422);
xor U4599 (N_4599,N_4435,N_4426);
nor U4600 (N_4600,N_4534,N_4529);
xnor U4601 (N_4601,N_4569,N_4542);
nor U4602 (N_4602,N_4530,N_4547);
and U4603 (N_4603,N_4531,N_4502);
and U4604 (N_4604,N_4535,N_4588);
and U4605 (N_4605,N_4571,N_4519);
xnor U4606 (N_4606,N_4532,N_4562);
nand U4607 (N_4607,N_4559,N_4503);
xnor U4608 (N_4608,N_4567,N_4574);
or U4609 (N_4609,N_4584,N_4554);
nand U4610 (N_4610,N_4596,N_4586);
nor U4611 (N_4611,N_4582,N_4512);
or U4612 (N_4612,N_4589,N_4594);
and U4613 (N_4613,N_4555,N_4515);
and U4614 (N_4614,N_4599,N_4557);
xor U4615 (N_4615,N_4551,N_4597);
or U4616 (N_4616,N_4598,N_4539);
nor U4617 (N_4617,N_4556,N_4509);
or U4618 (N_4618,N_4540,N_4505);
xor U4619 (N_4619,N_4507,N_4537);
or U4620 (N_4620,N_4544,N_4566);
nand U4621 (N_4621,N_4548,N_4501);
nor U4622 (N_4622,N_4518,N_4520);
and U4623 (N_4623,N_4521,N_4587);
xnor U4624 (N_4624,N_4591,N_4572);
nand U4625 (N_4625,N_4590,N_4527);
nand U4626 (N_4626,N_4583,N_4514);
nand U4627 (N_4627,N_4565,N_4549);
or U4628 (N_4628,N_4538,N_4593);
and U4629 (N_4629,N_4592,N_4504);
or U4630 (N_4630,N_4513,N_4550);
xor U4631 (N_4631,N_4546,N_4561);
nand U4632 (N_4632,N_4516,N_4552);
and U4633 (N_4633,N_4575,N_4536);
xor U4634 (N_4634,N_4508,N_4500);
or U4635 (N_4635,N_4580,N_4577);
nand U4636 (N_4636,N_4522,N_4564);
nor U4637 (N_4637,N_4506,N_4573);
nand U4638 (N_4638,N_4560,N_4524);
nor U4639 (N_4639,N_4543,N_4533);
or U4640 (N_4640,N_4510,N_4528);
or U4641 (N_4641,N_4558,N_4578);
xor U4642 (N_4642,N_4570,N_4526);
nand U4643 (N_4643,N_4568,N_4595);
nand U4644 (N_4644,N_4553,N_4579);
nand U4645 (N_4645,N_4545,N_4576);
nand U4646 (N_4646,N_4511,N_4517);
nand U4647 (N_4647,N_4581,N_4523);
nor U4648 (N_4648,N_4525,N_4585);
nand U4649 (N_4649,N_4541,N_4563);
nor U4650 (N_4650,N_4529,N_4524);
xnor U4651 (N_4651,N_4530,N_4545);
nand U4652 (N_4652,N_4533,N_4573);
xnor U4653 (N_4653,N_4593,N_4565);
nand U4654 (N_4654,N_4594,N_4598);
xor U4655 (N_4655,N_4596,N_4504);
or U4656 (N_4656,N_4533,N_4519);
xnor U4657 (N_4657,N_4505,N_4560);
and U4658 (N_4658,N_4549,N_4558);
nand U4659 (N_4659,N_4590,N_4557);
xnor U4660 (N_4660,N_4545,N_4562);
and U4661 (N_4661,N_4532,N_4585);
nor U4662 (N_4662,N_4520,N_4535);
and U4663 (N_4663,N_4597,N_4534);
xor U4664 (N_4664,N_4574,N_4588);
xor U4665 (N_4665,N_4580,N_4552);
nand U4666 (N_4666,N_4556,N_4576);
xor U4667 (N_4667,N_4581,N_4522);
and U4668 (N_4668,N_4520,N_4599);
nand U4669 (N_4669,N_4508,N_4595);
and U4670 (N_4670,N_4547,N_4536);
or U4671 (N_4671,N_4580,N_4526);
and U4672 (N_4672,N_4549,N_4593);
nand U4673 (N_4673,N_4513,N_4530);
xor U4674 (N_4674,N_4529,N_4560);
and U4675 (N_4675,N_4527,N_4519);
or U4676 (N_4676,N_4563,N_4514);
nor U4677 (N_4677,N_4586,N_4539);
xnor U4678 (N_4678,N_4547,N_4546);
xor U4679 (N_4679,N_4562,N_4533);
nand U4680 (N_4680,N_4531,N_4589);
xor U4681 (N_4681,N_4562,N_4535);
xor U4682 (N_4682,N_4598,N_4550);
xnor U4683 (N_4683,N_4579,N_4545);
nor U4684 (N_4684,N_4574,N_4503);
xor U4685 (N_4685,N_4534,N_4501);
xor U4686 (N_4686,N_4575,N_4547);
nand U4687 (N_4687,N_4561,N_4542);
or U4688 (N_4688,N_4570,N_4517);
nand U4689 (N_4689,N_4540,N_4594);
xor U4690 (N_4690,N_4534,N_4554);
or U4691 (N_4691,N_4543,N_4529);
and U4692 (N_4692,N_4564,N_4568);
xor U4693 (N_4693,N_4532,N_4595);
and U4694 (N_4694,N_4533,N_4528);
nor U4695 (N_4695,N_4599,N_4507);
nand U4696 (N_4696,N_4543,N_4535);
nand U4697 (N_4697,N_4585,N_4542);
or U4698 (N_4698,N_4515,N_4582);
and U4699 (N_4699,N_4530,N_4540);
and U4700 (N_4700,N_4637,N_4616);
xor U4701 (N_4701,N_4643,N_4681);
and U4702 (N_4702,N_4673,N_4697);
xnor U4703 (N_4703,N_4610,N_4683);
xnor U4704 (N_4704,N_4630,N_4600);
or U4705 (N_4705,N_4639,N_4680);
nor U4706 (N_4706,N_4664,N_4641);
nand U4707 (N_4707,N_4679,N_4677);
and U4708 (N_4708,N_4621,N_4696);
and U4709 (N_4709,N_4634,N_4650);
or U4710 (N_4710,N_4688,N_4635);
or U4711 (N_4711,N_4676,N_4661);
nor U4712 (N_4712,N_4628,N_4686);
and U4713 (N_4713,N_4606,N_4694);
xor U4714 (N_4714,N_4674,N_4655);
and U4715 (N_4715,N_4605,N_4658);
or U4716 (N_4716,N_4678,N_4645);
nand U4717 (N_4717,N_4654,N_4648);
nor U4718 (N_4718,N_4690,N_4636);
or U4719 (N_4719,N_4602,N_4623);
or U4720 (N_4720,N_4624,N_4663);
or U4721 (N_4721,N_4659,N_4604);
and U4722 (N_4722,N_4699,N_4662);
and U4723 (N_4723,N_4622,N_4614);
nand U4724 (N_4724,N_4617,N_4631);
or U4725 (N_4725,N_4692,N_4633);
xnor U4726 (N_4726,N_4649,N_4612);
and U4727 (N_4727,N_4651,N_4611);
and U4728 (N_4728,N_4665,N_4618);
nor U4729 (N_4729,N_4670,N_4625);
and U4730 (N_4730,N_4669,N_4619);
or U4731 (N_4731,N_4620,N_4672);
or U4732 (N_4732,N_4685,N_4693);
or U4733 (N_4733,N_4629,N_4608);
or U4734 (N_4734,N_4627,N_4647);
and U4735 (N_4735,N_4646,N_4640);
nor U4736 (N_4736,N_4603,N_4684);
nor U4737 (N_4737,N_4644,N_4660);
xor U4738 (N_4738,N_4638,N_4698);
xnor U4739 (N_4739,N_4607,N_4613);
or U4740 (N_4740,N_4615,N_4695);
xor U4741 (N_4741,N_4653,N_4682);
and U4742 (N_4742,N_4667,N_4668);
xor U4743 (N_4743,N_4657,N_4652);
xnor U4744 (N_4744,N_4689,N_4656);
and U4745 (N_4745,N_4632,N_4626);
and U4746 (N_4746,N_4609,N_4666);
nor U4747 (N_4747,N_4691,N_4687);
or U4748 (N_4748,N_4671,N_4675);
nor U4749 (N_4749,N_4601,N_4642);
xnor U4750 (N_4750,N_4626,N_4623);
and U4751 (N_4751,N_4619,N_4615);
nand U4752 (N_4752,N_4698,N_4610);
xor U4753 (N_4753,N_4605,N_4602);
nor U4754 (N_4754,N_4687,N_4620);
nand U4755 (N_4755,N_4602,N_4688);
or U4756 (N_4756,N_4651,N_4661);
nor U4757 (N_4757,N_4623,N_4622);
nor U4758 (N_4758,N_4692,N_4652);
xor U4759 (N_4759,N_4698,N_4637);
nand U4760 (N_4760,N_4627,N_4675);
xnor U4761 (N_4761,N_4664,N_4646);
and U4762 (N_4762,N_4612,N_4650);
nand U4763 (N_4763,N_4623,N_4662);
xnor U4764 (N_4764,N_4662,N_4663);
nor U4765 (N_4765,N_4625,N_4685);
xor U4766 (N_4766,N_4672,N_4668);
xor U4767 (N_4767,N_4680,N_4683);
xnor U4768 (N_4768,N_4667,N_4695);
and U4769 (N_4769,N_4683,N_4686);
xor U4770 (N_4770,N_4669,N_4617);
nor U4771 (N_4771,N_4637,N_4614);
or U4772 (N_4772,N_4665,N_4650);
and U4773 (N_4773,N_4645,N_4698);
nand U4774 (N_4774,N_4611,N_4629);
and U4775 (N_4775,N_4643,N_4667);
nor U4776 (N_4776,N_4611,N_4668);
nand U4777 (N_4777,N_4629,N_4631);
xnor U4778 (N_4778,N_4691,N_4619);
and U4779 (N_4779,N_4667,N_4604);
xor U4780 (N_4780,N_4638,N_4667);
nor U4781 (N_4781,N_4624,N_4646);
or U4782 (N_4782,N_4663,N_4685);
or U4783 (N_4783,N_4635,N_4606);
nor U4784 (N_4784,N_4637,N_4660);
and U4785 (N_4785,N_4674,N_4688);
xor U4786 (N_4786,N_4688,N_4643);
and U4787 (N_4787,N_4651,N_4662);
nor U4788 (N_4788,N_4619,N_4672);
nand U4789 (N_4789,N_4673,N_4605);
nor U4790 (N_4790,N_4632,N_4695);
nor U4791 (N_4791,N_4605,N_4685);
xnor U4792 (N_4792,N_4653,N_4600);
xnor U4793 (N_4793,N_4645,N_4658);
xor U4794 (N_4794,N_4645,N_4653);
nand U4795 (N_4795,N_4641,N_4653);
and U4796 (N_4796,N_4689,N_4608);
xnor U4797 (N_4797,N_4610,N_4625);
xnor U4798 (N_4798,N_4635,N_4659);
nor U4799 (N_4799,N_4655,N_4616);
nand U4800 (N_4800,N_4728,N_4712);
or U4801 (N_4801,N_4772,N_4770);
xor U4802 (N_4802,N_4727,N_4701);
or U4803 (N_4803,N_4721,N_4738);
xnor U4804 (N_4804,N_4799,N_4763);
nor U4805 (N_4805,N_4777,N_4754);
nor U4806 (N_4806,N_4761,N_4776);
xnor U4807 (N_4807,N_4756,N_4765);
and U4808 (N_4808,N_4719,N_4704);
xor U4809 (N_4809,N_4710,N_4767);
nand U4810 (N_4810,N_4771,N_4709);
and U4811 (N_4811,N_4794,N_4706);
nand U4812 (N_4812,N_4781,N_4746);
and U4813 (N_4813,N_4720,N_4736);
or U4814 (N_4814,N_4755,N_4744);
xor U4815 (N_4815,N_4766,N_4733);
and U4816 (N_4816,N_4786,N_4737);
or U4817 (N_4817,N_4768,N_4792);
and U4818 (N_4818,N_4787,N_4796);
and U4819 (N_4819,N_4743,N_4739);
and U4820 (N_4820,N_4708,N_4785);
or U4821 (N_4821,N_4747,N_4769);
and U4822 (N_4822,N_4780,N_4742);
xor U4823 (N_4823,N_4791,N_4764);
or U4824 (N_4824,N_4758,N_4723);
and U4825 (N_4825,N_4741,N_4749);
nand U4826 (N_4826,N_4762,N_4711);
xnor U4827 (N_4827,N_4788,N_4734);
xor U4828 (N_4828,N_4798,N_4782);
and U4829 (N_4829,N_4774,N_4773);
or U4830 (N_4830,N_4797,N_4789);
and U4831 (N_4831,N_4750,N_4730);
xor U4832 (N_4832,N_4700,N_4795);
nor U4833 (N_4833,N_4790,N_4783);
and U4834 (N_4834,N_4724,N_4775);
nor U4835 (N_4835,N_4705,N_4725);
nand U4836 (N_4836,N_4760,N_4703);
nand U4837 (N_4837,N_4726,N_4716);
xor U4838 (N_4838,N_4793,N_4759);
nand U4839 (N_4839,N_4715,N_4748);
xnor U4840 (N_4840,N_4784,N_4740);
nand U4841 (N_4841,N_4702,N_4757);
xnor U4842 (N_4842,N_4717,N_4729);
and U4843 (N_4843,N_4752,N_4731);
nand U4844 (N_4844,N_4735,N_4707);
xnor U4845 (N_4845,N_4718,N_4779);
nand U4846 (N_4846,N_4778,N_4722);
nor U4847 (N_4847,N_4714,N_4751);
or U4848 (N_4848,N_4732,N_4713);
xor U4849 (N_4849,N_4753,N_4745);
and U4850 (N_4850,N_4766,N_4736);
nand U4851 (N_4851,N_4765,N_4791);
and U4852 (N_4852,N_4751,N_4735);
nor U4853 (N_4853,N_4796,N_4788);
and U4854 (N_4854,N_4734,N_4711);
or U4855 (N_4855,N_4702,N_4776);
or U4856 (N_4856,N_4718,N_4787);
nor U4857 (N_4857,N_4714,N_4767);
or U4858 (N_4858,N_4715,N_4704);
or U4859 (N_4859,N_4714,N_4754);
nand U4860 (N_4860,N_4788,N_4785);
nand U4861 (N_4861,N_4775,N_4741);
and U4862 (N_4862,N_4794,N_4757);
or U4863 (N_4863,N_4750,N_4721);
and U4864 (N_4864,N_4735,N_4785);
or U4865 (N_4865,N_4700,N_4737);
and U4866 (N_4866,N_4721,N_4764);
xor U4867 (N_4867,N_4717,N_4724);
or U4868 (N_4868,N_4794,N_4723);
nand U4869 (N_4869,N_4764,N_4794);
and U4870 (N_4870,N_4777,N_4769);
xnor U4871 (N_4871,N_4770,N_4771);
or U4872 (N_4872,N_4720,N_4724);
or U4873 (N_4873,N_4750,N_4746);
nand U4874 (N_4874,N_4739,N_4735);
or U4875 (N_4875,N_4731,N_4764);
or U4876 (N_4876,N_4704,N_4772);
or U4877 (N_4877,N_4730,N_4773);
nand U4878 (N_4878,N_4713,N_4720);
xnor U4879 (N_4879,N_4769,N_4798);
nor U4880 (N_4880,N_4700,N_4753);
and U4881 (N_4881,N_4726,N_4710);
nor U4882 (N_4882,N_4764,N_4744);
or U4883 (N_4883,N_4716,N_4746);
nor U4884 (N_4884,N_4791,N_4730);
xor U4885 (N_4885,N_4702,N_4724);
or U4886 (N_4886,N_4730,N_4716);
xnor U4887 (N_4887,N_4745,N_4744);
or U4888 (N_4888,N_4739,N_4736);
and U4889 (N_4889,N_4758,N_4713);
nand U4890 (N_4890,N_4736,N_4706);
nand U4891 (N_4891,N_4738,N_4723);
or U4892 (N_4892,N_4783,N_4767);
nand U4893 (N_4893,N_4745,N_4708);
xnor U4894 (N_4894,N_4701,N_4720);
or U4895 (N_4895,N_4713,N_4709);
or U4896 (N_4896,N_4770,N_4769);
and U4897 (N_4897,N_4718,N_4701);
and U4898 (N_4898,N_4727,N_4774);
xnor U4899 (N_4899,N_4709,N_4784);
xnor U4900 (N_4900,N_4835,N_4883);
and U4901 (N_4901,N_4879,N_4800);
nor U4902 (N_4902,N_4896,N_4876);
xor U4903 (N_4903,N_4836,N_4801);
nor U4904 (N_4904,N_4814,N_4869);
and U4905 (N_4905,N_4893,N_4823);
and U4906 (N_4906,N_4887,N_4899);
nor U4907 (N_4907,N_4813,N_4855);
or U4908 (N_4908,N_4840,N_4810);
and U4909 (N_4909,N_4870,N_4812);
xnor U4910 (N_4910,N_4862,N_4880);
xnor U4911 (N_4911,N_4820,N_4839);
or U4912 (N_4912,N_4856,N_4828);
and U4913 (N_4913,N_4849,N_4817);
nand U4914 (N_4914,N_4873,N_4838);
nand U4915 (N_4915,N_4807,N_4891);
and U4916 (N_4916,N_4890,N_4809);
nand U4917 (N_4917,N_4844,N_4898);
and U4918 (N_4918,N_4845,N_4832);
or U4919 (N_4919,N_4819,N_4818);
nor U4920 (N_4920,N_4826,N_4874);
xor U4921 (N_4921,N_4853,N_4863);
and U4922 (N_4922,N_4829,N_4857);
xnor U4923 (N_4923,N_4847,N_4867);
nand U4924 (N_4924,N_4894,N_4827);
or U4925 (N_4925,N_4802,N_4866);
nor U4926 (N_4926,N_4861,N_4831);
nor U4927 (N_4927,N_4804,N_4884);
xor U4928 (N_4928,N_4878,N_4882);
and U4929 (N_4929,N_4875,N_4850);
xor U4930 (N_4930,N_4892,N_4825);
and U4931 (N_4931,N_4868,N_4822);
xnor U4932 (N_4932,N_4834,N_4842);
and U4933 (N_4933,N_4803,N_4841);
xor U4934 (N_4934,N_4877,N_4888);
nand U4935 (N_4935,N_4886,N_4889);
nand U4936 (N_4936,N_4897,N_4806);
nand U4937 (N_4937,N_4895,N_4881);
xor U4938 (N_4938,N_4852,N_4864);
nand U4939 (N_4939,N_4808,N_4815);
and U4940 (N_4940,N_4830,N_4824);
xor U4941 (N_4941,N_4860,N_4837);
or U4942 (N_4942,N_4843,N_4858);
xor U4943 (N_4943,N_4854,N_4821);
nand U4944 (N_4944,N_4816,N_4885);
or U4945 (N_4945,N_4848,N_4851);
or U4946 (N_4946,N_4871,N_4805);
nor U4947 (N_4947,N_4865,N_4833);
nor U4948 (N_4948,N_4811,N_4859);
nor U4949 (N_4949,N_4872,N_4846);
or U4950 (N_4950,N_4826,N_4894);
nand U4951 (N_4951,N_4851,N_4887);
nand U4952 (N_4952,N_4824,N_4890);
nand U4953 (N_4953,N_4827,N_4888);
xnor U4954 (N_4954,N_4817,N_4868);
or U4955 (N_4955,N_4871,N_4878);
and U4956 (N_4956,N_4858,N_4837);
nand U4957 (N_4957,N_4875,N_4811);
xor U4958 (N_4958,N_4826,N_4865);
xor U4959 (N_4959,N_4857,N_4813);
or U4960 (N_4960,N_4897,N_4880);
or U4961 (N_4961,N_4848,N_4801);
and U4962 (N_4962,N_4829,N_4867);
and U4963 (N_4963,N_4868,N_4838);
nand U4964 (N_4964,N_4809,N_4817);
and U4965 (N_4965,N_4887,N_4876);
nand U4966 (N_4966,N_4866,N_4814);
nor U4967 (N_4967,N_4849,N_4889);
and U4968 (N_4968,N_4802,N_4820);
xor U4969 (N_4969,N_4851,N_4853);
and U4970 (N_4970,N_4840,N_4828);
or U4971 (N_4971,N_4809,N_4878);
and U4972 (N_4972,N_4852,N_4838);
nand U4973 (N_4973,N_4891,N_4852);
or U4974 (N_4974,N_4887,N_4866);
or U4975 (N_4975,N_4880,N_4867);
nor U4976 (N_4976,N_4844,N_4861);
nor U4977 (N_4977,N_4821,N_4896);
nor U4978 (N_4978,N_4800,N_4885);
and U4979 (N_4979,N_4826,N_4809);
and U4980 (N_4980,N_4847,N_4846);
or U4981 (N_4981,N_4805,N_4883);
or U4982 (N_4982,N_4819,N_4862);
xor U4983 (N_4983,N_4866,N_4811);
nand U4984 (N_4984,N_4857,N_4865);
and U4985 (N_4985,N_4894,N_4882);
xor U4986 (N_4986,N_4826,N_4851);
or U4987 (N_4987,N_4880,N_4839);
nand U4988 (N_4988,N_4863,N_4852);
nor U4989 (N_4989,N_4802,N_4876);
nor U4990 (N_4990,N_4888,N_4868);
or U4991 (N_4991,N_4834,N_4833);
xnor U4992 (N_4992,N_4838,N_4893);
nor U4993 (N_4993,N_4848,N_4871);
xor U4994 (N_4994,N_4833,N_4887);
nand U4995 (N_4995,N_4819,N_4864);
or U4996 (N_4996,N_4823,N_4832);
or U4997 (N_4997,N_4865,N_4839);
xor U4998 (N_4998,N_4889,N_4852);
or U4999 (N_4999,N_4876,N_4817);
nand UO_0 (O_0,N_4910,N_4943);
or UO_1 (O_1,N_4906,N_4962);
nand UO_2 (O_2,N_4963,N_4969);
nand UO_3 (O_3,N_4980,N_4995);
nand UO_4 (O_4,N_4998,N_4970);
and UO_5 (O_5,N_4994,N_4948);
xnor UO_6 (O_6,N_4939,N_4964);
and UO_7 (O_7,N_4988,N_4984);
or UO_8 (O_8,N_4904,N_4940);
and UO_9 (O_9,N_4932,N_4934);
nand UO_10 (O_10,N_4944,N_4954);
nor UO_11 (O_11,N_4938,N_4945);
nor UO_12 (O_12,N_4991,N_4999);
or UO_13 (O_13,N_4900,N_4976);
xnor UO_14 (O_14,N_4979,N_4966);
xnor UO_15 (O_15,N_4931,N_4975);
xor UO_16 (O_16,N_4981,N_4930);
nor UO_17 (O_17,N_4937,N_4909);
xnor UO_18 (O_18,N_4918,N_4953);
xor UO_19 (O_19,N_4901,N_4917);
nand UO_20 (O_20,N_4986,N_4926);
nand UO_21 (O_21,N_4974,N_4983);
nand UO_22 (O_22,N_4946,N_4957);
or UO_23 (O_23,N_4989,N_4961);
xor UO_24 (O_24,N_4990,N_4915);
and UO_25 (O_25,N_4982,N_4914);
or UO_26 (O_26,N_4920,N_4960);
xnor UO_27 (O_27,N_4923,N_4958);
or UO_28 (O_28,N_4959,N_4922);
or UO_29 (O_29,N_4967,N_4933);
or UO_30 (O_30,N_4992,N_4965);
nand UO_31 (O_31,N_4955,N_4908);
and UO_32 (O_32,N_4993,N_4942);
nand UO_33 (O_33,N_4925,N_4985);
xnor UO_34 (O_34,N_4949,N_4972);
or UO_35 (O_35,N_4935,N_4977);
nor UO_36 (O_36,N_4996,N_4950);
nand UO_37 (O_37,N_4978,N_4916);
and UO_38 (O_38,N_4951,N_4905);
xnor UO_39 (O_39,N_4952,N_4936);
and UO_40 (O_40,N_4997,N_4902);
nand UO_41 (O_41,N_4912,N_4956);
nand UO_42 (O_42,N_4911,N_4924);
nor UO_43 (O_43,N_4941,N_4913);
nand UO_44 (O_44,N_4919,N_4987);
or UO_45 (O_45,N_4921,N_4927);
and UO_46 (O_46,N_4947,N_4903);
xor UO_47 (O_47,N_4971,N_4928);
or UO_48 (O_48,N_4929,N_4907);
or UO_49 (O_49,N_4968,N_4973);
or UO_50 (O_50,N_4958,N_4943);
xor UO_51 (O_51,N_4949,N_4956);
nand UO_52 (O_52,N_4929,N_4945);
or UO_53 (O_53,N_4922,N_4917);
nor UO_54 (O_54,N_4908,N_4927);
nand UO_55 (O_55,N_4908,N_4946);
nand UO_56 (O_56,N_4997,N_4916);
nand UO_57 (O_57,N_4997,N_4975);
and UO_58 (O_58,N_4967,N_4927);
or UO_59 (O_59,N_4901,N_4996);
and UO_60 (O_60,N_4998,N_4954);
or UO_61 (O_61,N_4975,N_4900);
nand UO_62 (O_62,N_4900,N_4952);
and UO_63 (O_63,N_4902,N_4905);
nand UO_64 (O_64,N_4910,N_4964);
nand UO_65 (O_65,N_4934,N_4993);
nor UO_66 (O_66,N_4909,N_4927);
xor UO_67 (O_67,N_4981,N_4959);
xor UO_68 (O_68,N_4935,N_4985);
or UO_69 (O_69,N_4980,N_4929);
xnor UO_70 (O_70,N_4968,N_4946);
nand UO_71 (O_71,N_4903,N_4978);
or UO_72 (O_72,N_4965,N_4956);
and UO_73 (O_73,N_4914,N_4919);
or UO_74 (O_74,N_4965,N_4918);
nor UO_75 (O_75,N_4993,N_4950);
nand UO_76 (O_76,N_4951,N_4965);
nand UO_77 (O_77,N_4923,N_4953);
and UO_78 (O_78,N_4961,N_4942);
xor UO_79 (O_79,N_4993,N_4918);
or UO_80 (O_80,N_4913,N_4975);
nand UO_81 (O_81,N_4913,N_4925);
nand UO_82 (O_82,N_4960,N_4987);
nor UO_83 (O_83,N_4903,N_4929);
nor UO_84 (O_84,N_4996,N_4932);
nor UO_85 (O_85,N_4961,N_4974);
or UO_86 (O_86,N_4948,N_4944);
nor UO_87 (O_87,N_4943,N_4934);
nor UO_88 (O_88,N_4948,N_4901);
nor UO_89 (O_89,N_4944,N_4989);
nor UO_90 (O_90,N_4937,N_4968);
or UO_91 (O_91,N_4958,N_4966);
nor UO_92 (O_92,N_4934,N_4958);
nor UO_93 (O_93,N_4977,N_4920);
xnor UO_94 (O_94,N_4971,N_4913);
nor UO_95 (O_95,N_4911,N_4985);
xnor UO_96 (O_96,N_4918,N_4968);
and UO_97 (O_97,N_4962,N_4964);
or UO_98 (O_98,N_4926,N_4991);
xor UO_99 (O_99,N_4935,N_4950);
nand UO_100 (O_100,N_4900,N_4931);
nor UO_101 (O_101,N_4999,N_4993);
xor UO_102 (O_102,N_4939,N_4945);
nor UO_103 (O_103,N_4997,N_4981);
nor UO_104 (O_104,N_4960,N_4916);
or UO_105 (O_105,N_4980,N_4951);
nand UO_106 (O_106,N_4976,N_4996);
nor UO_107 (O_107,N_4961,N_4971);
and UO_108 (O_108,N_4924,N_4962);
and UO_109 (O_109,N_4996,N_4965);
and UO_110 (O_110,N_4968,N_4912);
xor UO_111 (O_111,N_4927,N_4905);
nand UO_112 (O_112,N_4941,N_4998);
or UO_113 (O_113,N_4997,N_4924);
and UO_114 (O_114,N_4962,N_4972);
and UO_115 (O_115,N_4930,N_4903);
nor UO_116 (O_116,N_4915,N_4948);
xor UO_117 (O_117,N_4947,N_4951);
or UO_118 (O_118,N_4965,N_4947);
or UO_119 (O_119,N_4918,N_4913);
nand UO_120 (O_120,N_4973,N_4950);
nor UO_121 (O_121,N_4918,N_4998);
or UO_122 (O_122,N_4991,N_4912);
nand UO_123 (O_123,N_4938,N_4982);
and UO_124 (O_124,N_4929,N_4947);
and UO_125 (O_125,N_4999,N_4931);
and UO_126 (O_126,N_4921,N_4932);
or UO_127 (O_127,N_4973,N_4966);
or UO_128 (O_128,N_4982,N_4947);
xor UO_129 (O_129,N_4948,N_4909);
nor UO_130 (O_130,N_4903,N_4925);
nor UO_131 (O_131,N_4900,N_4948);
and UO_132 (O_132,N_4958,N_4974);
nor UO_133 (O_133,N_4940,N_4951);
nor UO_134 (O_134,N_4909,N_4951);
nor UO_135 (O_135,N_4945,N_4908);
and UO_136 (O_136,N_4945,N_4953);
nand UO_137 (O_137,N_4950,N_4924);
xnor UO_138 (O_138,N_4901,N_4974);
xnor UO_139 (O_139,N_4910,N_4946);
nor UO_140 (O_140,N_4985,N_4987);
nand UO_141 (O_141,N_4974,N_4992);
xnor UO_142 (O_142,N_4946,N_4954);
and UO_143 (O_143,N_4998,N_4990);
and UO_144 (O_144,N_4919,N_4966);
nand UO_145 (O_145,N_4982,N_4944);
and UO_146 (O_146,N_4944,N_4932);
nand UO_147 (O_147,N_4908,N_4991);
and UO_148 (O_148,N_4935,N_4922);
nand UO_149 (O_149,N_4920,N_4990);
xnor UO_150 (O_150,N_4954,N_4929);
and UO_151 (O_151,N_4922,N_4907);
xor UO_152 (O_152,N_4936,N_4909);
nand UO_153 (O_153,N_4998,N_4983);
or UO_154 (O_154,N_4909,N_4900);
nand UO_155 (O_155,N_4927,N_4932);
nor UO_156 (O_156,N_4990,N_4911);
or UO_157 (O_157,N_4994,N_4992);
or UO_158 (O_158,N_4917,N_4914);
and UO_159 (O_159,N_4992,N_4922);
nand UO_160 (O_160,N_4954,N_4919);
xor UO_161 (O_161,N_4968,N_4910);
or UO_162 (O_162,N_4937,N_4990);
nand UO_163 (O_163,N_4964,N_4932);
nand UO_164 (O_164,N_4938,N_4998);
nand UO_165 (O_165,N_4939,N_4996);
nor UO_166 (O_166,N_4986,N_4954);
or UO_167 (O_167,N_4918,N_4982);
and UO_168 (O_168,N_4942,N_4979);
xor UO_169 (O_169,N_4959,N_4975);
or UO_170 (O_170,N_4967,N_4966);
and UO_171 (O_171,N_4977,N_4979);
or UO_172 (O_172,N_4989,N_4996);
xnor UO_173 (O_173,N_4906,N_4908);
nor UO_174 (O_174,N_4988,N_4929);
nand UO_175 (O_175,N_4923,N_4950);
nand UO_176 (O_176,N_4976,N_4994);
nand UO_177 (O_177,N_4974,N_4967);
nor UO_178 (O_178,N_4906,N_4919);
or UO_179 (O_179,N_4951,N_4989);
xor UO_180 (O_180,N_4998,N_4930);
xor UO_181 (O_181,N_4991,N_4979);
nor UO_182 (O_182,N_4960,N_4904);
nor UO_183 (O_183,N_4990,N_4924);
xor UO_184 (O_184,N_4942,N_4998);
nand UO_185 (O_185,N_4942,N_4932);
and UO_186 (O_186,N_4909,N_4999);
nor UO_187 (O_187,N_4959,N_4937);
nand UO_188 (O_188,N_4922,N_4963);
or UO_189 (O_189,N_4996,N_4991);
nor UO_190 (O_190,N_4922,N_4931);
nor UO_191 (O_191,N_4927,N_4930);
nor UO_192 (O_192,N_4929,N_4981);
or UO_193 (O_193,N_4969,N_4952);
nand UO_194 (O_194,N_4943,N_4993);
nand UO_195 (O_195,N_4977,N_4985);
nand UO_196 (O_196,N_4904,N_4924);
or UO_197 (O_197,N_4977,N_4997);
nand UO_198 (O_198,N_4912,N_4970);
nor UO_199 (O_199,N_4940,N_4921);
nand UO_200 (O_200,N_4979,N_4957);
xnor UO_201 (O_201,N_4963,N_4949);
nor UO_202 (O_202,N_4989,N_4974);
xor UO_203 (O_203,N_4946,N_4905);
or UO_204 (O_204,N_4907,N_4941);
nor UO_205 (O_205,N_4987,N_4926);
xnor UO_206 (O_206,N_4960,N_4941);
nor UO_207 (O_207,N_4906,N_4939);
or UO_208 (O_208,N_4923,N_4948);
and UO_209 (O_209,N_4911,N_4947);
or UO_210 (O_210,N_4932,N_4998);
nand UO_211 (O_211,N_4916,N_4945);
nand UO_212 (O_212,N_4961,N_4958);
xor UO_213 (O_213,N_4963,N_4967);
and UO_214 (O_214,N_4922,N_4911);
or UO_215 (O_215,N_4942,N_4917);
xor UO_216 (O_216,N_4920,N_4963);
xnor UO_217 (O_217,N_4918,N_4920);
xnor UO_218 (O_218,N_4969,N_4908);
and UO_219 (O_219,N_4947,N_4986);
or UO_220 (O_220,N_4902,N_4926);
nor UO_221 (O_221,N_4941,N_4943);
nand UO_222 (O_222,N_4990,N_4994);
or UO_223 (O_223,N_4974,N_4937);
and UO_224 (O_224,N_4995,N_4966);
nor UO_225 (O_225,N_4915,N_4926);
nand UO_226 (O_226,N_4902,N_4979);
and UO_227 (O_227,N_4996,N_4975);
and UO_228 (O_228,N_4932,N_4967);
xnor UO_229 (O_229,N_4969,N_4970);
xor UO_230 (O_230,N_4901,N_4934);
nand UO_231 (O_231,N_4963,N_4930);
and UO_232 (O_232,N_4930,N_4989);
and UO_233 (O_233,N_4975,N_4983);
xnor UO_234 (O_234,N_4901,N_4918);
nand UO_235 (O_235,N_4984,N_4993);
and UO_236 (O_236,N_4907,N_4972);
and UO_237 (O_237,N_4980,N_4993);
nand UO_238 (O_238,N_4960,N_4980);
and UO_239 (O_239,N_4930,N_4906);
or UO_240 (O_240,N_4927,N_4929);
nand UO_241 (O_241,N_4960,N_4953);
or UO_242 (O_242,N_4969,N_4932);
nor UO_243 (O_243,N_4915,N_4979);
xor UO_244 (O_244,N_4906,N_4924);
and UO_245 (O_245,N_4977,N_4992);
xor UO_246 (O_246,N_4998,N_4940);
nand UO_247 (O_247,N_4989,N_4945);
or UO_248 (O_248,N_4929,N_4908);
and UO_249 (O_249,N_4971,N_4914);
and UO_250 (O_250,N_4917,N_4996);
nand UO_251 (O_251,N_4954,N_4928);
nor UO_252 (O_252,N_4946,N_4928);
or UO_253 (O_253,N_4979,N_4992);
nor UO_254 (O_254,N_4984,N_4974);
nor UO_255 (O_255,N_4912,N_4992);
or UO_256 (O_256,N_4922,N_4927);
and UO_257 (O_257,N_4931,N_4929);
nand UO_258 (O_258,N_4999,N_4992);
xnor UO_259 (O_259,N_4947,N_4932);
xor UO_260 (O_260,N_4922,N_4980);
and UO_261 (O_261,N_4999,N_4959);
and UO_262 (O_262,N_4938,N_4946);
xor UO_263 (O_263,N_4997,N_4983);
or UO_264 (O_264,N_4975,N_4923);
or UO_265 (O_265,N_4965,N_4983);
and UO_266 (O_266,N_4947,N_4978);
and UO_267 (O_267,N_4976,N_4919);
or UO_268 (O_268,N_4959,N_4954);
nand UO_269 (O_269,N_4900,N_4964);
or UO_270 (O_270,N_4980,N_4973);
xnor UO_271 (O_271,N_4978,N_4992);
or UO_272 (O_272,N_4953,N_4935);
nor UO_273 (O_273,N_4970,N_4973);
and UO_274 (O_274,N_4974,N_4912);
nand UO_275 (O_275,N_4998,N_4994);
nor UO_276 (O_276,N_4947,N_4930);
xor UO_277 (O_277,N_4923,N_4952);
xnor UO_278 (O_278,N_4984,N_4991);
and UO_279 (O_279,N_4995,N_4949);
nor UO_280 (O_280,N_4928,N_4963);
xnor UO_281 (O_281,N_4955,N_4925);
nand UO_282 (O_282,N_4945,N_4998);
or UO_283 (O_283,N_4962,N_4993);
xor UO_284 (O_284,N_4975,N_4999);
nor UO_285 (O_285,N_4929,N_4970);
and UO_286 (O_286,N_4969,N_4916);
or UO_287 (O_287,N_4966,N_4916);
nand UO_288 (O_288,N_4941,N_4915);
and UO_289 (O_289,N_4944,N_4947);
nand UO_290 (O_290,N_4959,N_4942);
nor UO_291 (O_291,N_4987,N_4996);
xnor UO_292 (O_292,N_4916,N_4943);
nor UO_293 (O_293,N_4943,N_4923);
or UO_294 (O_294,N_4932,N_4950);
nand UO_295 (O_295,N_4990,N_4979);
and UO_296 (O_296,N_4936,N_4917);
and UO_297 (O_297,N_4938,N_4960);
xor UO_298 (O_298,N_4961,N_4943);
or UO_299 (O_299,N_4904,N_4964);
and UO_300 (O_300,N_4967,N_4934);
nand UO_301 (O_301,N_4948,N_4978);
nand UO_302 (O_302,N_4988,N_4908);
xor UO_303 (O_303,N_4946,N_4901);
nand UO_304 (O_304,N_4905,N_4931);
nand UO_305 (O_305,N_4990,N_4945);
nand UO_306 (O_306,N_4917,N_4982);
or UO_307 (O_307,N_4994,N_4932);
nand UO_308 (O_308,N_4962,N_4983);
nor UO_309 (O_309,N_4907,N_4923);
or UO_310 (O_310,N_4953,N_4910);
and UO_311 (O_311,N_4964,N_4918);
nor UO_312 (O_312,N_4916,N_4902);
nor UO_313 (O_313,N_4988,N_4920);
nand UO_314 (O_314,N_4910,N_4907);
or UO_315 (O_315,N_4961,N_4903);
and UO_316 (O_316,N_4918,N_4911);
or UO_317 (O_317,N_4918,N_4932);
xnor UO_318 (O_318,N_4923,N_4927);
and UO_319 (O_319,N_4986,N_4950);
nand UO_320 (O_320,N_4913,N_4933);
xor UO_321 (O_321,N_4957,N_4930);
nand UO_322 (O_322,N_4927,N_4968);
nor UO_323 (O_323,N_4904,N_4953);
nor UO_324 (O_324,N_4989,N_4915);
nand UO_325 (O_325,N_4973,N_4981);
nor UO_326 (O_326,N_4961,N_4960);
xnor UO_327 (O_327,N_4979,N_4969);
nand UO_328 (O_328,N_4939,N_4908);
or UO_329 (O_329,N_4917,N_4925);
nor UO_330 (O_330,N_4953,N_4948);
xor UO_331 (O_331,N_4900,N_4982);
nor UO_332 (O_332,N_4907,N_4917);
or UO_333 (O_333,N_4981,N_4995);
and UO_334 (O_334,N_4977,N_4990);
or UO_335 (O_335,N_4987,N_4972);
nand UO_336 (O_336,N_4954,N_4962);
and UO_337 (O_337,N_4933,N_4940);
nand UO_338 (O_338,N_4917,N_4934);
or UO_339 (O_339,N_4994,N_4937);
or UO_340 (O_340,N_4967,N_4976);
nand UO_341 (O_341,N_4941,N_4927);
xor UO_342 (O_342,N_4920,N_4970);
nor UO_343 (O_343,N_4948,N_4904);
nor UO_344 (O_344,N_4983,N_4917);
and UO_345 (O_345,N_4994,N_4945);
or UO_346 (O_346,N_4927,N_4971);
nor UO_347 (O_347,N_4966,N_4930);
nor UO_348 (O_348,N_4920,N_4945);
xor UO_349 (O_349,N_4996,N_4937);
xnor UO_350 (O_350,N_4989,N_4966);
nand UO_351 (O_351,N_4931,N_4942);
xnor UO_352 (O_352,N_4990,N_4959);
or UO_353 (O_353,N_4996,N_4902);
nor UO_354 (O_354,N_4919,N_4925);
nor UO_355 (O_355,N_4987,N_4944);
xnor UO_356 (O_356,N_4980,N_4937);
nand UO_357 (O_357,N_4917,N_4966);
xor UO_358 (O_358,N_4902,N_4948);
nor UO_359 (O_359,N_4962,N_4938);
nand UO_360 (O_360,N_4903,N_4906);
or UO_361 (O_361,N_4974,N_4903);
nand UO_362 (O_362,N_4906,N_4938);
xor UO_363 (O_363,N_4906,N_4941);
xor UO_364 (O_364,N_4911,N_4980);
xor UO_365 (O_365,N_4910,N_4909);
xor UO_366 (O_366,N_4987,N_4945);
nand UO_367 (O_367,N_4961,N_4940);
nor UO_368 (O_368,N_4914,N_4996);
nor UO_369 (O_369,N_4926,N_4953);
nand UO_370 (O_370,N_4921,N_4952);
nand UO_371 (O_371,N_4970,N_4949);
or UO_372 (O_372,N_4905,N_4900);
and UO_373 (O_373,N_4968,N_4938);
xor UO_374 (O_374,N_4993,N_4947);
and UO_375 (O_375,N_4980,N_4931);
nor UO_376 (O_376,N_4992,N_4915);
nor UO_377 (O_377,N_4938,N_4932);
nand UO_378 (O_378,N_4901,N_4936);
xor UO_379 (O_379,N_4933,N_4906);
nor UO_380 (O_380,N_4962,N_4974);
and UO_381 (O_381,N_4994,N_4930);
or UO_382 (O_382,N_4936,N_4965);
nand UO_383 (O_383,N_4923,N_4986);
nand UO_384 (O_384,N_4957,N_4941);
nand UO_385 (O_385,N_4984,N_4919);
and UO_386 (O_386,N_4966,N_4942);
and UO_387 (O_387,N_4981,N_4943);
nor UO_388 (O_388,N_4989,N_4982);
and UO_389 (O_389,N_4923,N_4910);
nand UO_390 (O_390,N_4955,N_4904);
nor UO_391 (O_391,N_4928,N_4966);
xor UO_392 (O_392,N_4985,N_4947);
xor UO_393 (O_393,N_4970,N_4988);
nand UO_394 (O_394,N_4998,N_4909);
and UO_395 (O_395,N_4969,N_4902);
nor UO_396 (O_396,N_4912,N_4941);
or UO_397 (O_397,N_4914,N_4936);
nor UO_398 (O_398,N_4989,N_4903);
and UO_399 (O_399,N_4953,N_4905);
or UO_400 (O_400,N_4965,N_4954);
nor UO_401 (O_401,N_4982,N_4990);
and UO_402 (O_402,N_4975,N_4960);
and UO_403 (O_403,N_4995,N_4936);
and UO_404 (O_404,N_4909,N_4993);
xnor UO_405 (O_405,N_4958,N_4986);
nand UO_406 (O_406,N_4972,N_4904);
and UO_407 (O_407,N_4978,N_4985);
or UO_408 (O_408,N_4951,N_4935);
nand UO_409 (O_409,N_4926,N_4932);
or UO_410 (O_410,N_4996,N_4973);
nor UO_411 (O_411,N_4941,N_4949);
nor UO_412 (O_412,N_4928,N_4987);
xnor UO_413 (O_413,N_4934,N_4915);
xor UO_414 (O_414,N_4942,N_4992);
or UO_415 (O_415,N_4991,N_4943);
or UO_416 (O_416,N_4947,N_4988);
xnor UO_417 (O_417,N_4994,N_4922);
xnor UO_418 (O_418,N_4905,N_4915);
nor UO_419 (O_419,N_4902,N_4931);
xor UO_420 (O_420,N_4969,N_4993);
and UO_421 (O_421,N_4937,N_4933);
and UO_422 (O_422,N_4916,N_4964);
or UO_423 (O_423,N_4937,N_4934);
xnor UO_424 (O_424,N_4909,N_4967);
nand UO_425 (O_425,N_4944,N_4908);
and UO_426 (O_426,N_4983,N_4992);
or UO_427 (O_427,N_4970,N_4976);
and UO_428 (O_428,N_4912,N_4930);
xor UO_429 (O_429,N_4998,N_4922);
xor UO_430 (O_430,N_4956,N_4936);
and UO_431 (O_431,N_4954,N_4970);
or UO_432 (O_432,N_4951,N_4906);
nand UO_433 (O_433,N_4976,N_4940);
xnor UO_434 (O_434,N_4945,N_4917);
nand UO_435 (O_435,N_4936,N_4957);
nand UO_436 (O_436,N_4999,N_4927);
nand UO_437 (O_437,N_4924,N_4975);
nand UO_438 (O_438,N_4964,N_4976);
nand UO_439 (O_439,N_4988,N_4943);
xnor UO_440 (O_440,N_4998,N_4974);
or UO_441 (O_441,N_4949,N_4953);
nor UO_442 (O_442,N_4906,N_4991);
or UO_443 (O_443,N_4948,N_4930);
xnor UO_444 (O_444,N_4924,N_4927);
and UO_445 (O_445,N_4939,N_4952);
nor UO_446 (O_446,N_4970,N_4979);
nand UO_447 (O_447,N_4921,N_4957);
or UO_448 (O_448,N_4905,N_4960);
xor UO_449 (O_449,N_4984,N_4997);
and UO_450 (O_450,N_4966,N_4934);
xnor UO_451 (O_451,N_4962,N_4987);
or UO_452 (O_452,N_4934,N_4908);
or UO_453 (O_453,N_4973,N_4951);
nand UO_454 (O_454,N_4906,N_4942);
and UO_455 (O_455,N_4958,N_4914);
nand UO_456 (O_456,N_4958,N_4993);
nor UO_457 (O_457,N_4943,N_4932);
nor UO_458 (O_458,N_4920,N_4939);
nand UO_459 (O_459,N_4928,N_4948);
nor UO_460 (O_460,N_4959,N_4963);
or UO_461 (O_461,N_4945,N_4970);
or UO_462 (O_462,N_4940,N_4941);
or UO_463 (O_463,N_4932,N_4995);
xnor UO_464 (O_464,N_4975,N_4902);
nor UO_465 (O_465,N_4983,N_4956);
nand UO_466 (O_466,N_4906,N_4909);
xor UO_467 (O_467,N_4908,N_4941);
and UO_468 (O_468,N_4946,N_4918);
or UO_469 (O_469,N_4908,N_4935);
nor UO_470 (O_470,N_4944,N_4929);
nor UO_471 (O_471,N_4901,N_4903);
or UO_472 (O_472,N_4983,N_4976);
nand UO_473 (O_473,N_4912,N_4950);
xor UO_474 (O_474,N_4939,N_4921);
nand UO_475 (O_475,N_4985,N_4951);
and UO_476 (O_476,N_4920,N_4940);
and UO_477 (O_477,N_4916,N_4949);
or UO_478 (O_478,N_4972,N_4952);
and UO_479 (O_479,N_4957,N_4919);
nand UO_480 (O_480,N_4999,N_4938);
or UO_481 (O_481,N_4981,N_4961);
and UO_482 (O_482,N_4925,N_4910);
nand UO_483 (O_483,N_4993,N_4982);
and UO_484 (O_484,N_4904,N_4978);
and UO_485 (O_485,N_4960,N_4908);
nand UO_486 (O_486,N_4976,N_4980);
and UO_487 (O_487,N_4981,N_4988);
and UO_488 (O_488,N_4983,N_4921);
nor UO_489 (O_489,N_4941,N_4968);
xor UO_490 (O_490,N_4917,N_4960);
nor UO_491 (O_491,N_4965,N_4977);
nand UO_492 (O_492,N_4968,N_4950);
nor UO_493 (O_493,N_4903,N_4907);
xnor UO_494 (O_494,N_4915,N_4976);
or UO_495 (O_495,N_4986,N_4973);
nand UO_496 (O_496,N_4957,N_4985);
nand UO_497 (O_497,N_4999,N_4979);
nor UO_498 (O_498,N_4971,N_4998);
or UO_499 (O_499,N_4962,N_4992);
xnor UO_500 (O_500,N_4909,N_4972);
nor UO_501 (O_501,N_4910,N_4942);
or UO_502 (O_502,N_4942,N_4987);
nand UO_503 (O_503,N_4937,N_4947);
nand UO_504 (O_504,N_4967,N_4990);
nor UO_505 (O_505,N_4985,N_4901);
nor UO_506 (O_506,N_4958,N_4975);
and UO_507 (O_507,N_4976,N_4916);
and UO_508 (O_508,N_4974,N_4935);
xnor UO_509 (O_509,N_4978,N_4967);
nor UO_510 (O_510,N_4964,N_4934);
nand UO_511 (O_511,N_4939,N_4941);
nor UO_512 (O_512,N_4937,N_4929);
or UO_513 (O_513,N_4901,N_4959);
nor UO_514 (O_514,N_4951,N_4943);
and UO_515 (O_515,N_4902,N_4974);
or UO_516 (O_516,N_4970,N_4967);
nor UO_517 (O_517,N_4900,N_4965);
and UO_518 (O_518,N_4934,N_4960);
xnor UO_519 (O_519,N_4988,N_4966);
xnor UO_520 (O_520,N_4974,N_4980);
xnor UO_521 (O_521,N_4983,N_4967);
nor UO_522 (O_522,N_4925,N_4997);
nand UO_523 (O_523,N_4964,N_4984);
nand UO_524 (O_524,N_4968,N_4954);
or UO_525 (O_525,N_4999,N_4964);
nor UO_526 (O_526,N_4985,N_4973);
and UO_527 (O_527,N_4972,N_4924);
nand UO_528 (O_528,N_4973,N_4953);
and UO_529 (O_529,N_4974,N_4970);
xnor UO_530 (O_530,N_4903,N_4920);
xor UO_531 (O_531,N_4914,N_4930);
or UO_532 (O_532,N_4902,N_4999);
nor UO_533 (O_533,N_4926,N_4930);
nand UO_534 (O_534,N_4916,N_4954);
xnor UO_535 (O_535,N_4943,N_4939);
and UO_536 (O_536,N_4923,N_4997);
and UO_537 (O_537,N_4924,N_4907);
xnor UO_538 (O_538,N_4925,N_4930);
nor UO_539 (O_539,N_4905,N_4925);
xnor UO_540 (O_540,N_4961,N_4922);
nor UO_541 (O_541,N_4931,N_4960);
xnor UO_542 (O_542,N_4930,N_4917);
nor UO_543 (O_543,N_4931,N_4944);
and UO_544 (O_544,N_4972,N_4997);
or UO_545 (O_545,N_4940,N_4967);
xor UO_546 (O_546,N_4970,N_4948);
or UO_547 (O_547,N_4937,N_4905);
xor UO_548 (O_548,N_4909,N_4963);
or UO_549 (O_549,N_4980,N_4971);
xor UO_550 (O_550,N_4998,N_4962);
and UO_551 (O_551,N_4988,N_4990);
or UO_552 (O_552,N_4957,N_4927);
or UO_553 (O_553,N_4937,N_4960);
nand UO_554 (O_554,N_4942,N_4972);
and UO_555 (O_555,N_4991,N_4914);
nor UO_556 (O_556,N_4977,N_4975);
nor UO_557 (O_557,N_4965,N_4950);
xnor UO_558 (O_558,N_4961,N_4900);
and UO_559 (O_559,N_4915,N_4966);
xor UO_560 (O_560,N_4949,N_4969);
nand UO_561 (O_561,N_4904,N_4922);
nand UO_562 (O_562,N_4975,N_4990);
or UO_563 (O_563,N_4945,N_4926);
and UO_564 (O_564,N_4922,N_4979);
nand UO_565 (O_565,N_4918,N_4933);
nor UO_566 (O_566,N_4907,N_4937);
xnor UO_567 (O_567,N_4945,N_4948);
nor UO_568 (O_568,N_4958,N_4956);
xor UO_569 (O_569,N_4956,N_4907);
nor UO_570 (O_570,N_4932,N_4960);
and UO_571 (O_571,N_4961,N_4905);
nor UO_572 (O_572,N_4995,N_4950);
nand UO_573 (O_573,N_4991,N_4970);
and UO_574 (O_574,N_4987,N_4905);
or UO_575 (O_575,N_4963,N_4938);
nor UO_576 (O_576,N_4976,N_4920);
xor UO_577 (O_577,N_4946,N_4961);
xor UO_578 (O_578,N_4949,N_4903);
nand UO_579 (O_579,N_4917,N_4968);
and UO_580 (O_580,N_4989,N_4952);
xnor UO_581 (O_581,N_4931,N_4998);
nand UO_582 (O_582,N_4918,N_4939);
nor UO_583 (O_583,N_4983,N_4923);
nor UO_584 (O_584,N_4971,N_4957);
xor UO_585 (O_585,N_4995,N_4952);
xnor UO_586 (O_586,N_4964,N_4997);
nor UO_587 (O_587,N_4951,N_4944);
xor UO_588 (O_588,N_4935,N_4976);
xor UO_589 (O_589,N_4949,N_4954);
and UO_590 (O_590,N_4933,N_4921);
or UO_591 (O_591,N_4905,N_4982);
nand UO_592 (O_592,N_4925,N_4970);
or UO_593 (O_593,N_4986,N_4936);
and UO_594 (O_594,N_4925,N_4998);
and UO_595 (O_595,N_4930,N_4991);
nor UO_596 (O_596,N_4991,N_4955);
nand UO_597 (O_597,N_4985,N_4965);
nand UO_598 (O_598,N_4949,N_4984);
nor UO_599 (O_599,N_4962,N_4947);
or UO_600 (O_600,N_4924,N_4913);
or UO_601 (O_601,N_4936,N_4943);
xnor UO_602 (O_602,N_4923,N_4994);
and UO_603 (O_603,N_4922,N_4970);
xor UO_604 (O_604,N_4918,N_4934);
xor UO_605 (O_605,N_4916,N_4908);
or UO_606 (O_606,N_4993,N_4976);
or UO_607 (O_607,N_4957,N_4960);
and UO_608 (O_608,N_4961,N_4950);
and UO_609 (O_609,N_4975,N_4928);
nand UO_610 (O_610,N_4901,N_4935);
nand UO_611 (O_611,N_4923,N_4956);
or UO_612 (O_612,N_4926,N_4921);
and UO_613 (O_613,N_4963,N_4900);
nor UO_614 (O_614,N_4980,N_4909);
and UO_615 (O_615,N_4928,N_4958);
and UO_616 (O_616,N_4954,N_4996);
xnor UO_617 (O_617,N_4968,N_4997);
or UO_618 (O_618,N_4962,N_4921);
and UO_619 (O_619,N_4906,N_4973);
nor UO_620 (O_620,N_4923,N_4919);
nor UO_621 (O_621,N_4953,N_4965);
or UO_622 (O_622,N_4954,N_4900);
and UO_623 (O_623,N_4963,N_4946);
xnor UO_624 (O_624,N_4997,N_4905);
or UO_625 (O_625,N_4923,N_4941);
nand UO_626 (O_626,N_4953,N_4985);
nand UO_627 (O_627,N_4970,N_4907);
xor UO_628 (O_628,N_4970,N_4999);
or UO_629 (O_629,N_4958,N_4980);
nor UO_630 (O_630,N_4932,N_4983);
or UO_631 (O_631,N_4943,N_4933);
nand UO_632 (O_632,N_4994,N_4987);
nor UO_633 (O_633,N_4990,N_4914);
xor UO_634 (O_634,N_4987,N_4900);
nand UO_635 (O_635,N_4909,N_4912);
and UO_636 (O_636,N_4971,N_4959);
nand UO_637 (O_637,N_4944,N_4911);
or UO_638 (O_638,N_4935,N_4927);
nor UO_639 (O_639,N_4911,N_4958);
nand UO_640 (O_640,N_4946,N_4984);
nor UO_641 (O_641,N_4994,N_4929);
or UO_642 (O_642,N_4997,N_4992);
xor UO_643 (O_643,N_4909,N_4982);
nand UO_644 (O_644,N_4998,N_4958);
nand UO_645 (O_645,N_4979,N_4924);
or UO_646 (O_646,N_4947,N_4969);
xor UO_647 (O_647,N_4952,N_4974);
and UO_648 (O_648,N_4990,N_4931);
nand UO_649 (O_649,N_4950,N_4955);
xnor UO_650 (O_650,N_4943,N_4983);
nand UO_651 (O_651,N_4979,N_4980);
nor UO_652 (O_652,N_4999,N_4982);
xor UO_653 (O_653,N_4936,N_4988);
nand UO_654 (O_654,N_4969,N_4974);
xor UO_655 (O_655,N_4951,N_4969);
and UO_656 (O_656,N_4950,N_4947);
or UO_657 (O_657,N_4982,N_4926);
xnor UO_658 (O_658,N_4953,N_4977);
nand UO_659 (O_659,N_4963,N_4989);
nor UO_660 (O_660,N_4969,N_4997);
nand UO_661 (O_661,N_4991,N_4904);
nor UO_662 (O_662,N_4979,N_4918);
or UO_663 (O_663,N_4966,N_4959);
nand UO_664 (O_664,N_4943,N_4909);
nand UO_665 (O_665,N_4918,N_4986);
nor UO_666 (O_666,N_4996,N_4977);
and UO_667 (O_667,N_4978,N_4986);
xor UO_668 (O_668,N_4978,N_4927);
or UO_669 (O_669,N_4985,N_4912);
nor UO_670 (O_670,N_4977,N_4952);
xnor UO_671 (O_671,N_4941,N_4996);
nand UO_672 (O_672,N_4906,N_4910);
xor UO_673 (O_673,N_4978,N_4917);
and UO_674 (O_674,N_4957,N_4909);
nor UO_675 (O_675,N_4977,N_4927);
nand UO_676 (O_676,N_4944,N_4957);
and UO_677 (O_677,N_4981,N_4917);
nand UO_678 (O_678,N_4913,N_4990);
or UO_679 (O_679,N_4986,N_4934);
nand UO_680 (O_680,N_4978,N_4964);
nand UO_681 (O_681,N_4936,N_4908);
or UO_682 (O_682,N_4976,N_4901);
nor UO_683 (O_683,N_4994,N_4995);
or UO_684 (O_684,N_4909,N_4978);
nor UO_685 (O_685,N_4965,N_4906);
and UO_686 (O_686,N_4943,N_4906);
nor UO_687 (O_687,N_4993,N_4926);
nand UO_688 (O_688,N_4946,N_4927);
nand UO_689 (O_689,N_4964,N_4941);
nand UO_690 (O_690,N_4947,N_4957);
nand UO_691 (O_691,N_4958,N_4907);
xor UO_692 (O_692,N_4915,N_4980);
and UO_693 (O_693,N_4928,N_4907);
xnor UO_694 (O_694,N_4928,N_4910);
nand UO_695 (O_695,N_4934,N_4974);
nor UO_696 (O_696,N_4972,N_4945);
nand UO_697 (O_697,N_4960,N_4955);
or UO_698 (O_698,N_4925,N_4978);
xnor UO_699 (O_699,N_4903,N_4939);
or UO_700 (O_700,N_4969,N_4959);
xor UO_701 (O_701,N_4913,N_4966);
nor UO_702 (O_702,N_4982,N_4937);
and UO_703 (O_703,N_4931,N_4988);
nand UO_704 (O_704,N_4924,N_4912);
nor UO_705 (O_705,N_4918,N_4973);
or UO_706 (O_706,N_4943,N_4989);
or UO_707 (O_707,N_4916,N_4933);
nor UO_708 (O_708,N_4993,N_4930);
and UO_709 (O_709,N_4928,N_4923);
nand UO_710 (O_710,N_4982,N_4922);
nand UO_711 (O_711,N_4911,N_4925);
xnor UO_712 (O_712,N_4921,N_4947);
or UO_713 (O_713,N_4940,N_4926);
nor UO_714 (O_714,N_4959,N_4958);
or UO_715 (O_715,N_4994,N_4913);
xnor UO_716 (O_716,N_4940,N_4989);
and UO_717 (O_717,N_4926,N_4928);
xnor UO_718 (O_718,N_4972,N_4992);
nand UO_719 (O_719,N_4959,N_4992);
and UO_720 (O_720,N_4983,N_4946);
and UO_721 (O_721,N_4976,N_4990);
xnor UO_722 (O_722,N_4972,N_4923);
nor UO_723 (O_723,N_4951,N_4968);
nand UO_724 (O_724,N_4940,N_4925);
nand UO_725 (O_725,N_4921,N_4950);
and UO_726 (O_726,N_4941,N_4916);
and UO_727 (O_727,N_4948,N_4958);
xor UO_728 (O_728,N_4928,N_4967);
xnor UO_729 (O_729,N_4977,N_4948);
or UO_730 (O_730,N_4970,N_4923);
or UO_731 (O_731,N_4919,N_4929);
or UO_732 (O_732,N_4953,N_4992);
and UO_733 (O_733,N_4951,N_4975);
or UO_734 (O_734,N_4967,N_4921);
and UO_735 (O_735,N_4919,N_4938);
and UO_736 (O_736,N_4907,N_4980);
nor UO_737 (O_737,N_4989,N_4986);
xnor UO_738 (O_738,N_4983,N_4986);
nand UO_739 (O_739,N_4927,N_4906);
or UO_740 (O_740,N_4928,N_4935);
or UO_741 (O_741,N_4907,N_4902);
nor UO_742 (O_742,N_4953,N_4966);
nand UO_743 (O_743,N_4994,N_4925);
or UO_744 (O_744,N_4963,N_4923);
or UO_745 (O_745,N_4995,N_4992);
xnor UO_746 (O_746,N_4955,N_4924);
or UO_747 (O_747,N_4906,N_4918);
nor UO_748 (O_748,N_4999,N_4951);
nand UO_749 (O_749,N_4930,N_4913);
xor UO_750 (O_750,N_4955,N_4999);
or UO_751 (O_751,N_4937,N_4943);
xor UO_752 (O_752,N_4917,N_4937);
nor UO_753 (O_753,N_4955,N_4951);
nand UO_754 (O_754,N_4951,N_4939);
nor UO_755 (O_755,N_4969,N_4920);
and UO_756 (O_756,N_4958,N_4932);
or UO_757 (O_757,N_4941,N_4954);
nor UO_758 (O_758,N_4928,N_4997);
nor UO_759 (O_759,N_4976,N_4985);
and UO_760 (O_760,N_4990,N_4987);
nor UO_761 (O_761,N_4902,N_4960);
nand UO_762 (O_762,N_4905,N_4919);
nor UO_763 (O_763,N_4958,N_4963);
and UO_764 (O_764,N_4928,N_4981);
or UO_765 (O_765,N_4906,N_4996);
nand UO_766 (O_766,N_4923,N_4902);
xnor UO_767 (O_767,N_4957,N_4912);
nand UO_768 (O_768,N_4919,N_4961);
xor UO_769 (O_769,N_4907,N_4967);
nand UO_770 (O_770,N_4989,N_4981);
xor UO_771 (O_771,N_4917,N_4993);
nor UO_772 (O_772,N_4971,N_4905);
nor UO_773 (O_773,N_4987,N_4916);
or UO_774 (O_774,N_4947,N_4998);
nor UO_775 (O_775,N_4904,N_4936);
and UO_776 (O_776,N_4960,N_4947);
xor UO_777 (O_777,N_4984,N_4929);
nand UO_778 (O_778,N_4936,N_4933);
nand UO_779 (O_779,N_4943,N_4978);
and UO_780 (O_780,N_4979,N_4952);
nor UO_781 (O_781,N_4969,N_4992);
and UO_782 (O_782,N_4914,N_4906);
xor UO_783 (O_783,N_4908,N_4930);
or UO_784 (O_784,N_4935,N_4906);
nand UO_785 (O_785,N_4988,N_4914);
or UO_786 (O_786,N_4937,N_4916);
xnor UO_787 (O_787,N_4913,N_4964);
or UO_788 (O_788,N_4974,N_4932);
nor UO_789 (O_789,N_4952,N_4912);
or UO_790 (O_790,N_4925,N_4992);
or UO_791 (O_791,N_4921,N_4959);
nand UO_792 (O_792,N_4913,N_4979);
or UO_793 (O_793,N_4933,N_4980);
or UO_794 (O_794,N_4979,N_4923);
nor UO_795 (O_795,N_4926,N_4964);
and UO_796 (O_796,N_4983,N_4966);
xnor UO_797 (O_797,N_4929,N_4975);
or UO_798 (O_798,N_4944,N_4991);
or UO_799 (O_799,N_4905,N_4993);
xor UO_800 (O_800,N_4964,N_4908);
nand UO_801 (O_801,N_4978,N_4942);
or UO_802 (O_802,N_4995,N_4977);
nand UO_803 (O_803,N_4929,N_4926);
nor UO_804 (O_804,N_4995,N_4985);
nand UO_805 (O_805,N_4990,N_4992);
and UO_806 (O_806,N_4985,N_4918);
or UO_807 (O_807,N_4973,N_4975);
xor UO_808 (O_808,N_4972,N_4912);
xnor UO_809 (O_809,N_4925,N_4967);
or UO_810 (O_810,N_4900,N_4922);
nand UO_811 (O_811,N_4960,N_4956);
and UO_812 (O_812,N_4982,N_4980);
and UO_813 (O_813,N_4985,N_4940);
nand UO_814 (O_814,N_4933,N_4997);
nor UO_815 (O_815,N_4972,N_4918);
nand UO_816 (O_816,N_4911,N_4986);
nor UO_817 (O_817,N_4968,N_4913);
and UO_818 (O_818,N_4949,N_4976);
xor UO_819 (O_819,N_4947,N_4931);
and UO_820 (O_820,N_4921,N_4905);
or UO_821 (O_821,N_4945,N_4991);
xnor UO_822 (O_822,N_4910,N_4956);
nand UO_823 (O_823,N_4952,N_4996);
and UO_824 (O_824,N_4955,N_4996);
xor UO_825 (O_825,N_4939,N_4931);
and UO_826 (O_826,N_4994,N_4942);
nor UO_827 (O_827,N_4954,N_4903);
or UO_828 (O_828,N_4917,N_4903);
xnor UO_829 (O_829,N_4995,N_4915);
and UO_830 (O_830,N_4925,N_4964);
or UO_831 (O_831,N_4965,N_4944);
nand UO_832 (O_832,N_4904,N_4949);
or UO_833 (O_833,N_4970,N_4931);
xor UO_834 (O_834,N_4941,N_4973);
nor UO_835 (O_835,N_4998,N_4993);
xnor UO_836 (O_836,N_4923,N_4908);
or UO_837 (O_837,N_4969,N_4966);
nor UO_838 (O_838,N_4993,N_4978);
or UO_839 (O_839,N_4920,N_4953);
nor UO_840 (O_840,N_4979,N_4903);
xor UO_841 (O_841,N_4969,N_4926);
nand UO_842 (O_842,N_4979,N_4929);
nor UO_843 (O_843,N_4993,N_4929);
xnor UO_844 (O_844,N_4998,N_4986);
nor UO_845 (O_845,N_4959,N_4947);
nor UO_846 (O_846,N_4942,N_4975);
nand UO_847 (O_847,N_4976,N_4962);
xor UO_848 (O_848,N_4955,N_4940);
and UO_849 (O_849,N_4965,N_4973);
or UO_850 (O_850,N_4917,N_4954);
or UO_851 (O_851,N_4943,N_4949);
nor UO_852 (O_852,N_4957,N_4974);
nand UO_853 (O_853,N_4946,N_4980);
nor UO_854 (O_854,N_4978,N_4949);
nor UO_855 (O_855,N_4910,N_4949);
and UO_856 (O_856,N_4953,N_4997);
or UO_857 (O_857,N_4906,N_4940);
or UO_858 (O_858,N_4918,N_4950);
and UO_859 (O_859,N_4923,N_4940);
and UO_860 (O_860,N_4969,N_4954);
nor UO_861 (O_861,N_4964,N_4922);
and UO_862 (O_862,N_4981,N_4966);
and UO_863 (O_863,N_4959,N_4941);
nand UO_864 (O_864,N_4919,N_4913);
xnor UO_865 (O_865,N_4916,N_4903);
and UO_866 (O_866,N_4994,N_4980);
or UO_867 (O_867,N_4930,N_4974);
xor UO_868 (O_868,N_4932,N_4981);
xor UO_869 (O_869,N_4904,N_4999);
nor UO_870 (O_870,N_4961,N_4929);
or UO_871 (O_871,N_4979,N_4972);
nor UO_872 (O_872,N_4913,N_4915);
nor UO_873 (O_873,N_4922,N_4966);
nor UO_874 (O_874,N_4969,N_4935);
nor UO_875 (O_875,N_4926,N_4948);
and UO_876 (O_876,N_4972,N_4938);
nor UO_877 (O_877,N_4929,N_4969);
nor UO_878 (O_878,N_4988,N_4923);
nor UO_879 (O_879,N_4928,N_4938);
nor UO_880 (O_880,N_4922,N_4926);
nand UO_881 (O_881,N_4914,N_4924);
or UO_882 (O_882,N_4963,N_4976);
or UO_883 (O_883,N_4950,N_4985);
xnor UO_884 (O_884,N_4990,N_4951);
nand UO_885 (O_885,N_4939,N_4972);
nor UO_886 (O_886,N_4913,N_4922);
nor UO_887 (O_887,N_4975,N_4971);
or UO_888 (O_888,N_4984,N_4990);
or UO_889 (O_889,N_4986,N_4915);
nand UO_890 (O_890,N_4951,N_4950);
nor UO_891 (O_891,N_4968,N_4934);
nor UO_892 (O_892,N_4940,N_4935);
xor UO_893 (O_893,N_4919,N_4934);
nand UO_894 (O_894,N_4953,N_4962);
or UO_895 (O_895,N_4946,N_4976);
and UO_896 (O_896,N_4915,N_4902);
nor UO_897 (O_897,N_4962,N_4933);
nand UO_898 (O_898,N_4923,N_4984);
or UO_899 (O_899,N_4982,N_4985);
nand UO_900 (O_900,N_4998,N_4917);
and UO_901 (O_901,N_4960,N_4974);
nor UO_902 (O_902,N_4933,N_4926);
or UO_903 (O_903,N_4928,N_4982);
nand UO_904 (O_904,N_4983,N_4949);
nand UO_905 (O_905,N_4934,N_4996);
xor UO_906 (O_906,N_4929,N_4918);
nor UO_907 (O_907,N_4971,N_4933);
and UO_908 (O_908,N_4941,N_4976);
nand UO_909 (O_909,N_4958,N_4981);
and UO_910 (O_910,N_4970,N_4942);
xnor UO_911 (O_911,N_4919,N_4979);
nor UO_912 (O_912,N_4937,N_4915);
nand UO_913 (O_913,N_4929,N_4985);
and UO_914 (O_914,N_4950,N_4917);
and UO_915 (O_915,N_4972,N_4947);
nand UO_916 (O_916,N_4969,N_4978);
nor UO_917 (O_917,N_4969,N_4938);
xnor UO_918 (O_918,N_4943,N_4987);
and UO_919 (O_919,N_4930,N_4960);
and UO_920 (O_920,N_4900,N_4966);
xor UO_921 (O_921,N_4919,N_4968);
nor UO_922 (O_922,N_4908,N_4951);
and UO_923 (O_923,N_4980,N_4925);
and UO_924 (O_924,N_4992,N_4923);
or UO_925 (O_925,N_4934,N_4942);
nand UO_926 (O_926,N_4900,N_4938);
nor UO_927 (O_927,N_4986,N_4942);
or UO_928 (O_928,N_4909,N_4968);
xnor UO_929 (O_929,N_4934,N_4972);
nor UO_930 (O_930,N_4933,N_4973);
nor UO_931 (O_931,N_4943,N_4938);
nor UO_932 (O_932,N_4906,N_4969);
nor UO_933 (O_933,N_4942,N_4949);
and UO_934 (O_934,N_4944,N_4935);
nor UO_935 (O_935,N_4912,N_4960);
and UO_936 (O_936,N_4933,N_4963);
nand UO_937 (O_937,N_4937,N_4965);
xnor UO_938 (O_938,N_4905,N_4904);
or UO_939 (O_939,N_4919,N_4927);
and UO_940 (O_940,N_4945,N_4927);
nor UO_941 (O_941,N_4941,N_4971);
xor UO_942 (O_942,N_4949,N_4911);
xor UO_943 (O_943,N_4996,N_4924);
nand UO_944 (O_944,N_4987,N_4955);
nor UO_945 (O_945,N_4926,N_4904);
nand UO_946 (O_946,N_4974,N_4956);
nand UO_947 (O_947,N_4914,N_4976);
and UO_948 (O_948,N_4957,N_4955);
and UO_949 (O_949,N_4996,N_4918);
nor UO_950 (O_950,N_4936,N_4970);
or UO_951 (O_951,N_4962,N_4934);
or UO_952 (O_952,N_4923,N_4944);
xor UO_953 (O_953,N_4970,N_4947);
nand UO_954 (O_954,N_4918,N_4952);
or UO_955 (O_955,N_4908,N_4980);
and UO_956 (O_956,N_4980,N_4944);
nor UO_957 (O_957,N_4985,N_4927);
or UO_958 (O_958,N_4952,N_4915);
or UO_959 (O_959,N_4916,N_4968);
or UO_960 (O_960,N_4960,N_4989);
nor UO_961 (O_961,N_4932,N_4931);
xnor UO_962 (O_962,N_4914,N_4950);
xor UO_963 (O_963,N_4985,N_4983);
xor UO_964 (O_964,N_4911,N_4948);
xor UO_965 (O_965,N_4903,N_4991);
or UO_966 (O_966,N_4910,N_4990);
nor UO_967 (O_967,N_4991,N_4960);
xnor UO_968 (O_968,N_4901,N_4988);
nand UO_969 (O_969,N_4996,N_4923);
xnor UO_970 (O_970,N_4968,N_4948);
xnor UO_971 (O_971,N_4947,N_4956);
nor UO_972 (O_972,N_4957,N_4961);
xor UO_973 (O_973,N_4960,N_4972);
and UO_974 (O_974,N_4904,N_4984);
or UO_975 (O_975,N_4956,N_4950);
nand UO_976 (O_976,N_4950,N_4940);
nor UO_977 (O_977,N_4969,N_4958);
nand UO_978 (O_978,N_4954,N_4931);
nand UO_979 (O_979,N_4930,N_4941);
nor UO_980 (O_980,N_4919,N_4910);
xor UO_981 (O_981,N_4968,N_4980);
nor UO_982 (O_982,N_4930,N_4987);
and UO_983 (O_983,N_4926,N_4949);
nor UO_984 (O_984,N_4955,N_4930);
nor UO_985 (O_985,N_4992,N_4936);
or UO_986 (O_986,N_4945,N_4903);
or UO_987 (O_987,N_4914,N_4977);
and UO_988 (O_988,N_4981,N_4993);
and UO_989 (O_989,N_4927,N_4947);
or UO_990 (O_990,N_4995,N_4923);
or UO_991 (O_991,N_4992,N_4987);
nor UO_992 (O_992,N_4972,N_4968);
xor UO_993 (O_993,N_4991,N_4931);
nand UO_994 (O_994,N_4956,N_4948);
nand UO_995 (O_995,N_4938,N_4996);
or UO_996 (O_996,N_4984,N_4939);
or UO_997 (O_997,N_4954,N_4927);
xnor UO_998 (O_998,N_4939,N_4937);
or UO_999 (O_999,N_4966,N_4975);
endmodule